// Benchmark "dalu" written by ABC on Sun Apr 22 21:43:02 2018

module dalu ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461;
  assign n92 = ~pi66 & ~pi67;
  assign n93 = pi33 & pi70;
  assign n94 = ~pi70 & pi71;
  assign n95 = pi01 & n94;
  assign n96 = ~pi71 & n93;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~pi69 & ~n97;
  assign n99 = pi68 & n98;
  assign n100 = pi32 & pi70;
  assign n101 = pi00 & n94;
  assign n102 = ~pi71 & n100;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~pi69 & ~n103;
  assign n105 = pi68 & n104;
  assign n106 = ~n99 & n105;
  assign n107 = n99 & ~n105;
  assign n108 = ~n106 & ~n107;
  assign n109 = pi34 & pi70;
  assign n110 = pi02 & n94;
  assign n111 = ~pi71 & n109;
  assign n112 = ~n110 & ~n111;
  assign n113 = ~pi69 & ~n112;
  assign n114 = pi68 & n113;
  assign n115 = n105 & ~n114;
  assign n116 = ~n105 & n114;
  assign n117 = ~n115 & ~n116;
  assign n118 = pi35 & pi70;
  assign n119 = pi03 & n94;
  assign n120 = ~pi71 & n118;
  assign n121 = ~n119 & ~n120;
  assign n122 = ~pi69 & ~n121;
  assign n123 = pi68 & n122;
  assign n124 = n105 & ~n123;
  assign n125 = ~n105 & n123;
  assign n126 = ~n124 & ~n125;
  assign n127 = pi40 & pi70;
  assign n128 = pi08 & n94;
  assign n129 = ~pi71 & n127;
  assign n130 = ~n128 & ~n129;
  assign n131 = ~pi69 & ~n130;
  assign n132 = pi68 & n131;
  assign n133 = n105 & ~n132;
  assign n134 = ~n105 & n132;
  assign n135 = ~n133 & ~n134;
  assign n136 = pi41 & pi70;
  assign n137 = pi09 & n94;
  assign n138 = ~pi71 & n136;
  assign n139 = ~n137 & ~n138;
  assign n140 = ~pi69 & ~n139;
  assign n141 = pi68 & n140;
  assign n142 = n105 & ~n141;
  assign n143 = ~n105 & n141;
  assign n144 = ~n142 & ~n143;
  assign n145 = pi42 & pi70;
  assign n146 = pi10 & n94;
  assign n147 = ~pi71 & n145;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~pi69 & ~n148;
  assign n150 = pi68 & n149;
  assign n151 = n105 & ~n150;
  assign n152 = ~n105 & n150;
  assign n153 = ~n151 & ~n152;
  assign n154 = pi43 & pi70;
  assign n155 = pi11 & n94;
  assign n156 = ~pi71 & n154;
  assign n157 = ~n155 & ~n156;
  assign n158 = ~pi69 & ~n157;
  assign n159 = pi68 & n158;
  assign n160 = n105 & ~n159;
  assign n161 = ~n105 & n159;
  assign n162 = ~n160 & ~n161;
  assign n163 = ~n135 & ~n144;
  assign n164 = ~n153 & ~n162;
  assign n165 = n163 & n164;
  assign n166 = pi36 & pi70;
  assign n167 = pi04 & n94;
  assign n168 = ~pi71 & n166;
  assign n169 = ~n167 & ~n168;
  assign n170 = ~pi69 & ~n169;
  assign n171 = pi68 & n170;
  assign n172 = n105 & ~n171;
  assign n173 = ~n105 & n171;
  assign n174 = ~n172 & ~n173;
  assign n175 = pi37 & pi70;
  assign n176 = pi05 & n94;
  assign n177 = ~pi71 & n175;
  assign n178 = ~n176 & ~n177;
  assign n179 = ~pi69 & ~n178;
  assign n180 = pi68 & n179;
  assign n181 = n105 & ~n180;
  assign n182 = ~n105 & n180;
  assign n183 = ~n181 & ~n182;
  assign n184 = pi38 & pi70;
  assign n185 = pi06 & n94;
  assign n186 = ~pi71 & n184;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~pi69 & ~n187;
  assign n189 = pi68 & n188;
  assign n190 = n105 & ~n189;
  assign n191 = ~n105 & n189;
  assign n192 = ~n190 & ~n191;
  assign n193 = pi39 & pi70;
  assign n194 = pi07 & n94;
  assign n195 = ~pi71 & n193;
  assign n196 = ~n194 & ~n195;
  assign n197 = ~pi69 & ~n196;
  assign n198 = pi68 & n197;
  assign n199 = n105 & ~n198;
  assign n200 = ~n105 & n198;
  assign n201 = ~n199 & ~n200;
  assign n202 = ~n174 & ~n183;
  assign n203 = ~n192 & ~n201;
  assign n204 = n202 & n203;
  assign n205 = pi44 & pi70;
  assign n206 = pi12 & n94;
  assign n207 = ~pi71 & n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~pi69 & ~n208;
  assign n210 = pi68 & n209;
  assign n211 = n105 & ~n210;
  assign n212 = ~n105 & n210;
  assign n213 = ~n211 & ~n212;
  assign n214 = pi45 & pi70;
  assign n215 = pi13 & n94;
  assign n216 = ~pi71 & n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = ~pi69 & ~n217;
  assign n219 = pi68 & n218;
  assign n220 = n105 & ~n219;
  assign n221 = ~n105 & n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = pi46 & pi70;
  assign n224 = pi14 & n94;
  assign n225 = ~pi71 & n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~pi69 & ~n226;
  assign n228 = pi68 & n227;
  assign n229 = n105 & ~n228;
  assign n230 = ~n105 & n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = pi47 & pi70;
  assign n233 = pi15 & n94;
  assign n234 = ~pi71 & n232;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~pi69 & ~n235;
  assign n237 = pi68 & n236;
  assign n238 = n105 & ~n237;
  assign n239 = ~n105 & n237;
  assign n240 = ~n238 & ~n239;
  assign n241 = ~n213 & ~n222;
  assign n242 = ~n231 & ~n240;
  assign n243 = n241 & n242;
  assign n244 = n165 & n204;
  assign n245 = n105 & n244;
  assign n246 = n243 & n245;
  assign n247 = ~n108 & ~n117;
  assign n248 = ~n126 & n246;
  assign n249 = n247 & n248;
  assign n250 = pi48 & pi70;
  assign n251 = pi70 & ~pi71;
  assign n252 = ~n94 & ~n251;
  assign n253 = pi71 & n250;
  assign n254 = pi16 & ~n252;
  assign n255 = ~n253 & ~n254;
  assign n256 = ~pi68 & pi69;
  assign n257 = ~pi70 & ~pi71;
  assign n258 = ~pi69 & n257;
  assign n259 = pi48 & pi68;
  assign n260 = n258 & n259;
  assign n261 = ~n255 & n256;
  assign n262 = ~n260 & ~n261;
  assign n263 = pi65 & ~n262;
  assign n264 = ~pi65 & n249;
  assign n265 = ~n263 & ~n264;
  assign n266 = pi65 & n92;
  assign n267 = n249 & n266;
  assign n268 = ~n92 & ~n265;
  assign n269 = ~n267 & ~n268;
  assign n270 = pi00 & ~pi70;
  assign n271 = ~n100 & ~n270;
  assign n272 = ~pi69 & ~n271;
  assign n273 = pi71 & n272;
  assign n274 = pi69 & ~pi70;
  assign n275 = pi48 & n274;
  assign n276 = ~pi69 & pi70;
  assign n277 = pi16 & n276;
  assign n278 = ~n275 & ~n277;
  assign n279 = ~pi71 & ~n278;
  assign n280 = ~n273 & ~n279;
  assign n281 = ~pi68 & ~n280;
  assign n282 = pi32 & pi68;
  assign n283 = ~pi69 & n282;
  assign n284 = ~pi70 & n283;
  assign n285 = ~pi71 & n284;
  assign n286 = pi71 & n100;
  assign n287 = pi00 & ~n252;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~pi68 & ~n288;
  assign n290 = pi69 & n289;
  assign n291 = ~n285 & ~n290;
  assign n292 = ~pi64 & ~pi66;
  assign n293 = ~pi65 & pi66;
  assign n294 = ~n292 & ~n293;
  assign n295 = pi64 & pi65;
  assign n296 = ~pi67 & n294;
  assign n297 = ~n295 & n296;
  assign n298 = n291 & n297;
  assign n299 = ~n291 & ~n297;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~n281 & ~n300;
  assign n302 = n281 & n300;
  assign n303 = ~n301 & ~n302;
  assign n304 = pi33 & pi68;
  assign n305 = ~pi69 & n304;
  assign n306 = ~pi70 & n305;
  assign n307 = ~pi71 & n306;
  assign n308 = pi71 & n93;
  assign n309 = pi01 & ~n252;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~pi68 & ~n310;
  assign n312 = pi69 & n311;
  assign n313 = ~n307 & ~n312;
  assign n314 = n297 & n313;
  assign n315 = ~n297 & ~n313;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi01 & ~pi70;
  assign n318 = ~n93 & ~n317;
  assign n319 = ~pi69 & ~n318;
  assign n320 = pi71 & n319;
  assign n321 = pi49 & n274;
  assign n322 = pi17 & n276;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~pi71 & ~n323;
  assign n325 = ~n320 & ~n324;
  assign n326 = ~pi68 & ~n325;
  assign n327 = ~n316 & n326;
  assign n328 = pi34 & pi68;
  assign n329 = ~pi69 & n328;
  assign n330 = ~pi70 & n329;
  assign n331 = ~pi71 & n330;
  assign n332 = pi71 & n109;
  assign n333 = pi02 & ~n252;
  assign n334 = ~n332 & ~n333;
  assign n335 = ~pi68 & ~n334;
  assign n336 = pi69 & n335;
  assign n337 = ~n331 & ~n336;
  assign n338 = n297 & n337;
  assign n339 = ~n297 & ~n337;
  assign n340 = ~n338 & ~n339;
  assign n341 = pi02 & ~pi70;
  assign n342 = ~n109 & ~n341;
  assign n343 = ~pi69 & ~n342;
  assign n344 = pi71 & n343;
  assign n345 = pi50 & n274;
  assign n346 = pi18 & n276;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~pi71 & ~n347;
  assign n349 = ~n344 & ~n348;
  assign n350 = ~pi68 & ~n349;
  assign n351 = ~n340 & n350;
  assign n352 = pi35 & pi68;
  assign n353 = ~pi69 & n352;
  assign n354 = ~pi70 & n353;
  assign n355 = ~pi71 & n354;
  assign n356 = pi71 & n118;
  assign n357 = pi03 & ~n252;
  assign n358 = ~n356 & ~n357;
  assign n359 = ~pi68 & ~n358;
  assign n360 = pi69 & n359;
  assign n361 = ~n355 & ~n360;
  assign n362 = n297 & n361;
  assign n363 = ~n297 & ~n361;
  assign n364 = ~n362 & ~n363;
  assign n365 = pi03 & ~pi70;
  assign n366 = ~n118 & ~n365;
  assign n367 = ~pi69 & ~n366;
  assign n368 = pi71 & n367;
  assign n369 = pi51 & n274;
  assign n370 = pi19 & n276;
  assign n371 = ~n369 & ~n370;
  assign n372 = ~pi71 & ~n371;
  assign n373 = ~n368 & ~n372;
  assign n374 = ~pi68 & ~n373;
  assign n375 = ~n364 & n374;
  assign n376 = ~pi65 & ~pi66;
  assign n377 = pi64 & n376;
  assign n378 = ~pi64 & pi66;
  assign n379 = pi65 & n378;
  assign n380 = ~n377 & ~n379;
  assign n381 = ~pi67 & ~n380;
  assign n382 = pi12 & ~pi70;
  assign n383 = ~n205 & ~n382;
  assign n384 = ~pi69 & ~n383;
  assign n385 = pi71 & n384;
  assign n386 = pi60 & n274;
  assign n387 = pi28 & n276;
  assign n388 = ~n386 & ~n387;
  assign n389 = ~pi71 & ~n388;
  assign n390 = ~n385 & ~n389;
  assign n391 = ~pi68 & ~n390;
  assign n392 = pi44 & pi68;
  assign n393 = ~pi69 & n392;
  assign n394 = ~pi70 & n393;
  assign n395 = ~pi71 & n394;
  assign n396 = pi71 & n205;
  assign n397 = pi12 & ~n252;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~pi68 & ~n398;
  assign n400 = pi69 & n399;
  assign n401 = ~n395 & ~n400;
  assign n402 = n297 & n401;
  assign n403 = ~n297 & ~n401;
  assign n404 = ~n402 & ~n403;
  assign n405 = pi13 & ~pi70;
  assign n406 = ~n214 & ~n405;
  assign n407 = ~pi69 & ~n406;
  assign n408 = pi71 & n407;
  assign n409 = pi61 & n274;
  assign n410 = pi29 & n276;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~pi71 & ~n411;
  assign n413 = ~n408 & ~n412;
  assign n414 = ~pi68 & ~n413;
  assign n415 = pi45 & pi68;
  assign n416 = ~pi69 & n415;
  assign n417 = ~pi70 & n416;
  assign n418 = ~pi71 & n417;
  assign n419 = pi71 & n214;
  assign n420 = pi13 & ~n252;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~pi68 & ~n421;
  assign n423 = pi69 & n422;
  assign n424 = ~n418 & ~n423;
  assign n425 = n297 & n424;
  assign n426 = ~n297 & ~n424;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~n391 & n404;
  assign n429 = ~n414 & n427;
  assign n430 = ~n428 & ~n429;
  assign n431 = pi14 & ~pi70;
  assign n432 = ~n223 & ~n431;
  assign n433 = ~pi69 & ~n432;
  assign n434 = pi71 & n433;
  assign n435 = pi62 & n274;
  assign n436 = pi30 & n276;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~pi71 & ~n437;
  assign n439 = ~n434 & ~n438;
  assign n440 = ~pi68 & ~n439;
  assign n441 = pi46 & pi68;
  assign n442 = ~pi69 & n441;
  assign n443 = ~pi70 & n442;
  assign n444 = ~pi71 & n443;
  assign n445 = pi71 & n223;
  assign n446 = pi14 & ~n252;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~pi68 & ~n447;
  assign n449 = pi69 & n448;
  assign n450 = ~n444 & ~n449;
  assign n451 = n297 & n450;
  assign n452 = ~n297 & ~n450;
  assign n453 = ~n451 & ~n452;
  assign n454 = pi15 & ~pi70;
  assign n455 = ~n232 & ~n454;
  assign n456 = ~pi69 & ~n455;
  assign n457 = pi71 & n456;
  assign n458 = pi63 & n274;
  assign n459 = pi31 & n276;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~pi71 & ~n460;
  assign n462 = ~n457 & ~n461;
  assign n463 = ~pi68 & ~n462;
  assign n464 = pi47 & pi68;
  assign n465 = ~pi69 & n464;
  assign n466 = ~pi70 & n465;
  assign n467 = ~pi71 & n466;
  assign n468 = pi71 & n232;
  assign n469 = pi15 & ~n252;
  assign n470 = ~n468 & ~n469;
  assign n471 = ~pi68 & ~n470;
  assign n472 = pi69 & n471;
  assign n473 = ~n467 & ~n472;
  assign n474 = n297 & n473;
  assign n475 = ~n297 & ~n473;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n440 & n453;
  assign n478 = ~n463 & n476;
  assign n479 = ~n477 & ~n478;
  assign n480 = n430 & n479;
  assign n481 = n381 & n480;
  assign n482 = n463 & ~n476;
  assign n483 = n440 & ~n453;
  assign n484 = ~n477 & n482;
  assign n485 = ~n483 & ~n484;
  assign n486 = ~n429 & ~n485;
  assign n487 = n414 & ~n427;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~n428 & ~n488;
  assign n490 = n391 & ~n404;
  assign n491 = ~n489 & ~n490;
  assign n492 = ~n481 & n491;
  assign n493 = pi08 & ~pi70;
  assign n494 = ~n127 & ~n493;
  assign n495 = ~pi69 & ~n494;
  assign n496 = pi71 & n495;
  assign n497 = pi56 & n274;
  assign n498 = pi24 & n276;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~pi71 & ~n499;
  assign n501 = ~n496 & ~n500;
  assign n502 = ~pi68 & ~n501;
  assign n503 = pi40 & pi68;
  assign n504 = ~pi69 & n503;
  assign n505 = ~pi70 & n504;
  assign n506 = ~pi71 & n505;
  assign n507 = pi71 & n127;
  assign n508 = pi08 & ~n252;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~pi68 & ~n509;
  assign n511 = pi69 & n510;
  assign n512 = ~n506 & ~n511;
  assign n513 = n297 & n512;
  assign n514 = ~n297 & ~n512;
  assign n515 = ~n513 & ~n514;
  assign n516 = pi09 & ~pi70;
  assign n517 = ~n136 & ~n516;
  assign n518 = ~pi69 & ~n517;
  assign n519 = pi71 & n518;
  assign n520 = pi57 & n274;
  assign n521 = pi25 & n276;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~pi71 & ~n522;
  assign n524 = ~n519 & ~n523;
  assign n525 = ~pi68 & ~n524;
  assign n526 = pi41 & pi68;
  assign n527 = ~pi69 & n526;
  assign n528 = ~pi70 & n527;
  assign n529 = ~pi71 & n528;
  assign n530 = pi71 & n136;
  assign n531 = pi09 & ~n252;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~pi68 & ~n532;
  assign n534 = pi69 & n533;
  assign n535 = ~n529 & ~n534;
  assign n536 = n297 & n535;
  assign n537 = ~n297 & ~n535;
  assign n538 = ~n536 & ~n537;
  assign n539 = ~n502 & n515;
  assign n540 = ~n525 & n538;
  assign n541 = ~n539 & ~n540;
  assign n542 = pi10 & ~pi70;
  assign n543 = ~n145 & ~n542;
  assign n544 = ~pi69 & ~n543;
  assign n545 = pi71 & n544;
  assign n546 = pi58 & n274;
  assign n547 = pi26 & n276;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~pi71 & ~n548;
  assign n550 = ~n545 & ~n549;
  assign n551 = ~pi68 & ~n550;
  assign n552 = pi42 & pi68;
  assign n553 = ~pi69 & n552;
  assign n554 = ~pi70 & n553;
  assign n555 = ~pi71 & n554;
  assign n556 = pi71 & n145;
  assign n557 = pi10 & ~n252;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~pi68 & ~n558;
  assign n560 = pi69 & n559;
  assign n561 = ~n555 & ~n560;
  assign n562 = n297 & n561;
  assign n563 = ~n297 & ~n561;
  assign n564 = ~n562 & ~n563;
  assign n565 = pi11 & ~pi70;
  assign n566 = ~n154 & ~n565;
  assign n567 = ~pi69 & ~n566;
  assign n568 = pi71 & n567;
  assign n569 = pi59 & n274;
  assign n570 = pi27 & n276;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~pi71 & ~n571;
  assign n573 = ~n568 & ~n572;
  assign n574 = ~pi68 & ~n573;
  assign n575 = pi43 & pi68;
  assign n576 = ~pi69 & n575;
  assign n577 = ~pi70 & n576;
  assign n578 = ~pi71 & n577;
  assign n579 = pi71 & n154;
  assign n580 = pi11 & ~n252;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~pi68 & ~n581;
  assign n583 = pi69 & n582;
  assign n584 = ~n578 & ~n583;
  assign n585 = n297 & n584;
  assign n586 = ~n297 & ~n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n551 & n564;
  assign n589 = ~n574 & n587;
  assign n590 = ~n588 & ~n589;
  assign n591 = n541 & n590;
  assign n592 = n574 & ~n587;
  assign n593 = n551 & ~n564;
  assign n594 = ~n588 & n592;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n540 & ~n595;
  assign n597 = n525 & ~n538;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~n539 & ~n598;
  assign n600 = n502 & ~n515;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n492 & n591;
  assign n603 = n601 & ~n602;
  assign n604 = pi04 & ~pi70;
  assign n605 = ~n166 & ~n604;
  assign n606 = ~pi69 & ~n605;
  assign n607 = pi71 & n606;
  assign n608 = pi52 & n274;
  assign n609 = pi20 & n276;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~pi71 & ~n610;
  assign n612 = ~n607 & ~n611;
  assign n613 = ~pi68 & ~n612;
  assign n614 = pi36 & pi68;
  assign n615 = ~pi69 & n614;
  assign n616 = ~pi70 & n615;
  assign n617 = ~pi71 & n616;
  assign n618 = pi71 & n166;
  assign n619 = pi04 & ~n252;
  assign n620 = ~n618 & ~n619;
  assign n621 = ~pi68 & ~n620;
  assign n622 = pi69 & n621;
  assign n623 = ~n617 & ~n622;
  assign n624 = n297 & n623;
  assign n625 = ~n297 & ~n623;
  assign n626 = ~n624 & ~n625;
  assign n627 = pi05 & ~pi70;
  assign n628 = ~n175 & ~n627;
  assign n629 = ~pi69 & ~n628;
  assign n630 = pi71 & n629;
  assign n631 = pi53 & n274;
  assign n632 = pi21 & n276;
  assign n633 = ~n631 & ~n632;
  assign n634 = ~pi71 & ~n633;
  assign n635 = ~n630 & ~n634;
  assign n636 = ~pi68 & ~n635;
  assign n637 = pi37 & pi68;
  assign n638 = ~pi69 & n637;
  assign n639 = ~pi70 & n638;
  assign n640 = ~pi71 & n639;
  assign n641 = pi71 & n175;
  assign n642 = pi05 & ~n252;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~pi68 & ~n643;
  assign n645 = pi69 & n644;
  assign n646 = ~n640 & ~n645;
  assign n647 = n297 & n646;
  assign n648 = ~n297 & ~n646;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n613 & n626;
  assign n651 = ~n636 & n649;
  assign n652 = ~n650 & ~n651;
  assign n653 = pi06 & ~pi70;
  assign n654 = ~n184 & ~n653;
  assign n655 = ~pi69 & ~n654;
  assign n656 = pi71 & n655;
  assign n657 = pi54 & n274;
  assign n658 = pi22 & n276;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~pi71 & ~n659;
  assign n661 = ~n656 & ~n660;
  assign n662 = ~pi68 & ~n661;
  assign n663 = pi38 & pi68;
  assign n664 = ~pi69 & n663;
  assign n665 = ~pi70 & n664;
  assign n666 = ~pi71 & n665;
  assign n667 = pi71 & n184;
  assign n668 = pi06 & ~n252;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~pi68 & ~n669;
  assign n671 = pi69 & n670;
  assign n672 = ~n666 & ~n671;
  assign n673 = n297 & n672;
  assign n674 = ~n297 & ~n672;
  assign n675 = ~n673 & ~n674;
  assign n676 = pi07 & ~pi70;
  assign n677 = ~n193 & ~n676;
  assign n678 = ~pi69 & ~n677;
  assign n679 = pi71 & n678;
  assign n680 = pi55 & n274;
  assign n681 = pi23 & n276;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~pi71 & ~n682;
  assign n684 = ~n679 & ~n683;
  assign n685 = ~pi68 & ~n684;
  assign n686 = pi39 & pi68;
  assign n687 = ~pi69 & n686;
  assign n688 = ~pi70 & n687;
  assign n689 = ~pi71 & n688;
  assign n690 = pi71 & n193;
  assign n691 = pi07 & ~n252;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~pi68 & ~n692;
  assign n694 = pi69 & n693;
  assign n695 = ~n689 & ~n694;
  assign n696 = n297 & n695;
  assign n697 = ~n297 & ~n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~n662 & n675;
  assign n700 = ~n685 & n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n603 & n652;
  assign n703 = n701 & n702;
  assign n704 = n685 & ~n698;
  assign n705 = ~n699 & n704;
  assign n706 = n662 & ~n675;
  assign n707 = ~n705 & ~n706;
  assign n708 = ~n651 & ~n707;
  assign n709 = n636 & ~n649;
  assign n710 = ~n708 & ~n709;
  assign n711 = ~n650 & ~n710;
  assign n712 = n613 & ~n626;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n703 & n713;
  assign n715 = n364 & ~n374;
  assign n716 = ~n375 & n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = n340 & ~n350;
  assign n719 = ~n351 & ~n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = n316 & ~n326;
  assign n722 = ~n327 & ~n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~n714 & ~n715;
  assign n725 = ~n375 & ~n724;
  assign n726 = ~n718 & ~n725;
  assign n727 = ~n351 & ~n726;
  assign n728 = ~n721 & ~n727;
  assign n729 = ~n327 & ~n728;
  assign n730 = n303 & ~n729;
  assign n731 = ~n303 & ~n723;
  assign n732 = ~n730 & ~n731;
  assign n733 = pi66 & ~pi67;
  assign n734 = ~pi66 & pi67;
  assign n735 = ~n733 & ~n734;
  assign n736 = n92 & ~n262;
  assign n737 = ~n732 & ~n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~pi65 & ~n738;
  assign n740 = pi64 & n739;
  assign n741 = ~pi64 & ~n269;
  assign po00 = n740 | n741;
  assign n743 = pi49 & pi70;
  assign n744 = pi71 & n743;
  assign n745 = pi17 & ~n252;
  assign n746 = ~n744 & ~n745;
  assign n747 = pi49 & pi68;
  assign n748 = n258 & n747;
  assign n749 = n256 & ~n746;
  assign n750 = ~n748 & ~n749;
  assign n751 = pi72 & ~pi74;
  assign n752 = ~pi73 & pi74;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~pi72 & pi73;
  assign n755 = n753 & ~n754;
  assign n756 = ~n262 & ~n755;
  assign n757 = ~n750 & n755;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n117 & n246;
  assign n760 = ~n126 & n759;
  assign n761 = ~n108 & ~n760;
  assign n762 = n108 & n760;
  assign n763 = ~n761 & ~n762;
  assign n764 = pi65 & ~n758;
  assign n765 = ~pi65 & ~n763;
  assign n766 = ~n764 & ~n765;
  assign n767 = pi65 & ~n763;
  assign n768 = n92 & n767;
  assign n769 = ~n92 & ~n766;
  assign n770 = ~n768 & ~n769;
  assign n771 = n316 & n326;
  assign n772 = ~n316 & ~n326;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~n727 & n773;
  assign n775 = ~n720 & ~n773;
  assign n776 = ~n774 & ~n775;
  assign n777 = n92 & ~n758;
  assign n778 = ~n735 & ~n776;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~pi65 & ~n779;
  assign n781 = pi64 & n780;
  assign n782 = ~pi64 & ~n770;
  assign po01 = n781 | n782;
  assign n784 = pi72 & pi74;
  assign n785 = pi50 & pi70;
  assign n786 = pi71 & n785;
  assign n787 = pi18 & ~n252;
  assign n788 = ~n786 & ~n787;
  assign n789 = pi50 & pi68;
  assign n790 = n258 & n789;
  assign n791 = n256 & ~n788;
  assign n792 = ~n790 & ~n791;
  assign n793 = pi73 & ~n792;
  assign n794 = pi73 & ~n784;
  assign n795 = pi72 & ~pi73;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~pi74 & ~n792;
  assign n798 = pi74 & ~n750;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~pi72 & ~pi73;
  assign n801 = ~n262 & ~n796;
  assign n802 = ~n799 & n800;
  assign n803 = ~n801 & ~n802;
  assign n804 = n784 & n793;
  assign n805 = n803 & ~n804;
  assign n806 = ~n117 & ~n248;
  assign n807 = n117 & n248;
  assign n808 = ~n806 & ~n807;
  assign n809 = pi65 & ~n805;
  assign n810 = ~pi65 & ~n808;
  assign n811 = ~n809 & ~n810;
  assign n812 = pi65 & ~n808;
  assign n813 = n92 & n812;
  assign n814 = ~n92 & ~n811;
  assign n815 = ~n813 & ~n814;
  assign n816 = n340 & n350;
  assign n817 = ~n340 & ~n350;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n725 & n818;
  assign n820 = ~n717 & ~n818;
  assign n821 = ~n819 & ~n820;
  assign n822 = n92 & ~n805;
  assign n823 = ~n735 & ~n821;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~pi65 & ~n824;
  assign n826 = pi64 & n825;
  assign n827 = ~pi64 & ~n815;
  assign po02 = n826 | n827;
  assign n829 = pi51 & pi70;
  assign n830 = pi71 & n829;
  assign n831 = pi19 & ~n252;
  assign n832 = ~n830 & ~n831;
  assign n833 = pi51 & pi68;
  assign n834 = n258 & n833;
  assign n835 = n256 & ~n832;
  assign n836 = ~n834 & ~n835;
  assign n837 = pi73 & pi74;
  assign n838 = ~n836 & n837;
  assign n839 = ~n262 & ~n837;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~pi73 & ~n836;
  assign n842 = pi73 & ~n750;
  assign n843 = ~n841 & ~n842;
  assign n844 = n752 & ~n792;
  assign n845 = ~n262 & n837;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~pi74 & ~n843;
  assign n848 = n846 & ~n847;
  assign n849 = pi72 & ~n840;
  assign n850 = ~pi72 & ~n848;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n364 & ~n374;
  assign n853 = n364 & n374;
  assign n854 = ~n852 & ~n853;
  assign n855 = ~n714 & n854;
  assign n856 = n714 & ~n854;
  assign n857 = ~n855 & ~n856;
  assign n858 = n92 & ~n851;
  assign n859 = ~n735 & ~n857;
  assign n860 = ~n858 & ~n859;
  assign n861 = pi64 & ~pi65;
  assign n862 = ~n126 & ~n246;
  assign n863 = n126 & n246;
  assign n864 = ~n862 & ~n863;
  assign n865 = pi65 & ~n851;
  assign n866 = ~pi65 & ~n864;
  assign n867 = ~n865 & ~n866;
  assign n868 = pi65 & ~n864;
  assign n869 = n92 & n868;
  assign n870 = ~n92 & ~n867;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n860 & n861;
  assign n873 = ~pi64 & ~n871;
  assign po03 = n872 | n873;
  assign n875 = pi52 & pi70;
  assign n876 = pi71 & n875;
  assign n877 = pi20 & ~n252;
  assign n878 = ~n876 & ~n877;
  assign n879 = pi52 & pi68;
  assign n880 = n258 & n879;
  assign n881 = n256 & ~n878;
  assign n882 = ~n880 & ~n881;
  assign n883 = ~pi72 & ~n750;
  assign n884 = pi72 & ~n882;
  assign n885 = ~n883 & ~n884;
  assign n886 = pi72 & ~n262;
  assign n887 = ~pi73 & ~n882;
  assign n888 = ~n793 & ~n887;
  assign n889 = n752 & ~n836;
  assign n890 = ~pi74 & ~n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n837 & n886;
  assign n893 = ~pi72 & ~n891;
  assign n894 = ~n892 & ~n893;
  assign n895 = n837 & ~n885;
  assign n896 = n894 & ~n895;
  assign n897 = n204 & n243;
  assign n898 = n105 & n897;
  assign n899 = ~n183 & ~n192;
  assign n900 = ~n201 & n898;
  assign n901 = n899 & n900;
  assign n902 = ~n174 & ~n901;
  assign n903 = n174 & n901;
  assign n904 = ~n902 & ~n903;
  assign n905 = pi65 & ~n896;
  assign n906 = ~pi65 & ~n904;
  assign n907 = ~n905 & ~n906;
  assign n908 = pi65 & ~n904;
  assign n909 = n92 & n908;
  assign n910 = ~n92 & ~n907;
  assign n911 = ~n909 & ~n910;
  assign n912 = n613 & n626;
  assign n913 = ~n613 & ~n626;
  assign n914 = ~n912 & ~n913;
  assign n915 = n603 & ~n704;
  assign n916 = ~n700 & ~n915;
  assign n917 = ~n706 & ~n916;
  assign n918 = ~n699 & ~n917;
  assign n919 = ~n709 & ~n918;
  assign n920 = ~n651 & ~n919;
  assign n921 = ~n603 & ~n700;
  assign n922 = ~n704 & ~n921;
  assign n923 = ~n699 & ~n922;
  assign n924 = ~n706 & ~n923;
  assign n925 = ~n651 & ~n924;
  assign n926 = ~n709 & ~n925;
  assign n927 = n914 & ~n926;
  assign n928 = ~n914 & ~n920;
  assign n929 = ~n927 & ~n928;
  assign n930 = n92 & ~n896;
  assign n931 = ~n735 & ~n929;
  assign n932 = ~n930 & ~n931;
  assign n933 = ~pi65 & ~n932;
  assign n934 = pi64 & n933;
  assign n935 = ~pi64 & ~n911;
  assign po04 = n934 | n935;
  assign n937 = pi53 & pi70;
  assign n938 = pi71 & n937;
  assign n939 = pi21 & ~n252;
  assign n940 = ~n938 & ~n939;
  assign n941 = pi53 & pi68;
  assign n942 = n258 & n941;
  assign n943 = n256 & ~n940;
  assign n944 = ~n942 & ~n943;
  assign n945 = pi72 & ~n944;
  assign n946 = ~pi72 & ~n792;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~pi72 & ~n882;
  assign n949 = ~n886 & ~n948;
  assign n950 = pi73 & ~n947;
  assign n951 = ~pi73 & ~n949;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~pi72 & ~n836;
  assign n954 = ~n886 & ~n953;
  assign n955 = ~pi72 & ~n944;
  assign n956 = pi72 & ~n750;
  assign n957 = ~n955 & ~n956;
  assign n958 = pi73 & ~n954;
  assign n959 = ~pi73 & ~n957;
  assign n960 = ~n958 & ~n959;
  assign n961 = pi74 & ~n952;
  assign n962 = ~pi74 & ~n960;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~n192 & n898;
  assign n965 = ~n201 & n964;
  assign n966 = ~n183 & ~n965;
  assign n967 = n183 & n965;
  assign n968 = ~n966 & ~n967;
  assign n969 = pi65 & ~n963;
  assign n970 = ~pi65 & ~n968;
  assign n971 = ~n969 & ~n970;
  assign n972 = pi65 & ~n968;
  assign n973 = n92 & n972;
  assign n974 = ~n92 & ~n971;
  assign n975 = ~n973 & ~n974;
  assign n976 = n636 & n649;
  assign n977 = ~n636 & ~n649;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n924 & n978;
  assign n980 = ~n918 & ~n978;
  assign n981 = ~n979 & ~n980;
  assign n982 = n92 & ~n963;
  assign n983 = ~n735 & ~n981;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~pi65 & ~n984;
  assign n986 = pi64 & n985;
  assign n987 = ~pi64 & ~n975;
  assign po05 = n986 | n987;
  assign n989 = pi54 & pi70;
  assign n990 = pi71 & n989;
  assign n991 = pi22 & ~n252;
  assign n992 = ~n990 & ~n991;
  assign n993 = pi54 & pi68;
  assign n994 = n258 & n993;
  assign n995 = n256 & ~n992;
  assign n996 = ~n994 & ~n995;
  assign n997 = pi72 & ~n996;
  assign n998 = ~n953 & ~n997;
  assign n999 = pi73 & ~n998;
  assign n1000 = ~n959 & ~n999;
  assign n1001 = ~pi72 & ~n996;
  assign n1002 = pi72 & ~n792;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = pi73 & ~n949;
  assign n1005 = ~pi73 & ~n1003;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = pi74 & ~n1000;
  assign n1008 = ~pi74 & ~n1006;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = ~n192 & ~n900;
  assign n1011 = n192 & n900;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = pi65 & ~n1009;
  assign n1014 = ~pi65 & ~n1012;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = pi65 & ~n1012;
  assign n1017 = n92 & n1016;
  assign n1018 = ~n92 & ~n1015;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n662 & n675;
  assign n1021 = ~n662 & ~n675;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n922 & n1022;
  assign n1024 = ~n916 & ~n1022;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n92 & ~n1009;
  assign n1027 = ~n735 & ~n1025;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~pi65 & ~n1028;
  assign n1030 = pi64 & n1029;
  assign n1031 = ~pi64 & ~n1019;
  assign po06 = n1030 | n1031;
  assign n1033 = pi55 & pi70;
  assign n1034 = pi71 & n1033;
  assign n1035 = pi23 & ~n252;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = pi55 & pi68;
  assign n1038 = n258 & n1037;
  assign n1039 = n256 & ~n1036;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = pi72 & ~n1040;
  assign n1042 = ~n948 & ~n1041;
  assign n1043 = pi73 & ~n1042;
  assign n1044 = ~n1005 & ~n1043;
  assign n1045 = ~n886 & ~n955;
  assign n1046 = ~pi72 & ~n1040;
  assign n1047 = pi72 & ~n836;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = pi73 & ~n1045;
  assign n1050 = ~pi73 & ~n1048;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = pi74 & ~n1044;
  assign n1053 = ~pi74 & ~n1051;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = n685 & n698;
  assign n1056 = ~n685 & ~n698;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = ~n603 & n1057;
  assign n1059 = n603 & ~n1057;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = n92 & ~n1054;
  assign n1062 = ~n735 & ~n1060;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n201 & ~n898;
  assign n1065 = n201 & n898;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = pi65 & ~n1054;
  assign n1068 = ~pi65 & ~n1066;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = pi65 & ~n1066;
  assign n1071 = n92 & n1070;
  assign n1072 = ~n92 & ~n1069;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = n861 & ~n1063;
  assign n1075 = ~pi64 & ~n1073;
  assign po07 = n1074 | n1075;
  assign n1077 = pi56 & pi70;
  assign n1078 = pi71 & n1077;
  assign n1079 = pi24 & ~n252;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = pi56 & pi68;
  assign n1082 = n258 & n1081;
  assign n1083 = n256 & ~n1080;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = pi72 & ~n1084;
  assign n1086 = ~n955 & ~n1085;
  assign n1087 = pi73 & ~n1086;
  assign n1088 = ~n1050 & ~n1087;
  assign n1089 = ~n886 & ~n1001;
  assign n1090 = ~pi72 & ~n1084;
  assign n1091 = ~n884 & ~n1090;
  assign n1092 = pi73 & ~n1089;
  assign n1093 = ~pi73 & ~n1091;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = pi74 & ~n1088;
  assign n1096 = ~pi74 & ~n1094;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = n105 & n243;
  assign n1099 = ~n144 & ~n153;
  assign n1100 = ~n162 & n1098;
  assign n1101 = n1099 & n1100;
  assign n1102 = ~n135 & ~n1101;
  assign n1103 = n135 & n1101;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = pi65 & ~n1097;
  assign n1106 = ~pi65 & ~n1104;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = pi65 & ~n1104;
  assign n1109 = n92 & n1108;
  assign n1110 = ~n92 & ~n1107;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = n502 & n515;
  assign n1113 = ~n502 & ~n515;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = n492 & ~n592;
  assign n1116 = ~n589 & ~n1115;
  assign n1117 = ~n593 & ~n1116;
  assign n1118 = ~n588 & ~n1117;
  assign n1119 = ~n597 & ~n1118;
  assign n1120 = ~n540 & ~n1119;
  assign n1121 = ~n492 & ~n589;
  assign n1122 = ~n592 & ~n1121;
  assign n1123 = ~n588 & ~n1122;
  assign n1124 = ~n593 & ~n1123;
  assign n1125 = ~n540 & ~n1124;
  assign n1126 = ~n597 & ~n1125;
  assign n1127 = n1114 & ~n1126;
  assign n1128 = ~n1114 & ~n1120;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = n92 & ~n1097;
  assign n1131 = ~n735 & ~n1129;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~pi65 & ~n1132;
  assign n1134 = pi64 & n1133;
  assign n1135 = ~pi64 & ~n1111;
  assign po08 = n1134 | n1135;
  assign n1137 = pi57 & pi70;
  assign n1138 = pi71 & n1137;
  assign n1139 = pi25 & ~n252;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = pi57 & pi68;
  assign n1142 = n258 & n1141;
  assign n1143 = n256 & ~n1140;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = pi72 & ~n1144;
  assign n1146 = ~n1001 & ~n1145;
  assign n1147 = pi73 & ~n1146;
  assign n1148 = ~n1093 & ~n1147;
  assign n1149 = ~n956 & ~n1046;
  assign n1150 = ~pi72 & ~n1144;
  assign n1151 = ~n945 & ~n1150;
  assign n1152 = pi73 & ~n1149;
  assign n1153 = ~pi73 & ~n1151;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = pi74 & ~n1148;
  assign n1156 = ~pi74 & ~n1154;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n153 & n1098;
  assign n1159 = ~n162 & n1158;
  assign n1160 = ~n144 & ~n1159;
  assign n1161 = n144 & n1159;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = pi65 & ~n1157;
  assign n1164 = ~pi65 & ~n1162;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = pi65 & ~n1162;
  assign n1167 = n92 & n1166;
  assign n1168 = ~n92 & ~n1165;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = n525 & n538;
  assign n1171 = ~n525 & ~n538;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n1124 & n1172;
  assign n1174 = ~n1118 & ~n1172;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = n92 & ~n1157;
  assign n1177 = ~n735 & ~n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~pi65 & ~n1178;
  assign n1180 = pi64 & n1179;
  assign n1181 = ~pi64 & ~n1169;
  assign po09 = n1180 | n1181;
  assign n1183 = pi58 & pi70;
  assign n1184 = pi71 & n1183;
  assign n1185 = pi26 & ~n252;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = pi58 & pi68;
  assign n1188 = n258 & n1187;
  assign n1189 = n256 & ~n1186;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = pi72 & ~n1190;
  assign n1192 = ~n1046 & ~n1191;
  assign n1193 = pi73 & ~n1192;
  assign n1194 = ~n1153 & ~n1193;
  assign n1195 = ~n1002 & ~n1090;
  assign n1196 = ~pi72 & ~n1190;
  assign n1197 = ~n997 & ~n1196;
  assign n1198 = pi73 & ~n1195;
  assign n1199 = ~pi73 & ~n1197;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = pi74 & ~n1194;
  assign n1202 = ~pi74 & ~n1200;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~n153 & ~n1100;
  assign n1205 = n153 & n1100;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = pi65 & ~n1203;
  assign n1208 = ~pi65 & ~n1206;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = pi65 & ~n1206;
  assign n1211 = n92 & n1210;
  assign n1212 = ~n92 & ~n1209;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = n551 & n564;
  assign n1215 = ~n551 & ~n564;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1122 & n1216;
  assign n1218 = ~n1116 & ~n1216;
  assign n1219 = ~n1217 & ~n1218;
  assign n1220 = n92 & ~n1203;
  assign n1221 = ~n735 & ~n1219;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~pi65 & ~n1222;
  assign n1224 = pi64 & n1223;
  assign n1225 = ~pi64 & ~n1213;
  assign po10 = n1224 | n1225;
  assign n1227 = pi59 & pi70;
  assign n1228 = pi71 & n1227;
  assign n1229 = pi27 & ~n252;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = pi59 & pi68;
  assign n1232 = n258 & n1231;
  assign n1233 = n256 & ~n1230;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = pi72 & ~n1234;
  assign n1236 = ~n1090 & ~n1235;
  assign n1237 = pi73 & ~n1236;
  assign n1238 = ~n1199 & ~n1237;
  assign n1239 = ~n1047 & ~n1150;
  assign n1240 = ~pi72 & ~n1234;
  assign n1241 = ~n1041 & ~n1240;
  assign n1242 = pi73 & ~n1239;
  assign n1243 = ~pi73 & ~n1241;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = pi74 & ~n1238;
  assign n1246 = ~pi74 & ~n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n574 & ~n587;
  assign n1249 = n574 & n587;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~n492 & n1250;
  assign n1252 = n492 & ~n1250;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = n92 & ~n1247;
  assign n1255 = ~n735 & ~n1253;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n162 & ~n1098;
  assign n1258 = n162 & n1098;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = pi65 & ~n1247;
  assign n1261 = ~pi65 & ~n1259;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = pi65 & ~n1259;
  assign n1264 = n92 & n1263;
  assign n1265 = ~n92 & ~n1262;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n861 & ~n1256;
  assign n1268 = ~pi64 & ~n1266;
  assign po11 = n1267 | n1268;
  assign n1270 = pi60 & pi70;
  assign n1271 = pi71 & n1270;
  assign n1272 = pi28 & ~n252;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = pi60 & pi68;
  assign n1275 = n258 & n1274;
  assign n1276 = n256 & ~n1273;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = pi72 & ~n1277;
  assign n1279 = ~n1150 & ~n1278;
  assign n1280 = pi73 & ~n1279;
  assign n1281 = ~n1243 & ~n1280;
  assign n1282 = ~n884 & ~n1196;
  assign n1283 = ~pi72 & ~n1277;
  assign n1284 = ~n1085 & ~n1283;
  assign n1285 = pi73 & ~n1282;
  assign n1286 = ~pi73 & ~n1284;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = pi74 & ~n1281;
  assign n1289 = ~pi74 & ~n1287;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n222 & ~n231;
  assign n1292 = n105 & ~n240;
  assign n1293 = n1291 & n1292;
  assign n1294 = ~n213 & ~n1293;
  assign n1295 = n213 & n1293;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = pi65 & ~n1290;
  assign n1298 = ~pi65 & ~n1296;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = pi65 & ~n1296;
  assign n1301 = n92 & n1300;
  assign n1302 = ~n92 & ~n1299;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = n391 & n404;
  assign n1305 = ~n391 & ~n404;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = ~n381 & ~n482;
  assign n1308 = ~n478 & ~n1307;
  assign n1309 = ~n483 & ~n1308;
  assign n1310 = ~n477 & ~n1309;
  assign n1311 = ~n487 & ~n1310;
  assign n1312 = ~n429 & ~n1311;
  assign n1313 = n381 & ~n478;
  assign n1314 = ~n482 & ~n1313;
  assign n1315 = ~n477 & ~n1314;
  assign n1316 = ~n483 & ~n1315;
  assign n1317 = ~n429 & ~n1316;
  assign n1318 = ~n487 & ~n1317;
  assign n1319 = n1306 & ~n1318;
  assign n1320 = ~n1306 & ~n1312;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n92 & ~n1290;
  assign n1323 = ~n735 & ~n1321;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~pi65 & ~n1324;
  assign n1326 = pi64 & n1325;
  assign n1327 = ~pi64 & ~n1303;
  assign po12 = n1326 | n1327;
  assign n1329 = pi61 & pi70;
  assign n1330 = pi71 & n1329;
  assign n1331 = pi29 & ~n252;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = pi61 & pi68;
  assign n1334 = n258 & n1333;
  assign n1335 = n256 & ~n1332;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = pi72 & ~n1336;
  assign n1338 = ~n1196 & ~n1337;
  assign n1339 = pi73 & ~n1338;
  assign n1340 = ~n1286 & ~n1339;
  assign n1341 = ~n945 & ~n1240;
  assign n1342 = ~pi72 & ~n1336;
  assign n1343 = ~n1145 & ~n1342;
  assign n1344 = pi73 & ~n1341;
  assign n1345 = ~pi73 & ~n1343;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = pi74 & ~n1340;
  assign n1348 = ~pi74 & ~n1346;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = n105 & ~n231;
  assign n1351 = ~n240 & n1350;
  assign n1352 = ~n222 & ~n1351;
  assign n1353 = n222 & n1351;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = pi65 & ~n1349;
  assign n1356 = ~pi65 & ~n1354;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = pi65 & ~n1354;
  assign n1359 = n92 & n1358;
  assign n1360 = ~n92 & ~n1357;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = n414 & n427;
  assign n1363 = ~n414 & ~n427;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~n1316 & n1364;
  assign n1366 = ~n1310 & ~n1364;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = n92 & ~n1349;
  assign n1369 = ~n735 & ~n1367;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~pi65 & ~n1370;
  assign n1372 = pi64 & n1371;
  assign n1373 = ~pi64 & ~n1361;
  assign po13 = n1372 | n1373;
  assign n1375 = pi62 & pi70;
  assign n1376 = pi71 & n1375;
  assign n1377 = pi30 & ~n252;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = pi62 & pi68;
  assign n1380 = n258 & n1379;
  assign n1381 = n256 & ~n1378;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = pi72 & ~n1382;
  assign n1384 = ~n1240 & ~n1383;
  assign n1385 = pi73 & ~n1384;
  assign n1386 = ~n1345 & ~n1385;
  assign n1387 = ~n997 & ~n1283;
  assign n1388 = ~pi72 & ~n1382;
  assign n1389 = ~n1191 & ~n1388;
  assign n1390 = pi73 & ~n1387;
  assign n1391 = ~pi73 & ~n1389;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = pi74 & ~n1386;
  assign n1394 = ~pi74 & ~n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = ~n231 & ~n1292;
  assign n1397 = n231 & n1292;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = pi65 & ~n1395;
  assign n1400 = ~pi65 & ~n1398;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = pi65 & ~n1398;
  assign n1403 = n92 & n1402;
  assign n1404 = ~n92 & ~n1401;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = n440 & n453;
  assign n1407 = ~n440 & ~n453;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = ~n1314 & n1408;
  assign n1410 = ~n1308 & ~n1408;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = n92 & ~n1395;
  assign n1413 = ~n735 & ~n1411;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~pi65 & ~n1414;
  assign n1416 = pi64 & n1415;
  assign n1417 = ~pi64 & ~n1405;
  assign po14 = n1416 | n1417;
  assign n1419 = pi63 & pi70;
  assign n1420 = pi71 & n1419;
  assign n1421 = pi31 & ~n252;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = pi63 & pi68;
  assign n1424 = n258 & n1423;
  assign n1425 = n256 & ~n1422;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = pi72 & ~n1426;
  assign n1428 = ~n1283 & ~n1427;
  assign n1429 = pi73 & ~n1428;
  assign n1430 = ~n1391 & ~n1429;
  assign n1431 = ~n1041 & ~n1342;
  assign n1432 = ~pi72 & ~n1426;
  assign n1433 = ~n1235 & ~n1432;
  assign n1434 = pi73 & ~n1431;
  assign n1435 = ~pi73 & ~n1433;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = pi74 & ~n1430;
  assign n1438 = ~pi74 & ~n1436;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~n105 & ~n240;
  assign n1441 = n105 & n240;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = pi65 & ~n1439;
  assign n1444 = ~pi65 & ~n1442;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = pi65 & ~n1442;
  assign n1447 = n92 & n1446;
  assign n1448 = ~n92 & ~n1445;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~n463 & ~n476;
  assign n1451 = n463 & n476;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = n381 & n1452;
  assign n1454 = ~n381 & ~n1452;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = n92 & ~n1439;
  assign n1457 = ~n735 & ~n1455;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~pi65 & ~n1458;
  assign n1460 = pi64 & n1459;
  assign n1461 = ~pi64 & ~n1449;
  assign po15 = n1460 | n1461;
endmodule



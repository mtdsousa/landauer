// written by CirKit Wed Nov  2 14:26:17 2016

module arbiter_best_speed_2015.1.blif_ (
        pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, 
        po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178;
assign w0 = pi049 & ~pi177;
assign w1 = pi050 & ~pi178;
assign w2 = (~pi178 & w0) | (~pi178 & w1) | (w0 & w1);
assign w3 = ~pi052 & pi179;
assign w4 = pi051 & ~pi179;
assign w5 = ~pi052 & ~w4;
assign w6 = (~w2 & w3) | (~w2 & w5) | (w3 & w5);
assign w7 = ~pi180 & ~pi181;
assign w8 = ~pi182 & ~pi183;
assign w9 = w7 & w8;
assign w10 = ~w6 & w9;
assign w11 = pi053 & ~pi181;
assign w12 = pi054 & ~pi183;
assign w13 = (~pi183 & w11) | (~pi183 & w12) | (w11 & w12);
assign w14 = ~pi182 & w13;
assign w15 = pi055 & ~pi183;
assign w16 = ~pi056 & ~w15;
assign w17 = ~w14 & w16;
assign w18 = ~w10 & w17;
assign w19 = ~pi192 & ~pi193;
assign w20 = ~pi194 & ~pi195;
assign w21 = w19 & w20;
assign w22 = ~pi196 & ~pi197;
assign w23 = ~pi198 & ~pi199;
assign w24 = w22 & w23;
assign w25 = w21 & w24;
assign w26 = ~pi188 & ~pi189;
assign w27 = ~pi190 & ~pi191;
assign w28 = w26 & w27;
assign w29 = ~pi184 & ~pi185;
assign w30 = ~pi186 & ~pi187;
assign w31 = w29 & w30;
assign w32 = w28 & w31;
assign w33 = w25 & w32;
assign w34 = ~w18 & w33;
assign w35 = pi057 & ~pi185;
assign w36 = pi058 & ~pi186;
assign w37 = (~pi186 & w35) | (~pi186 & w36) | (w35 & w36);
assign w38 = ~pi060 & pi187;
assign w39 = pi059 & ~pi187;
assign w40 = ~pi060 & ~w39;
assign w41 = (~w37 & w38) | (~w37 & w40) | (w38 & w40);
assign w42 = w28 & ~w41;
assign w43 = pi061 & ~pi189;
assign w44 = pi062 & ~pi190;
assign w45 = (~pi190 & w43) | (~pi190 & w44) | (w43 & w44);
assign w46 = ~pi064 & pi191;
assign w47 = pi063 & ~pi191;
assign w48 = ~pi064 & ~w47;
assign w49 = (~w45 & w46) | (~w45 & w48) | (w46 & w48);
assign w50 = w25 & ~w49;
assign w51 = (w25 & w42) | (w25 & w50) | (w42 & w50);
assign w52 = pi065 & ~pi193;
assign w53 = pi066 & ~pi194;
assign w54 = (~pi194 & w52) | (~pi194 & w53) | (w52 & w53);
assign w55 = ~pi068 & pi195;
assign w56 = pi067 & ~pi195;
assign w57 = ~pi068 & ~w56;
assign w58 = (~w54 & w55) | (~w54 & w57) | (w55 & w57);
assign w59 = w24 & ~w58;
assign w60 = pi069 & ~pi197;
assign w61 = pi070 & ~pi198;
assign w62 = (~pi198 & w60) | (~pi198 & w61) | (w60 & w61);
assign w63 = ~pi072 & pi199;
assign w64 = pi071 & ~pi199;
assign w65 = ~pi072 & ~w64;
assign w66 = (~w62 & w63) | (~w62 & w65) | (w63 & w65);
assign w67 = ~w59 & w66;
assign w68 = ~w51 & w67;
assign w69 = ~w34 & w68;
assign w70 = pi041 & ~pi169;
assign w71 = ~pi042 & ~w70;
assign w72 = ~pi170 & ~pi171;
assign w73 = ~pi172 & ~pi173;
assign w74 = w72 & w73;
assign w75 = ~pi174 & ~pi175;
assign w76 = w74 & w75;
assign w77 = ~w71 & w76;
assign w78 = pi043 & ~pi171;
assign w79 = ~pi044 & ~w78;
assign w80 = w73 & w75;
assign w81 = ~w79 & w80;
assign w82 = ~pi048 & ~w81;
assign w83 = ~w77 & w82;
assign w84 = pi045 & ~pi173;
assign w85 = pi046 & ~pi174;
assign w86 = (~pi174 & w84) | (~pi174 & w85) | (w84 & w85);
assign w87 = pi047 & ~pi175;
assign w88 = (~pi175 & w86) | (~pi175 & w87) | (w86 & w87);
assign w89 = w83 & ~w88;
assign w90 = ~pi176 & ~pi177;
assign w91 = ~pi178 & ~pi179;
assign w92 = w90 & w91;
assign w93 = w9 & w92;
assign w94 = w33 & w93;
assign w95 = ~w89 & w94;
assign w96 = w69 & ~w95;
assign w97 = ~pi226 & ~pi233;
assign w98 = ~pi234 & ~pi235;
assign w99 = w97 & w98;
assign w100 = ~pi236 & w99;
assign w101 = ~pi227 & ~pi228;
assign w102 = ~pi229 & ~pi230;
assign w103 = w101 & w102;
assign w104 = ~pi231 & ~pi232;
assign w105 = w103 & w104;
assign w106 = w100 & w105;
assign w107 = ~pi220 & ~pi223;
assign w108 = ~pi224 & ~pi225;
assign w109 = w107 & w108;
assign w110 = w106 & w109;
assign w111 = ~pi247 & ~pi248;
assign w112 = ~pi249 & ~pi250;
assign w113 = w111 & w112;
assign w114 = ~pi245 & ~pi246;
assign w115 = ~pi251 & w114;
assign w116 = w113 & w115;
assign w117 = ~pi240 & ~pi241;
assign w118 = ~pi242 & ~pi243;
assign w119 = w117 & w118;
assign w120 = ~pi244 & w119;
assign w121 = w116 & w120;
assign w122 = ~pi221 & ~pi222;
assign w123 = ~pi238 & ~pi239;
assign w124 = w122 & w123;
assign w125 = ~pi237 & w124;
assign w126 = w121 & w125;
assign w127 = w110 & w126;
assign w128 = ~pi211 & ~pi212;
assign w129 = ~pi213 & ~pi214;
assign w130 = w128 & w129;
assign w131 = ~pi215 & ~pi219;
assign w132 = w130 & w131;
assign w133 = ~pi208 & ~pi209;
assign w134 = ~pi210 & ~pi216;
assign w135 = w133 & w134;
assign w136 = ~pi217 & ~pi218;
assign w137 = w135 & w136;
assign w138 = w132 & w137;
assign w139 = ~pi203 & ~pi204;
assign w140 = ~pi205 & ~pi206;
assign w141 = w139 & w140;
assign w142 = ~pi207 & w141;
assign w143 = ~pi200 & ~pi201;
assign w144 = ~pi202 & w143;
assign w145 = w142 & w144;
assign w146 = w138 & w145;
assign w147 = w127 & w146;
assign w148 = ~w96 & w147;
assign w149 = pi099 & w104;
assign w150 = w103 & w149;
assign w151 = ~pi106 & ~pi107;
assign w152 = ~w150 & w151;
assign w153 = pi101 & ~pi229;
assign w154 = pi102 & ~pi230;
assign w155 = (~pi230 & w153) | (~pi230 & w154) | (w153 & w154);
assign w156 = ~pi103 & ~w155;
assign w157 = pi100 & ~pi228;
assign w158 = w102 & w157;
assign w159 = ~pi104 & ~pi105;
assign w160 = ~w158 & w159;
assign w161 = w156 & w160;
assign w162 = w152 & w161;
assign w163 = ~pi235 & ~pi236;
assign w164 = ~pi237 & w163;
assign w165 = ~pi104 & pi231;
assign w166 = ~pi105 & pi232;
assign w167 = (~pi105 & w165) | (~pi105 & w166) | (w165 & w166);
assign w168 = pi106 & ~pi234;
assign w169 = ~pi106 & pi233;
assign w170 = ~pi234 & ~w169;
assign w171 = (~w167 & w168) | (~w167 & w170) | (w168 & w170);
assign w172 = pi107 & ~pi237;
assign w173 = w163 & w172;
assign w174 = (w164 & w171) | (w164 & w173) | (w171 & w173);
assign w175 = ~w162 & w174;
assign w176 = pi108 & ~pi236;
assign w177 = pi109 & ~pi237;
assign w178 = (~pi237 & w176) | (~pi237 & w177) | (w176 & w177);
assign w179 = pi094 & ~pi222;
assign w180 = ~pi095 & ~pi098;
assign w181 = ~w179 & w180;
assign w182 = ~pi096 & ~pi097;
assign w183 = w181 & w182;
assign w184 = pi093 & ~pi221;
assign w185 = ~pi222 & w184;
assign w186 = w183 & ~w185;
assign w187 = ~pi096 & pi223;
assign w188 = ~pi097 & pi224;
assign w189 = (~pi097 & w187) | (~pi097 & w188) | (w187 & w188);
assign w190 = ~pi098 & pi225;
assign w191 = (~pi098 & w189) | (~pi098 & w190) | (w189 & w190);
assign w192 = w105 & ~w191;
assign w193 = ~w186 & w192;
assign w194 = ~pi236 & ~pi237;
assign w195 = w99 & w194;
assign w196 = ~w178 & ~w195;
assign w197 = (~w178 & ~w193) | (~w178 & w196) | (~w193 & w196);
assign w198 = ~w175 & w197;
assign w199 = w121 & w123;
assign w200 = ~w198 & w199;
assign w201 = pi089 & ~pi217;
assign w202 = pi090 & ~pi218;
assign w203 = (~pi218 & w201) | (~pi218 & w202) | (w201 & w202);
assign w204 = ~pi091 & ~w203;
assign w205 = ~pi092 & pi219;
assign w206 = ~pi216 & ~pi217;
assign w207 = ~pi218 & ~pi219;
assign w208 = w206 & w207;
assign w209 = ~pi092 & ~w208;
assign w210 = (w204 & w205) | (w204 & w209) | (w205 & w209);
assign w211 = pi085 & ~pi213;
assign w212 = pi086 & ~pi214;
assign w213 = (~pi214 & w211) | (~pi214 & w212) | (w211 & w212);
assign w214 = pi087 & ~pi215;
assign w215 = (~pi215 & w213) | (~pi215 & w214) | (w213 & w214);
assign w216 = ~pi089 & ~pi090;
assign w217 = ~pi091 & ~pi092;
assign w218 = w216 & w217;
assign w219 = ~pi088 & w218;
assign w220 = ~w215 & w219;
assign w221 = pi084 & ~pi212;
assign w222 = w129 & w221;
assign w223 = ~pi215 & w222;
assign w224 = w220 & ~w223;
assign w225 = ~pi215 & w130;
assign w226 = pi081 & ~pi209;
assign w227 = pi082 & ~pi210;
assign w228 = (~pi210 & w226) | (~pi210 & w227) | (w226 & w227);
assign w229 = ~pi083 & ~w228;
assign w230 = w225 & ~w229;
assign w231 = ~w210 & w230;
assign w232 = (~w210 & ~w224) | (~w210 & w231) | (~w224 & w231);
assign w233 = pi078 & ~pi206;
assign w234 = pi079 & ~pi207;
assign w235 = (~pi207 & w233) | (~pi207 & w234) | (w233 & w234);
assign w236 = ~pi080 & ~w235;
assign w237 = pi076 & ~pi204;
assign w238 = pi077 & ~pi207;
assign w239 = (~pi207 & w237) | (~pi207 & w238) | (w237 & w238);
assign w240 = w140 & w239;
assign w241 = w236 & ~w240;
assign w242 = pi073 & ~pi201;
assign w243 = pi074 & ~pi202;
assign w244 = (~pi202 & w242) | (~pi202 & w243) | (w242 & w243);
assign w245 = ~pi075 & ~w244;
assign w246 = w142 & ~w245;
assign w247 = w241 & ~w246;
assign w248 = w138 & ~w247;
assign w249 = ~w232 & ~w248;
assign w250 = w127 & ~w249;
assign w251 = ~w200 & ~w250;
assign w252 = ~w148 & w251;
assign w253 = ~pi125 & pi252;
assign w254 = ~pi126 & pi253;
assign w255 = (~pi126 & w253) | (~pi126 & w254) | (w253 & w254);
assign w256 = ~pi127 & pi254;
assign w257 = (~pi127 & w255) | (~pi127 & w256) | (w255 & w256);
assign w258 = w94 & w146;
assign w259 = w127 & w258;
assign w260 = ~pi252 & ~pi253;
assign w261 = ~pi254 & w260;
assign w262 = ~pi168 & ~pi169;
assign w263 = w261 & w262;
assign w264 = w76 & w263;
assign w265 = ~pi160 & ~pi161;
assign w266 = ~pi162 & w265;
assign w267 = ~pi163 & ~pi164;
assign w268 = ~pi165 & ~pi166;
assign w269 = w267 & w268;
assign w270 = ~pi167 & w269;
assign w271 = w266 & w270;
assign w272 = w264 & w271;
assign w273 = ~pi156 & ~pi157;
assign w274 = ~pi158 & ~pi159;
assign w275 = w273 & w274;
assign w276 = w272 & w275;
assign w277 = ~pi149 & ~pi150;
assign w278 = ~pi151 & w277;
assign w279 = ~pi153 & ~pi154;
assign w280 = ~pi155 & w279;
assign w281 = w278 & w280;
assign w282 = ~pi147 & ~pi148;
assign w283 = w281 & w282;
assign w284 = ~pi141 & ~pi142;
assign w285 = ~pi143 & ~pi144;
assign w286 = w284 & w285;
assign w287 = ~pi145 & ~pi146;
assign w288 = ~pi152 & w287;
assign w289 = w286 & w288;
assign w290 = w283 & w289;
assign w291 = w276 & w290;
assign w292 = w259 & w291;
assign w293 = pi011 & ~pi139;
assign w294 = pi012 & ~pi140;
assign w295 = (~pi140 & w293) | (~pi140 & w294) | (w293 & w294);
assign w296 = ~pi013 & ~w295;
assign w297 = ~pi136 & ~pi137;
assign w298 = ~pi135 & w297;
assign w299 = pi006 & ~pi134;
assign w300 = ~pi010 & ~w299;
assign w301 = (~pi010 & ~w298) | (~pi010 & w300) | (~w298 & w300);
assign w302 = pi007 & ~pi135;
assign w303 = pi008 & ~pi136;
assign w304 = (~pi136 & w302) | (~pi136 & w303) | (w302 & w303);
assign w305 = pi009 & ~pi137;
assign w306 = (~pi137 & w304) | (~pi137 & w305) | (w304 & w305);
assign w307 = w301 & ~w306;
assign w308 = ~pi138 & ~pi139;
assign w309 = ~pi140 & w308;
assign w310 = w296 & ~w309;
assign w311 = (w296 & w307) | (w296 & w310) | (w307 & w310);
assign w312 = w257 & w311;
assign w313 = (w257 & ~w292) | (w257 & w312) | (~w292 & w312);
assign w314 = w292 & ~w311;
assign w315 = pi125 & ~pi253;
assign w316 = pi126 & ~pi254;
assign w317 = (~pi254 & w315) | (~pi254 & w316) | (w315 & w316);
assign w318 = ~pi127 & ~w317;
assign w319 = pi113 & ~pi241;
assign w320 = pi114 & ~pi242;
assign w321 = (~pi242 & w319) | (~pi242 & w320) | (w319 & w320);
assign w322 = ~pi116 & pi243;
assign w323 = pi115 & ~pi243;
assign w324 = ~pi116 & ~w323;
assign w325 = (~w321 & w322) | (~w321 & w324) | (w322 & w324);
assign w326 = ~pi117 & pi244;
assign w327 = (~pi117 & w325) | (~pi117 & w326) | (w325 & w326);
assign w328 = pi110 & ~pi238;
assign w329 = pi111 & ~pi239;
assign w330 = (~pi239 & w328) | (~pi239 & w329) | (w328 & w329);
assign w331 = ~pi112 & ~w330;
assign w332 = w120 & ~w331;
assign w333 = w327 & ~w332;
assign w334 = ~w116 & w318;
assign w335 = (w318 & w333) | (w318 & w334) | (w333 & w334);
assign w336 = ~pi251 & w113;
assign w337 = pi118 & ~pi246;
assign w338 = ~pi119 & ~w337;
assign w339 = w336 & ~w338;
assign w340 = pi120 & ~pi248;
assign w341 = pi121 & ~pi249;
assign w342 = (~pi249 & w340) | (~pi249 & w341) | (w340 & w341);
assign w343 = ~pi123 & pi250;
assign w344 = pi122 & ~pi250;
assign w345 = ~pi123 & ~w344;
assign w346 = (~w342 & w343) | (~w342 & w345) | (w343 & w345);
assign w347 = ~pi251 & ~w346;
assign w348 = ~w339 & ~w347;
assign w349 = ~pi124 & w348;
assign w350 = w335 & w349;
assign w351 = ~w257 & ~w350;
assign w352 = ~w314 & ~w351;
assign w353 = (w252 & w313) | (w252 & w352) | (w313 & w352);
assign w354 = ~pi130 & ~pi131;
assign w355 = ~pi132 & w354;
assign w356 = pi001 & ~pi129;
assign w357 = ~pi002 & ~w356;
assign w358 = w355 & ~w357;
assign w359 = pi003 & ~pi131;
assign w360 = pi004 & ~pi132;
assign w361 = (~pi132 & w359) | (~pi132 & w360) | (w359 & w360);
assign w362 = ~pi005 & ~w361;
assign w363 = ~w358 & w362;
assign w364 = ~pi133 & ~pi134;
assign w365 = ~pi135 & ~pi136;
assign w366 = w364 & w365;
assign w367 = ~pi137 & ~pi255;
assign w368 = w366 & w367;
assign w369 = w309 & w368;
assign w370 = ~w363 & w369;
assign w371 = ~pi000 & ~w370;
assign w372 = (~pi000 & ~w292) | (~pi000 & w371) | (~w292 & w371);
assign w373 = pi255 & w372;
assign w374 = w259 & w276;
assign w375 = pi017 & ~pi145;
assign w376 = ~pi142 & ~pi143;
assign w377 = ~pi144 & ~pi145;
assign w378 = w376 & w377;
assign w379 = ~pi014 & ~w375;
assign w380 = (~w375 & ~w378) | (~w375 & w379) | (~w378 & w379);
assign w381 = pi015 & ~pi143;
assign w382 = pi016 & ~pi145;
assign w383 = (~pi145 & w381) | (~pi145 & w382) | (w381 & w382);
assign w384 = ~pi144 & w383;
assign w385 = w380 & ~w384;
assign w386 = ~pi018 & w385;
assign w387 = ~pi146 & w282;
assign w388 = w278 & w387;
assign w389 = ~pi027 & pi152;
assign w390 = (~pi027 & ~w388) | (~pi027 & w389) | (~w388 & w389);
assign w391 = (~pi027 & w386) | (~pi027 & w390) | (w386 & w390);
assign w392 = pi028 & w275;
assign w393 = pi031 & ~pi159;
assign w394 = ~pi032 & ~w393;
assign w395 = ~w392 & w394;
assign w396 = pi029 & ~pi157;
assign w397 = pi030 & ~pi159;
assign w398 = (~pi159 & w396) | (~pi159 & w397) | (w396 & w397);
assign w399 = ~pi158 & w398;
assign w400 = w266 & w399;
assign w401 = (w266 & ~w395) | (w266 & w400) | (~w395 & w400);
assign w402 = pi033 & ~pi161;
assign w403 = pi034 & ~pi162;
assign w404 = (~pi162 & w402) | (~pi162 & w403) | (w402 & w403);
assign w405 = ~pi035 & ~pi036;
assign w406 = ~w404 & w405;
assign w407 = ~w401 & w406;
assign w408 = w391 & w407;
assign w409 = pi019 & ~pi147;
assign w410 = pi020 & ~pi148;
assign w411 = (~pi148 & w409) | (~pi148 & w410) | (w409 & w410);
assign w412 = ~pi021 & ~w411;
assign w413 = w278 & ~w412;
assign w414 = ~pi025 & pi152;
assign w415 = w280 & ~w414;
assign w416 = pi022 & ~pi150;
assign w417 = pi023 & ~pi151;
assign w418 = (~pi151 & w416) | (~pi151 & w417) | (w416 & w417);
assign w419 = pi024 & ~pi152;
assign w420 = ~pi025 & ~w419;
assign w421 = (w414 & ~w418) | (w414 & w420) | (~w418 & w420);
assign w422 = w280 & ~w421;
assign w423 = (w413 & w415) | (w413 & w422) | (w415 & w422);
assign w424 = pi026 & ~pi154;
assign w425 = pi027 & ~pi155;
assign w426 = (~pi155 & w424) | (~pi155 & w425) | (w424 & w425);
assign w427 = ~pi028 & ~w426;
assign w428 = ~pi146 & ~pi152;
assign w429 = w282 & w428;
assign w430 = w281 & w429;
assign w431 = w427 & ~w430;
assign w432 = ~w423 & w431;
assign w433 = ~w423 & w427;
assign w434 = pi037 & ~pi165;
assign w435 = pi038 & ~pi166;
assign w436 = (~pi166 & w434) | (~pi166 & w435) | (w434 & w435);
assign w437 = ~pi040 & pi167;
assign w438 = pi039 & ~pi167;
assign w439 = ~pi040 & ~w438;
assign w440 = (~w436 & w437) | (~w436 & w439) | (w437 & w439);
assign w441 = w414 & w440;
assign w442 = w421 & w440;
assign w443 = (~w413 & w441) | (~w413 & w442) | (w441 & w442);
assign w444 = w430 & ~w443;
assign w445 = w433 & ~w444;
assign w446 = (w408 & w432) | (w408 & w445) | (w432 & w445);
assign w447 = w374 & ~w446;
assign w448 = w266 & ~w394;
assign w449 = (w266 & w399) | (w266 & w448) | (w399 & w448);
assign w450 = ~pi036 & pi163;
assign w451 = pi035 & ~pi163;
assign w452 = ~pi036 & ~w451;
assign w453 = (~w404 & w450) | (~w404 & w452) | (w450 & w452);
assign w454 = (~w449 & w450) | (~w449 & w453) | (w450 & w453);
assign w455 = w264 & ~w440;
assign w456 = ~pi164 & ~pi165;
assign w457 = ~pi166 & ~pi167;
assign w458 = w456 & w457;
assign w459 = w440 & ~w458;
assign w460 = w264 & ~w459;
assign w461 = (~w454 & w455) | (~w454 & w460) | (w455 & w460);
assign w462 = ~pi255 & w461;
assign w463 = w259 & w462;
assign w464 = ~pi255 & w264;
assign w465 = w259 & w464;
assign w466 = (w447 & w463) | (w447 & w465) | (w463 & w465);
assign w467 = w372 & ~w466;
assign w468 = (w353 & w373) | (w353 & w467) | (w373 & w467);
assign w469 = pi128 & ~w468;
assign w470 = ~pi001 & pi128;
assign w471 = pi000 & ~pi128;
assign w472 = ~pi001 & ~w471;
assign w473 = ~pi128 & ~w371;
assign w474 = ~pi001 & ~w473;
assign w475 = (~w292 & w472) | (~w292 & w474) | (w472 & w474);
assign w476 = (pi255 & w470) | (pi255 & w475) | (w470 & w475);
assign w477 = (~w466 & w470) | (~w466 & w475) | (w470 & w475);
assign w478 = (w353 & w476) | (w353 & w477) | (w476 & w477);
assign w479 = pi129 & ~w478;
assign w480 = ~pi000 & ~pi127;
assign w481 = ~pi000 & w256;
assign w482 = (w255 & w480) | (w255 & w481) | (w480 & w481);
assign w483 = w309 & ~w362;
assign w484 = w368 & w483;
assign w485 = w311 & ~w484;
assign w486 = ~pi000 & w257;
assign w487 = w485 & w486;
assign w488 = (~w292 & w482) | (~w292 & w487) | (w482 & w487);
assign w489 = ~pi000 & w485;
assign w490 = (~pi000 & ~w292) | (~pi000 & w489) | (~w292 & w489);
assign w491 = ~w351 & w490;
assign w492 = (w252 & w488) | (w252 & w491) | (w488 & w491);
assign w493 = ~pi000 & pi255;
assign w494 = ~pi128 & ~pi129;
assign w495 = ~w493 & w494;
assign w496 = w357 & ~w495;
assign w497 = w461 & w495;
assign w498 = w259 & w497;
assign w499 = w264 & w495;
assign w500 = w259 & w499;
assign w501 = (w447 & w498) | (w447 & w500) | (w498 & w500);
assign w502 = w357 & ~w501;
assign w503 = (w492 & w496) | (w492 & w502) | (w496 & w502);
assign w504 = pi130 & ~w503;
assign w505 = ~pi003 & pi130;
assign w506 = pi002 & ~pi130;
assign w507 = (~pi130 & w356) | (~pi130 & w506) | (w356 & w506);
assign w508 = ~pi003 & ~w507;
assign w509 = (~w495 & w505) | (~w495 & w508) | (w505 & w508);
assign w510 = (~w501 & w505) | (~w501 & w508) | (w505 & w508);
assign w511 = (w492 & w509) | (w492 & w510) | (w509 & w510);
assign w512 = pi131 & ~w511;
assign w513 = ~pi004 & pi131;
assign w514 = ~pi004 & ~w359;
assign w515 = (~w507 & w513) | (~w507 & w514) | (w513 & w514);
assign w516 = pi005 & w367;
assign w517 = w366 & w516;
assign w518 = w309 & w517;
assign w519 = w515 & ~w518;
assign w520 = (~w292 & w515) | (~w292 & w519) | (w515 & w519);
assign w521 = w493 & w520;
assign w522 = (~pi000 & ~w264) | (~pi000 & w493) | (~w264 & w493);
assign w523 = (~pi000 & ~w259) | (~pi000 & w522) | (~w259 & w522);
assign w524 = ~pi000 & ~w463;
assign w525 = (~w447 & w523) | (~w447 & w524) | (w523 & w524);
assign w526 = w520 & w525;
assign w527 = (w353 & w521) | (w353 & w526) | (w521 & w526);
assign w528 = w354 & w494;
assign w529 = pi132 & w528;
assign w530 = (pi132 & ~w515) | (pi132 & w529) | (~w515 & w529);
assign w531 = ~w527 & w530;
assign w532 = ~pi132 & ~w493;
assign w533 = w528 & w532;
assign w534 = ~pi132 & w528;
assign w535 = ~w525 & w534;
assign w536 = (~w353 & w533) | (~w353 & w535) | (w533 & w535);
assign w537 = w363 & ~w536;
assign w538 = pi133 & ~w537;
assign w539 = ~pi132 & ~pi133;
assign w540 = ~pi255 & w539;
assign w541 = w528 & w540;
assign w542 = ~w493 & w541;
assign w543 = ~w525 & w541;
assign w544 = (~w353 & w542) | (~w353 & w543) | (w542 & w543);
assign w545 = (~pi129 & w356) | (~pi129 & w471) | (w356 & w471);
assign w546 = ~pi002 & ~w545;
assign w547 = w355 & ~w546;
assign w548 = ~pi006 & pi133;
assign w549 = pi005 & ~pi133;
assign w550 = ~pi006 & ~w549;
assign w551 = (~w361 & w548) | (~w361 & w550) | (w548 & w550);
assign w552 = (~w547 & w548) | (~w547 & w551) | (w548 & w551);
assign w553 = ~w544 & w552;
assign w554 = pi134 & ~w553;
assign w555 = ~pi010 & ~w305;
assign w556 = w309 & ~w555;
assign w557 = w296 & ~w556;
assign w558 = w257 & w557;
assign w559 = (w257 & ~w292) | (w257 & w558) | (~w292 & w558);
assign w560 = w292 & ~w557;
assign w561 = ~w351 & ~w560;
assign w562 = (w252 & w559) | (w252 & w561) | (w559 & w561);
assign w563 = ~pi007 & pi134;
assign w564 = pi008 & w309;
assign w565 = w541 & w564;
assign w566 = w297 & w565;
assign w567 = ~pi134 & w566;
assign w568 = ~pi007 & ~w567;
assign w569 = (~pi007 & ~w292) | (~pi007 & w568) | (~w292 & w568);
assign w570 = ~w541 & w548;
assign w571 = ~w541 & w551;
assign w572 = (~w547 & w570) | (~w547 & w571) | (w570 & w571);
assign w573 = (w563 & w569) | (w563 & w572) | (w569 & w572);
assign w574 = w264 & w541;
assign w575 = w552 & ~w574;
assign w576 = (~w259 & w552) | (~w259 & w575) | (w552 & w575);
assign w577 = w461 & w541;
assign w578 = w259 & w577;
assign w579 = w552 & ~w578;
assign w580 = (~w447 & w576) | (~w447 & w579) | (w576 & w579);
assign w581 = (w563 & w569) | (w563 & w580) | (w569 & w580);
assign w582 = (w562 & w573) | (w562 & w581) | (w573 & w581);
assign w583 = pi135 & ~w582;
assign w584 = ~pi008 & pi135;
assign w585 = (~pi008 & w563) | (~pi008 & w584) | (w563 & w584);
assign w586 = ~pi134 & ~w548;
assign w587 = ~pi134 & ~w551;
assign w588 = (w547 & w586) | (w547 & w587) | (w586 & w587);
assign w589 = ~pi008 & ~w302;
assign w590 = (w584 & ~w588) | (w584 & w589) | (~w588 & w589);
assign w591 = (~w541 & w585) | (~w541 & w590) | (w585 & w590);
assign w592 = w259 & w574;
assign w593 = (w447 & w578) | (w447 & w592) | (w578 & w592);
assign w594 = (w585 & w590) | (w585 & ~w593) | (w590 & ~w593);
assign w595 = (w562 & w591) | (w562 & w594) | (w591 & w594);
assign w596 = pi136 & ~w595;
assign w597 = ~pi009 & ~w304;
assign w598 = ~pi134 & ~pi135;
assign w599 = ~pi136 & w598;
assign w600 = ~w572 & w599;
assign w601 = ~w580 & w599;
assign w602 = (~w562 & w600) | (~w562 & w601) | (w600 & w601);
assign w603 = w597 & ~w602;
assign w604 = pi137 & ~w603;
assign w605 = w368 & w534;
assign w606 = ~w493 & w605;
assign w607 = ~w525 & w605;
assign w608 = (~w353 & w606) | (~w353 & w607) | (w606 & w607);
assign w609 = ~pi137 & w366;
assign w610 = ~w362 & w609;
assign w611 = (w547 & w609) | (w547 & w610) | (w609 & w610);
assign w612 = w307 & ~w611;
assign w613 = ~w608 & w612;
assign w614 = pi138 & ~w613;
assign w615 = (~w252 & ~w257) | (~w252 & w351) | (~w257 & w351);
assign w616 = w259 & w264;
assign w617 = w259 & w461;
assign w618 = (w447 & w616) | (w447 & w617) | (w616 & w617);
assign w619 = ~pi013 & ~w294;
assign w620 = w307 & w619;
assign w621 = ~w611 & w620;
assign w622 = (~w292 & w612) | (~w292 & w621) | (w612 & w621);
assign w623 = ~w618 & w622;
assign w624 = ~w615 & w623;
assign w625 = w307 & ~w605;
assign w626 = ~w611 & w625;
assign w627 = ~pi011 & pi138;
assign w628 = (~pi011 & w626) | (~pi011 & w627) | (w626 & w627);
assign w629 = (~pi011 & w624) | (~pi011 & w628) | (w624 & w628);
assign w630 = pi139 & ~w629;
assign w631 = ~pi011 & ~pi012;
assign w632 = ~pi012 & pi138;
assign w633 = ~pi011 & w632;
assign w634 = (w626 & w631) | (w626 & w633) | (w631 & w633);
assign w635 = (w624 & w631) | (w624 & w634) | (w631 & w634);
assign w636 = ~pi012 & pi139;
assign w637 = pi140 & ~w636;
assign w638 = ~w635 & w637;
assign w639 = ~w307 & w309;
assign w640 = (w309 & w611) | (w309 & w639) | (w611 & w639);
assign w641 = w296 & ~w640;
assign w642 = (w310 & ~w605) | (w310 & w641) | (~w605 & w641);
assign w643 = w605 & w617;
assign w644 = w605 & w616;
assign w645 = (w447 & w643) | (w447 & w644) | (w643 & w644);
assign w646 = (w310 & w641) | (w310 & ~w645) | (w641 & ~w645);
assign w647 = (~w615 & w642) | (~w615 & w646) | (w642 & w646);
assign w648 = pi141 & ~w647;
assign w649 = ~pi140 & ~pi141;
assign w650 = w308 & w649;
assign w651 = w605 & w650;
assign w652 = w276 & w651;
assign w653 = w259 & w652;
assign w654 = pi144 & ~w375;
assign w655 = (~w375 & ~w383) | (~w375 & w654) | (~w383 & w654);
assign w656 = ~pi018 & w655;
assign w657 = w430 & ~w656;
assign w658 = w653 & w657;
assign w659 = ~w307 & w650;
assign w660 = (w611 & w650) | (w611 & w659) | (w650 & w659);
assign w661 = ~pi014 & pi141;
assign w662 = pi013 & ~pi141;
assign w663 = ~pi014 & ~w662;
assign w664 = (~w295 & w661) | (~w295 & w663) | (w661 & w663);
assign w665 = ~w650 & w664;
assign w666 = (~w605 & w664) | (~w605 & w665) | (w664 & w665);
assign w667 = ~w660 & w666;
assign w668 = ~w658 & w667;
assign w669 = w276 & ~w433;
assign w670 = w259 & w669;
assign w671 = ~w617 & ~w670;
assign w672 = ~w660 & w664;
assign w673 = ~w667 & ~w672;
assign w674 = (~w667 & ~w671) | (~w667 & w673) | (~w671 & w673);
assign w675 = ~w658 & ~w674;
assign w676 = (~w615 & w668) | (~w615 & w675) | (w668 & w675);
assign w677 = pi142 & ~w676;
assign w678 = pi016 & ~pi144;
assign w679 = (~pi145 & w375) | (~pi145 & w678) | (w375 & w678);
assign w680 = ~pi018 & ~w679;
assign w681 = w430 & ~w680;
assign w682 = w666 & ~w681;
assign w683 = ~w660 & w682;
assign w684 = (~w653 & w667) | (~w653 & w683) | (w667 & w683);
assign w685 = w653 & w681;
assign w686 = ~w674 & ~w685;
assign w687 = (~w615 & w684) | (~w615 & w686) | (w684 & w686);
assign w688 = ~pi015 & pi142;
assign w689 = (~pi015 & w687) | (~pi015 & w688) | (w687 & w688);
assign w690 = pi143 & ~w689;
assign w691 = ~pi016 & pi143;
assign w692 = (~pi016 & w688) | (~pi016 & w691) | (w688 & w691);
assign w693 = ~pi015 & ~pi016;
assign w694 = ~w692 & ~w693;
assign w695 = ~pi016 & ~pi018;
assign w696 = ~w679 & w695;
assign w697 = ~pi015 & w696;
assign w698 = (~w430 & w693) | (~w430 & w697) | (w693 & w697);
assign w699 = ~w692 & ~w698;
assign w700 = (w653 & w694) | (w653 & w699) | (w694 & w699);
assign w701 = (~w667 & ~w692) | (~w667 & w700) | (~w692 & w700);
assign w702 = (w674 & ~w692) | (w674 & w700) | (~w692 & w700);
assign w703 = (w615 & w701) | (w615 & w702) | (w701 & w702);
assign w704 = pi144 & w703;
assign w705 = ~pi017 & pi144;
assign w706 = (~pi017 & w692) | (~pi017 & w705) | (w692 & w705);
assign w707 = ~pi144 & w694;
assign w708 = ~pi017 & ~w707;
assign w709 = ~pi144 & w699;
assign w710 = ~pi017 & ~w709;
assign w711 = (~w653 & w708) | (~w653 & w710) | (w708 & w710);
assign w712 = (w667 & w706) | (w667 & w711) | (w706 & w711);
assign w713 = (~w674 & w706) | (~w674 & w711) | (w706 & w711);
assign w714 = (~w615 & w712) | (~w615 & w713) | (w712 & w713);
assign w715 = pi145 & ~w714;
assign w716 = w378 & ~w666;
assign w717 = (w378 & w660) | (w378 & w716) | (w660 & w716);
assign w718 = w656 & ~w717;
assign w719 = w378 & ~w667;
assign w720 = w378 & w673;
assign w721 = (~w671 & w719) | (~w671 & w720) | (w719 & w720);
assign w722 = w656 & ~w721;
assign w723 = (~w615 & w718) | (~w615 & w722) | (w718 & w722);
assign w724 = pi146 & ~w723;
assign w725 = ~pi146 & ~pi155;
assign w726 = w279 & w725;
assign w727 = ~pi152 & w726;
assign w728 = w275 & w727;
assign w729 = w272 & w728;
assign w730 = w259 & w729;
assign w731 = ~pi018 & ~w378;
assign w732 = w655 & w731;
assign w733 = ~pi146 & ~w732;
assign w734 = w378 & ~w664;
assign w735 = w656 & ~w734;
assign w736 = ~pi146 & ~w735;
assign w737 = (w660 & w733) | (w660 & w736) | (w733 & w736);
assign w738 = ~pi019 & ~w737;
assign w739 = ~pi145 & w286;
assign w740 = w309 & w739;
assign w741 = w605 & w740;
assign w742 = (~w413 & w414) | (~w413 & w421) | (w414 & w421);
assign w743 = w741 & ~w742;
assign w744 = ~pi019 & ~w743;
assign w745 = ~w737 & w744;
assign w746 = (~w730 & w738) | (~w730 & w745) | (w738 & w745);
assign w747 = pi025 & ~pi155;
assign w748 = w279 & w747;
assign w749 = w275 & w748;
assign w750 = (w275 & ~w427) | (w275 & w749) | (~w427 & w749);
assign w751 = w272 & w750;
assign w752 = w259 & w751;
assign w753 = ~w617 & ~w752;
assign w754 = w350 & w753;
assign w755 = w252 & w754;
assign w756 = pi127 & ~pi146;
assign w757 = ~pi146 & ~w256;
assign w758 = (~w255 & w756) | (~w255 & w757) | (w756 & w757);
assign w759 = w741 & w758;
assign w760 = w746 & ~w759;
assign w761 = (w746 & w755) | (w746 & w760) | (w755 & w760);
assign w762 = pi147 & ~w761;
assign w763 = ~pi147 & w759;
assign w764 = (~pi147 & ~w746) | (~pi147 & w763) | (~w746 & w763);
assign w765 = ~pi020 & ~w764;
assign w766 = ~pi147 & ~w746;
assign w767 = ~pi020 & ~w766;
assign w768 = (w755 & w765) | (w755 & w767) | (w765 & w767);
assign w769 = pi148 & ~w768;
assign w770 = w412 & ~w727;
assign w771 = w412 | w770;
assign w772 = (w412 & ~w741) | (w412 & w771) | (~w741 & w771);
assign w773 = (w412 & ~w741) | (w412 & w770) | (~w741 & w770);
assign w774 = pi024 & w282;
assign w775 = (w282 & w418) | (w282 & w774) | (w418 & w774);
assign w776 = w275 & w775;
assign w777 = w272 & w776;
assign w778 = (w412 & w773) | (w412 & ~w777) | (w773 & ~w777);
assign w779 = (~w259 & w772) | (~w259 & w778) | (w772 & w778);
assign w780 = w387 & ~w735;
assign w781 = w387 & ~w732;
assign w782 = (w660 & w780) | (w660 & w781) | (w780 & w781);
assign w783 = w779 & ~w782;
assign w784 = ~w257 & w387;
assign w785 = w741 & w784;
assign w786 = ~w782 & ~w785;
assign w787 = w779 & w786;
assign w788 = (w755 & w783) | (w755 & w787) | (w783 & w787);
assign w789 = pi149 & ~w788;
assign w790 = ~pi149 & w782;
assign w791 = (~pi149 & ~w779) | (~pi149 & w790) | (~w779 & w790);
assign w792 = ~pi022 & ~w791;
assign w793 = ~pi149 & ~w787;
assign w794 = ~pi022 & ~w793;
assign w795 = (w755 & w792) | (w755 & w794) | (w792 & w794);
assign w796 = pi150 & ~w795;
assign w797 = ~pi023 & pi150;
assign w798 = ~pi023 & ~w416;
assign w799 = (~w791 & w797) | (~w791 & w798) | (w797 & w798);
assign w800 = (~w793 & w797) | (~w793 & w798) | (w797 & w798);
assign w801 = (w755 & w799) | (w755 & w800) | (w799 & w800);
assign w802 = pi151 & ~w801;
assign w803 = ~pi024 & ~w418;
assign w804 = w278 & ~w783;
assign w805 = w803 & ~w804;
assign w806 = w278 & ~w787;
assign w807 = w803 & ~w806;
assign w808 = (w755 & w805) | (w755 & w807) | (w805 & w807);
assign w809 = pi152 & ~w808;
assign w810 = w275 & ~w427;
assign w811 = w272 & w810;
assign w812 = w259 & w811;
assign w813 = w257 & ~w461;
assign w814 = (w257 & ~w259) | (w257 & w813) | (~w259 & w813);
assign w815 = ~w812 & w814;
assign w816 = ~w351 & ~w617;
assign w817 = ~w812 & w816;
assign w818 = (w252 & w815) | (w252 & w817) | (w815 & w817);
assign w819 = ~pi152 & w388;
assign w820 = (~w660 & w732) | (~w660 & w735) | (w732 & w735);
assign w821 = w819 & ~w820;
assign w822 = w742 & ~w821;
assign w823 = ~w741 & w820;
assign w824 = w819 & ~w823;
assign w825 = w742 & ~w824;
assign w826 = (w818 & w822) | (w818 & w825) | (w822 & w825);
assign w827 = pi153 & ~w826;
assign w828 = ~w656 & w819;
assign w829 = ~pi153 & w828;
assign w830 = (~pi153 & ~w742) | (~pi153 & w829) | (~w742 & w829);
assign w831 = w278 & w282;
assign w832 = ~pi146 & w378;
assign w833 = w831 & w832;
assign w834 = ~pi152 & ~pi153;
assign w835 = ~w664 & w834;
assign w836 = w833 & w835;
assign w837 = ~pi026 & ~w836;
assign w838 = ~pi026 & ~w834;
assign w839 = (~pi026 & ~w833) | (~pi026 & w838) | (~w833 & w838);
assign w840 = (~w660 & w837) | (~w660 & w839) | (w837 & w839);
assign w841 = ~w830 & w840;
assign w842 = w388 & w834;
assign w843 = w741 & w842;
assign w844 = w841 & ~w843;
assign w845 = (w818 & w841) | (w818 & w844) | (w841 & w844);
assign w846 = pi154 & ~w845;
assign w847 = pi028 & w276;
assign w848 = w259 & w847;
assign w849 = w814 & ~w848;
assign w850 = w816 & ~w848;
assign w851 = (w252 & w849) | (w252 & w850) | (w849 & w850);
assign w852 = ~pi154 & ~w841;
assign w853 = ~pi027 & ~w852;
assign w854 = ~pi154 & ~w844;
assign w855 = ~pi027 & ~w854;
assign w856 = (w851 & w853) | (w851 & w855) | (w853 & w855);
assign w857 = pi155 & ~w856;
assign w858 = w430 & w741;
assign w859 = ~w816 & w858;
assign w860 = ~w814 & w858;
assign w861 = (~w252 & w859) | (~w252 & w860) | (w859 & w860);
assign w862 = ~pi027 & pi154;
assign w863 = ~pi028 & pi155;
assign w864 = (~pi028 & w862) | (~pi028 & w863) | (w862 & w863);
assign w865 = ~pi027 & ~pi028;
assign w866 = w840 & w865;
assign w867 = ~pi153 & ~w864;
assign w868 = ~w414 & ~w864;
assign w869 = ~w421 & ~w864;
assign w870 = (w413 & w868) | (w413 & w869) | (w868 & w869);
assign w871 = (w829 & w867) | (w829 & w870) | (w867 & w870);
assign w872 = (~w864 & ~w866) | (~w864 & w871) | (~w866 & w871);
assign w873 = ~w861 & ~w872;
assign w874 = pi156 & ~w873;
assign w875 = ~pi029 & pi156;
assign w876 = ~pi156 & ~w864;
assign w877 = ~pi029 & ~w876;
assign w878 = ~pi156 & w867;
assign w879 = ~pi156 & w870;
assign w880 = (w829 & w878) | (w829 & w879) | (w878 & w879);
assign w881 = ~pi029 & ~w880;
assign w882 = (w866 & w877) | (w866 & w881) | (w877 & w881);
assign w883 = (~w861 & w875) | (~w861 & w882) | (w875 & w882);
assign w884 = pi157 & ~w883;
assign w885 = ~pi030 & pi157;
assign w886 = (~pi030 & w875) | (~pi030 & w885) | (w875 & w885);
assign w887 = (~pi030 & w882) | (~pi030 & w885) | (w882 & w885);
assign w888 = (~w861 & w886) | (~w861 & w887) | (w886 & w887);
assign w889 = pi158 & ~w888;
assign w890 = pi030 & ~pi158;
assign w891 = (~pi158 & w396) | (~pi158 & w890) | (w396 & w890);
assign w892 = ~pi031 & ~w891;
assign w893 = ~pi157 & ~pi158;
assign w894 = ~pi156 & w893;
assign w895 = w892 & ~w894;
assign w896 = (~w866 & w876) | (~w866 & w880) | (w876 & w880);
assign w897 = w893 & w896;
assign w898 = w892 & ~w897;
assign w899 = (~w861 & w895) | (~w861 & w898) | (w895 & w898);
assign w900 = pi159 & ~w899;
assign w901 = w275 & w429;
assign w902 = w281 & w901;
assign w903 = w741 & w902;
assign w904 = ~w814 & w903;
assign w905 = ~w816 & w903;
assign w906 = (~w252 & w904) | (~w252 & w905) | (w904 & w905);
assign w907 = w394 & w864;
assign w908 = ~w399 & w907;
assign w909 = w394 & ~w399;
assign w910 = (~w275 & w908) | (~w275 & w909) | (w908 & w909);
assign w911 = ~pi153 & w275;
assign w912 = (w908 & w909) | (w908 & ~w911) | (w909 & ~w911);
assign w913 = w275 & ~w414;
assign w914 = w275 & ~w421;
assign w915 = (w413 & w913) | (w413 & w914) | (w913 & w914);
assign w916 = (w908 & w909) | (w908 & ~w915) | (w909 & ~w915);
assign w917 = (~w829 & w912) | (~w829 & w916) | (w912 & w916);
assign w918 = (w866 & w910) | (w866 & w917) | (w910 & w917);
assign w919 = ~w906 & w918;
assign w920 = pi160 & ~w919;
assign w921 = ~pi035 & ~w403;
assign w922 = w270 & ~w921;
assign w923 = pi036 & w458;
assign w924 = w440 & ~w923;
assign w925 = ~w922 & w924;
assign w926 = w264 & ~w925;
assign w927 = w259 & w926;
assign w928 = ~w351 & ~w927;
assign w929 = w903 & ~w928;
assign w930 = ~w257 & w902;
assign w931 = w741 & w930;
assign w932 = w257 & ~w264;
assign w933 = (w257 & w925) | (w257 & w932) | (w925 & w932);
assign w934 = w903 & ~w933;
assign w935 = (w259 & w931) | (w259 & w934) | (w931 & w934);
assign w936 = (~w252 & w929) | (~w252 & w935) | (w929 & w935);
assign w937 = ~pi033 & pi160;
assign w938 = ~pi160 & ~w910;
assign w939 = ~pi160 & ~w917;
assign w940 = (~w866 & w938) | (~w866 & w939) | (w938 & w939);
assign w941 = ~pi033 & ~w940;
assign w942 = (~w936 & w937) | (~w936 & w941) | (w937 & w941);
assign w943 = pi161 & ~w942;
assign w944 = ~pi034 & pi161;
assign w945 = ~pi034 & ~w402;
assign w946 = (pi160 & w944) | (pi160 & w945) | (w944 & w945);
assign w947 = (~w940 & w944) | (~w940 & w945) | (w944 & w945);
assign w948 = (~w936 & w946) | (~w936 & w947) | (w946 & w947);
assign w949 = pi162 & ~w948;
assign w950 = ~pi035 & ~w404;
assign w951 = ~w266 & w950;
assign w952 = w266 & ~w918;
assign w953 = w950 & ~w952;
assign w954 = (~w936 & w951) | (~w936 & w953) | (w951 & w953);
assign w955 = pi163 & ~w954;
assign w956 = w266 & w429;
assign w957 = w281 & w956;
assign w958 = ~pi163 & w275;
assign w959 = w957 & w958;
assign w960 = w741 & w959;
assign w961 = w259 & w455;
assign w962 = ~w351 & ~w961;
assign w963 = w960 & ~w962;
assign w964 = w257 & ~w961;
assign w965 = w960 & ~w964;
assign w966 = (~w252 & w963) | (~w252 & w965) | (w963 & w965);
assign w967 = ~w449 & w950;
assign w968 = w266 & w275;
assign w969 = ~pi163 & ~w864;
assign w970 = w968 & w969;
assign w971 = ~pi036 & ~w970;
assign w972 = (w450 & w967) | (w450 & w971) | (w967 & w971);
assign w973 = (~pi163 & ~w967) | (~pi163 & w970) | (~w967 & w970);
assign w974 = w450 & w865;
assign w975 = pi163 & w865;
assign w976 = ~w451 & w865;
assign w977 = (~w404 & w975) | (~w404 & w976) | (w975 & w976);
assign w978 = ~pi036 & w977;
assign w979 = (~w449 & w974) | (~w449 & w978) | (w974 & w978);
assign w980 = (~pi036 & ~w973) | (~pi036 & w979) | (~w973 & w979);
assign w981 = (w841 & w972) | (w841 & w980) | (w972 & w980);
assign w982 = ~w966 & w981;
assign w983 = pi164 & ~w982;
assign w984 = w264 & ~w439;
assign w985 = w259 & w984;
assign w986 = ~w351 & ~w985;
assign w987 = w960 & ~w986;
assign w988 = ~w257 & w960;
assign w989 = w257 & w439;
assign w990 = (w257 & ~w264) | (w257 & w989) | (~w264 & w989);
assign w991 = w960 & ~w990;
assign w992 = (w259 & w988) | (w259 & w991) | (w988 & w991);
assign w993 = (~w252 & w987) | (~w252 & w992) | (w987 & w992);
assign w994 = w264 & w960;
assign w995 = w259 & w994;
assign w996 = ~pi167 & w435;
assign w997 = w995 & w996;
assign w998 = w981 & ~w997;
assign w999 = ~pi164 & ~w998;
assign w1000 = (~pi164 & w993) | (~pi164 & w999) | (w993 & w999);
assign w1001 = ~pi037 & ~w1000;
assign w1002 = pi165 & ~w1001;
assign w1003 = ~pi038 & ~w434;
assign w1004 = ~w456 & w1003;
assign w1005 = w456 & ~w972;
assign w1006 = w456 & ~w980;
assign w1007 = (~w841 & w1005) | (~w841 & w1006) | (w1005 & w1006);
assign w1008 = w1003 & ~w1007;
assign w1009 = (~w993 & w1004) | (~w993 & w1008) | (w1004 & w1008);
assign w1010 = pi166 & ~w1009;
assign w1011 = ~pi039 & pi166;
assign w1012 = (~pi039 & w1004) | (~pi039 & w1011) | (w1004 & w1011);
assign w1013 = (~pi039 & w1008) | (~pi039 & w1011) | (w1008 & w1011);
assign w1014 = (~w993 & w1012) | (~w993 & w1013) | (w1012 & w1013);
assign w1015 = pi167 & ~w1014;
assign w1016 = w408 & w443;
assign w1017 = ~pi026 & pi153;
assign w1018 = (~pi027 & w862) | (~pi027 & w1017) | (w862 & w1017);
assign w1019 = ~pi155 & ~w1018;
assign w1020 = w968 & w1019;
assign w1021 = w406 & ~w1020;
assign w1022 = ~w401 & w1021;
assign w1023 = ~w450 & w458;
assign w1024 = w440 & ~w1023;
assign w1025 = (w440 & w1022) | (w440 & w1024) | (w1022 & w1024);
assign w1026 = ~w840 & ~w1025;
assign w1027 = (~w1016 & ~w1025) | (~w1016 & w1026) | (~w1025 & w1026);
assign w1028 = w270 & w968;
assign w1029 = w430 & w1028;
assign w1030 = w741 & w1029;
assign w1031 = ~w257 & w1030;
assign w1032 = ~w1027 & ~w1031;
assign w1033 = ~w350 & w1031;
assign w1034 = ~w1027 & ~w1033;
assign w1035 = (w252 & w1032) | (w252 & w1034) | (w1032 & w1034);
assign w1036 = pi168 & ~w1035;
assign w1037 = ~pi041 & pi168;
assign w1038 = (~pi041 & w1035) | (~pi041 & w1037) | (w1035 & w1037);
assign w1039 = pi169 & ~w1038;
assign w1040 = ~w69 & w147;
assign w1041 = ~w250 & ~w1040;
assign w1042 = ~w200 & w350;
assign w1043 = w1041 & w1042;
assign w1044 = w261 & w1030;
assign w1045 = w259 & w1044;
assign w1046 = ~pi041 & ~pi042;
assign w1047 = ~w1031 & w1046;
assign w1048 = ~w88 & w1046;
assign w1049 = w82 & w1048;
assign w1050 = ~w1031 & w1049;
assign w1051 = (~w1045 & w1047) | (~w1045 & w1050) | (w1047 & w1050);
assign w1052 = ~w1027 & w1051;
assign w1053 = (~w1045 & w1046) | (~w1045 & w1049) | (w1046 & w1049);
assign w1054 = ~w1027 & w1053;
assign w1055 = (w1043 & w1052) | (w1043 & w1054) | (w1052 & w1054);
assign w1056 = pi170 & ~w1055;
assign w1057 = ~pi042 & pi169;
assign w1058 = (~pi042 & w1037) | (~pi042 & w1057) | (w1037 & w1057);
assign w1059 = w1056 & ~w1058;
assign w1060 = (w1043 & w1051) | (w1043 & w1053) | (w1051 & w1053);
assign w1061 = ~pi170 & pi171;
assign w1062 = ~w1058 & w1061;
assign w1063 = w1027 & ~w1058;
assign w1064 = w1061 & w1063;
assign w1065 = (~w1060 & w1062) | (~w1060 & w1064) | (w1062 & w1064);
assign w1066 = pi043 & pi171;
assign w1067 = ~w1065 & ~w1066;
assign w1068 = ~w1027 & w1046;
assign w1069 = ~pi127 & w1046;
assign w1070 = w256 & w1046;
assign w1071 = (w255 & w1069) | (w255 & w1070) | (w1069 & w1070);
assign w1072 = (~w1030 & w1046) | (~w1030 & w1071) | (w1046 & w1071);
assign w1073 = ~w1027 & w1072;
assign w1074 = (w1043 & w1068) | (w1043 & w1073) | (w1068 & w1073);
assign w1075 = w72 & w262;
assign w1076 = ~pi175 & w1075;
assign w1077 = ~pi047 & ~w86;
assign w1078 = w1076 & ~w1077;
assign w1079 = w1045 & w1078;
assign w1080 = ~pi043 & pi170;
assign w1081 = ~pi171 & ~w1080;
assign w1082 = (w78 & ~w1058) | (w78 & w1081) | (~w1058 & w1081);
assign w1083 = ~pi044 & ~w1082;
assign w1084 = ~w1079 & w1083;
assign w1085 = pi048 & w259;
assign w1086 = ~pi043 & ~pi044;
assign w1087 = pi044 & ~w1086;
assign w1088 = (w1082 & ~w1086) | (w1082 & w1087) | (~w1086 & w1087);
assign w1089 = ~pi044 & pi254;
assign w1090 = (~pi044 & ~w260) | (~pi044 & w1089) | (~w260 & w1089);
assign w1091 = ~pi043 & w1090;
assign w1092 = ~w1083 & ~w1091;
assign w1093 = (w1030 & w1088) | (w1030 & w1092) | (w1088 & w1092);
assign w1094 = (w1085 & w1088) | (w1085 & w1093) | (w1088 & w1093);
assign w1095 = ~w1079 & ~w1094;
assign w1096 = (w1074 & w1084) | (w1074 & w1095) | (w1084 & w1095);
assign w1097 = pi172 & ~w1096;
assign w1098 = ~pi045 & pi172;
assign w1099 = ~pi172 & w1078;
assign w1100 = ~pi045 & ~w1099;
assign w1101 = (~pi045 & ~w1045) | (~pi045 & w1100) | (~w1045 & w1100);
assign w1102 = (w1083 & w1098) | (w1083 & w1101) | (w1098 & w1101);
assign w1103 = (~w1094 & w1098) | (~w1094 & w1101) | (w1098 & w1101);
assign w1104 = (w1074 & w1102) | (w1074 & w1103) | (w1102 & w1103);
assign w1105 = pi173 & ~w1104;
assign w1106 = ~pi045 & ~pi046;
assign w1107 = w87 & w1075;
assign w1108 = w1083 & ~w1107;
assign w1109 = (~w1045 & w1083) | (~w1045 & w1108) | (w1083 & w1108);
assign w1110 = w1106 & w1109;
assign w1111 = w1045 & w1107;
assign w1112 = ~w1094 & ~w1111;
assign w1113 = w1106 & w1112;
assign w1114 = (w1074 & w1110) | (w1074 & w1113) | (w1110 & w1113);
assign w1115 = ~pi046 & pi173;
assign w1116 = (~pi046 & w1098) | (~pi046 & w1115) | (w1098 & w1115);
assign w1117 = pi174 & ~w1116;
assign w1118 = ~w1114 & w1117;
assign w1119 = ~pi173 & ~pi174;
assign w1120 = ~pi172 & w1119;
assign w1121 = pi044 & ~pi172;
assign w1122 = w1119 & w1121;
assign w1123 = (w1082 & w1120) | (w1082 & w1122) | (w1120 & w1122);
assign w1124 = w1077 & ~w1123;
assign w1125 = ~pi172 & w1088;
assign w1126 = ~pi172 & w1093;
assign w1127 = (w1085 & w1125) | (w1085 & w1126) | (w1125 & w1126);
assign w1128 = w1119 & w1127;
assign w1129 = w1077 & ~w1128;
assign w1130 = (w1074 & w1124) | (w1074 & w1129) | (w1124 & w1129);
assign w1131 = pi175 & ~w1130;
assign w1132 = (~w1027 & w1032) | (~w1027 & w1043) | (w1032 & w1043);
assign w1133 = w75 & w262;
assign w1134 = w74 & w1133;
assign w1135 = w89 & ~w1134;
assign w1136 = (w89 & w1132) | (w89 & w1135) | (w1132 & w1135);
assign w1137 = pi176 & ~w1136;
assign w1138 = w272 & w902;
assign w1139 = w741 & w1138;
assign w1140 = w147 & w1139;
assign w1141 = (~pi179 & w1) | (~pi179 & w4) | (w1 & w4);
assign w1142 = ~pi052 & ~w1141;
assign w1143 = w9 & ~w1142;
assign w1144 = w17 & ~w1143;
assign w1145 = w33 & ~w1144;
assign w1146 = w1140 & w1145;
assign w1147 = ~w88 & w440;
assign w1148 = w83 & w1147;
assign w1149 = w979 & w1148;
assign w1150 = w841 & w1149;
assign w1151 = w89 & ~w973;
assign w1152 = ~pi036 & w440;
assign w1153 = w1151 & w1152;
assign w1154 = ~w459 & w1134;
assign w1155 = w89 & ~w1154;
assign w1156 = ~w1153 & ~w1155;
assign w1157 = ~w1150 & w1156;
assign w1158 = ~w1146 & ~w1157;
assign w1159 = ~w68 & w147;
assign w1160 = ~w200 & ~w1159;
assign w1161 = ~w250 & w350;
assign w1162 = w1160 & w1161;
assign w1163 = w1028 & w1134;
assign w1164 = w430 & w1163;
assign w1165 = ~w257 & w741;
assign w1166 = w1164 & w1165;
assign w1167 = ~w1162 & w1166;
assign w1168 = w1158 & ~w1167;
assign w1169 = ~pi049 & pi176;
assign w1170 = (~pi049 & w1168) | (~pi049 & w1169) | (w1168 & w1169);
assign w1171 = pi177 & ~w1170;
assign w1172 = ~pi049 & ~pi050;
assign w1173 = pi176 & w1172;
assign w1174 = (w1168 & w1172) | (w1168 & w1173) | (w1172 & w1173);
assign w1175 = ~pi050 & pi177;
assign w1176 = pi178 & ~w1175;
assign w1177 = ~w1174 & w1176;
assign w1178 = ~pi051 & ~w2;
assign w1179 = ~pi178 & w90;
assign w1180 = w1178 & ~w1179;
assign w1181 = (w1168 & w1178) | (w1168 & w1180) | (w1178 & w1180);
assign w1182 = pi179 & ~w1181;
assign w1183 = w6 & ~w1179;
assign w1184 = (w6 & w1168) | (w6 & w1183) | (w1168 & w1183);
assign w1185 = pi180 & ~w3;
assign w1186 = ~w1184 & w1185;
assign w1187 = pi054 & w8;
assign w1188 = w16 & ~w1187;
assign w1189 = w33 & ~w1188;
assign w1190 = w1140 & w1189;
assign w1191 = ~w1157 & ~w1190;
assign w1192 = ~w1167 & w1191;
assign w1193 = ~pi053 & pi180;
assign w1194 = (~pi053 & w6) | (~pi053 & w1193) | (w6 & w1193);
assign w1195 = ~pi180 & w92;
assign w1196 = (~pi180 & ~w6) | (~pi180 & w1195) | (~w6 & w1195);
assign w1197 = ~pi053 & ~w1196;
assign w1198 = (w1192 & w1194) | (w1192 & w1197) | (w1194 & w1197);
assign w1199 = pi181 & ~w1198;
assign w1200 = ~pi054 & ~w11;
assign w1201 = w6 & w1200;
assign w1202 = ~w92 & w1200;
assign w1203 = w6 & w1202;
assign w1204 = (w1192 & w1201) | (w1192 & w1203) | (w1201 & w1203);
assign w1205 = pi182 & w7;
assign w1206 = (pi182 & ~w1200) | (pi182 & w1205) | (~w1200 & w1205);
assign w1207 = ~w1204 & w1206;
assign w1208 = w92 & w1157;
assign w1209 = (w92 & w1167) | (w92 & w1208) | (w1167 & w1208);
assign w1210 = ~pi054 & ~pi055;
assign w1211 = ~w11 & w1210;
assign w1212 = w6 & w1211;
assign w1213 = pi056 & w92;
assign w1214 = w1200 & ~w1213;
assign w1215 = (~w33 & w1200) | (~w33 & w1214) | (w1200 & w1214);
assign w1216 = ~pi055 & w6;
assign w1217 = w1215 & w1216;
assign w1218 = (~w1140 & w1212) | (~w1140 & w1217) | (w1212 & w1217);
assign w1219 = ~w1209 & w1218;
assign w1220 = ~pi182 & w7;
assign w1221 = (~pi182 & ~w1200) | (~pi182 & w1220) | (~w1200 & w1220);
assign w1222 = pi055 & pi183;
assign w1223 = (pi183 & w1221) | (pi183 & w1222) | (w1221 & w1222);
assign w1224 = ~w1219 & w1223;
assign w1225 = w116 & ~w333;
assign w1226 = w349 & ~w1225;
assign w1227 = w318 & w1226;
assign w1228 = w1166 & ~w1227;
assign w1229 = (~w251 & w1166) | (~w251 & w1228) | (w1166 & w1228);
assign w1230 = ~w1157 & ~w1229;
assign w1231 = w147 & w1138;
assign w1232 = w93 & w741;
assign w1233 = w18 & w67;
assign w1234 = (w18 & ~w1232) | (w18 & w1233) | (~w1232 & w1233);
assign w1235 = (w18 & ~w1231) | (w18 & w1234) | (~w1231 & w1234);
assign w1236 = w25 & w93;
assign w1237 = w741 & w1236;
assign w1238 = ~w68 & w1237;
assign w1239 = w1231 & w1238;
assign w1240 = w1235 & ~w1239;
assign w1241 = ~w93 & ~w1238;
assign w1242 = (~w93 & ~w1231) | (~w93 & w1241) | (~w1231 & w1241);
assign w1243 = w1235 & w1242;
assign w1244 = (w1230 & w1240) | (w1230 & w1243) | (w1240 & w1243);
assign w1245 = pi184 & ~w1244;
assign w1246 = ~pi057 & pi184;
assign w1247 = (~pi057 & w1243) | (~pi057 & w1246) | (w1243 & w1246);
assign w1248 = (~pi057 & w1240) | (~pi057 & w1246) | (w1240 & w1246);
assign w1249 = (w1230 & w1247) | (w1230 & w1248) | (w1247 & w1248);
assign w1250 = pi185 & ~w1249;
assign w1251 = ~pi058 & pi185;
assign w1252 = (~pi058 & w1246) | (~pi058 & w1251) | (w1246 & w1251);
assign w1253 = ~pi058 & ~w35;
assign w1254 = (w1243 & w1252) | (w1243 & w1253) | (w1252 & w1253);
assign w1255 = (w1240 & w1252) | (w1240 & w1253) | (w1252 & w1253);
assign w1256 = (w1230 & w1254) | (w1230 & w1255) | (w1254 & w1255);
assign w1257 = pi186 & ~w1256;
assign w1258 = ~pi059 & ~w37;
assign w1259 = ~pi184 & ~w1243;
assign w1260 = ~pi184 & ~w1240;
assign w1261 = (~w1230 & w1259) | (~w1230 & w1260) | (w1259 & w1260);
assign w1262 = ~pi185 & ~pi186;
assign w1263 = ~pi059 & ~w1262;
assign w1264 = ~w37 & w1263;
assign w1265 = (w1258 & ~w1261) | (w1258 & w1264) | (~w1261 & w1264);
assign w1266 = pi187 & ~w1265;
assign w1267 = w1138 & w1237;
assign w1268 = w147 & w1267;
assign w1269 = ~w49 & w1268;
assign w1270 = w1235 & ~w1269;
assign w1271 = w31 & ~w1270;
assign w1272 = w18 & ~w93;
assign w1273 = ~w93 & w1234;
assign w1274 = (~w1231 & w1272) | (~w1231 & w1273) | (w1272 & w1273);
assign w1275 = ~w1269 & w1274;
assign w1276 = w31 & ~w1275;
assign w1277 = (~w1230 & w1271) | (~w1230 & w1276) | (w1271 & w1276);
assign w1278 = w41 & ~w1277;
assign w1279 = pi188 & ~w1278;
assign w1280 = w31 & w93;
assign w1281 = (~w18 & w31) | (~w18 & w1280) | (w31 & w1280);
assign w1282 = w25 & ~w48;
assign w1283 = w67 & ~w1282;
assign w1284 = w18 & w1283;
assign w1285 = (w18 & ~w1140) | (w18 & w1284) | (~w1140 & w1284);
assign w1286 = ~w1157 & w1285;
assign w1287 = w1229 & w1281;
assign w1288 = (w1281 & ~w1286) | (w1281 & w1287) | (~w1286 & w1287);
assign w1289 = ~pi061 & pi188;
assign w1290 = (~pi061 & w41) | (~pi061 & w1289) | (w41 & w1289);
assign w1291 = pi062 & w27;
assign w1292 = w31 & w1291;
assign w1293 = w41 & ~w1292;
assign w1294 = (~pi061 & w1289) | (~pi061 & w1293) | (w1289 & w1293);
assign w1295 = (~w1268 & w1290) | (~w1268 & w1294) | (w1290 & w1294);
assign w1296 = (~w1288 & w1289) | (~w1288 & w1295) | (w1289 & w1295);
assign w1297 = pi189 & ~w1296;
assign w1298 = ~pi062 & pi189;
assign w1299 = (~pi062 & w1289) | (~pi062 & w1298) | (w1289 & w1298);
assign w1300 = ~pi061 & ~pi062;
assign w1301 = ~w31 & w1300;
assign w1302 = w41 & w1301;
assign w1303 = w41 & w1300;
assign w1304 = ~w1280 & w1303;
assign w1305 = (w18 & w1302) | (w18 & w1304) | (w1302 & w1304);
assign w1306 = ~w1299 & ~w1305;
assign w1307 = ~w18 & w1281;
assign w1308 = w1281 & ~w1284;
assign w1309 = (w1140 & w1307) | (w1140 & w1308) | (w1307 & w1308);
assign w1310 = w1303 & ~w1309;
assign w1311 = ~w1299 & ~w1310;
assign w1312 = (~w1230 & w1306) | (~w1230 & w1311) | (w1306 & w1311);
assign w1313 = pi190 & w1312;
assign w1314 = ~pi063 & pi190;
assign w1315 = (~pi063 & w1299) | (~pi063 & w1314) | (w1299 & w1314);
assign w1316 = (~pi063 & w1305) | (~pi063 & w1315) | (w1305 & w1315);
assign w1317 = (~pi063 & w1310) | (~pi063 & w1315) | (w1310 & w1315);
assign w1318 = (w1230 & w1316) | (w1230 & w1317) | (w1316 & w1317);
assign w1319 = pi191 & ~w1318;
assign w1320 = ~w28 & w49;
assign w1321 = ~w42 & w49;
assign w1322 = ~w18 & w31;
assign w1323 = w31 & ~w1234;
assign w1324 = (w1231 & w1322) | (w1231 & w1323) | (w1322 & w1323);
assign w1325 = (w1320 & w1321) | (w1320 & ~w1324) | (w1321 & ~w1324);
assign w1326 = w31 & ~w1274;
assign w1327 = (w1320 & w1321) | (w1320 & ~w1326) | (w1321 & ~w1326);
assign w1328 = (w1230 & w1325) | (w1230 & w1327) | (w1325 & w1327);
assign w1329 = pi192 & ~w1328;
assign w1330 = w41 & w49;
assign w1331 = w18 & w1330;
assign w1332 = ~w1157 & w1331;
assign w1333 = (~pi195 & w53) | (~pi195 & w56) | (w53 & w56);
assign w1334 = ~pi068 & ~w1333;
assign w1335 = w24 & ~w1334;
assign w1336 = w66 & ~w1335;
assign w1337 = w1140 & ~w1336;
assign w1338 = ~w1229 & ~w1337;
assign w1339 = w1332 & w1338;
assign w1340 = ~w31 & w41;
assign w1341 = w41 & ~w1280;
assign w1342 = (w18 & w1340) | (w18 & w1341) | (w1340 & w1341);
assign w1343 = ~pi192 & w28;
assign w1344 = (~pi192 & ~w49) | (~pi192 & w1343) | (~w49 & w1343);
assign w1345 = ~pi065 & ~w1344;
assign w1346 = ~pi065 & pi192;
assign w1347 = (~pi065 & w49) | (~pi065 & w1346) | (w49 & w1346);
assign w1348 = (w1342 & w1345) | (w1342 & w1347) | (w1345 & w1347);
assign w1349 = (~pi065 & w1339) | (~pi065 & w1348) | (w1339 & w1348);
assign w1350 = pi193 & ~w1349;
assign w1351 = ~pi066 & ~w52;
assign w1352 = ~pi066 & pi193;
assign w1353 = (~pi066 & w1346) | (~pi066 & w1352) | (w1346 & w1352);
assign w1354 = (w49 & w1351) | (w49 & w1353) | (w1351 & w1353);
assign w1355 = (~w1344 & w1351) | (~w1344 & w1352) | (w1351 & w1352);
assign w1356 = (w1342 & w1354) | (w1342 & w1355) | (w1354 & w1355);
assign w1357 = (w1339 & w1351) | (w1339 & w1356) | (w1351 & w1356);
assign w1358 = pi194 & ~w1357;
assign w1359 = ~pi067 & ~w54;
assign w1360 = pi065 & ~pi194;
assign w1361 = ~pi193 & w1360;
assign w1362 = w1359 & ~w1361;
assign w1363 = ~pi067 & pi193;
assign w1364 = ~w54 & w1363;
assign w1365 = ~pi194 & ~w1346;
assign w1366 = (~w49 & w1360) | (~w49 & w1365) | (w1360 & w1365);
assign w1367 = (w1359 & w1364) | (w1359 & ~w1366) | (w1364 & ~w1366);
assign w1368 = (pi194 & w1359) | (pi194 & w1364) | (w1359 & w1364);
assign w1369 = (w1359 & ~w1360) | (w1359 & w1364) | (~w1360 & w1364);
assign w1370 = (~w1344 & w1368) | (~w1344 & w1369) | (w1368 & w1369);
assign w1371 = (w1342 & w1367) | (w1342 & w1370) | (w1367 & w1370);
assign w1372 = (w1339 & w1362) | (w1339 & w1371) | (w1362 & w1371);
assign w1373 = pi195 & ~w1372;
assign w1374 = w21 & ~w49;
assign w1375 = w58 & ~w1374;
assign w1376 = ~pi193 & w20;
assign w1377 = w58 & ~w1376;
assign w1378 = (w58 & ~w1344) | (w58 & w1377) | (~w1344 & w1377);
assign w1379 = (w1342 & w1375) | (w1342 & w1378) | (w1375 & w1378);
assign w1380 = w58 & w66;
assign w1381 = w1330 & w1380;
assign w1382 = w18 & w1381;
assign w1383 = ~w1379 & ~w1382;
assign w1384 = w58 & w1330;
assign w1385 = w18 & w1384;
assign w1386 = ~w1379 & ~w1385;
assign w1387 = (w1140 & w1383) | (w1140 & w1386) | (w1383 & w1386);
assign w1388 = (~w1230 & ~w1379) | (~w1230 & w1387) | (~w1379 & w1387);
assign w1389 = pi196 & w1388;
assign w1390 = ~pi196 & ~w1379;
assign w1391 = ~pi069 & ~w1390;
assign w1392 = ~pi196 & w1387;
assign w1393 = ~pi069 & ~w1392;
assign w1394 = (w1230 & w1391) | (w1230 & w1393) | (w1391 & w1393);
assign w1395 = pi197 & ~w1394;
assign w1396 = ~pi069 & pi196;
assign w1397 = ~pi197 & ~w1396;
assign w1398 = ~pi069 & w1378;
assign w1399 = ~pi069 & w1375;
assign w1400 = (w1342 & w1398) | (w1342 & w1399) | (w1398 & w1399);
assign w1401 = w1397 & ~w1400;
assign w1402 = ~pi070 & ~w1401;
assign w1403 = pi069 & w1397;
assign w1404 = (w1387 & w1397) | (w1387 & w1403) | (w1397 & w1403);
assign w1405 = ~pi070 & ~w1404;
assign w1406 = (w1230 & w1402) | (w1230 & w1405) | (w1402 & w1405);
assign w1407 = pi198 & ~w1406;
assign w1408 = ~pi071 & ~w62;
assign w1409 = ~pi198 & w22;
assign w1410 = ~w58 & w1409;
assign w1411 = (w1374 & w1409) | (w1374 & w1410) | (w1409 & w1410);
assign w1412 = w1344 & w1376;
assign w1413 = (w1409 & w1410) | (w1409 & w1412) | (w1410 & w1412);
assign w1414 = (~w1342 & w1411) | (~w1342 & w1413) | (w1411 & w1413);
assign w1415 = ~w1379 & w1414;
assign w1416 = w1408 & ~w1415;
assign w1417 = w1387 & w1414;
assign w1418 = w1408 & ~w1417;
assign w1419 = (w1230 & w1416) | (w1230 & w1418) | (w1416 & w1418);
assign w1420 = pi199 & ~w1419;
assign w1421 = w94 & w1154;
assign w1422 = (~w89 & w94) | (~w89 & w1421) | (w94 & w1421);
assign w1423 = w69 & ~w1422;
assign w1424 = w1229 & ~w1423;
assign w1425 = (~w1332 & ~w1423) | (~w1332 & w1424) | (~w1423 & w1424);
assign w1426 = w67 & ~w1425;
assign w1427 = pi200 & ~w1426;
assign w1428 = w830 & ~w1153;
assign w1429 = ~w318 & w741;
assign w1430 = w18 & ~w1029;
assign w1431 = (w18 & ~w1429) | (w18 & w1430) | (~w1429 & w1430);
assign w1432 = w68 & w89;
assign w1433 = w1431 & w1432;
assign w1434 = w1153 & w1433;
assign w1435 = w840 & w1149;
assign w1436 = w1433 & w1435;
assign w1437 = (~w1428 & w1434) | (~w1428 & w1436) | (w1434 & w1436);
assign w1438 = w1274 & w1437;
assign w1439 = w1235 & w1437;
assign w1440 = (w1230 & w1438) | (w1230 & w1439) | (w1438 & w1439);
assign w1441 = ~pi073 & pi200;
assign w1442 = (~pi073 & w1423) | (~pi073 & w1441) | (w1423 & w1441);
assign w1443 = (~pi073 & w1440) | (~pi073 & w1442) | (w1440 & w1442);
assign w1444 = pi201 & ~w1443;
assign w1445 = (~w1153 & w1428) | (~w1153 & ~w1435) | (w1428 & ~w1435);
assign w1446 = w94 & w127;
assign w1447 = w1139 & w1446;
assign w1448 = pi075 & ~pi207;
assign w1449 = w141 & w1448;
assign w1450 = w241 & ~w1449;
assign w1451 = w138 & ~w1450;
assign w1452 = w1447 & w1451;
assign w1453 = w1423 & ~w1452;
assign w1454 = ~w1423 & ~w1433;
assign w1455 = ~w1452 & ~w1454;
assign w1456 = (~w1445 & w1453) | (~w1445 & w1455) | (w1453 & w1455);
assign w1457 = ~pi074 & pi201;
assign w1458 = ~pi074 & ~w242;
assign w1459 = (pi200 & w1457) | (pi200 & w1458) | (w1457 & w1458);
assign w1460 = w94 & w430;
assign w1461 = w276 & w1460;
assign w1462 = w741 & w1461;
assign w1463 = w200 & w1462;
assign w1464 = ~pi200 & w1462;
assign w1465 = w127 & w232;
assign w1466 = w1226 & ~w1465;
assign w1467 = ~pi200 & ~w1466;
assign w1468 = (w1463 & w1464) | (w1463 & w1467) | (w1464 & w1467);
assign w1469 = (w1457 & w1458) | (w1457 & ~w1468) | (w1458 & ~w1468);
assign w1470 = (w1456 & w1459) | (w1456 & w1469) | (w1459 & w1469);
assign w1471 = pi202 & ~w1470;
assign w1472 = (~w1423 & w1445) | (~w1423 & w1454) | (w1445 & w1454);
assign w1473 = ~w144 & w245;
assign w1474 = w144 & w741;
assign w1475 = w1461 & w1474;
assign w1476 = w144 & ~w1466;
assign w1477 = (w1463 & w1475) | (w1463 & w1476) | (w1475 & w1476);
assign w1478 = w245 & ~w1477;
assign w1479 = (~w1472 & w1473) | (~w1472 & w1478) | (w1473 & w1478);
assign w1480 = w138 & w741;
assign w1481 = w1138 & w1480;
assign w1482 = w1446 & w1481;
assign w1483 = w144 & ~w241;
assign w1484 = w1482 & w1483;
assign w1485 = w1479 & ~w1484;
assign w1486 = pi203 & ~w1485;
assign w1487 = ~w1477 & ~w1484;
assign w1488 = (~w144 & ~w1472) | (~w144 & w1487) | (~w1472 & w1487);
assign w1489 = ~pi076 & pi203;
assign w1490 = pi075 & ~pi203;
assign w1491 = ~pi076 & ~w1490;
assign w1492 = (~w244 & w1489) | (~w244 & w1491) | (w1489 & w1491);
assign w1493 = (w1488 & w1489) | (w1488 & w1492) | (w1489 & w1492);
assign w1494 = pi204 & ~w1493;
assign w1495 = w1138 & w1446;
assign w1496 = ~pi076 & w1489;
assign w1497 = (~pi075 & ~pi076) | (~pi075 & w1489) | (~pi076 & w1489);
assign w1498 = (~w244 & w1496) | (~w244 & w1497) | (w1496 & w1497);
assign w1499 = (~w144 & w1489) | (~w144 & w1498) | (w1489 & w1498);
assign w1500 = w138 & ~w236;
assign w1501 = w741 & w1500;
assign w1502 = (~pi076 & ~w144) | (~pi076 & w1489) | (~w144 & w1489);
assign w1503 = (w245 & w1496) | (w245 & w1502) | (w1496 & w1502);
assign w1504 = (~w144 & w1489) | (~w144 & w1503) | (w1489 & w1503);
assign w1505 = (w1499 & ~w1501) | (w1499 & w1504) | (~w1501 & w1504);
assign w1506 = (~w1495 & w1499) | (~w1495 & w1505) | (w1499 & w1505);
assign w1507 = (w1498 & ~w1501) | (w1498 & w1503) | (~w1501 & w1503);
assign w1508 = (~w1495 & w1498) | (~w1495 & w1507) | (w1498 & w1507);
assign w1509 = (~w1477 & w1489) | (~w1477 & w1508) | (w1489 & w1508);
assign w1510 = (~w1472 & w1506) | (~w1472 & w1509) | (w1506 & w1509);
assign w1511 = ~pi077 & pi204;
assign w1512 = (~pi077 & w1510) | (~pi077 & w1511) | (w1510 & w1511);
assign w1513 = pi205 & ~w1512;
assign w1514 = ~pi076 & ~pi077;
assign w1515 = ~pi075 & w1514;
assign w1516 = ~w244 & w1515;
assign w1517 = ~w144 & w1516;
assign w1518 = ~pi080 & ~w234;
assign w1519 = w144 & ~w1518;
assign w1520 = w1514 & ~w1519;
assign w1521 = (~w138 & w1514) | (~w138 & w1520) | (w1514 & w1520);
assign w1522 = w1473 & w1521;
assign w1523 = (~w1447 & w1517) | (~w1447 & w1522) | (w1517 & w1522);
assign w1524 = w245 & w1521;
assign w1525 = (~w1447 & w1516) | (~w1447 & w1524) | (w1516 & w1524);
assign w1526 = ~w1477 & w1525;
assign w1527 = (~w1472 & w1523) | (~w1472 & w1526) | (w1523 & w1526);
assign w1528 = (~pi077 & w1489) | (~pi077 & w1511) | (w1489 & w1511);
assign w1529 = ~pi078 & pi205;
assign w1530 = (~pi078 & w1528) | (~pi078 & w1529) | (w1528 & w1529);
assign w1531 = (~pi078 & w1527) | (~pi078 & w1530) | (w1527 & w1530);
assign w1532 = pi206 & ~w1531;
assign w1533 = ~pi079 & ~w233;
assign w1534 = ~pi206 & ~w1529;
assign w1535 = (w233 & ~w1528) | (w233 & w1534) | (~w1528 & w1534);
assign w1536 = ~pi079 & ~w1535;
assign w1537 = (w1527 & w1533) | (w1527 & w1536) | (w1533 & w1536);
assign w1538 = pi207 & ~w1537;
assign w1539 = ~pi088 & pi215;
assign w1540 = ~pi088 & ~w214;
assign w1541 = (~w213 & w1539) | (~w213 & w1540) | (w1539 & w1540);
assign w1542 = ~w223 & w1541;
assign w1543 = ~pi218 & w206;
assign w1544 = w204 & ~w1543;
assign w1545 = (w204 & w1542) | (w204 & w1544) | (w1542 & w1544);
assign w1546 = pi092 & ~pi202;
assign w1547 = w143 & w1546;
assign w1548 = w142 & w1547;
assign w1549 = w144 & ~w205;
assign w1550 = w142 & w1549;
assign w1551 = (~w1545 & w1548) | (~w1545 & w1550) | (w1548 & w1550);
assign w1552 = w1447 & w1551;
assign w1553 = w144 & w208;
assign w1554 = w142 & w1553;
assign w1555 = w230 & w1554;
assign w1556 = w1447 & w1555;
assign w1557 = ~w1552 & ~w1556;
assign w1558 = w142 & ~w1473;
assign w1559 = w241 & ~w1558;
assign w1560 = w1557 & w1559;
assign w1561 = ~w200 & w1226;
assign w1562 = w241 & w245;
assign w1563 = ~w1559 & ~w1562;
assign w1564 = ~w741 & w1562;
assign w1565 = ~w1559 & ~w1564;
assign w1566 = (w1461 & w1563) | (w1461 & w1565) | (w1563 & w1565);
assign w1567 = (~w1561 & w1563) | (~w1561 & w1566) | (w1563 & w1566);
assign w1568 = w1557 & ~w1567;
assign w1569 = (~w1472 & w1560) | (~w1472 & w1568) | (w1560 & w1568);
assign w1570 = pi208 & ~w1569;
assign w1571 = (w1472 & ~w1559) | (w1472 & w1567) | (~w1559 & w1567);
assign w1572 = ~pi081 & pi208;
assign w1573 = (~pi081 & w1557) | (~pi081 & w1572) | (w1557 & w1572);
assign w1574 = (~w1571 & w1572) | (~w1571 & w1573) | (w1572 & w1573);
assign w1575 = pi209 & ~w1574;
assign w1576 = ~w1551 & w1559;
assign w1577 = (~w1447 & w1559) | (~w1447 & w1576) | (w1559 & w1576);
assign w1578 = ~w1552 & ~w1567;
assign w1579 = (~w1472 & w1577) | (~w1472 & w1578) | (w1577 & w1578);
assign w1580 = ~pi081 & ~pi082;
assign w1581 = pi083 & ~pi215;
assign w1582 = ~pi082 & ~w1581;
assign w1583 = (~pi082 & ~w130) | (~pi082 & w1582) | (~w130 & w1582);
assign w1584 = ~pi081 & w1583;
assign w1585 = (~w1554 & w1580) | (~w1554 & w1584) | (w1580 & w1584);
assign w1586 = (~w1447 & w1580) | (~w1447 & w1585) | (w1580 & w1585);
assign w1587 = w1579 & w1586;
assign w1588 = ~pi082 & pi209;
assign w1589 = (~pi082 & w1572) | (~pi082 & w1588) | (w1572 & w1588);
assign w1590 = pi210 & ~w1589;
assign w1591 = ~w1587 & w1590;
assign w1592 = ~pi210 & w133;
assign w1593 = w229 & ~w1592;
assign w1594 = (w229 & w1579) | (w229 & w1593) | (w1579 & w1593);
assign w1595 = pi211 & ~w1594;
assign w1596 = ~pi210 & ~pi211;
assign w1597 = w133 & w1596;
assign w1598 = ~w1541 & w1597;
assign w1599 = w1554 & w1598;
assign w1600 = w1447 & w1599;
assign w1601 = ~pi083 & ~pi084;
assign w1602 = ~w228 & w1601;
assign w1603 = w241 & w1602;
assign w1604 = ~w1558 & w1603;
assign w1605 = pi091 & ~pi219;
assign w1606 = ~pi092 & ~w1605;
assign w1607 = (~w203 & w205) | (~w203 & w1606) | (w205 & w1606);
assign w1608 = ~pi084 & w1607;
assign w1609 = (~pi084 & ~w145) | (~pi084 & w1608) | (~w145 & w1608);
assign w1610 = w229 & w1609;
assign w1611 = w1559 & w1610;
assign w1612 = (~w1447 & w1604) | (~w1447 & w1611) | (w1604 & w1611);
assign w1613 = (~w1447 & w1602) | (~w1447 & w1610) | (w1602 & w1610);
assign w1614 = w1612 & w1613;
assign w1615 = (~w1461 & w1562) | (~w1461 & w1564) | (w1562 & w1564);
assign w1616 = (w1561 & w1562) | (w1561 & w1615) | (w1562 & w1615);
assign w1617 = (w1612 & w1613) | (w1612 & w1616) | (w1613 & w1616);
assign w1618 = (~w1472 & w1614) | (~w1472 & w1617) | (w1614 & w1617);
assign w1619 = ~pi084 & pi211;
assign w1620 = ~pi084 & ~w1597;
assign w1621 = (w229 & w1619) | (w229 & w1620) | (w1619 & w1620);
assign w1622 = ~w1599 & w1621;
assign w1623 = (~w1447 & w1621) | (~w1447 & w1622) | (w1621 & w1622);
assign w1624 = (~w1600 & w1618) | (~w1600 & w1623) | (w1618 & w1623);
assign w1625 = pi212 & ~w1624;
assign w1626 = ~w1472 & w1616;
assign w1627 = (~pi215 & w212) | (~pi215 & w214) | (w212 & w214);
assign w1628 = ~pi088 & ~w1627;
assign w1629 = w1554 & ~w1628;
assign w1630 = w1447 & w1629;
assign w1631 = w1612 & ~w1630;
assign w1632 = (~pi211 & ~pi212) | (~pi211 & w221) | (~pi212 & w221);
assign w1633 = (~pi212 & w221) | (~pi212 & w1597) | (w221 & w1597);
assign w1634 = (~w229 & w1632) | (~w229 & w1633) | (w1632 & w1633);
assign w1635 = ~pi085 & ~w1634;
assign w1636 = (~pi085 & w1631) | (~pi085 & w1635) | (w1631 & w1635);
assign w1637 = w1613 & ~w1630;
assign w1638 = (~pi085 & w1635) | (~pi085 & w1637) | (w1635 & w1637);
assign w1639 = (w1626 & w1636) | (w1626 & w1638) | (w1636 & w1638);
assign w1640 = pi213 & ~w1639;
assign w1641 = ~pi086 & pi213;
assign w1642 = ~pi086 & ~w211;
assign w1643 = w1641 | w1642;
assign w1644 = (~w1634 & w1641) | (~w1634 & w1642) | (w1641 & w1642);
assign w1645 = (w1631 & w1643) | (w1631 & w1644) | (w1643 & w1644);
assign w1646 = (w1637 & w1643) | (w1637 & w1644) | (w1643 & w1644);
assign w1647 = (w1626 & w1645) | (w1626 & w1646) | (w1645 & w1646);
assign w1648 = pi214 & ~w1647;
assign w1649 = ~pi087 & ~w213;
assign w1650 = ~pi087 & ~pi088;
assign w1651 = (~pi087 & ~w1597) | (~pi087 & w1650) | (~w1597 & w1650);
assign w1652 = ~w213 & w1651;
assign w1653 = (~w1554 & w1649) | (~w1554 & w1652) | (w1649 & w1652);
assign w1654 = (~w1447 & w1649) | (~w1447 & w1653) | (w1649 & w1653);
assign w1655 = w1621 & w1649;
assign w1656 = pi088 & w1597;
assign w1657 = w1554 & w1656;
assign w1658 = ~pi087 & w1621;
assign w1659 = ~w1657 & w1658;
assign w1660 = ~w213 & w1659;
assign w1661 = (~w1447 & w1655) | (~w1447 & w1660) | (w1655 & w1660);
assign w1662 = (w1618 & w1654) | (w1618 & w1661) | (w1654 & w1661);
assign w1663 = ~pi212 & pi215;
assign w1664 = w129 & w1663;
assign w1665 = (pi215 & ~w1649) | (pi215 & w1664) | (~w1649 & w1664);
assign w1666 = ~w1662 & w1665;
assign w1667 = ~pi212 & ~pi213;
assign w1668 = ~pi214 & ~pi215;
assign w1669 = w1667 & w1668;
assign w1670 = w1541 & ~w1669;
assign w1671 = (w1541 & w1621) | (w1541 & w1670) | (w1621 & w1670);
assign w1672 = (w1541 & w1618) | (w1541 & w1671) | (w1618 & w1671);
assign w1673 = pi216 & ~w1672;
assign w1674 = w225 & w1592;
assign w1675 = ~w230 & w1542;
assign w1676 = w1559 & w1675;
assign w1677 = w144 & ~w1606;
assign w1678 = w142 & w1677;
assign w1679 = w1674 & w1678;
assign w1680 = w1675 & ~w1679;
assign w1681 = w1559 & w1680;
assign w1682 = (~w1447 & w1676) | (~w1447 & w1681) | (w1676 & w1681);
assign w1683 = (~w1447 & w1675) | (~w1447 & w1680) | (w1675 & w1680);
assign w1684 = (~w1674 & w1682) | (~w1674 & w1683) | (w1682 & w1683);
assign w1685 = ~w1562 & w1674;
assign w1686 = ~w1564 & w1674;
assign w1687 = (w1461 & w1685) | (w1461 & w1686) | (w1685 & w1686);
assign w1688 = (~w1561 & w1685) | (~w1561 & w1687) | (w1685 & w1687);
assign w1689 = (w1682 & w1683) | (w1682 & ~w1688) | (w1683 & ~w1688);
assign w1690 = (~w1472 & w1684) | (~w1472 & w1689) | (w1684 & w1689);
assign w1691 = ~pi089 & pi216;
assign w1692 = w145 & w1674;
assign w1693 = ~pi216 & ~pi219;
assign w1694 = w202 & w1693;
assign w1695 = ~pi089 & ~w1694;
assign w1696 = (~pi089 & ~w1692) | (~pi089 & w1695) | (~w1692 & w1695);
assign w1697 = (~pi089 & ~w1447) | (~pi089 & w1696) | (~w1447 & w1696);
assign w1698 = (w1690 & w1691) | (w1690 & w1697) | (w1691 & w1697);
assign w1699 = pi217 & ~w1698;
assign w1700 = (~pi089 & w1675) | (~pi089 & w1691) | (w1675 & w1691);
assign w1701 = (~pi089 & w1680) | (~pi089 & w1691) | (w1680 & w1691);
assign w1702 = (~w1447 & w1700) | (~w1447 & w1701) | (w1700 & w1701);
assign w1703 = ~pi216 & ~w1681;
assign w1704 = ~pi216 & ~w1675;
assign w1705 = (~pi216 & ~w1559) | (~pi216 & w1704) | (~w1559 & w1704);
assign w1706 = (w1447 & w1703) | (w1447 & w1705) | (w1703 & w1705);
assign w1707 = ~pi089 & ~w1706;
assign w1708 = (~w1674 & w1702) | (~w1674 & w1707) | (w1702 & w1707);
assign w1709 = (~w1688 & w1702) | (~w1688 & w1707) | (w1702 & w1707);
assign w1710 = (~w1472 & w1708) | (~w1472 & w1709) | (w1708 & w1709);
assign w1711 = ~pi090 & pi217;
assign w1712 = (~pi090 & w1710) | (~pi090 & w1711) | (w1710 & w1711);
assign w1713 = pi218 & ~w1712;
assign w1714 = (w204 & w1544) | (w204 & w1690) | (w1544 & w1690);
assign w1715 = pi219 & ~w1714;
assign w1716 = ~w146 & w249;
assign w1717 = w146 & ~w1562;
assign w1718 = w146 & ~w1615;
assign w1719 = (~w1561 & w1717) | (~w1561 & w1718) | (w1717 & w1718);
assign w1720 = w249 & ~w1719;
assign w1721 = (~w1472 & w1716) | (~w1472 & w1720) | (w1716 & w1720);
assign w1722 = pi220 & ~w1721;
assign w1723 = ~pi220 & w146;
assign w1724 = w76 & ~w1058;
assign w1725 = w82 & ~w1724;
assign w1726 = ~w88 & w1725;
assign w1727 = w94 & ~w1726;
assign w1728 = w34 & w1723;
assign w1729 = (w1723 & w1727) | (w1723 & w1728) | (w1727 & w1728);
assign w1730 = w89 & w1431;
assign w1731 = w1729 & ~w1730;
assign w1732 = (w1027 & w1729) | (w1027 & w1731) | (w1729 & w1731);
assign w1733 = ~w68 & w146;
assign w1734 = w249 & ~w1733;
assign w1735 = ~pi093 & pi220;
assign w1736 = (~pi093 & w1734) | (~pi093 & w1735) | (w1734 & w1735);
assign w1737 = ~w1732 & w1736;
assign w1738 = w741 & w1723;
assign w1739 = w1461 & w1738;
assign w1740 = ~w1561 & w1739;
assign w1741 = w1737 & ~w1740;
assign w1742 = pi221 & ~w1741;
assign w1743 = ~pi094 & pi221;
assign w1744 = ~pi221 & w1739;
assign w1745 = ~w1561 & w1744;
assign w1746 = ~pi094 & ~w1745;
assign w1747 = (w1737 & w1743) | (w1737 & w1746) | (w1743 & w1746);
assign w1748 = pi222 & ~w1747;
assign w1749 = ~pi221 & ~w1736;
assign w1750 = (~pi221 & w1732) | (~pi221 & w1749) | (w1732 & w1749);
assign w1751 = w122 & w1739;
assign w1752 = ~pi110 & ~w178;
assign w1753 = ~w174 & w1752;
assign w1754 = (w162 & w1752) | (w162 & w1753) | (w1752 & w1753);
assign w1755 = pi096 & ~pi224;
assign w1756 = pi097 & ~pi225;
assign w1757 = (~pi225 & w1755) | (~pi225 & w1756) | (w1755 & w1756);
assign w1758 = ~pi098 & ~w1757;
assign w1759 = w105 & w195;
assign w1760 = ~w1758 & w1759;
assign w1761 = w199 & w1760;
assign w1762 = (w199 & ~w1754) | (w199 & w1761) | (~w1754 & w1761);
assign w1763 = ~pi112 & ~w329;
assign w1764 = w120 & ~w1763;
assign w1765 = w327 & ~w1764;
assign w1766 = w116 & ~w1765;
assign w1767 = w349 & ~w1766;
assign w1768 = ~w1762 & w1767;
assign w1769 = ~pi095 & w1768;
assign w1770 = (~pi095 & ~w1751) | (~pi095 & w1769) | (~w1751 & w1769);
assign w1771 = pi222 & w1770;
assign w1772 = ~w179 & w1770;
assign w1773 = (~w1750 & w1771) | (~w1750 & w1772) | (w1771 & w1772);
assign w1774 = pi223 & ~w1773;
assign w1775 = pi093 & w122;
assign w1776 = w122 & ~w1735;
assign w1777 = (~w1734 & w1775) | (~w1734 & w1776) | (w1775 & w1776);
assign w1778 = (w122 & w1732) | (w122 & w1777) | (w1732 & w1777);
assign w1779 = ~pi095 & ~w179;
assign w1780 = ~pi098 & ~w1756;
assign w1781 = w1759 & ~w1780;
assign w1782 = w199 & w1781;
assign w1783 = (w199 & ~w1754) | (w199 & w1782) | (~w1754 & w1782);
assign w1784 = w1767 & ~w1783;
assign w1785 = w1779 & w1784;
assign w1786 = (~w1751 & w1779) | (~w1751 & w1785) | (w1779 & w1785);
assign w1787 = ~pi223 & ~w1786;
assign w1788 = (~pi223 & w1778) | (~pi223 & w1787) | (w1778 & w1787);
assign w1789 = ~pi096 & ~w1788;
assign w1790 = pi224 & ~w1789;
assign w1791 = w182 & ~w1788;
assign w1792 = pi225 & ~w188;
assign w1793 = ~w1791 & w1792;
assign w1794 = ~w122 & w183;
assign w1795 = w183 & ~w1777;
assign w1796 = (~w1732 & w1794) | (~w1732 & w1795) | (w1794 & w1795);
assign w1797 = ~w191 & ~w1770;
assign w1798 = (~w191 & ~w1796) | (~w191 & w1797) | (~w1796 & w1797);
assign w1799 = pi226 & w1798;
assign w1800 = w94 & w126;
assign w1801 = w276 & w1800;
assign w1802 = w858 & w1723;
assign w1803 = w1801 & w1802;
assign w1804 = ~pi098 & ~pi099;
assign w1805 = ~pi099 & w190;
assign w1806 = (w189 & w1804) | (w189 & w1805) | (w1804 & w1805);
assign w1807 = ~pi226 & ~w182;
assign w1808 = (~pi226 & ~w181) | (~pi226 & w1807) | (~w181 & w1807);
assign w1809 = (~pi099 & w1806) | (~pi099 & ~w1808) | (w1806 & ~w1808);
assign w1810 = (~pi106 & w167) | (~pi106 & w169) | (w167 & w169);
assign w1811 = (~pi106 & w161) | (~pi106 & w1810) | (w161 & w1810);
assign w1812 = pi107 & ~pi235;
assign w1813 = (~pi236 & w176) | (~pi236 & w1812) | (w176 & w1812);
assign w1814 = ~pi109 & ~w1813;
assign w1815 = w183 & w1814;
assign w1816 = ~pi234 & w163;
assign w1817 = w1814 & ~w1816;
assign w1818 = w183 & w1817;
assign w1819 = (w1811 & w1815) | (w1811 & w1818) | (w1815 & w1818);
assign w1820 = ~pi099 | w1806;
assign w1821 = (~pi099 & pi226) | (~pi099 & w1806) | (pi226 & w1806);
assign w1822 = (w1819 & w1820) | (w1819 & w1821) | (w1820 & w1821);
assign w1823 = (~w1803 & w1809) | (~w1803 & w1822) | (w1809 & w1822);
assign w1824 = ~w1226 & w1739;
assign w1825 = w1736 & ~w1824;
assign w1826 = ~w1732 & w1825;
assign w1827 = pi098 & w122;
assign w1828 = w122 & ~w190;
assign w1829 = (~w189 & w1827) | (~w189 & w1828) | (w1827 & w1828);
assign w1830 = ~pi226 & w1829;
assign w1831 = w1809 & ~w1830;
assign w1832 = w1821 & ~w1830;
assign w1833 = w1820 & ~w1830;
assign w1834 = (w1819 & w1832) | (w1819 & w1833) | (w1832 & w1833);
assign w1835 = (~w1803 & w1831) | (~w1803 & w1834) | (w1831 & w1834);
assign w1836 = (w1823 & w1826) | (w1823 & w1835) | (w1826 & w1835);
assign w1837 = pi227 & ~w1836;
assign w1838 = ~pi100 & pi227;
assign w1839 = (~pi100 & w1835) | (~pi100 & w1838) | (w1835 & w1838);
assign w1840 = (~pi100 & w1823) | (~pi100 & w1838) | (w1823 & w1838);
assign w1841 = (w1826 & w1839) | (w1826 & w1840) | (w1839 & w1840);
assign w1842 = pi228 & ~w1841;
assign w1843 = ~pi101 & pi228;
assign w1844 = (~pi101 & w1838) | (~pi101 & w1843) | (w1838 & w1843);
assign w1845 = ~pi101 & ~w157;
assign w1846 = (w1835 & w1844) | (w1835 & w1845) | (w1844 & w1845);
assign w1847 = (w1823 & w1844) | (w1823 & w1845) | (w1844 & w1845);
assign w1848 = (w1826 & w1846) | (w1826 & w1847) | (w1846 & w1847);
assign w1849 = pi229 & ~w1848;
assign w1850 = w122 & ~w1226;
assign w1851 = w1739 & w1850;
assign w1852 = w183 & ~w1851;
assign w1853 = ~pi099 & ~pi100;
assign w1854 = pi105 & ~pi233;
assign w1855 = ~pi106 & ~w1854;
assign w1856 = w1816 & ~w1855;
assign w1857 = w1814 & ~w1856;
assign w1858 = w1853 & w1857;
assign w1859 = (~w1803 & w1853) | (~w1803 & w1858) | (w1853 & w1858);
assign w1860 = w1852 & w1859;
assign w1861 = ~w1778 & w1860;
assign w1862 = w153 & ~w1843;
assign w1863 = ~pi102 & ~w1862;
assign w1864 = ~pi223 & ~pi224;
assign w1865 = ~pi225 & w1864;
assign w1866 = pi103 & ~pi231;
assign w1867 = ~pi104 & ~w1866;
assign w1868 = w1865 & ~w1867;
assign w1869 = ~pi227 & ~pi236;
assign w1870 = ~pi232 & w1869;
assign w1871 = w99 & w1870;
assign w1872 = w1868 & w1871;
assign w1873 = ~pi102 & pi229;
assign w1874 = (~pi102 & w1843) | (~pi102 & w1873) | (w1843 & w1873);
assign w1875 = (w1863 & ~w1872) | (w1863 & w1874) | (~w1872 & w1874);
assign w1876 = (~w1803 & w1863) | (~w1803 & w1875) | (w1863 & w1875);
assign w1877 = pi098 & ~pi226;
assign w1878 = ~pi226 & ~w190;
assign w1879 = (~w189 & w1877) | (~w189 & w1878) | (w1877 & w1878);
assign w1880 = ~pi229 & ~w1843;
assign w1881 = pi099 & ~pi227;
assign w1882 = ~pi100 & ~pi101;
assign w1883 = ~w1881 & w1882;
assign w1884 = w1880 & ~w1883;
assign w1885 = ~pi101 & w1838;
assign w1886 = w1880 & ~w1885;
assign w1887 = (w1879 & w1884) | (w1879 & w1886) | (w1884 & w1886);
assign w1888 = ~pi102 & ~w1887;
assign w1889 = (~w1879 & w1883) | (~w1879 & w1885) | (w1883 & w1885);
assign w1890 = ~w1872 & w1889;
assign w1891 = (~pi102 & w1874) | (~pi102 & w1890) | (w1874 & w1890);
assign w1892 = (~w1803 & w1888) | (~w1803 & w1891) | (w1888 & w1891);
assign w1893 = (w1861 & w1876) | (w1861 & w1892) | (w1876 & w1892);
assign w1894 = pi230 & ~w1893;
assign w1895 = ~pi228 & ~pi229;
assign w1896 = ~pi230 & w1895;
assign w1897 = w156 & ~w1896;
assign w1898 = (w156 & ~w1872) | (w156 & w1897) | (~w1872 & w1897);
assign w1899 = (w156 & ~w1803) | (w156 & w1898) | (~w1803 & w1898);
assign w1900 = ~w1838 & w1896;
assign w1901 = ~pi100 & ~w1881;
assign w1902 = w1896 & ~w1901;
assign w1903 = (w1879 & w1900) | (w1879 & w1902) | (w1900 & w1902);
assign w1904 = w156 & ~w1903;
assign w1905 = (w1838 & ~w1879) | (w1838 & w1901) | (~w1879 & w1901);
assign w1906 = ~w1872 & w1905;
assign w1907 = (w156 & w1897) | (w156 & w1906) | (w1897 & w1906);
assign w1908 = (~w1803 & w1904) | (~w1803 & w1907) | (w1904 & w1907);
assign w1909 = (w1861 & w1899) | (w1861 & w1908) | (w1899 & w1908);
assign w1910 = pi231 & ~w1909;
assign w1911 = (~w155 & w165) | (~w155 & w1867) | (w165 & w1867);
assign w1912 = (w165 & ~w1903) | (w165 & w1911) | (~w1903 & w1911);
assign w1913 = (w1861 & w1911) | (w1861 & w1912) | (w1911 & w1912);
assign w1914 = pi232 & ~w1913;
assign w1915 = ~w161 & ~w167;
assign w1916 = w105 & ~w1831;
assign w1917 = w105 & ~w1834;
assign w1918 = (w1803 & w1916) | (w1803 & w1917) | (w1916 & w1917);
assign w1919 = ~w1915 & ~w1918;
assign w1920 = w105 & ~w1809;
assign w1921 = w105 & ~w1822;
assign w1922 = (w1803 & w1920) | (w1803 & w1921) | (w1920 & w1921);
assign w1923 = ~w1915 & ~w1922;
assign w1924 = (w1826 & w1919) | (w1826 & w1923) | (w1919 & w1923);
assign w1925 = pi233 & ~w1924;
assign w1926 = ~w150 & w167;
assign w1927 = (~w150 & w161) | (~w150 & w1926) | (w161 & w1926);
assign w1928 = (~pi106 & w169) | (~pi106 & w1927) | (w169 & w1927);
assign w1929 = ~w1814 & w1865;
assign w1930 = w191 & ~w1929;
assign w1931 = (w191 & ~w1803) | (w191 & w1930) | (~w1803 & w1930);
assign w1932 = w1803 & w1929;
assign w1933 = ~w183 & ~w191;
assign w1934 = (~w191 & w1851) | (~w191 & w1933) | (w1851 & w1933);
assign w1935 = ~w1932 & ~w1934;
assign w1936 = (~w1778 & w1931) | (~w1778 & w1935) | (w1931 & w1935);
assign w1937 = ~pi226 & w104;
assign w1938 = w103 & w1937;
assign w1939 = (~pi106 & w169) | (~pi106 & ~w1938) | (w169 & ~w1938);
assign w1940 = pi233 & w169;
assign w1941 = (w169 & ~w1938) | (w169 & w1940) | (~w1938 & w1940);
assign w1942 = (w1927 & w1939) | (w1927 & w1941) | (w1939 & w1941);
assign w1943 = (w1928 & w1936) | (w1928 & w1942) | (w1936 & w1942);
assign w1944 = pi234 & ~w1943;
assign w1945 = ~pi107 & ~w171;
assign w1946 = ~w162 & ~w1945;
assign w1947 = ~pi233 & ~pi234;
assign w1948 = w1938 & w1947;
assign w1949 = ~w1823 & w1948;
assign w1950 = ~w1946 & ~w1949;
assign w1951 = ~w1835 & w1948;
assign w1952 = ~w1946 & ~w1951;
assign w1953 = (w1826 & w1950) | (w1826 & w1952) | (w1950 & w1952);
assign w1954 = pi235 & ~w1953;
assign w1955 = pi109 & ~pi225;
assign w1956 = w1864 & w1955;
assign w1957 = w191 & ~w1956;
assign w1958 = (w191 & ~w1803) | (w191 & w1957) | (~w1803 & w1957);
assign w1959 = w1803 & w1956;
assign w1960 = ~w1934 & ~w1959;
assign w1961 = (~w1778 & w1958) | (~w1778 & w1960) | (w1958 & w1960);
assign w1962 = ~pi107 & ~pi108;
assign w1963 = ~w171 & w1962;
assign w1964 = (~pi108 & w162) | (~pi108 & w1963) | (w162 & w1963);
assign w1965 = w1961 & w1964;
assign w1966 = w1945 & ~w1948;
assign w1967 = (w162 & ~w1948) | (w162 & w1966) | (~w1948 & w1966);
assign w1968 = pi108 & pi236;
assign w1969 = ~pi108 & pi235;
assign w1970 = pi236 & ~w1969;
assign w1971 = (~w1967 & w1968) | (~w1967 & w1970) | (w1968 & w1970);
assign w1972 = ~w1965 & w1971;
assign w1973 = ~w163 & w1814;
assign w1974 = (w1814 & w1967) | (w1814 & w1973) | (w1967 & w1973);
assign w1975 = w163 & ~w1945;
assign w1976 = ~w162 & w1975;
assign w1977 = w1814 & ~w1976;
assign w1978 = (w191 & w1974) | (w191 & w1977) | (w1974 & w1977);
assign w1979 = (~w1934 & w1974) | (~w1934 & w1977) | (w1974 & w1977);
assign w1980 = (~w1778 & w1978) | (~w1778 & w1979) | (w1978 & w1979);
assign w1981 = pi237 & ~w1980;
assign w1982 = ~w191 & w1759;
assign w1983 = w1754 & ~w1982;
assign w1984 = w1759 & w1933;
assign w1985 = (w1851 & w1982) | (w1851 & w1984) | (w1982 & w1984);
assign w1986 = w1754 & ~w1985;
assign w1987 = (~w1778 & w1983) | (~w1778 & w1986) | (w1983 & w1986);
assign w1988 = pi238 & ~w1987;
assign w1989 = ~pi111 & pi238;
assign w1990 = (~pi111 & w1754) | (~pi111 & w1989) | (w1754 & w1989);
assign w1991 = (~w1982 & w1989) | (~w1982 & w1990) | (w1989 & w1990);
assign w1992 = (~w1985 & w1989) | (~w1985 & w1990) | (w1989 & w1990);
assign w1993 = (~w1778 & w1991) | (~w1778 & w1992) | (w1991 & w1992);
assign w1994 = pi239 & ~w1993;
assign w1995 = w105 & w124;
assign w1996 = ~pi223 & w194;
assign w1997 = w99 & w1996;
assign w1998 = w108 & w1997;
assign w1999 = w1995 & w1998;
assign w2000 = w1739 & w1999;
assign w2001 = ~w1767 & w2000;
assign w2002 = w105 & ~w183;
assign w2003 = ~w191 & w195;
assign w2004 = w2002 & w2003;
assign w2005 = w1752 & ~w2004;
assign w2006 = ~w175 & w2005;
assign w2007 = w124 & ~w191;
assign w2008 = w1759 & w2007;
assign w2009 = w1763 & ~w2008;
assign w2010 = ~w123 & w1763;
assign w2011 = ~w2008 & w2010;
assign w2012 = (w2006 & w2009) | (w2006 & w2011) | (w2009 & w2011);
assign w2013 = (w1763 & w2006) | (w1763 & w2010) | (w2006 & w2010);
assign w2014 = pi093 & w2008;
assign w2015 = ~w1735 & w2008;
assign w2016 = (~w1734 & w2014) | (~w1734 & w2015) | (w2014 & w2015);
assign w2017 = w2013 & ~w2016;
assign w2018 = (~w1732 & w2012) | (~w1732 & w2017) | (w2012 & w2017);
assign w2019 = ~w2001 & w2018;
assign w2020 = pi240 & ~w2019;
assign w2021 = (w1732 & w2008) | (w1732 & w2016) | (w2008 & w2016);
assign w2022 = ~pi113 & pi240;
assign w2023 = pi116 & ~pi244;
assign w2024 = ~pi117 & ~pi124;
assign w2025 = ~w2023 & w2024;
assign w2026 = (~pi124 & ~w116) | (~pi124 & w2025) | (~w116 & w2025);
assign w2027 = pi115 & ~pi244;
assign w2028 = (~pi244 & w320) | (~pi244 & w2027) | (w320 & w2027);
assign w2029 = ~pi243 & w2028;
assign w2030 = w116 & w2029;
assign w2031 = w2026 & ~w2030;
assign w2032 = w348 & w2031;
assign w2033 = w1999 & ~w2032;
assign w2034 = w1739 & w2033;
assign w2035 = ~pi240 & ~w1763;
assign w2036 = ~pi240 & ~w2010;
assign w2037 = (~w2006 & w2035) | (~w2006 & w2036) | (w2035 & w2036);
assign w2038 = (~pi240 & w2034) | (~pi240 & w2037) | (w2034 & w2037);
assign w2039 = ~pi113 & ~w2038;
assign w2040 = (~w2021 & w2022) | (~w2021 & w2039) | (w2022 & w2039);
assign w2041 = pi241 & ~w2040;
assign w2042 = ~pi113 & ~pi114;
assign w2043 = pi240 & w2042;
assign w2044 = ~w2038 & w2042;
assign w2045 = (~w2021 & w2043) | (~w2021 & w2044) | (w2043 & w2044);
assign w2046 = ~pi114 & pi241;
assign w2047 = pi242 & ~w2046;
assign w2048 = ~w2045 & w2047;
assign w2049 = ~pi115 & ~w321;
assign w2050 = ~pi242 & w117;
assign w2051 = w2049 & ~w2050;
assign w2052 = w348 & w2026;
assign w2053 = w1999 & ~w2052;
assign w2054 = w2050 & w2053;
assign w2055 = w1739 & w2054;
assign w2056 = w2049 & ~w2055;
assign w2057 = (w2018 & w2051) | (w2018 & w2056) | (w2051 & w2056);
assign w2058 = pi243 & ~w2057;
assign w2059 = ~pi115 & ~pi116;
assign w2060 = ~w321 & w2059;
assign w2061 = ~w2050 & w2060;
assign w2062 = ~w2055 & w2060;
assign w2063 = (w2018 & w2061) | (w2018 & w2062) | (w2061 & w2062);
assign w2064 = pi244 & ~w322;
assign w2065 = ~w2063 & w2064;
assign w2066 = ~w120 & w327;
assign w2067 = w120 & w2053;
assign w2068 = w1739 & w2067;
assign w2069 = w327 & ~w2068;
assign w2070 = (w2018 & w2066) | (w2018 & w2069) | (w2066 & w2069);
assign w2071 = pi245 & ~w2070;
assign w2072 = ~pi117 & ~pi118;
assign w2073 = ~pi118 & w326;
assign w2074 = (w325 & w2072) | (w325 & w2073) | (w2072 & w2073);
assign w2075 = ~w120 & w2074;
assign w2076 = ~w2068 & w2074;
assign w2077 = (w2018 & w2075) | (w2018 & w2076) | (w2075 & w2076);
assign w2078 = ~pi118 & pi245;
assign w2079 = pi246 & ~w2078;
assign w2080 = ~w2077 & w2079;
assign w2081 = w114 & w1999;
assign w2082 = ~pi124 & pi251;
assign w2083 = (~pi124 & w346) | (~pi124 & w2082) | (w346 & w2082);
assign w2084 = w120 & ~w2083;
assign w2085 = w2081 & w2084;
assign w2086 = ~pi119 & ~w2085;
assign w2087 = (~pi119 & ~w1739) | (~pi119 & w2086) | (~w1739 & w2086);
assign w2088 = w1763 & w2072;
assign w2089 = w1763 & w2073;
assign w2090 = (w325 & w2088) | (w325 & w2089) | (w2088 & w2089);
assign w2091 = w2010 & w2074;
assign w2092 = (w2006 & w2090) | (w2006 & w2091) | (w2090 & w2091);
assign w2093 = w1736 & w2092;
assign w2094 = ~w1732 & w2093;
assign w2095 = pi117 & ~pi245;
assign w2096 = ~pi118 & ~w2095;
assign w2097 = (~pi118 & w326) | (~pi118 & w2078) | (w326 & w2078);
assign w2098 = (w325 & w2096) | (w325 & w2097) | (w2096 & w2097);
assign w2099 = (~w120 & w2078) | (~w120 & w2098) | (w2078 & w2098);
assign w2100 = w120 & ~w2010;
assign w2101 = (w2078 & w2098) | (w2078 & ~w2100) | (w2098 & ~w2100);
assign w2102 = (~w2008 & w2099) | (~w2008 & w2101) | (w2099 & w2101);
assign w2103 = ~pi246 & ~w2102;
assign w2104 = (~w1764 & w2078) | (~w1764 & w2098) | (w2078 & w2098);
assign w2105 = (~w2008 & w2099) | (~w2008 & w2104) | (w2099 & w2104);
assign w2106 = ~pi246 & ~w2105;
assign w2107 = (~w2006 & w2103) | (~w2006 & w2106) | (w2103 & w2106);
assign w2108 = w2087 & ~w2107;
assign w2109 = (w2087 & w2094) | (w2087 & w2108) | (w2094 & w2108);
assign w2110 = pi247 & ~w2109;
assign w2111 = ~pi119 & pi246;
assign w2112 = ~pi120 & pi247;
assign w2113 = (~pi120 & w2111) | (~pi120 & w2112) | (w2111 & w2112);
assign w2114 = ~pi119 & ~pi120;
assign w2115 = ~pi244 & w114;
assign w2116 = w119 & w2115;
assign w2117 = ~w2083 & w2116;
assign w2118 = w1999 & w2117;
assign w2119 = w2114 & ~w2118;
assign w2120 = (~w1739 & w2114) | (~w1739 & w2119) | (w2114 & w2119);
assign w2121 = ~w2113 & ~w2120;
assign w2122 = (w2006 & w2102) | (w2006 & w2105) | (w2102 & w2105);
assign w2123 = w2120 & w2122;
assign w2124 = ~w2113 & ~w2123;
assign w2125 = (~w2094 & w2121) | (~w2094 & w2124) | (w2121 & w2124);
assign w2126 = pi248 & w2125;
assign w2127 = ~pi121 & pi248;
assign w2128 = (~pi121 & w2113) | (~pi121 & w2127) | (w2113 & w2127);
assign w2129 = (~pi121 & w2120) | (~pi121 & w2128) | (w2120 & w2128);
assign w2130 = (~pi121 & w2123) | (~pi121 & w2128) | (w2123 & w2128);
assign w2131 = (w2094 & w2129) | (w2094 & w2130) | (w2129 & w2130);
assign w2132 = pi249 & ~w2131;
assign w2133 = ~pi122 & ~w341;
assign w2134 = ~pi249 & ~w2127;
assign w2135 = (w341 & ~w2113) | (w341 & w2134) | (~w2113 & w2134);
assign w2136 = ~pi122 & ~w2135;
assign w2137 = (w2120 & w2133) | (w2120 & w2136) | (w2133 & w2136);
assign w2138 = (w2123 & w2133) | (w2123 & w2136) | (w2133 & w2136);
assign w2139 = (w2094 & w2137) | (w2094 & w2138) | (w2137 & w2138);
assign w2140 = pi250 & ~w2139;
assign w2141 = ~w113 & w346;
assign w2142 = w114 & w120;
assign w2143 = pi124 & w2142;
assign w2144 = w1999 & w2143;
assign w2145 = ~pi119 & ~w2144;
assign w2146 = (~pi119 & ~w1739) | (~pi119 & w2145) | (~w1739 & w2145);
assign w2147 = (w346 & w2141) | (w346 & w2146) | (w2141 & w2146);
assign w2148 = w1739 & w2144;
assign w2149 = ~pi119 & ~w2107;
assign w2150 = ~w2148 & w2149;
assign w2151 = (w346 & w2141) | (w346 & w2150) | (w2141 & w2150);
assign w2152 = (w2094 & w2147) | (w2094 & w2151) | (w2147 & w2151);
assign w2153 = pi251 & ~w2152;
assign w2154 = pi119 & w336;
assign w2155 = w2083 & ~w2154;
assign w2156 = w336 & ~w2149;
assign w2157 = w2083 & ~w2156;
assign w2158 = (w2094 & w2155) | (w2094 & w2157) | (w2155 & w2157);
assign w2159 = pi252 & ~w2158;
assign w2160 = ~pi127 & ~w316;
assign w2161 = w1134 & ~w2160;
assign w2162 = w1030 & w2161;
assign w2163 = w259 & w2162;
assign w2164 = (w259 & w1157) | (w259 & w2163) | (w1157 & w2163);
assign w2165 = w1041 & w1561;
assign w2166 = ~pi252 & ~w2165;
assign w2167 = (~pi252 & w2164) | (~pi252 & w2166) | (w2164 & w2166);
assign w2168 = ~pi125 & ~w2167;
assign w2169 = pi253 & ~w2168;
assign w2170 = ~pi126 & ~w315;
assign w2171 = (w254 & ~w2167) | (w254 & w2170) | (~w2167 & w2170);
assign w2172 = pi254 & ~w2171;
assign w2173 = w259 & w1157;
assign w2174 = w261 & ~w2165;
assign w2175 = (w261 & w2173) | (w261 & w2174) | (w2173 & w2174);
assign w2176 = w318 & ~w2175;
assign w2177 = pi255 & ~w2176;
assign w2178 = w1045 & w1134;
assign one = 1;
assign po000 = w469;
assign po001 = w479;
assign po002 = w504;
assign po003 = w512;
assign po004 = w531;
assign po005 = w538;
assign po006 = w554;
assign po007 = w583;
assign po008 = w596;
assign po009 = w604;
assign po010 = w614;
assign po011 = w630;
assign po012 = w638;
assign po013 = w648;
assign po014 = w677;
assign po015 = w690;
assign po016 = w704;
assign po017 = w715;
assign po018 = w724;
assign po019 = w762;
assign po020 = w769;
assign po021 = w789;
assign po022 = w796;
assign po023 = w802;
assign po024 = w809;
assign po025 = w827;
assign po026 = w846;
assign po027 = w857;
assign po028 = w874;
assign po029 = w884;
assign po030 = w889;
assign po031 = w900;
assign po032 = w920;
assign po033 = w943;
assign po034 = w949;
assign po035 = w955;
assign po036 = w983;
assign po037 = w1002;
assign po038 = w1010;
assign po039 = w1015;
assign po040 = w1036;
assign po041 = w1039;
assign po042 = w1059;
assign po043 = ~w1067;
assign po044 = w1097;
assign po045 = w1105;
assign po046 = w1118;
assign po047 = w1131;
assign po048 = w1137;
assign po049 = w1171;
assign po050 = w1177;
assign po051 = w1182;
assign po052 = w1186;
assign po053 = w1199;
assign po054 = w1207;
assign po055 = w1224;
assign po056 = w1245;
assign po057 = w1250;
assign po058 = w1257;
assign po059 = w1266;
assign po060 = w1279;
assign po061 = w1297;
assign po062 = w1313;
assign po063 = w1319;
assign po064 = w1329;
assign po065 = w1350;
assign po066 = w1358;
assign po067 = w1373;
assign po068 = w1389;
assign po069 = w1395;
assign po070 = w1407;
assign po071 = w1420;
assign po072 = w1427;
assign po073 = w1444;
assign po074 = w1471;
assign po075 = w1486;
assign po076 = w1494;
assign po077 = w1513;
assign po078 = w1532;
assign po079 = w1538;
assign po080 = w1570;
assign po081 = w1575;
assign po082 = w1591;
assign po083 = w1595;
assign po084 = w1625;
assign po085 = w1640;
assign po086 = w1648;
assign po087 = w1666;
assign po088 = w1673;
assign po089 = w1699;
assign po090 = w1713;
assign po091 = w1715;
assign po092 = w1722;
assign po093 = w1742;
assign po094 = w1748;
assign po095 = w1774;
assign po096 = w1790;
assign po097 = w1793;
assign po098 = w1799;
assign po099 = w1837;
assign po100 = w1842;
assign po101 = w1849;
assign po102 = w1894;
assign po103 = w1910;
assign po104 = w1914;
assign po105 = w1925;
assign po106 = w1944;
assign po107 = w1954;
assign po108 = w1972;
assign po109 = w1981;
assign po110 = w1988;
assign po111 = w1994;
assign po112 = w2020;
assign po113 = w2041;
assign po114 = w2048;
assign po115 = w2058;
assign po116 = w2065;
assign po117 = w2071;
assign po118 = w2080;
assign po119 = w2110;
assign po120 = w2126;
assign po121 = w2132;
assign po122 = w2140;
assign po123 = w2153;
assign po124 = w2159;
assign po125 = w2169;
assign po126 = w2172;
assign po127 = w2177;
assign po128 = ~w2178;
endmodule

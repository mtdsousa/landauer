// Benchmark "k2" written by ABC on Sun Apr 22 21:43:06 2018

module k2 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n136, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n431, n432, n433, n434, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n449, n450,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n572, n573, n574, n575, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088,
    n1089, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1395, n1396, n1397, n1398, n1399, n1401, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1433, n1434, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1551,
    n1552, n1553, n1554, n1556, n1557, n1558, n1560, n1561, n1562, n1563,
    n1564, n1565, n1567, n1568, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2084, n2085, n2086, n2087, n2088;
  assign n92 = ~pi00 & ~pi18;
  assign n93 = ~pi19 & n92;
  assign n94 = pi20 & n93;
  assign n95 = pi21 & n94;
  assign n96 = pi24 & n95;
  assign n97 = ~pi29 & n96;
  assign n98 = pi30 & n97;
  assign n99 = ~pi18 & pi19;
  assign n100 = pi21 & n99;
  assign n101 = pi24 & n100;
  assign n102 = ~pi28 & n101;
  assign n103 = ~pi29 & n102;
  assign n104 = pi30 & n103;
  assign n105 = pi10 & ~pi18;
  assign n106 = pi19 & n105;
  assign n107 = pi21 & n106;
  assign n108 = pi25 & n107;
  assign n109 = ~pi28 & n108;
  assign n110 = ~pi29 & n109;
  assign n111 = pi30 & n110;
  assign n112 = pi26 & n100;
  assign n113 = ~pi28 & n112;
  assign n114 = ~pi29 & n113;
  assign n115 = pi30 & n114;
  assign n116 = ~pi00 & pi18;
  assign n117 = ~pi19 & n116;
  assign n118 = ~pi20 & n117;
  assign n119 = pi21 & n118;
  assign n120 = ~pi28 & n119;
  assign n121 = ~pi29 & n120;
  assign n122 = pi30 & n121;
  assign n123 = pi19 & n116;
  assign n124 = pi20 & n123;
  assign n125 = pi21 & n124;
  assign n126 = pi24 & n125;
  assign n127 = ~pi29 & n126;
  assign n128 = pi30 & n127;
  assign n129 = ~n115 & ~n122;
  assign n130 = ~n128 & n129;
  assign n131 = ~n98 & ~n104;
  assign n132 = ~n111 & n131;
  assign po00 = ~n130 | ~n132;
  assign po01 = n98 | n128;
  assign po03 = n111 | n115;
  assign n136 = ~n104 & ~n115;
  assign po04 = n128 | ~n136;
  assign n138 = pi00 & ~pi18;
  assign n139 = ~pi19 & n138;
  assign n140 = pi20 & n139;
  assign n141 = pi21 & n140;
  assign n142 = pi24 & n141;
  assign n143 = ~pi29 & n142;
  assign n144 = pi30 & n143;
  assign n145 = pi19 & n138;
  assign n146 = pi21 & n145;
  assign n147 = pi28 & n146;
  assign n148 = ~pi29 & n147;
  assign n149 = pi30 & n148;
  assign n150 = pi00 & pi18;
  assign n151 = ~pi19 & n150;
  assign n152 = ~pi20 & n151;
  assign n153 = pi21 & n152;
  assign n154 = ~pi28 & n153;
  assign n155 = ~pi29 & n154;
  assign n156 = pi30 & n155;
  assign n157 = pi19 & n150;
  assign n158 = pi20 & n157;
  assign n159 = pi21 & n158;
  assign n160 = ~pi29 & n159;
  assign n161 = pi30 & n160;
  assign n162 = ~n144 & ~n149;
  assign n163 = ~n156 & ~n161;
  assign po05 = ~n162 | ~n163;
  assign n165 = pi22 & n141;
  assign n166 = ~pi29 & n165;
  assign n167 = pi30 & n166;
  assign n168 = pi00 & pi10;
  assign n169 = ~pi11 & n168;
  assign n170 = ~pi18 & n169;
  assign n171 = ~pi19 & n170;
  assign n172 = pi20 & n171;
  assign n173 = pi21 & n172;
  assign n174 = pi25 & n173;
  assign n175 = ~pi29 & n174;
  assign n176 = pi30 & n175;
  assign n177 = pi11 & n168;
  assign n178 = ~pi18 & n177;
  assign n179 = ~pi19 & n178;
  assign n180 = pi20 & n179;
  assign n181 = pi21 & n180;
  assign n182 = pi25 & n181;
  assign n183 = ~pi29 & n182;
  assign n184 = pi30 & n183;
  assign n185 = pi00 & ~pi11;
  assign n186 = ~pi18 & n185;
  assign n187 = ~pi19 & n186;
  assign n188 = pi20 & n187;
  assign n189 = pi21 & n188;
  assign n190 = pi26 & n189;
  assign n191 = ~pi29 & n190;
  assign n192 = pi30 & n191;
  assign n193 = pi00 & pi11;
  assign n194 = ~pi18 & n193;
  assign n195 = ~pi19 & n194;
  assign n196 = pi20 & n195;
  assign n197 = pi21 & n196;
  assign n198 = pi26 & n197;
  assign n199 = ~pi29 & n198;
  assign n200 = pi30 & n199;
  assign n201 = pi00 & ~pi05;
  assign n202 = ~pi15 & n201;
  assign n203 = ~pi18 & n202;
  assign n204 = pi19 & n203;
  assign n205 = pi20 & n204;
  assign n206 = pi21 & n205;
  assign n207 = pi22 & n206;
  assign n208 = ~pi28 & n207;
  assign n209 = ~pi29 & n208;
  assign po41 = pi30 & n209;
  assign n211 = pi18 & n202;
  assign n212 = ~pi19 & n211;
  assign n213 = pi20 & n212;
  assign n214 = pi21 & n213;
  assign n215 = pi22 & n214;
  assign n216 = ~pi28 & n215;
  assign n217 = ~pi29 & n216;
  assign n218 = pi30 & n217;
  assign n219 = pi10 & n201;
  assign n220 = ~pi11 & n219;
  assign n221 = ~pi15 & n220;
  assign n222 = pi18 & n221;
  assign n223 = ~pi19 & n222;
  assign n224 = pi20 & n223;
  assign n225 = pi21 & n224;
  assign n226 = pi25 & n225;
  assign n227 = ~pi28 & n226;
  assign n228 = ~pi29 & n227;
  assign n229 = pi30 & n228;
  assign n230 = pi11 & n219;
  assign n231 = ~pi15 & n230;
  assign n232 = pi18 & n231;
  assign n233 = ~pi19 & n232;
  assign n234 = pi20 & n233;
  assign n235 = pi21 & n234;
  assign n236 = pi25 & n235;
  assign n237 = ~pi28 & n236;
  assign n238 = ~pi29 & n237;
  assign n239 = pi30 & n238;
  assign n240 = ~pi11 & n201;
  assign n241 = ~pi15 & n240;
  assign n242 = pi18 & n241;
  assign n243 = ~pi19 & n242;
  assign n244 = pi20 & n243;
  assign n245 = pi21 & n244;
  assign n246 = pi26 & n245;
  assign n247 = ~pi28 & n246;
  assign n248 = ~pi29 & n247;
  assign n249 = pi30 & n248;
  assign n250 = pi11 & n201;
  assign n251 = ~pi15 & n250;
  assign n252 = pi18 & n251;
  assign n253 = ~pi19 & n252;
  assign n254 = pi20 & n253;
  assign n255 = pi21 & n254;
  assign n256 = pi26 & n255;
  assign n257 = ~pi28 & n256;
  assign n258 = ~pi29 & n257;
  assign n259 = pi30 & n258;
  assign n260 = pi00 & ~pi03;
  assign n261 = ~pi05 & n260;
  assign n262 = ~pi18 & n261;
  assign n263 = ~pi19 & n262;
  assign n264 = ~pi20 & n263;
  assign n265 = ~pi21 & n264;
  assign n266 = ~pi28 & n265;
  assign n267 = pi29 & n266;
  assign n268 = ~pi30 & n267;
  assign n269 = pi00 & pi02;
  assign n270 = ~pi03 & n269;
  assign n271 = ~pi18 & n270;
  assign n272 = ~pi19 & n271;
  assign n273 = ~pi20 & n272;
  assign n274 = ~pi21 & n273;
  assign n275 = pi28 & n274;
  assign n276 = ~pi29 & n275;
  assign n277 = pi30 & n276;
  assign n278 = ~pi21 & n140;
  assign n279 = pi23 & n278;
  assign n280 = ~pi28 & n279;
  assign n281 = pi29 & n280;
  assign n282 = ~pi30 & n281;
  assign n283 = pi00 & ~pi02;
  assign n284 = ~pi03 & n283;
  assign n285 = ~pi18 & n284;
  assign n286 = ~pi19 & n285;
  assign n287 = pi20 & n286;
  assign n288 = ~pi21 & n287;
  assign n289 = pi28 & n288;
  assign n290 = ~pi29 & n289;
  assign n291 = pi30 & n290;
  assign n292 = ~pi18 & n201;
  assign n293 = pi19 & n292;
  assign n294 = pi20 & n293;
  assign n295 = ~pi21 & n294;
  assign n296 = pi22 & n295;
  assign n297 = ~pi28 & n296;
  assign n298 = pi29 & n297;
  assign n299 = ~pi30 & n298;
  assign n300 = pi20 & n145;
  assign n301 = ~pi21 & n300;
  assign n302 = pi22 & n301;
  assign n303 = pi28 & n302;
  assign n304 = pi29 & n303;
  assign n305 = ~pi30 & n304;
  assign n306 = pi00 & pi17;
  assign n307 = pi18 & n306;
  assign n308 = ~pi19 & n307;
  assign n309 = pi20 & n308;
  assign n310 = ~pi21 & n309;
  assign n311 = pi26 & n310;
  assign n312 = ~pi28 & n311;
  assign n313 = pi29 & n312;
  assign n314 = ~pi30 & n313;
  assign n315 = pi00 & ~pi17;
  assign n316 = pi18 & n315;
  assign n317 = ~pi19 & n316;
  assign n318 = pi20 & n317;
  assign n319 = ~pi21 & n318;
  assign n320 = pi26 & n319;
  assign n321 = ~pi28 & n320;
  assign n322 = pi29 & n321;
  assign n323 = ~pi30 & n322;
  assign n324 = pi18 & n185;
  assign n325 = ~pi19 & n324;
  assign n326 = pi20 & n325;
  assign n327 = ~pi21 & n326;
  assign n328 = pi26 & n327;
  assign n329 = pi28 & n328;
  assign n330 = ~pi29 & n329;
  assign n331 = pi30 & n330;
  assign n332 = pi18 & n193;
  assign n333 = ~pi19 & n332;
  assign n334 = pi20 & n333;
  assign n335 = ~pi21 & n334;
  assign n336 = pi26 & n335;
  assign n337 = pi28 & n336;
  assign n338 = ~pi29 & n337;
  assign n339 = pi30 & n338;
  assign n340 = ~pi20 & n157;
  assign n341 = ~pi21 & n340;
  assign n342 = pi22 & n341;
  assign n343 = pi29 & n342;
  assign n344 = ~pi30 & n343;
  assign n345 = pi18 & n177;
  assign n346 = pi19 & n345;
  assign n347 = ~pi20 & n346;
  assign n348 = ~pi21 & n347;
  assign n349 = pi25 & n348;
  assign n350 = pi29 & n349;
  assign n351 = ~pi30 & n350;
  assign n352 = pi18 & n169;
  assign n353 = pi19 & n352;
  assign n354 = ~pi20 & n353;
  assign n355 = ~pi21 & n354;
  assign n356 = pi25 & n355;
  assign n357 = pi29 & n356;
  assign n358 = ~pi30 & n357;
  assign n359 = pi26 & n341;
  assign n360 = ~pi28 & n359;
  assign n361 = pi29 & n360;
  assign n362 = ~pi30 & n361;
  assign n363 = pi19 & n332;
  assign n364 = ~pi20 & n363;
  assign n365 = ~pi21 & n364;
  assign n366 = pi26 & n365;
  assign n367 = pi28 & n366;
  assign n368 = ~pi29 & n367;
  assign n369 = pi30 & n368;
  assign n370 = pi19 & n324;
  assign n371 = ~pi20 & n370;
  assign n372 = ~pi21 & n371;
  assign n373 = pi26 & n372;
  assign n374 = pi28 & n373;
  assign n375 = ~pi29 & n374;
  assign n376 = pi30 & n375;
  assign n377 = pi18 & n201;
  assign n378 = pi19 & n377;
  assign n379 = pi20 & n378;
  assign n380 = ~pi21 & n379;
  assign n381 = ~pi27 & n380;
  assign n382 = ~pi28 & n381;
  assign n383 = pi29 & n382;
  assign n384 = pi30 & n383;
  assign n385 = ~pi00 & ~pi04;
  assign n386 = pi18 & n385;
  assign n387 = pi19 & n386;
  assign n388 = pi20 & n387;
  assign n389 = ~pi21 & n388;
  assign n390 = ~pi27 & n389;
  assign n391 = pi28 & n390;
  assign n392 = pi29 & n391;
  assign n393 = ~pi30 & n392;
  assign n394 = pi00 & pi03;
  assign n395 = pi18 & n394;
  assign n396 = pi19 & n395;
  assign n397 = pi20 & n396;
  assign n398 = ~pi21 & n397;
  assign n399 = pi27 & n398;
  assign n400 = ~pi29 & n399;
  assign n401 = ~pi30 & n400;
  assign n402 = ~n384 & ~n393;
  assign n403 = ~n401 & n402;
  assign n404 = ~n369 & ~n376;
  assign n405 = ~n358 & ~n362;
  assign n406 = n404 & n405;
  assign n407 = n403 & n406;
  assign n408 = ~n344 & ~n351;
  assign n409 = ~n331 & ~n339;
  assign n410 = n408 & n409;
  assign n411 = ~n314 & ~n323;
  assign n412 = ~n299 & ~n305;
  assign n413 = n411 & n412;
  assign n414 = n410 & n413;
  assign n415 = n407 & n414;
  assign n416 = ~n277 & ~n282;
  assign n417 = ~n291 & n416;
  assign n418 = ~n259 & ~n268;
  assign n419 = ~n239 & ~n249;
  assign n420 = n418 & n419;
  assign n421 = n417 & n420;
  assign n422 = ~n167 & ~n176;
  assign n423 = ~n184 & ~n192;
  assign n424 = n422 & n423;
  assign n425 = ~n218 & ~n229;
  assign n426 = ~n200 & ~po41;
  assign n427 = n425 & n426;
  assign n428 = n424 & n427;
  assign n429 = n421 & n428;
  assign po06 = ~n415 | ~n429;
  assign n431 = ~n239 & ~n351;
  assign n432 = ~n358 & n431;
  assign n433 = ~n176 & ~n184;
  assign n434 = ~n229 & n433;
  assign po07 = ~n432 | ~n434;
  assign n436 = ~n358 & ~n376;
  assign n437 = ~n393 & n436;
  assign n438 = ~n339 & ~n344;
  assign n439 = ~n291 & ~n305;
  assign n440 = n438 & n439;
  assign n441 = n437 & n440;
  assign n442 = ~n192 & ~po41;
  assign n443 = n422 & n442;
  assign n444 = ~n249 & ~n268;
  assign n445 = n425 & n444;
  assign n446 = n443 & n445;
  assign po08 = ~n441 | ~n446;
  assign po09 = n401 | ~n416;
  assign n449 = ~pi18 & ~pi19;
  assign n450 = pi20 & n449;
  assign n451 = pi21 & n450;
  assign n452 = ~pi26 & n451;
  assign n453 = pi29 & n452;
  assign n454 = ~pi30 & n453;
  assign n455 = pi26 & n451;
  assign n456 = pi29 & n455;
  assign n457 = ~pi30 & n456;
  assign n458 = pi30 & n456;
  assign n459 = pi24 & n451;
  assign n460 = pi29 & n459;
  assign n461 = ~pi30 & n460;
  assign n462 = pi01 & ~pi18;
  assign n463 = pi19 & n462;
  assign n464 = ~pi20 & n463;
  assign n465 = pi21 & n464;
  assign n466 = pi22 & n465;
  assign n467 = ~pi28 & n466;
  assign n468 = ~pi29 & n467;
  assign n469 = pi30 & n468;
  assign n470 = pi23 & n465;
  assign n471 = ~pi28 & n470;
  assign n472 = ~pi29 & n471;
  assign n473 = pi30 & n472;
  assign n474 = pi28 & n100;
  assign n475 = pi29 & n474;
  assign n476 = ~pi30 & n475;
  assign n477 = pi20 & n99;
  assign n478 = pi21 & n477;
  assign n479 = pi22 & n478;
  assign n480 = ~pi28 & n479;
  assign n481 = pi29 & n480;
  assign n482 = ~pi30 & n481;
  assign n483 = pi18 & ~pi19;
  assign n484 = ~pi20 & n483;
  assign n485 = pi21 & n484;
  assign n486 = ~pi28 & n485;
  assign n487 = pi29 & n486;
  assign n488 = ~pi30 & n487;
  assign n489 = pi20 & n483;
  assign n490 = pi21 & n489;
  assign n491 = pi22 & n490;
  assign n492 = ~pi28 & n491;
  assign n493 = pi29 & n492;
  assign n494 = ~pi30 & n493;
  assign n495 = ~pi11 & pi18;
  assign n496 = ~pi19 & n495;
  assign n497 = pi20 & n496;
  assign n498 = pi21 & n497;
  assign n499 = pi25 & n498;
  assign n500 = ~pi28 & n499;
  assign n501 = pi29 & n500;
  assign n502 = ~pi30 & n501;
  assign n503 = pi11 & pi18;
  assign n504 = ~pi19 & n503;
  assign n505 = pi20 & n504;
  assign n506 = pi21 & n505;
  assign n507 = pi25 & n506;
  assign n508 = ~pi28 & n507;
  assign n509 = pi29 & n508;
  assign n510 = ~pi30 & n509;
  assign n511 = pi26 & n498;
  assign n512 = ~pi28 & n511;
  assign n513 = pi29 & n512;
  assign n514 = ~pi30 & n513;
  assign n515 = pi30 & n513;
  assign n516 = pi26 & n506;
  assign n517 = ~pi28 & n516;
  assign n518 = pi29 & n517;
  assign n519 = ~pi30 & n518;
  assign n520 = pi30 & n518;
  assign n521 = pi18 & pi19;
  assign n522 = pi20 & n521;
  assign n523 = pi21 & n522;
  assign n524 = pi29 & n523;
  assign n525 = ~pi30 & n524;
  assign n526 = ~pi20 & n449;
  assign n527 = ~pi21 & n526;
  assign n528 = ~pi28 & n527;
  assign n529 = pi29 & n528;
  assign n530 = pi30 & n529;
  assign n531 = pi28 & n527;
  assign n532 = pi29 & n531;
  assign n533 = ~pi30 & n532;
  assign n534 = ~pi21 & n450;
  assign n535 = ~pi28 & n534;
  assign n536 = pi29 & n535;
  assign n537 = pi30 & n536;
  assign n538 = pi28 & n534;
  assign n539 = pi29 & n538;
  assign n540 = ~pi30 & n539;
  assign n541 = ~pi21 & n464;
  assign n542 = pi22 & n541;
  assign n543 = pi29 & n542;
  assign n544 = ~pi30 & n543;
  assign n545 = pi23 & n541;
  assign n546 = pi29 & n545;
  assign n547 = ~pi30 & n546;
  assign n548 = ~pi21 & n477;
  assign n549 = pi22 & n548;
  assign n550 = ~pi28 & n549;
  assign n551 = pi29 & n550;
  assign n552 = pi30 & n551;
  assign n553 = pi28 & n549;
  assign n554 = pi29 & n553;
  assign n555 = pi30 & n554;
  assign n556 = pi17 & pi18;
  assign n557 = ~pi19 & n556;
  assign n558 = pi20 & n557;
  assign n559 = ~pi21 & n558;
  assign n560 = pi26 & n559;
  assign n561 = ~pi28 & n560;
  assign n562 = pi29 & n561;
  assign n563 = ~pi30 & n562;
  assign n564 = ~pi17 & pi18;
  assign n565 = ~pi19 & n564;
  assign n566 = pi20 & n565;
  assign n567 = ~pi21 & n566;
  assign n568 = pi26 & n567;
  assign n569 = ~pi28 & n568;
  assign n570 = pi29 & n569;
  assign po20 = pi30 & n570;
  assign n572 = ~pi21 & n489;
  assign n573 = pi26 & n572;
  assign n574 = pi28 & n573;
  assign n575 = pi29 & n574;
  assign po21 = ~pi30 & n575;
  assign n577 = ~pi20 & n521;
  assign n578 = ~pi21 & n577;
  assign n579 = pi22 & n578;
  assign n580 = pi29 & n579;
  assign n581 = pi30 & n580;
  assign n582 = pi25 & n578;
  assign n583 = pi29 & n582;
  assign n584 = pi30 & n583;
  assign n585 = pi26 & n578;
  assign n586 = ~pi28 & n585;
  assign n587 = pi29 & n586;
  assign n588 = pi30 & n587;
  assign n589 = pi28 & n585;
  assign n590 = pi29 & n589;
  assign n591 = ~pi30 & n590;
  assign n592 = ~pi21 & n522;
  assign n593 = ~pi27 & n592;
  assign n594 = pi28 & n593;
  assign n595 = ~pi29 & n594;
  assign n596 = ~pi30 & n595;
  assign n597 = pi29 & n594;
  assign n598 = pi30 & n597;
  assign n599 = pi27 & n592;
  assign n600 = ~pi29 & n599;
  assign n601 = pi30 & n600;
  assign n602 = ~pi09 & ~pi18;
  assign n603 = ~pi19 & n602;
  assign n604 = ~pi20 & n603;
  assign n605 = pi21 & n604;
  assign n606 = pi22 & n605;
  assign n607 = ~pi28 & n606;
  assign n608 = ~pi29 & n607;
  assign n609 = pi30 & n608;
  assign n610 = pi09 & ~pi18;
  assign n611 = ~pi19 & n610;
  assign n612 = ~pi20 & n611;
  assign n613 = pi21 & n612;
  assign n614 = pi22 & n613;
  assign n615 = ~pi28 & n614;
  assign n616 = ~pi29 & n615;
  assign n617 = pi30 & n616;
  assign n618 = ~pi31 & n617;
  assign n619 = ~pi33 & n618;
  assign n620 = pi39 & n619;
  assign n621 = pi29 & n607;
  assign n622 = ~pi30 & n621;
  assign n623 = pi38 & n622;
  assign n624 = ~pi38 & n622;
  assign n625 = pi41 & n624;
  assign n626 = ~pi39 & n624;
  assign n627 = ~pi41 & n626;
  assign n628 = pi42 & n627;
  assign n629 = pi39 & n624;
  assign n630 = ~pi41 & n629;
  assign n631 = ~pi42 & n630;
  assign n632 = pi42 & n630;
  assign n633 = pi21 & n526;
  assign n634 = pi22 & n633;
  assign n635 = ~pi28 & n634;
  assign n636 = pi29 & n635;
  assign n637 = pi30 & n636;
  assign n638 = ~pi40 & n626;
  assign n639 = ~pi41 & n638;
  assign n640 = ~pi42 & n639;
  assign n641 = ~pi43 & n640;
  assign n642 = pi44 & n641;
  assign n643 = ~n637 & ~n642;
  assign n644 = ~n628 & ~n631;
  assign n645 = ~n632 & n644;
  assign n646 = n643 & n645;
  assign n647 = ~n620 & ~n623;
  assign n648 = ~n625 & n647;
  assign n649 = ~n598 & ~n601;
  assign n650 = ~n609 & n649;
  assign n651 = n648 & n650;
  assign n652 = n646 & n651;
  assign n653 = ~n591 & ~n596;
  assign n654 = ~n581 & ~n584;
  assign n655 = ~n588 & n654;
  assign n656 = n653 & n655;
  assign n657 = ~n563 & ~po20;
  assign n658 = ~po21 & n657;
  assign n659 = ~n547 & ~n552;
  assign n660 = ~n555 & n659;
  assign n661 = n658 & n660;
  assign n662 = n656 & n661;
  assign n663 = n652 & n662;
  assign n664 = ~n540 & ~n544;
  assign n665 = ~n530 & ~n533;
  assign n666 = ~n537 & n665;
  assign n667 = n664 & n666;
  assign n668 = ~n519 & ~n520;
  assign n669 = ~n525 & n668;
  assign n670 = ~n510 & ~n514;
  assign n671 = ~n515 & n670;
  assign n672 = n669 & n671;
  assign n673 = n667 & n672;
  assign n674 = ~n461 & ~n469;
  assign n675 = ~n473 & n674;
  assign n676 = ~n454 & ~n457;
  assign n677 = ~n458 & n676;
  assign n678 = n675 & n677;
  assign n679 = ~n494 & ~n502;
  assign n680 = ~n476 & ~n482;
  assign n681 = ~n488 & n680;
  assign n682 = n679 & n681;
  assign n683 = n678 & n682;
  assign n684 = n673 & n683;
  assign po10 = ~n663 | ~n684;
  assign n686 = pi30 & n453;
  assign n687 = pi30 & n460;
  assign n688 = ~pi20 & n99;
  assign n689 = pi21 & n688;
  assign n690 = pi22 & n689;
  assign n691 = ~pi28 & n690;
  assign n692 = pi29 & n691;
  assign n693 = ~pi30 & n692;
  assign n694 = pi23 & n689;
  assign n695 = ~pi28 & n694;
  assign n696 = pi29 & n695;
  assign n697 = ~pi30 & n696;
  assign n698 = pi30 & n475;
  assign n699 = pi30 & n481;
  assign n700 = pi30 & n487;
  assign n701 = pi30 & n493;
  assign n702 = pi30 & n501;
  assign n703 = pi30 & n509;
  assign n704 = pi28 & n560;
  assign n705 = ~pi29 & n704;
  assign n706 = ~pi30 & n705;
  assign n707 = ~pi29 & n589;
  assign n708 = ~pi30 & n707;
  assign n709 = ~pi03 & pi18;
  assign n710 = pi19 & n709;
  assign n711 = pi20 & n710;
  assign n712 = ~pi21 & n711;
  assign n713 = pi27 & n712;
  assign n714 = ~pi29 & n713;
  assign n715 = ~pi30 & n714;
  assign n716 = pi43 & n640;
  assign n717 = ~pi44 & n716;
  assign n718 = ~n601 & ~n717;
  assign n719 = ~n596 & ~n715;
  assign n720 = n718 & n719;
  assign n721 = ~n588 & ~n708;
  assign n722 = ~n552 & ~n563;
  assign n723 = ~n706 & n722;
  assign n724 = n721 & n723;
  assign n725 = n720 & n724;
  assign n726 = ~n537 & ~n540;
  assign n727 = ~n525 & ~n530;
  assign n728 = ~n533 & n727;
  assign n729 = n726 & n728;
  assign n730 = ~n514 & ~n703;
  assign n731 = ~n515 & n730;
  assign n732 = n668 & n731;
  assign n733 = n729 & n732;
  assign n734 = n725 & n733;
  assign n735 = ~n502 & ~n702;
  assign n736 = ~n494 & ~n700;
  assign n737 = ~n701 & n736;
  assign n738 = n735 & n737;
  assign n739 = ~n488 & ~n699;
  assign n740 = ~n476 & ~n698;
  assign n741 = ~n482 & n740;
  assign n742 = n739 & n741;
  assign n743 = n738 & n742;
  assign n744 = ~n693 & ~n697;
  assign n745 = ~n469 & ~n687;
  assign n746 = ~n473 & n745;
  assign n747 = n744 & n746;
  assign n748 = ~n458 & ~n461;
  assign n749 = ~n454 & ~n686;
  assign n750 = ~n457 & n749;
  assign n751 = n748 & n750;
  assign n752 = n747 & n751;
  assign n753 = n743 & n752;
  assign po11 = ~n734 | ~n753;
  assign n755 = pi10 & pi18;
  assign n756 = pi19 & n755;
  assign n757 = ~pi20 & n756;
  assign n758 = pi21 & n757;
  assign n759 = pi25 & n758;
  assign n760 = pi30 & n759;
  assign n761 = pi21 & n577;
  assign n762 = pi26 & n761;
  assign n763 = pi30 & n762;
  assign n764 = pi30 & n524;
  assign n765 = ~pi44 & n641;
  assign n766 = ~n609 & ~n642;
  assign n767 = ~n765 & n766;
  assign n768 = ~n598 & ~n715;
  assign n769 = ~n601 & n768;
  assign n770 = n767 & n769;
  assign n771 = ~n591 & ~n708;
  assign n772 = ~n596 & n771;
  assign n773 = ~po21 & ~n581;
  assign n774 = ~n584 & ~n588;
  assign n775 = n773 & n774;
  assign n776 = n772 & n775;
  assign n777 = n770 & n776;
  assign n778 = ~n563 & ~n706;
  assign n779 = ~po20 & n778;
  assign n780 = n660 & n779;
  assign n781 = ~n544 & n726;
  assign n782 = ~n525 & ~n764;
  assign n783 = n665 & n782;
  assign n784 = n781 & n783;
  assign n785 = n780 & n784;
  assign n786 = n777 & n785;
  assign n787 = ~n514 & ~n515;
  assign n788 = ~n519 & n787;
  assign n789 = ~n520 & ~n760;
  assign n790 = ~n763 & n789;
  assign n791 = n788 & n790;
  assign n792 = ~n510 & ~n702;
  assign n793 = ~n703 & n792;
  assign n794 = ~n502 & ~n701;
  assign n795 = n736 & n794;
  assign n796 = n793 & n795;
  assign n797 = n791 & n796;
  assign n798 = ~n482 & ~n699;
  assign n799 = ~n488 & n798;
  assign n800 = ~n476 & ~n697;
  assign n801 = ~n698 & n800;
  assign n802 = n799 & n801;
  assign n803 = ~n457 & ~n458;
  assign n804 = n749 & n803;
  assign n805 = ~n461 & ~n687;
  assign n806 = ~n693 & n805;
  assign n807 = n804 & n806;
  assign n808 = n802 & n807;
  assign n809 = n797 & n808;
  assign po12 = ~n786 | ~n809;
  assign n811 = pi14 & ~pi27;
  assign n812 = ~pi28 & n811;
  assign n813 = ~pi29 & n812;
  assign n814 = ~pi30 & n813;
  assign n815 = pi13 & ~pi14;
  assign n816 = pi21 & n815;
  assign n817 = ~pi27 & n816;
  assign n818 = ~pi28 & n817;
  assign n819 = ~pi29 & n818;
  assign n820 = ~pi30 & n819;
  assign n821 = ~pi29 & n528;
  assign n822 = pi30 & n821;
  assign n823 = pi23 & n534;
  assign n824 = ~pi28 & n823;
  assign n825 = ~pi29 & n824;
  assign n826 = pi30 & n825;
  assign n827 = ~pi21 & n688;
  assign n828 = pi22 & n827;
  assign n829 = ~pi29 & n828;
  assign n830 = pi30 & n829;
  assign n831 = pi23 & n827;
  assign n832 = ~pi29 & n831;
  assign n833 = pi30 & n832;
  assign n834 = ~pi29 & n550;
  assign n835 = pi30 & n834;
  assign n836 = pi23 & n548;
  assign n837 = ~pi28 & n836;
  assign n838 = ~pi29 & n837;
  assign n839 = pi30 & n838;
  assign n840 = pi26 & n548;
  assign n841 = ~pi28 & n840;
  assign n842 = ~pi29 & n841;
  assign n843 = pi30 & n842;
  assign n844 = pi03 & ~pi18;
  assign n845 = pi19 & n844;
  assign n846 = pi20 & n845;
  assign n847 = ~pi21 & n846;
  assign n848 = pi22 & n847;
  assign n849 = pi28 & n848;
  assign n850 = ~pi29 & n849;
  assign n851 = pi30 & n850;
  assign n852 = ~pi02 & ~pi03;
  assign n853 = ~pi18 & n852;
  assign n854 = pi19 & n853;
  assign n855 = pi20 & n854;
  assign n856 = ~pi21 & n855;
  assign n857 = pi22 & n856;
  assign n858 = pi28 & n857;
  assign n859 = ~pi29 & n858;
  assign n860 = pi30 & n859;
  assign n861 = pi22 & n572;
  assign n862 = pi30 & n861;
  assign n863 = pi23 & n572;
  assign n864 = pi30 & n863;
  assign n865 = ~pi29 & n561;
  assign n866 = pi30 & n865;
  assign n867 = ~pi29 & n569;
  assign n868 = pi30 & n867;
  assign n869 = ~pi29 & n579;
  assign n870 = pi30 & n869;
  assign n871 = ~pi21 & n757;
  assign n872 = pi25 & n871;
  assign n873 = ~pi29 & n872;
  assign n874 = pi30 & n873;
  assign n875 = ~pi29 & n586;
  assign n876 = pi30 & n875;
  assign n877 = ~pi28 & n593;
  assign n878 = ~pi29 & n877;
  assign n879 = pi30 & n878;
  assign n880 = ~n862 & ~n864;
  assign n881 = ~n555 & ~n851;
  assign n882 = ~n860 & n881;
  assign n883 = n880 & n882;
  assign n884 = ~n835 & ~n839;
  assign n885 = ~n843 & n884;
  assign n886 = ~n544 & ~n833;
  assign n887 = ~n547 & n886;
  assign n888 = n885 & n887;
  assign n889 = n883 & n888;
  assign n890 = ~n473 & ~n510;
  assign n891 = ~n760 & n890;
  assign n892 = ~n814 & ~n820;
  assign n893 = ~n469 & n892;
  assign n894 = n891 & n893;
  assign n895 = ~n826 & ~n830;
  assign n896 = ~n763 & ~n764;
  assign n897 = ~n822 & n896;
  assign n898 = n895 & n897;
  assign n899 = n894 & n898;
  assign n900 = n889 & n899;
  assign n901 = ~n708 & ~n876;
  assign n902 = ~n581 & ~n874;
  assign n903 = ~n584 & n902;
  assign n904 = n901 & n903;
  assign n905 = ~po20 & ~po21;
  assign n906 = ~n870 & n905;
  assign n907 = ~n866 & ~n868;
  assign n908 = ~n706 & n907;
  assign n909 = n906 & n908;
  assign n910 = n904 & n909;
  assign n911 = ~n620 & ~n715;
  assign n912 = ~n591 & ~n879;
  assign n913 = ~n598 & n912;
  assign n914 = n911 & n913;
  assign n915 = n646 & n914;
  assign n916 = n910 & n915;
  assign po13 = ~n900 | ~n916;
  assign n918 = pi33 & n617;
  assign n919 = pi40 & n626;
  assign n920 = ~pi41 & n919;
  assign n921 = ~pi42 & n920;
  assign n922 = ~n631 & ~n637;
  assign n923 = ~n921 & n922;
  assign n924 = ~n620 & ~n625;
  assign n925 = ~n715 & ~n918;
  assign n926 = n924 & n925;
  assign n927 = n923 & n926;
  assign n928 = ~n598 & n771;
  assign n929 = n654 & n905;
  assign n930 = n928 & n929;
  assign n931 = n927 & n930;
  assign n932 = ~n458 & ~n473;
  assign n933 = ~n698 & ~n699;
  assign n934 = n932 & n933;
  assign n935 = ~n510 & ~n515;
  assign n936 = ~n520 & n935;
  assign n937 = n934 & n936;
  assign n938 = ~n555 & ~n860;
  assign n939 = ~n706 & n938;
  assign n940 = ~n547 & ~n851;
  assign n941 = ~n544 & ~n763;
  assign n942 = n940 & n941;
  assign n943 = n939 & n942;
  assign n944 = n937 & n943;
  assign po14 = ~n931 | ~n944;
  assign n946 = pi28 & n485;
  assign n947 = ~pi29 & n946;
  assign n948 = ~pi30 & n947;
  assign n949 = ~pi19 & n844;
  assign n950 = ~pi20 & n949;
  assign n951 = ~pi21 & n950;
  assign n952 = ~pi28 & n951;
  assign n953 = pi29 & n952;
  assign n954 = ~pi30 & n953;
  assign n955 = ~pi03 & pi05;
  assign n956 = ~pi18 & n955;
  assign n957 = ~pi19 & n956;
  assign n958 = ~pi20 & n957;
  assign n959 = ~pi21 & n958;
  assign n960 = ~pi28 & n959;
  assign n961 = pi29 & n960;
  assign n962 = ~pi30 & n961;
  assign n963 = pi24 & n534;
  assign n964 = ~pi29 & n963;
  assign n965 = pi30 & n964;
  assign n966 = pi03 & pi06;
  assign n967 = ~pi18 & n966;
  assign n968 = ~pi19 & n967;
  assign n969 = pi20 & n968;
  assign n970 = ~pi21 & n969;
  assign n971 = pi28 & n970;
  assign n972 = ~pi29 & n971;
  assign n973 = pi30 & n972;
  assign n974 = pi06 & n852;
  assign n975 = ~pi18 & n974;
  assign n976 = ~pi19 & n975;
  assign n977 = pi20 & n976;
  assign n978 = ~pi21 & n977;
  assign n979 = pi28 & n978;
  assign n980 = ~pi29 & n979;
  assign n981 = pi30 & n980;
  assign n982 = pi05 & ~pi18;
  assign n983 = pi19 & n982;
  assign n984 = pi20 & n983;
  assign n985 = ~pi21 & n984;
  assign n986 = pi22 & n985;
  assign n987 = ~pi28 & n986;
  assign n988 = pi29 & n987;
  assign n989 = ~pi30 & n988;
  assign n990 = pi02 & ~pi03;
  assign n991 = ~pi18 & n990;
  assign n992 = pi19 & n991;
  assign n993 = pi20 & n992;
  assign n994 = ~pi21 & n993;
  assign n995 = pi22 & n994;
  assign n996 = pi28 & n995;
  assign n997 = ~pi29 & n996;
  assign n998 = pi30 & n997;
  assign n999 = pi05 & pi18;
  assign n1000 = pi19 & n999;
  assign n1001 = pi20 & n1000;
  assign n1002 = ~pi21 & n1001;
  assign n1003 = ~pi27 & n1002;
  assign n1004 = ~pi28 & n1003;
  assign n1005 = pi29 & n1004;
  assign n1006 = pi30 & n1005;
  assign n1007 = pi04 & pi18;
  assign n1008 = pi19 & n1007;
  assign n1009 = pi20 & n1008;
  assign n1010 = ~pi21 & n1009;
  assign n1011 = ~pi27 & n1010;
  assign n1012 = pi28 & n1011;
  assign n1013 = pi29 & n1012;
  assign n1014 = ~pi30 & n1013;
  assign n1015 = ~pi28 & n599;
  assign n1016 = pi29 & n1015;
  assign n1017 = ~pi30 & n1016;
  assign n1018 = pi28 & n634;
  assign n1019 = pi30 & n1018;
  assign n1020 = pi23 & n633;
  assign n1021 = ~pi29 & n1020;
  assign n1022 = pi30 & n1021;
  assign n1023 = pi29 & n1020;
  assign n1024 = ~pi30 & n1023;
  assign n1025 = pi31 & n1024;
  assign n1026 = ~pi31 & n1024;
  assign n1027 = pi32 & n1026;
  assign n1028 = ~pi32 & n1026;
  assign n1029 = ~pi33 & n1028;
  assign n1030 = pi34 & n1029;
  assign n1031 = ~pi34 & n1029;
  assign n1032 = pi35 & n1031;
  assign n1033 = ~pi35 & n1031;
  assign n1034 = ~pi36 & n1033;
  assign n1035 = pi37 & n1034;
  assign n1036 = ~n291 & ~n540;
  assign n1037 = ~n830 & n1036;
  assign n1038 = ~n973 & ~n981;
  assign n1039 = ~n537 & ~n965;
  assign n1040 = n1038 & n1039;
  assign n1041 = n1037 & n1040;
  assign n1042 = ~n277 & ~n533;
  assign n1043 = ~n530 & ~n962;
  assign n1044 = n1042 & n1043;
  assign n1045 = ~n525 & ~n954;
  assign n1046 = ~n514 & ~n519;
  assign n1047 = n1045 & n1046;
  assign n1048 = n1044 & n1047;
  assign n1049 = n1041 & n1048;
  assign n1050 = ~n510 & n679;
  assign n1051 = ~n488 & ~n948;
  assign n1052 = ~n156 & ~n482;
  assign n1053 = n1051 & n1052;
  assign n1054 = n1050 & n1053;
  assign n1055 = n676 & n892;
  assign n1056 = ~n473 & ~n476;
  assign n1057 = n674 & n1056;
  assign n1058 = n1055 & n1057;
  assign n1059 = n1054 & n1058;
  assign n1060 = n1049 & n1059;
  assign n1061 = ~n1030 & ~n1032;
  assign n1062 = ~n1035 & n1061;
  assign n1063 = ~n1025 & ~n1027;
  assign n1064 = ~n717 & ~n1022;
  assign n1065 = n1063 & n1064;
  assign n1066 = n1062 & n1065;
  assign n1067 = ~n401 & ~n601;
  assign n1068 = ~n1017 & ~n1019;
  assign n1069 = n1067 & n1068;
  assign n1070 = ~n598 & ~n1014;
  assign n1071 = ~n596 & ~n1006;
  assign n1072 = n1070 & n1071;
  assign n1073 = n1069 & n1072;
  assign n1074 = n1066 & n1073;
  assign n1075 = ~n588 & ~n876;
  assign n1076 = ~n591 & n1075;
  assign n1077 = n929 & n1076;
  assign n1078 = ~n563 & ~n866;
  assign n1079 = ~n555 & ~n998;
  assign n1080 = n1078 & n1079;
  assign n1081 = ~n544 & ~n547;
  assign n1082 = ~n552 & ~n989;
  assign n1083 = n1081 & n1082;
  assign n1084 = n1080 & n1083;
  assign n1085 = n1077 & n1084;
  assign n1086 = n1074 & n1085;
  assign po15 = ~n1060 | ~n1086;
  assign n1088 = pi22 & n534;
  assign n1089 = ~pi29 & n1088;
  assign po24 = pi30 & n1089;
  assign n1091 = pi29 & n963;
  assign n1092 = ~pi30 & n1091;
  assign n1093 = pi29 & n877;
  assign n1094 = ~pi30 & n1093;
  assign n1095 = ~n632 & ~n637;
  assign n1096 = ~n642 & n1095;
  assign n1097 = ~n625 & ~n628;
  assign n1098 = ~n631 & n1097;
  assign n1099 = n1096 & n1098;
  assign n1100 = ~n609 & ~n620;
  assign n1101 = ~n623 & n1100;
  assign n1102 = ~n401 & ~n1017;
  assign n1103 = n768 & n1102;
  assign n1104 = n1101 & n1103;
  assign n1105 = n1099 & n1104;
  assign n1106 = ~n1014 & n1071;
  assign n1107 = ~n879 & ~n1094;
  assign n1108 = n771 & n1107;
  assign n1109 = n1106 & n1108;
  assign n1110 = ~n584 & ~n874;
  assign n1111 = ~n876 & n1110;
  assign n1112 = ~n581 & ~n870;
  assign n1113 = n905 & n1112;
  assign n1114 = n1111 & n1113;
  assign n1115 = n1109 & n1114;
  assign n1116 = n1105 & n1115;
  assign n1117 = ~n457 & ~n510;
  assign n1118 = n892 & n1117;
  assign n1119 = ~n954 & n1046;
  assign n1120 = n1118 & n1119;
  assign n1121 = ~n291 & n1038;
  assign n1122 = ~po24 & ~n1092;
  assign n1123 = ~n277 & ~n962;
  assign n1124 = n1122 & n1123;
  assign n1125 = n1121 & n1124;
  assign n1126 = n1120 & n1125;
  assign n1127 = ~n851 & ~n989;
  assign n1128 = ~n555 & n1127;
  assign n1129 = ~n839 & ~n843;
  assign n1130 = n1081 & n1129;
  assign n1131 = n1128 & n1130;
  assign n1132 = ~n860 & ~n998;
  assign n1133 = ~n862 & n1132;
  assign n1134 = n908 & n1133;
  assign n1135 = n1131 & n1134;
  assign n1136 = n1126 & n1135;
  assign po16 = ~n1116 | ~n1136;
  assign n1138 = pi30 & n947;
  assign n1139 = pi22 & n761;
  assign n1140 = pi30 & n1139;
  assign n1141 = pi36 & n1033;
  assign n1142 = ~n1035 & ~n1141;
  assign n1143 = n1064 & n1142;
  assign n1144 = ~n765 & ~n921;
  assign n1145 = ~n918 & ~n1019;
  assign n1146 = n1144 & n1145;
  assign n1147 = n1143 & n1146;
  assign n1148 = ~n601 & ~n1017;
  assign n1149 = ~n598 & ~n1094;
  assign n1150 = n1148 & n1149;
  assign n1151 = ~n584 & ~n876;
  assign n1152 = ~n588 & n1151;
  assign n1153 = n771 & n1152;
  assign n1154 = n1150 & n1153;
  assign n1155 = n1147 & n1154;
  assign n1156 = ~po20 & ~n706;
  assign n1157 = n773 & n1156;
  assign n1158 = n880 & n1078;
  assign n1159 = n1157 & n1158;
  assign n1160 = ~n552 & ~n851;
  assign n1161 = n938 & n1160;
  assign n1162 = ~n830 & ~n839;
  assign n1163 = ~n540 & n1039;
  assign n1164 = n1162 & n1163;
  assign n1165 = n1161 & n1164;
  assign n1166 = n1159 & n1165;
  assign n1167 = n1155 & n1166;
  assign n1168 = ~n760 & ~n763;
  assign n1169 = ~n520 & ~n1140;
  assign n1170 = n1168 & n1169;
  assign n1171 = n783 & n1170;
  assign n1172 = ~n700 & ~n1138;
  assign n1173 = ~n494 & n1172;
  assign n1174 = n794 & n1173;
  assign n1175 = ~n515 & ~n703;
  assign n1176 = n792 & n1175;
  assign n1177 = n1174 & n1176;
  assign n1178 = n1171 & n1177;
  assign n1179 = ~n482 & ~n698;
  assign n1180 = n739 & n1179;
  assign n1181 = ~n473 & ~n693;
  assign n1182 = n800 & n1181;
  assign n1183 = n1180 & n1182;
  assign n1184 = ~n457 & ~n686;
  assign n1185 = ~n454 & n892;
  assign n1186 = n1184 & n1185;
  assign n1187 = n745 & n748;
  assign n1188 = n1186 & n1187;
  assign n1189 = n1183 & n1188;
  assign n1190 = n1178 & n1189;
  assign po17 = ~n1167 | ~n1190;
  assign n1192 = ~pi19 & n755;
  assign n1193 = ~pi20 & n1192;
  assign n1194 = ~pi21 & n1193;
  assign n1195 = pi25 & n1194;
  assign n1196 = pi30 & n1195;
  assign n1197 = ~n1017 & ~n1030;
  assign n1198 = ~n1032 & n1197;
  assign n1199 = n1142 & n1198;
  assign n1200 = ~n715 & ~n879;
  assign n1201 = ~n601 & n1200;
  assign n1202 = ~n870 & ~n874;
  assign n1203 = ~n588 & n1202;
  assign n1204 = n1201 & n1203;
  assign n1205 = n1199 & n1204;
  assign n1206 = ~n563 & ~n868;
  assign n1207 = ~n552 & ~n1196;
  assign n1208 = ~n862 & n1207;
  assign n1209 = n1206 & n1208;
  assign n1210 = n888 & n1209;
  assign n1211 = n1205 & n1210;
  assign n1212 = ~n540 & ~n830;
  assign n1213 = ~n826 & ~n965;
  assign n1214 = ~n537 & n1213;
  assign n1215 = n1212 & n1214;
  assign n1216 = ~n530 & ~n822;
  assign n1217 = ~n533 & n1216;
  assign n1218 = ~n525 & n679;
  assign n1219 = n1217 & n1218;
  assign n1220 = n1215 & n1219;
  assign n1221 = n675 & n1185;
  assign n1222 = ~n488 & ~n1138;
  assign n1223 = ~n156 & n680;
  assign n1224 = n1222 & n1223;
  assign n1225 = n1221 & n1224;
  assign n1226 = n1220 & n1225;
  assign po18 = ~n1211 | ~n1226;
  assign n1228 = pi33 & n1028;
  assign n1229 = ~n1027 & ~n1228;
  assign n1230 = ~n1032 & n1229;
  assign n1231 = ~n717 & n1068;
  assign n1232 = n1230 & n1231;
  assign n1233 = n721 & ~n879;
  assign n1234 = ~n601 & n719;
  assign n1235 = n1233 & n1234;
  assign n1236 = n1232 & n1235;
  assign n1237 = ~n876 & n1202;
  assign n1238 = ~n706 & n1206;
  assign n1239 = n1237 & n1238;
  assign n1240 = ~n860 & ~n864;
  assign n1241 = ~n866 & n1240;
  assign n1242 = n884 & n1160;
  assign n1243 = n1241 & n1242;
  assign n1244 = n1239 & n1243;
  assign n1245 = n1236 & n1244;
  assign n1246 = ~n502 & ~n514;
  assign n1247 = ~n519 & n1246;
  assign n1248 = ~n156 & ~n488;
  assign n1249 = ~n494 & n1248;
  assign n1250 = n1247 & n1249;
  assign n1251 = n674 & n676;
  assign n1252 = ~n482 & n1056;
  assign n1253 = n1251 & n1252;
  assign n1254 = n1250 & n1253;
  assign n1255 = ~n830 & ~n833;
  assign n1256 = ~n547 & n1255;
  assign n1257 = ~n537 & ~n826;
  assign n1258 = ~n540 & n1257;
  assign n1259 = n1256 & n1258;
  assign n1260 = ~n533 & ~po24;
  assign n1261 = ~n1092 & n1260;
  assign n1262 = ~n525 & ~n822;
  assign n1263 = ~n530 & n1262;
  assign n1264 = n1261 & n1263;
  assign n1265 = n1259 & n1264;
  assign n1266 = n1254 & n1265;
  assign po19 = ~n1245 | ~n1266;
  assign n1268 = ~pi10 & ~pi18;
  assign n1269 = ~pi19 & n1268;
  assign n1270 = pi20 & n1269;
  assign n1271 = pi21 & n1270;
  assign n1272 = pi25 & n1271;
  assign n1273 = pi19 & n1268;
  assign n1274 = pi21 & n1273;
  assign n1275 = pi25 & n1274;
  assign n1276 = ~pi28 & n1275;
  assign n1277 = ~pi29 & n1276;
  assign n1278 = pi30 & n1277;
  assign n1279 = pi05 & ~pi10;
  assign n1280 = pi18 & n1279;
  assign n1281 = ~pi19 & n1280;
  assign n1282 = pi20 & n1281;
  assign n1283 = pi21 & n1282;
  assign n1284 = pi25 & n1283;
  assign n1285 = ~pi28 & n1284;
  assign n1286 = ~pi29 & n1285;
  assign n1287 = pi30 & n1286;
  assign n1288 = ~pi10 & n201;
  assign n1289 = ~pi15 & n1288;
  assign n1290 = pi18 & n1289;
  assign n1291 = ~pi19 & n1290;
  assign n1292 = pi20 & n1291;
  assign n1293 = pi21 & n1292;
  assign n1294 = pi25 & n1293;
  assign n1295 = ~pi28 & n1294;
  assign n1296 = ~pi29 & n1295;
  assign n1297 = pi30 & n1296;
  assign n1298 = ~pi10 & pi18;
  assign n1299 = pi19 & n1298;
  assign n1300 = ~pi20 & n1299;
  assign n1301 = pi21 & n1300;
  assign n1302 = pi25 & n1301;
  assign n1303 = pi30 & n1302;
  assign n1304 = ~pi19 & n1298;
  assign n1305 = ~pi20 & n1304;
  assign n1306 = ~pi21 & n1305;
  assign n1307 = pi25 & n1306;
  assign n1308 = pi30 & n1307;
  assign n1309 = ~pi21 & n1300;
  assign n1310 = pi25 & n1309;
  assign n1311 = ~pi29 & n1310;
  assign n1312 = pi30 & n1311;
  assign n1313 = ~n1032 & ~n1141;
  assign n1314 = ~n1035 & n1313;
  assign n1315 = ~n1030 & ~n1228;
  assign n1316 = n1063 & n1315;
  assign n1317 = n1314 & n1316;
  assign n1318 = ~n717 & ~n765;
  assign n1319 = ~n1022 & n1318;
  assign n1320 = ~n642 & ~n921;
  assign n1321 = ~n637 & ~n1019;
  assign n1322 = n1320 & n1321;
  assign n1323 = n1319 & n1322;
  assign n1324 = n1317 & n1323;
  assign n1325 = ~n623 & ~n625;
  assign n1326 = ~n620 & ~n918;
  assign n1327 = n1325 & n1326;
  assign n1328 = n645 & n1327;
  assign n1329 = ~n609 & ~n1017;
  assign n1330 = n1067 & n1329;
  assign n1331 = ~n596 & ~n1014;
  assign n1332 = n768 & n1331;
  assign n1333 = n1330 & n1332;
  assign n1334 = n1328 & n1333;
  assign n1335 = n1324 & n1334;
  assign n1336 = ~n1006 & n1107;
  assign n1337 = n771 & n1075;
  assign n1338 = n1336 & n1337;
  assign n1339 = ~n874 & ~n1312;
  assign n1340 = ~n584 & n1339;
  assign n1341 = n1113 & n1340;
  assign n1342 = n1338 & n1341;
  assign n1343 = ~n864 & ~n866;
  assign n1344 = ~n862 & ~n1308;
  assign n1345 = n1343 & n1344;
  assign n1346 = n1238 & n1345;
  assign n1347 = ~n998 & ~n1196;
  assign n1348 = n938 & n1347;
  assign n1349 = ~n843 & ~n989;
  assign n1350 = n1160 & n1349;
  assign n1351 = n1348 & n1350;
  assign n1352 = n1346 & n1351;
  assign n1353 = n1342 & n1352;
  assign n1354 = n1335 & n1353;
  assign n1355 = ~n502 & ~n1297;
  assign n1356 = ~n701 & ~n1287;
  assign n1357 = n1355 & n1356;
  assign n1358 = n793 & n1357;
  assign n1359 = ~n494 & ~n1138;
  assign n1360 = ~n700 & ~n948;
  assign n1361 = n1359 & n1360;
  assign n1362 = n798 & n1248;
  assign n1363 = n1361 & n1362;
  assign n1364 = n1358 & n1363;
  assign n1365 = ~n693 & ~n1278;
  assign n1366 = ~n469 & ~n473;
  assign n1367 = n1365 & n1366;
  assign n1368 = n801 & n1367;
  assign n1369 = ~n454 & ~n814;
  assign n1370 = ~n686 & ~n1272;
  assign n1371 = n1369 & n1370;
  assign n1372 = n803 & n805;
  assign n1373 = n1371 & n1372;
  assign n1374 = n1368 & n1373;
  assign n1375 = n1364 & n1374;
  assign n1376 = ~n277 & n1043;
  assign n1377 = ~n822 & ~n954;
  assign n1378 = n782 & n1377;
  assign n1379 = n1376 & n1378;
  assign n1380 = ~n763 & ~n1303;
  assign n1381 = ~n760 & ~n1140;
  assign n1382 = n1380 & n1381;
  assign n1383 = n668 & n787;
  assign n1384 = n1382 & n1383;
  assign n1385 = n1379 & n1384;
  assign n1386 = ~n547 & ~n835;
  assign n1387 = ~n839 & n1386;
  assign n1388 = ~n291 & ~n830;
  assign n1389 = n886 & n1388;
  assign n1390 = n1387 & n1389;
  assign n1391 = ~n537 & ~n973;
  assign n1392 = ~n981 & n1391;
  assign n1393 = ~n826 & ~n1092;
  assign po43 = n965 | po24;
  assign n1395 = n1393 & ~po43;
  assign n1396 = n1392 & n1395;
  assign n1397 = n1390 & n1396;
  assign n1398 = n1385 & n1397;
  assign n1399 = n1375 & n1398;
  assign po22 = ~n1354 | ~n1399;
  assign n1401 = ~n457 & ~n514;
  assign po23 = n519 | ~n1401;
  assign n1403 = pi22 & n523;
  assign n1404 = pi30 & n1403;
  assign n1405 = pi26 & n534;
  assign n1406 = ~pi29 & n1405;
  assign n1407 = pi30 & n1406;
  assign n1408 = ~pi21 & n484;
  assign n1409 = pi22 & n1408;
  assign n1410 = pi30 & n1409;
  assign n1411 = ~n876 & ~n879;
  assign n1412 = ~n1022 & n1411;
  assign n1413 = ~n868 & ~n870;
  assign n1414 = n1339 & n1413;
  assign n1415 = n1412 & n1414;
  assign n1416 = ~n1196 & ~n1410;
  assign n1417 = n1129 & n1416;
  assign n1418 = n1345 & n1417;
  assign n1419 = n1415 & n1418;
  assign n1420 = ~n835 & n1255;
  assign n1421 = ~n826 & ~n1407;
  assign n1422 = ~po43 & n1421;
  assign n1423 = n1420 & n1422;
  assign n1424 = ~n820 & ~n1272;
  assign n1425 = ~n1278 & ~n1287;
  assign n1426 = n1424 & n1425;
  assign n1427 = ~n822 & ~n1404;
  assign n1428 = ~n1297 & ~n1303;
  assign n1429 = n1427 & n1428;
  assign n1430 = n1426 & n1429;
  assign n1431 = n1423 & n1430;
  assign po25 = ~n1419 | ~n1431;
  assign n1433 = ~n822 & ~n826;
  assign n1434 = ~n835 & ~n879;
  assign po26 = ~n1433 | ~n1434;
  assign n1436 = ~n954 & ~n962;
  assign n1437 = ~n277 & n1436;
  assign n1438 = n1121 & n1437;
  assign n1439 = ~n401 & ~n1014;
  assign n1440 = ~n989 & ~n998;
  assign n1441 = ~n1006 & n1440;
  assign n1442 = n1439 & n1441;
  assign po27 = ~n1438 | ~n1442;
  assign n1444 = pi21 & n984;
  assign n1445 = pi22 & n1444;
  assign n1446 = ~pi28 & n1445;
  assign n1447 = ~pi29 & n1446;
  assign n1448 = pi30 & n1447;
  assign n1449 = pi08 & pi16;
  assign n1450 = ~pi18 & n1449;
  assign n1451 = pi19 & n1450;
  assign n1452 = pi20 & n1451;
  assign n1453 = pi21 & n1452;
  assign n1454 = pi22 & n1453;
  assign n1455 = pi28 & n1454;
  assign n1456 = ~pi29 & n1455;
  assign n1457 = ~pi30 & n1456;
  assign n1458 = pi07 & ~pi16;
  assign n1459 = ~pi18 & n1458;
  assign n1460 = pi19 & n1459;
  assign n1461 = pi20 & n1460;
  assign n1462 = pi21 & n1461;
  assign n1463 = pi22 & n1462;
  assign n1464 = pi28 & n1463;
  assign n1465 = ~pi29 & n1464;
  assign n1466 = ~pi30 & n1465;
  assign n1467 = ~pi19 & n999;
  assign n1468 = pi20 & n1467;
  assign n1469 = pi21 & n1468;
  assign n1470 = ~pi25 & n1469;
  assign n1471 = ~pi28 & n1470;
  assign n1472 = ~pi29 & n1471;
  assign n1473 = pi30 & n1472;
  assign n1474 = pi05 & pi10;
  assign n1475 = pi18 & n1474;
  assign n1476 = ~pi19 & n1475;
  assign n1477 = pi20 & n1476;
  assign n1478 = pi21 & n1477;
  assign n1479 = pi25 & n1478;
  assign n1480 = ~pi28 & n1479;
  assign n1481 = ~pi29 & n1480;
  assign n1482 = pi30 & n1481;
  assign n1483 = pi18 & n1449;
  assign n1484 = ~pi19 & n1483;
  assign n1485 = pi20 & n1484;
  assign n1486 = pi21 & n1485;
  assign n1487 = pi28 & n1486;
  assign n1488 = pi18 & n1458;
  assign n1489 = ~pi19 & n1488;
  assign n1490 = pi20 & n1489;
  assign n1491 = pi21 & n1490;
  assign n1492 = pi28 & n1491;
  assign n1493 = ~pi37 & n1034;
  assign n1494 = ~n1035 & ~n1493;
  assign n1495 = n1061 & ~n1141;
  assign n1496 = n1494 & n1495;
  assign n1497 = ~n765 & ~n1019;
  assign n1498 = ~n1025 & n1497;
  assign n1499 = n1229 & n1498;
  assign n1500 = n1496 & n1499;
  assign n1501 = ~n764 & ~n1404;
  assign n1502 = ~po24 & n1501;
  assign n1503 = n1168 & ~n1303;
  assign n1504 = n1502 & n1503;
  assign n1505 = ~n1092 & ~n1407;
  assign n1506 = ~n1410 & n1505;
  assign n1507 = ~n1196 & ~n1308;
  assign n1508 = n1506 & n1507;
  assign n1509 = n1504 & n1508;
  assign n1510 = n1500 & n1509;
  assign n1511 = ~n687 & ~n1278;
  assign n1512 = ~n693 & n1511;
  assign n1513 = ~n458 & n1370;
  assign n1514 = n1512 & n1513;
  assign n1515 = ~n1457 & ~n1466;
  assign n1516 = ~n697 & ~n698;
  assign n1517 = ~n1448 & n1516;
  assign n1518 = n1515 & n1517;
  assign n1519 = n1514 & n1518;
  assign n1520 = ~n1487 & ~n1492;
  assign n1521 = ~n703 & n1520;
  assign n1522 = n1169 & n1521;
  assign n1523 = ~n1287 & ~n1297;
  assign n1524 = ~n1138 & ~n1473;
  assign n1525 = ~n1482 & n1524;
  assign n1526 = n1523 & n1525;
  assign n1527 = n1522 & n1526;
  assign n1528 = n1519 & n1527;
  assign po28 = ~n1510 | ~n1528;
  assign n1530 = ~n291 & ~n299;
  assign n1531 = ~n314 & n1530;
  assign n1532 = ~n362 & ~n384;
  assign n1533 = ~n401 & n1532;
  assign n1534 = n1531 & n1533;
  assign n1535 = ~n249 & ~n259;
  assign n1536 = ~n161 & n1535;
  assign n1537 = ~n268 & ~n277;
  assign n1538 = ~n282 & n1537;
  assign n1539 = n1536 & n1538;
  assign n1540 = n1534 & n1539;
  assign n1541 = ~n192 & ~n200;
  assign n1542 = ~n144 & n1541;
  assign n1543 = ~n184 & n422;
  assign n1544 = n1542 & n1543;
  assign n1545 = ~n149 & ~po41;
  assign n1546 = ~n156 & n1545;
  assign n1547 = ~n239 & n425;
  assign n1548 = n1546 & n1547;
  assign n1549 = n1544 & n1548;
  assign po29 = ~n1540 | ~n1549;
  assign n1551 = ~n351 & ~n358;
  assign n1552 = ~n393 & n1551;
  assign n1553 = ~n305 & ~n323;
  assign n1554 = ~n344 & n1553;
  assign po30 = ~n1552 | ~n1554;
  assign n1556 = ~n393 & n404;
  assign n1557 = ~n305 & ~n331;
  assign n1558 = ~n339 & n1557;
  assign po31 = ~n1556 | ~n1558;
  assign n1560 = ~pi12 & ~pi13;
  assign n1561 = ~pi14 & n1560;
  assign n1562 = pi21 & n1561;
  assign n1563 = ~pi27 & n1562;
  assign n1564 = ~pi28 & n1563;
  assign n1565 = ~pi29 & n1564;
  assign po32 = ~pi30 & n1565;
  assign n1567 = ~n1006 & ~n1014;
  assign n1568 = ~n598 & n1567;
  assign po33 = ~n1067 | ~n1568;
  assign n1570 = ~pi29 & n531;
  assign n1571 = ~pi30 & n1570;
  assign n1572 = ~pi29 & n538;
  assign n1573 = ~pi30 & n1572;
  assign n1574 = ~pi29 & n553;
  assign n1575 = ~pi30 & n1574;
  assign n1576 = pi30 & n595;
  assign n1577 = pi31 & n617;
  assign n1578 = ~pi39 & n619;
  assign n1579 = ~n642 & ~n717;
  assign n1580 = n923 & n1579;
  assign n1581 = ~n628 & n1325;
  assign n1582 = ~n1577 & ~n1578;
  assign n1583 = ~n620 & n1582;
  assign n1584 = n1581 & n1583;
  assign n1585 = n1580 & n1584;
  assign n1586 = ~n393 & ~n1576;
  assign n1587 = ~n918 & n1586;
  assign n1588 = ~n376 & ~n384;
  assign n1589 = ~n596 & n1588;
  assign n1590 = n1587 & n1589;
  assign n1591 = ~n331 & ~n706;
  assign n1592 = ~n339 & n1591;
  assign n1593 = ~n369 & n721;
  assign n1594 = n1592 & n1593;
  assign n1595 = n1590 & n1594;
  assign n1596 = n1585 & n1595;
  assign n1597 = ~n149 & ~n476;
  assign n1598 = ~n699 & n1597;
  assign n1599 = ~n104 & ~n111;
  assign n1600 = ~n115 & n1599;
  assign n1601 = n1598 & n1600;
  assign n1602 = ~n701 & n1360;
  assign n1603 = ~n515 & ~n702;
  assign n1604 = ~n530 & n1603;
  assign n1605 = n1602 & n1604;
  assign n1606 = n1601 & n1605;
  assign n1607 = ~n277 & ~n1571;
  assign n1608 = ~n537 & n1607;
  assign n1609 = ~n291 & ~n1573;
  assign n1610 = ~n552 & n1609;
  assign n1611 = n1608 & n1610;
  assign n1612 = ~n563 & ~n860;
  assign n1613 = ~n851 & ~n1575;
  assign n1614 = ~n305 & n1613;
  assign n1615 = n1612 & n1614;
  assign n1616 = n1611 & n1615;
  assign n1617 = n1606 & n1616;
  assign po34 = ~n1596 | ~n1617;
  assign n1619 = ~pi19 & n853;
  assign n1620 = ~pi20 & n1619;
  assign n1621 = ~pi21 & n1620;
  assign n1622 = pi28 & n1621;
  assign n1623 = ~pi29 & n1622;
  assign n1624 = pi30 & n1623;
  assign n1625 = pi03 & ~pi06;
  assign n1626 = ~pi18 & n1625;
  assign n1627 = ~pi19 & n1626;
  assign n1628 = pi20 & n1627;
  assign n1629 = ~pi21 & n1628;
  assign n1630 = pi28 & n1629;
  assign n1631 = ~pi29 & n1630;
  assign n1632 = pi30 & n1631;
  assign n1633 = ~pi06 & n852;
  assign n1634 = ~pi18 & n1633;
  assign n1635 = ~pi19 & n1634;
  assign n1636 = pi20 & n1635;
  assign n1637 = ~pi21 & n1636;
  assign n1638 = pi28 & n1637;
  assign n1639 = ~pi29 & n1638;
  assign n1640 = pi30 & n1639;
  assign n1641 = ~n632 & ~n1022;
  assign n1642 = ~n601 & ~n609;
  assign n1643 = n1641 & n1642;
  assign n1644 = ~n393 & ~n715;
  assign n1645 = ~n1006 & ~n1576;
  assign n1646 = ~n1014 & n1645;
  assign n1647 = n1644 & n1646;
  assign n1648 = n1643 & n1647;
  assign n1649 = n404 & n1107;
  assign n1650 = ~n362 & ~n876;
  assign n1651 = ~n351 & ~n874;
  assign n1652 = ~n358 & n1651;
  assign n1653 = n1650 & n1652;
  assign n1654 = n1649 & n1653;
  assign n1655 = n1648 & n1654;
  assign n1656 = ~n344 & ~n870;
  assign n1657 = n409 & n1656;
  assign n1658 = ~n860 & ~n866;
  assign n1659 = ~n868 & n1658;
  assign n1660 = n411 & n1659;
  assign n1661 = n1657 & n1660;
  assign n1662 = ~n833 & ~n835;
  assign n1663 = ~n291 & ~n1640;
  assign n1664 = ~n830 & n1663;
  assign n1665 = n1662 & n1664;
  assign n1666 = ~n299 & ~n851;
  assign n1667 = ~n305 & ~n555;
  assign n1668 = n1666 & n1667;
  assign n1669 = n1665 & n1668;
  assign n1670 = n1661 & n1669;
  assign n1671 = n1655 & n1670;
  assign n1672 = ~n277 & ~n1624;
  assign n1673 = ~n268 & n1262;
  assign n1674 = n1672 & n1673;
  assign n1675 = ~n282 & ~n1632;
  assign n1676 = n1213 & n1675;
  assign n1677 = n1674 & n1676;
  assign n1678 = ~n161 & ~n519;
  assign n1679 = ~n259 & ~n514;
  assign n1680 = n1678 & n1679;
  assign n1681 = ~n249 & ~n510;
  assign n1682 = ~n229 & ~n502;
  assign n1683 = ~n239 & n1682;
  assign n1684 = n1681 & n1683;
  assign n1685 = n1680 & n1684;
  assign n1686 = n1677 & n1685;
  assign n1687 = ~n200 & ~n457;
  assign n1688 = ~n144 & n1687;
  assign n1689 = n674 & n1688;
  assign n1690 = ~n167 & ~n454;
  assign n1691 = ~n176 & n1690;
  assign n1692 = n423 & n1691;
  assign n1693 = n1689 & n1692;
  assign n1694 = ~n218 & ~n494;
  assign n1695 = n1248 & n1694;
  assign n1696 = ~po41 & ~n482;
  assign n1697 = ~n149 & ~n473;
  assign n1698 = ~n476 & n1697;
  assign n1699 = n1696 & n1698;
  assign n1700 = n1695 & n1699;
  assign n1701 = n1693 & n1700;
  assign n1702 = n1686 & n1701;
  assign po35 = ~n1671 | ~n1702;
  assign n1704 = ~pi14 & ~pi18;
  assign n1705 = ~pi19 & n1704;
  assign n1706 = pi20 & n1705;
  assign n1707 = ~pi21 & n1706;
  assign n1708 = ~pi23 & n1707;
  assign n1709 = ~pi27 & n1708;
  assign n1710 = ~pi28 & n1709;
  assign n1711 = ~pi29 & n1710;
  assign n1712 = ~pi30 & n1711;
  assign n1713 = ~pi14 & pi18;
  assign n1714 = ~pi19 & n1713;
  assign n1715 = ~pi20 & n1714;
  assign n1716 = ~pi21 & n1715;
  assign n1717 = ~pi27 & n1716;
  assign n1718 = ~pi28 & n1717;
  assign n1719 = ~pi29 & n1718;
  assign n1720 = ~pi30 & n1719;
  assign n1721 = ~pi21 & n815;
  assign n1722 = ~pi27 & n1721;
  assign n1723 = ~pi28 & n1722;
  assign n1724 = ~pi29 & n1723;
  assign n1725 = ~pi30 & n1724;
  assign n1726 = ~pi05 & pi15;
  assign n1727 = ~pi18 & n1726;
  assign n1728 = pi19 & n1727;
  assign n1729 = pi20 & n1728;
  assign n1730 = pi21 & n1729;
  assign n1731 = pi22 & n1730;
  assign n1732 = ~pi28 & n1731;
  assign n1733 = ~pi29 & n1732;
  assign n1734 = pi30 & n1733;
  assign n1735 = ~pi08 & pi16;
  assign n1736 = ~pi18 & n1735;
  assign n1737 = pi19 & n1736;
  assign n1738 = pi20 & n1737;
  assign n1739 = pi21 & n1738;
  assign n1740 = pi22 & n1739;
  assign n1741 = pi28 & n1740;
  assign n1742 = ~pi29 & n1741;
  assign n1743 = ~pi30 & n1742;
  assign n1744 = ~pi07 & ~pi16;
  assign n1745 = ~pi18 & n1744;
  assign n1746 = pi19 & n1745;
  assign n1747 = pi20 & n1746;
  assign n1748 = pi21 & n1747;
  assign n1749 = pi22 & n1748;
  assign n1750 = pi28 & n1749;
  assign n1751 = ~pi29 & n1750;
  assign n1752 = ~pi30 & n1751;
  assign n1753 = pi18 & n1726;
  assign n1754 = ~pi19 & n1753;
  assign n1755 = pi20 & n1754;
  assign n1756 = pi21 & n1755;
  assign n1757 = ~pi28 & n1756;
  assign n1758 = ~pi29 & n1757;
  assign n1759 = pi30 & n1758;
  assign n1760 = pi18 & n1744;
  assign n1761 = ~pi19 & n1760;
  assign n1762 = pi20 & n1761;
  assign n1763 = pi21 & n1762;
  assign n1764 = pi28 & n1763;
  assign n1765 = pi18 & n1735;
  assign n1766 = ~pi19 & n1765;
  assign n1767 = pi20 & n1766;
  assign n1768 = pi21 & n1767;
  assign n1769 = pi28 & n1768;
  assign n1770 = ~n632 & ~n918;
  assign n1771 = ~n921 & n1770;
  assign n1772 = ~n401 & n1644;
  assign n1773 = n1771 & n1772;
  assign n1774 = ~n362 & n1551;
  assign n1775 = ~n708 & ~n1094;
  assign n1776 = ~n596 & n1775;
  assign n1777 = n1774 & n1776;
  assign n1778 = n1773 & n1777;
  assign n1779 = ~n323 & ~n706;
  assign n1780 = ~n344 & n1779;
  assign n1781 = ~n305 & ~n1575;
  assign n1782 = ~n314 & n1781;
  assign n1783 = n1780 & n1782;
  assign n1784 = ~n282 & ~n1573;
  assign n1785 = ~n299 & n1784;
  assign n1786 = ~n268 & ~n1571;
  assign n1787 = ~n519 & ~n525;
  assign n1788 = n1786 & n1787;
  assign n1789 = n1785 & n1788;
  assign n1790 = n1783 & n1789;
  assign n1791 = n1778 & n1790;
  assign n1792 = ~n476 & ~n1734;
  assign n1793 = ~n482 & n1792;
  assign n1794 = n1600 & n1793;
  assign n1795 = ~n1712 & ~n1720;
  assign n1796 = ~po32 & ~n1725;
  assign n1797 = n1795 & n1796;
  assign n1798 = ~n461 & n676;
  assign n1799 = n1797 & n1798;
  assign n1800 = n1794 & n1799;
  assign n1801 = ~n514 & n792;
  assign n1802 = ~n1764 & ~n1769;
  assign n1803 = ~n502 & n1802;
  assign n1804 = n1801 & n1803;
  assign n1805 = ~n494 & ~n948;
  assign n1806 = ~n1759 & n1805;
  assign n1807 = ~n1743 & ~n1752;
  assign n1808 = ~n488 & n1807;
  assign n1809 = n1806 & n1808;
  assign n1810 = n1804 & n1809;
  assign n1811 = n1800 & n1810;
  assign po36 = ~n1791 | ~n1811;
  assign n1813 = n1063 & ~n1228;
  assign n1814 = n1319 & n1813;
  assign n1815 = n1496 & n1814;
  assign n1816 = ~n1019 & n1095;
  assign n1817 = n1320 & n1816;
  assign n1818 = ~n620 & ~n1578;
  assign n1819 = ~n623 & n1818;
  assign n1820 = n1098 & n1819;
  assign n1821 = n1817 & n1820;
  assign n1822 = n1815 & n1821;
  assign n1823 = ~n918 & ~n1577;
  assign n1824 = ~n609 & n1148;
  assign n1825 = n1823 & n1824;
  assign n1826 = ~n401 & n768;
  assign n1827 = ~n1014 & ~n1576;
  assign n1828 = ~n393 & n1827;
  assign n1829 = n1826 & n1828;
  assign n1830 = n1825 & n1829;
  assign n1831 = ~n384 & ~n1006;
  assign n1832 = ~n596 & n1831;
  assign n1833 = n912 & ~n1094;
  assign n1834 = n1832 & n1833;
  assign n1835 = ~n369 & ~n708;
  assign n1836 = ~n376 & n1835;
  assign n1837 = ~n588 & n1650;
  assign n1838 = n1836 & n1837;
  assign n1839 = n1834 & n1838;
  assign n1840 = n1830 & n1839;
  assign n1841 = n1822 & n1840;
  assign n1842 = ~n358 & ~n584;
  assign n1843 = ~n351 & n1339;
  assign n1844 = n1842 & n1843;
  assign n1845 = ~n581 & n1656;
  assign n1846 = n409 & ~po21;
  assign n1847 = n1845 & n1846;
  assign n1848 = n1844 & n1847;
  assign n1849 = ~po20 & n1779;
  assign n1850 = ~n314 & ~n868;
  assign n1851 = ~n563 & n1850;
  assign n1852 = n1849 & n1851;
  assign n1853 = ~n1308 & n1416;
  assign n1854 = ~n866 & n880;
  assign n1855 = n1853 & n1854;
  assign n1856 = n1852 & n1855;
  assign n1857 = n1848 & n1856;
  assign n1858 = ~n305 & ~n851;
  assign n1859 = ~n555 & n1858;
  assign n1860 = n1132 & n1859;
  assign n1861 = ~n299 & ~n552;
  assign n1862 = ~n1575 & n1861;
  assign n1863 = ~n989 & n1129;
  assign n1864 = n1862 & n1863;
  assign n1865 = n1860 & n1864;
  assign n1866 = ~n547 & ~n833;
  assign n1867 = ~n835 & n1866;
  assign n1868 = ~n544 & n1212;
  assign n1869 = n1867 & n1868;
  assign n1870 = ~n1573 & ~n1632;
  assign n1871 = ~n1640 & n1870;
  assign n1872 = n1121 & n1871;
  assign n1873 = n1869 & n1872;
  assign n1874 = n1865 & n1873;
  assign n1875 = n1857 & n1874;
  assign n1876 = n1841 & n1875;
  assign n1877 = ~n282 & ~n537;
  assign n1878 = ~n826 & n1505;
  assign n1879 = n1877 & n1878;
  assign n1880 = ~n965 & n1260;
  assign n1881 = ~n1571 & ~n1624;
  assign n1882 = ~n277 & n1881;
  assign n1883 = n1880 & n1882;
  assign n1884 = n1879 & n1883;
  assign n1885 = ~n268 & ~n962;
  assign n1886 = ~n530 & n1885;
  assign n1887 = ~n764 & ~n822;
  assign n1888 = ~n954 & n1887;
  assign n1889 = n1886 & n1888;
  assign n1890 = ~n161 & ~n1404;
  assign n1891 = ~n525 & n1890;
  assign n1892 = n1503 & n1891;
  assign n1893 = n1889 & n1892;
  assign n1894 = n1884 & n1893;
  assign n1895 = ~n259 & ~n515;
  assign n1896 = ~n519 & n1895;
  assign n1897 = n1169 & n1896;
  assign n1898 = ~n239 & ~n702;
  assign n1899 = ~n510 & n1898;
  assign n1900 = ~n249 & ~n703;
  assign n1901 = ~n514 & n1900;
  assign n1902 = n1899 & n1901;
  assign n1903 = n1897 & n1902;
  assign n1904 = ~n1297 & ~n1487;
  assign n1905 = ~n1492 & n1904;
  assign n1906 = ~n229 & ~n1769;
  assign n1907 = ~n502 & n1906;
  assign n1908 = n1905 & n1907;
  assign n1909 = ~n1473 & ~n1482;
  assign n1910 = ~n1287 & n1909;
  assign n1911 = ~n701 & ~n1759;
  assign n1912 = ~n1764 & n1911;
  assign n1913 = n1910 & n1912;
  assign n1914 = n1908 & n1913;
  assign n1915 = n1903 & n1914;
  assign n1916 = n1894 & n1915;
  assign n1917 = ~n1138 & n1360;
  assign n1918 = n1694 & n1917;
  assign n1919 = ~n1457 & ~n1743;
  assign n1920 = ~n1752 & n1919;
  assign n1921 = ~n156 & ~n1466;
  assign n1922 = ~n488 & n1921;
  assign n1923 = n1920 & n1922;
  assign n1924 = n1918 & n1923;
  assign n1925 = ~n149 & ~n697;
  assign n1926 = ~n476 & n1925;
  assign n1927 = ~n473 & ~n1278;
  assign n1928 = ~n693 & n1927;
  assign n1929 = n1926 & n1928;
  assign n1930 = ~n698 & ~n1448;
  assign n1931 = ~n1734 & n1930;
  assign n1932 = ~n699 & n1696;
  assign n1933 = n1931 & n1932;
  assign n1934 = n1929 & n1933;
  assign n1935 = n1924 & n1934;
  assign n1936 = ~n115 & ~n469;
  assign n1937 = ~n104 & ~n687;
  assign n1938 = ~n111 & n1937;
  assign n1939 = n1936 & n1938;
  assign n1940 = ~n144 & ~n458;
  assign n1941 = ~n461 & n1940;
  assign n1942 = ~n457 & n1541;
  assign n1943 = n1941 & n1942;
  assign n1944 = n1939 & n1943;
  assign n1945 = ~n686 & n1690;
  assign n1946 = ~n176 & ~n1272;
  assign n1947 = ~n184 & n1946;
  assign n1948 = n1945 & n1947;
  assign n1949 = ~n1720 & ~n1725;
  assign n1950 = ~po32 & n1949;
  assign n1951 = pi19 & pi20;
  assign n1952 = pi18 & n1951;
  assign n1953 = pi26 & pi30;
  assign n1954 = pi21 & n1953;
  assign n1955 = n1952 & n1954;
  assign n1956 = ~n814 & ~n1955;
  assign n1957 = ~n1712 & n1956;
  assign n1958 = n1950 & n1957;
  assign n1959 = n1948 & n1958;
  assign n1960 = n1944 & n1959;
  assign n1961 = n1935 & n1960;
  assign n1962 = n1916 & n1961;
  assign po37 = ~n1876 | ~n1962;
  assign n1964 = ~pi19 & pi20;
  assign n1965 = ~pi18 & n1964;
  assign n1966 = ~pi29 & pi30;
  assign n1967 = pi21 & n1966;
  assign n1968 = n1965 & n1967;
  assign n1969 = pi19 & ~pi20;
  assign n1970 = pi18 & n1969;
  assign n1971 = pi29 & ~pi30;
  assign n1972 = ~pi21 & n1971;
  assign n1973 = n1970 & n1972;
  assign n1974 = ~n1968 & ~n1973;
  assign n1975 = ~pi22 & ~pi25;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~pi05 & ~pi28;
  assign n1978 = ~pi28 & ~n1977;
  assign n1979 = pi22 & ~n1978;
  assign n1980 = pi19 & n1979;
  assign n1981 = pi23 & ~pi28;
  assign n1982 = ~pi19 & n1981;
  assign n1983 = ~n1980 & ~n1982;
  assign n1984 = ~pi18 & ~n1983;
  assign n1985 = pi26 & ~pi28;
  assign n1986 = ~pi19 & n1985;
  assign n1987 = ~pi04 & ~pi27;
  assign n1988 = pi19 & pi28;
  assign n1989 = n1987 & n1988;
  assign n1990 = ~n1986 & ~n1989;
  assign n1991 = pi18 & ~n1990;
  assign n1992 = ~n1984 & ~n1991;
  assign n1993 = ~pi30 & ~n1992;
  assign n1994 = pi19 & ~pi28;
  assign n1995 = pi18 & n1994;
  assign n1996 = ~pi05 & ~pi27;
  assign n1997 = pi30 & n1996;
  assign n1998 = n1995 & n1997;
  assign n1999 = ~n1993 & ~n1998;
  assign n2000 = pi29 & ~n1999;
  assign n2001 = ~pi19 & pi28;
  assign n2002 = pi11 & pi26;
  assign n2003 = pi30 & n2002;
  assign n2004 = n2001 & n2003;
  assign n2005 = pi03 & pi27;
  assign n2006 = pi19 & n2005;
  assign n2007 = ~n2004 & ~n2006;
  assign n2008 = pi18 & ~n2007;
  assign n2009 = ~pi18 & n2001;
  assign n2010 = pi30 & n990;
  assign n2011 = n2009 & n2010;
  assign n2012 = ~n2008 & ~n2011;
  assign n2013 = ~pi29 & ~n2012;
  assign n2014 = ~n2000 & ~n2013;
  assign n2015 = pi20 & ~n2014;
  assign n2016 = pi28 & n1966;
  assign n2017 = ~pi28 & n1971;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = pi26 & ~n2018;
  assign n2020 = pi19 & n2019;
  assign n2021 = pi18 & n2020;
  assign n2022 = ~pi28 & pi29;
  assign n2023 = ~pi05 & ~pi30;
  assign n2024 = n2022 & n2023;
  assign n2025 = pi28 & ~pi29;
  assign n2026 = ~pi02 & pi30;
  assign n2027 = n2025 & n2026;
  assign n2028 = ~n2024 & ~n2027;
  assign n2029 = ~pi03 & ~n2028;
  assign n2030 = ~pi19 & n2029;
  assign n2031 = ~pi18 & n2030;
  assign n2032 = ~n2021 & ~n2031;
  assign n2033 = ~pi20 & ~n2032;
  assign n2034 = ~n2015 & ~n2033;
  assign n2035 = ~pi21 & ~n2034;
  assign n2036 = pi20 & pi22;
  assign n2037 = ~pi05 & ~pi15;
  assign n2038 = ~pi28 & n2037;
  assign n2039 = n2036 & n2038;
  assign n2040 = ~pi28 & ~n2039;
  assign n2041 = pi19 & ~n2040;
  assign n2042 = pi20 & pi26;
  assign n2043 = ~pi19 & n2042;
  assign n2044 = ~n2041 & ~n2043;
  assign n2045 = ~pi18 & ~n2044;
  assign n2046 = pi18 & n1964;
  assign n2047 = n2038 & n2046;
  assign n2048 = ~n2045 & ~n2047;
  assign n2049 = pi30 & ~n2048;
  assign n2050 = ~pi29 & n2049;
  assign n2051 = pi21 & n2050;
  assign n2052 = ~n2035 & ~n2051;
  assign n2053 = ~n1976 & n2052;
  assign n2054 = ~pi00 & ~n2053;
  assign n2055 = ~pi22 & ~pi23;
  assign n2056 = pi21 & ~pi28;
  assign n2057 = n1966 & n2056;
  assign n2058 = ~n1972 & ~n2057;
  assign n2059 = ~n2055 & ~n2058;
  assign n2060 = ~pi20 & n2059;
  assign n2061 = pi19 & n2060;
  assign n2062 = ~pi18 & n2061;
  assign n2063 = ~pi01 & n2062;
  assign n2064 = ~n122 & ~n128;
  assign n2065 = ~n98 & n2064;
  assign n2066 = ~n2063 & n2065;
  assign po38 = n2054 | ~n2066;
  assign n2068 = ~n591 & ~n1014;
  assign n2069 = ~n601 & n2068;
  assign n2070 = n929 & n2069;
  assign n2071 = ~n547 & ~n989;
  assign n2072 = ~n998 & n2071;
  assign n2073 = ~n533 & ~n537;
  assign n2074 = n664 & n2073;
  assign n2075 = n2072 & n2074;
  assign n2076 = n2070 & n2075;
  assign n2077 = ~n525 & n1046;
  assign n2078 = ~n502 & ~n510;
  assign n2079 = ~n488 & ~n494;
  assign n2080 = n2078 & n2079;
  assign n2081 = n2077 & n2080;
  assign n2082 = n1253 & n2081;
  assign po39 = ~n2076 | ~n2082;
  assign n2084 = ~n1448 & ~n1473;
  assign n2085 = ~n954 & ~n1482;
  assign n2086 = n2084 & n2085;
  assign n2087 = ~n962 & ~n989;
  assign n2088 = ~n1006 & n2087;
  assign po40 = ~n2086 | ~n2088;
  assign po02 = 1'b0;
  assign po42 = 1'b0;
  assign po44 = po24;
endmodule



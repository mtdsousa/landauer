module top (
            a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, 
            sin_0, sin_1, sin_2, sin_3, sin_4, sin_5, sin_6, sin_7, sin_8, sin_9, sin_10, sin_11, sin_12, sin_13, sin_14, sin_15, sin_16, sin_17, sin_18, sin_19, sin_20, sin_21, sin_22, sin_23, sin_24);
input a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23;
output sin_0, sin_1, sin_2, sin_3, sin_4, sin_5, sin_6, sin_7, sin_8, sin_9, sin_10, sin_11, sin_12, sin_13, sin_14, sin_15, sin_16, sin_17, sin_18, sin_19, sin_20, sin_21, sin_22, sin_23, sin_24;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894;
assign w0 = ~a_0 & ~a_1;
assign w1 = ~a_2 & ~a_3;
assign w2 = w0 & w1;
assign w3 = ~a_4 & ~a_5;
assign w4 = ~a_6 & w3;
assign w5 = w2 & w4;
assign w6 = ~a_7 & ~a_8;
assign w7 = ~a_9 & w6;
assign w8 = ~a_10 & ~a_11;
assign w9 = ~a_12 & w8;
assign w10 = w7 & w9;
assign w11 = w5 & w10;
assign w12 = ~a_13 & ~a_14;
assign w13 = ~a_15 & w12;
assign w14 = w11 & w13;
assign w15 = ~a_16 & ~a_17;
assign w16 = ~a_22 & w15;
assign w17 = (w16 & ~w11) | (w16 & w5433) | (~w11 & w5433);
assign w18 = a_16 & ~a_17;
assign w19 = ~a_22 & w18;
assign w20 = w13 & w19;
assign w21 = a_16 & a_17;
assign w22 = a_22 & w21;
assign w23 = (~w22 & ~w11) | (~w22 & w5434) | (~w11 & w5434);
assign w24 = ~w17 & w23;
assign w25 = ~a_22 & w12;
assign w26 = ~a_15 & ~a_22;
assign w27 = a_15 & a_22;
assign w28 = ~w26 & ~w27;
assign w29 = (w28 & ~w11) | (w28 & w5435) | (~w11 & w5435);
assign w30 = ~w14 & ~w29;
assign w31 = ~w24 & w30;
assign w32 = w13 & w15;
assign w33 = ~a_18 & ~a_19;
assign w34 = ~a_22 & w33;
assign w35 = (w34 & ~w11) | (w34 & w5436) | (~w11 & w5436);
assign w36 = w13 & w16;
assign w37 = a_18 & ~a_19;
assign w38 = w36 & w37;
assign w39 = w11 & w38;
assign w40 = a_18 & a_19;
assign w41 = a_22 & w40;
assign w42 = ~w39 & ~w41;
assign w43 = ~w35 & w42;
assign w44 = w15 & w33;
assign w45 = w13 & w44;
assign w46 = ~a_20 & ~a_21;
assign w47 = ~a_22 & w46;
assign w48 = (w47 & ~w11) | (w47 & w5437) | (~w11 & w5437);
assign w49 = a_20 & ~a_21;
assign w50 = ~a_22 & w49;
assign w51 = w45 & w50;
assign w52 = w11 & w51;
assign w53 = a_20 & a_21;
assign w54 = a_22 & w53;
assign w55 = ~w52 & ~w54;
assign w56 = ~w48 & w55;
assign w57 = ~w43 & ~w56;
assign w58 = w31 & w57;
assign w59 = ~a_22 & ~w37;
assign w60 = (w59 & ~w11) | (w59 & w5438) | (~w11 & w5438);
assign w61 = ~a_18 & a_19;
assign w62 = w13 & w5439;
assign w63 = a_22 & ~w61;
assign w64 = (~w63 & ~w11) | (~w63 & w5440) | (~w11 & w5440);
assign w65 = ~w60 & w64;
assign w66 = ~a_22 & w21;
assign w67 = (w66 & ~w11) | (w66 & w5441) | (~w11 & w5441);
assign w68 = a_22 & w15;
assign w69 = (~w68 & ~w11) | (~w68 & w5442) | (~w11 & w5442);
assign w70 = ~w67 & w69;
assign w71 = w65 & ~w70;
assign w72 = ~a_22 & w53;
assign w73 = (w72 & ~w11) | (w72 & w5443) | (~w11 & w5443);
assign w74 = a_22 & w46;
assign w75 = w45 & w46;
assign w76 = w11 & w75;
assign w77 = ~w74 & ~w76;
assign w78 = ~w73 & w77;
assign w79 = ~w30 & ~w78;
assign w80 = w71 & w79;
assign w81 = (w19 & ~w11) | (w19 & w5444) | (~w11 & w5444);
assign w82 = ~a_16 & a_17;
assign w83 = a_22 & w82;
assign w84 = w13 & w82;
assign w85 = (~w83 & ~w11) | (~w83 & w5445) | (~w11 & w5445);
assign w86 = ~w81 & w85;
assign w87 = w30 & ~w86;
assign w88 = ~w43 & ~w78;
assign w89 = w87 & w88;
assign w90 = ~w30 & ~w70;
assign w91 = ~a_22 & ~w40;
assign w92 = (w91 & ~w11) | (w91 & w5446) | (~w11 & w5446);
assign w93 = w13 & w5447;
assign w94 = a_22 & ~w33;
assign w95 = (~w94 & ~w11) | (~w94 & w5448) | (~w11 & w5448);
assign w96 = ~w92 & w95;
assign w97 = ~a_20 & a_21;
assign w98 = ~a_22 & w97;
assign w99 = (w98 & ~w11) | (w98 & w5449) | (~w11 & w5449);
assign w100 = w45 & w72;
assign w101 = w11 & w100;
assign w102 = a_22 & w49;
assign w103 = ~w101 & ~w102;
assign w104 = ~w99 & w103;
assign w105 = w96 & ~w104;
assign w106 = w90 & w105;
assign w107 = ~w89 & ~w106;
assign w108 = ~w56 & w96;
assign w109 = w87 & w108;
assign w110 = ~a_22 & w61;
assign w111 = (w110 & ~w11) | (w110 & w5450) | (~w11 & w5450);
assign w112 = w36 & w40;
assign w113 = w11 & w112;
assign w114 = a_22 & w37;
assign w115 = ~w113 & ~w114;
assign w116 = ~w111 & w115;
assign w117 = ~w56 & ~w116;
assign w118 = w30 & ~w70;
assign w119 = w117 & w118;
assign w120 = ~w109 & ~w119;
assign w121 = ~w78 & ~w116;
assign w122 = w31 & w121;
assign w123 = ~w56 & w65;
assign w124 = w31 & w123;
assign w125 = (w50 & ~w11) | (w50 & w5451) | (~w11 & w5451);
assign w126 = a_22 & w97;
assign w127 = w45 & w97;
assign w128 = w11 & w127;
assign w129 = ~w126 & ~w128;
assign w130 = ~w125 & w129;
assign w131 = ~w116 & ~w130;
assign w132 = ~w30 & ~w86;
assign w133 = w131 & w132;
assign w134 = ~a_22 & w82;
assign w135 = (w134 & ~w11) | (w134 & w5452) | (~w11 & w5452);
assign w136 = w13 & w66;
assign w137 = a_22 & w18;
assign w138 = (~w137 & ~w11) | (~w137 & w5453) | (~w11 & w5453);
assign w139 = ~w135 & w138;
assign w140 = ~w30 & ~w139;
assign w141 = w131 & w140;
assign w142 = ~w133 & ~w141;
assign w143 = ~w122 & ~w124;
assign w144 = w107 & w143;
assign w145 = w120 & w142;
assign w146 = w144 & w145;
assign w147 = w90 & w117;
assign w148 = ~w30 & ~w56;
assign w149 = ~w24 & w96;
assign w150 = w148 & w149;
assign w151 = ~w147 & ~w150;
assign w152 = w65 & ~w104;
assign w153 = w132 & w152;
assign w154 = w30 & ~w139;
assign w155 = w131 & w154;
assign w156 = ~w153 & ~w155;
assign w157 = ~w24 & w65;
assign w158 = w148 & w157;
assign w159 = w57 & w87;
assign w160 = w108 & w154;
assign w161 = ~w159 & ~w160;
assign w162 = ~w158 & w161;
assign w163 = w123 & w132;
assign w164 = w121 & w140;
assign w165 = ~w163 & ~w164;
assign w166 = w57 & w132;
assign w167 = ~w24 & ~w116;
assign w168 = ~w104 & w167;
assign w169 = ~w166 & ~w168;
assign w170 = w151 & w169;
assign w171 = w156 & w165;
assign w172 = w170 & w171;
assign w173 = w162 & w172;
assign w174 = ~w58 & ~w80;
assign w175 = w146 & w174;
assign w176 = w173 & w175;
assign w177 = ~w56 & w5454;
assign w178 = w105 & w118;
assign w179 = w121 & w132;
assign w180 = w117 & w132;
assign w181 = w118 & w121;
assign w182 = ~w43 & ~w86;
assign w183 = w79 & w182;
assign w184 = ~w181 & ~w183;
assign w185 = ~w180 & w184;
assign w186 = w87 & w117;
assign w187 = w118 & w152;
assign w188 = ~w104 & ~w116;
assign w189 = w132 & w188;
assign w190 = ~w187 & ~w189;
assign w191 = ~w177 & ~w178;
assign w192 = ~w179 & ~w186;
assign w193 = w191 & w192;
assign w194 = w190 & w193;
assign w195 = w185 & w194;
assign w196 = w108 & w118;
assign w197 = w117 & w140;
assign w198 = ~w196 & ~w197;
assign w199 = w31 & w117;
assign w200 = w152 & w154;
assign w201 = ~w199 & ~w200;
assign w202 = w198 & w201;
assign w203 = ~w30 & ~w104;
assign w204 = w71 & w203;
assign w205 = w108 & w140;
assign w206 = w71 & w148;
assign w207 = ~w204 & ~w205;
assign w208 = ~w206 & w207;
assign w209 = w96 & ~w130;
assign w210 = w118 & w209;
assign w211 = w121 & w154;
assign w212 = ~w210 & ~w211;
assign w213 = w88 & w118;
assign w214 = ~w30 & ~w130;
assign w215 = w149 & w214;
assign w216 = ~w213 & ~w215;
assign w217 = w118 & w131;
assign w218 = w90 & w121;
assign w219 = ~w217 & ~w218;
assign w220 = w212 & w216;
assign w221 = w219 & w220;
assign w222 = w202 & w208;
assign w223 = w221 & w222;
assign w224 = w195 & w223;
assign w225 = w176 & w224;
assign w226 = w154 & w209;
assign w227 = w87 & w123;
assign w228 = w132 & w209;
assign w229 = ~w227 & ~w228;
assign w230 = w31 & w108;
assign w231 = w108 & w132;
assign w232 = ~w230 & ~w231;
assign w233 = w229 & w232;
assign w234 = w140 & w209;
assign w235 = w117 & w154;
assign w236 = w57 & w140;
assign w237 = w87 & w121;
assign w238 = w31 & w88;
assign w239 = ~w24 & ~w43;
assign w240 = w30 & ~w130;
assign w241 = w239 & w240;
assign w242 = ~w238 & ~w241;
assign w243 = ~w234 & ~w235;
assign w244 = ~w236 & ~w237;
assign w245 = w243 & w244;
assign w246 = w242 & w245;
assign w247 = ~w226 & w233;
assign w248 = w246 & w247;
assign w249 = w87 & w188;
assign w250 = w148 & w239;
assign w251 = ~w249 & ~w250;
assign w252 = w87 & w209;
assign w253 = w140 & w152;
assign w254 = w57 & w154;
assign w255 = ~w253 & ~w254;
assign w256 = w57 & w118;
assign w257 = w214 & w239;
assign w258 = w90 & w108;
assign w259 = ~w257 & ~w258;
assign w260 = ~w256 & w259;
assign w261 = w251 & ~w252;
assign w262 = w255 & w261;
assign w263 = w260 & w262;
assign w264 = w90 & w131;
assign w265 = w57 & w90;
assign w266 = ~w264 & ~w265;
assign w267 = w154 & w188;
assign w268 = w149 & w240;
assign w269 = ~w267 & ~w268;
assign w270 = w118 & w123;
assign w271 = w148 & w167;
assign w272 = ~w270 & ~w271;
assign w273 = w88 & w154;
assign w274 = w272 & ~w273;
assign w275 = w90 & w209;
assign w276 = ~w43 & ~w139;
assign w277 = w79 & w276;
assign w278 = ~w275 & ~w277;
assign w279 = w79 & w239;
assign w280 = w79 & w167;
assign w281 = ~w279 & ~w280;
assign w282 = w266 & w281;
assign w283 = w269 & w278;
assign w284 = w282 & w283;
assign w285 = w274 & w284;
assign w286 = w248 & w285;
assign w287 = w263 & w286;
assign w288 = w225 & w287;
assign w289 = w65 & ~w130;
assign w290 = w87 & w289;
assign w291 = w182 & w214;
assign w292 = ~w80 & ~w290;
assign w293 = ~w291 & w292;
assign w294 = w156 & w293;
assign w295 = w65 & ~w78;
assign w296 = w87 & w295;
assign w297 = w118 & w188;
assign w298 = ~w250 & ~w297;
assign w299 = ~w204 & ~w253;
assign w300 = ~w296 & w299;
assign w301 = w298 & w300;
assign w302 = ~w206 & ~w268;
assign w303 = w157 & w240;
assign w304 = ~w217 & ~w303;
assign w305 = ~w186 & w304;
assign w306 = ~w43 & ~w104;
assign w307 = w31 & w306;
assign w308 = ~w43 & ~w70;
assign w309 = w79 & w308;
assign w310 = ~w307 & ~w309;
assign w311 = w302 & w310;
assign w312 = w305 & w311;
assign w313 = ~w78 & w96;
assign w314 = w31 & w313;
assign w315 = w31 & w105;
assign w316 = ~w238 & ~w314;
assign w317 = ~w315 & w316;
assign w318 = ~w58 & ~w124;
assign w319 = ~w227 & w318;
assign w320 = ~w178 & ~w254;
assign w321 = w79 & w157;
assign w322 = ~w200 & ~w321;
assign w323 = w57 & ~w70;
assign w324 = w157 & w214;
assign w325 = ~w264 & ~w323;
assign w326 = ~w324 & w325;
assign w327 = w320 & w322;
assign w328 = w326 & w327;
assign w329 = w87 & w313;
assign w330 = ~w179 & ~w329;
assign w331 = ~w279 & w330;
assign w332 = w117 & ~w139;
assign w333 = w330 & w5455;
assign w334 = ~w130 & w276;
assign w335 = ~w133 & ~w166;
assign w336 = w31 & w295;
assign w337 = w132 & w313;
assign w338 = ~w334 & ~w336;
assign w339 = ~w337 & w338;
assign w340 = w335 & w339;
assign w341 = w317 & w319;
assign w342 = w340 & w341;
assign w343 = w328 & w333;
assign w344 = w342 & w343;
assign w345 = ~w158 & ~w163;
assign w346 = w140 & w188;
assign w347 = w87 & w306;
assign w348 = ~w346 & ~w347;
assign w349 = ~w122 & ~w159;
assign w350 = w345 & w348;
assign w351 = w349 & w350;
assign w352 = w182 & w203;
assign w353 = ~w236 & ~w352;
assign w354 = w24 & ~w132;
assign w355 = w117 & ~w354;
assign w356 = w182 & w240;
assign w357 = ~w177 & ~w237;
assign w358 = ~w356 & w357;
assign w359 = w353 & ~w355;
assign w360 = w358 & w359;
assign w361 = w351 & w360;
assign w362 = w90 & w188;
assign w363 = ~w270 & ~w362;
assign w364 = w361 & w363;
assign w365 = w154 & w306;
assign w366 = w214 & w308;
assign w367 = ~w141 & ~w215;
assign w368 = ~w365 & ~w366;
assign w369 = w367 & w368;
assign w370 = ~w106 & ~w187;
assign w371 = w203 & w239;
assign w372 = w240 & w308;
assign w373 = w79 & w149;
assign w374 = ~w372 & ~w373;
assign w375 = ~w280 & ~w371;
assign w376 = w370 & w375;
assign w377 = w374 & w376;
assign w378 = w369 & w377;
assign w379 = w294 & w301;
assign w380 = w312 & w379;
assign w381 = w378 & w380;
assign w382 = w344 & w364;
assign w383 = w381 & w382;
assign w384 = w288 & w383;
assign w385 = ~w288 & ~w383;
assign w386 = ~w384 & ~w385;
assign w387 = ~a_22 & ~w0;
assign w388 = a_2 & ~a_22;
assign w389 = (a_3 & w387) | (a_3 & w5860) | (w387 & w5860);
assign w390 = ~w387 & w5861;
assign w391 = ~w389 & ~w390;
assign w392 = w386 & w391;
assign w393 = ~w118 & w139;
assign w394 = w306 & ~w393;
assign w395 = ~w104 & w157;
assign w396 = ~w347 & ~w395;
assign w397 = ~w394 & w396;
assign w398 = ~w133 & ~w371;
assign w399 = w397 & w398;
assign w400 = ~w210 & ~w268;
assign w401 = ~w228 & ~w275;
assign w402 = w203 & w308;
assign w403 = ~w226 & ~w402;
assign w404 = ~w252 & w400;
assign w405 = w401 & w403;
assign w406 = w404 & w405;
assign w407 = w399 & w406;
assign w408 = w295 & ~w393;
assign w409 = w132 & w295;
assign w410 = ~w307 & ~w352;
assign w411 = w87 & w152;
assign w412 = ~w215 & ~w234;
assign w413 = ~w411 & w412;
assign w414 = w410 & w413;
assign w415 = ~w213 & ~w273;
assign w416 = ~w155 & ~w217;
assign w417 = ~w141 & ~w264;
assign w418 = w416 & w417;
assign w419 = w88 & ~w354;
assign w420 = ~w178 & ~w277;
assign w421 = w107 & w420;
assign w422 = w415 & ~w419;
assign w423 = w421 & w422;
assign w424 = w418 & w423;
assign w425 = ~w309 & ~w321;
assign w426 = ~w296 & ~w336;
assign w427 = w425 & w426;
assign w428 = w423 & w5456;
assign w429 = ~w408 & ~w409;
assign w430 = w413 & w5457;
assign w431 = w407 & w430;
assign w432 = w428 & w431;
assign w433 = ~w385 & ~w432;
assign w434 = ~w392 & w433;
assign w435 = w167 & w214;
assign w436 = ~w296 & ~w435;
assign w437 = w276 & w214;
assign w438 = ~w58 & ~w147;
assign w439 = ~w205 & ~w270;
assign w440 = w438 & w439;
assign w441 = ~w437 & w440;
assign w442 = ~w104 & w5862;
assign w443 = ~w133 & ~w442;
assign w444 = w348 & w443;
assign w445 = ~w253 & ~w277;
assign w446 = ~w215 & w445;
assign w447 = ~w210 & ~w291;
assign w448 = ~w337 & w447;
assign w449 = ~w250 & ~w256;
assign w450 = ~w307 & w449;
assign w451 = w436 & w450;
assign w452 = w444 & w446;
assign w453 = w448 & w452;
assign w454 = w441 & w451;
assign w455 = w453 & w454;
assign w456 = w87 & w105;
assign w457 = w154 & w289;
assign w458 = w90 & w313;
assign w459 = ~w457 & ~w458;
assign w460 = w203 & w276;
assign w461 = ~w130 & w5863;
assign w462 = ~w89 & ~w411;
assign w463 = ~w297 & w5864;
assign w464 = w462 & w463;
assign w465 = w105 & w132;
assign w466 = ~w254 & ~w465;
assign w467 = w118 & w313;
assign w468 = w118 & w295;
assign w469 = ~w366 & ~w468;
assign w470 = w31 & w188;
assign w471 = ~w228 & ~w268;
assign w472 = ~w196 & ~w467;
assign w473 = ~w470 & w472;
assign w474 = w466 & w469;
assign w475 = w471 & w474;
assign w476 = w473 & w475;
assign w477 = w118 & w289;
assign w478 = ~w180 & ~w477;
assign w479 = ~w150 & ~w280;
assign w480 = w154 & w295;
assign w481 = ~w218 & ~w480;
assign w482 = ~w249 & ~w402;
assign w483 = ~w211 & ~w252;
assign w484 = w118 & w306;
assign w485 = ~w187 & ~w484;
assign w486 = w140 & w289;
assign w487 = ~w199 & ~w217;
assign w488 = ~w336 & ~w486;
assign w489 = w487 & w488;
assign w490 = w266 & w482;
assign w491 = w483 & w485;
assign w492 = w490 & w491;
assign w493 = w489 & w492;
assign w494 = ~w356 & ~w456;
assign w495 = ~w460 & w494;
assign w496 = w120 & w459;
assign w497 = w478 & w479;
assign w498 = w481 & w497;
assign w499 = w495 & w496;
assign w500 = w498 & w499;
assign w501 = w333 & w464;
assign w502 = w500 & w501;
assign w503 = w476 & w493;
assign w504 = w502 & w503;
assign w505 = w455 & w504;
assign w506 = (~a_22 & ~w5) | (~a_22 & w5865) | (~w5 & w5865);
assign w507 = (w5 & w7274) | (w5 & w7275) | (w7274 & w7275);
assign w508 = (w5 & w7276) | (w5 & w7277) | (w7276 & w7277);
assign w509 = (w506 & w5868) | (w506 & w5869) | (w5868 & w5869);
assign w510 = ~a_12 & w7864;
assign w511 = ~w509 & ~w510;
assign w512 = (~w511 & ~w504) | (~w511 & w5458) | (~w504 & w5458);
assign w513 = w149 & w203;
assign w514 = w132 & w289;
assign w515 = ~w513 & ~w514;
assign w516 = ~w186 & w515;
assign w517 = w90 & w289;
assign w518 = ~w356 & ~w517;
assign w519 = ~w196 & ~w206;
assign w520 = ~w279 & ~w315;
assign w521 = w519 & w520;
assign w522 = w161 & w278;
assign w523 = ~w437 & w518;
assign w524 = w522 & w523;
assign w525 = w369 & w521;
assign w526 = w516 & w525;
assign w527 = w524 & w526;
assign w528 = w140 & w313;
assign w529 = ~w267 & ~w528;
assign w530 = ~w265 & ~w297;
assign w531 = ~w106 & ~w253;
assign w532 = ~w122 & ~w153;
assign w533 = ~w178 & ~w213;
assign w534 = ~w458 & w533;
assign w535 = w400 & w532;
assign w536 = w531 & w535;
assign w537 = w534 & w536;
assign w538 = w240 & w276;
assign w539 = ~w150 & ~w372;
assign w540 = ~w227 & ~w538;
assign w541 = w345 & w540;
assign w542 = w539 & w541;
assign w543 = ~w337 & ~w373;
assign w544 = ~w307 & ~w324;
assign w545 = ~w226 & ~w252;
assign w546 = ~w457 & w545;
assign w547 = ~w235 & ~w371;
assign w548 = ~w280 & w543;
assign w549 = w544 & w547;
assign w550 = w548 & w549;
assign w551 = w546 & w550;
assign w552 = ~w197 & ~w211;
assign w553 = ~w218 & ~w230;
assign w554 = w552 & w553;
assign w555 = w184 & w529;
assign w556 = w530 & w555;
assign w557 = w554 & w556;
assign w558 = w542 & w557;
assign w559 = w537 & w551;
assign w560 = w558 & w559;
assign w561 = w527 & w560;
assign w562 = ~w505 & ~w561;
assign w563 = (~w512 & w562) | (~w512 & w5459) | (w562 & w5459);
assign w564 = a_11 & w7865;
assign w565 = ~w508 & ~w564;
assign w566 = (~w565 & ~w504) | (~w565 & w5460) | (~w504 & w5460);
assign w567 = w561 & ~w566;
assign w568 = ~w563 & ~w567;
assign w569 = w434 & w568;
assign w570 = ~w434 & ~w568;
assign w571 = ~w569 & ~w570;
assign w572 = (a_4 & w2) | (a_4 & w5870) | (w2 & w5870);
assign w573 = ~w2 & w5871;
assign w574 = ~w572 & ~w573;
assign w575 = w431 & w5872;
assign w576 = (~w574 & ~w431) | (~w574 & w5873) | (~w431 & w5873);
assign w577 = ~w575 & ~w576;
assign w578 = w386 & w577;
assign w579 = w288 & ~w432;
assign w580 = ~w385 & ~w579;
assign w581 = ~w383 & ~w391;
assign w582 = (w391 & ~w431) | (w391 & w5874) | (~w431 & w5874);
assign w583 = (~w582 & w383) | (~w582 & w5875) | (w383 & w5875);
assign w584 = ~w580 & w583;
assign w585 = ~w578 & ~w584;
assign w586 = w571 & ~w585;
assign w587 = ~w571 & w585;
assign w588 = w154 & w313;
assign w589 = ~w196 & ~w588;
assign w590 = ~w280 & ~w486;
assign w591 = ~w309 & ~w324;
assign w592 = ~w133 & ~w160;
assign w593 = w259 & w592;
assign w594 = w589 & w590;
assign w595 = w591 & w594;
assign w596 = w593 & w595;
assign w597 = ~w409 & ~w477;
assign w598 = w518 & w597;
assign w599 = ~w458 & ~w528;
assign w600 = ~w122 & ~w336;
assign w601 = ~w155 & ~w181;
assign w602 = ~w334 & ~w467;
assign w603 = w304 & w602;
assign w604 = w599 & w600;
assign w605 = w601 & w604;
assign w606 = w598 & w603;
assign w607 = w605 & w606;
assign w608 = w596 & w607;
assign w609 = w105 & w140;
assign w610 = ~w394 & ~w609;
assign w611 = ~w147 & ~w352;
assign w612 = ~w197 & ~w402;
assign w613 = w611 & w612;
assign w614 = ~w153 & ~w470;
assign w615 = w167 & w203;
assign w616 = ~w106 & ~w615;
assign w617 = ~w362 & ~w465;
assign w618 = w269 & w617;
assign w619 = w616 & w618;
assign w620 = w123 & w140;
assign w621 = ~w180 & ~w620;
assign w622 = ~w277 & ~w307;
assign w623 = ~w119 & ~w159;
assign w624 = ~w80 & w623;
assign w625 = ~w200 & ~w250;
assign w626 = w624 & w625;
assign w627 = w167 & w240;
assign w628 = ~w235 & ~w627;
assign w629 = ~w256 & w481;
assign w630 = ~w58 & ~w186;
assign w631 = w546 & w630;
assign w632 = w629 & w631;
assign w633 = ~w166 & ~w275;
assign w634 = ~w513 & w633;
assign w635 = w165 & w628;
assign w636 = w634 & w635;
assign w637 = w274 & w636;
assign w638 = w464 & w626;
assign w639 = w637 & w638;
assign w640 = w632 & w639;
assign w641 = ~w158 & ~w230;
assign w642 = w614 & w641;
assign w643 = w621 & w622;
assign w644 = w642 & w643;
assign w645 = w610 & w613;
assign w646 = w644 & w645;
assign w647 = w619 & w646;
assign w648 = w608 & w647;
assign w649 = w640 & w648;
assign w650 = ~w505 & ~w649;
assign w651 = w505 & w649;
assign w652 = ~w650 & ~w651;
assign w653 = ~w228 & ~w371;
assign w654 = w140 & w295;
assign w655 = ~w468 & ~w654;
assign w656 = w653 & w655;
assign w657 = ~w435 & ~w620;
assign w658 = w71 & ~w130;
assign w659 = ~w199 & ~w658;
assign w660 = ~w153 & ~w227;
assign w661 = ~w279 & ~w373;
assign w662 = w660 & w661;
assign w663 = w659 & w662;
assign w664 = ~w346 & ~w486;
assign w665 = ~w230 & w255;
assign w666 = w657 & w664;
assign w667 = w665 & w666;
assign w668 = w317 & w656;
assign w669 = w667 & w668;
assign w670 = w663 & w669;
assign w671 = ~w213 & ~w264;
assign w672 = ~w290 & ~w356;
assign w673 = ~w366 & w672;
assign w674 = w589 & w671;
assign w675 = w673 & w674;
assign w676 = ~w252 & ~w609;
assign w677 = ~w241 & ~w297;
assign w678 = w157 & w203;
assign w679 = ~w58 & ~w678;
assign w680 = ~w89 & w679;
assign w681 = ~w210 & ~w329;
assign w682 = ~w460 & w681;
assign w683 = ~w336 & w353;
assign w684 = w682 & w683;
assign w685 = ~w205 & ~w467;
assign w686 = ~w514 & w591;
assign w687 = w685 & w686;
assign w688 = w105 & w154;
assign w689 = ~w24 & w121;
assign w690 = ~w257 & ~w513;
assign w691 = w87 & w131;
assign w692 = ~w109 & ~w166;
assign w693 = ~w691 & w692;
assign w694 = ~w204 & ~w307;
assign w695 = w628 & w694;
assign w696 = w690 & w695;
assign w697 = w693 & w696;
assign w698 = ~w158 & ~w372;
assign w699 = ~w402 & ~w470;
assign w700 = ~w688 & ~w689;
assign w701 = w699 & w700;
assign w702 = w251 & w698;
assign w703 = w701 & w702;
assign w704 = w684 & w703;
assign w705 = w687 & w704;
assign w706 = w697 & w705;
assign w707 = ~w337 & ~w528;
assign w708 = w459 & w707;
assign w709 = w676 & w677;
assign w710 = w708 & w709;
assign w711 = w305 & w624;
assign w712 = w680 & w711;
assign w713 = w675 & w710;
assign w714 = w712 & w713;
assign w715 = w670 & w714;
assign w716 = w706 & w715;
assign w717 = (w5 & w6596) | (w5 & w6597) | (w6596 & w6597);
assign w718 = ~a_9 & w7866;
assign w719 = (w5 & w6598) | (w5 & w6599) | (w6598 & w6599);
assign w720 = ~w718 & ~w719;
assign w721 = ~w716 & ~w720;
assign w722 = w716 & w720;
assign w723 = ~w721 & ~w722;
assign w724 = w652 & ~w723;
assign w725 = a_8 & w7746;
assign w726 = ~w717 & ~w725;
assign w727 = w716 & w726;
assign w728 = w650 & ~w727;
assign w729 = ~w716 & ~w726;
assign w730 = w651 & ~w729;
assign w731 = ~w728 & ~w730;
assign w732 = ~w724 & w731;
assign w733 = (~w566 & w562) | (~w566 & w5461) | (w562 & w5461);
assign w734 = a_10 & w506;
assign w735 = ~w507 & ~w734;
assign w736 = (~w735 & ~w504) | (~w735 & w5462) | (~w504 & w5462);
assign w737 = w561 & ~w736;
assign w738 = ~w733 & ~w737;
assign w739 = w732 & w738;
assign w740 = ~w732 & ~w738;
assign w741 = ~w291 & ~w460;
assign w742 = ~w241 & w741;
assign w743 = ~w234 & w320;
assign w744 = w742 & w743;
assign w745 = w441 & w744;
assign w746 = ~w186 & ~w231;
assign w747 = ~w408 & w746;
assign w748 = w653 & w747;
assign w749 = ~w166 & ~w250;
assign w750 = ~w365 & w749;
assign w751 = ~w80 & ~w206;
assign w752 = ~w280 & ~w323;
assign w753 = w751 & w752;
assign w754 = w750 & w753;
assign w755 = w748 & w754;
assign w756 = w745 & w755;
assign w757 = ~w249 & ~w678;
assign w758 = ~w324 & w757;
assign w759 = ~w217 & ~w321;
assign w760 = w758 & w759;
assign w761 = ~w210 & ~w236;
assign w762 = ~w238 & ~w513;
assign w763 = ~w409 & w436;
assign w764 = w518 & w761;
assign w765 = w762 & w764;
assign w766 = w763 & w765;
assign w767 = ~w366 & ~w514;
assign w768 = ~w315 & ~w362;
assign w769 = w31 & w152;
assign w770 = ~w200 & ~w268;
assign w771 = ~w769 & w770;
assign w772 = ~w159 & ~w615;
assign w773 = w767 & w772;
assign w774 = w768 & w773;
assign w775 = w771 & w774;
assign w776 = ~w253 & ~w279;
assign w777 = ~w486 & w776;
assign w778 = w621 & w777;
assign w779 = w146 & w778;
assign w780 = w760 & w779;
assign w781 = w766 & w775;
assign w782 = w780 & w781;
assign w783 = w756 & w782;
assign w784 = ~w716 & ~w783;
assign w785 = w716 & w783;
assign w786 = ~w784 & ~w785;
assign w787 = ~w178 & w416;
assign w788 = ~w303 & ~w588;
assign w789 = ~w153 & ~w457;
assign w790 = w788 & w789;
assign w791 = ~w183 & ~w329;
assign w792 = ~w89 & ~w688;
assign w793 = ~w189 & ~w253;
assign w794 = w751 & w793;
assign w795 = w792 & w794;
assign w796 = ~w456 & ~w484;
assign w797 = ~w470 & ~w620;
assign w798 = w791 & w797;
assign w799 = w796 & w798;
assign w800 = w787 & w790;
assign w801 = w799 & w800;
assign w802 = w795 & w801;
assign w803 = ~w130 & w182;
assign w804 = ~w409 & ~w460;
assign w805 = ~w230 & ~w258;
assign w806 = ~w309 & ~w362;
assign w807 = w685 & w806;
assign w808 = w804 & w805;
assign w809 = w807 & w808;
assign w810 = ~w314 & ~w627;
assign w811 = ~w234 & ~w252;
assign w812 = ~w119 & ~w196;
assign w813 = ~w249 & w812;
assign w814 = ~w199 & ~w321;
assign w815 = w762 & ~w769;
assign w816 = w814 & w815;
assign w817 = ~w187 & ~w237;
assign w818 = ~w133 & ~w346;
assign w819 = w272 & w767;
assign w820 = w818 & w819;
assign w821 = ~w211 & ~w264;
assign w822 = ~w181 & w821;
assign w823 = ~w277 & ~w517;
assign w824 = ~w654 & w823;
assign w825 = w410 & w479;
assign w826 = w817 & w825;
assign w827 = w822 & w824;
assign w828 = w826 & w827;
assign w829 = w820 & w828;
assign w830 = ~w147 & ~w538;
assign w831 = ~w803 & w830;
assign w832 = w810 & w811;
assign w833 = w831 & w832;
assign w834 = w813 & w833;
assign w835 = w809 & w816;
assign w836 = w834 & w835;
assign w837 = w802 & w836;
assign w838 = w829 & w837;
assign w839 = w716 & ~w838;
assign w840 = ~w716 & w838;
assign w841 = ~w839 & ~w840;
assign w842 = ~w786 & ~w841;
assign w843 = a_5 & ~a_22;
assign w844 = (w2 & w5879) | (w2 & w5880) | (w5879 & w5880);
assign w845 = a_6 & ~w844;
assign w846 = ~a_6 & w844;
assign w847 = ~w845 & ~w846;
assign w848 = w716 & w847;
assign w849 = ~w716 & ~w847;
assign w850 = ~w848 & ~w849;
assign w851 = w842 & w850;
assign w852 = ~w5 & w5881;
assign w853 = (a_7 & w5) | (a_7 & w5882) | (w5 & w5882);
assign w854 = ~w852 & ~w853;
assign w855 = w837 & w5463;
assign w856 = (~w854 & ~w837) | (~w854 & w5883) | (~w837 & w5883);
assign w857 = ~w855 & ~w856;
assign w858 = w786 & w857;
assign w859 = ~w851 & ~w858;
assign w860 = ~w740 & ~w859;
assign w861 = ~w739 & ~w860;
assign w862 = ~w587 & ~w861;
assign w863 = ~w586 & ~w862;
assign w864 = w383 & w574;
assign w865 = ~w383 & ~w574;
assign w866 = ~w864 & ~w865;
assign w867 = w577 & ~w866;
assign w868 = ~w386 & ~w867;
assign w869 = ~a_5 & w7747;
assign w870 = (w2 & w5884) | (w2 & w5885) | (w5884 & w5885);
assign w871 = ~w869 & ~w870;
assign w872 = w431 & w5886;
assign w873 = ~w384 & ~w872;
assign w874 = (w871 & ~w431) | (w871 & w5887) | (~w431 & w5887);
assign w875 = ~w385 & ~w874;
assign w876 = w873 & w875;
assign w877 = ~w868 & ~w876;
assign w878 = (~a_13 & w11) | (~a_13 & w5888) | (w11 & w5888);
assign w879 = ~w11 & w5889;
assign w880 = ~w878 & ~w879;
assign w881 = (~w880 & ~w504) | (~w880 & w5464) | (~w504 & w5464);
assign w882 = (~w881 & w562) | (~w881 & w5465) | (w562 & w5465);
assign w883 = ~w512 & w561;
assign w884 = ~w882 & ~w883;
assign w885 = w565 & ~w716;
assign w886 = ~w565 & w716;
assign w887 = ~w885 & ~w886;
assign w888 = w652 & w887;
assign w889 = w649 & ~w716;
assign w890 = ~w650 & ~w889;
assign w891 = ~w716 & w735;
assign w892 = ~w736 & ~w891;
assign w893 = ~w890 & w892;
assign w894 = ~w888 & ~w893;
assign w895 = w884 & ~w894;
assign w896 = ~w884 & w894;
assign w897 = ~w895 & ~w896;
assign w898 = ~w877 & w897;
assign w899 = w877 & ~w897;
assign w900 = ~w898 & ~w899;
assign w901 = ~w863 & ~w900;
assign w902 = w863 & w900;
assign w903 = ~w901 & ~w902;
assign w904 = ~w297 & ~w442;
assign w905 = ~w465 & ~w513;
assign w906 = w904 & w905;
assign w907 = ~w456 & w768;
assign w908 = w906 & w907;
assign w909 = ~w200 & ~w204;
assign w910 = ~w267 & ~w615;
assign w911 = ~w249 & ~w253;
assign w912 = w190 & w911;
assign w913 = w614 & w909;
assign w914 = w910 & w913;
assign w915 = w912 & w914;
assign w916 = ~w346 & w908;
assign w917 = w915 & w916;
assign w918 = w414 & w418;
assign w919 = w407 & w918;
assign w920 = (w919 & ~w432) | (w919 & w5466) | (~w432 & w5466);
assign w921 = w391 & w920;
assign w922 = ~w373 & ~w528;
assign w923 = w348 & w922;
assign w924 = ~w226 & ~w409;
assign w925 = w483 & w924;
assign w926 = w923 & w925;
assign w927 = w796 & w926;
assign w928 = ~w273 & ~w314;
assign w929 = w741 & w928;
assign w930 = ~w256 & ~w457;
assign w931 = ~w486 & ~w538;
assign w932 = ~w236 & ~w477;
assign w933 = ~w254 & w515;
assign w934 = ~w265 & ~w437;
assign w935 = w123 & w154;
assign w936 = ~w371 & ~w480;
assign w937 = ~w200 & ~w372;
assign w938 = ~w183 & ~w356;
assign w939 = ~w402 & ~w935;
assign w940 = w938 & w939;
assign w941 = w310 & w936;
assign w942 = w937 & w941;
assign w943 = w233 & w940;
assign w944 = w933 & w934;
assign w945 = w943 & w944;
assign w946 = w942 & w945;
assign w947 = ~w178 & ~w336;
assign w948 = ~w465 & ~w588;
assign w949 = w947 & w948;
assign w950 = w298 & w930;
assign w951 = w931 & w932;
assign w952 = w950 & w951;
assign w953 = w929 & w949;
assign w954 = w952 & w953;
assign w955 = w927 & w954;
assign w956 = w176 & w955;
assign w957 = w946 & w956;
assign w958 = ~w838 & ~w957;
assign w959 = w838 & w957;
assign w960 = ~w958 & ~w959;
assign w961 = w383 & w847;
assign w962 = ~w383 & ~w847;
assign w963 = ~w961 & ~w962;
assign w964 = w960 & w963;
assign w965 = w383 & ~w871;
assign w966 = w958 & ~w965;
assign w967 = ~w383 & w871;
assign w968 = w959 & ~w967;
assign w969 = ~w966 & ~w968;
assign w970 = ~w964 & w969;
assign w971 = w716 & ~w735;
assign w972 = ~w891 & ~w971;
assign w973 = w652 & w972;
assign w974 = (w720 & ~w504) | (w720 & w5467) | (~w504 & w5467);
assign w975 = ~w721 & ~w974;
assign w976 = ~w890 & w975;
assign w977 = ~w973 & ~w976;
assign w978 = ~w970 & w977;
assign w979 = (~w726 & ~w837) | (~w726 & w5468) | (~w837 & w5468);
assign w980 = w837 & w5469;
assign w981 = ~w979 & ~w980;
assign w982 = w786 & ~w981;
assign w983 = w716 & w854;
assign w984 = ~w716 & ~w854;
assign w985 = ~w983 & ~w984;
assign w986 = w842 & ~w985;
assign w987 = ~w982 & ~w986;
assign w988 = w970 & ~w977;
assign w989 = w987 & ~w988;
assign w990 = (~w921 & w989) | (~w921 & w5470) | (w989 & w5470);
assign w991 = ~w989 & w5471;
assign w992 = ~w990 & ~w991;
assign w993 = w383 & ~w854;
assign w994 = ~w383 & w854;
assign w995 = ~w993 & ~w994;
assign w996 = w960 & w995;
assign w997 = w958 & ~w961;
assign w998 = w959 & ~w962;
assign w999 = ~w997 & ~w998;
assign w1000 = ~w996 & w999;
assign w1001 = w837 & w5472;
assign w1002 = (~w720 & ~w837) | (~w720 & w5473) | (~w837 & w5473);
assign w1003 = ~w1001 & ~w1002;
assign w1004 = w786 & ~w1003;
assign w1005 = w784 & ~w980;
assign w1006 = w785 & ~w979;
assign w1007 = ~w1005 & ~w1006;
assign w1008 = ~w1004 & w1007;
assign w1009 = ~w1000 & ~w1008;
assign w1010 = w1000 & w1008;
assign w1011 = ~w1009 & ~w1010;
assign w1012 = w569 & ~w1011;
assign w1013 = ~w569 & w1011;
assign w1014 = ~w1012 & ~w1013;
assign w1015 = ~w992 & w1014;
assign w1016 = w992 & ~w1014;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = w903 & w1017;
assign w1019 = (~w901 & ~w903) | (~w901 & w5890) | (~w903 & w5890);
assign w1020 = (~w11 & w5891) | (~w11 & w5892) | (w5891 & w5892);
assign w1021 = (w11 & w5893) | (w11 & w5894) | (w5893 & w5894);
assign w1022 = ~w1020 & ~w1021;
assign w1023 = (w1022 & ~w504) | (w1022 & w5474) | (~w504 & w5474);
assign w1024 = ~w562 & ~w1022;
assign w1025 = (~w1023 & w562) | (~w1023 & w5475) | (w562 & w5475);
assign w1026 = ~w147 & ~w186;
assign w1027 = ~w271 & ~w486;
assign w1028 = w1026 & w1027;
assign w1029 = ~w119 & ~w457;
assign w1030 = w659 & w1029;
assign w1031 = w1028 & w1030;
assign w1032 = ~w124 & ~w257;
assign w1033 = ~w323 & ~w803;
assign w1034 = w1032 & w1033;
assign w1035 = ~w56 & w5476;
assign w1036 = ~w24 & w57;
assign w1037 = ~w461 & w628;
assign w1038 = ~w435 & ~w691;
assign w1039 = ~w180 & w1038;
assign w1040 = ~w206 & ~w620;
assign w1041 = ~w324 & w1040;
assign w1042 = ~w197 & ~w270;
assign w1043 = ~w303 & w1042;
assign w1044 = w1037 & w1043;
assign w1045 = w1039 & w1041;
assign w1046 = w1044 & w1045;
assign w1047 = ~w230 & ~w366;
assign w1048 = ~w437 & w1047;
assign w1049 = w542 & w1048;
assign w1050 = ~w241 & ~w258;
assign w1051 = ~w166 & w1050;
assign w1052 = ~w56 & w276;
assign w1053 = ~w196 & ~w205;
assign w1054 = ~w935 & ~w1052;
assign w1055 = w1053 & w1054;
assign w1056 = w1051 & w1055;
assign w1057 = w1049 & w1056;
assign w1058 = ~w1035 & ~w1036;
assign w1059 = w161 & w1058;
assign w1060 = w1034 & w1059;
assign w1061 = w1031 & w1060;
assign w1062 = w1046 & w1061;
assign w1063 = w1057 & w1062;
assign w1064 = w561 & ~w881;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = ~w1025 & w1065;
assign w1067 = w1063 & w1064;
assign w1068 = ~w1023 & w1063;
assign w1069 = ~w1024 & w1068;
assign w1070 = ~w1067 & ~w1069;
assign w1071 = ~w1066 & w1070;
assign w1072 = w511 & ~w716;
assign w1073 = ~w511 & w716;
assign w1074 = ~w1072 & ~w1073;
assign w1075 = w652 & w1074;
assign w1076 = ~w566 & ~w885;
assign w1077 = ~w890 & w1076;
assign w1078 = ~w1075 & ~w1077;
assign w1079 = ~w391 & w1063;
assign w1080 = w432 & w5895;
assign w1081 = ~w920 & ~w1079;
assign w1082 = ~w1080 & w1081;
assign w1083 = ~w574 & ~w1063;
assign w1084 = w574 & w1063;
assign w1085 = ~w1083 & ~w1084;
assign w1086 = w920 & w1085;
assign w1087 = ~w1082 & ~w1086;
assign w1088 = ~w1078 & ~w1087;
assign w1089 = w1078 & w1087;
assign w1090 = ~w1088 & ~w1089;
assign w1091 = w1071 & ~w1090;
assign w1092 = ~w1071 & w1090;
assign w1093 = ~w1091 & ~w1092;
assign w1094 = (~w991 & w1014) | (~w991 & w5477) | (w1014 & w5477);
assign w1095 = ~w1093 & ~w1094;
assign w1096 = w1093 & w1094;
assign w1097 = ~w1095 & ~w1096;
assign w1098 = w837 & w5478;
assign w1099 = (~w735 & ~w837) | (~w735 & w5479) | (~w837 & w5479);
assign w1100 = ~w1098 & ~w1099;
assign w1101 = w786 & ~w1100;
assign w1102 = w842 & w1003;
assign w1103 = ~w1101 & ~w1102;
assign w1104 = ~w383 & w726;
assign w1105 = w383 & ~w726;
assign w1106 = ~w1104 & ~w1105;
assign w1107 = w960 & w1106;
assign w1108 = ~w383 & w957;
assign w1109 = ~w958 & ~w1108;
assign w1110 = ~w855 & ~w993;
assign w1111 = ~w1109 & ~w1110;
assign w1112 = ~w1107 & ~w1111;
assign w1113 = w431 & w5896;
assign w1114 = (~w847 & ~w431) | (~w847 & w5897) | (~w431 & w5897);
assign w1115 = ~w1113 & ~w1114;
assign w1116 = w386 & ~w1115;
assign w1117 = ~w873 & ~w875;
assign w1118 = ~w1116 & ~w1117;
assign w1119 = ~w1112 & ~w1118;
assign w1120 = w1112 & w1118;
assign w1121 = ~w1119 & ~w1120;
assign w1122 = w1103 & ~w1121;
assign w1123 = ~w1103 & ~w1120;
assign w1124 = ~w1119 & w1123;
assign w1125 = ~w1122 & ~w1124;
assign w1126 = ~w569 & ~w1010;
assign w1127 = ~w1009 & ~w1126;
assign w1128 = ~w877 & ~w895;
assign w1129 = ~w896 & ~w1128;
assign w1130 = w1127 & w1129;
assign w1131 = ~w1127 & ~w1129;
assign w1132 = ~w1130 & ~w1131;
assign w1133 = ~w1125 & w1132;
assign w1134 = w1125 & ~w1132;
assign w1135 = ~w1133 & ~w1134;
assign w1136 = w1097 & ~w1135;
assign w1137 = ~w1097 & w1135;
assign w1138 = ~w1136 & ~w1137;
assign w1139 = w1019 & ~w1138;
assign w1140 = w391 & w960;
assign w1141 = ~w383 & ~w958;
assign w1142 = ~w1140 & w1141;
assign w1143 = (~w736 & w562) | (~w736 & w5480) | (w562 & w5480);
assign w1144 = w561 & ~w974;
assign w1145 = ~w1143 & ~w1144;
assign w1146 = w1142 & w1145;
assign w1147 = ~w965 & ~w967;
assign w1148 = w960 & ~w1147;
assign w1149 = w383 & w958;
assign w1150 = ~w1141 & ~w1149;
assign w1151 = w837 & w5481;
assign w1152 = (~w574 & ~w837) | (~w574 & w5482) | (~w837 & w5482);
assign w1153 = ~w1151 & ~w1152;
assign w1154 = ~w960 & ~w1153;
assign w1155 = ~w1150 & w1154;
assign w1156 = ~w1148 & ~w1155;
assign w1157 = w1146 & ~w1156;
assign w1158 = ~w1146 & w1156;
assign w1159 = ~w1157 & ~w1158;
assign w1160 = w392 & w1159;
assign w1161 = (~w1157 & ~w1159) | (~w1157 & w5483) | (~w1159 & w5483);
assign w1162 = ~w978 & ~w988;
assign w1163 = w987 & ~w1162;
assign w1164 = ~w987 & w1162;
assign w1165 = ~w1163 & ~w1164;
assign w1166 = ~w1161 & w1165;
assign w1167 = w1161 & ~w1165;
assign w1168 = ~w1166 & ~w1167;
assign w1169 = ~w586 & ~w587;
assign w1170 = w861 & w1169;
assign w1171 = ~w861 & ~w1169;
assign w1172 = ~w1170 & ~w1171;
assign w1173 = w1168 & ~w1172;
assign w1174 = ~w1166 & ~w1173;
assign w1175 = ~w903 & ~w1017;
assign w1176 = ~w1018 & ~w1175;
assign w1177 = w1174 & ~w1176;
assign w1178 = ~w1139 & ~w1177;
assign w1179 = ~w1095 & ~w1136;
assign w1180 = w432 & w5898;
assign w1181 = w871 & w1063;
assign w1182 = ~w871 & ~w1063;
assign w1183 = ~w1181 & ~w1182;
assign w1184 = ~w920 & w1084;
assign w1185 = (~w1180 & w1183) | (~w1180 & w5899) | (w1183 & w5899);
assign w1186 = ~w1184 & w1185;
assign w1187 = w1066 & w1186;
assign w1188 = ~w1066 & ~w1186;
assign w1189 = ~w1187 & ~w1188;
assign w1190 = ~w1119 & ~w1123;
assign w1191 = (w1189 & w1123) | (w1189 & w5900) | (w1123 & w5900);
assign w1192 = ~w1123 & w5901;
assign w1193 = ~w1191 & ~w1192;
assign w1194 = ~w1125 & ~w1130;
assign w1195 = ~w1194 & w5902;
assign w1196 = (~w1193 & w1194) | (~w1193 & w5903) | (w1194 & w5903);
assign w1197 = ~w1195 & ~w1196;
assign w1198 = (~w565 & ~w837) | (~w565 & w5484) | (~w837 & w5484);
assign w1199 = w837 & w5485;
assign w1200 = ~w1198 & ~w1199;
assign w1201 = w786 & ~w1200;
assign w1202 = ~w785 & ~w1098;
assign w1203 = ~w784 & ~w1099;
assign w1204 = ~w1202 & ~w1203;
assign w1205 = ~w1201 & ~w1204;
assign w1206 = ~w383 & w720;
assign w1207 = w383 & ~w720;
assign w1208 = ~w1206 & ~w1207;
assign w1209 = w960 & ~w1208;
assign w1210 = ~w979 & ~w1104;
assign w1211 = ~w1109 & w1210;
assign w1212 = ~w1209 & ~w1211;
assign w1213 = w1205 & w1212;
assign w1214 = ~w1205 & ~w1212;
assign w1215 = ~w1213 & ~w1214;
assign w1216 = w431 & w5904;
assign w1217 = (~w854 & ~w431) | (~w854 & w5905) | (~w431 & w5905);
assign w1218 = ~w1216 & ~w1217;
assign w1219 = w386 & w1218;
assign w1220 = ~w386 & ~w1115;
assign w1221 = w963 & w1220;
assign w1222 = ~w1219 & ~w1221;
assign w1223 = w1215 & w1222;
assign w1224 = ~w1215 & ~w1222;
assign w1225 = ~w1223 & ~w1224;
assign w1226 = w391 & ~w1063;
assign w1227 = (w1226 & w562) | (w1226 & w5486) | (w562 & w5486);
assign w1228 = ~w562 & w5487;
assign w1229 = ~w1227 & ~w1228;
assign w1230 = w716 & ~w880;
assign w1231 = ~w716 & w880;
assign w1232 = ~w1230 & ~w1231;
assign w1233 = w652 & w1232;
assign w1234 = ~w512 & ~w1072;
assign w1235 = ~w890 & w1234;
assign w1236 = ~w1233 & ~w1235;
assign w1237 = w1229 & ~w1236;
assign w1238 = ~w1229 & w1236;
assign w1239 = ~w1237 & ~w1238;
assign w1240 = ~w1071 & ~w1088;
assign w1241 = ~w1089 & ~w1240;
assign w1242 = w1239 & w1241;
assign w1243 = ~w1239 & ~w1241;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = w1225 & ~w1244;
assign w1246 = ~w1225 & w1244;
assign w1247 = ~w1245 & ~w1246;
assign w1248 = w1197 & w1247;
assign w1249 = ~w1197 & ~w1247;
assign w1250 = ~w1248 & ~w1249;
assign w1251 = ~w1179 & w1250;
assign w1252 = ~w1019 & w1138;
assign w1253 = ~w1251 & ~w1252;
assign w1254 = ~w1178 & w1253;
assign w1255 = w1179 & ~w1250;
assign w1256 = (~w1195 & ~w1197) | (~w1195 & w5488) | (~w1197 & w5488);
assign w1257 = (~w1213 & ~w1215) | (~w1213 & w5489) | (~w1215 & w5489);
assign w1258 = (~w1227 & w1236) | (~w1227 & w5490) | (w1236 & w5490);
assign w1259 = w847 & ~w1063;
assign w1260 = ~w847 & w1063;
assign w1261 = ~w1259 & ~w1260;
assign w1262 = w920 & w1261;
assign w1263 = ~w872 & ~w1181;
assign w1264 = ~w920 & w1263;
assign w1265 = ~w1262 & ~w1264;
assign w1266 = w1258 & w1265;
assign w1267 = ~w1258 & ~w1265;
assign w1268 = ~w1266 & ~w1267;
assign w1269 = w1257 & ~w1268;
assign w1270 = ~w1257 & w1268;
assign w1271 = ~w1269 & ~w1270;
assign w1272 = w1225 & ~w1242;
assign w1273 = ~w1243 & ~w1272;
assign w1274 = ~w1271 & w1273;
assign w1275 = w1271 & ~w1273;
assign w1276 = ~w1274 & ~w1275;
assign w1277 = (~w1187 & w1190) | (~w1187 & w5491) | (w1190 & w5491);
assign w1278 = w505 & w716;
assign w1279 = ~w505 & ~w716;
assign w1280 = ~w1278 & ~w1279;
assign w1281 = w1232 & w1280;
assign w1282 = ~w652 & ~w1281;
assign w1283 = w505 & ~w1083;
assign w1284 = ~w505 & w1083;
assign w1285 = ~w1283 & ~w1284;
assign w1286 = w716 & w1022;
assign w1287 = ~w716 & ~w1022;
assign w1288 = ~w1286 & ~w1287;
assign w1289 = w652 & ~w1288;
assign w1290 = w1285 & ~w1289;
assign w1291 = ~w1282 & w1290;
assign w1292 = (~w1285 & w1282) | (~w1285 & w5906) | (w1282 & w5906);
assign w1293 = ~w1291 & ~w1292;
assign w1294 = w383 & ~w735;
assign w1295 = ~w383 & w735;
assign w1296 = ~w1294 & ~w1295;
assign w1297 = w960 & w1296;
assign w1298 = ~w1001 & ~w1207;
assign w1299 = ~w1109 & ~w1298;
assign w1300 = ~w1297 & ~w1299;
assign w1301 = w837 & w5492;
assign w1302 = (~w511 & ~w837) | (~w511 & w5493) | (~w837 & w5493);
assign w1303 = ~w1301 & ~w1302;
assign w1304 = w786 & ~w1303;
assign w1305 = ~w785 & ~w1199;
assign w1306 = ~w784 & ~w1198;
assign w1307 = ~w1305 & ~w1306;
assign w1308 = ~w1304 & ~w1307;
assign w1309 = ~w1300 & ~w1308;
assign w1310 = w1300 & w1308;
assign w1311 = ~w1309 & ~w1310;
assign w1312 = w431 & w5907;
assign w1313 = (w726 & ~w431) | (w726 & w5908) | (~w431 & w5908);
assign w1314 = ~w1312 & ~w1313;
assign w1315 = w386 & w1314;
assign w1316 = ~w386 & w1218;
assign w1317 = w995 & w1316;
assign w1318 = ~w1315 & ~w1317;
assign w1319 = ~w1311 & w1318;
assign w1320 = w1311 & ~w1318;
assign w1321 = ~w1319 & ~w1320;
assign w1322 = w1293 & w1321;
assign w1323 = ~w1293 & ~w1321;
assign w1324 = ~w1322 & ~w1323;
assign w1325 = w1277 & ~w1324;
assign w1326 = ~w1277 & w1324;
assign w1327 = ~w1325 & ~w1326;
assign w1328 = w1276 & w1327;
assign w1329 = ~w1276 & ~w1327;
assign w1330 = ~w1328 & ~w1329;
assign w1331 = ~w1256 & w1330;
assign w1332 = w1256 & ~w1330;
assign w1333 = ~w1331 & ~w1332;
assign w1334 = ~w1255 & w1333;
assign w1335 = ~w784 & ~w838;
assign w1336 = w391 & w786;
assign w1337 = w1335 & ~w1336;
assign w1338 = (~w726 & ~w504) | (~w726 & w5909) | (~w504 & w5909);
assign w1339 = (~w1338 & w562) | (~w1338 & w5910) | (w562 & w5910);
assign w1340 = (w854 & ~w504) | (w854 & w6600) | (~w504 & w6600);
assign w1341 = w561 & ~w1340;
assign w1342 = ~w1339 & ~w1341;
assign w1343 = w1337 & w1342;
assign w1344 = w1337 & w5911;
assign w1345 = (~w1140 & ~w1337) | (~w1140 & w5912) | (~w1337 & w5912);
assign w1346 = ~w1344 & ~w1345;
assign w1347 = w652 & ~w850;
assign w1348 = ~w652 & w1280;
assign w1349 = w716 & w871;
assign w1350 = ~w716 & ~w871;
assign w1351 = ~w1349 & ~w1350;
assign w1352 = w1348 & w1351;
assign w1353 = ~w1347 & ~w1352;
assign w1354 = w786 & w1153;
assign w1355 = w391 & w716;
assign w1356 = ~w391 & ~w716;
assign w1357 = ~w1355 & ~w1356;
assign w1358 = w842 & w1357;
assign w1359 = ~w1354 & ~w1358;
assign w1360 = ~w1353 & ~w1359;
assign w1361 = w1353 & w1359;
assign w1362 = ~w1337 & ~w1342;
assign w1363 = ~w1343 & ~w1362;
assign w1364 = ~w1361 & w1363;
assign w1365 = (w1346 & w1364) | (w1346 & w5913) | (w1364 & w5913);
assign w1366 = ~w1364 & w5914;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = (~w974 & w562) | (~w974 & w5915) | (w562 & w5915);
assign w1369 = w561 & ~w1338;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = w652 & w985;
assign w1372 = ~w850 & w1348;
assign w1373 = (w1370 & w1372) | (w1370 & w5916) | (w1372 & w5916);
assign w1374 = ~w1372 & w5917;
assign w1375 = ~w1373 & ~w1374;
assign w1376 = w786 & ~w838;
assign w1377 = w786 & w5918;
assign w1378 = w786 & w5919;
assign w1379 = w574 & w716;
assign w1380 = ~w574 & ~w716;
assign w1381 = ~w1379 & ~w1380;
assign w1382 = w1153 & ~w1381;
assign w1383 = ~w786 & ~w1382;
assign w1384 = ~w1377 & ~w1378;
assign w1385 = ~w1383 & w1384;
assign w1386 = w1375 & w1385;
assign w1387 = ~w1375 & ~w1385;
assign w1388 = ~w1386 & ~w1387;
assign w1389 = w1367 & w1388;
assign w1390 = ~w562 & ~w854;
assign w1391 = (~w847 & ~w504) | (~w847 & w5920) | (~w504 & w5920);
assign w1392 = w561 & ~w1391;
assign w1393 = (~w1392 & w1390) | (~w1392 & w5921) | (w1390 & w5921);
assign w1394 = w652 & w1351;
assign w1395 = w1348 & w1381;
assign w1396 = (w1393 & w1395) | (w1393 & w5922) | (w1395 & w5922);
assign w1397 = (~w1391 & w562) | (~w1391 & w5923) | (w562 & w5923);
assign w1398 = (w871 & ~w504) | (w871 & w6601) | (~w504 & w6601);
assign w1399 = w561 & ~w1398;
assign w1400 = ~w1397 & ~w1399;
assign w1401 = w391 & w652;
assign w1402 = ~w650 & ~w716;
assign w1403 = ~w1401 & w1402;
assign w1404 = w1400 & w1403;
assign w1405 = ~w1395 & w5924;
assign w1406 = ~w1396 & ~w1405;
assign w1407 = w1404 & w1406;
assign w1408 = (~w1396 & ~w1406) | (~w1396 & w5494) | (~w1406 & w5494);
assign w1409 = ~w1360 & ~w1361;
assign w1410 = ~w1363 & w1409;
assign w1411 = w1363 & ~w1409;
assign w1412 = ~w1410 & ~w1411;
assign w1413 = ~w1408 & ~w1412;
assign w1414 = ~w1404 & ~w1406;
assign w1415 = ~w1407 & ~w1414;
assign w1416 = w1336 & w1415;
assign w1417 = ~w1336 & ~w1415;
assign w1418 = w652 & w1381;
assign w1419 = w1348 & ~w1357;
assign w1420 = ~w1418 & ~w1419;
assign w1421 = ~w1400 & ~w1403;
assign w1422 = ~w1404 & ~w1421;
assign w1423 = w391 & ~w652;
assign w1424 = (w574 & ~w504) | (w574 & w5925) | (~w504 & w5925);
assign w1425 = (~w1424 & ~w652) | (~w1424 & w5927) | (~w652 & w5927);
assign w1426 = (~w1398 & w562) | (~w1398 & w6602) | (w562 & w6602);
assign w1427 = ~w1423 & ~w1426;
assign w1428 = ~w1425 & w1427;
assign w1429 = (~w1420 & w1422) | (~w1420 & w5928) | (w1422 & w5928);
assign w1430 = w1422 & w1428;
assign w1431 = ~w1429 & ~w1430;
assign w1432 = ~w1417 & ~w1431;
assign w1433 = ~w1413 & ~w1416;
assign w1434 = ~w1432 & w1433;
assign w1435 = ~w1367 & ~w1388;
assign w1436 = w1408 & w1412;
assign w1437 = ~w1435 & ~w1436;
assign w1438 = (~w1389 & w1434) | (~w1389 & w5929) | (w1434 & w5929);
assign w1439 = ~w1344 & ~w1365;
assign w1440 = ~w1142 & ~w1145;
assign w1441 = ~w1146 & ~w1440;
assign w1442 = (~w1373 & ~w1375) | (~w1373 & w5495) | (~w1375 & w5495);
assign w1443 = w1441 & ~w1442;
assign w1444 = ~w1441 & w1442;
assign w1445 = ~w1443 & ~w1444;
assign w1446 = ~w727 & ~w729;
assign w1447 = w652 & ~w1446;
assign w1448 = w985 & w1348;
assign w1449 = ~w1447 & ~w1448;
assign w1450 = w786 & w5496;
assign w1451 = w786 & w5497;
assign w1452 = ~w841 & ~w1351;
assign w1453 = ~w786 & ~w1452;
assign w1454 = ~w1450 & ~w1451;
assign w1455 = ~w1453 & w1454;
assign w1456 = ~w1449 & w1455;
assign w1457 = w1449 & ~w1455;
assign w1458 = ~w1456 & ~w1457;
assign w1459 = w958 & w5930;
assign w1460 = w866 & w960;
assign w1461 = w581 & w959;
assign w1462 = ~w1459 & ~w1461;
assign w1463 = ~w1460 & w1462;
assign w1464 = w1458 & ~w1463;
assign w1465 = ~w1458 & w1463;
assign w1466 = ~w1464 & ~w1465;
assign w1467 = w1445 & w1466;
assign w1468 = ~w1445 & ~w1466;
assign w1469 = ~w1467 & ~w1468;
assign w1470 = w1439 & ~w1469;
assign w1471 = ~w1438 & ~w1470;
assign w1472 = ~w1439 & w1469;
assign w1473 = ~w1443 & ~w1467;
assign w1474 = ~w739 & ~w740;
assign w1475 = ~w859 & w1474;
assign w1476 = w859 & ~w1474;
assign w1477 = ~w1475 & ~w1476;
assign w1478 = ~w1457 & ~w1463;
assign w1479 = ~w1456 & ~w1478;
assign w1480 = w1477 & ~w1479;
assign w1481 = ~w1477 & w1479;
assign w1482 = ~w1480 & ~w1481;
assign w1483 = ~w392 & ~w1159;
assign w1484 = ~w1160 & ~w1483;
assign w1485 = w1482 & w1484;
assign w1486 = ~w1482 & ~w1484;
assign w1487 = ~w1485 & ~w1486;
assign w1488 = ~w1473 & w1487;
assign w1489 = ~w1472 & ~w1488;
assign w1490 = w1473 & ~w1487;
assign w1491 = (~w1480 & ~w1482) | (~w1480 & w5931) | (~w1482 & w5931);
assign w1492 = ~w1168 & w1172;
assign w1493 = ~w1173 & ~w1492;
assign w1494 = w1491 & ~w1493;
assign w1495 = ~w1490 & ~w1494;
assign w1496 = (w1495 & w1471) | (w1495 & w5498) | (w1471 & w5498);
assign w1497 = ~w1491 & w1493;
assign w1498 = ~w1174 & w1176;
assign w1499 = ~w1497 & ~w1498;
assign w1500 = ~w1252 & w1499;
assign w1501 = w1499 & w1253;
assign w1502 = ~w1496 & w1501;
assign w1503 = ~w1254 & w1334;
assign w1504 = ~w206 & ~w234;
assign w1505 = ~w336 & ~w365;
assign w1506 = ~w197 & ~w935;
assign w1507 = ~w254 & ~w267;
assign w1508 = ~w228 & ~w237;
assign w1509 = ~w257 & w1508;
assign w1510 = w1507 & w1509;
assign w1511 = ~w56 & w157;
assign w1512 = ~w371 & w478;
assign w1513 = ~w179 & ~w1511;
assign w1514 = w1512 & w1513;
assign w1515 = ~w215 & ~w226;
assign w1516 = ~w362 & ~w689;
assign w1517 = w1515 & w1516;
assign w1518 = w1510 & w1517;
assign w1519 = w1514 & w1518;
assign w1520 = ~w164 & ~w296;
assign w1521 = w482 & w657;
assign w1522 = w909 & w1520;
assign w1523 = w1521 & w1522;
assign w1524 = w822 & w1523;
assign w1525 = ~w290 & ~w457;
assign w1526 = ~w654 & w1525;
assign w1527 = w462 & w616;
assign w1528 = w928 & w1504;
assign w1529 = w1505 & w1506;
assign w1530 = w1528 & w1529;
assign w1531 = w1526 & w1527;
assign w1532 = w742 & w1531;
assign w1533 = w1530 & w1532;
assign w1534 = w1524 & w1533;
assign w1535 = w1519 & w1534;
assign w1536 = w1503 & w5932;
assign w1537 = ~w1496 & w1500;
assign w1538 = ~w1251 & ~w1255;
assign w1539 = ~w1178 & ~w1252;
assign w1540 = w1538 & ~w1539;
assign w1541 = ~w1537 & w1540;
assign w1542 = ~w1251 & ~w1333;
assign w1543 = ~w1333 & w5933;
assign w1544 = ~w1541 & w1543;
assign w1545 = ~w1536 & ~w1544;
assign w1546 = (~w1538 & w1537) | (~w1538 & w5934) | (w1537 & w5934);
assign w1547 = ~w627 & ~w654;
assign w1548 = ~w164 & ~w204;
assign w1549 = ~w249 & ~w460;
assign w1550 = w1548 & w1549;
assign w1551 = w400 & w1547;
assign w1552 = w1550 & w1551;
assign w1553 = w319 & w1028;
assign w1554 = w1552 & w1553;
assign w1555 = w184 & ~w465;
assign w1556 = w749 & w5935;
assign w1557 = ~w267 & ~w517;
assign w1558 = ~w352 & ~w356;
assign w1559 = w1557 & w1558;
assign w1560 = ~w106 & ~w484;
assign w1561 = w198 & w1560;
assign w1562 = ~w122 & ~w258;
assign w1563 = w443 & w1562;
assign w1564 = w817 & w1563;
assign w1565 = w787 & w1559;
assign w1566 = w1561 & w1565;
assign w1567 = w1556 & w1564;
assign w1568 = w1566 & w1567;
assign w1569 = w330 & w1568;
assign w1570 = ~w290 & ~w678;
assign w1571 = ~w334 & w811;
assign w1572 = w1570 & w1571;
assign w1573 = w446 & w629;
assign w1574 = w790 & w1555;
assign w1575 = w1573 & w1574;
assign w1576 = w687 & w1572;
assign w1577 = w1575 & w1576;
assign w1578 = w1554 & w1577;
assign w1579 = w1569 & w1578;
assign w1580 = ~w1541 & w1579;
assign w1581 = ~w1546 & w1580;
assign w1582 = ~w1541 & w1542;
assign w1583 = (w1535 & ~w1503) | (w1535 & w5936) | (~w1503 & w5936);
assign w1584 = ~w1582 & w1583;
assign w1585 = ~w1581 & ~w1584;
assign w1586 = w1545 & ~w1585;
assign w1587 = (~w1331 & ~w1503) | (~w1331 & w5937) | (~w1503 & w5937);
assign w1588 = ~w1274 & ~w1328;
assign w1589 = w505 & ~w1182;
assign w1590 = ~w505 & w1182;
assign w1591 = ~w1589 & ~w1590;
assign w1592 = w1288 & w1348;
assign w1593 = w652 & ~w716;
assign w1594 = (w1591 & w1592) | (w1591 & w5499) | (w1592 & w5499);
assign w1595 = ~w1592 & w5938;
assign w1596 = ~w1594 & ~w1595;
assign w1597 = ~w1099 & ~w1295;
assign w1598 = ~w1109 & w1597;
assign w1599 = w383 & ~w565;
assign w1600 = ~w383 & w565;
assign w1601 = ~w1599 & ~w1600;
assign w1602 = w960 & w1601;
assign w1603 = ~w1598 & ~w1602;
assign w1604 = w837 & w5500;
assign w1605 = (w880 & ~w837) | (w880 & w5501) | (~w837 & w5501);
assign w1606 = ~w1604 & ~w1605;
assign w1607 = w786 & w1606;
assign w1608 = ~w785 & ~w1301;
assign w1609 = ~w784 & ~w1302;
assign w1610 = ~w1608 & ~w1609;
assign w1611 = ~w1607 & ~w1610;
assign w1612 = w1603 & w1611;
assign w1613 = ~w1603 & ~w1611;
assign w1614 = ~w1612 & ~w1613;
assign w1615 = w431 & w5939;
assign w1616 = (~w720 & ~w431) | (~w720 & w5940) | (~w431 & w5940);
assign w1617 = ~w1615 & ~w1616;
assign w1618 = w386 & w1617;
assign w1619 = ~w386 & w1314;
assign w1620 = ~w1106 & w1619;
assign w1621 = ~w1618 & ~w1620;
assign w1622 = w1614 & w1621;
assign w1623 = ~w1614 & ~w1621;
assign w1624 = ~w1622 & ~w1623;
assign w1625 = w1596 & ~w1624;
assign w1626 = ~w1596 & w1624;
assign w1627 = ~w1625 & ~w1626;
assign w1628 = ~w1266 & ~w1270;
assign w1629 = w1627 & w1628;
assign w1630 = ~w1627 & ~w1628;
assign w1631 = ~w1629 & ~w1630;
assign w1632 = w1277 & ~w1322;
assign w1633 = ~w854 & ~w1063;
assign w1634 = w854 & w1063;
assign w1635 = ~w1633 & ~w1634;
assign w1636 = w920 & w1635;
assign w1637 = w917 & w1113;
assign w1638 = ~w920 & ~w1260;
assign w1639 = ~w1637 & w1638;
assign w1640 = ~w1636 & ~w1639;
assign w1641 = ~w1291 & w5502;
assign w1642 = (~w1640 & w1291) | (~w1640 & w5941) | (w1291 & w5941);
assign w1643 = ~w1641 & ~w1642;
assign w1644 = ~w1310 & ~w1318;
assign w1645 = ~w1309 & ~w1644;
assign w1646 = ~w1643 & w1645;
assign w1647 = ~w1645 & w1643;
assign w1648 = ~w1646 & ~w1647;
assign w1649 = (~w1648 & w1632) | (~w1648 & w5942) | (w1632 & w5942);
assign w1650 = ~w1632 & w5943;
assign w1651 = ~w1649 & ~w1650;
assign w1652 = w1631 & ~w1651;
assign w1653 = ~w1631 & w1651;
assign w1654 = ~w1652 & ~w1653;
assign w1655 = w1588 & w1654;
assign w1656 = ~w1588 & ~w1654;
assign w1657 = ~w1655 & ~w1656;
assign w1658 = ~w80 & ~w470;
assign w1659 = w440 & w5944;
assign w1660 = ~w187 & ~w297;
assign w1661 = ~w279 & ~w411;
assign w1662 = w417 & w1661;
assign w1663 = w1050 & w1660;
assign w1664 = w1662 & w1663;
assign w1665 = ~w280 & ~w769;
assign w1666 = ~w189 & ~w588;
assign w1667 = ~w275 & ~w467;
assign w1668 = w910 & w1667;
assign w1669 = w1666 & w1668;
assign w1670 = ~w277 & ~w362;
assign w1671 = ~w238 & ~w296;
assign w1672 = ~w218 & ~w337;
assign w1673 = ~w402 & ~w609;
assign w1674 = w1672 & w1673;
assign w1675 = ~w480 & w928;
assign w1676 = w1505 & w1665;
assign w1677 = w1670 & w1671;
assign w1678 = w1676 & w1677;
assign w1679 = w656 & w1675;
assign w1680 = w1555 & w1674;
assign w1681 = w1679 & w1680;
assign w1682 = w1669 & w1678;
assign w1683 = w1681 & w1682;
assign w1684 = ~w196 & ~w231;
assign w1685 = ~w324 & ~w329;
assign w1686 = ~w517 & w1685;
assign w1687 = w302 & w1684;
assign w1688 = w459 & w931;
assign w1689 = w1687 & w1688;
assign w1690 = w1686 & w1689;
assign w1691 = w1664 & w1690;
assign w1692 = w361 & w697;
assign w1693 = w1659 & w1692;
assign w1694 = w1683 & w1691;
assign w1695 = w1693 & w1694;
assign w1696 = w1657 & ~w1695;
assign w1697 = ~w1657 & w1695;
assign w1698 = ~w1696 & ~w1697;
assign w1699 = w1587 & ~w1698;
assign w1700 = ~w1587 & w1698;
assign w1701 = ~w1699 & ~w1700;
assign w1702 = ~w1586 & ~w1701;
assign w1703 = w1586 & w1701;
assign w1704 = ~w1702 & ~w1703;
assign w1705 = w1545 & ~w1584;
assign w1706 = w1541 & ~w1579;
assign w1707 = ~w1538 & ~w1579;
assign w1708 = (w1707 & w1537) | (w1707 & w5945) | (w1537 & w5945);
assign w1709 = ~w1706 & ~w1708;
assign w1710 = ~w1581 & w1709;
assign w1711 = ~w1705 & w1710;
assign w1712 = ~w1704 & w1711;
assign w1713 = w1581 & ~w1705;
assign w1714 = w1545 & w1585;
assign w1715 = ~w1713 & ~w1714;
assign w1716 = (w1715 & w1704) | (w1715 & w5503) | (w1704 & w5503);
assign w1717 = (w1503 & w6584) | (w1503 & w6585) | (w6584 & w6585);
assign w1718 = (w5504 & ~w1503) | (w5504 & w6586) | (~w1503 & w6586);
assign w1719 = ~w1717 & ~w1718;
assign w1720 = w1503 & w5946;
assign w1721 = w1331 & ~w1655;
assign w1722 = ~w1656 & ~w1721;
assign w1723 = (~w1642 & w1645) | (~w1642 & w5947) | (w1645 & w5947);
assign w1724 = w431 & w6603;
assign w1725 = (~w735 & ~w431) | (~w735 & w5948) | (~w431 & w5948);
assign w1726 = ~w1724 & ~w1725;
assign w1727 = w386 & ~w1726;
assign w1728 = (~w1616 & w383) | (~w1616 & w5949) | (w383 & w5949);
assign w1729 = ~w580 & w1728;
assign w1730 = ~w1727 & ~w1729;
assign w1731 = w432 & w5950;
assign w1732 = w726 & ~w1063;
assign w1733 = ~w726 & w1063;
assign w1734 = ~w1732 & ~w1733;
assign w1735 = w920 & ~w1734;
assign w1736 = ~w920 & w1634;
assign w1737 = ~w1735 & w5505;
assign w1738 = w1730 & ~w1737;
assign w1739 = ~w1730 & w1737;
assign w1740 = ~w1738 & ~w1739;
assign w1741 = ~w1232 & w1606;
assign w1742 = ~w786 & ~w1741;
assign w1743 = w837 & w5506;
assign w1744 = ~w785 & ~w1743;
assign w1745 = (w1022 & ~w837) | (w1022 & w5507) | (~w837 & w5507);
assign w1746 = ~w784 & ~w1745;
assign w1747 = w1744 & w1746;
assign w1748 = ~w1742 & ~w1747;
assign w1749 = w1740 & w1748;
assign w1750 = ~w1740 & ~w1748;
assign w1751 = ~w1749 & ~w1750;
assign w1752 = (~w1612 & ~w1614) | (~w1612 & w5508) | (~w1614 & w5508);
assign w1753 = ~w1751 & ~w1752;
assign w1754 = w1751 & w1752;
assign w1755 = ~w1753 & ~w1754;
assign w1756 = w1723 & ~w1755;
assign w1757 = ~w1723 & w1755;
assign w1758 = ~w1756 & ~w1757;
assign w1759 = ~w1590 & ~w1594;
assign w1760 = (w1259 & w1280) | (w1259 & w5509) | (w1280 & w5509);
assign w1761 = ~w1280 & w5510;
assign w1762 = ~w1760 & ~w1761;
assign w1763 = w383 & ~w511;
assign w1764 = ~w383 & w511;
assign w1765 = ~w1763 & ~w1764;
assign w1766 = w960 & w1765;
assign w1767 = ~w960 & w1200;
assign w1768 = w1601 & w1767;
assign w1769 = ~w1766 & ~w1768;
assign w1770 = w1762 & ~w1769;
assign w1771 = ~w1762 & w1769;
assign w1772 = ~w1770 & ~w1771;
assign w1773 = ~w1759 & w1772;
assign w1774 = w1759 & ~w1772;
assign w1775 = ~w1773 & ~w1774;
assign w1776 = w1627 & w5511;
assign w1777 = ~w1625 & ~w1775;
assign w1778 = w1625 & w1775;
assign w1779 = ~w1777 & ~w1778;
assign w1780 = ~w1629 & w1779;
assign w1781 = ~w1776 & ~w1780;
assign w1782 = ~w1758 & ~w1781;
assign w1783 = w1758 & w1781;
assign w1784 = ~w1782 & ~w1783;
assign w1785 = w1631 & ~w1649;
assign w1786 = (~w1650 & ~w1631) | (~w1650 & w5951) | (~w1631 & w5951);
assign w1787 = ~w315 & ~w372;
assign w1788 = ~w179 & ~w480;
assign w1789 = ~w270 & ~w291;
assign w1790 = ~w213 & ~w230;
assign w1791 = ~w336 & ~w477;
assign w1792 = w1790 & w1791;
assign w1793 = w1787 & w1788;
assign w1794 = w1789 & w1793;
assign w1795 = w923 & w1792;
assign w1796 = w1794 & w1795;
assign w1797 = w1556 & w1664;
assign w1798 = w1796 & w1797;
assign w1799 = w1554 & w1798;
assign w1800 = w802 & w1799;
assign w1801 = ~w1785 & w5512;
assign w1802 = (w1800 & w1785) | (w1800 & w5513) | (w1785 & w5513);
assign w1803 = ~w1801 & ~w1802;
assign w1804 = w1784 & w1803;
assign w1805 = ~w1784 & ~w1803;
assign w1806 = ~w1804 & ~w1805;
assign w1807 = w1722 & w1806;
assign w1808 = ~w1722 & ~w1806;
assign w1809 = ~w1807 & ~w1808;
assign w1810 = w1720 & ~w1809;
assign w1811 = ~w1720 & w1809;
assign w1812 = ~w1810 & ~w1811;
assign w1813 = w1719 & ~w1812;
assign w1814 = ~w1719 & w1812;
assign w1815 = ~w1813 & ~w1814;
assign w1816 = w1703 & w1815;
assign w1817 = ~w1703 & ~w1815;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = ~w1716 & w1818;
assign w1820 = ~w1586 & w5514;
assign w1821 = ~w1816 & ~w1820;
assign w1822 = ~w1819 & w1821;
assign w1823 = ~w1702 & w1815;
assign w1824 = ~w1820 & ~w1823;
assign w1825 = ~w1254 & ~w1502;
assign w1826 = w1333 & w5952;
assign w1827 = w1825 & w1826;
assign w1828 = w1722 & w5515;
assign w1829 = ~w1827 & w1828;
assign w1830 = ~w1784 & ~w1786;
assign w1831 = w1784 & w1786;
assign w1832 = ~w1830 & ~w1831;
assign w1833 = w1800 & ~w1832;
assign w1834 = w1826 & w1833;
assign w1835 = w1825 & w1834;
assign w1836 = ~w1722 & w1833;
assign w1837 = ~w1835 & ~w1836;
assign w1838 = ~w1829 & w1837;
assign w1839 = ~w1813 & w1838;
assign w1840 = ~w1701 & w1838;
assign w1841 = ~w1586 & w1840;
assign w1842 = ~w1839 & ~w1841;
assign w1843 = (~w1770 & ~w1772) | (~w1770 & w5693) | (~w1772 & w5693);
assign w1844 = w1723 & ~w1754;
assign w1845 = (w1843 & w1844) | (w1843 & w5516) | (w1844 & w5516);
assign w1846 = ~w1844 & w5517;
assign w1847 = ~w1845 & ~w1846;
assign w1848 = (~w1739 & ~w1740) | (~w1739 & w5518) | (~w1740 & w5518);
assign w1849 = ~w1744 & ~w1746;
assign w1850 = ~w1376 & ~w1849;
assign w1851 = ~w1633 & ~w1850;
assign w1852 = w1633 & w1850;
assign w1853 = ~w1851 & ~w1852;
assign w1854 = w383 & w880;
assign w1855 = ~w383 & ~w880;
assign w1856 = ~w1854 & ~w1855;
assign w1857 = w960 & ~w1856;
assign w1858 = ~w960 & w1303;
assign w1859 = w1765 & w1858;
assign w1860 = ~w1857 & ~w1859;
assign w1861 = ~w1853 & w1860;
assign w1862 = w1853 & ~w1860;
assign w1863 = ~w1861 & ~w1862;
assign w1864 = ~w1848 & w1863;
assign w1865 = w1848 & ~w1863;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = ~w1278 & ~w1760;
assign w1868 = (~w1724 & ~w383) | (~w1724 & w6604) | (~w383 & w6604);
assign w1869 = ~w580 & ~w1868;
assign w1870 = w431 & w5953;
assign w1871 = (~w565 & ~w431) | (~w565 & w5954) | (~w431 & w5954);
assign w1872 = ~w1870 & ~w1871;
assign w1873 = w386 & ~w1872;
assign w1874 = ~w1869 & ~w1873;
assign w1875 = w432 & w5955;
assign w1876 = w720 & w1063;
assign w1877 = ~w720 & ~w1063;
assign w1878 = ~w1876 & ~w1877;
assign w1879 = w920 & ~w1878;
assign w1880 = ~w920 & w1733;
assign w1881 = ~w1879 & w5519;
assign w1882 = w1874 & ~w1881;
assign w1883 = ~w1874 & w1881;
assign w1884 = ~w1882 & ~w1883;
assign w1885 = ~w1867 & ~w1884;
assign w1886 = w1867 & w1884;
assign w1887 = ~w1885 & ~w1886;
assign w1888 = w1866 & ~w1887;
assign w1889 = ~w1866 & w1887;
assign w1890 = ~w1888 & ~w1889;
assign w1891 = w1847 & ~w1890;
assign w1892 = ~w1847 & w1890;
assign w1893 = ~w1891 & ~w1892;
assign w1894 = ~w1629 & w1777;
assign w1895 = (~w1894 & w1781) | (~w1894 & w5520) | (w1781 & w5520);
assign w1896 = ~w1893 & w1895;
assign w1897 = ~w1830 & ~w1896;
assign w1898 = w1722 & w1897;
assign w1899 = ~w241 & ~w365;
assign w1900 = ~w160 & ~w314;
assign w1901 = ~w179 & ~w435;
assign w1902 = w142 & w1901;
assign w1903 = w479 & w1899;
assign w1904 = w1900 & w1903;
assign w1905 = w1902 & w1904;
assign w1906 = w684 & w1905;
assign w1907 = ~w337 & ~w437;
assign w1908 = ~w620 & ~w627;
assign w1909 = ~w180 & ~w257;
assign w1910 = w462 & w1909;
assign w1911 = w1910 & w5956;
assign w1912 = ~w279 & ~w409;
assign w1913 = w229 & w1912;
assign w1914 = ~w324 & ~w347;
assign w1915 = ~w356 & ~w480;
assign w1916 = w1914 & w1915;
assign w1917 = w184 & w1916;
assign w1918 = w1913 & w1917;
assign w1919 = w294 & w619;
assign w1920 = w1918 & w1919;
assign w1921 = w349 & ~w514;
assign w1922 = w1920 & w1921;
assign w1923 = ~w395 & ~w1036;
assign w1924 = w304 & w1923;
assign w1925 = w445 & w547;
assign w1926 = w817 & w1925;
assign w1927 = w1924 & w1926;
assign w1928 = w1911 & w1927;
assign w1929 = w1906 & w1928;
assign w1930 = w1922 & w1929;
assign w1931 = w1893 & ~w1895;
assign w1932 = ~w1896 & ~w1931;
assign w1933 = ~w1831 & w1932;
assign w1934 = ~w1930 & w1933;
assign w1935 = (w1934 & w1827) | (w1934 & w5521) | (w1827 & w5521);
assign w1936 = w1334 & w5694;
assign w1937 = w1825 & w1936;
assign w1938 = (~w1831 & w1721) | (~w1831 & w5695) | (w1721 & w5695);
assign w1939 = ~w1830 & ~w1932;
assign w1940 = ~w1930 & w1939;
assign w1941 = ~w1937 & w5522;
assign w1942 = ~w1935 & ~w1941;
assign w1943 = w1930 & ~w1933;
assign w1944 = (w1930 & w1784) | (w1930 & w5957) | (w1784 & w5957);
assign w1945 = w1722 & w1944;
assign w1946 = (~w1943 & w1827) | (~w1943 & w5523) | (w1827 & w5523);
assign w1947 = (w5696 & w5958) | (w5696 & w5959) | (w5958 & w5959);
assign w1948 = ~w1946 & ~w1947;
assign w1949 = w1942 & ~w1948;
assign w1950 = (w1949 & w1841) | (w1949 & w5960) | (w1841 & w5960);
assign w1951 = ~w1841 & w5961;
assign w1952 = ~w1950 & ~w1951;
assign w1953 = ~w1824 & ~w1952;
assign w1954 = w1824 & w1952;
assign w1955 = ~w1953 & ~w1954;
assign w1956 = ~w1822 & w1955;
assign w1957 = ~w720 & ~w726;
assign w1958 = w720 & w726;
assign w1959 = ~w1957 & ~w1958;
assign w1960 = w565 & ~w735;
assign w1961 = ~w565 & w735;
assign w1962 = ~w1960 & ~w1961;
assign w1963 = ~w1959 & ~w1962;
assign w1964 = w1955 & w5524;
assign w1965 = ~w1816 & w5962;
assign w1966 = ~w1819 & w1965;
assign w1967 = ~w1955 & w1966;
assign w1968 = ~w1959 & w1962;
assign w1969 = w1952 & w1968;
assign w1970 = w720 & w735;
assign w1971 = ~w720 & ~w735;
assign w1972 = ~w1970 & ~w1971;
assign w1973 = w1959 & ~w1962;
assign w1974 = w1972 & w1973;
assign w1975 = w1704 & w1974;
assign w1976 = w1959 & ~w1972;
assign w1977 = ~w1823 & w5525;
assign w1978 = ~w1975 & ~w1977;
assign w1979 = ~w1969 & w1978;
assign w1980 = ~w1967 & w1979;
assign w1981 = ~w511 & w565;
assign w1982 = w511 & ~w565;
assign w1983 = ~w1981 & ~w1982;
assign w1984 = w880 & w1022;
assign w1985 = ~w880 & ~w1022;
assign w1986 = ~w1984 & ~w1985;
assign w1987 = ~w1983 & w1986;
assign w1988 = ~w511 & ~w880;
assign w1989 = w511 & w880;
assign w1990 = ~w1988 & ~w1989;
assign w1991 = w1983 & w1990;
assign w1992 = ~w1710 & w1991;
assign w1993 = (~w1992 & ~w1715) | (~w1992 & w5526) | (~w1715 & w5526);
assign w1994 = ~w1983 & ~w1986;
assign w1995 = ~w1705 & w1709;
assign w1996 = w1705 & ~w1709;
assign w1997 = ~w1995 & ~w1996;
assign w1998 = w1994 & ~w1997;
assign w1999 = w1993 & ~w1998;
assign w2000 = ~w1710 & w1982;
assign w2001 = ~w1710 & w1981;
assign w2002 = ~w2000 & ~w2001;
assign w2003 = ~w1022 & ~w2002;
assign w2004 = ~w1999 & w2003;
assign w2005 = w1999 & ~w2003;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = w565 & w2006;
assign w2008 = w1980 & w5527;
assign w2009 = ~w565 & w2006;
assign w2010 = (w2009 & ~w1980) | (w2009 & w5528) | (~w1980 & w5528);
assign w2011 = ~w2008 & ~w2010;
assign w2012 = w565 & ~w2006;
assign w2013 = (w2012 & ~w1980) | (w2012 & w5529) | (~w1980 & w5529);
assign w2014 = (~w565 & w2002) | (~w565 & w5963) | (w2002 & w5963);
assign w2015 = w1999 & w2014;
assign w2016 = ~w1710 & w5964;
assign w2017 = ~w1999 & w2016;
assign w2018 = ~w2015 & ~w2017;
assign w2019 = w1979 & ~w2018;
assign w2020 = ~w1967 & w2019;
assign w2021 = ~w1964 & w2020;
assign w2022 = ~w2013 & ~w2021;
assign w2023 = w2011 & w2022;
assign w2024 = w1716 & ~w1818;
assign w2025 = w1963 & w2024;
assign w2026 = w1818 & w1963;
assign w2027 = ~w1716 & w2026;
assign w2028 = ~w1823 & w5530;
assign w2029 = w1704 & w1976;
assign w2030 = w1715 & w1974;
assign w2031 = ~w2029 & ~w2030;
assign w2032 = ~w2028 & w2031;
assign w2033 = ~w2027 & w2032;
assign w2034 = ~w2025 & w2033;
assign w2035 = w1704 & ~w1711;
assign w2036 = ~w1712 & ~w2035;
assign w2037 = w1963 & ~w2036;
assign w2038 = w1704 & w1968;
assign w2039 = ~w1710 & w1974;
assign w2040 = (~w2039 & ~w1715) | (~w2039 & w5531) | (~w1715 & w5531);
assign w2041 = ~w2038 & w2040;
assign w2042 = ~w1710 & w1976;
assign w2043 = (~w2042 & ~w1715) | (~w2042 & w5532) | (~w1715 & w5532);
assign w2044 = w1963 & ~w1997;
assign w2045 = ~w1710 & ~w1959;
assign w2046 = (w565 & w1710) | (w565 & w5965) | (w1710 & w5965);
assign w2047 = (w2046 & w1997) | (w2046 & w5533) | (w1997 & w5533);
assign w2048 = w2043 & w2047;
assign w2049 = w2041 & w2048;
assign w2050 = ~w2037 & w2049;
assign w2051 = ~w2001 & ~w2050;
assign w2052 = w2034 & ~w2051;
assign w2053 = (w2000 & ~w2033) | (w2000 & w5534) | (~w2033 & w5534);
assign w2054 = ~w2052 & ~w2053;
assign w2055 = ~w2023 & w2054;
assign w2056 = w2023 & ~w2054;
assign w2057 = ~w2055 & ~w2056;
assign w2058 = ~w1845 & ~w1891;
assign w2059 = w383 & w1022;
assign w2060 = ~w383 & ~w1022;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = w960 & w2061;
assign w2063 = ~w1604 & ~w1854;
assign w2064 = ~w1109 & ~w2063;
assign w2065 = ~w2062 & ~w2064;
assign w2066 = w431 & w5966;
assign w2067 = (w511 & ~w431) | (w511 & w5967) | (~w431 & w5967);
assign w2068 = ~w2066 & ~w2067;
assign w2069 = w386 & w2068;
assign w2070 = (~w1870 & ~w383) | (~w1870 & w5968) | (~w383 & w5968);
assign w2071 = ~w580 & ~w2070;
assign w2072 = ~w2069 & ~w2071;
assign w2073 = w2065 & w2072;
assign w2074 = ~w2065 & ~w2072;
assign w2075 = ~w2073 & ~w2074;
assign w2076 = ~w920 & w1876;
assign w2077 = ~w735 & w1063;
assign w2078 = w735 & ~w1063;
assign w2079 = ~w2077 & ~w2078;
assign w2080 = w920 & ~w2079;
assign w2081 = w432 & w5969;
assign w2082 = ~w2076 & ~w2081;
assign w2083 = ~w2080 & w2082;
assign w2084 = w2075 & ~w2083;
assign w2085 = ~w2075 & w2083;
assign w2086 = ~w2084 & ~w2085;
assign w2087 = ~w1865 & ~w1887;
assign w2088 = (~w2086 & w2087) | (~w2086 & w5535) | (w2087 & w5535);
assign w2089 = ~w2087 & w5536;
assign w2090 = ~w2088 & ~w2089;
assign w2091 = ~w1852 & ~w1860;
assign w2092 = ~w1851 & ~w2091;
assign w2093 = ~w1867 & ~w1882;
assign w2094 = ~w1883 & ~w2093;
assign w2095 = ~w2092 & ~w2094;
assign w2096 = w2092 & w2094;
assign w2097 = ~w2095 & ~w2096;
assign w2098 = (w1633 & w784) | (w1633 & w5537) | (w784 & w5537);
assign w2099 = ~w838 & ~w1633;
assign w2100 = ~w784 & w2099;
assign w2101 = ~w2098 & ~w2100;
assign w2102 = ~w1732 & w2101;
assign w2103 = w1732 & ~w2101;
assign w2104 = ~w2102 & ~w2103;
assign w2105 = ~w2097 & w2104;
assign w2106 = w2097 & ~w2104;
assign w2107 = ~w2105 & ~w2106;
assign w2108 = w2090 & w2107;
assign w2109 = ~w2090 & ~w2107;
assign w2110 = ~w2108 & ~w2109;
assign w2111 = w2058 & w2110;
assign w2112 = ~w1896 & ~w2111;
assign w2113 = ~w1830 & w2112;
assign w2114 = w1722 & w2113;
assign w2115 = ~w1827 & w2114;
assign w2116 = ~w1831 & ~w1931;
assign w2117 = w2112 & ~w2116;
assign w2118 = ~w2058 & ~w2110;
assign w2119 = (~w2118 & w2116) | (~w2118 & w5970) | (w2116 & w5970);
assign w2120 = w1732 & ~w2100;
assign w2121 = ~w2098 & ~w2120;
assign w2122 = w432 & w5971;
assign w2123 = ~w565 & w1063;
assign w2124 = w565 & ~w1063;
assign w2125 = ~w2123 & ~w2124;
assign w2126 = w920 & ~w2125;
assign w2127 = ~w920 & w2077;
assign w2128 = ~w2126 & w5538;
assign w2129 = ~w2121 & w2128;
assign w2130 = w2121 & ~w2128;
assign w2131 = ~w2129 & ~w2130;
assign w2132 = ~w2073 & w2131;
assign w2133 = ~w2084 & w2132;
assign w2134 = (~w2073 & ~w2075) | (~w2073 & w5972) | (~w2075 & w5972);
assign w2135 = ~w2131 & ~w2134;
assign w2136 = ~w2133 & ~w2135;
assign w2137 = ~w960 & ~w2061;
assign w2138 = ~w1150 & ~w2137;
assign w2139 = ~w1877 & w2138;
assign w2140 = w1877 & ~w2138;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = w431 & w5973;
assign w2143 = (w880 & ~w431) | (w880 & w5974) | (~w431 & w5974);
assign w2144 = ~w2142 & ~w2143;
assign w2145 = w386 & w2144;
assign w2146 = ~w386 & w2068;
assign w2147 = ~w1765 & w2146;
assign w2148 = ~w2145 & ~w2147;
assign w2149 = w2141 & ~w2148;
assign w2150 = ~w2141 & w2148;
assign w2151 = ~w2149 & ~w2150;
assign w2152 = ~w2095 & w2104;
assign w2153 = (~w2151 & w2152) | (~w2151 & w5539) | (w2152 & w5539);
assign w2154 = ~w2152 & w5540;
assign w2155 = ~w2153 & ~w2154;
assign w2156 = w2136 & ~w2155;
assign w2157 = ~w2136 & w2155;
assign w2158 = ~w2156 & ~w2157;
assign w2159 = ~w2088 & ~w2107;
assign w2160 = ~w2089 & ~w2159;
assign w2161 = ~w2158 & w2160;
assign w2162 = w2158 & ~w2160;
assign w2163 = ~w2161 & ~w2162;
assign w2164 = ~w227 & ~w409;
assign w2165 = ~w218 & w278;
assign w2166 = ~w180 & ~w226;
assign w2167 = w936 & w2166;
assign w2168 = ~w769 & w1040;
assign w2169 = w2164 & w2168;
assign w2170 = w2165 & w2167;
assign w2171 = w2169 & w2170;
assign w2172 = w675 & w2171;
assign w2173 = ~w124 & ~w457;
assign w2174 = ~w271 & ~w615;
assign w2175 = ~w153 & ~w315;
assign w2176 = ~w178 & ~w321;
assign w2177 = w2173 & w2176;
assign w2178 = w2174 & w2175;
assign w2179 = w2177 & w2178;
assign w2180 = ~w164 & ~w183;
assign w2181 = w705 & w5975;
assign w2182 = ~w211 & ~w296;
assign w2183 = ~w155 & ~w347;
assign w2184 = ~w270 & w2182;
assign w2185 = w2183 & w2184;
assign w2186 = ~w147 & ~w160;
assign w2187 = ~w365 & ~w654;
assign w2188 = w2186 & w2187;
assign w2189 = w232 & w485;
assign w2190 = w2188 & w2189;
assign w2191 = w2179 & w2190;
assign w2192 = w2185 & w2191;
assign w2193 = w2172 & w2192;
assign w2194 = w2181 & w2193;
assign w2195 = ~w2163 & w2194;
assign w2196 = w2163 & ~w2194;
assign w2197 = ~w2195 & ~w2196;
assign w2198 = w2119 & ~w2197;
assign w2199 = ~w2115 & w2198;
assign w2200 = w1722 & w5541;
assign w2201 = ~w1827 & w2200;
assign w2202 = ~w2119 & w2197;
assign w2203 = ~w2201 & ~w2202;
assign w2204 = ~w2199 & w2203;
assign w2205 = (~w1896 & w1831) | (~w1896 & w5542) | (w1831 & w5542);
assign w2206 = (~w2205 & ~w1722) | (~w2205 & w5543) | (~w1722 & w5543);
assign w2207 = w1826 & ~w2205;
assign w2208 = w1825 & w2207;
assign w2209 = ~w2111 & ~w2118;
assign w2210 = ~w2208 & w5544;
assign w2211 = (w2209 & w2208) | (w2209 & w5545) | (w2208 & w5545);
assign w2212 = ~w2210 & ~w2211;
assign w2213 = ~w133 & ~w271;
assign w2214 = w216 & w2213;
assign w2215 = w530 & w791;
assign w2216 = w792 & w2183;
assign w2217 = w2215 & w2216;
assign w2218 = w162 & w2214;
assign w2219 = w750 & w1037;
assign w2220 = w2218 & w2219;
assign w2221 = w663 & w2217;
assign w2222 = w748 & w1669;
assign w2223 = w2221 & w2222;
assign w2224 = w745 & w2220;
assign w2225 = w1524 & w2224;
assign w2226 = w2223 & w2225;
assign w2227 = w2212 & w2226;
assign w2228 = w1949 & ~w2227;
assign w2229 = (w2228 & w1841) | (w2228 & w6587) | (w1841 & w6587);
assign w2230 = ~w2209 & w2226;
assign w2231 = w2209 & ~w2226;
assign w2232 = ~w2230 & ~w2231;
assign w2233 = ~w2208 & w5546;
assign w2234 = (~w2232 & w2208) | (~w2232 & w5547) | (w2208 & w5547);
assign w2235 = ~w2233 & ~w2234;
assign w2236 = w1942 & w2235;
assign w2237 = ~w2227 & ~w2236;
assign w2238 = (~w2237 & w1842) | (~w2237 & w5697) | (w1842 & w5697);
assign w2239 = (w2204 & w2229) | (w2204 & w5548) | (w2229 & w5548);
assign w2240 = ~w2229 & w5549;
assign w2241 = ~w2239 & ~w2240;
assign w2242 = ~w1942 & ~w2235;
assign w2243 = ~w2236 & ~w2242;
assign w2244 = (w2243 & w1842) | (w2243 & w5550) | (w1842 & w5550);
assign w2245 = w2235 & w1949;
assign w2246 = (w2245 & w1841) | (w2245 & w5976) | (w1841 & w5976);
assign w2247 = ~w2244 & ~w2246;
assign w2248 = ~w2241 & ~w2247;
assign w2249 = ~w2194 & ~w2204;
assign w2250 = ~w958 & w5977;
assign w2251 = (w1877 & w958) | (w1877 & w5978) | (w958 & w5978);
assign w2252 = ~w2250 & ~w2251;
assign w2253 = w2078 & w2252;
assign w2254 = ~w2078 & ~w2252;
assign w2255 = ~w2253 & ~w2254;
assign w2256 = ~w2133 & w5551;
assign w2257 = (w2255 & w2133) | (w2255 & w5552) | (w2133 & w5552);
assign w2258 = ~w2256 & ~w2257;
assign w2259 = (~w2139 & ~w2141) | (~w2139 & w5979) | (~w2141 & w5979);
assign w2260 = w432 & w5980;
assign w2261 = ~w511 & w1063;
assign w2262 = w511 & ~w1063;
assign w2263 = ~w2261 & ~w2262;
assign w2264 = ~w920 & w2123;
assign w2265 = (~w2260 & w2263) | (~w2260 & w5981) | (w2263 & w5981);
assign w2266 = ~w2264 & w2265;
assign w2267 = w1856 & w2144;
assign w2268 = ~w386 & ~w2267;
assign w2269 = (w1022 & ~w431) | (w1022 & w5982) | (~w431 & w5982);
assign w2270 = w431 & w5983;
assign w2271 = ~w2269 & ~w2270;
assign w2272 = w386 & w2271;
assign w2273 = ~w2268 & w5984;
assign w2274 = (~w2266 & w2268) | (~w2266 & w5985) | (w2268 & w5985);
assign w2275 = ~w2273 & ~w2274;
assign w2276 = ~w2259 & w2275;
assign w2277 = w2259 & ~w2275;
assign w2278 = ~w2276 & ~w2277;
assign w2279 = w2258 & w2278;
assign w2280 = ~w2258 & ~w2278;
assign w2281 = ~w2279 & ~w2280;
assign w2282 = ~w2136 & ~w2154;
assign w2283 = ~w2153 & ~w2282;
assign w2284 = w2281 & w2283;
assign w2285 = ~w2281 & ~w2283;
assign w2286 = ~w2284 & ~w2285;
assign w2287 = w2161 & w2286;
assign w2288 = ~w2118 & ~w2162;
assign w2289 = ~w2118 & w5986;
assign w2290 = w2162 & ~w2286;
assign w2291 = ~w337 & ~w615;
assign w2292 = w664 & w937;
assign w2293 = w2291 & w2292;
assign w2294 = w2167 & w2293;
assign w2295 = ~w141 & ~w231;
assign w2296 = ~w241 & w2295;
assign w2297 = ~w468 & ~w935;
assign w2298 = ~w89 & ~w315;
assign w2299 = ~w235 & ~w538;
assign w2300 = w156 & w2298;
assign w2301 = w2299 & w2300;
assign w2302 = ~w58 & ~w230;
assign w2303 = ~w456 & w2302;
assign w2304 = w259 & w483;
assign w2305 = w2297 & w2304;
assign w2306 = w293 & w2303;
assign w2307 = w1559 & w2296;
assign w2308 = w2306 & w2307;
assign w2309 = w2301 & w2305;
assign w2310 = w2308 & w2309;
assign w2311 = ~w158 & ~w181;
assign w2312 = ~w336 & w2311;
assign w2313 = w2310 & w2312;
assign w2314 = ~w130 & w149;
assign w2315 = ~w189 & ~w238;
assign w2316 = ~w265 & w2315;
assign w2317 = ~w150 & ~w166;
assign w2318 = ~w279 & ~w362;
assign w2319 = w2317 & w2318;
assign w2320 = w610 & w2319;
assign w2321 = w1041 & w2316;
assign w2322 = w2320 & w2321;
assign w2323 = ~w205 & ~w218;
assign w2324 = ~w303 & ~w2314;
assign w2325 = w2323 & w2324;
assign w2326 = w459 & w810;
assign w2327 = w1026 & w1665;
assign w2328 = w2326 & w2327;
assign w2329 = w933 & w2325;
assign w2330 = w2328 & w2329;
assign w2331 = w2294 & w2330;
assign w2332 = w2322 & w2331;
assign w2333 = w2313 & w2332;
assign w2334 = ~w2290 & w2333;
assign w2335 = (w2117 & w5987) | (w2117 & w5988) | (w5987 & w5988);
assign w2336 = ~w1830 & ~w2287;
assign w2337 = w2112 & w2336;
assign w2338 = w1722 & w2337;
assign w2339 = w2337 & w5989;
assign w2340 = ~w1827 & w2339;
assign w2341 = ~w2335 & ~w2340;
assign w2342 = ~w2161 & ~w2286;
assign w2343 = ~w2119 & w2342;
assign w2344 = w1722 & w5554;
assign w2345 = ~w1827 & w2344;
assign w2346 = ~w2343 & ~w2345;
assign w2347 = ~w2341 & w2346;
assign w2348 = (w2288 & w2116) | (w2288 & w5698) | (w2116 & w5698);
assign w2349 = (w2348 & w1827) | (w2348 & w5555) | (w1827 & w5555);
assign w2350 = ~w2333 & w2342;
assign w2351 = ~w2349 & w2350;
assign w2352 = ~w1827 & w2338;
assign w2353 = ~w2333 & w7748;
assign w2354 = ~w2352 & w2353;
assign w2355 = ~w2351 & ~w2354;
assign w2356 = ~w2347 & w2355;
assign w2357 = w2249 & ~w2356;
assign w2358 = ~w2249 & w2355;
assign w2359 = ~w2249 & w2356;
assign w2360 = ~w2357 & ~w2359;
assign w2361 = ~w2238 & ~w2360;
assign w2362 = w2194 & ~w2204;
assign w2363 = ~w2356 & ~w2362;
assign w2364 = w2356 & w2362;
assign w2365 = ~w2363 & ~w2364;
assign w2366 = w2238 & w2365;
assign w2367 = ~w2361 & ~w2366;
assign w2368 = ~w2248 & w2367;
assign w2369 = w1948 & ~w2235;
assign w2370 = ~w1948 & w2235;
assign w2371 = ~w2369 & ~w2370;
assign w2372 = w1842 & ~w2371;
assign w2373 = ~w1842 & ~w2243;
assign w2374 = ~w2372 & ~w2373;
assign w2375 = ~w1953 & w2374;
assign w2376 = ~w1956 & w2375;
assign w2377 = w1952 & ~w2243;
assign w2378 = ~w2212 & ~w2226;
assign w2379 = ~w2204 & ~w2378;
assign w2380 = w2204 & w2378;
assign w2381 = ~w2379 & ~w2380;
assign w2382 = ~w2244 & w5990;
assign w2383 = ~w2377 & ~w2382;
assign w2384 = (w2383 & w1956) | (w2383 & w5556) | (w1956 & w5556);
assign w2385 = w2368 & ~w2384;
assign w2386 = w2248 & ~w2367;
assign w2387 = ~w2367 & w2383;
assign w2388 = ~w2376 & w2387;
assign w2389 = (~w2386 & w2376) | (~w2386 & w5557) | (w2376 & w5557);
assign w2390 = ~w2385 & w2389;
assign w2391 = ~w726 & ~w854;
assign w2392 = w847 & w871;
assign w2393 = ~w2392 & w7376;
assign w2394 = w2391 & ~w2393;
assign w2395 = w726 & w854;
assign w2396 = ~w2393 & w2395;
assign w2397 = (w726 & w2393) | (w726 & w6605) | (w2393 & w6605);
assign w2398 = ~w2394 & ~w2397;
assign w2399 = w847 & ~w854;
assign w2400 = ~w847 & w854;
assign w2401 = ~w2399 & ~w2400;
assign w2402 = w2393 & w2401;
assign w2403 = ~w2391 & ~w2395;
assign w2404 = w2393 & ~w2401;
assign w2405 = ~w2403 & w2404;
assign w2406 = ~w2244 & w5991;
assign w2407 = w2359 & ~w2239;
assign w2408 = (w2204 & w2236) | (w2204 & w6606) | (w2236 & w6606);
assign w2409 = (w2363 & w2229) | (w2363 & w5699) | (w2229 & w5699);
assign w2410 = ~w2407 & ~w2409;
assign w2411 = ~w2393 & w2403;
assign w2412 = (~w2406 & ~w2241) | (~w2406 & w5992) | (~w2241 & w5992);
assign w2413 = w2412 & w6607;
assign w2414 = (w726 & ~w2412) | (w726 & w6608) | (~w2412 & w6608);
assign w2415 = w2412 & w6609;
assign w2416 = (w2415 & ~w2389) | (w2415 & w5993) | (~w2389 & w5993);
assign w2417 = (~w2414 & ~w2390) | (~w2414 & w5700) | (~w2390 & w5700);
assign w2418 = ~w2416 & w2417;
assign w2419 = w2057 & w2418;
assign w2420 = w1952 & w2405;
assign w2421 = ~w2244 & w5994;
assign w2422 = ~w2420 & ~w2421;
assign w2423 = ~w2229 & w5558;
assign w2424 = ~w2204 & w2411;
assign w2425 = (w2424 & w2229) | (w2424 & w5559) | (w2229 & w5559);
assign w2426 = ~w2423 & ~w2425;
assign w2427 = w726 & w2426;
assign w2428 = w2422 & w2427;
assign w2429 = (~w2377 & w1956) | (~w2377 & w5560) | (w1956 & w5560);
assign w2430 = (~w2382 & w2241) | (~w2382 & w5995) | (w2241 & w5995);
assign w2431 = w2429 & ~w2430;
assign w2432 = w2429 & w5701;
assign w2433 = w2428 & w2430;
assign w2434 = ~w2429 & w2433;
assign w2435 = (~w726 & ~w2422) | (~w726 & w5702) | (~w2422 & w5702);
assign w2436 = ~w2393 & ~w2403;
assign w2437 = w2427 & w5996;
assign w2438 = ~w2435 & ~w2437;
assign w2439 = ~w2434 & w2438;
assign w2440 = ~w2432 & w2439;
assign w2441 = ~w2248 & w5703;
assign w2442 = w2429 & w2441;
assign w2443 = (w2394 & w2248) | (w2394 & w5704) | (w2248 & w5704);
assign w2444 = ~w2429 & w2443;
assign w2445 = ~w2442 & ~w2444;
assign w2446 = (w565 & w1710) | (w565 & w5997) | (w1710 & w5997);
assign w2447 = ~w2000 & ~w2446;
assign w2448 = ~w2050 & ~w2447;
assign w2449 = w2043 & ~w2044;
assign w2450 = ~w6000 & w2449;
assign w2451 = w2449 & w5998;
assign w2452 = ~w2037 & w5999;
assign w2453 = ~w2448 & ~w2452;
assign w2454 = ~w2034 & w2453;
assign w2455 = w2034 & ~w2453;
assign w2456 = ~w2454 & ~w2455;
assign w2457 = (~w2456 & ~w2440) | (~w2456 & w5705) | (~w2440 & w5705);
assign w2458 = w1953 & ~w2374;
assign w2459 = ~w2375 & ~w2458;
assign w2460 = ~w1956 & w2459;
assign w2461 = w1955 & w5561;
assign w2462 = ~w2460 & ~w2461;
assign w2463 = (w2394 & w2460) | (w2394 & w5562) | (w2460 & w5562);
assign w2464 = (w565 & ~w2449) | (w565 & w6000) | (~w2449 & w6000);
assign w2465 = (w2464 & w2037) | (w2464 & w6001) | (w2037 & w6001);
assign w2466 = ~w2037 & w6002;
assign w2467 = ~w2465 & ~w2466;
assign w2468 = w2463 & w2467;
assign w2469 = (w2396 & w2460) | (w2396 & w5563) | (w2460 & w5563);
assign w2470 = ~w1823 & w6003;
assign w2471 = (~w2470 & ~w1952) | (~w2470 & w6004) | (~w1952 & w6004);
assign w2472 = w2471 & w5564;
assign w2473 = (w726 & ~w2471) | (w726 & w5565) | (~w2471 & w5565);
assign w2474 = ~w2472 & ~w2473;
assign w2475 = w2467 & w2474;
assign w2476 = ~w2469 & w2475;
assign w2477 = ~w2468 & ~w2476;
assign w2478 = ~w2036 & w2436;
assign w2479 = ~w1710 & w2405;
assign w2480 = w1704 & w2411;
assign w2481 = (~w2479 & ~w1715) | (~w2479 & w6005) | (~w1715 & w6005);
assign w2482 = ~w2480 & w2481;
assign w2483 = ~w1710 & w2392;
assign w2484 = w6555 & ~w2483;
assign w2485 = ~w1710 & w2402;
assign w2486 = w1715 & w2411;
assign w2487 = (~w2485 & w1997) | (~w2485 & w5566) | (w1997 & w5566);
assign w2488 = ~w2486 & w2487;
assign w2489 = ~w6620 & w2488;
assign w2490 = (w2478 & w6588) | (w2478 & w6589) | (w6588 & w6589);
assign w2491 = ~w1818 & w2436;
assign w2492 = w1716 & w2491;
assign w2493 = ~w1823 & w5568;
assign w2494 = w1704 & w2402;
assign w2495 = w1715 & w2405;
assign w2496 = ~w2494 & ~w2495;
assign w2497 = ~w2493 & w2496;
assign w2498 = ~w2492 & w2497;
assign w2499 = w2498 & w5569;
assign w2500 = ~w2490 & w2499;
assign w2501 = ~w2478 & w6590;
assign w2502 = ~w1710 & w1957;
assign w2503 = (w2502 & ~w2498) | (w2502 & w5571) | (~w2498 & w5571);
assign w2504 = ~w2501 & ~w2503;
assign w2505 = ~w2500 & w2504;
assign w2506 = w6000 & ~w2449;
assign w2507 = ~w2450 & ~w2506;
assign w2508 = ~w2505 & w2507;
assign w2509 = w2505 & ~w2507;
assign w2510 = ~w1816 & w6006;
assign w2511 = ~w1819 & w2510;
assign w2512 = ~w1955 & w2511;
assign w2513 = ~w1823 & w6007;
assign w2514 = w1704 & w2405;
assign w2515 = w1952 & w2411;
assign w2516 = ~w2513 & ~w2514;
assign w2517 = ~w2515 & w2516;
assign w2518 = ~w2512 & w2517;
assign w2519 = w2518 & w5572;
assign w2520 = (w726 & ~w2518) | (w726 & w5573) | (~w2518 & w5573);
assign w2521 = ~w2519 & ~w2520;
assign w2522 = ~w2509 & w2521;
assign w2523 = ~w2508 & ~w2522;
assign w2524 = w2477 & w2523;
assign w2525 = w2445 & w2456;
assign w2526 = w2440 & w2525;
assign w2527 = ~w2469 & w2474;
assign w2528 = ~w2463 & ~w2467;
assign w2529 = ~w2527 & w2528;
assign w2530 = (~w2529 & ~w2440) | (~w2529 & w6008) | (~w2440 & w6008);
assign w2531 = ~w2524 & w2530;
assign w2532 = ~w2457 & ~w2531;
assign w2533 = ~w2057 & ~w2418;
assign w2534 = ~w2419 & ~w2533;
assign w2535 = ~w2532 & w2534;
assign w2536 = ~w2419 & ~w2535;
assign w2537 = ~w2021 & ~w2054;
assign w2538 = ~w2013 & w2537;
assign w2539 = w2011 & ~w2538;
assign w2540 = (w2002 & w1997) | (w2002 & w5574) | (w1997 & w5574);
assign w2541 = w1993 & w2540;
assign w2542 = (~w1022 & ~w2540) | (~w1022 & w6009) | (~w2540 & w6009);
assign w2543 = w1994 & ~w2036;
assign w2544 = w1704 & w1987;
assign w2545 = w1983 & ~w1986;
assign w2546 = ~w1990 & w2545;
assign w2547 = ~w1710 & w2546;
assign w2548 = (~w2547 & ~w1715) | (~w2547 & w5575) | (~w1715 & w5575);
assign w2549 = ~w2544 & w2548;
assign w2550 = (w2542 & w2543) | (w2542 & w5576) | (w2543 & w5576);
assign w2551 = ~w2543 & w5577;
assign w2552 = ~w2550 & ~w2551;
assign w2553 = (w1968 & w1842) | (w1968 & w5578) | (w1842 & w5578);
assign w2554 = ~w2244 & w2553;
assign w2555 = ~w1823 & w5579;
assign w2556 = ~w1948 & w5580;
assign w2557 = ~w1841 & w6010;
assign w2558 = (w1976 & w1948) | (w1976 & w5581) | (w1948 & w5581);
assign w2559 = (~w2558 & w1841) | (~w2558 & w6011) | (w1841 & w6011);
assign w2560 = ~w2557 & ~w2559;
assign w2561 = ~w2555 & ~w2560;
assign w2562 = (w565 & ~w2561) | (w565 & w5582) | (~w2561 & w5582);
assign w2563 = ~w1959 & w1960;
assign w2564 = ~w2563 & ~w6968;
assign w2565 = w2561 & w5583;
assign w2566 = ~w2562 & ~w2565;
assign w2567 = w2552 & ~w2566;
assign w2568 = ~w2552 & w2566;
assign w2569 = ~w2567 & ~w2568;
assign w2570 = ~w2462 & ~w2569;
assign w2571 = w2561 & w5584;
assign w2572 = ~w2562 & ~w2571;
assign w2573 = ~w2552 & ~w2572;
assign w2574 = w2552 & w2572;
assign w2575 = w2462 & w5585;
assign w2576 = ~w2570 & ~w2575;
assign w2577 = w2539 & w2576;
assign w2578 = ~w2539 & ~w2576;
assign w2579 = ~w2577 & ~w2578;
assign w2580 = w2241 & ~w2360;
assign w2581 = ~w2368 & ~w2580;
assign w2582 = w2383 & ~w2580;
assign w2583 = ~w2376 & w2582;
assign w2584 = ~w2581 & ~w2583;
assign w2585 = (~w2284 & w1654) | (~w2284 & w5586) | (w1654 & w5586);
assign w2586 = ~w1721 & w2585;
assign w2587 = w2337 & w2586;
assign w2588 = ~w1827 & w2587;
assign w2589 = ~w2284 & ~w2287;
assign w2590 = (~w2257 & ~w2258) | (~w2257 & w6012) | (~w2258 & w6012);
assign w2591 = w385 & w2270;
assign w2592 = ~w433 & ~w2591;
assign w2593 = (w2124 & w2592) | (w2124 & w6013) | (w2592 & w6013);
assign w2594 = ~w2592 & w6014;
assign w2595 = ~w2593 & ~w2594;
assign w2596 = ~w920 & w2261;
assign w2597 = w880 & ~w1063;
assign w2598 = ~w880 & w1063;
assign w2599 = ~w2597 & ~w2598;
assign w2600 = w920 & ~w2599;
assign w2601 = w432 & w6015;
assign w2602 = ~w2596 & ~w2601;
assign w2603 = ~w2600 & w2602;
assign w2604 = w2595 & w2603;
assign w2605 = ~w2595 & ~w2603;
assign w2606 = ~w2604 & ~w2605;
assign w2607 = (~w2251 & ~w2252) | (~w2251 & w6016) | (~w2252 & w6016);
assign w2608 = (~w2273 & w2259) | (~w2273 & w6017) | (w2259 & w6017);
assign w2609 = ~w2607 & ~w2608;
assign w2610 = w2607 & w2608;
assign w2611 = ~w2609 & ~w2610;
assign w2612 = w2606 & w2611;
assign w2613 = ~w2606 & ~w2611;
assign w2614 = ~w2612 & ~w2613;
assign w2615 = w2590 & ~w2614;
assign w2616 = ~w2590 & w2614;
assign w2617 = ~w2615 & ~w2616;
assign w2618 = ~w179 & w349;
assign w2619 = ~w109 & ~w249;
assign w2620 = ~w346 & ~w769;
assign w2621 = ~w234 & ~w402;
assign w2622 = w2620 & w2621;
assign w2623 = w682 & w2622;
assign w2624 = ~w437 & ~w588;
assign w2625 = w2173 & w2624;
assign w2626 = w202 & w2625;
assign w2627 = w301 & w2623;
assign w2628 = w2626 & w2627;
assign w2629 = w278 & ~w477;
assign w2630 = w415 & w1547;
assign w2631 = w2619 & w2630;
assign w2632 = w2316 & w2629;
assign w2633 = w2618 & w2632;
assign w2634 = w312 & w2631;
assign w2635 = w2633 & w2634;
assign w2636 = w2310 & w2635;
assign w2637 = w2628 & w2636;
assign w2638 = ~w2617 & w2637;
assign w2639 = w2617 & ~w2637;
assign w2640 = ~w2638 & ~w2639;
assign w2641 = w2640 & w7749;
assign w2642 = ~w2588 & w2641;
assign w2643 = w2337 & w6018;
assign w2644 = ~w1827 & w2643;
assign w2645 = (w2117 & w6019) | (w2117 & w6020) | (w6019 & w6020);
assign w2646 = ~w2644 & ~w2645;
assign w2647 = ~w2642 & w2646;
assign w2648 = (~w2347 & w2249) | (~w2347 & w5588) | (w2249 & w5588);
assign w2649 = ~w2647 & ~w2648;
assign w2650 = w2204 & ~w2347;
assign w2651 = (~w2229 & w6021) | (~w2229 & w6022) | (w6021 & w6022);
assign w2652 = w2647 & w2648;
assign w2653 = w2647 & w2650;
assign w2654 = (~w2229 & w6023) | (~w2229 & w6024) | (w6023 & w6024);
assign w2655 = ~w2651 & w2654;
assign w2656 = w2410 & w2655;
assign w2657 = ~w2355 & ~w2647;
assign w2658 = w2355 & w2647;
assign w2659 = ~w2657 & ~w2658;
assign w2660 = ~w2410 & w2659;
assign w2661 = ~w2656 & ~w2660;
assign w2662 = (w2661 & w2583) | (w2661 & w5591) | (w2583 & w5591);
assign w2663 = ~w2583 & w5592;
assign w2664 = ~w2662 & ~w2663;
assign w2665 = w2411 & ~w2655;
assign w2666 = w2241 & w2405;
assign w2667 = ~w2665 & w7278;
assign w2668 = (w2665 & w726) | (w2665 & w7279) | (w726 & w7279);
assign w2669 = ~w2665 & w7280;
assign w2670 = w2664 & w2669;
assign w2671 = (~w2668 & w2664) | (~w2668 & w5706) | (w2664 & w5706);
assign w2672 = ~w2670 & w2671;
assign w2673 = ~w2579 & ~w2672;
assign w2674 = w2579 & w2672;
assign w2675 = ~w2673 & ~w2674;
assign w2676 = (~w2609 & ~w2611) | (~w2609 & w6028) | (~w2611 & w6028);
assign w2677 = (~w2594 & ~w2595) | (~w2594 & w6029) | (~w2595 & w6029);
assign w2678 = w1022 & w1063;
assign w2679 = ~w1022 & ~w1063;
assign w2680 = ~w2678 & ~w2679;
assign w2681 = w920 & ~w2680;
assign w2682 = ~w920 & w2598;
assign w2683 = w432 & w6030;
assign w2684 = ~w2681 & w6031;
assign w2685 = w2677 & ~w2684;
assign w2686 = ~w2677 & w2684;
assign w2687 = ~w2685 & ~w2686;
assign w2688 = (~w2124 & w385) | (~w2124 & w6032) | (w385 & w6032);
assign w2689 = w2262 & ~w2688;
assign w2690 = ~w2262 & w2688;
assign w2691 = ~w2689 & ~w2690;
assign w2692 = w2687 & ~w2691;
assign w2693 = ~w2687 & w2691;
assign w2694 = ~w2692 & ~w2693;
assign w2695 = ~w2676 & w2694;
assign w2696 = w2676 & ~w2694;
assign w2697 = ~w2695 & ~w2696;
assign w2698 = ~w314 & ~w484;
assign w2699 = w107 & w259;
assign w2700 = w353 & w403;
assign w2701 = w425 & w466;
assign w2702 = w2698 & w2701;
assign w2703 = w2699 & w2700;
assign w2704 = w693 & w790;
assign w2705 = w2703 & w2704;
assign w2706 = w2702 & w2705;
assign w2707 = w195 & w775;
assign w2708 = w2706 & w2707;
assign w2709 = w455 & w2708;
assign w2710 = ~w2697 & ~w2709;
assign w2711 = ~w2284 & ~w2616;
assign w2712 = ~w2615 & ~w2711;
assign w2713 = w2710 & ~w2712;
assign w2714 = (w2713 & w2352) | (w2713 & w5593) | (w2352 & w5593);
assign w2715 = w2337 & w6033;
assign w2716 = ~w1827 & w2715;
assign w2717 = (w2117 & w5707) | (w2117 & w5708) | (w5707 & w5708);
assign w2718 = (~w2709 & w2614) | (~w2709 & w6034) | (w2614 & w6034);
assign w2719 = w2697 & w2718;
assign w2720 = ~w2716 & w5594;
assign w2721 = ~w2714 & ~w2720;
assign w2722 = ~w2695 & w2711;
assign w2723 = w2337 & w6035;
assign w2724 = ~w1827 & w2723;
assign w2725 = (~w2695 & w2615) | (~w2695 & w6036) | (w2615 & w6036);
assign w2726 = ~w2124 & ~w2262;
assign w2727 = w917 & w2270;
assign w2728 = w2597 & w2727;
assign w2729 = w919 & w1063;
assign w2730 = ~w2597 & ~w2678;
assign w2731 = w2730 & w6037;
assign w2732 = (w2726 & w2731) | (w2726 & w6038) | (w2731 & w6038);
assign w2733 = ~w2731 & w6039;
assign w2734 = ~w2732 & ~w2733;
assign w2735 = (w2687 & w7281) | (w2687 & w7282) | (w7281 & w7282);
assign w2736 = (w6040 & ~w2687) | (w6040 & w7283) | (~w2687 & w7283);
assign w2737 = ~w2735 & ~w2736;
assign w2738 = ~w264 & ~w477;
assign w2739 = ~w470 & ~w627;
assign w2740 = ~w291 & ~w465;
assign w2741 = ~w141 & ~w164;
assign w2742 = ~w213 & ~w234;
assign w2743 = w2741 & w2742;
assign w2744 = ~w366 & ~w373;
assign w2745 = ~w456 & ~w678;
assign w2746 = w2744 & w2745;
assign w2747 = w622 & w788;
assign w2748 = w2740 & w2747;
assign w2749 = w2743 & w2746;
assign w2750 = w2748 & w2749;
assign w2751 = ~w236 & w1038;
assign w2752 = ~w181 & ~w270;
assign w2753 = w232 & w2752;
assign w2754 = w345 & w2297;
assign w2755 = w2738 & w2739;
assign w2756 = w2754 & w2755;
assign w2757 = w331 & w2753;
assign w2758 = w2751 & w2757;
assign w2759 = w816 & w2756;
assign w2760 = w2758 & w2759;
assign w2761 = w2294 & w2750;
assign w2762 = w2760 & w2761;
assign w2763 = w1568 & w2762;
assign w2764 = w2737 & w2763;
assign w2765 = ~w2737 & ~w2763;
assign w2766 = ~w2764 & ~w2765;
assign w2767 = ~w2724 & w5709;
assign w2768 = (w2766 & w2724) | (w2766 & w5710) | (w2724 & w5710);
assign w2769 = ~w2767 & ~w2768;
assign w2770 = w2721 & w2769;
assign w2771 = ~w2721 & ~w2769;
assign w2772 = ~w2770 & ~w2771;
assign w2773 = w2655 & ~w2772;
assign w2774 = w2697 & w2709;
assign w2775 = ~w2712 & w2774;
assign w2776 = (w2775 & w2352) | (w2775 & w5596) | (w2352 & w5596);
assign w2777 = (w2709 & w2614) | (w2709 & w6041) | (w2614 & w6041);
assign w2778 = ~w2697 & w2777;
assign w2779 = ~w2716 & w5597;
assign w2780 = ~w2776 & ~w2779;
assign w2781 = w2721 & w2780;
assign w2782 = w2637 & w2647;
assign w2783 = (~w2782 & w2648) | (~w2782 & w5711) | (w2648 & w5711);
assign w2784 = w2650 & ~w2782;
assign w2785 = (w2784 & w2229) | (w2784 & w5598) | (w2229 & w5598);
assign w2786 = ~w2785 & w5712;
assign w2787 = (w2781 & w2785) | (w2781 & w5713) | (w2785 & w5713);
assign w2788 = ~w2786 & ~w2787;
assign w2789 = ~w2773 & w2788;
assign w2790 = ~w2781 & ~w2782;
assign w2791 = w2781 & w2782;
assign w2792 = ~w2790 & ~w2791;
assign w2793 = (w5715 & w6611) | (w5715 & w6612) | (w6611 & w6612);
assign w2794 = ~w2637 & w2647;
assign w2795 = ~w2781 & w2794;
assign w2796 = w2781 & ~w2794;
assign w2797 = ~w2795 & ~w2796;
assign w2798 = w2797 & w7750;
assign w2799 = ~w2793 & ~w2798;
assign w2800 = ~w2656 & ~w2799;
assign w2801 = ~w2789 & ~w2800;
assign w2802 = w2661 & ~w2789;
assign w2803 = (~w2801 & w2584) | (~w2801 & w5599) | (w2584 & w5599);
assign w2804 = ~w2763 & w2769;
assign w2805 = ~w2347 & ~w2647;
assign w2806 = w2780 & w2805;
assign w2807 = w2805 & w5600;
assign w2808 = (w2807 & w2229) | (w2807 & w5601) | (w2229 & w5601);
assign w2809 = (w2780 & w2794) | (w2780 & w5602) | (w2794 & w5602);
assign w2810 = ~w2358 & w2806;
assign w2811 = ~w2810 & w5603;
assign w2812 = ~w2808 & w2811;
assign w2813 = (~w2804 & w2808) | (~w2804 & w6042) | (w2808 & w6042);
assign w2814 = (~w2763 & ~w5709) | (~w2763 & w6043) | (~w5709 & w6043);
assign w2815 = ~w2810 & w5604;
assign w2816 = ~w2725 & w2737;
assign w2817 = ~w517 & ~w528;
assign w2818 = ~w164 & ~w435;
assign w2819 = ~w321 & w2818;
assign w2820 = w2296 & w2819;
assign w2821 = ~w150 & ~w206;
assign w2822 = ~w256 & ~w477;
assign w2823 = ~w609 & w2822;
assign w2824 = w2821 & w2823;
assign w2825 = ~w163 & ~w467;
assign w2826 = w216 & w398;
assign w2827 = w459 & w1506;
assign w2828 = w2817 & w2825;
assign w2829 = w2827 & w2828;
assign w2830 = w2826 & w2829;
assign w2831 = w2820 & w2824;
assign w2832 = w2830 & w2831;
assign w2833 = w493 & w697;
assign w2834 = w2832 & w2833;
assign w2835 = w1922 & w2834;
assign w2836 = w919 & ~w1986;
assign w2837 = ~w919 & w1986;
assign w2838 = ~w1063 & ~w2836;
assign w2839 = ~w2837 & w2838;
assign w2840 = ~w2835 & w2839;
assign w2841 = w2835 & ~w2839;
assign w2842 = ~w2840 & ~w2841;
assign w2843 = (w2687 & w7284) | (w2687 & w7285) | (w7284 & w7285);
assign w2844 = ~w2731 & ~w2733;
assign w2845 = (w6045 & w6046) | (w6045 & ~w2692) | (w6046 & ~w2692);
assign w2846 = ~w2843 & ~w2845;
assign w2847 = w2842 & w2846;
assign w2848 = ~w2842 & ~w2846;
assign w2849 = ~w2847 & ~w2848;
assign w2850 = ~w2724 & w5716;
assign w2851 = (~w2849 & w2724) | (~w2849 & w5717) | (w2724 & w5717);
assign w2852 = ~w2850 & ~w2851;
assign w2853 = ~w2767 & ~w2852;
assign w2854 = (w2853 & w2808) | (w2853 & w6047) | (w2808 & w6047);
assign w2855 = ~w2813 & w2854;
assign w2856 = ~w2808 & w6048;
assign w2857 = ~w2804 & w2852;
assign w2858 = (w2857 & w2808) | (w2857 & w6049) | (w2808 & w6049);
assign w2859 = ~w2856 & ~w2858;
assign w2860 = ~w2855 & w2859;
assign w2861 = ~w2803 & ~w2860;
assign w2862 = (~w2769 & w2810) | (~w2769 & w5606) | (w2810 & w5606);
assign w2863 = ~w2769 & w2807;
assign w2864 = ~w2238 & w2863;
assign w2865 = ~w2862 & ~w2864;
assign w2866 = ~w2812 & w2865;
assign w2867 = ~w2788 & ~w2866;
assign w2868 = ~w2860 & ~w2867;
assign w2869 = ~w2789 & w2860;
assign w2870 = ~w2868 & ~w2869;
assign w2871 = w2800 & w2860;
assign w2872 = ~w2867 & w2871;
assign w2873 = (~w2870 & w2662) | (~w2870 & w6050) | (w2662 & w6050);
assign w2874 = ~w2861 & w2873;
assign w2875 = w574 & ~w871;
assign w2876 = (a_2 & w0) | (a_2 & w6051) | (w0 & w6051);
assign w2877 = ~w0 & w6052;
assign w2878 = ~w2876 & ~w2877;
assign w2879 = w391 & ~w2878;
assign w2880 = ~w391 & w2878;
assign w2881 = ~w2879 & ~w2880;
assign w2882 = w2875 & w2881;
assign w2883 = ~w2874 & w2882;
assign w2884 = ~w574 & w871;
assign w2885 = w2881 & w2884;
assign w2886 = w391 & w574;
assign w2887 = ~w391 & ~w574;
assign w2888 = ~w2886 & ~w2887;
assign w2889 = ~w2875 & ~w2884;
assign w2890 = ~w2881 & w2888;
assign w2891 = ~w2889 & w2890;
assign w2892 = w2788 & w2891;
assign w2893 = ~w2881 & ~w2888;
assign w2894 = w2865 & w6613;
assign w2895 = ~w2769 & ~w2852;
assign w2896 = (w2895 & w2810) | (w2895 & w5607) | (w2810 & w5607);
assign w2897 = w2807 & w2895;
assign w2898 = ~w2238 & w2897;
assign w2899 = ~w2896 & ~w2898;
assign w2900 = w2804 & ~w2852;
assign w2901 = (~w2900 & ~w5608) | (~w2900 & w5718) | (~w5608 & w5718);
assign w2902 = w2899 & w2901;
assign w2903 = w2881 & w2889;
assign w2904 = w2901 & w6053;
assign w2905 = ~w2892 & ~w2894;
assign w2906 = (w871 & ~w2905) | (w871 & w6054) | (~w2905 & w6054);
assign w2907 = w2905 & w6055;
assign w2908 = ~w2906 & ~w2907;
assign w2909 = (w2908 & w2874) | (w2908 & w5719) | (w2874 & w5719);
assign w2910 = ~w2883 & ~w2909;
assign w2911 = w2675 & w2910;
assign w2912 = w2536 & w2911;
assign w2913 = ~w2675 & w2910;
assign w2914 = ~w2536 & w2913;
assign w2915 = ~w2912 & ~w2914;
assign w2916 = w2536 & w2675;
assign w2917 = (~w2910 & w2536) | (~w2910 & w5720) | (w2536 & w5720);
assign w2918 = ~w2916 & w2917;
assign w2919 = w2915 & ~w2918;
assign w2920 = (~w2529 & ~w2523) | (~w2529 & w5721) | (~w2523 & w5721);
assign w2921 = ~w2457 & ~w2526;
assign w2922 = ~w2920 & w2921;
assign w2923 = w2920 & ~w2921;
assign w2924 = ~w2922 & ~w2923;
assign w2925 = w2800 & ~w2662;
assign w2926 = w2656 & w2799;
assign w2927 = ~w2580 & ~w2660;
assign w2928 = w2799 & w2927;
assign w2929 = (~w2926 & w2385) | (~w2926 & w6614) | (w2385 & w6614);
assign w2930 = ~w2925 & w2929;
assign w2931 = ~w2925 & w6615;
assign w2932 = ~w2655 & w2893;
assign w2933 = ~w2410 & w2891;
assign w2934 = ~w2932 & ~w2933;
assign w2935 = (w871 & ~w2934) | (w871 & w6616) | (~w2934 & w6616);
assign w2936 = w2934 & w6617;
assign w2937 = ~w2935 & ~w2936;
assign w2938 = (w2937 & ~w2930) | (w2937 & w6056) | (~w2930 & w6056);
assign w2939 = ~w2931 & ~w2938;
assign w2940 = ~w2924 & w2939;
assign w2941 = ~w2664 & w2882;
assign w2942 = ~w2410 & w2893;
assign w2943 = w2241 & w2891;
assign w2944 = ~w2942 & ~w2943;
assign w2945 = (w871 & ~w2944) | (w871 & w6057) | (~w2944 & w6057);
assign w2946 = w2944 & w6058;
assign w2947 = ~w2945 & ~w2946;
assign w2948 = (w2947 & w2664) | (w2947 & w5722) | (w2664 & w5722);
assign w2949 = ~w2941 & ~w2948;
assign w2950 = w2477 & ~w2529;
assign w2951 = w2523 & ~w2950;
assign w2952 = ~w2523 & w2950;
assign w2953 = ~w2951 & ~w2952;
assign w2954 = ~w2949 & ~w2953;
assign w2955 = ~w2244 & w6059;
assign w2956 = (~w2955 & ~w2241) | (~w2955 & w6060) | (~w2241 & w6060);
assign w2957 = w2956 & w6618;
assign w2958 = (~w2882 & w6062) | (~w2882 & w7867) | (w6062 & w7867);
assign w2959 = w2390 & ~w2958;
assign w2960 = (~w871 & ~w2956) | (~w871 & w6619) | (~w2956 & w6619);
assign w2961 = ~w2960 & w7751;
assign w2962 = ~w2959 & w2961;
assign w2963 = ~w2508 & ~w2509;
assign w2964 = w2521 & w2963;
assign w2965 = ~w2521 & ~w2963;
assign w2966 = ~w2964 & ~w2965;
assign w2967 = ~w2962 & ~w2966;
assign w2968 = ~w2248 & w5723;
assign w2969 = w2429 & w2968;
assign w2970 = (w2882 & w2248) | (w2882 & w5724) | (w2248 & w5724);
assign w2971 = ~w2429 & w2970;
assign w2972 = ~w2969 & ~w2971;
assign w2973 = ~w2248 & w5725;
assign w2974 = w2429 & w2973;
assign w2975 = w2241 & w2903;
assign w2976 = w1952 & w2891;
assign w2977 = ~w2244 & w6064;
assign w2978 = ~w2976 & ~w2977;
assign w2979 = ~w2975 & w6065;
assign w2980 = (~w871 & w2975) | (~w871 & w6066) | (w2975 & w6066);
assign w2981 = ~w2979 & ~w2980;
assign w2982 = w2885 & ~w2430;
assign w2983 = ~w2429 & w2982;
assign w2984 = ~w2974 & ~w2981;
assign w2985 = ~w2983 & w2984;
assign w2986 = ~w2490 & ~w2501;
assign w2987 = (~w726 & ~w2498) | (~w726 & w5609) | (~w2498 & w5609);
assign w2988 = ~w2499 & ~w2987;
assign w2989 = w2986 & ~w2988;
assign w2990 = ~w2986 & w2988;
assign w2991 = ~w2989 & ~w2990;
assign w2992 = (~w2991 & w2985) | (~w2991 & w6067) | (w2985 & w6067);
assign w2993 = (w726 & ~w2488) | (w726 & w6620) | (~w2488 & w6620);
assign w2994 = (w2993 & w2478) | (w2993 & w6621) | (w2478 & w6621);
assign w2995 = ~w2478 & w6622;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = (w2882 & w2460) | (w2882 & w5726) | (w2460 & w5726);
assign w2998 = (w2885 & w2460) | (w2885 & w5610) | (w2460 & w5610);
assign w2999 = ~w1823 & w6068;
assign w3000 = ~w2244 & w6069;
assign w3001 = (~w2999 & ~w1952) | (~w2999 & w6070) | (~w1952 & w6070);
assign w3002 = (w871 & ~w3001) | (w871 & w5727) | (~w3001 & w5727);
assign w3003 = w3001 & w5728;
assign w3004 = ~w3002 & ~w3003;
assign w3005 = ~w2998 & w3004;
assign w3006 = (~w2996 & w3005) | (~w2996 & w5729) | (w3005 & w5729);
assign w3007 = w6620 & ~w2488;
assign w3008 = ~w2489 & ~w3007;
assign w3009 = w2881 & ~w2889;
assign w3010 = w1819 & w3009;
assign w3011 = ~w1818 & w3009;
assign w3012 = w1716 & w3011;
assign w3013 = ~w1823 & w5611;
assign w3014 = w1704 & w2893;
assign w3015 = w1715 & w2891;
assign w3016 = ~w3014 & ~w3015;
assign w3017 = ~w3013 & w3016;
assign w3018 = ~w3012 & w3017;
assign w3019 = ~w3010 & w3018;
assign w3020 = ~w2036 & w3009;
assign w3021 = ~w1710 & w2891;
assign w3022 = w1704 & w2903;
assign w3023 = (~w3021 & ~w1715) | (~w3021 & w6071) | (~w1715 & w6071);
assign w3024 = ~w3022 & w3023;
assign w3025 = ~w1710 & w2881;
assign w3026 = ~w1710 & w3009;
assign w3027 = ~w1715 & w3026;
assign w3028 = ~w1710 & w2893;
assign w3029 = ~w1705 & w5612;
assign w3030 = ~w3028 & ~w3029;
assign w3031 = ~w3027 & w3030;
assign w3032 = w3031 & w5613;
assign w3033 = (w3020 & w6623) | (w3020 & w6624) | (w6623 & w6624);
assign w3034 = w3019 & ~w3033;
assign w3035 = ~w3020 & w7628;
assign w3036 = (w2483 & ~w3018) | (w2483 & w5730) | (~w3018 & w5730);
assign w3037 = ~w3035 & ~w3036;
assign w3038 = ~w3034 & w3037;
assign w3039 = w3008 & ~w3038;
assign w3040 = w3037 & w5616;
assign w3041 = ~w1816 & w6073;
assign w3042 = ~w1819 & w3041;
assign w3043 = ~w1955 & w3042;
assign w3044 = ~w1823 & w6074;
assign w3045 = w1704 & w2891;
assign w3046 = w1952 & w2903;
assign w3047 = ~w3044 & ~w3045;
assign w3048 = ~w3046 & w3047;
assign w3049 = ~w3043 & w3048;
assign w3050 = w3049 & w5617;
assign w3051 = (~w871 & ~w3049) | (~w871 & w5618) | (~w3049 & w5618);
assign w3052 = ~w3050 & ~w3051;
assign w3053 = ~w3040 & w3052;
assign w3054 = ~w3039 & ~w3053;
assign w3055 = ~w3006 & ~w3054;
assign w3056 = w2972 & w2991;
assign w3057 = ~w2985 & w3056;
assign w3058 = ~w3005 & w5731;
assign w3059 = ~w3057 & ~w3058;
assign w3060 = ~w3055 & w3059;
assign w3061 = ~w2992 & ~w3060;
assign w3062 = ~w2967 & w3061;
assign w3063 = w2962 & w2966;
assign w3064 = w2949 & w2953;
assign w3065 = ~w3063 & ~w3064;
assign w3066 = ~w3062 & w3065;
assign w3067 = ~w2954 & ~w3066;
assign w3068 = (~w2940 & w3066) | (~w2940 & w5732) | (w3066 & w5732);
assign w3069 = w2924 & ~w2939;
assign w3070 = w2532 & ~w2534;
assign w3071 = ~w2535 & ~w3070;
assign w3072 = w2772 & w2788;
assign w3073 = ~w2867 & ~w3072;
assign w3074 = ~w2655 & w2788;
assign w3075 = (w5591 & w6075) | (w5591 & w6076) | (w6075 & w6076);
assign w3076 = w3073 & ~w3075;
assign w3077 = ~w3073 & w3075;
assign w3078 = ~w3076 & ~w3077;
assign w3079 = w2882 & w3078;
assign w3080 = ~w2655 & w2891;
assign w3081 = w2865 & w6625;
assign w3082 = ~w3080 & ~w3081;
assign w3083 = (w871 & ~w3082) | (w871 & w6077) | (~w3082 & w6077);
assign w3084 = w3082 & w6078;
assign w3085 = ~w3083 & ~w3084;
assign w3086 = (w3085 & ~w3078) | (w3085 & w6079) | (~w3078 & w6079);
assign w3087 = ~w3079 & ~w3086;
assign w3088 = ~w3071 & ~w3087;
assign w3089 = (~w3069 & w3071) | (~w3069 & w5734) | (w3071 & w5734);
assign w3090 = ~w3068 & w3089;
assign w3091 = w3071 & w3087;
assign w3092 = ~w3090 & ~w3091;
assign w3093 = ~w2919 & w3092;
assign w3094 = w2919 & ~w3092;
assign w3095 = ~w3093 & ~w3094;
assign w3096 = ~w2835 & w2852;
assign w3097 = ~w124 & ~w265;
assign w3098 = ~w409 & ~w935;
assign w3099 = w3097 & w3098;
assign w3100 = w151 & w544;
assign w3101 = w3099 & w3100;
assign w3102 = w229 & ~w231;
assign w3103 = w415 & w590;
assign w3104 = w679 & w1788;
assign w3105 = w3103 & w3104;
assign w3106 = w444 & w3102;
assign w3107 = w3105 & w3106;
assign w3108 = w246 & w3101;
assign w3109 = w3107 & w3108;
assign w3110 = w1524 & w3109;
assign w3111 = w527 & w3110;
assign w3112 = (w3111 & ~w2852) | (w3111 & w6080) | (~w2852 & w6080);
assign w3113 = ~w2900 & w3112;
assign w3114 = ~w163 & ~w372;
assign w3115 = ~w197 & ~w456;
assign w3116 = ~w691 & w3115;
assign w3117 = ~w252 & w932;
assign w3118 = w932 & w6081;
assign w3119 = ~w183 & ~w204;
assign w3120 = ~w213 & ~w609;
assign w3121 = ~w217 & ~w769;
assign w3122 = ~w160 & ~w250;
assign w3123 = w1570 & w3122;
assign w3124 = w401 & w805;
assign w3125 = w2297 & w2740;
assign w3126 = w3119 & w3120;
assign w3127 = w3121 & w3126;
assign w3128 = w3124 & w3125;
assign w3129 = w3123 & w3128;
assign w3130 = w3118 & w3127;
assign w3131 = w3129 & w3130;
assign w3132 = ~w124 & ~w186;
assign w3133 = ~w210 & ~w273;
assign w3134 = w3132 & w3133;
assign w3135 = w1507 & w1899;
assign w3136 = w3114 & w3135;
assign w3137 = w2618 & w3134;
assign w3138 = w3116 & w3137;
assign w3139 = w795 & w3136;
assign w3140 = w3138 & w3139;
assign w3141 = w829 & w3140;
assign w3142 = w3131 & w3141;
assign w3143 = ~w2900 & w6082;
assign w3144 = ~w2898 & w6083;
assign w3145 = ~w2898 & w5619;
assign w3146 = (~w3142 & ~w5619) | (~w3142 & w5735) | (~w5619 & w5735);
assign w3147 = ~w3144 & ~w3146;
assign w3148 = ~a_0 & a_1;
assign w3149 = (w3148 & w3146) | (w3148 & w6084) | (w3146 & w6084);
assign w3150 = ~w226 & ~w373;
assign w3151 = ~w307 & ~w470;
assign w3152 = w599 & w3151;
assign w3153 = w757 & w1672;
assign w3154 = w2698 & w3150;
assign w3155 = w3153 & w3154;
assign w3156 = w3152 & w3155;
assign w3157 = w1031 & w1669;
assign w3158 = w2623 & w3157;
assign w3159 = w424 & w3156;
assign w3160 = w3158 & w3159;
assign w3161 = w1057 & w3160;
assign w3162 = ~w2898 & w6626;
assign w3163 = (w2898 & w6627) | (w2898 & w6628) | (w6627 & w6628);
assign w3164 = ~w3162 & ~w3163;
assign w3165 = ~a_0 & ~a_22;
assign w3166 = ~w3165 & w6085;
assign w3167 = (a_2 & w3165) | (a_2 & w6086) | (w3165 & w6086);
assign w3168 = ~w3166 & ~w3167;
assign w3169 = a_0 & w3168;
assign w3170 = ~w2900 & ~w3096;
assign w3171 = (~w3111 & ~w5622) | (~w3111 & w5736) | (~w5622 & w5736);
assign w3172 = ~w3145 & ~w3171;
assign w3173 = a_2 & w0;
assign w3174 = (w3173 & w3171) | (w3173 & w6087) | (w3171 & w6087);
assign w3175 = a_0 & ~w3168;
assign w3176 = w2852 & w6088;
assign w3177 = ~w3112 & ~w3176;
assign w3178 = w5608 & w5737;
assign w3179 = (w3177 & ~w5608) | (w3177 & w5738) | (~w5608 & w5738);
assign w3180 = ~w3178 & ~w3179;
assign w3181 = ~w2902 & w3180;
assign w3182 = w2868 & ~w3181;
assign w3183 = w2803 & w3182;
assign w3184 = ~w3147 & ~w3172;
assign w3185 = w3164 & w3184;
assign w3186 = w2866 & w2901;
assign w3187 = ~w3180 & ~w3186;
assign w3188 = w2901 & w7752;
assign w3189 = ~w3185 & ~w3188;
assign w3190 = (~w5736 & w6089) | (~w5736 & w6090) | (w6089 & w6090);
assign w3191 = (w5736 & w6091) | (w5736 & w6092) | (w6091 & w6092);
assign w3192 = ~w3190 & ~w3191;
assign w3193 = (~w5735 & w5687) | (~w5735 & w6093) | (w5687 & w6093);
assign w3194 = (w5735 & w5688) | (w5735 & w6094) | (w5688 & w6094);
assign w3195 = ~w3193 & ~w3194;
assign w3196 = ~w3192 & w3195;
assign w3197 = ~w3185 & ~w3196;
assign w3198 = ~w3197 & w7753;
assign w3199 = ~w3184 & ~w3195;
assign w3200 = ~w3184 & w6097;
assign w3201 = ~w3188 & w3199;
assign w3202 = (~w5740 & w6098) | (~w5740 & w6099) | (w6098 & w6099);
assign w3203 = ~w3198 & w3202;
assign w3204 = w6100 & w7754;
assign w3205 = (w3203 & w6629) | (w3203 & w6630) | (w6629 & w6630);
assign w3206 = ~w3204 & ~w3205;
assign w3207 = w3095 & w3206;
assign w3208 = ~w3095 & ~w3206;
assign w3209 = ~w3207 & ~w3208;
assign w3210 = ~w2967 & ~w3063;
assign w3211 = w3061 & ~w3210;
assign w3212 = ~w3061 & w3210;
assign w3213 = ~w3211 & ~w3212;
assign w3214 = w2788 & w3148;
assign w3215 = w2865 & w6631;
assign w3216 = ~w3214 & ~w3215;
assign w3217 = (w3078 & w6632) | (w3078 & w6633) | (w6632 & w6633);
assign w3218 = (~w2878 & w2655) | (~w2878 & w6101) | (w2655 & w6101);
assign w3219 = w3216 & w7755;
assign w3220 = ~w3217 & ~w3219;
assign w3221 = ~w3213 & ~w3220;
assign w3222 = w2901 & w6102;
assign w3223 = w2865 & w6634;
assign w3224 = w2788 & w3173;
assign w3225 = ~w3223 & ~w3224;
assign w3226 = (w2874 & w6635) | (w2874 & w6636) | (w6635 & w6636);
assign w3227 = (~w2874 & w6104) | (~w2874 & w6105) | (w6104 & w6105);
assign w3228 = ~w3226 & ~w3227;
assign w3229 = (~w3063 & ~w3061) | (~w3063 & w6106) | (~w3061 & w6106);
assign w3230 = ~w2954 & ~w3064;
assign w3231 = w3229 & w3230;
assign w3232 = ~w3229 & ~w3230;
assign w3233 = ~w3231 & ~w3232;
assign w3234 = w3228 & ~w3233;
assign w3235 = (~w3058 & w3054) | (~w3058 & w6107) | (w3054 & w6107);
assign w3236 = ~w2992 & ~w3057;
assign w3237 = ~w3235 & w3236;
assign w3238 = w3235 & ~w3236;
assign w3239 = ~w3237 & ~w3238;
assign w3240 = w2788 & w3169;
assign w3241 = ~w2655 & w3148;
assign w3242 = ~w2410 & w3173;
assign w3243 = ~w3241 & ~w3242;
assign w3244 = (w2925 & w6637) | (w2925 & w6638) | (w6637 & w6638);
assign w3245 = w2878 & w3244;
assign w3246 = (~w2878 & ~w3243) | (~w2878 & w7868) | (~w3243 & w7868);
assign w3247 = ~w3245 & ~w3246;
assign w3248 = ~w3239 & ~w3247;
assign w3249 = w3239 & w3247;
assign w3250 = ~w2655 & w3169;
assign w3251 = ~w2410 & w3148;
assign w3252 = (w2878 & w3250) | (w2878 & w7756) | (w3250 & w7756);
assign w3253 = (~w2878 & ~w2241) | (~w2878 & w6101) | (~w2241 & w6101);
assign w3254 = (w2664 & w6639) | (w2664 & w6640) | (w6639 & w6640);
assign w3255 = ~w3252 & ~w3254;
assign w3256 = ~w3006 & ~w3058;
assign w3257 = w3054 & ~w3256;
assign w3258 = ~w3054 & w3256;
assign w3259 = ~w3257 & ~w3258;
assign w3260 = ~w3255 & w3259;
assign w3261 = (w871 & w1710) | (w871 & w6108) | (w1710 & w6108);
assign w3262 = (w3020 & w7629) | (w3020 & w7630) | (w7629 & w7630);
assign w3263 = ~w3035 & ~w3262;
assign w3264 = ~w3019 & w3263;
assign w3265 = w3019 & ~w3263;
assign w3266 = ~w3264 & ~w3265;
assign w3267 = ~w2244 & w6109;
assign w3268 = ~w2429 & w2430;
assign w3269 = ~w2431 & ~w3268;
assign w3270 = w1952 & w3173;
assign w3271 = w2241 & w3169;
assign w3272 = ~w3267 & ~w3270;
assign w3273 = ~w3271 & w3272;
assign w3274 = w3273 & w7757;
assign w3275 = (w3266 & w3274) | (w3266 & w6112) | (w3274 & w6112);
assign w3276 = ~w2244 & w6113;
assign w3277 = ~w1823 & w6114;
assign w3278 = (w3175 & w2460) | (w3175 & w6115) | (w2460 & w6115);
assign w3279 = (~w3277 & ~w1952) | (~w3277 & w6116) | (~w1952 & w6116);
assign w3280 = ~w3276 & w3279;
assign w3281 = (~w2878 & w3278) | (~w2878 & w6117) | (w3278 & w6117);
assign w3282 = ~w3278 & w6118;
assign w3283 = ~w3281 & ~w3282;
assign w3284 = (~w871 & ~w3031) | (~w871 & w6119) | (~w3031 & w6119);
assign w3285 = (w3284 & w3020) | (w3284 & w6120) | (w3020 & w6120);
assign w3286 = ~w3020 & w6121;
assign w3287 = ~w3285 & ~w3286;
assign w3288 = ~w3283 & ~w3287;
assign w3289 = w3283 & w3287;
assign w3290 = (w6925 & ~w3031) | (w6925 & w6122) | (~w3031 & w6122);
assign w3291 = ~w3032 & ~w3290;
assign w3292 = ~w1823 & w6123;
assign w3293 = ~w1819 & ~w2024;
assign w3294 = w1704 & w3148;
assign w3295 = ~w3292 & ~w3294;
assign w3296 = (w3295 & w3293) | (w3295 & w6124) | (w3293 & w6124);
assign w3297 = (~w2878 & ~w1715) | (~w2878 & w6101) | (~w1715 & w6101);
assign w3298 = w3296 & ~w3297;
assign w3299 = a_0 & w1704;
assign w3300 = (~w0 & w3168) | (~w0 & w6125) | (w3168 & w6125);
assign w3301 = w1715 & w3300;
assign w3302 = w1710 & ~w2878;
assign w3303 = (w3302 & w1997) | (w3302 & w6126) | (w1997 & w6126);
assign w3304 = ~w3301 & w3303;
assign w3305 = ~w3299 & w3304;
assign w3306 = ~w3025 & ~w3305;
assign w3307 = (~w3306 & w3296) | (~w3306 & w6127) | (w3296 & w6127);
assign w3308 = ~w3298 & w3307;
assign w3309 = ~w3291 & ~w3308;
assign w3310 = w3291 & w3308;
assign w3311 = w1952 & w3169;
assign w3312 = w1704 & w3173;
assign w3313 = ~w1823 & w6128;
assign w3314 = w1822 & ~w1955;
assign w3315 = ~w1956 & ~w3314;
assign w3316 = ~w3312 & ~w3313;
assign w3317 = (~w3315 & w6641) | (~w3315 & w6642) | (w6641 & w6642);
assign w3318 = (w3315 & w6130) | (w3315 & w6131) | (w6130 & w6131);
assign w3319 = (~w3309 & ~w6132) | (~w3309 & w6643) | (~w6132 & w6643);
assign w3320 = ~w3289 & ~w3319;
assign w3321 = ~w3320 & w7733;
assign w3322 = ~w2244 & w6133;
assign w3323 = (~w3322 & ~w2241) | (~w3322 & w6135) | (~w2241 & w6135);
assign w3324 = (w6134 & w6644) | (w6134 & w6645) | (w6644 & w6645);
assign w3325 = (w6137 & ~w6134) | (w6137 & w6646) | (~w6134 & w6646);
assign w3326 = ~w3324 & ~w3325;
assign w3327 = ~w3039 & ~w3040;
assign w3328 = w3052 & w3327;
assign w3329 = ~w3052 & ~w3327;
assign w3330 = ~w3328 & ~w3329;
assign w3331 = ~w3274 & w6138;
assign w3332 = (~w3331 & ~w3330) | (~w3331 & w7734) | (~w3330 & w7734);
assign w3333 = ~w3321 & w3332;
assign w3334 = ~w3326 & ~w3330;
assign w3335 = (~w3334 & ~w3255) | (~w3334 & w6139) | (~w3255 & w6139);
assign w3336 = ~w3333 & w3335;
assign w3337 = ~w3249 & ~w3260;
assign w3338 = ~w3336 & w3337;
assign w3339 = (~w3248 & ~w3213) | (~w3248 & w6140) | (~w3213 & w6140);
assign w3340 = ~w3338 & w3339;
assign w3341 = ~w3221 & ~w3234;
assign w3342 = ~w3340 & w3341;
assign w3343 = ~w3069 & ~w3068;
assign w3344 = ~w3088 & ~w3091;
assign w3345 = (~w3188 & ~w2803) | (~w3188 & w5741) | (~w2803 & w5741);
assign w3346 = ~w3192 & w3345;
assign w3347 = w3192 & ~w3345;
assign w3348 = ~w3346 & ~w3347;
assign w3349 = (w3169 & w3146) | (w3169 & w6141) | (w3146 & w6141);
assign w3350 = (w3148 & w3171) | (w3148 & w6142) | (w3171 & w6142);
assign w3351 = w2901 & w6143;
assign w3352 = ~w3349 & ~w3350;
assign w3353 = (~w2878 & ~w3352) | (~w2878 & w7758) | (~w3352 & w7758);
assign w3354 = (w3348 & w6144) | (w3348 & w6145) | (w6144 & w6145);
assign w3355 = ~w3353 & ~w3354;
assign w3356 = w3344 & ~w3355;
assign w3357 = ~w3228 & w3233;
assign w3358 = (w3169 & w3171) | (w3169 & w6146) | (w3171 & w6146);
assign w3359 = w2901 & w6147;
assign w3360 = (w3187 & ~w2803) | (w3187 & w5742) | (~w2803 & w5742);
assign w3361 = (w2803 & w6148) | (w2803 & w6149) | (w6148 & w6149);
assign w3362 = ~w3360 & ~w3361;
assign w3363 = ~w3358 & ~w3359;
assign w3364 = (w2878 & w3358) | (w2878 & w7759) | (w3358 & w7759);
assign w3365 = (~w2878 & w6101) | (~w2878 & ~w2866) | (w6101 & ~w2866);
assign w3366 = (w3362 & w6647) | (w3362 & w6648) | (w6647 & w6648);
assign w3367 = ~w3364 & ~w3366;
assign w3368 = ~w2940 & ~w3069;
assign w3369 = w3067 & ~w3368;
assign w3370 = ~w3067 & w3368;
assign w3371 = ~w3369 & ~w3370;
assign w3372 = w3367 & w3371;
assign w3373 = ~w3344 & ~w3355;
assign w3374 = ~w3343 & w3373;
assign w3375 = (~w3357 & ~w3356) | (~w3357 & w6150) | (~w3356 & w6150);
assign w3376 = ~w3372 & ~w3374;
assign w3377 = w3376 & w6151;
assign w3378 = (~w3355 & w3371) | (~w3355 & w6152) | (w3371 & w6152);
assign w3379 = ~w3371 & w5743;
assign w3380 = w3343 & ~w3344;
assign w3381 = ~w3343 & w3344;
assign w3382 = ~w3380 & ~w3381;
assign w3383 = ~w3379 & w3382;
assign w3384 = ~w3378 & ~w3383;
assign w3385 = ~w3377 & ~w3384;
assign w3386 = w3209 & ~w3385;
assign w3387 = w2901 & w6153;
assign w3388 = w2865 & w6649;
assign w3389 = (w2903 & w3171) | (w2903 & w6154) | (w3171 & w6154);
assign w3390 = ~w3387 & ~w3388;
assign w3391 = ~w3389 & w3390;
assign w3392 = (~w871 & ~w3391) | (~w871 & w7760) | (~w3391 & w7760);
assign w3393 = (w3362 & w6155) | (w3362 & w6156) | (w6155 & w6156);
assign w3394 = ~w3392 & ~w3393;
assign w3395 = ~w2419 & ~w2674;
assign w3396 = ~w2535 & w3395;
assign w3397 = ~w2673 & ~w3396;
assign w3398 = ~w2925 & w6650;
assign w3399 = w2402 & ~w2655;
assign w3400 = w2405 & ~w2410;
assign w3401 = ~w3399 & ~w3400;
assign w3402 = w3401 & w6651;
assign w3403 = (w726 & ~w3401) | (w726 & w6652) | (~w3401 & w6652);
assign w3404 = ~w3402 & ~w3403;
assign w3405 = (w3404 & ~w2930) | (w3404 & w6157) | (~w2930 & w6157);
assign w3406 = ~w3398 & ~w3405;
assign w3407 = w2552 & w2576;
assign w3408 = ~w2578 & ~w3407;
assign w3409 = w2563 & w3269;
assign w3410 = w1952 & w1974;
assign w3411 = ~w2244 & w6158;
assign w3412 = ~w3410 & ~w3411;
assign w3413 = ~w2229 & w5623;
assign w3414 = w1968 & ~w2204;
assign w3415 = (w3414 & w2229) | (w3414 & w5624) | (w2229 & w5624);
assign w3416 = ~w3413 & ~w3415;
assign w3417 = ~w565 & w3416;
assign w3418 = w3412 & w3417;
assign w3419 = w2429 & w5744;
assign w3420 = w2430 & w3418;
assign w3421 = ~w2429 & w3420;
assign w3422 = w3412 & w5745;
assign w3423 = (w565 & ~w3412) | (w565 & w5746) | (~w3412 & w5746);
assign w3424 = ~w3422 & ~w3423;
assign w3425 = ~w3421 & w3424;
assign w3426 = ~w3419 & w3425;
assign w3427 = w2541 & w2549;
assign w3428 = ~w2543 & w3427;
assign w3429 = ~w1022 & w1710;
assign w3430 = ~w3428 & w3429;
assign w3431 = w3428 & w5625;
assign w3432 = ~w3430 & ~w3431;
assign w3433 = w1994 & ~w3293;
assign w3434 = w1715 & w2546;
assign w3435 = ~w1823 & w6159;
assign w3436 = w1704 & w1991;
assign w3437 = ~w3434 & ~w3436;
assign w3438 = ~w3435 & w3437;
assign w3439 = ~w3433 & w3438;
assign w3440 = ~w3432 & w3439;
assign w3441 = w3432 & ~w3439;
assign w3442 = ~w3440 & ~w3441;
assign w3443 = (w3442 & ~w3426) | (w3442 & w6160) | (~w3426 & w6160);
assign w3444 = w3426 & w6161;
assign w3445 = ~w3443 & ~w3444;
assign w3446 = w3408 & w3445;
assign w3447 = ~w3408 & ~w3445;
assign w3448 = ~w3446 & ~w3447;
assign w3449 = ~w3406 & ~w3448;
assign w3450 = w3406 & w3448;
assign w3451 = ~w3449 & ~w3450;
assign w3452 = w3397 & ~w3451;
assign w3453 = ~w3397 & w3451;
assign w3454 = ~w3452 & ~w3453;
assign w3455 = w3394 & ~w3454;
assign w3456 = ~w3394 & w3454;
assign w3457 = ~w3455 & ~w3456;
assign w3458 = w2915 & ~w3091;
assign w3459 = (~w2918 & ~w3458) | (~w2918 & w5747) | (~w3458 & w5747);
assign w3460 = w3457 & w3459;
assign w3461 = ~w3457 & ~w3459;
assign w3462 = ~w3460 & ~w3461;
assign w3463 = ~w119 & w628;
assign w3464 = w613 & ~w935;
assign w3465 = w1034 & w1039;
assign w3466 = w3463 & w3465;
assign w3467 = w399 & w3464;
assign w3468 = w908 & w3467;
assign w3469 = w424 & w3466;
assign w3470 = w1049 & w3469;
assign w3471 = w3468 & w3470;
assign w3472 = ~w2898 & w6653;
assign w3473 = (w2898 & ~w3471) | (w2898 & w6654) | (~w3471 & w6654);
assign w3474 = ~w3472 & ~w3473;
assign w3475 = (w3173 & w3146) | (w3173 & w6164) | (w3146 & w6164);
assign w3476 = w3148 & ~w3164;
assign w3477 = ~w3147 & ~w3164;
assign w3478 = w3164 & w3471;
assign w3479 = ~w3164 & ~w3474;
assign w3480 = ~w3478 & ~w3479;
assign w3481 = (w6096 & w7287) | (w6096 & w7288) | (w7287 & w7288);
assign w3482 = w6166 & w7761;
assign w3483 = ~w3481 & ~w3482;
assign w3484 = ~w3475 & ~w3476;
assign w3485 = (w3483 & w6655) | (w3483 & w6656) | (w6655 & w6656);
assign w3486 = w3484 & w7762;
assign w3487 = ~w3485 & ~w3486;
assign w3488 = w3462 & w3487;
assign w3489 = (~w3207 & ~w3462) | (~w3207 & w5748) | (~w3462 & w5748);
assign w3490 = ~w3386 & w3489;
assign w3491 = ~w3462 & ~w3487;
assign w3492 = (~w3455 & ~w3457) | (~w3455 & w5749) | (~w3457 & w5749);
assign w3493 = ~w3397 & ~w3449;
assign w3494 = (~w3450 & w3397) | (~w3450 & w5750) | (w3397 & w5750);
assign w3495 = ~w1022 & ~w1715;
assign w3496 = ~w1823 & w6167;
assign w3497 = w1704 & w2546;
assign w3498 = w1952 & w1987;
assign w3499 = ~w3496 & ~w3497;
assign w3500 = (w3495 & w3498) | (w3495 & w6168) | (w3498 & w6168);
assign w3501 = ~w3498 & w6169;
assign w3502 = ~w3500 & ~w3501;
assign w3503 = (~w3502 & w3315) | (~w3502 & w6170) | (w3315 & w6170);
assign w3504 = (~w1022 & w3428) | (~w1022 & w5625) | (w3428 & w5625);
assign w3505 = w3439 & w3504;
assign w3506 = ~w1715 & w5775;
assign w3507 = ~w3315 & w3506;
assign w3508 = w3505 & ~w3507;
assign w3509 = ~w3503 & w3508;
assign w3510 = (~w3505 & w3503) | (~w3505 & w5626) | (w3503 & w5626);
assign w3511 = ~w3509 & ~w3510;
assign w3512 = ~w2244 & w6171;
assign w3513 = (~w3512 & ~w2241) | (~w3512 & w6172) | (~w2241 & w6172);
assign w3514 = (~w565 & ~w3513) | (~w565 & w5751) | (~w3513 & w5751);
assign w3515 = w3513 & w5752;
assign w3516 = ~w3514 & ~w3515;
assign w3517 = ~w2390 & w3516;
assign w3518 = w3513 & w5753;
assign w3519 = ~w3514 & ~w3518;
assign w3520 = w2390 & w3519;
assign w3521 = ~w3517 & ~w3520;
assign w3522 = w3511 & w3521;
assign w3523 = ~w3511 & ~w3521;
assign w3524 = ~w3522 & ~w3523;
assign w3525 = w3408 & ~w3444;
assign w3526 = (~w3443 & ~w3408) | (~w3443 & w5627) | (~w3408 & w5627);
assign w3527 = w3524 & ~w3526;
assign w3528 = ~w3524 & w3526;
assign w3529 = ~w3527 & ~w3528;
assign w3530 = w2394 & w3078;
assign w3531 = w2405 & ~w2655;
assign w3532 = w2865 & w6657;
assign w3533 = ~w3531 & ~w3532;
assign w3534 = (w726 & ~w3533) | (w726 & w6173) | (~w3533 & w6173);
assign w3535 = w3533 & w6174;
assign w3536 = ~w3534 & ~w3535;
assign w3537 = (w3536 & ~w3078) | (w3536 & w6175) | (~w3078 & w6175);
assign w3538 = ~w3530 & ~w3537;
assign w3539 = ~w3529 & ~w3538;
assign w3540 = w3529 & w3538;
assign w3541 = ~w3539 & ~w3540;
assign w3542 = w3494 & ~w3541;
assign w3543 = ~w3494 & w3541;
assign w3544 = ~w3542 & ~w3543;
assign w3545 = ~w133 & ~w411;
assign w3546 = ~w56 & w149;
assign w3547 = w3545 & ~w3546;
assign w3548 = w1031 & w3547;
assign w3549 = w1046 & w3548;
assign w3550 = w917 & w3549;
assign w3551 = w424 & w3550;
assign w3552 = ~w3471 & ~w3551;
assign w3553 = (w2898 & w3552) | (w2898 & w6658) | (w3552 & w6658);
assign w3554 = w3471 & w3550;
assign w3555 = (~w3554 & ~w3164) | (~w3554 & w6177) | (~w3164 & w6177);
assign w3556 = ~w3553 & w3555;
assign w3557 = (w3556 & w3185) | (w3556 & w6178) | (w3185 & w6178);
assign w3558 = ~w3553 & ~w3554;
assign w3559 = ~w3161 & w3471;
assign w3560 = (~w5735 & w6181) | (~w5735 & w6182) | (w6181 & w6182);
assign w3561 = ~w3164 & ~w3560;
assign w3562 = w3558 & ~w3561;
assign w3563 = ~w3558 & w3561;
assign w3564 = ~w3562 & ~w3563;
assign w3565 = ~w3564 & w7763;
assign w3566 = ~w3478 & ~w3558;
assign w3567 = (w6096 & w7289) | (w6096 & w7290) | (w7289 & w7290);
assign w3568 = ~w3565 & ~w3567;
assign w3569 = ~w3472 & w6183;
assign w3570 = ~w3164 & w3173;
assign w3571 = ~w3569 & ~w3570;
assign w3572 = (w3568 & w6659) | (w3568 & w6660) | (w6659 & w6660);
assign w3573 = (~w2878 & ~w3571) | (~w2878 & w7764) | (~w3571 & w7764);
assign w3574 = ~w3572 & ~w3573;
assign w3575 = w2882 & ~w3348;
assign w3576 = (w2893 & w3171) | (w2893 & w6184) | (w3171 & w6184);
assign w3577 = (w2903 & w3146) | (w2903 & w6185) | (w3146 & w6185);
assign w3578 = w2901 & w6186;
assign w3579 = ~w3576 & ~w3577;
assign w3580 = (w871 & ~w3579) | (w871 & w6187) | (~w3579 & w6187);
assign w3581 = w3579 & w6188;
assign w3582 = ~w3580 & ~w3581;
assign w3583 = (w3582 & w3348) | (w3582 & w6189) | (w3348 & w6189);
assign w3584 = ~w3575 & ~w3583;
assign w3585 = ~w3584 & w3574;
assign w3586 = (w3584 & w3572) | (w3584 & w6190) | (w3572 & w6190);
assign w3587 = ~w3585 & ~w3586;
assign w3588 = w3544 & ~w3587;
assign w3589 = ~w3544 & w3587;
assign w3590 = ~w3588 & ~w3589;
assign w3591 = w3492 & w3590;
assign w3592 = ~w3492 & ~w3590;
assign w3593 = ~w3591 & ~w3592;
assign w3594 = ~w3491 & w3593;
assign w3595 = ~w3490 & w3594;
assign w3596 = ~w3593 & w7765;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = w304 & ~w460;
assign w3599 = w539 & w3598;
assign w3600 = w3123 & w3599;
assign w3601 = w328 & w3600;
assign w3602 = ~w275 & ~w307;
assign w3603 = ~w181 & ~w205;
assign w3604 = ~w314 & ~w329;
assign w3605 = ~w124 & ~w411;
assign w3606 = ~w480 & w3605;
assign w3607 = w1789 & w3606;
assign w3608 = ~w186 & w1047;
assign w3609 = w3603 & w3604;
assign w3610 = w3608 & w3609;
assign w3611 = w2301 & w3610;
assign w3612 = w3607 & w3611;
assign w3613 = ~w196 & w3602;
assign w3614 = w3611 & w6191;
assign w3615 = w2817 & w3116;
assign w3616 = ~w166 & ~w211;
assign w3617 = ~w227 & ~w457;
assign w3618 = w677 & w3617;
assign w3619 = w2621 & w3119;
assign w3620 = w3616 & w3619;
assign w3621 = w3618 & w3620;
assign w3622 = w3615 & w3621;
assign w3623 = w361 & w3622;
assign w3624 = w3623 & w6192;
assign w3625 = ~w3597 & w3624;
assign w3626 = w928 & w1665;
assign w3627 = w2751 & w3626;
assign w3628 = w2179 & w3627;
assign w3629 = ~w159 & ~w199;
assign w3630 = w926 & w3629;
assign w3631 = w2824 & w3630;
assign w3632 = w216 & w531;
assign w3633 = ~w163 & ~w258;
assign w3634 = ~w324 & w3633;
assign w3635 = w471 & w1047;
assign w3636 = w1505 & w1658;
assign w3637 = w2619 & w3636;
assign w3638 = w3634 & w3635;
assign w3639 = w3632 & w3638;
assign w3640 = w3637 & w3639;
assign w3641 = w1911 & w3628;
assign w3642 = w3640 & w3641;
assign w3643 = w3631 & w3642;
assign w3644 = ~w3209 & w3385;
assign w3645 = (~w3643 & ~w3209) | (~w3643 & w6193) | (~w3209 & w6193);
assign w3646 = w600 & w1666;
assign w3647 = ~w362 & w931;
assign w3648 = w1558 & w1908;
assign w3649 = w3114 & w3119;
assign w3650 = w3648 & w3649;
assign w3651 = w3646 & w3647;
assign w3652 = w3650 & w3651;
assign w3653 = ~w147 & ~w210;
assign w3654 = ~w484 & w3653;
assign w3655 = ~w654 & ~w688;
assign w3656 = w242 & w601;
assign w3657 = w614 & w3655;
assign w3658 = w3656 & w3657;
assign w3659 = w1913 & w3658;
assign w3660 = w632 & w3659;
assign w3661 = w929 & w6194;
assign w3662 = w3660 & w3661;
assign w3663 = ~w347 & ~w435;
assign w3664 = ~w205 & ~w309;
assign w3665 = ~w199 & ~w234;
assign w3666 = w3120 & w3665;
assign w3667 = w3663 & w3664;
assign w3668 = w3666 & w3667;
assign w3669 = w3654 & w3668;
assign w3670 = w1514 & w3669;
assign w3671 = w3652 & w3670;
assign w3672 = w3662 & w3671;
assign w3673 = w3645 & w6661;
assign w3674 = (w3672 & ~w3645) | (w3672 & w6662) | (~w3645 & w6662);
assign w3675 = (~w3207 & ~w3209) | (~w3207 & w6195) | (~w3209 & w6195);
assign w3676 = ~w3488 & ~w3491;
assign w3677 = ~w3675 & w3676;
assign w3678 = w3675 & ~w3676;
assign w3679 = ~w3677 & ~w3678;
assign w3680 = (~w3673 & ~w3679) | (~w3673 & w6663) | (~w3679 & w6663);
assign w3681 = ~w3625 & ~w3680;
assign w3682 = w3597 & ~w3624;
assign w3683 = w3574 & ~w3593;
assign w3684 = (~w3683 & w3490) | (~w3683 & w5755) | (w3490 & w5755);
assign w3685 = w3544 & ~w3584;
assign w3686 = w3543 & w3584;
assign w3687 = ~w3541 & w3584;
assign w3688 = w3494 & w3687;
assign w3689 = ~w3455 & ~w3688;
assign w3690 = ~w3686 & w3689;
assign w3691 = ~w3460 & w3690;
assign w3692 = ~w3450 & ~w3540;
assign w3693 = ~w3493 & w3692;
assign w3694 = ~w3539 & ~w3693;
assign w3695 = w2882 & w3203;
assign w3696 = w2885 & ~w3200;
assign w3697 = w3696 & w7766;
assign w3698 = ~w3198 & w3697;
assign w3699 = (w2893 & w3146) | (w2893 & w6196) | (w3146 & w6196);
assign w3700 = (w2891 & w3171) | (w2891 & w6197) | (w3171 & w6197);
assign w3701 = (w871 & ~w6198) | (w871 & w6664) | (~w6198 & w6664);
assign w3702 = w6198 & w6665;
assign w3703 = ~w3701 & ~w3702;
assign w3704 = ~w3698 & w3703;
assign w3705 = ~w3695 & ~w3704;
assign w3706 = w2394 & ~w2874;
assign w3707 = w2405 & w2788;
assign w3708 = w2865 & w6666;
assign w3709 = w2901 & w6199;
assign w3710 = ~w3707 & ~w3708;
assign w3711 = w3710 & w6200;
assign w3712 = (w726 & ~w3710) | (w726 & w6201) | (~w3710 & w6201);
assign w3713 = ~w3711 & ~w3712;
assign w3714 = (w3713 & w2874) | (w3713 & w6202) | (w2874 & w6202);
assign w3715 = ~w3706 & ~w3714;
assign w3716 = ~w3705 & ~w3715;
assign w3717 = w3705 & w3715;
assign w3718 = ~w3716 & ~w3717;
assign w3719 = ~w3443 & ~w3523;
assign w3720 = (~w3522 & w3525) | (~w3522 & w5628) | (w3525 & w5628);
assign w3721 = ~w1022 & w3501;
assign w3722 = (w3721 & w3315) | (w3721 & w6203) | (w3315 & w6203);
assign w3723 = (~w3722 & ~w3508) | (~w3722 & w6591) | (~w3508 & w6591);
assign w3724 = (w1994 & w2460) | (w1994 & w5629) | (w2460 & w5629);
assign w3725 = ~w1022 & ~w1704;
assign w3726 = ~w1823 & w6204;
assign w3727 = ~w2244 & w6205;
assign w3728 = (~w3726 & ~w1952) | (~w3726 & w6206) | (~w1952 & w6206);
assign w3729 = ~w3727 & w3728;
assign w3730 = ~w3725 & ~w3729;
assign w3731 = w3725 & w3729;
assign w3732 = ~w3730 & ~w3731;
assign w3733 = ~w3724 & w3732;
assign w3734 = w3724 & w3725;
assign w3735 = ~w3733 & ~w3734;
assign w3736 = w3723 & ~w3735;
assign w3737 = ~w3723 & w3735;
assign w3738 = ~w3736 & ~w3737;
assign w3739 = w1968 & ~w2655;
assign w3740 = w1974 & w2241;
assign w3741 = (w3739 & w7291) | (w3739 & w7292) | (w7291 & w7292);
assign w3742 = ~w3739 & w7293;
assign w3743 = ~w3741 & ~w3742;
assign w3744 = w2664 & w3743;
assign w3745 = ~w3739 & w7294;
assign w3746 = ~w3741 & ~w3745;
assign w3747 = ~w2664 & w3746;
assign w3748 = ~w3744 & ~w3747;
assign w3749 = w3738 & ~w3748;
assign w3750 = ~w3738 & w3748;
assign w3751 = ~w3749 & ~w3750;
assign w3752 = w3720 & w3751;
assign w3753 = ~w3720 & ~w3751;
assign w3754 = ~w3752 & ~w3753;
assign w3755 = w3718 & ~w3754;
assign w3756 = ~w3718 & w3754;
assign w3757 = ~w3755 & ~w3756;
assign w3758 = w3694 & w3757;
assign w3759 = ~w3694 & ~w3757;
assign w3760 = ~w3758 & ~w3759;
assign w3761 = (~w3760 & w3691) | (~w3760 & w5756) | (w3691 & w5756);
assign w3762 = ~w3685 & w3760;
assign w3763 = ~w3691 & w3762;
assign w3764 = ~w3761 & ~w3763;
assign w3765 = ~w296 & ~w457;
assign w3766 = ~w514 & ~w691;
assign w3767 = w3765 & w3766;
assign w3768 = w374 & w1547;
assign w3769 = w3604 & w3768;
assign w3770 = w3767 & w3769;
assign w3771 = ~w109 & ~w205;
assign w3772 = ~w237 & w3771;
assign w3773 = w469 & w821;
assign w3774 = w1672 & w1788;
assign w3775 = w3773 & w3774;
assign w3776 = w293 & w3772;
assign w3777 = w3775 & w3776;
assign w3778 = w2820 & w3777;
assign w3779 = w3770 & w3778;
assign w3780 = w608 & w3779;
assign w3781 = (w3169 & ~w3779) | (w3169 & w6210) | (~w3779 & w6210);
assign w3782 = ~w3472 & w6211;
assign w3783 = (w3780 & w3472) | (w3780 & w6212) | (w3472 & w6212);
assign w3784 = ~w3782 & ~w3783;
assign w3785 = w3555 & ~w3562;
assign w3786 = ~w3557 & ~w3785;
assign w3787 = w3189 & ~w3785;
assign w3788 = ~w3183 & w3787;
assign w3789 = (w3784 & w5757) | (w3784 & w3788) | (w5757 & w3788);
assign w3790 = ~w3788 & w6213;
assign w3791 = (~w3781 & w3474) | (~w3781 & w6214) | (w3474 & w6214);
assign w3792 = w3791 & w7869;
assign w3793 = (w3790 & w7295) | (w3790 & w7296) | (w7295 & w7296);
assign w3794 = ~w3792 & ~w3793;
assign w3795 = ~w241 & ~w467;
assign w3796 = ~w538 & w3795;
assign w3797 = w664 & w3604;
assign w3798 = w3796 & w3797;
assign w3799 = w448 & w516;
assign w3800 = w3116 & w3799;
assign w3801 = w146 & w3798;
assign w3802 = w3800 & w3801;
assign w3803 = w173 & w263;
assign w3804 = w3802 & w3803;
assign w3805 = w2172 & w3804;
assign w3806 = ~w3792 & w6215;
assign w3807 = (w3805 & w3792) | (w3805 & w6216) | (w3792 & w6216);
assign w3808 = ~w3806 & ~w3807;
assign w3809 = w3764 & ~w3808;
assign w3810 = ~w3764 & w3808;
assign w3811 = ~w3809 & ~w3810;
assign w3812 = w3684 & w3811;
assign w3813 = ~w3684 & ~w3811;
assign w3814 = ~w3812 & ~w3813;
assign w3815 = ~w3682 & w3814;
assign w3816 = ~w3681 & w3815;
assign w3817 = ~w3681 & ~w3682;
assign w3818 = ~w3814 & ~w3817;
assign w3819 = ~w3816 & ~w3818;
assign w3820 = ~w3625 & ~w3682;
assign w3821 = w3680 & ~w3820;
assign w3822 = ~w3680 & w3820;
assign w3823 = ~w3821 & ~w3822;
assign w3824 = ~w3819 & w3823;
assign w3825 = w3819 & ~w3823;
assign w3826 = ~w3824 & ~w3825;
assign w3827 = ~a_22 & ~a_23;
assign w3828 = a_22 & a_23;
assign w3829 = ~w3827 & ~w3828;
assign w3830 = w3826 & w3829;
assign w3831 = w3805 & ~w3814;
assign w3832 = ~w3816 & ~w3831;
assign w3833 = ~w3764 & ~w3794;
assign w3834 = ~w3763 & w3794;
assign w3835 = ~w3761 & w3834;
assign w3836 = ~w3683 & ~w3835;
assign w3837 = (~w3833 & ~w3836) | (~w3833 & w6592) | (~w3836 & w6592);
assign w3838 = ~w180 & w529;
assign w3839 = ~w271 & w3663;
assign w3840 = ~w237 & ~w654;
assign w3841 = w219 & w3840;
assign w3842 = w623 & w1660;
assign w3843 = w3841 & w3842;
assign w3844 = w260 & w3116;
assign w3845 = w3838 & w3839;
assign w3846 = w3844 & w3845;
assign w3847 = w3118 & w3843;
assign w3848 = w3846 & w3847;
assign w3849 = w2322 & w3848;
assign w3850 = w3612 & w3849;
assign w3851 = w3705 & ~w3760;
assign w3852 = ~w3763 & ~w3851;
assign w3853 = w3715 & w3754;
assign w3854 = (~w3539 & w3754) | (~w3539 & w6217) | (w3754 & w6217);
assign w3855 = ~w3693 & w3854;
assign w3856 = (~w3853 & w3693) | (~w3853 & w6595) | (w3693 & w6595);
assign w3857 = w3524 & ~w3750;
assign w3858 = w3526 & w3857;
assign w3859 = (w3522 & w3738) | (w3522 & w5630) | (w3738 & w5630);
assign w3860 = ~w3749 & ~w3859;
assign w3861 = ~w3858 & w3860;
assign w3862 = (w1963 & w2656) | (w1963 & w6667) | (w2656 & w6667);
assign w3863 = w1963 & w2927;
assign w3864 = ~w2385 & w3863;
assign w3865 = (~w3862 & w2385) | (~w3862 & w6668) | (w2385 & w6668);
assign w3866 = w2929 & ~w3865;
assign w3867 = w1976 & ~w2655;
assign w3868 = w1974 & ~w2410;
assign w3869 = ~w3867 & ~w3868;
assign w3870 = (w565 & w3866) | (w565 & w6218) | (w3866 & w6218);
assign w3871 = ~w3866 & w6219;
assign w3872 = ~w3870 & ~w3871;
assign w3873 = ~w1022 & w1704;
assign w3874 = w3729 & w3873;
assign w3875 = ~w3724 & w3874;
assign w3876 = (~w3875 & w3723) | (~w3875 & w5631) | (w3723 & w5631);
assign w3877 = ~w2248 & w5758;
assign w3878 = w2429 & w3877;
assign w3879 = (w1994 & w2248) | (w1994 & w5759) | (w2248 & w5759);
assign w3880 = ~w2429 & w3879;
assign w3881 = ~w3878 & ~w3880;
assign w3882 = (~w1022 & w1823) | (~w1022 & w6220) | (w1823 & w6220);
assign w3883 = ~w2244 & w6221;
assign w3884 = w1952 & w2546;
assign w3885 = w1987 & w2241;
assign w3886 = ~w3883 & ~w3884;
assign w3887 = (~w3882 & w3885) | (~w3882 & w6222) | (w3885 & w6222);
assign w3888 = ~w3885 & w6223;
assign w3889 = ~w3887 & ~w3888;
assign w3890 = w3881 & w3889;
assign w3891 = ~w3881 & w3882;
assign w3892 = ~w3890 & ~w3891;
assign w3893 = w3876 & ~w3892;
assign w3894 = ~w3876 & w3892;
assign w3895 = ~w3893 & ~w3894;
assign w3896 = w3872 & w3895;
assign w3897 = ~w3872 & ~w3895;
assign w3898 = ~w3896 & ~w3897;
assign w3899 = w3861 & ~w3898;
assign w3900 = ~w3861 & w3898;
assign w3901 = ~w3899 & ~w3900;
assign w3902 = (w2411 & w3171) | (w2411 & w6224) | (w3171 & w6224);
assign w3903 = w2865 & w6669;
assign w3904 = w2901 & w6225;
assign w3905 = ~w3902 & ~w3903;
assign w3906 = (w726 & ~w3905) | (w726 & w7768) | (~w3905 & w7768);
assign w3907 = (w3362 & w6226) | (w3362 & w6227) | (w6226 & w6227);
assign w3908 = ~w3906 & ~w3907;
assign w3909 = w3901 & w3908;
assign w3910 = ~w3901 & ~w3908;
assign w3911 = ~w3909 & ~w3910;
assign w3912 = w3856 & w3911;
assign w3913 = ~w3856 & ~w3911;
assign w3914 = ~w3912 & ~w3913;
assign w3915 = w2893 & ~w3164;
assign w3916 = (w2891 & w3146) | (w2891 & w6228) | (w3146 & w6228);
assign w3917 = ~w3915 & ~w3916;
assign w3918 = w3917 & w7769;
assign w3919 = (w3483 & w6229) | (w3483 & w6230) | (w6229 & w6230);
assign w3920 = ~w3918 & ~w3919;
assign w3921 = ~w237 & ~w460;
assign w3922 = w322 & w3921;
assign w3923 = w1658 & w1660;
assign w3924 = w2298 & w3923;
assign w3925 = w3922 & w3924;
assign w3926 = w414 & w3925;
assign w3927 = ~w204 & ~w513;
assign w3928 = w757 & w3927;
assign w3929 = ~w164 & ~w309;
assign w3930 = ~w688 & w3929;
assign w3931 = w331 & w3930;
assign w3932 = w3928 & w3931;
assign w3933 = w537 & w3932;
assign w3934 = w927 & w3933;
assign w3935 = w1683 & w3926;
assign w3936 = w3934 & w3935;
assign w3937 = (w3936 & w3472) | (w3936 & w6231) | (w3472 & w6231);
assign w3938 = ~w3472 & w6232;
assign w3939 = ~w3937 & ~w3938;
assign w3940 = ~w3789 & w6233;
assign w3941 = (w3939 & w3789) | (w3939 & w6234) | (w3789 & w6234);
assign w3942 = ~w3940 & ~w3941;
assign w3943 = w3169 & ~w3936;
assign w3944 = (w3148 & ~w3779) | (w3148 & w6235) | (~w3779 & w6235);
assign w3945 = (w6238 & ~w3942) | (w6238 & w6670) | (~w3942 & w6670);
assign w3946 = (w3942 & w6671) | (w3942 & w6672) | (w6671 & w6672);
assign w3947 = ~w3945 & ~w3946;
assign w3948 = w3920 & ~w3947;
assign w3949 = ~w3920 & w3947;
assign w3950 = ~w3948 & ~w3949;
assign w3951 = w3914 & ~w3950;
assign w3952 = ~w3914 & w3950;
assign w3953 = ~w3951 & ~w3952;
assign w3954 = w3852 & w3953;
assign w3955 = ~w3852 & ~w3953;
assign w3956 = ~w3954 & ~w3955;
assign w3957 = ~w3850 & w3956;
assign w3958 = w3850 & ~w3956;
assign w3959 = ~w3957 & ~w3958;
assign w3960 = w3837 & w3959;
assign w3961 = ~w3837 & ~w3959;
assign w3962 = ~w3960 & ~w3961;
assign w3963 = ~w3816 & w6239;
assign w3964 = (~w3962 & w3816) | (~w3962 & w6240) | (w3816 & w6240);
assign w3965 = ~w3963 & ~w3964;
assign w3966 = w3826 & w6241;
assign w3967 = w3824 & ~w3965;
assign w3968 = ~w3824 & w3965;
assign w3969 = ~w3967 & ~w3968;
assign w3970 = ~w3830 & w3969;
assign w3971 = ~w3966 & ~w3970;
assign w3972 = ~w3805 & ~w3814;
assign w3973 = ~w3850 & ~w3956;
assign w3974 = ~w3837 & ~w3973;
assign w3975 = w3837 & ~w3957;
assign w3976 = ~w3974 & ~w3975;
assign w3977 = ~w3972 & ~w3976;
assign w3978 = w3850 & w3956;
assign w3979 = ~w3837 & ~w3978;
assign w3980 = w3837 & ~w3958;
assign w3981 = ~w3979 & ~w3980;
assign w3982 = ~w3977 & ~w3981;
assign w3983 = w3814 & ~w3981;
assign w3984 = ~w3817 & w3983;
assign w3985 = ~w3982 & ~w3984;
assign w3986 = ~w3947 & w3956;
assign w3987 = w3837 & ~w3986;
assign w3988 = ~w3914 & ~w3920;
assign w3989 = ~w3911 & w3920;
assign w3990 = w3856 & w3989;
assign w3991 = w3911 & w3920;
assign w3992 = ~w3856 & w3991;
assign w3993 = ~w3990 & ~w3992;
assign w3994 = ~w3851 & w3993;
assign w3995 = (~w3988 & ~w3994) | (~w3988 & w5632) | (~w3994 & w5632);
assign w3996 = ~w3853 & ~w3910;
assign w3997 = (~w3909 & ~w3996) | (~w3909 & w5633) | (~w3996 & w5633);
assign w3998 = (~w3896 & w3861) | (~w3896 & w5760) | (w3861 & w5760);
assign w3999 = ~w1823 & w6242;
assign w4000 = ~w3885 & w6243;
assign w4001 = w3881 & w4000;
assign w4002 = ~w3892 & ~w4001;
assign w4003 = ~w3875 & ~w4001;
assign w4004 = ~w3737 & w4003;
assign w4005 = ~w4002 & ~w4004;
assign w4006 = ~w1022 & ~w1952;
assign w4007 = (w1994 & ~w2248) | (w1994 & w6244) | (~w2248 & w6244);
assign w4008 = ~w2388 & w4007;
assign w4009 = ~w2244 & w6245;
assign w4010 = w1987 & ~w2410;
assign w4011 = (~w4009 & ~w2241) | (~w4009 & w6246) | (~w2241 & w6246);
assign w4012 = ~w4010 & w4011;
assign w4013 = (w4012 & ~w4008) | (w4012 & w5634) | (~w4008 & w5634);
assign w4014 = w4006 & ~w4013;
assign w4015 = ~w4006 & w4013;
assign w4016 = ~w4014 & ~w4015;
assign w4017 = (w4016 & w4004) | (w4016 & w5635) | (w4004 & w5635);
assign w4018 = ~w4004 & w5636;
assign w4019 = ~w4017 & ~w4018;
assign w4020 = (w1963 & w2867) | (w1963 & w6673) | (w2867 & w6673);
assign w4021 = ~w3075 & w4020;
assign w4022 = ~w2789 & ~w2867;
assign w4023 = (w4022 & w3864) | (w4022 & w5761) | (w3864 & w5761);
assign w4024 = w1974 & ~w2655;
assign w4025 = w2865 & w6674;
assign w4026 = w1976 & w2788;
assign w4027 = ~w4024 & ~w4025;
assign w4028 = ~w4026 & w4027;
assign w4029 = ~w4023 & w4028;
assign w4030 = ~w4021 & w4029;
assign w4031 = ~w565 & w4030;
assign w4032 = w565 & ~w4030;
assign w4033 = ~w4031 & ~w4032;
assign w4034 = ~w4019 & w4033;
assign w4035 = w4019 & ~w4033;
assign w4036 = ~w4034 & ~w4035;
assign w4037 = w2396 & ~w3348;
assign w4038 = (w2402 & w3171) | (w2402 & w6247) | (w3171 & w6247);
assign w4039 = (w2411 & w3146) | (w2411 & w6248) | (w3146 & w6248);
assign w4040 = w2901 & w6249;
assign w4041 = ~w4038 & ~w4039;
assign w4042 = (~w726 & ~w4041) | (~w726 & w6250) | (~w4041 & w6250);
assign w4043 = w4041 & w6251;
assign w4044 = ~w4042 & ~w4043;
assign w4045 = (w4044 & w3348) | (w4044 & w6252) | (w3348 & w6252);
assign w4046 = ~w4037 & ~w4045;
assign w4047 = w4036 & ~w4046;
assign w4048 = ~w4036 & w4046;
assign w4049 = ~w4047 & ~w4048;
assign w4050 = w3998 & ~w4049;
assign w4051 = ~w3998 & w4049;
assign w4052 = ~w4050 & ~w4051;
assign w4053 = ~w3472 & w6253;
assign w4054 = w2891 & ~w3164;
assign w4055 = ~w4053 & ~w4054;
assign w4056 = (w871 & ~w4055) | (w871 & w6254) | (~w4055 & w6254);
assign w4057 = w4055 & w6255;
assign w4058 = (w4057 & w3568) | (w4057 & w6675) | (w3568 & w6675);
assign w4059 = (~w4056 & w3568) | (~w4056 & w6256) | (w3568 & w6256);
assign w4060 = ~w4058 & w4059;
assign w4061 = w4052 & ~w4060;
assign w4062 = ~w4052 & w4060;
assign w4063 = ~w4061 & ~w4062;
assign w4064 = w3997 & w4063;
assign w4065 = ~w3997 & ~w4063;
assign w4066 = ~w4064 & ~w4065;
assign w4067 = ~w3780 & w3936;
assign w4068 = (~w3788 & w7531) | (~w3788 & w7297) | (w7531 & w7297);
assign w4069 = w3780 & ~w3936;
assign w4070 = (w4069 & w3788) | (w4069 & w7298) | (w3788 & w7298);
assign w4071 = ~w4068 & ~w4070;
assign w4072 = w3148 & ~w3936;
assign w4073 = (w0 & ~w3779) | (w0 & w6676) | (~w3779 & w6676);
assign w4074 = (~w2878 & w6965) | (~w2878 & w7770) | (w6965 & w7770);
assign w4075 = (w4071 & w6677) | (w4071 & w6678) | (w6677 & w6678);
assign w4076 = ~w4074 & ~w4075;
assign w4077 = ~w4066 & w4076;
assign w4078 = w3995 & w4077;
assign w4079 = w4066 & w4076;
assign w4080 = ~w3995 & w4079;
assign w4081 = ~w4078 & ~w4080;
assign w4082 = w4066 & ~w4076;
assign w4083 = w3995 & w4082;
assign w4084 = ~w4066 & ~w4076;
assign w4085 = ~w3995 & w4084;
assign w4086 = ~w4083 & ~w4085;
assign w4087 = w4081 & w4086;
assign w4088 = ~w237 & ~w270;
assign w4089 = w611 & w4088;
assign w4090 = w2825 & w4089;
assign w4091 = w531 & w3628;
assign w4092 = ~w164 & ~w226;
assign w4093 = ~w347 & w4092;
assign w4094 = w190 & w2739;
assign w4095 = w4093 & w4094;
assign w4096 = w208 & w1051;
assign w4097 = w4095 & w4096;
assign w4098 = w4090 & w4097;
assign w4099 = w946 & w4098;
assign w4100 = w4091 & w4099;
assign w4101 = ~w3988 & w3993;
assign w4102 = ~w3852 & ~w4101;
assign w4103 = w3852 & w4101;
assign w4104 = ~w4102 & ~w4103;
assign w4105 = w3947 & ~w4104;
assign w4106 = (w4100 & w4104) | (w4100 & w5762) | (w4104 & w5762);
assign w4107 = ~w4087 & w4106;
assign w4108 = ~w3987 & w4107;
assign w4109 = (~w4105 & ~w3837) | (~w4105 & w5763) | (~w3837 & w5763);
assign w4110 = w4087 & w4100;
assign w4111 = ~w4109 & w4110;
assign w4112 = ~w4108 & ~w4111;
assign w4113 = (~w4100 & w4104) | (~w4100 & w5764) | (w4104 & w5764);
assign w4114 = w4087 & w4113;
assign w4115 = ~w3987 & w4114;
assign w4116 = ~w4087 & ~w4100;
assign w4117 = ~w4109 & w4116;
assign w4118 = ~w4115 & ~w4117;
assign w4119 = w4112 & w4118;
assign w4120 = w3985 & ~w4119;
assign w4121 = ~w3985 & w4119;
assign w4122 = ~w4120 & ~w4121;
assign w4123 = ~w3967 & ~w4122;
assign w4124 = w3967 & w4122;
assign w4125 = ~w4123 & ~w4124;
assign w4126 = ~w3826 & ~w3969;
assign w4127 = w4125 & ~w6258;
assign w4128 = ~w4125 & w6258;
assign w4129 = ~w4127 & ~w4128;
assign w4130 = ~w4125 & w4126;
assign w4131 = (w3829 & w4125) | (w3829 & w6258) | (w4125 & w6258);
assign w4132 = ~w3976 & ~w4115;
assign w4133 = ~w4117 & w4132;
assign w4134 = w4112 & ~w4133;
assign w4135 = ~w3962 & ~w4108;
assign w4136 = ~w4111 & w4135;
assign w4137 = w3832 & w4136;
assign w4138 = ~w4134 & ~w4137;
assign w4139 = w4081 & ~w4105;
assign w4140 = w4086 & ~w4139;
assign w4141 = ~w3956 & w4086;
assign w4142 = w3837 & w4141;
assign w4143 = ~w4140 & ~w4142;
assign w4144 = w3995 & w4066;
assign w4145 = ~w4060 & ~w4066;
assign w4146 = ~w4144 & ~w4145;
assign w4147 = ~w3896 & ~w4034;
assign w4148 = ~w3900 & w4147;
assign w4149 = (~w4035 & w3900) | (~w4035 & w5637) | (w3900 & w5637);
assign w4150 = w1974 & w2788;
assign w4151 = w2865 & w6679;
assign w4152 = w2901 & w6259;
assign w4153 = ~w4150 & ~w4151;
assign w4154 = (w2874 & w6260) | (w2874 & w6261) | (w6260 & w6261);
assign w4155 = (~w2874 & w6262) | (~w2874 & w6263) | (w6262 & w6263);
assign w4156 = ~w4154 & ~w4155;
assign w4157 = w1022 & w4013;
assign w4158 = ~w4014 & ~w4157;
assign w4159 = (w1994 & w2656) | (w1994 & w6680) | (w2656 & w6680);
assign w4160 = ~w2583 & w6681;
assign w4161 = ~w2656 & w6682;
assign w4162 = (w4161 & w2583) | (w4161 & w6683) | (w2583 & w6683);
assign w4163 = ~w4160 & ~w4162;
assign w4164 = (~w1022 & w2244) | (~w1022 & w6264) | (w2244 & w6264);
assign w4165 = w1991 & ~w2410;
assign w4166 = w2241 & w2546;
assign w4167 = ~w4165 & ~w4166;
assign w4168 = (w4164 & ~w4167) | (w4164 & w6265) | (~w4167 & w6265);
assign w4169 = w4167 & w6266;
assign w4170 = ~w4168 & ~w4169;
assign w4171 = ~w4163 & ~w4170;
assign w4172 = w4163 & w4170;
assign w4173 = ~w4171 & ~w4172;
assign w4174 = w4158 & ~w4173;
assign w4175 = ~w4158 & w4173;
assign w4176 = ~w4174 & ~w4175;
assign w4177 = ~w4017 & w4176;
assign w4178 = w4017 & ~w4176;
assign w4179 = ~w4177 & ~w4178;
assign w4180 = w4156 & ~w4179;
assign w4181 = ~w4156 & w4179;
assign w4182 = ~w4180 & ~w4181;
assign w4183 = (w2405 & w3171) | (w2405 & w6267) | (w3171 & w6267);
assign w4184 = (w2402 & w3146) | (w2402 & w6268) | (w3146 & w6268);
assign w4185 = (w726 & ~w6269) | (w726 & w6684) | (~w6269 & w6684);
assign w4186 = w6269 & w7771;
assign w4187 = (~w4185 & ~w3203) | (~w4185 & w6686) | (~w3203 & w6686);
assign w4188 = ~w4186 & w4187;
assign w4189 = ~w4182 & w4188;
assign w4190 = w4149 & w4189;
assign w4191 = w4182 & w4188;
assign w4192 = ~w4149 & w4191;
assign w4193 = ~w4190 & ~w4192;
assign w4194 = w4182 & ~w4188;
assign w4195 = w4149 & w4194;
assign w4196 = ~w4182 & ~w4188;
assign w4197 = ~w4149 & w4196;
assign w4198 = ~w4195 & ~w4197;
assign w4199 = w4193 & w4198;
assign w4200 = (w2903 & ~w3779) | (w2903 & w6271) | (~w3779 & w6271);
assign w4201 = w2891 & ~w3474;
assign w4202 = (w3790 & w7299) | (w3790 & w7300) | (w7299 & w7300);
assign w4203 = ~w4201 & w7870;
assign w4204 = ~w4202 & ~w4203;
assign w4205 = w3173 & ~w3936;
assign w4206 = (w3780 & w3472) | (w3780 & w6273) | (w3472 & w6273);
assign w4207 = w3555 & ~w4206;
assign w4208 = w3175 & ~w3936;
assign w4209 = (w6096 & w7301) | (w6096 & w7302) | (w7301 & w7302);
assign w4210 = (w6096 & w7303) | (w6096 & w7304) | (w7303 & w7304);
assign w4211 = ~w4209 & w4210;
assign w4212 = ~w4204 & ~w4211;
assign w4213 = w4204 & w4211;
assign w4214 = ~w4212 & ~w4213;
assign w4215 = w4199 & w4214;
assign w4216 = ~w4199 & ~w4214;
assign w4217 = ~w4215 & ~w4216;
assign w4218 = (w5638 & w3861) | (w5638 & w6278) | (w3861 & w6278);
assign w4219 = ~w4047 & ~w4218;
assign w4220 = ~w4050 & ~w4219;
assign w4221 = (~w4220 & ~w3997) | (~w4220 & w6279) | (~w3997 & w6279);
assign w4222 = ~w4217 & w4221;
assign w4223 = w4217 & ~w4221;
assign w4224 = ~w4222 & ~w4223;
assign w4225 = (~w4224 & w4144) | (~w4224 & w6691) | (w4144 & w6691);
assign w4226 = ~w4145 & w4224;
assign w4227 = ~w4144 & w4226;
assign w4228 = ~w4225 & ~w4227;
assign w4229 = ~w4143 & w4228;
assign w4230 = w4143 & ~w4228;
assign w4231 = ~w4229 & ~w4230;
assign w4232 = ~w329 & ~w691;
assign w4233 = ~w109 & ~w204;
assign w4234 = ~w228 & ~w256;
assign w4235 = ~w402 & ~w528;
assign w4236 = w4234 & w4235;
assign w4237 = w4232 & w4233;
assign w4238 = w4236 & w4237;
assign w4239 = w680 & w3646;
assign w4240 = w3839 & w4239;
assign w4241 = w294 & w4238;
assign w4242 = w809 & w4241;
assign w4243 = w2294 & w4240;
assign w4244 = w4242 & w4243;
assign w4245 = w527 & w4244;
assign w4246 = w4231 & ~w4245;
assign w4247 = ~w4231 & w4245;
assign w4248 = ~w4246 & ~w4247;
assign w4249 = ~w4138 & w4248;
assign w4250 = w4138 & ~w4248;
assign w4251 = ~w4249 & ~w4250;
assign w4252 = w4124 & w4251;
assign w4253 = ~w4124 & ~w4251;
assign w4254 = ~w4252 & ~w4253;
assign w4255 = ~w4131 & w4254;
assign w4256 = w4131 & ~w4254;
assign w4257 = ~w4255 & ~w4256;
assign w4258 = w4138 & ~w4246;
assign w4259 = w4198 & ~w4220;
assign w4260 = w4193 & ~w4259;
assign w4261 = ~w4052 & w4193;
assign w4262 = w3997 & w4261;
assign w4263 = ~w4260 & ~w4262;
assign w4264 = ~w2244 & w6280;
assign w4265 = w4167 & w6281;
assign w4266 = w4163 & w4265;
assign w4267 = w4016 & ~w4266;
assign w4268 = ~w4005 & w4267;
assign w4269 = (w1994 & ~w2656) | (w1994 & w6692) | (~w2656 & w6692);
assign w4270 = (w4269 & w2385) | (w4269 & w6693) | (w2385 & w6693);
assign w4271 = ~w2925 & w4270;
assign w4272 = ~w2410 & w2546;
assign w4273 = w1991 & ~w2655;
assign w4274 = w1987 & w2788;
assign w4275 = ~w4272 & ~w4273;
assign w4276 = ~w4274 & w4275;
assign w4277 = (~w2878 & w2241) | (~w2878 & w6282) | (w2241 & w6282);
assign w4278 = ~w2241 & w6283;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = (~w2925 & w6694) | (~w2925 & w6695) | (w6694 & w6695);
assign w4281 = (w5766 & w2925) | (w5766 & w6696) | (w2925 & w6696);
assign w4282 = ~w4280 & ~w4281;
assign w4283 = ~w4268 & w5640;
assign w4284 = (w4282 & w4268) | (w4282 & w5641) | (w4268 & w5641);
assign w4285 = ~w4283 & ~w4284;
assign w4286 = (w1968 & w3171) | (w1968 & w6284) | (w3171 & w6284);
assign w4287 = w2865 & w6697;
assign w4288 = w2901 & w6285;
assign w4289 = ~w4286 & ~w4287;
assign w4290 = ~w4286 & w7305;
assign w4291 = (w2803 & w6286) | (w2803 & w6287) | (w6286 & w6287);
assign w4292 = ~w3361 & w4291;
assign w4293 = ~w4292 & w6288;
assign w4294 = (w565 & w4292) | (w565 & w6289) | (w4292 & w6289);
assign w4295 = ~w4293 & ~w4294;
assign w4296 = w4285 & ~w4295;
assign w4297 = ~w4285 & w4295;
assign w4298 = ~w4296 & ~w4297;
assign w4299 = w2396 & w3483;
assign w4300 = (w2405 & w3146) | (w2405 & w6290) | (w3146 & w6290);
assign w4301 = w2402 & ~w3164;
assign w4302 = ~w4300 & ~w4301;
assign w4303 = (~w726 & ~w4302) | (~w726 & w6291) | (~w4302 & w6291);
assign w4304 = w4302 & w6292;
assign w4305 = ~w4303 & ~w4304;
assign w4306 = (w4305 & ~w3483) | (w4305 & w6293) | (~w3483 & w6293);
assign w4307 = ~w4299 & ~w4306;
assign w4308 = w4298 & w4307;
assign w4309 = ~w4298 & ~w4307;
assign w4310 = ~w4308 & ~w4309;
assign w4311 = (~w4035 & ~w4179) | (~w4035 & w5642) | (~w4179 & w5642);
assign w4312 = (~w4180 & w4148) | (~w4180 & w5643) | (w4148 & w5643);
assign w4313 = ~w4067 & ~w4069;
assign w4314 = w3009 & ~w4313;
assign w4315 = w2903 & ~w3936;
assign w4316 = (w2893 & ~w3779) | (w2893 & w6295) | (~w3779 & w6295);
assign w4317 = ~w4315 & ~w4316;
assign w4318 = (w4317 & w3472) | (w4317 & w6297) | (w3472 & w6297);
assign w4319 = (w6698 & w6699) | (w6698 & w7871) | (w6699 & w7871);
assign w4320 = (~w871 & ~w4319) | (~w871 & w6298) | (~w4319 & w6298);
assign w4321 = w4319 & w6299;
assign w4322 = ~w4320 & ~w4321;
assign w4323 = w4312 & ~w4322;
assign w4324 = ~w4312 & w4322;
assign w4325 = ~w4323 & ~w4324;
assign w4326 = w4310 & w4325;
assign w4327 = ~w4310 & ~w4325;
assign w4328 = ~w4326 & ~w4327;
assign w4329 = w4263 & w4328;
assign w4330 = ~w4263 & ~w4328;
assign w4331 = ~w4329 & ~w4330;
assign w4332 = (~w4212 & ~w4199) | (~w4212 & w5644) | (~w4199 & w5644);
assign w4333 = w4221 & ~w4332;
assign w4334 = (~w4213 & ~w4199) | (~w4213 & w5645) | (~w4199 & w5645);
assign w4335 = ~w4221 & w4334;
assign w4336 = ~w4333 & ~w4335;
assign w4337 = w4331 & w4336;
assign w4338 = ~w4331 & ~w4336;
assign w4339 = ~w4337 & ~w4338;
assign w4340 = ~w160 & ~w211;
assign w4341 = w530 & w4340;
assign w4342 = w543 & w676;
assign w4343 = w2825 & w4342;
assign w4344 = w2165 & w4341;
assign w4345 = w4343 & w4344;
assign w4346 = w766 & w4345;
assign w4347 = w802 & w4346;
assign w4348 = w1519 & w4347;
assign w4349 = w4339 & ~w4348;
assign w4350 = ~w4339 & w4348;
assign w4351 = ~w4349 & ~w4350;
assign w4352 = w4227 & w4351;
assign w4353 = ~w4225 & w4351;
assign w4354 = w4143 & w4353;
assign w4355 = ~w4352 & ~w4354;
assign w4356 = w4143 & ~w4225;
assign w4357 = ~w4227 & ~w4351;
assign w4358 = ~w4356 & w4357;
assign w4359 = w4355 & ~w4358;
assign w4360 = ~w4247 & w4359;
assign w4361 = ~w4258 & w4360;
assign w4362 = ~w4138 & ~w4247;
assign w4363 = ~w4246 & ~w4359;
assign w4364 = ~w4362 & w4363;
assign w4365 = ~w4361 & ~w4364;
assign w4366 = ~w4252 & w4365;
assign w4367 = w4252 & ~w4365;
assign w4368 = ~w4366 & ~w4367;
assign w4369 = w4130 & ~w4254;
assign w4370 = (w3829 & w4254) | (w3829 & w6700) | (w4254 & w6700);
assign w4371 = w4368 & ~w4370;
assign w4372 = ~w4368 & w4370;
assign w4373 = ~w4371 & ~w4372;
assign w4374 = ~w4227 & w4339;
assign w4375 = ~w4348 & ~w4374;
assign w4376 = (~w4348 & w4146) | (~w4348 & w6300) | (w4146 & w6300);
assign w4377 = (~w4375 & ~w4143) | (~w4375 & w6701) | (~w4143 & w6701);
assign w4378 = w4355 & w5646;
assign w4379 = ~w4225 & w4374;
assign w4380 = w4143 & w4379;
assign w4381 = ~w4337 & ~w4374;
assign w4382 = (w2891 & ~w3779) | (w2891 & w6301) | (~w3779 & w6301);
assign w4383 = w2893 & ~w3936;
assign w4384 = (~w871 & w4383) | (~w871 & w6302) | (w4383 & w6302);
assign w4385 = ~w4383 & w6303;
assign w4386 = (w4385 & w4071) | (w4385 & w6702) | (w4071 & w6702);
assign w4387 = (~w4384 & w4071) | (~w4384 & w6304) | (w4071 & w6304);
assign w4388 = ~w4386 & w4387;
assign w4389 = ~w4309 & ~w4312;
assign w4390 = (w4388 & w4389) | (w4388 & w5767) | (w4389 & w5767);
assign w4391 = ~w4389 & w5768;
assign w4392 = ~w4390 & ~w4391;
assign w4393 = (~w4283 & ~w4285) | (~w4283 & w5769) | (~w4285 & w5769);
assign w4394 = w2402 & ~w3474;
assign w4395 = w2405 & ~w3164;
assign w4396 = ~w4394 & ~w4395;
assign w4397 = (w726 & ~w4396) | (w726 & w7772) | (~w4396 & w7772);
assign w4398 = (w3568 & w6305) | (w3568 & w6306) | (w6305 & w6306);
assign w4399 = ~w4397 & ~w4398;
assign w4400 = ~w4393 & w4399;
assign w4401 = w4393 & ~w4399;
assign w4402 = ~w4400 & ~w4401;
assign w4403 = (w2878 & w2410) | (w2878 & w6307) | (w2410 & w6307);
assign w4404 = ~w2410 & w6308;
assign w4405 = ~w4403 & ~w4404;
assign w4406 = (~w2925 & w6703) | (~w2925 & w6704) | (w6703 & w6704);
assign w4407 = (~w1022 & w2241) | (~w1022 & w6309) | (w2241 & w6309);
assign w4408 = (w5771 & w2925) | (w5771 & w6705) | (w2925 & w6705);
assign w4409 = ~w4406 & ~w4408;
assign w4410 = ~w4405 & ~w4409;
assign w4411 = ~w4403 & w4407;
assign w4412 = (w6310 & w2925) | (w6310 & w6706) | (w2925 & w6706);
assign w4413 = (w2925 & w7306) | (w2925 & w7307) | (w7306 & w7307);
assign w4414 = ~w4412 & w4413;
assign w4415 = ~w4410 & ~w4414;
assign w4416 = w2546 & ~w2655;
assign w4417 = w2865 & w6707;
assign w4418 = ~w4416 & ~w4417;
assign w4419 = (w1022 & ~w4418) | (w1022 & w6312) | (~w4418 & w6312);
assign w4420 = w4418 & w6313;
assign w4421 = ~w4419 & ~w4420;
assign w4422 = (w4421 & ~w3078) | (w4421 & w6314) | (~w3078 & w6314);
assign w4423 = w3078 & w5775;
assign w4424 = ~w4422 & ~w4423;
assign w4425 = ~w4415 & ~w4424;
assign w4426 = w4415 & w4424;
assign w4427 = ~w4425 & ~w4426;
assign w4428 = w2563 & ~w3348;
assign w4429 = ~w1959 & w1961;
assign w4430 = (w1976 & w3171) | (w1976 & w6315) | (w3171 & w6315);
assign w4431 = (w1968 & w3146) | (w1968 & w6316) | (w3146 & w6316);
assign w4432 = w2901 & w6317;
assign w4433 = ~w4430 & ~w4431;
assign w4434 = (~w565 & ~w4433) | (~w565 & w6318) | (~w4433 & w6318);
assign w4435 = w4433 & w6319;
assign w4436 = ~w4434 & ~w4435;
assign w4437 = (w4436 & w3348) | (w4436 & w6320) | (w3348 & w6320);
assign w4438 = ~w4428 & ~w4437;
assign w4439 = ~w4427 & w4438;
assign w4440 = w4427 & ~w4438;
assign w4441 = ~w4439 & ~w4440;
assign w4442 = w4402 & ~w4441;
assign w4443 = ~w4402 & w4441;
assign w4444 = ~w4442 & ~w4443;
assign w4445 = w4392 & w4444;
assign w4446 = ~w4392 & ~w4444;
assign w4447 = ~w4445 & ~w4446;
assign w4448 = w4322 & ~w4328;
assign w4449 = (w4447 & w4329) | (w4447 & w5772) | (w4329 & w5772);
assign w4450 = ~w4329 & w5773;
assign w4451 = ~w4449 & ~w4450;
assign w4452 = w539 & w2164;
assign w4453 = ~w109 & w1670;
assign w4454 = ~w314 & ~w486;
assign w4455 = w930 & w4454;
assign w4456 = w934 & w4455;
assign w4457 = w3463 & w3838;
assign w4458 = w4452 & w4453;
assign w4459 = w4457 & w4458;
assign w4460 = w2185 & w4456;
assign w4461 = w4459 & w4460;
assign w4462 = w3131 & w4461;
assign w4463 = w3926 & w4462;
assign w4464 = ~w4451 & w4463;
assign w4465 = w4451 & ~w4463;
assign w4466 = ~w4464 & ~w4465;
assign w4467 = ~w4381 & ~w4466;
assign w4468 = w4381 & w4466;
assign w4469 = ~w4467 & ~w4468;
assign w4470 = ~w4380 & ~w4469;
assign w4471 = w4143 & w6708;
assign w4472 = ~w4470 & ~w4471;
assign w4473 = ~w4378 & ~w4472;
assign w4474 = w4355 & ~w4377;
assign w4475 = ~w4246 & ~w4474;
assign w4476 = ~w4362 & w4475;
assign w4477 = w4473 & ~w4476;
assign w4478 = w4378 & w4472;
assign w4479 = w4472 & w4475;
assign w4480 = (~w4478 & ~w4479) | (~w4478 & w5647) | (~w4479 & w5647);
assign w4481 = ~w4477 & w4480;
assign w4482 = ~w4367 & ~w4481;
assign w4483 = w4367 & w4481;
assign w4484 = ~w4482 & ~w4483;
assign w4485 = ~w4368 & w4369;
assign w4486 = w3829 & ~w4485;
assign w4487 = ~w4484 & w4486;
assign w4488 = w4484 & ~w4486;
assign w4489 = ~w4487 & ~w4488;
assign w4490 = ~w4470 & w5648;
assign w4491 = (~w4490 & w4378) | (~w4490 & w6709) | (w4378 & w6709);
assign w4492 = w4475 & ~w4490;
assign w4493 = ~w4249 & w4492;
assign w4494 = ~w4337 & ~w4449;
assign w4495 = ~w4225 & w4494;
assign w4496 = w4143 & w4495;
assign w4497 = ~w273 & ~w347;
assign w4498 = w349 & w4497;
assign w4499 = w370 & w2164;
assign w4500 = w2174 & w4499;
assign w4501 = w1512 & w4498;
assign w4502 = w1674 & w3928;
assign w4503 = w4501 & w4502;
assign w4504 = w4500 & w4503;
assign w4505 = ~w119 & ~w935;
assign w4506 = ~w206 & w4505;
assign w4507 = ~w163 & ~w178;
assign w4508 = ~w200 & ~w238;
assign w4509 = w4507 & w4508;
assign w4510 = w2182 & w2620;
assign w4511 = w4509 & w4510;
assign w4512 = w4506 & w4511;
assign w4513 = w1510 & w4512;
assign w4514 = w4504 & w4513;
assign w4515 = w3614 & w4514;
assign w4516 = ~w4374 & w4494;
assign w4517 = (~w4390 & ~w4392) | (~w4390 & w6321) | (~w4392 & w6321);
assign w4518 = (w6096 & w7308) | (w6096 & w7309) | (w7308 & w7309);
assign w4519 = (~w871 & w6325) | (~w871 & w7872) | (w6325 & w7872);
assign w4520 = ~w4518 & ~w4519;
assign w4521 = ~w4401 & ~w4441;
assign w4522 = (~w4520 & w4521) | (~w4520 & w6326) | (w4521 & w6326);
assign w4523 = ~w4521 & w6327;
assign w4524 = ~w4522 & ~w4523;
assign w4525 = (w2878 & w2655) | (w2878 & w6307) | (w2655 & w6307);
assign w4526 = ~w2655 & w6308;
assign w4527 = ~w4525 & ~w4526;
assign w4528 = ~w4277 & ~w4404;
assign w4529 = ~w4527 & ~w4528;
assign w4530 = w4527 & w4528;
assign w4531 = ~w4529 & ~w4530;
assign w4532 = (w4531 & w4271) | (w4531 & w6328) | (w4271 & w6328);
assign w4533 = ~w4411 & w4527;
assign w4534 = w4411 & ~w4527;
assign w4535 = ~w4533 & ~w4534;
assign w4536 = ~w4271 & w6329;
assign w4537 = ~w4532 & ~w4536;
assign w4538 = w2546 & w2788;
assign w4539 = w2865 & w6712;
assign w4540 = w2901 & w6330;
assign w4541 = ~w4538 & ~w4539;
assign w4542 = (w1022 & ~w4541) | (w1022 & w6331) | (~w4541 & w6331);
assign w4543 = w4541 & w6332;
assign w4544 = ~w4542 & ~w4543;
assign w4545 = (w4544 & w2874) | (w4544 & w5774) | (w2874 & w5774);
assign w4546 = ~w2874 & w5775;
assign w4547 = ~w4545 & ~w4546;
assign w4548 = ~w4537 & ~w4547;
assign w4549 = w4537 & w4547;
assign w4550 = ~w4548 & ~w4549;
assign w4551 = w2563 & w3203;
assign w4552 = (w1976 & w3146) | (w1976 & w6333) | (w3146 & w6333);
assign w4553 = (w1974 & w3171) | (w1974 & w6334) | (w3171 & w6334);
assign w4554 = ~w4552 & ~w4553;
assign w4555 = (~w565 & ~w4554) | (~w565 & w6713) | (~w4554 & w6713);
assign w4556 = w4554 & w6714;
assign w4557 = ~w4555 & ~w4556;
assign w4558 = (w4557 & ~w3203) | (w4557 & w6335) | (~w3203 & w6335);
assign w4559 = ~w4551 & ~w4558;
assign w4560 = w4550 & ~w4559;
assign w4561 = ~w4550 & w4559;
assign w4562 = ~w4560 & ~w4561;
assign w4563 = ~w4426 & ~w4438;
assign w4564 = ~w4425 & ~w4563;
assign w4565 = ~w4562 & w4564;
assign w4566 = w4562 & ~w4564;
assign w4567 = ~w4565 & ~w4566;
assign w4568 = (w2411 & ~w3779) | (w2411 & w6337) | (~w3779 & w6337);
assign w4569 = w2405 & ~w3474;
assign w4570 = (w3790 & w7310) | (w3790 & w7311) | (w7310 & w7311);
assign w4571 = ~w4569 & w7873;
assign w4572 = ~w4570 & ~w4571;
assign w4573 = ~w4567 & w4572;
assign w4574 = w4567 & ~w4572;
assign w4575 = ~w4573 & ~w4574;
assign w4576 = ~w4524 & w4575;
assign w4577 = w4524 & ~w4575;
assign w4578 = ~w4576 & ~w4577;
assign w4579 = ~w4517 & w4578;
assign w4580 = w4517 & ~w4578;
assign w4581 = ~w4579 & ~w4580;
assign w4582 = ~w4450 & w4581;
assign w4583 = (w4582 & w4374) | (w4582 & w5649) | (w4374 & w5649);
assign w4584 = w4515 & w4583;
assign w4585 = ~w4496 & w4584;
assign w4586 = w4515 & ~w4581;
assign w4587 = (~w4374 & w5832) | (~w4374 & w5833) | (w5832 & w5833);
assign w4588 = w4495 & w4586;
assign w4589 = (~w4587 & ~w4143) | (~w4587 & w7262) | (~w4143 & w7262);
assign w4590 = ~w4585 & w4589;
assign w4591 = (w4143 & w7263) | (w4143 & w7264) | (w7263 & w7264);
assign w4592 = (~w4515 & w4496) | (~w4515 & w5777) | (w4496 & w5777);
assign w4593 = ~w4591 & w4592;
assign w4594 = w4590 & ~w4593;
assign w4595 = (w4594 & w4493) | (w4594 & w5651) | (w4493 & w5651);
assign w4596 = ~w4493 & w5652;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = ~w4483 & w4597;
assign w4599 = w4483 & ~w4597;
assign w4600 = ~w4598 & ~w4599;
assign w4601 = ~w4484 & w4485;
assign w4602 = w3829 & ~w4601;
assign w4603 = w4600 & ~w4602;
assign w4604 = ~w4600 & w4602;
assign w4605 = ~w4603 & ~w4604;
assign w4606 = (~w4572 & w4562) | (~w4572 & w6715) | (w4562 & w6715);
assign w4607 = w2396 & w3942;
assign w4608 = w2411 & ~w3936;
assign w4609 = (w2402 & ~w3779) | (w2402 & w6339) | (~w3779 & w6339);
assign w4610 = (~w3472 & w6716) | (~w3472 & w6717) | (w6716 & w6717);
assign w4611 = (w3472 & w6342) | (w3472 & w6343) | (w6342 & w6343);
assign w4612 = ~w4610 & ~w4611;
assign w4613 = (w4612 & ~w3942) | (w4612 & w6344) | (~w3942 & w6344);
assign w4614 = ~w4607 & ~w4613;
assign w4615 = (w4614 & ~w4562) | (w4614 & w6718) | (~w4562 & w6718);
assign w4616 = ~w4606 & w4615;
assign w4617 = (w4572 & ~w4562) | (w4572 & w6719) | (~w4562 & w6719);
assign w4618 = (~w4614 & w4562) | (~w4614 & w6720) | (w4562 & w6720);
assign w4619 = ~w4617 & w4618;
assign w4620 = ~w4616 & ~w4619;
assign w4621 = (~w4548 & ~w4550) | (~w4548 & w6345) | (~w4550 & w6345);
assign w4622 = (w1987 & w3171) | (w1987 & w6346) | (w3171 & w6346);
assign w4623 = w2865 & w6721;
assign w4624 = w2901 & w6347;
assign w4625 = ~w4622 & ~w4623;
assign w4626 = ~w4622 & w7312;
assign w4627 = w4625 & w6348;
assign w4628 = (w2803 & w6349) | (w2803 & w6350) | (w6349 & w6350);
assign w4629 = ~w3361 & w4628;
assign w4630 = ~w871 & ~w2878;
assign w4631 = w871 & w2878;
assign w4632 = ~w4630 & ~w4631;
assign w4633 = w2788 & w4632;
assign w4634 = (~w1022 & w2788) | (~w1022 & w6351) | (w2788 & w6351);
assign w4635 = ~w4633 & w4634;
assign w4636 = w1022 & ~w4632;
assign w4637 = ~w4635 & ~w4636;
assign w4638 = ~w4629 & w6352;
assign w4639 = (w4637 & w4629) | (w4637 & w6353) | (w4629 & w6353);
assign w4640 = ~w4638 & ~w4639;
assign w4641 = (~w4525 & ~w4537) | (~w4525 & w6354) | (~w4537 & w6354);
assign w4642 = ~w4640 & w4641;
assign w4643 = w4640 & ~w4641;
assign w4644 = ~w4642 & ~w4643;
assign w4645 = w2563 & w3483;
assign w4646 = w1976 & ~w3164;
assign w4647 = (w1974 & w3146) | (w1974 & w6355) | (w3146 & w6355);
assign w4648 = ~w4646 & ~w4647;
assign w4649 = (~w565 & ~w4648) | (~w565 & w6356) | (~w4648 & w6356);
assign w4650 = w4648 & w6357;
assign w4651 = ~w4649 & ~w4650;
assign w4652 = (w4651 & ~w3483) | (w4651 & w6358) | (~w3483 & w6358);
assign w4653 = ~w4645 & ~w4652;
assign w4654 = ~w4644 & ~w4653;
assign w4655 = w4644 & w4653;
assign w4656 = ~w4654 & ~w4655;
assign w4657 = ~w4621 & w4656;
assign w4658 = w4621 & ~w4656;
assign w4659 = ~w4657 & ~w4658;
assign w4660 = w4620 & ~w4659;
assign w4661 = ~w4620 & w4659;
assign w4662 = ~w4660 & ~w4661;
assign w4663 = (~w4523 & ~w4575) | (~w4523 & w6359) | (~w4575 & w6359);
assign w4664 = w4662 & w4663;
assign w4665 = ~w4662 & ~w4663;
assign w4666 = ~w4664 & ~w4665;
assign w4667 = ~w4579 & ~w4666;
assign w4668 = ~w4583 & w4667;
assign w4669 = w4495 & w4667;
assign w4670 = w4143 & w4669;
assign w4671 = ~w4668 & ~w4670;
assign w4672 = w4579 & w4666;
assign w4673 = ~w4450 & w5653;
assign w4674 = (w4673 & w4374) | (w4673 & w5778) | (w4374 & w5778);
assign w4675 = (~w4374 & w5779) | (~w4374 & w5780) | (w5779 & w5780);
assign w4676 = w4495 & ~w4672;
assign w4677 = (~w4675 & ~w4143) | (~w4675 & w7265) | (~w4143 & w7265);
assign w4678 = ~w160 & ~w366;
assign w4679 = w335 & w657;
assign w4680 = w814 & w3150;
assign w4681 = w3655 & w4678;
assign w4682 = w4680 & w4681;
assign w4683 = w4453 & w4679;
assign w4684 = w4682 & w4683;
assign w4685 = w4504 & w4684;
assign w4686 = w2313 & w4685;
assign w4687 = (w4686 & ~w4671) | (w4686 & w7266) | (~w4671 & w7266);
assign w4688 = (~w4686 & ~w4666) | (~w4686 & w6360) | (~w4666 & w6360);
assign w4689 = (~w4374 & w5781) | (~w4374 & w5782) | (w5781 & w5782);
assign w4690 = w4495 & w4688;
assign w4691 = (~w4689 & ~w4143) | (~w4689 & w7267) | (~w4143 & w7267);
assign w4692 = w4671 & ~w4691;
assign w4693 = ~w4687 & ~w4692;
assign w4694 = w4594 & w4693;
assign w4695 = (w4694 & w4493) | (w4694 & w5654) | (w4493 & w5654);
assign w4696 = w4590 & ~w4692;
assign w4697 = ~w4687 & w4696;
assign w4698 = (~w4590 & w4687) | (~w4590 & w6361) | (w4687 & w6361);
assign w4699 = ~w4697 & ~w4698;
assign w4700 = w4699 & ~w4595;
assign w4701 = ~w4695 & ~w4700;
assign w4702 = w4599 & ~w4701;
assign w4703 = ~w4599 & w4701;
assign w4704 = ~w4702 & ~w4703;
assign w4705 = ~w4600 & w4601;
assign w4706 = w3829 & ~w4705;
assign w4707 = w4704 & ~w4706;
assign w4708 = ~w4704 & w4706;
assign w4709 = ~w4707 & ~w4708;
assign w4710 = ~w4704 & w4705;
assign w4711 = (~w4664 & ~w4666) | (~w4664 & w6362) | (~w4666 & w6362);
assign w4712 = (~w4374 & w5783) | (~w4374 & w5784) | (w5783 & w5784);
assign w4713 = w4495 & w4711;
assign w4714 = w4143 & w4713;
assign w4715 = (~w4616 & ~w4620) | (~w4616 & w6363) | (~w4620 & w6363);
assign w4716 = w2563 & ~w3568;
assign w4717 = ~w3472 & w6364;
assign w4718 = w1974 & ~w3164;
assign w4719 = ~w4717 & ~w4718;
assign w4720 = (~w565 & ~w4719) | (~w565 & w6365) | (~w4719 & w6365);
assign w4721 = w4719 & w6366;
assign w4722 = ~w4720 & ~w4721;
assign w4723 = (w4722 & w3568) | (w4722 & w6367) | (w3568 & w6367);
assign w4724 = ~w4716 & ~w4723;
assign w4725 = (~w1022 & ~w2865) | (~w1022 & w6722) | (~w2865 & w6722);
assign w4726 = (~w4631 & ~w2788) | (~w4631 & w6368) | (~w2788 & w6368);
assign w4727 = w4725 & ~w4726;
assign w4728 = ~w4725 & w4726;
assign w4729 = ~w4727 & ~w4728;
assign w4730 = (w1987 & w3146) | (w1987 & w6369) | (w3146 & w6369);
assign w4731 = (w1991 & w3171) | (w1991 & w6370) | (w3171 & w6370);
assign w4732 = w2901 & w6371;
assign w4733 = ~w4730 & ~w4731;
assign w4734 = ~w4732 & w4733;
assign w4735 = w4729 & w7773;
assign w4736 = (w3348 & w6373) | (w3348 & w6374) | (w6373 & w6374);
assign w4737 = ~w4735 & ~w4736;
assign w4738 = ~w4724 & w4737;
assign w4739 = w4724 & ~w4737;
assign w4740 = ~w4738 & ~w4739;
assign w4741 = w1022 & w4632;
assign w4742 = ~w4629 & w6375;
assign w4743 = (w4635 & w4629) | (w4635 & w6376) | (w4629 & w6376);
assign w4744 = ~w4742 & ~w4743;
assign w4745 = ~w4642 & w4744;
assign w4746 = w4740 & w4745;
assign w4747 = ~w4740 & ~w4745;
assign w4748 = ~w4746 & ~w4747;
assign w4749 = w2402 & ~w3936;
assign w4750 = (w2405 & ~w3779) | (w2405 & w6377) | (~w3779 & w6377);
assign w4751 = (w4071 & w6723) | (w4071 & w6724) | (w6723 & w6724);
assign w4752 = (~w4071 & w6379) | (~w4071 & w6380) | (w6379 & w6380);
assign w4753 = ~w4751 & ~w4752;
assign w4754 = w4748 & ~w4753;
assign w4755 = ~w4748 & w4753;
assign w4756 = ~w4754 & ~w4755;
assign w4757 = (~w4654 & ~w4656) | (~w4654 & w6381) | (~w4656 & w6381);
assign w4758 = w4756 & w4757;
assign w4759 = ~w4756 & ~w4757;
assign w4760 = ~w4758 & ~w4759;
assign w4761 = ~w4715 & w4760;
assign w4762 = w4715 & ~w4760;
assign w4763 = ~w4761 & ~w4762;
assign w4764 = ~w303 & ~w402;
assign w4765 = w120 & w4764;
assign w4766 = w212 & w805;
assign w4767 = w2299 & w4766;
assign w4768 = w1561 & w4765;
assign w4769 = w4767 & w4768;
assign w4770 = w361 & w4769;
assign w4771 = ~w147 & ~w183;
assign w4772 = w1520 & w4771;
assign w4773 = w1557 & w3545;
assign w4774 = w4232 & w4773;
assign w4775 = w771 & w4772;
assign w4776 = w4774 & w4775;
assign w4777 = w760 & w4776;
assign w4778 = w4770 & w4777;
assign w4779 = w3662 & w4778;
assign w4780 = ~w4763 & ~w4779;
assign w4781 = ~w4714 & w5785;
assign w4782 = w4763 & ~w4779;
assign w4783 = (w4782 & w4714) | (w4782 & w5786) | (w4714 & w5786);
assign w4784 = ~w4781 & ~w4783;
assign w4785 = w4763 & w4779;
assign w4786 = ~w4714 & w5787;
assign w4787 = ~w4763 & w4779;
assign w4788 = (w4787 & w4714) | (w4787 & w5788) | (w4714 & w5788);
assign w4789 = ~w4786 & ~w4788;
assign w4790 = w4784 & w4789;
assign w4791 = (w4790 & w4697) | (w4790 & w5789) | (w4697 & w5789);
assign w4792 = ~w4697 & w5790;
assign w4793 = ~w4791 & ~w4792;
assign w4794 = w4695 & w4793;
assign w4795 = ~w4695 & ~w4793;
assign w4796 = ~w4794 & ~w4795;
assign w4797 = w4599 & w7268;
assign w4798 = (~w4796 & ~w4599) | (~w4796 & w7269) | (~w4599 & w7269);
assign w4799 = ~w4797 & ~w4798;
assign w4800 = ~w4710 & w7313;
assign w4801 = (w4799 & w4710) | (w4799 & w7314) | (w4710 & w7314);
assign w4802 = ~w4800 & ~w4801;
assign w4803 = ~w4692 & w4784;
assign w4804 = ~w4490 & ~w4593;
assign w4805 = w4803 & w4804;
assign w4806 = (w4805 & w4476) | (w4805 & w6725) | (w4476 & w6725);
assign w4807 = ~w4697 & w4803;
assign w4808 = ~w4664 & ~w4761;
assign w4809 = (~w4762 & w4672) | (~w4762 & w6382) | (w4672 & w6382);
assign w4810 = ~w4450 & w6726;
assign w4811 = w4495 & ~w4809;
assign w4812 = w4143 & w4811;
assign w4813 = (~w4738 & ~w4740) | (~w4738 & w6383) | (~w4740 & w6383);
assign w4814 = (w6096 & w7315) | (w6096 & w7316) | (w7315 & w7316);
assign w4815 = (w726 & w6387) | (w726 & w7874) | (w6387 & w7874);
assign w4816 = ~w4814 & ~w4815;
assign w4817 = w4813 & ~w4816;
assign w4818 = ~w4813 & w4816;
assign w4819 = ~w4817 & ~w4818;
assign w4820 = ~w1022 & w2860;
assign w4821 = w1987 & ~w3164;
assign w4822 = (w2546 & w3171) | (w2546 & w6388) | (w3171 & w6388);
assign w4823 = (w1991 & w3146) | (w1991 & w6389) | (w3146 & w6389);
assign w4824 = ~w4821 & w6390;
assign w4825 = w4824 & w7774;
assign w4826 = (w3203 & w6729) | (w3203 & w6730) | (w6729 & w6730);
assign w4827 = ~w4825 & ~w4826;
assign w4828 = (w3348 & w6391) | (w3348 & w6392) | (w6391 & w6392);
assign w4829 = ~w1022 & ~w4727;
assign w4830 = ~w4829 & w7773;
assign w4831 = ~w4828 & ~w4830;
assign w4832 = w4827 & w4831;
assign w4833 = ~w4827 & ~w4831;
assign w4834 = ~w4832 & ~w4833;
assign w4835 = (w1968 & ~w3779) | (w1968 & w6394) | (~w3779 & w6394);
assign w4836 = w1974 & ~w3474;
assign w4837 = (w3790 & w7317) | (w3790 & w7318) | (w7317 & w7318);
assign w4838 = ~w4836 & w7875;
assign w4839 = ~w4837 & ~w4838;
assign w4840 = w4834 & ~w4839;
assign w4841 = ~w4834 & w4839;
assign w4842 = ~w4840 & ~w4841;
assign w4843 = w4819 & ~w4842;
assign w4844 = ~w4819 & w4842;
assign w4845 = ~w4843 & ~w4844;
assign w4846 = (~w4755 & ~w4756) | (~w4755 & w6396) | (~w4756 & w6396);
assign w4847 = w4845 & ~w4846;
assign w4848 = ~w4845 & w4846;
assign w4849 = ~w4847 & ~w4848;
assign w4850 = ~w106 & ~w356;
assign w4851 = ~w538 & w4850;
assign w4852 = w2175 & w2818;
assign w4853 = w3150 & w4852;
assign w4854 = w3117 & w4851;
assign w4855 = w4506 & w4854;
assign w4856 = w820 & w4853;
assign w4857 = w4855 & w4856;
assign w4858 = w1683 & w4857;
assign w4859 = w3601 & w4858;
assign w4860 = w4849 & ~w4859;
assign w4861 = ~w4849 & w4859;
assign w4862 = ~w4860 & ~w4861;
assign w4863 = ~w4812 & w6731;
assign w4864 = (~w4862 & w4812) | (~w4862 & w6732) | (w4812 & w6732);
assign w4865 = ~w4863 & ~w4864;
assign w4866 = w4789 & w4865;
assign w4867 = (w4866 & w4697) | (w4866 & w6733) | (w4697 & w6733);
assign w4868 = ~w4806 & w4867;
assign w4869 = (w4789 & w4697) | (w4789 & w5791) | (w4697 & w5791);
assign w4870 = ~w4865 & ~w4869;
assign w4871 = w4804 & w5792;
assign w4872 = ~w4477 & w4871;
assign w4873 = ~w4870 & ~w4872;
assign w4874 = ~w4868 & w4873;
assign w4875 = w4796 & w4874;
assign w4876 = w4702 & w4875;
assign w4877 = (~w4874 & ~w4702) | (~w4874 & w5793) | (~w4702 & w5793);
assign w4878 = ~w4876 & ~w4877;
assign w4879 = w4710 & ~w4799;
assign w4880 = ~w4879 & w6397;
assign w4881 = (w4878 & w4879) | (w4878 & w6398) | (w4879 & w6398);
assign w4882 = ~w4880 & ~w4881;
assign w4883 = ~w4672 & w6399;
assign w4884 = w4495 & w4883;
assign w4885 = w4143 & w4884;
assign w4886 = (~w1022 & w3171) | (~w1022 & w6400) | (w3171 & w6400);
assign w4887 = w726 & ~w4886;
assign w4888 = ~w1022 & w7775;
assign w4889 = ~w4887 & ~w4888;
assign w4890 = w2865 & w6734;
assign w4891 = w4889 & ~w4890;
assign w4892 = ~w4889 & w4890;
assign w4893 = ~w4891 & ~w4892;
assign w4894 = w2902 & w4725;
assign w4895 = w4893 & ~w4894;
assign w4896 = ~w4827 & w4895;
assign w4897 = w4889 & w4894;
assign w4898 = ~w1022 & ~w2860;
assign w4899 = ~w4893 & ~w4898;
assign w4900 = (~w4897 & ~w4893) | (~w4897 & w6402) | (~w4893 & w6402);
assign w4901 = (w4900 & ~w4827) | (w4900 & w6735) | (~w4827 & w6735);
assign w4902 = (w2546 & w3146) | (w2546 & w6403) | (w3146 & w6403);
assign w4903 = w1991 & ~w3164;
assign w4904 = ~w4902 & ~w4903;
assign w4905 = (w3483 & w6736) | (w3483 & w6737) | (w6736 & w6737);
assign w4906 = w4904 & w7776;
assign w4907 = ~w4905 & ~w4906;
assign w4908 = w4901 & w6404;
assign w4909 = (~w4907 & ~w4901) | (~w4907 & w6405) | (~w4901 & w6405);
assign w4910 = ~w4908 & ~w4909;
assign w4911 = (~w4832 & ~w4834) | (~w4832 & w6406) | (~w4834 & w6406);
assign w4912 = w2563 & w3942;
assign w4913 = w1968 & ~w3936;
assign w4914 = (w1976 & ~w3779) | (w1976 & w6407) | (~w3779 & w6407);
assign w4915 = (~w3472 & w6738) | (~w3472 & w6739) | (w6738 & w6739);
assign w4916 = (w3472 & w6410) | (w3472 & w6411) | (w6410 & w6411);
assign w4917 = ~w4915 & ~w4916;
assign w4918 = (w4917 & ~w3942) | (w4917 & w6412) | (~w3942 & w6412);
assign w4919 = ~w4912 & ~w4918;
assign w4920 = w4911 & w4919;
assign w4921 = ~w4911 & ~w4919;
assign w4922 = ~w4920 & ~w4921;
assign w4923 = w4910 & w4922;
assign w4924 = ~w4910 & ~w4922;
assign w4925 = ~w4923 & ~w4924;
assign w4926 = (~w4817 & ~w4819) | (~w4817 & w6413) | (~w4819 & w6413);
assign w4927 = w4925 & ~w4926;
assign w4928 = ~w4925 & w4926;
assign w4929 = ~w4927 & ~w4928;
assign w4930 = (~w4848 & ~w4762) | (~w4848 & w6414) | (~w4762 & w6414);
assign w4931 = w4929 & w4930;
assign w4932 = ~w290 & w614;
assign w4933 = w690 & w4505;
assign w4934 = w4932 & w4933;
assign w4935 = w758 & w787;
assign w4936 = w4934 & w4935;
assign w4937 = w3615 & w4936;
assign w4938 = w248 & w3652;
assign w4939 = w4937 & w4938;
assign w4940 = w455 & w4939;
assign w4941 = ~w4885 & w6740;
assign w4942 = ~w4929 & w4940;
assign w4943 = (w4885 & w4942) | (w4885 & w6741) | (w4942 & w6741);
assign w4944 = ~w4941 & ~w4943;
assign w4945 = (w4885 & ~w4929) | (w4885 & w6742) | (~w4929 & w6742);
assign w4946 = (w4885 & ~w4940) | (w4885 & w6743) | (~w4940 & w6743);
assign w4947 = ~w4945 & w4946;
assign w4948 = w4944 & ~w4947;
assign w4949 = ~w4859 & ~w4865;
assign w4950 = w4805 & ~w4949;
assign w4951 = ~w4477 & w4950;
assign w4952 = ~w4951 & w5797;
assign w4953 = (w4948 & w4951) | (w4948 & w5798) | (w4951 & w5798);
assign w4954 = ~w4952 & ~w4953;
assign w4955 = w4876 & ~w4954;
assign w4956 = ~w4876 & w4954;
assign w4957 = ~w4955 & ~w4956;
assign w4958 = ~w4878 & w4879;
assign w4959 = (w3829 & ~w4879) | (w3829 & w6415) | (~w4879 & w6415);
assign w4960 = w4957 & ~w4959;
assign w4961 = ~w4957 & w4959;
assign w4962 = ~w4960 & ~w4961;
assign w4963 = w4866 & w4944;
assign w4964 = ~w4807 & w4963;
assign w4965 = ~w4806 & w4964;
assign w4966 = (~w4920 & ~w4922) | (~w4920 & w6416) | (~w4922 & w6416);
assign w4967 = (w4827 & w6744) | (w4827 & w6745) | (w6744 & w6745);
assign w4968 = (~w4967 & ~w6404) | (~w4967 & w7320) | (~w6404 & w7320);
assign w4969 = (~w1022 & w3146) | (~w1022 & w6417) | (w3146 & w6417);
assign w4970 = (~w4887 & ~w4889) | (~w4887 & w6418) | (~w4889 & w6418);
assign w4971 = w4969 & ~w4970;
assign w4972 = (~w1022 & ~w4970) | (~w1022 & w6419) | (~w4970 & w6419);
assign w4973 = ~w4971 & w4972;
assign w4974 = w1991 & ~w3474;
assign w4975 = w2546 & ~w3164;
assign w4976 = ~w3472 & w6420;
assign w4977 = ~w4974 & ~w4975;
assign w4978 = ~w4976 & w4977;
assign w4979 = w4973 & w7777;
assign w4980 = (w3568 & w6422) | (w3568 & w6423) | (w6422 & w6423);
assign w4981 = ~w4979 & ~w4980;
assign w4982 = w1976 & ~w3936;
assign w4983 = (w1974 & ~w3779) | (w1974 & w6424) | (~w3779 & w6424);
assign w4984 = (~w4071 & w6746) | (~w4071 & w6747) | (w6746 & w6747);
assign w4985 = (w4071 & w6426) | (w4071 & w6427) | (w6426 & w6427);
assign w4986 = ~w4984 & ~w4985;
assign w4987 = w4981 & ~w4986;
assign w4988 = ~w4981 & w4986;
assign w4989 = ~w4987 & ~w4988;
assign w4990 = w4968 & w4989;
assign w4991 = ~w4968 & ~w4989;
assign w4992 = ~w4990 & ~w4991;
assign w4993 = ~w4966 & ~w4992;
assign w4994 = w4966 & w4992;
assign w4995 = ~w4993 & ~w4994;
assign w4996 = w397 & w591;
assign w4997 = w598 & w906;
assign w4998 = w4996 & w4997;
assign w4999 = w3770 & w4998;
assign w5000 = w225 & w4999;
assign w5001 = ~w4995 & w5000;
assign w5002 = (w4885 & w5835) | (w4885 & w6748) | (w5835 & w6748);
assign w5003 = w4995 & w5000;
assign w5004 = (~w4885 & w6749) | (~w4885 & w6750) | (w6749 & w6750);
assign w5005 = ~w5002 & ~w5004;
assign w5006 = w4995 & ~w5000;
assign w5007 = (w4885 & w5839) | (w4885 & w6751) | (w5839 & w6751);
assign w5008 = ~w4995 & ~w5000;
assign w5009 = (~w4885 & w6752) | (~w4885 & w6753) | (w6752 & w6753);
assign w5010 = ~w5007 & ~w5009;
assign w5011 = w5005 & w5010;
assign w5012 = w4944 & w4949;
assign w5013 = (~w4947 & ~w4949) | (~w4947 & w6428) | (~w4949 & w6428);
assign w5014 = ~w5011 & w5013;
assign w5015 = (w5014 & w4806) | (w5014 & w6429) | (w4806 & w6429);
assign w5016 = ~w4807 & w6754;
assign w5017 = ~w4806 & w5016;
assign w5018 = w5011 & ~w5013;
assign w5019 = ~w5017 & ~w5018;
assign w5020 = ~w5015 & w5019;
assign w5021 = ~w4954 & w5020;
assign w5022 = w4876 & w5021;
assign w5023 = (~w5020 & ~w4876) | (~w5020 & w5799) | (~w4876 & w5799);
assign w5024 = ~w5022 & ~w5023;
assign w5025 = ~w4957 & w4958;
assign w5026 = (w3829 & ~w4958) | (w3829 & w6430) | (~w4958 & w6430);
assign w5027 = ~w5024 & ~w5026;
assign w5028 = w5024 & w5026;
assign w5029 = ~w5027 & ~w5028;
assign w5030 = ~w5012 & w5800;
assign w5031 = ~w4927 & ~w4993;
assign w5032 = (~w4994 & w4927) | (~w4994 & w6431) | (w4927 & w6431);
assign w5033 = w4929 & ~w4994;
assign w5034 = (~w5032 & ~w4930) | (~w5032 & w6755) | (~w4930 & w6755);
assign w5035 = w4883 & w5031;
assign w5036 = (~w5034 & ~w4883) | (~w5034 & w6756) | (~w4883 & w6756);
assign w5037 = (w6096 & w7321) | (w6096 & w7322) | (w7321 & w7322);
assign w5038 = (w565 & w6435) | (w565 & w7876) | (w6435 & w7876);
assign w5039 = ~w5037 & ~w5038;
assign w5040 = (w1987 & ~w3779) | (w1987 & w6436) | (~w3779 & w6436);
assign w5041 = (~w5040 & w3474) | (~w5040 & w6437) | (w3474 & w6437);
assign w5042 = (w3790 & w7323) | (w3790 & w7324) | (w7323 & w7324);
assign w5043 = w5041 & w7877;
assign w5044 = ~w5042 & ~w5043;
assign w5045 = w5039 & ~w5044;
assign w5046 = ~w5039 & w5044;
assign w5047 = ~w5045 & ~w5046;
assign w5048 = ~w1022 & w3195;
assign w5049 = (w6438 & w6759) | (w6438 & w6760) | (w6759 & w6760);
assign w5050 = (w6440 & ~w6438) | (w6440 & w6761) | (~w6438 & w6761);
assign w5051 = ~w5049 & ~w5050;
assign w5052 = w5047 & w5051;
assign w5053 = ~w5047 & ~w5051;
assign w5054 = ~w5052 & ~w5053;
assign w5055 = ~w4987 & ~w4990;
assign w5056 = w5054 & w5055;
assign w5057 = ~w5054 & ~w5055;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = ~w264 & ~w609;
assign w5060 = ~w691 & w5059;
assign w5061 = w1787 & w5060;
assign w5062 = ~w177 & w1900;
assign w5063 = w3616 & w5062;
assign w5064 = w680 & w5063;
assign w5065 = w4090 & w5061;
assign w5066 = w5064 & w5065;
assign w5067 = w1920 & w5066;
assign w5068 = w2628 & w5067;
assign w5069 = w5058 & ~w5068;
assign w5070 = ~w5058 & w5068;
assign w5071 = ~w5069 & ~w5070;
assign w5072 = (w5657 & w5801) | (w5657 & w5802) | (w5801 & w5802);
assign w5073 = (~w5657 & w5803) | (~w5657 & w5804) | (w5803 & w5804);
assign w5074 = ~w5072 & ~w5073;
assign w5075 = ~w5017 & w5805;
assign w5076 = (w5074 & w5017) | (w5074 & w5806) | (w5017 & w5806);
assign w5077 = ~w5075 & ~w5076;
assign w5078 = (~w5077 & ~w4876) | (~w5077 & w6762) | (~w4876 & w6762);
assign w5079 = w4876 & w6763;
assign w5080 = ~w5078 & ~w5079;
assign w5081 = (w5026 & w6442) | (w5026 & w6443) | (w6442 & w6443);
assign w5082 = ~w5080 & w7778;
assign w5083 = ~w5081 & ~w5082;
assign w5084 = (~w5046 & ~w5047) | (~w5046 & w7325) | (~w5047 & w7325);
assign w5085 = w3164 & w4969;
assign w5086 = (~w6438 & w6764) | (~w6438 & w6765) | (w6764 & w6765);
assign w5087 = (w565 & w3164) | (w565 & w6446) | (w3164 & w6446);
assign w5088 = ~w3164 & w6447;
assign w5089 = ~w5087 & ~w5088;
assign w5090 = ~w1022 & ~w3474;
assign w5091 = w5089 & w5090;
assign w5092 = ~w5089 & ~w5090;
assign w5093 = ~w5091 & ~w5092;
assign w5094 = (w1991 & ~w3779) | (w1991 & w6449) | (~w3779 & w6449);
assign w5095 = w1987 & ~w3936;
assign w5096 = (w6451 & ~w3942) | (w6451 & w6766) | (~w3942 & w6766);
assign w5097 = (w3942 & w6767) | (w3942 & w6768) | (w6767 & w6768);
assign w5098 = ~w5096 & ~w5097;
assign w5099 = w5093 & w5098;
assign w5100 = ~w5093 & ~w5098;
assign w5101 = ~w5099 & ~w5100;
assign w5102 = ~w5086 & w5101;
assign w5103 = w5086 & ~w5101;
assign w5104 = ~w5102 & ~w5103;
assign w5105 = ~w5084 & w5104;
assign w5106 = w5084 & ~w5104;
assign w5107 = ~w5105 & ~w5106;
assign w5108 = ~w5057 & w5107;
assign w5109 = (~w4496 & w6769) | (~w4496 & w6770) | (w6769 & w6770);
assign w5110 = ~w5056 & ~w5107;
assign w5111 = w5057 & ~w5107;
assign w5112 = (~w4496 & w6771) | (~w4496 & w6772) | (w6771 & w6772);
assign w5113 = ~w5109 & w5112;
assign w5114 = ~w58 & ~w160;
assign w5115 = ~w268 & w5114;
assign w5116 = w677 & w5115;
assign w5117 = ~w122 & ~w215;
assign w5118 = ~w517 & w5117;
assign w5119 = w611 & w3664;
assign w5120 = w5118 & w5119;
assign w5121 = w3838 & w5120;
assign w5122 = w626 & w5116;
assign w5123 = w5121 & w5122;
assign w5124 = w493 & w2750;
assign w5125 = w5123 & w5124;
assign w5126 = w4091 & w5125;
assign w5127 = w5113 & ~w5126;
assign w5128 = ~w5113 & w5126;
assign w5129 = ~w5127 & ~w5128;
assign w5130 = ~w5068 & ~w5074;
assign w5131 = w5129 & w5130;
assign w5132 = ~w5129 & ~w5130;
assign w5133 = ~w5131 & ~w5132;
assign w5134 = w5077 & w5133;
assign w5135 = w4876 & w6773;
assign w5136 = ~w5133 & ~w5076;
assign w5137 = (w5030 & w4806) | (w5030 & w5807) | (w4806 & w5807);
assign w5138 = w5005 & w5074;
assign w5139 = ~w5128 & w5138;
assign w5140 = (~w5807 & w6774) | (~w5807 & w6775) | (w6774 & w6775);
assign w5141 = w6452 & ~w5137;
assign w5142 = ~w5136 & ~w5141;
assign w5143 = (~w4876 & w6776) | (~w4876 & w6777) | (w6776 & w6777);
assign w5144 = ~w5135 & ~w5143;
assign w5145 = ~w5024 & ~w5080;
assign w5146 = w5025 & w5145;
assign w5147 = (w5025 & w6778) | (w5025 & w6779) | (w6778 & w6779);
assign w5148 = (w6454 & ~w5025) | (w6454 & w6780) | (~w5025 & w6780);
assign w5149 = ~w5147 & ~w5148;
assign w5150 = ~w5056 & ~w5105;
assign w5151 = (~w5105 & ~w5107) | (~w5105 & w6455) | (~w5107 & w6455);
assign w5152 = (~w5099 & ~w5101) | (~w5099 & w6456) | (~w5101 & w6456);
assign w5153 = ~w3472 & w6457;
assign w5154 = (~w5088 & ~w5089) | (~w5088 & w6458) | (~w5089 & w6458);
assign w5155 = ~w5153 & ~w5154;
assign w5156 = w5153 & w5154;
assign w5157 = ~w5155 & ~w5156;
assign w5158 = w1991 & ~w3936;
assign w5159 = (w2546 & ~w3779) | (w2546 & w6459) | (~w3779 & w6459);
assign w5160 = (~w4071 & w6781) | (~w4071 & w6782) | (w6781 & w6782);
assign w5161 = ~w5160 & w6463;
assign w5162 = (~w5157 & w5160) | (~w5157 & w6464) | (w5160 & w6464);
assign w5163 = ~w5161 & ~w5162;
assign w5164 = (w5101 & w7631) | (w5101 & w7632) | (w7631 & w7632);
assign w5165 = ~w5163 & w5152;
assign w5166 = ~w5164 & ~w5165;
assign w5167 = ~w189 & ~w254;
assign w5168 = ~w271 & w5167;
assign w5169 = w229 & w367;
assign w5170 = w1900 & w2738;
assign w5171 = w4505 & w5170;
assign w5172 = w5168 & w5169;
assign w5173 = w5171 & w5172;
assign w5174 = w551 & w5173;
assign w5175 = w775 & w1659;
assign w5176 = w5174 & w5175;
assign w5177 = w1569 & w5176;
assign w5178 = w5166 & w5177;
assign w5179 = (~w4496 & w6783) | (~w4496 & w6784) | (w6783 & w6784);
assign w5180 = ~w5166 & w5177;
assign w5181 = (w4496 & w6785) | (w4496 & w6786) | (w6785 & w6786);
assign w5182 = ~w5179 & ~w5181;
assign w5183 = (~w4496 & w6787) | (~w4496 & w6788) | (w6787 & w6788);
assign w5184 = (w4496 & w6789) | (w4496 & w6790) | (w6789 & w6790);
assign w5185 = ~w5183 & ~w5184;
assign w5186 = ~w5177 & ~w5185;
assign w5187 = w5182 & ~w5186;
assign w5188 = ~w5127 & ~w5130;
assign w5189 = ~w5128 & ~w5188;
assign w5190 = ~w5139 & ~w5189;
assign w5191 = w5030 & ~w5189;
assign w5192 = (~w5190 & w4965) | (~w5190 & w5809) | (w4965 & w5809);
assign w5193 = ~w5187 & w5192;
assign w5194 = w5187 & ~w5192;
assign w5195 = ~w5193 & ~w5194;
assign w5196 = w5022 & w5810;
assign w5197 = (w5195 & ~w5022) | (w5195 & w5811) | (~w5022 & w5811);
assign w5198 = ~w5196 & ~w5197;
assign w5199 = w5198 & w7779;
assign w5200 = (w5146 & w6791) | (w5146 & w6792) | (w6791 & w6792);
assign w5201 = ~w5199 & ~w5200;
assign w5202 = (w6096 & w7326) | (w6096 & w7327) | (w7326 & w7327);
assign w5203 = ~w3784 & w5262;
assign w5204 = ~w5202 & ~w5203;
assign w5205 = (w6469 & ~w6463) | (w6469 & w6795) | (~w6463 & w6795);
assign w5206 = (w6463 & w6796) | (w6463 & w6797) | (w6796 & w6797);
assign w5207 = ~w5205 & ~w5206;
assign w5208 = (w5207 & ~w5152) | (w5207 & w6471) | (~w5152 & w6471);
assign w5209 = w5152 & w6472;
assign w5210 = ~w5208 & ~w5209;
assign w5211 = ~w5166 & w5210;
assign w5212 = w5150 & ~w5211;
assign w5213 = w5151 & w5166;
assign w5214 = (w5210 & ~w5151) | (w5210 & w5211) | (~w5151 & w5211);
assign w5215 = (~w4496 & w6798) | (~w4496 & w6799) | (w6798 & w6799);
assign w5216 = w5150 & ~w5164;
assign w5217 = w5150 & w6473;
assign w5218 = w5151 & w6474;
assign w5219 = (~w4496 & w6800) | (~w4496 & w6801) | (w6800 & w6801);
assign w5220 = ~w5215 & w5219;
assign w5221 = ~w231 & w1504;
assign w5222 = w639 & w6475;
assign w5223 = ~w227 & ~w291;
assign w5224 = w416 & w5223;
assign w5225 = w1666 & w1671;
assign w5226 = w5224 & w5225;
assign w5227 = w3632 & w5226;
assign w5228 = w5061 & w5227;
assign w5229 = w476 & w5228;
assign w5230 = w1906 & w5229;
assign w5231 = w5222 & w5230;
assign w5232 = ~w5220 & ~w5231;
assign w5233 = w5220 & w5231;
assign w5234 = ~w5232 & ~w5233;
assign w5235 = ~w5186 & ~w5234;
assign w5236 = ~w5234 & w5847;
assign w5237 = w5139 & ~w5236;
assign w5238 = ~w5188 & w6476;
assign w5239 = w5235 & ~w5238;
assign w5240 = (w5239 & w5137) | (w5239 & w6477) | (w5137 & w6477);
assign w5241 = ~w5186 & ~w5232;
assign w5242 = ~w5189 & w5241;
assign w5243 = w5182 & ~w5233;
assign w5244 = ~w5232 & w5243;
assign w5245 = ~w5242 & w5244;
assign w5246 = w5139 & w5244;
assign w5247 = (~w5807 & w6802) | (~w5807 & w6803) | (w6802 & w6803);
assign w5248 = ~w5245 & ~w5247;
assign w5249 = ~w5240 & w5248;
assign w5250 = ~w5195 & w5249;
assign w5251 = w5135 & w5250;
assign w5252 = (~w5249 & ~w5022) | (~w5249 & w6804) | (~w5022 & w6804);
assign w5253 = ~w5251 & ~w5252;
assign w5254 = ~w5144 & ~w5198;
assign w5255 = w5146 & w5254;
assign w5256 = (w3829 & ~w5146) | (w3829 & w5848) | (~w5146 & w5848);
assign w5257 = (w5146 & w7328) | (w5146 & w7329) | (w7328 & w7329);
assign w5258 = w5253 & w5256;
assign w5259 = ~w5257 & ~w5258;
assign w5260 = (w5208 & ~w5151) | (w5208 & w6478) | (~w5151 & w6478);
assign w5261 = ~w1022 & ~w3939;
assign w5262 = (~w1022 & w3936) | (~w1022 & w7878) | (w3936 & w7878);
assign w5263 = ~w5202 & ~w5262;
assign w5264 = ~w3472 & w6479;
assign w5265 = ~w5263 & w6480;
assign w5266 = (w5261 & w5263) | (w5261 & w6481) | (w5263 & w6481);
assign w5267 = ~w5265 & ~w5266;
assign w5268 = ~w155 & ~w197;
assign w5269 = ~w273 & ~w538;
assign w5270 = w5268 & w5269;
assign w5271 = w255 & w3121;
assign w5272 = w5270 & w5271;
assign w5273 = w2316 & w5272;
assign w5274 = w3607 & w5116;
assign w5275 = w5273 & w5274;
assign w5276 = w3631 & w5275;
assign w5277 = w2181 & w5276;
assign w5278 = ~w5267 & ~w5277;
assign w5279 = (w4496 & w7518) | (w4496 & w7270) | (w7518 & w7270);
assign w5280 = w5267 & w5277;
assign w5281 = ~w5278 & ~w5280;
assign w5282 = (~w5277 & ~w5204) | (~w5277 & w7879) | (~w5204 & w7879);
assign w5283 = (~w4496 & w7522) | (~w4496 & w7271) | (w7522 & w7271);
assign w5284 = ~w5279 & ~w5283;
assign w5285 = ~w5247 & w5849;
assign w5286 = (w5284 & w5247) | (w5284 & w5850) | (w5247 & w5850);
assign w5287 = ~w5285 & ~w5286;
assign w5288 = w5135 & w5812;
assign w5289 = (~w5287 & ~w5135) | (~w5287 & w5813) | (~w5135 & w5813);
assign w5290 = ~w5288 & ~w5289;
assign w5291 = w5290 & w7780;
assign w5292 = (w5256 & w6485) | (w5256 & w6486) | (w6485 & w6486);
assign w5293 = ~w5291 & ~w5292;
assign w5294 = ~w5253 & ~w5290;
assign w5295 = w5146 & w6805;
assign w5296 = (~w4496 & w7330) | (~w4496 & w7331) | (w7330 & w7331);
assign w5297 = ~w5189 & w6593;
assign w5298 = ~w5232 & ~w5243;
assign w5299 = ~w620 & ~w691;
assign w5300 = w804 & w5299;
assign w5301 = w2817 & w3603;
assign w5302 = w5300 & w5301;
assign w5303 = w813 & w3654;
assign w5304 = w5302 & w5303;
assign w5305 = w351 & w5304;
assign w5306 = w344 & w5305;
assign w5307 = w3131 & w5306;
assign w5308 = (w6491 & w5243) | (w6491 & w7633) | (w5243 & w7633);
assign w5309 = (w5308 & w5140) | (w5308 & w6492) | (w5140 & w6492);
assign w5310 = (~w5243 & w7634) | (~w5243 & w7635) | (w7634 & w7635);
assign w5311 = ~w5189 & w6494;
assign w5312 = (~w5137 & w6806) | (~w5137 & w6807) | (w6806 & w6807);
assign w5313 = ~w5309 & w5312;
assign w5314 = w5288 & ~w5313;
assign w5315 = ~w5288 & w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = (w5255 & w6808) | (w5255 & w6809) | (w6808 & w6809);
assign w5318 = ~w5316 & w7781;
assign w5319 = ~w5317 & ~w5318;
assign w5320 = w5255 & w5814;
assign w5321 = ~w124 & w466;
assign w5322 = w2291 & w4232;
assign w5323 = w5321 & w5322;
assign w5324 = w208 & w2743;
assign w5325 = w5323 & w5324;
assign w5326 = w464 & w1556;
assign w5327 = w5325 & w5326;
assign w5328 = w596 & w5327;
assign w5329 = w364 & w3660;
assign w5330 = w5328 & w5329;
assign w5331 = (w5137 & w6810) | (w5137 & w6811) | (w6810 & w6811);
assign w5332 = (w5662 & w5140) | (w5662 & w6496) | (w5140 & w6496);
assign w5333 = w5284 & ~w5330;
assign w5334 = ~w5243 & w6497;
assign w5335 = (w5139 & ~w5298) | (w5139 & w5851) | (~w5298 & w5851);
assign w5336 = (~w5807 & w6812) | (~w5807 & w6813) | (w6812 & w6813);
assign w5337 = (w5333 & w5242) | (w5333 & w5334) | (w5242 & w5334);
assign w5338 = ~w5336 & w5337;
assign w5339 = ~w5284 & ~w5330;
assign w5340 = ~w5242 & w5663;
assign w5341 = ~w5298 & w5852;
assign w5342 = (~w5807 & w6814) | (~w5807 & w6815) | (w6814 & w6815);
assign w5343 = ~w5340 & ~w5342;
assign w5344 = ~w5338 & w5343;
assign w5345 = w5312 & ~w5344;
assign w5346 = w5135 & w5853;
assign w5347 = (~w5140 & w6816) | (~w5140 & w6817) | (w6816 & w6817);
assign w5348 = ~w5288 & w5347;
assign w5349 = ~w5331 & ~w5332;
assign w5350 = ~w5346 & w5349;
assign w5351 = ~w5348 & w5350;
assign w5352 = ~w5351 & w7782;
assign w5353 = (w5295 & w6498) | (w5295 & w6499) | (w6498 & w6499);
assign w5354 = ~w5352 & ~w5353;
assign w5355 = ~w158 & ~w187;
assign w5356 = w761 & w5355;
assign w5357 = w3115 & w5356;
assign w5358 = w185 & w4453;
assign w5359 = w5357 & w5358;
assign w5360 = w3101 & w5359;
assign w5361 = w670 & w5360;
assign w5362 = w5222 & w5361;
assign w5363 = (w5140 & w7332) | (w5140 & w7333) | (w7332 & w7333);
assign w5364 = (~w5140 & w7334) | (~w5140 & w7335) | (w7334 & w7335);
assign w5365 = ~w5363 & ~w5364;
assign w5366 = w5313 & ~w5344;
assign w5367 = w5251 & w5854;
assign w5368 = (~w5365 & ~w5251) | (~w5365 & w5855) | (~w5251 & w5855);
assign w5369 = ~w5367 & ~w5368;
assign w5370 = w3829 & w5351;
assign w5371 = (w5295 & ~w3829) | (w5295 & w5856) | (~w3829 & w5856);
assign w5372 = w5369 & ~w5371;
assign w5373 = ~w5369 & w5371;
assign w5374 = ~w5372 & ~w5373;
assign w5375 = ~w5351 & ~w5369;
assign w5376 = w5255 & w6818;
assign w5377 = ~w179 & w545;
assign w5378 = w1032 & w3602;
assign w5379 = w4678 & w5378;
assign w5380 = w4452 & w5377;
assign w5381 = w5379 & w5380;
assign w5382 = w908 & w5381;
assign w5383 = w756 & w5382;
assign w5384 = w4770 & w5383;
assign w5385 = ~w5362 & ~w5384;
assign w5386 = (~w5140 & w6500) | (~w5140 & w6501) | (w6500 & w6501);
assign w5387 = ~w5344 & w6502;
assign w5388 = w5135 & w6503;
assign w5389 = (~w5140 & w7336) | (~w5140 & w7337) | (w7336 & w7337);
assign w5390 = (w5665 & w5140) | (w5665 & w6505) | (w5140 & w6505);
assign w5391 = ~w5389 & ~w5390;
assign w5392 = (~w5388 & w5367) | (~w5388 & w5666) | (w5367 & w5666);
assign w5393 = (w5320 & w6819) | (w5320 & w6820) | (w6819 & w6820);
assign w5394 = (~w5320 & w5396) | (~w5320 & w6821) | (w5396 & w6821);
assign w5395 = ~w5393 & ~w5394;
assign w5396 = w3829 & ~w5392;
assign w5397 = w818 & ~w2314;
assign w5398 = w908 & w5397;
assign w5399 = w428 & w5398;
assign w5400 = w1063 & w5399;
assign w5401 = (w5857 & ~w5297) | (w5857 & w7783) | (~w5297 & w7783);
assign w5402 = (w5137 & w6823) | (w5137 & w6824) | (w6823 & w6824);
assign w5403 = ~w5401 & ~w5402;
assign w5404 = w5251 & w5815;
assign w5405 = (~w5403 & ~w5251) | (~w5403 & w5816) | (~w5251 & w5816);
assign w5406 = ~w5404 & ~w5405;
assign w5407 = w3829 & ~w5406;
assign w5408 = ~w3829 & w5406;
assign w5409 = ~w5407 & ~w5408;
assign w5410 = (w5409 & ~w5320) | (w5409 & w6825) | (~w5320 & w6825);
assign w5411 = ~w5392 & w5407;
assign w5412 = w5376 & w5411;
assign w5413 = ~w5410 & ~w5412;
assign w5414 = w1063 & w6506;
assign w5415 = (w5388 & w5817) | (w5388 & w5818) | (w5817 & w5818);
assign w5416 = (~w5388 & w5819) | (~w5388 & w5820) | (w5819 & w5820);
assign w5417 = ~w5415 & ~w5416;
assign w5418 = w3829 & ~w5417;
assign w5419 = ~w3829 & w5417;
assign w5420 = ~w5418 & ~w5419;
assign w5421 = (~w5420 & ~w5376) | (~w5420 & w6507) | (~w5376 & w6507);
assign w5422 = w5376 & w5668;
assign w5423 = ~w5421 & ~w5422;
assign w5424 = (w5320 & w6826) | (w5320 & w6827) | (w6826 & w6827);
assign w5425 = w11 & w6508;
assign w5426 = (w5388 & w7338) | (w5388 & w7339) | (w7338 & w7339);
assign w5427 = ~w5406 & ~w5425;
assign w5428 = w5427 & w6509;
assign w5429 = (~w5426 & ~w5376) | (~w5426 & w6510) | (~w5376 & w6510);
assign w5430 = ~w5424 & ~w5429;
assign w5431 = w5376 & w6511;
assign w5432 = w3829 & ~w5431;
assign w5433 = ~w13 & w16;
assign w5434 = ~w20 & ~w22;
assign w5435 = ~w25 & w28;
assign w5436 = ~w32 & w34;
assign w5437 = ~w45 & w47;
assign w5438 = ~w32 & w59;
assign w5439 = w15 & ~w61;
assign w5440 = ~w62 & ~w63;
assign w5441 = ~w13 & w66;
assign w5442 = ~w32 & ~w68;
assign w5443 = ~w45 & w72;
assign w5444 = ~w13 & w19;
assign w5445 = ~w84 & ~w83;
assign w5446 = ~w32 & w91;
assign w5447 = w15 & ~w33;
assign w5448 = ~w93 & ~w94;
assign w5449 = ~w45 & w98;
assign w5450 = ~w32 & w110;
assign w5451 = ~w45 & w50;
assign w5452 = ~w13 & w134;
assign w5453 = ~w136 & ~w137;
assign w5454 = w65 & ~w139;
assign w5455 = ~w279 & ~w332;
assign w5456 = w418 & w427;
assign w5457 = w410 & w429;
assign w5458 = ~w455 & ~w511;
assign w5459 = ~w511 & ~w512;
assign w5460 = ~w455 & ~w565;
assign w5461 = ~w565 & ~w566;
assign w5462 = ~w455 & ~w735;
assign w5463 = w828 & w6512;
assign w5464 = ~w455 & ~w880;
assign w5465 = ~w880 & ~w881;
assign w5466 = ~w917 & w919;
assign w5467 = ~w455 & w720;
assign w5468 = (~w726 & ~w828) | (~w726 & w6513) | (~w828 & w6513);
assign w5469 = w828 & w6514;
assign w5470 = w978 & ~w921;
assign w5471 = ~w978 & w921;
assign w5472 = w828 & w6515;
assign w5473 = (~w720 & ~w828) | (~w720 & w6516) | (~w828 & w6516);
assign w5474 = ~w455 & w1022;
assign w5475 = w1022 & ~w1023;
assign w5476 = w96 & ~w86;
assign w5477 = w990 & ~w991;
assign w5478 = w828 & w6517;
assign w5479 = (~w735 & ~w828) | (~w735 & w6518) | (~w828 & w6518);
assign w5480 = ~w735 & ~w736;
assign w5481 = w828 & w6519;
assign w5482 = (~w574 & ~w828) | (~w574 & w6520) | (~w828 & w6520);
assign w5483 = ~w392 & ~w1157;
assign w5484 = (~w565 & ~w828) | (~w565 & w6521) | (~w828 & w6521);
assign w5485 = w828 & w6522;
assign w5486 = w1023 & w1226;
assign w5487 = ~w1023 & ~w1226;
assign w5488 = ~w1247 & ~w1195;
assign w5489 = ~w1222 & ~w1213;
assign w5490 = ~w1229 & ~w1227;
assign w5491 = ~w1189 & ~w1187;
assign w5492 = w828 & w6523;
assign w5493 = (~w511 & ~w828) | (~w511 & w6524) | (~w828 & w6524);
assign w5494 = ~w1404 & ~w1396;
assign w5495 = ~w1385 & ~w1373;
assign w5496 = (w847 & ~w837) | (w847 & w6525) | (~w837 & w6525);
assign w5497 = w837 & w6526;
assign w5498 = ~w1489 & w1495;
assign w5499 = w1593 & w1591;
assign w5500 = w828 & w6527;
assign w5501 = (w880 & ~w828) | (w880 & w6528) | (~w828 & w6528);
assign w5502 = ~w1284 & w1640;
assign w5503 = ~w1711 & w1715;
assign w5504 = ~w1657 & w6530;
assign w5505 = ~w1731 & ~w1736;
assign w5506 = w828 & w6531;
assign w5507 = (w1022 & ~w828) | (w1022 & w6532) | (~w828 & w6532);
assign w5508 = ~w1621 & ~w1612;
assign w5509 = w650 & w1259;
assign w5510 = ~w650 & ~w1259;
assign w5511 = w1628 & ~w1775;
assign w5512 = ~w1650 & ~w1800;
assign w5513 = w1650 & w1800;
assign w5514 = ~w1701 & ~w1812;
assign w5515 = w1806 & w1800;
assign w5516 = w1753 & w1843;
assign w5517 = ~w1753 & ~w1843;
assign w5518 = ~w1748 & ~w1739;
assign w5519 = ~w1875 & ~w1880;
assign w5520 = w1758 & ~w1894;
assign w5521 = ~w1898 & w1934;
assign w5522 = ~w1938 & w1940;
assign w5523 = ~w1945 & ~w1943;
assign w5524 = (w1963 & w1819) | (w1963 & w5669) | (w1819 & w5669);
assign w5525 = ~w1820 & w1976;
assign w5526 = (~w1987 & w1710) | (~w1987 & w6533) | (w1710 & w6533);
assign w5527 = ~w1964 & w2007;
assign w5528 = w1964 & w2009;
assign w5529 = w1964 & w2012;
assign w5530 = ~w1820 & w1968;
assign w5531 = (~w1976 & w1710) | (~w1976 & w6534) | (w1710 & w6534);
assign w5532 = (~w1968 & w1710) | (~w1968 & w6535) | (w1710 & w6535);
assign w5533 = (w1710 & w6536) | (w1710 & w6537) | (w6536 & w6537);
assign w5534 = w2024 & w6538;
assign w5535 = w1864 & ~w2086;
assign w5536 = ~w1864 & w2086;
assign w5537 = w838 & w1633;
assign w5538 = ~w2122 & ~w2127;
assign w5539 = w2096 & ~w2151;
assign w5540 = ~w2096 & w2151;
assign w5541 = w2113 & w2197;
assign w5542 = w1931 & ~w1896;
assign w5543 = ~w1897 & ~w2205;
assign w5544 = (~w5543 & w6539) | (~w5543 & w6540) | (w6539 & w6540);
assign w5545 = (w5543 & w6541) | (w5543 & w6542) | (w6541 & w6542);
assign w5546 = ~w2206 & w2232;
assign w5547 = w2206 & ~w2232;
assign w5548 = ~w2236 & w6543;
assign w5549 = (~w2204 & w2236) | (~w2204 & w6544) | (w2236 & w6544);
assign w5550 = ~w1949 & w2243;
assign w5551 = ~w2129 & ~w2255;
assign w5552 = w2129 & w2255;
assign w5553 = (~w2287 & ~w2288) | (~w2287 & w5670) | (~w2288 & w5670);
assign w5554 = w2113 & w2342;
assign w5555 = ~w2114 & w2348;
assign w5556 = ~w2375 & w2383;
assign w5557 = ~w2387 & ~w2386;
assign w5558 = ~w2237 & w5671;
assign w5559 = w2237 & w2424;
assign w5560 = ~w2375 & ~w2377;
assign w5561 = ~w1822 & w2374;
assign w5562 = w2461 & w2394;
assign w5563 = w2461 & w2396;
assign w5564 = (w2244 & w6545) | (w2244 & w6546) | (w6545 & w6546);
assign w5565 = ~w2244 & w6547;
assign w5566 = (~w2436 & w1710) | (~w2436 & w6548) | (w1710 & w6548);
assign w5567 = (~w2045 & w5674) | (~w2045 & ~w2489) | (w5674 & ~w2489);
assign w5568 = ~w1820 & w2411;
assign w5569 = (w726 & ~w1819) | (w726 & w5675) | (~w1819 & w5675);
assign w5570 = w2488 & w6549;
assign w5571 = w1819 & w5822;
assign w5572 = (~w726 & ~w1955) | (~w726 & w5678) | (~w1955 & w5678);
assign w5573 = w1955 & w5679;
assign w5574 = ~w1994 & w2002;
assign w5575 = (~w1991 & w1710) | (~w1991 & w6550) | (w1710 & w6550);
assign w5576 = ~w2549 & w2542;
assign w5577 = w2549 & ~w2542;
assign w5578 = ~w2245 & w1968;
assign w5579 = ~w1820 & w1974;
assign w5580 = w1942 & w1976;
assign w5581 = ~w1942 & w1976;
assign w5582 = w2554 & w565;
assign w5583 = ~w2554 & ~w2564;
assign w5584 = ~w2554 & ~w565;
assign w5585 = ~w2573 & ~w2574;
assign w5586 = w1588 & ~w2284;
assign w5587 = ~w2289 & w2589;
assign w5588 = ~w2355 & ~w2347;
assign w5589 = w2237 & w2650;
assign w5590 = w2237 & w2653;
assign w5591 = w2581 & w2661;
assign w5592 = ~w2581 & ~w2661;
assign w5593 = (w2117 & w6551) | (w2117 & w6552) | (w6551 & w6552);
assign w5594 = ~w2717 & w2719;
assign w5595 = (~w2725 & w5680) | (~w2725 & w7748) | (w5680 & w7748);
assign w5596 = (w2117 & w6553) | (w2117 & w6554) | (w6553 & w6554);
assign w5597 = ~w2717 & w2778;
assign w5598 = w2237 & w2784;
assign w5599 = ~w2802 & ~w2801;
assign w5600 = w2780 & w2204;
assign w5601 = w2237 & w2807;
assign w5602 = ~w2721 & w2780;
assign w5603 = ~w2809 & w2769;
assign w5604 = ~w2809 & w2814;
assign w5605 = (w2816 & w5681) | (w2816 & w7748) | (w5681 & w7748);
assign w5606 = w2809 & ~w2769;
assign w5607 = w2809 & w2895;
assign w5608 = ~w2862 & w2857;
assign w5609 = w1819 & w5682;
assign w5610 = w2461 & w2885;
assign w5611 = ~w1820 & w2903;
assign w5612 = w1710 & w3009;
assign w5613 = (~w6925 & ~w1715) | (~w6925 & w5683) | (~w1715 & w5683);
assign w5614 = (~w3031 & w6555) | (~w3031 & w6556) | (w6555 & w6556);
assign w5615 = w3031 & w7340;
assign w5616 = (~w3008 & ~w3019) | (~w3008 & w6828) | (~w3019 & w6828);
assign w5617 = (w871 & ~w1955) | (w871 & w5685) | (~w1955 & w5685);
assign w5618 = w1955 & w5686;
assign w5619 = ~w2896 & w3113;
assign w5620 = ~w2900 & w6557;
assign w5621 = (w2900 & w7113) | (w2900 & w6558) | (w7113 & w6558);
assign w5622 = ~w2896 & w3170;
assign w5623 = ~w2237 & w5689;
assign w5624 = w2237 & w3414;
assign w5625 = ~w1710 & ~w1022;
assign w5626 = w3507 & ~w3505;
assign w5627 = w3444 & ~w3443;
assign w5628 = ~w3719 & ~w3522;
assign w5629 = w2461 & w1994;
assign w5630 = ~w3748 & w3522;
assign w5631 = ~w3735 & ~w3875;
assign w5632 = w3763 & ~w3988;
assign w5633 = w3855 & ~w3909;
assign w5634 = w2385 & w4012;
assign w5635 = w4002 & w4016;
assign w5636 = ~w4002 & ~w4016;
assign w5637 = ~w4147 & ~w4035;
assign w5638 = ~w3896 & ~w4046;
assign w5639 = ~w4158 & ~w4266;
assign w5640 = (~w5639 & w6829) | (~w5639 & w6830) | (w6829 & w6830);
assign w5641 = (w5639 & w6831) | (w5639 & w6832) | (w6831 & w6832);
assign w5642 = (w4156 & ~w4019) | (w4156 & w6559) | (~w4019 & w6559);
assign w5643 = ~w4311 & ~w4180;
assign w5644 = ~w4214 & ~w4212;
assign w5645 = ~w4214 & ~w4213;
assign w5646 = ~w4358 & w4377;
assign w5647 = w4249 & ~w4478;
assign w5648 = (~w4143 & ~w4463) | (~w4143 & w6833) | (~w4463 & w6833);
assign w5649 = ~w4494 & w4582;
assign w5650 = (~w4450 & w4337) | (~w4450 & w5823) | (w4337 & w5823);
assign w5651 = ~w4473 & w5824;
assign w5652 = (~w4594 & w4473) | (~w4594 & w5825) | (w4473 & w5825);
assign w5653 = ~w4580 & w4666;
assign w5654 = w4491 & w4694;
assign w5655 = ~w4673 & w4711;
assign w5656 = ~w4673 & w4883;
assign w5657 = w4143 & w6560;
assign w5658 = ~w5206 & ~w5278;
assign w5659 = ~w5282 & ~w5281;
assign w5660 = (w4496 & w7341) | (w4496 & w7342) | (w7341 & w7342);
assign w5661 = ~w5316 & w3829;
assign w5662 = (w6567 & w5243) | (w6567 & w7636) | (w5243 & w7636);
assign w5663 = (w5339 & w5243) | (w5339 & w6568) | (w5243 & w6568);
assign w5664 = (~w5243 & w7651) | (~w5243 & w7637) | (w7651 & w7637);
assign w5665 = (w6569 & w5243) | (w6569 & w7638) | (w5243 & w7638);
assign w5666 = w5391 & ~w5388;
assign w5667 = w5375 & w5396;
assign w5668 = w5407 & w6570;
assign w5669 = (w1963 & w1816) | (w1963 & w6571) | (w1816 & w6571);
assign w5670 = ~w2286 & ~w2287;
assign w5671 = w2204 & w2411;
assign w5672 = (~w726 & ~w2403) | (~w726 & w6572) | (~w2403 & w6572);
assign w5673 = w2403 & w6573;
assign w5674 = (~w726 & w1710) | (~w726 & w6574) | (w1710 & w6574);
assign w5675 = (w726 & w2403) | (w726 & w6575) | (w2403 & w6575);
assign w5676 = ~w1710 & w6576;
assign w5677 = (w2436 & w1816) | (w2436 & w6577) | (w1816 & w6577);
assign w5678 = ~w726 & w7784;
assign w5679 = (w1819 & w6579) | (w1819 & w6580) | (w6579 & w6580);
assign w5680 = ~w2722 & ~w2725;
assign w5681 = ~w2722 & w2816;
assign w5682 = ~w2403 & w6581;
assign w5683 = (~w2903 & w1710) | (~w2903 & w6582) | (w1710 & w6582);
assign w5684 = (w3009 & w1816) | (w3009 & w6583) | (w1816 & w6583);
assign w5685 = w871 & w7786;
assign w5686 = (w1819 & w6839) | (w1819 & w6840) | (w6839 & w6840);
assign w5687 = w3142 & w3161;
assign w5688 = ~w3142 & ~w3161;
assign w5689 = w2204 & w1968;
assign w5690 = ~w4466 & ~w4463;
assign w5691 = ~w5150 & ~w5151;
assign w5692 = ~w5217 & ~w5218;
assign w5693 = w1759 & ~w1770;
assign w5694 = ~w1655 & ~w1831;
assign w5695 = w1656 & ~w1831;
assign w5696 = ~w1936 & ~w1938;
assign w5697 = ~w2228 & ~w2237;
assign w5698 = ~w2112 & w2288;
assign w5699 = ~w2408 & w2363;
assign w5700 = ~w2413 & ~w2414;
assign w5701 = ~w2430 & w2428;
assign w5702 = ~w2426 & ~w726;
assign w5703 = ~w2382 & w2394;
assign w5704 = w2382 & w2394;
assign w5705 = ~w2445 & ~w2456;
assign w5706 = ~w2667 & ~w2668;
assign w5707 = w2711 & ~w2287;
assign w5708 = w2711 & w5553;
assign w5709 = w5595 & ~w2766;
assign w5710 = ~w5595 & w2766;
assign w5711 = w2647 & ~w2782;
assign w5712 = ~w2783 & ~w2781;
assign w5713 = w2783 & w2781;
assign w5714 = ~w2648 & ~w2650;
assign w5715 = ~w2648 & ~w5589;
assign w5716 = w5605 & w2849;
assign w5717 = ~w5605 & ~w2849;
assign w5718 = ~w2238 & w6842;
assign w5719 = ~w2885 & w2908;
assign w5720 = w2675 & ~w2910;
assign w5721 = ~w2477 & ~w2529;
assign w5722 = ~w2885 & w2947;
assign w5723 = ~w2382 & w2882;
assign w5724 = w2382 & w2882;
assign w5725 = ~w2382 & w2885;
assign w5726 = w2461 & w2882;
assign w5727 = w3000 & w871;
assign w5728 = ~w3000 & ~w871;
assign w5729 = w2997 & ~w2996;
assign w5730 = w1819 & w6843;
assign w5731 = ~w2997 & w2996;
assign w5732 = w2954 & ~w2940;
assign w5733 = ~w2800 & ~w3074;
assign w5734 = w3087 & ~w3069;
assign w5735 = ~w2238 & w6844;
assign w5736 = ~w2238 & w6845;
assign w5737 = (~w3177 & w2238) | (~w3177 & w6846) | (w2238 & w6846);
assign w5738 = ~w2238 & w6847;
assign w5739 = ~w3182 & w3189;
assign w5740 = ~w3182 & w3201;
assign w5741 = ~w3182 & ~w3188;
assign w5742 = ~w2868 & w3187;
assign w5743 = ~w3367 & w3355;
assign w5744 = ~w2430 & w3418;
assign w5745 = w3416 & w6968;
assign w5746 = ~w3416 & w565;
assign w5747 = w3090 & ~w2918;
assign w5748 = (~w3487 & ~w3095) | (~w3487 & w6848) | (~w3095 & w6848);
assign w5749 = ~w3459 & ~w3455;
assign w5750 = w3449 & ~w3450;
assign w5751 = ~w2410 & w6849;
assign w5752 = (w565 & w2410) | (w565 & w6850) | (w2410 & w6850);
assign w5753 = (w2564 & w2410) | (w2564 & w6851) | (w2410 & w6851);
assign w5754 = ~w3489 & ~w3491;
assign w5755 = ~w3594 & ~w3683;
assign w5756 = w3685 & ~w3760;
assign w5757 = ~w3557 & w6852;
assign w5758 = ~w2382 & w1994;
assign w5759 = w2382 & w1994;
assign w5760 = ~w3898 & ~w3896;
assign w5761 = w3862 & w4022;
assign w5762 = ~w3947 & w4100;
assign w5763 = w3986 & ~w4105;
assign w5764 = ~w3947 & ~w4100;
assign w5765 = (w4279 & ~w4275) | (w4279 & w6853) | (~w4275 & w6853);
assign w5766 = w4275 & w6854;
assign w5767 = w4298 & w6855;
assign w5768 = (~w4388 & ~w4298) | (~w4388 & w6856) | (~w4298 & w6856);
assign w5769 = w4295 & ~w4283;
assign w5770 = (~w4277 & ~w4275) | (~w4277 & w6857) | (~w4275 & w6857);
assign w5771 = w4275 & w6858;
assign w5772 = w4448 & w4447;
assign w5773 = ~w4448 & ~w4447;
assign w5774 = ~w1994 & w4544;
assign w5775 = w1994 & ~w1022;
assign w5776 = (~w4374 & w6859) | (~w4374 & w6860) | (w6859 & w6860);
assign w5777 = ~w4583 & ~w4515;
assign w5778 = ~w4494 & w4673;
assign w5779 = ~w4673 & ~w4672;
assign w5780 = (~w4672 & w5779) | (~w4672 & w4494) | (w5779 & w4494);
assign w5781 = ~w4673 & w4688;
assign w5782 = (w4688 & w5781) | (w4688 & w4494) | (w5781 & w4494);
assign w5783 = w5655 & w4711;
assign w5784 = (w4711 & w5655) | (w4711 & w4494) | (w5655 & w4494);
assign w5785 = ~w4712 & w4780;
assign w5786 = w4712 & w4782;
assign w5787 = ~w4712 & w4785;
assign w5788 = w4712 & w4787;
assign w5789 = w4692 & w4790;
assign w5790 = ~w4692 & ~w4790;
assign w5791 = ~w4803 & w4789;
assign w5792 = w4803 & ~w4865;
assign w5793 = ~w4796 & ~w4874;
assign w5794 = w4930 & w6861;
assign w5795 = ~w4930 & w4942;
assign w5796 = ~w4866 & ~w4949;
assign w5797 = ~w4948 & w7787;
assign w5798 = (w4807 & w6862) | (w4807 & w6863) | (w6862 & w6863);
assign w5799 = w4954 & ~w5020;
assign w5800 = ~w4947 & w5010;
assign w5801 = (~w6756 & w5829) | (~w6756 & w7343) | (w5829 & w7343);
assign w5802 = (~w5071 & ~w4674) | (~w5071 & w5829) | (~w4674 & w5829);
assign w5803 = (w6756 & w5830) | (w6756 & w7344) | (w5830 & w7344);
assign w5804 = w4674 & w5830;
assign w5805 = (~w5074 & w5831) | (~w5074 & w5030) | (w5831 & w5030);
assign w5806 = (w5138 & w5012) | (w5138 & w6864) | (w5012 & w6864);
assign w5807 = ~w4964 & w5030;
assign w5808 = ~w5077 & ~w5142;
assign w5809 = ~w5191 & ~w5190;
assign w5810 = w5134 & ~w5195;
assign w5811 = ~w5134 & w5195;
assign w5812 = w5250 & w5287;
assign w5813 = ~w5250 & ~w5287;
assign w5814 = w5294 & w5316;
assign w5815 = w5387 & w5403;
assign w5816 = ~w5387 & ~w5403;
assign w5817 = (~w5137 & w7735) | (~w5137 & w7736) | (w7735 & w7736);
assign w5818 = (~w5414 & w5403) | (~w5414 & w5817) | (w5403 & w5817);
assign w5819 = (w5137 & w7737) | (w5137 & w7738) | (w7737 & w7738);
assign w5820 = ~w5403 & w5819;
assign w5821 = (w5388 & w7345) | (w5388 & w7494) | (w7345 & w7494);
assign w5822 = ~w1710 & w6865;
assign w5823 = w4449 & ~w4450;
assign w5824 = ~w4490 & w4594;
assign w5825 = w4490 & ~w4594;
assign w5826 = ~w5110 & ~w5111;
assign w5827 = ~w5212 & w5214;
assign w5828 = w5385 & w6866;
assign w5829 = ~w5032 & w7788;
assign w5830 = w5071 & ~w5034;
assign w5831 = ~w5005 & ~w5074;
assign w5832 = w4586 & w4450;
assign w5833 = w4586 & ~w5650;
assign w5834 = ~w4930 & ~w4929;
assign w5835 = w5001 & ~w4927;
assign w5836 = ~w4931 & w5835;
assign w5837 = w5003 & w4927;
assign w5838 = (w5003 & w4931) | (w5003 & w5837) | (w4931 & w5837);
assign w5839 = w5006 & ~w4927;
assign w5840 = ~w4931 & w5839;
assign w5841 = w5008 & w4927;
assign w5842 = (w5008 & w4931) | (w5008 & w5841) | (w4931 & w5841);
assign w5843 = w5178 & ~w5151;
assign w5844 = w5180 & w5151;
assign w5845 = ~w5166 & ~w5151;
assign w5846 = (w5035 & w6871) | (w5035 & w6872) | (w6871 & w6872);
assign w5847 = ~w5186 & ~w5182;
assign w5848 = (w3829 & w5198) | (w3829 & w6454) | (w5198 & w6454);
assign w5849 = (w5242 & w6873) | (w5242 & w6874) | (w6873 & w6874);
assign w5850 = (~w5242 & w6875) | (~w5242 & w6876) | (w6875 & w6876);
assign w5851 = ~w5333 & w5139;
assign w5852 = w5139 & w5339;
assign w5853 = w5250 & w5345;
assign w5854 = w5366 & w5365;
assign w5855 = ~w5366 & ~w5365;
assign w5856 = ~w5370 & ~w5661;
assign w5857 = (w7347 & w5243) | (w7347 & w7639) | (w5243 & w7639);
assign w5858 = (~w5243 & w7640) | (~w5243 & w7641) | (w7640 & w7641);
assign w5859 = (~w4940 & ~w4930) | (~w4940 & w6877) | (~w4930 & w6877);
assign w5860 = w388 & a_3;
assign w5861 = ~w388 & ~a_3;
assign w5862 = w96 & ~w139;
assign w5863 = w65 & ~w86;
assign w5864 = ~w395 & ~w461;
assign w5865 = (~a_22 & ~w6) | (~a_22 & w6878) | (~w6 & w6878);
assign w5866 = a_10 & ~a_22;
assign w5867 = ~a_22 & w7789;
assign w5868 = ~w7276 & w6879;
assign w5869 = a_12 & w5867;
assign w5870 = a_22 & a_4;
assign w5871 = ~a_22 & ~a_4;
assign w5872 = w428 & w574;
assign w5873 = ~w428 & ~w574;
assign w5874 = ~w428 & w391;
assign w5875 = w391 & ~w582;
assign w5876 = a_7 & ~a_22;
assign w5877 = a_8 & ~a_22;
assign w5878 = a_4 & ~a_22;
assign w5879 = ~w843 & a_22;
assign w5880 = ~w843 & ~w5878;
assign w5881 = ~a_22 & ~a_7;
assign w5882 = a_22 & a_7;
assign w5883 = (~w854 & ~w828) | (~w854 & w6880) | (~w828 & w6880);
assign w5884 = a_5 & a_22;
assign w5885 = a_5 & ~w5878;
assign w5886 = w428 & ~w871;
assign w5887 = ~w428 & w871;
assign w5888 = a_22 & ~a_13;
assign w5889 = ~a_22 & a_13;
assign w5890 = ~w1017 & ~w901;
assign w5891 = ~a_14 & w5889;
assign w5892 = ~w5888 & w6881;
assign w5893 = a_14 & ~w5889;
assign w5894 = (a_14 & w5888) | (a_14 & w6882) | (w5888 & w6882);
assign w5895 = w917 & w391;
assign w5896 = w428 & w847;
assign w5897 = ~w428 & ~w847;
assign w5898 = w917 & ~w574;
assign w5899 = ~w920 & ~w1180;
assign w5900 = w1119 & w1189;
assign w5901 = ~w1119 & ~w1189;
assign w5902 = ~w1131 & w1193;
assign w5903 = w1131 & ~w1193;
assign w5904 = w428 & w854;
assign w5905 = ~w428 & ~w854;
assign w5906 = w1289 & ~w1285;
assign w5907 = w428 & ~w726;
assign w5908 = ~w428 & w726;
assign w5909 = ~w455 & ~w726;
assign w5910 = ~w726 & ~w1338;
assign w5911 = w1342 & w1140;
assign w5912 = ~w1342 & ~w1140;
assign w5913 = w1360 & w1346;
assign w5914 = ~w1360 & ~w1346;
assign w5915 = w720 & ~w974;
assign w5916 = w1371 & w1370;
assign w5917 = ~w1371 & ~w1370;
assign w5918 = (~w871 & ~w837) | (~w871 & w6883) | (~w837 & w6883);
assign w5919 = w837 & w6884;
assign w5920 = ~w455 & ~w847;
assign w5921 = w1340 & ~w1392;
assign w5922 = w1394 & w1393;
assign w5923 = ~w847 & ~w1391;
assign w5924 = ~w1394 & ~w1393;
assign w5925 = ~w455 & w574;
assign w5926 = (w391 & ~w560) | (w391 & w6885) | (~w560 & w6885);
assign w5927 = ~w5926 & ~w1424;
assign w5928 = w1428 & ~w1420;
assign w5929 = ~w1437 & ~w1389;
assign w5930 = w383 & w391;
assign w5931 = ~w1484 & ~w1480;
assign w5932 = ~w1502 & ~w1535;
assign w5933 = ~w1251 & ~w1535;
assign w5934 = w1539 & ~w1538;
assign w5935 = ~w365 & ~w265;
assign w5936 = w1502 & w1535;
assign w5937 = w1502 & ~w1331;
assign w5938 = ~w1593 & ~w1591;
assign w5939 = w428 & w720;
assign w5940 = ~w428 & ~w720;
assign w5941 = w1284 & ~w1640;
assign w5942 = w1323 & ~w1648;
assign w5943 = ~w1323 & w1648;
assign w5944 = ~w437 & w1658;
assign w5945 = w1539 & w1707;
assign w5946 = ~w1502 & w1657;
assign w5947 = w1641 & ~w1642;
assign w5948 = ~w428 & ~w735;
assign w5949 = ~w720 & ~w1616;
assign w5950 = w917 & ~w854;
assign w5951 = w1649 & ~w1650;
assign w5952 = ~w1255 & ~w1655;
assign w5953 = w428 & w565;
assign w5954 = ~w428 & ~w565;
assign w5955 = w917 & w726;
assign w5956 = w1908 & w1907;
assign w5957 = w1786 & w1930;
assign w5958 = w1939 & ~w1938;
assign w5959 = w1939 & ~w1825;
assign w5960 = w1839 & w1949;
assign w5961 = ~w1839 & ~w1949;
assign w5962 = ~w1820 & w1963;
assign w5963 = w1022 & ~w565;
assign w5964 = w1982 & ~w1022;
assign w5965 = w1959 & w565;
assign w5966 = w428 & ~w511;
assign w5967 = ~w428 & w511;
assign w5968 = w565 & ~w1870;
assign w5969 = w917 & ~w720;
assign w5970 = ~w2112 & ~w2118;
assign w5971 = w917 & w735;
assign w5972 = w2083 & ~w2073;
assign w5973 = w428 & ~w880;
assign w5974 = ~w428 & w880;
assign w5975 = w696 & w6886;
assign w5976 = w1839 & w2245;
assign w5977 = ~w383 & ~w1877;
assign w5978 = w383 & w1877;
assign w5979 = w2148 & ~w2139;
assign w5980 = w917 & w565;
assign w5981 = ~w920 & ~w2260;
assign w5982 = ~w428 & w1022;
assign w5983 = w428 & ~w1022;
assign w5984 = ~w2272 & w2266;
assign w5985 = w2272 & ~w2266;
assign w5986 = ~w2162 & w2286;
assign w5987 = w2334 & ~w2287;
assign w5988 = w2334 & w5553;
assign w5989 = w1722 & w2334;
assign w5990 = ~w2246 & w2381;
assign w5991 = ~w2246 & w2405;
assign w5992 = ~w2402 & ~w2406;
assign w5993 = w2385 & w2415;
assign w5994 = ~w2246 & w2402;
assign w5995 = w2247 & ~w2382;
assign w5996 = w2422 & ~w2436;
assign w5997 = w511 & w565;
assign w5998 = ~w6000 & ~w2002;
assign w5999 = w2041 & w2451;
assign w6000 = ~w1710 & w6887;
assign w6001 = ~w2041 & w2464;
assign w6002 = w2041 & ~w2464;
assign w6003 = ~w1820 & w2405;
assign w6004 = ~w2402 & ~w2470;
assign w6005 = (~w2402 & w1710) | (~w2402 & w6888) | (w1710 & w6888);
assign w6006 = ~w1820 & w2436;
assign w6007 = ~w1820 & w2402;
assign w6008 = ~w2525 & ~w2529;
assign w6009 = (w1715 & w6889) | (w1715 & w6890) | (w6889 & w6890);
assign w6010 = ~w1839 & ~w2556;
assign w6011 = w1839 & ~w2558;
assign w6012 = ~w2278 & ~w2257;
assign w6013 = w384 & w6891;
assign w6014 = (~w2124 & ~w384) | (~w2124 & w6892) | (~w384 & w6892);
assign w6015 = w917 & w511;
assign w6016 = ~w2078 & ~w2251;
assign w6017 = ~w2275 & ~w2273;
assign w6018 = w2586 & ~w2640;
assign w6019 = ~w2640 & w2589;
assign w6020 = ~w2640 & w5587;
assign w6021 = ~w2648 & w6893;
assign w6022 = w2649 & ~w5589;
assign w6023 = ~w2652 & ~w2653;
assign w6024 = ~w2652 & ~w5590;
assign w6025 = (w2398 & w2410) | (w2398 & w6894) | (w2410 & w6894);
assign w6026 = ~w2410 & w6895;
assign w6027 = (~w726 & w2410) | (~w726 & w6896) | (w2410 & w6896);
assign w6028 = (~w2606 & w2608) | (~w2606 & w7349) | (w2608 & w7349);
assign w6029 = ~w2603 & ~w2594;
assign w6030 = w917 & w880;
assign w6031 = ~w2683 & ~w2682;
assign w6032 = w432 & ~w2124;
assign w6033 = ~w1721 & w6897;
assign w6034 = ~w2590 & ~w2709;
assign w6035 = ~w1721 & w6898;
assign w6036 = w2696 & ~w2695;
assign w6037 = ~w2729 & ~w2727;
assign w6038 = w2728 & w2726;
assign w6039 = ~w2728 & ~w2726;
assign w6040 = (~w2734 & w2677) | (~w2734 & w6900) | (w2677 & w6900);
assign w6041 = ~w2590 & w2709;
assign w6042 = ~w2811 & ~w2804;
assign w6043 = w2724 & ~w2763;
assign w6044 = ~w2731 & w2734;
assign w6045 = ~w2844 & ~w2734;
assign w6046 = (~w2844 & w2677) | (~w2844 & w6902) | (w2677 & w6902);
assign w6047 = ~w2815 & w2853;
assign w6048 = w2815 & w2852;
assign w6049 = ~w2811 & w2857;
assign w6050 = ~w2872 & ~w2870;
assign w6051 = a_22 & a_2;
assign w6052 = ~a_22 & ~a_2;
assign w6053 = ~w2898 & w6903;
assign w6054 = w2904 & w871;
assign w6055 = ~w2904 & ~w871;
assign w6056 = ~w2885 & w2937;
assign w6057 = ~w2655 & w6904;
assign w6058 = (~w871 & w2655) | (~w871 & w6905) | (w2655 & w6905);
assign w6059 = ~w2246 & w2891;
assign w6060 = ~w2893 & ~w2955;
assign w6061 = (w871 & ~w2881) | (w871 & w6906) | (~w2881 & w6906);
assign w6062 = ~w6061 & ~w2882;
assign w6063 = w2385 & w2957;
assign w6064 = ~w2246 & w2893;
assign w6065 = w2978 & w871;
assign w6066 = ~w2978 & ~w871;
assign w6067 = ~w2972 & ~w2991;
assign w6068 = ~w1820 & w2891;
assign w6069 = ~w2246 & w2903;
assign w6070 = ~w2893 & ~w2999;
assign w6071 = (~w2893 & w1710) | (~w2893 & w6907) | (w1710 & w6907);
assign w6072 = (~w1715 & w6908) | (~w1715 & w6909) | (w6908 & w6909);
assign w6073 = ~w1820 & w3009;
assign w6074 = ~w1820 & w2893;
assign w6075 = (~w3074 & w5733) | (~w3074 & w2661) | (w5733 & w2661);
assign w6076 = (~w3074 & w5733) | (~w3074 & w2583) | (w5733 & w2583);
assign w6077 = w2788 & w6910;
assign w6078 = (~w871 & ~w2788) | (~w871 & w6911) | (~w2788 & w6911);
assign w6079 = ~w2885 & w3085;
assign w6080 = w2835 & w3111;
assign w6081 = ~w252 & ~w164;
assign w6082 = w3142 & w3112;
assign w6083 = ~w2896 & w3143;
assign w6084 = w3144 & w3148;
assign w6085 = a_1 & ~a_2;
assign w6086 = ~a_1 & a_2;
assign w6087 = w3145 & w3173;
assign w6088 = ~w2835 & ~w3111;
assign w6089 = ~w3142 & w3111;
assign w6090 = ~w2896 & w6912;
assign w6091 = w3142 & ~w3111;
assign w6092 = (w3142 & w2896) | (w3142 & w6913) | (w2896 & w6913);
assign w6093 = ~w2896 & w6914;
assign w6094 = (~w3161 & w2896) | (~w3161 & w6915) | (w2896 & w6915);
assign w6095 = ~w3197 & ~w3189;
assign w6096 = ~w3197 & w2803;
assign w6097 = ~w3195 & w3192;
assign w6098 = (~w3200 & w3188) | (~w3200 & w6916) | (w3188 & w6916);
assign w6099 = ~w3200 & w2803;
assign w6100 = ~w3149 & ~w3174;
assign w6101 = ~w0 & ~w2878;
assign w6102 = ~w2898 & w6918;
assign w6103 = w3225 & w6919;
assign w6104 = (~w2878 & ~w3225) | (~w2878 & w6920) | (~w3225 & w6920);
assign w6105 = ~w2878 & ~w6103;
assign w6106 = w2967 & ~w3063;
assign w6107 = w3006 & ~w3058;
assign w6108 = ~w847 & w871;
assign w6109 = ~w2246 & w3148;
assign w6110 = ~w2878 & ~w3273;
assign w6111 = (~w2878 & ~w3273) | (~w2878 & w7620) | (~w3273 & w7620);
assign w6112 = (w3269 & w7642) | (w3269 & w7643) | (w7642 & w7643);
assign w6113 = ~w2246 & w3169;
assign w6114 = ~w1820 & w3173;
assign w6115 = w2461 & w3175;
assign w6116 = ~w3148 & ~w3277;
assign w6117 = ~w3280 & ~w2878;
assign w6118 = w3280 & w2878;
assign w6119 = (w1715 & w6924) | (w1715 & w6925) | (w6924 & w6925);
assign w6120 = ~w3024 & w3284;
assign w6121 = w3024 & ~w3284;
assign w6122 = w1715 & w6926;
assign w6123 = ~w1820 & w3169;
assign w6124 = ~w3175 & w3295;
assign w6125 = ~a_0 & ~w0;
assign w6126 = w1710 & w6927;
assign w6127 = (w2878 & w3305) | (w2878 & w6928) | (w3305 & w6928);
assign w6128 = ~w1820 & w3148;
assign w6129 = ~w3311 & w6929;
assign w6130 = ~w3311 & w6930;
assign w6131 = ~w2878 & w6129;
assign w6132 = ~w3318 & ~w3310;
assign w6133 = ~w2246 & w3173;
assign w6134 = (w3175 & w2384) | (w3175 & w6931) | (w2384 & w6931);
assign w6135 = ~w3148 & ~w3322;
assign w6136 = (~w2878 & ~w3323) | (~w2878 & w7393) | (~w3323 & w7393);
assign w6137 = w3323 & w6932;
assign w6138 = ~w3266 & w7790;
assign w6139 = w3259 & ~w3334;
assign w6140 = ~w3220 & ~w3248;
assign w6141 = w3144 & w3169;
assign w6142 = w3145 & w3148;
assign w6143 = ~w2898 & w6933;
assign w6144 = w3352 & w6934;
assign w6145 = w3352 & w6935;
assign w6146 = w3145 & w3169;
assign w6147 = ~w2898 & w6936;
assign w6148 = w3180 & w3186;
assign w6149 = (w3180 & w2868) | (w3180 & w6148) | (w2868 & w6148);
assign w6150 = ~w3343 & ~w3357;
assign w6151 = w3375 & ~w3342;
assign w6152 = w3367 & ~w3355;
assign w6153 = ~w2898 & w6937;
assign w6154 = w3145 & w2903;
assign w6155 = w871 & w3391;
assign w6156 = w3391 & w6838;
assign w6157 = ~w2396 & w3404;
assign w6158 = ~w2246 & w1976;
assign w6159 = ~w1820 & w1987;
assign w6160 = w3409 & w3442;
assign w6161 = ~w3409 & ~w3442;
assign w6162 = ~w2900 & w7351;
assign w6163 = (~w3471 & w2900) | (~w3471 & w7352) | (w2900 & w7352);
assign w6164 = w3144 & w3173;
assign w6165 = w3477 & w3480;
assign w6166 = ~w3477 & ~w3480;
assign w6167 = ~w1820 & w1991;
assign w6168 = ~w3499 & w3495;
assign w6169 = w3499 & ~w3495;
assign w6170 = ~w1994 & ~w3502;
assign w6171 = ~w2246 & w1974;
assign w6172 = ~w1976 & ~w3512;
assign w6173 = w2788 & w6895;
assign w6174 = (~w726 & ~w2788) | (~w726 & w6896) | (~w2788 & w6896);
assign w6175 = ~w2396 & w3536;
assign w6176 = (w3552 & w2900) | (w3552 & w7354) | (w2900 & w7354);
assign w6177 = ~w3471 & ~w3554;
assign w6178 = w3196 & w3556;
assign w6179 = w3557 & ~w3189;
assign w6180 = w3557 & w2803;
assign w6181 = w3559 & w3142;
assign w6182 = ~w2896 & w6939;
assign w6183 = (w3169 & ~w3550) | (w3169 & w6940) | (~w3550 & w6940);
assign w6184 = w3145 & w2893;
assign w6185 = w3144 & w2903;
assign w6186 = ~w2898 & w6942;
assign w6187 = w3578 & w871;
assign w6188 = ~w3578 & ~w871;
assign w6189 = ~w2885 & w3582;
assign w6190 = w3573 & w3584;
assign w6191 = w3607 & w3613;
assign w6192 = w3601 & w3614;
assign w6193 = ~w3643 & w3385;
assign w6194 = ~w187 & w1907;
assign w6195 = ~w3207 & w3385;
assign w6196 = w3144 & w2893;
assign w6197 = w3145 & w2891;
assign w6198 = ~w3699 & ~w3700;
assign w6199 = ~w2898 & w6943;
assign w6200 = ~w3709 & ~w726;
assign w6201 = w3709 & w726;
assign w6202 = ~w2396 & w3713;
assign w6203 = w3501 & w6944;
assign w6204 = ~w1820 & w2546;
assign w6205 = ~w2246 & w1987;
assign w6206 = ~w1991 & ~w3726;
assign w6207 = ~w2410 & w6945;
assign w6208 = (~w565 & w2410) | (~w565 & w6946) | (w2410 & w6946);
assign w6209 = (~w2564 & w2410) | (~w2564 & w6947) | (w2410 & w6947);
assign w6210 = ~w608 & w3169;
assign w6211 = ~w3551 & ~w3780;
assign w6212 = w3551 & w3780;
assign w6213 = ~w3786 & ~w3784;
assign w6214 = ~w3173 & ~w3781;
assign w6215 = (w6950 & w6951) | (w6950 & w7767) | (w6951 & w7767);
assign w6216 = (w3790 & w7357) | (w3790 & w7358) | (w7357 & w7358);
assign w6217 = (w3715 & w3529) | (w3715 & w6594) | (w3529 & w6594);
assign w6218 = (w565 & ~w3869) | (w565 & w6952) | (~w3869 & w6952);
assign w6219 = w3869 & w6953;
assign w6220 = w1820 & ~w1022;
assign w6221 = ~w2246 & w1991;
assign w6222 = ~w3886 & ~w3882;
assign w6223 = w3886 & w3882;
assign w6224 = w3145 & w2411;
assign w6225 = ~w2898 & w6954;
assign w6226 = w3905 & w6955;
assign w6227 = w3905 & w6956;
assign w6228 = w3144 & w2891;
assign w6229 = (~w871 & ~w3917) | (~w871 & w6957) | (~w3917 & w6957);
assign w6230 = (~w871 & ~w3917) | (~w871 & w7359) | (~w3917 & w7359);
assign w6231 = w3551 & w3936;
assign w6232 = ~w3551 & ~w3936;
assign w6233 = ~w3782 & ~w3939;
assign w6234 = w3782 & w3939;
assign w6235 = ~w608 & w3148;
assign w6236 = (w3173 & ~w3550) | (w3173 & w6958) | (~w3550 & w6958);
assign w6237 = ~w3943 & w6959;
assign w6238 = (w3472 & w6960) | (w3472 & w6961) | (w6960 & w6961);
assign w6239 = ~w3831 & w3962;
assign w6240 = w3831 & ~w3962;
assign w6241 = w3829 & w3965;
assign w6242 = ~w1820 & ~w1022;
assign w6243 = w3886 & w3999;
assign w6244 = w2367 & w1994;
assign w6245 = ~w2246 & w2546;
assign w6246 = ~w1991 & ~w4009;
assign w6247 = w3145 & w2402;
assign w6248 = w3144 & w2411;
assign w6249 = ~w2898 & w6963;
assign w6250 = w4040 & ~w726;
assign w6251 = ~w4040 & w726;
assign w6252 = ~w2394 & w4044;
assign w6253 = (w2903 & ~w3550) | (w2903 & w6964) | (~w3550 & w6964);
assign w6254 = ~w3474 & w6910;
assign w6255 = (~w871 & w3474) | (~w871 & w6911) | (w3474 & w6911);
assign w6256 = (w4055 & w7360) | (w4055 & w7361) | (w7360 & w7361);
assign w6257 = (~w3175 & w3936) | (~w3175 & w7505) | (w3936 & w7505);
assign w6258 = (w3829 & w3969) | (w3829 & w3830) | (w3969 & w3830);
assign w6259 = ~w2898 & w6966;
assign w6260 = w4153 & w6967;
assign w6261 = w4153 & w7362;
assign w6262 = (w565 & ~w4153) | (w565 & w6969) | (~w4153 & w6969);
assign w6263 = (~w4153 & w7363) | (~w4153 & w7364) | (w7363 & w7364);
assign w6264 = w2246 & ~w1022;
assign w6265 = ~w2655 & w6971;
assign w6266 = (~w4164 & w2655) | (~w4164 & w6972) | (w2655 & w6972);
assign w6267 = w3145 & w2405;
assign w6268 = w3144 & w2402;
assign w6269 = ~w4183 & ~w4184;
assign w6270 = (w2893 & ~w3550) | (w2893 & w6973) | (~w3550 & w6973);
assign w6271 = ~w608 & w2903;
assign w6272 = ~w6270 & ~w4200;
assign w6273 = ~w6232 & w3780;
assign w6274 = w3936 & w3780;
assign w6275 = (w2878 & w3936) | (w2878 & w6976) | (w3936 & w6976);
assign w6276 = (~w3553 & w6977) | (~w3553 & w6978) | (w6977 & w6978);
assign w6277 = (w3553 & w6979) | (w3553 & w6980) | (w6979 & w6980);
assign w6278 = ~w3898 & w5638;
assign w6279 = w4052 & ~w4220;
assign w6280 = ~w2246 & ~w1022;
assign w6281 = (w4264 & w2655) | (w4264 & w6981) | (w2655 & w6981);
assign w6282 = w1022 & ~w2878;
assign w6283 = ~w1022 & w2878;
assign w6284 = w3145 & w1968;
assign w6285 = ~w2898 & w6982;
assign w6286 = w4290 & ~w3187;
assign w6287 = w4290 & ~w5742;
assign w6288 = (~w565 & ~w4289) | (~w565 & w6983) | (~w4289 & w6983);
assign w6289 = w4289 & w6984;
assign w6290 = w3144 & w2405;
assign w6291 = ~w3474 & w6985;
assign w6292 = (w726 & w3474) | (w726 & w6986) | (w3474 & w6986);
assign w6293 = ~w2394 & w4305;
assign w6294 = (w3472 & w6987) | (w3472 & w6988) | (w6987 & w6988);
assign w6295 = ~w608 & w2893;
assign w6296 = (w2891 & ~w3550) | (w2891 & w6989) | (~w3550 & w6989);
assign w6297 = ~w4315 & w6991;
assign w6298 = (~w3788 & w7367) | (~w3788 & w7368) | (w7367 & w7368);
assign w6299 = (w3788 & w7369) | (w3788 & w7370) | (w7369 & w7370);
assign w6300 = w4224 & ~w4348;
assign w6301 = ~w608 & w2891;
assign w6302 = w4382 & ~w871;
assign w6303 = ~w4382 & w871;
assign w6304 = ~w2882 & ~w4384;
assign w6305 = w4396 & w6995;
assign w6306 = w4396 & w6996;
assign w6307 = w1022 & w2878;
assign w6308 = ~w1022 & ~w2878;
assign w6309 = ~w6283 & ~w1022;
assign w6310 = w4275 & w6997;
assign w6311 = ~w4404 & w4277;
assign w6312 = w2788 & w6998;
assign w6313 = (~w1022 & ~w2788) | (~w1022 & w6999) | (~w2788 & w6999);
assign w6314 = ~w1994 & w4421;
assign w6315 = w3145 & w1976;
assign w6316 = w3144 & w1968;
assign w6317 = ~w2898 & w7000;
assign w6318 = w4432 & ~w565;
assign w6319 = ~w4432 & w565;
assign w6320 = ~w4429 & w4436;
assign w6321 = ~w4444 & ~w4390;
assign w6322 = ~w2891 & ~w3009;
assign w6323 = (~w3553 & w7002) | (~w3553 & w7003) | (w7002 & w7003);
assign w6324 = ~w3936 & w871;
assign w6325 = w3936 & ~w871;
assign w6326 = ~w4393 & w7004;
assign w6327 = (w4520 & w4393) | (w4520 & w7005) | (w4393 & w7005);
assign w6328 = ~w4276 & w4531;
assign w6329 = w4276 & w4535;
assign w6330 = ~w2898 & w7006;
assign w6331 = w4540 & w1022;
assign w6332 = ~w4540 & ~w1022;
assign w6333 = w3144 & w1976;
assign w6334 = w3145 & w1974;
assign w6335 = ~w4429 & w4557;
assign w6336 = (w2402 & ~w3550) | (w2402 & w7007) | (~w3550 & w7007);
assign w6337 = ~w608 & w2411;
assign w6338 = ~w6336 & ~w4568;
assign w6339 = ~w608 & w2402;
assign w6340 = (w2405 & ~w3550) | (w2405 & w7009) | (~w3550 & w7009);
assign w6341 = ~w4608 & w7010;
assign w6342 = ~w4608 & w7011;
assign w6343 = w726 & w6341;
assign w6344 = ~w2394 & w4612;
assign w6345 = w4559 & ~w4548;
assign w6346 = w3145 & w1987;
assign w6347 = ~w2898 & w7012;
assign w6348 = ~w4624 & ~w1994;
assign w6349 = w4626 & ~w3187;
assign w6350 = w4626 & ~w5742;
assign w6351 = w4632 & ~w1022;
assign w6352 = ~w4627 & ~w4637;
assign w6353 = w4627 & w4637;
assign w6354 = w4526 & ~w4525;
assign w6355 = w3144 & w1974;
assign w6356 = ~w3474 & w6849;
assign w6357 = (w565 & w3474) | (w565 & w6850) | (w3474 & w6850);
assign w6358 = ~w4429 & w4651;
assign w6359 = w4522 & ~w4523;
assign w6360 = (~w4686 & ~w4578) | (~w4686 & w7013) | (~w4578 & w7013);
assign w6361 = w4692 & ~w4590;
assign w6362 = ~w4579 & ~w4664;
assign w6363 = w4659 & ~w4616;
assign w6364 = (w1968 & ~w3550) | (w1968 & w7014) | (~w3550 & w7014);
assign w6365 = ~w3474 & w7015;
assign w6366 = (w565 & w3474) | (w565 & w7016) | (w3474 & w7016);
assign w6367 = ~w4429 & w4722;
assign w6368 = ~w6351 & ~w4631;
assign w6369 = w3144 & w1987;
assign w6370 = w3145 & w1991;
assign w6371 = ~w2898 & w7017;
assign w6372 = w4733 & w7018;
assign w6373 = ~w4729 & w4734;
assign w6374 = ~w4729 & w6372;
assign w6375 = (w4741 & ~w4625) | (w4741 & w7019) | (~w4625 & w7019);
assign w6376 = w4625 & w7020;
assign w6377 = ~w608 & w2405;
assign w6378 = ~w4749 & w7021;
assign w6379 = (w726 & w4749) | (w726 & w7022) | (w4749 & w7022);
assign w6380 = w726 & ~w6378;
assign w6381 = w4621 & ~w4654;
assign w6382 = ~w4808 & ~w4762;
assign w6383 = ~w4745 & ~w4738;
assign w6384 = ~w2405 & ~w2436;
assign w6385 = (~w3553 & w7024) | (~w3553 & w7025) | (w7024 & w7025);
assign w6386 = ~w3936 & ~w726;
assign w6387 = w3936 & w726;
assign w6388 = w3145 & w2546;
assign w6389 = w3144 & w1991;
assign w6390 = ~w4822 & ~w4823;
assign w6391 = w4733 & w7026;
assign w6392 = w4733 & w7027;
assign w6393 = (w1976 & ~w3550) | (w1976 & w7028) | (~w3550 & w7028);
assign w6394 = ~w608 & w1968;
assign w6395 = ~w6393 & ~w4835;
assign w6396 = (~w4757 & w4748) | (~w4757 & w7030) | (w4748 & w7030);
assign w6397 = w3829 & ~w4878;
assign w6398 = ~w3829 & w4878;
assign w6399 = ~w4761 & w7031;
assign w6400 = w3145 & ~w1022;
assign w6401 = ~w4894 & w4898;
assign w6402 = ~w6401 & ~w4897;
assign w6403 = w3144 & w2546;
assign w6404 = ~w4896 & w4907;
assign w6405 = w4896 & ~w4907;
assign w6406 = w4839 & ~w4832;
assign w6407 = ~w608 & w1976;
assign w6408 = (w1974 & ~w3550) | (w1974 & w7033) | (~w3550 & w7033);
assign w6409 = ~w4913 & w7034;
assign w6410 = ~w4913 & w7035;
assign w6411 = w565 & w6409;
assign w6412 = ~w4429 & w4917;
assign w6413 = w4842 & ~w4817;
assign w6414 = w4847 & ~w4848;
assign w6415 = w4878 & w3829;
assign w6416 = ~w4910 & ~w4920;
assign w6417 = w3144 & ~w1022;
assign w6418 = (w4890 & w4886) | (w4890 & w7036) | (w4886 & w7036);
assign w6419 = ~w1022 & w7791;
assign w6420 = (w1987 & ~w3550) | (w1987 & w7037) | (~w3550 & w7037);
assign w6421 = w4977 & w7038;
assign w6422 = ~w4973 & w4978;
assign w6423 = ~w4973 & w6421;
assign w6424 = ~w608 & w1974;
assign w6425 = ~w4982 & w7039;
assign w6426 = ~w4982 & w7040;
assign w6427 = ~w565 & w6425;
assign w6428 = ~w4944 & ~w4947;
assign w6429 = ~w4964 & w5014;
assign w6430 = w4957 & w3829;
assign w6431 = w4993 & ~w4994;
assign w6432 = ~w1974 & ~w1963;
assign w6433 = (~w3553 & w7042) | (~w3553 & w7043) | (w7042 & w7043);
assign w6434 = ~w3936 & ~w565;
assign w6435 = w3936 & w565;
assign w6436 = ~w608 & w1987;
assign w6437 = ~w2546 & ~w5040;
assign w6438 = ~w4971 & w7880;
assign w6439 = w4970 & w7045;
assign w6440 = (w5048 & ~w4970) | (w5048 & w7046) | (~w4970 & w7046);
assign w6441 = w5024 & w3829;
assign w6442 = w5080 & w3829;
assign w6443 = w5080 & w6441;
assign w6444 = ~w5085 & w5048;
assign w6445 = (~w5085 & ~w4970) | (~w5085 & w7047) | (~w4970 & w7047);
assign w6446 = w1022 & w565;
assign w6447 = ~w1022 & ~w565;
assign w6448 = (w2546 & ~w3550) | (w2546 & w7048) | (~w3550 & w7048);
assign w6449 = ~w608 & w1991;
assign w6450 = ~w5095 & w7049;
assign w6451 = (w3472 & w7050) | (w3472 & w7051) | (w7050 & w7051);
assign w6452 = w5139 & ~w5127;
assign w6453 = ~w3829 & ~w5144;
assign w6454 = w3829 & w5144;
assign w6455 = w5057 & ~w5105;
assign w6456 = (w5086 & ~w5098) | (w5086 & w7372) | (~w5098 & w7372);
assign w6457 = (~w1022 & ~w3550) | (~w1022 & w7053) | (~w3550 & w7053);
assign w6458 = ~w5090 & ~w5088;
assign w6459 = ~w608 & w2546;
assign w6460 = ~w5158 & w7054;
assign w6461 = ~w5158 & w7055;
assign w6462 = w1022 & w6460;
assign w6463 = w5157 & w7792;
assign w6464 = (w4071 & w7056) | (w4071 & w7057) | (w7056 & w7057);
assign w6465 = (w3553 & w7058) | (w3553 & w7490) | (w7058 & w7490);
assign w6466 = w2546 & ~w3936;
assign w6467 = (~w3936 & w3784) | (~w3936 & w7059) | (w3784 & w7059);
assign w6468 = (w6466 & w3784) | (w6466 & w7060) | (w3784 & w7060);
assign w6469 = ~w5155 & ~w5204;
assign w6470 = w5155 & w5204;
assign w6471 = w5163 & w5207;
assign w6472 = ~w5163 & ~w5207;
assign w6473 = ~w5164 & w5208;
assign w6474 = w5166 & w5207;
assign w6475 = w631 & w7061;
assign w6476 = ~w5128 & w5182;
assign w6477 = ~w5237 & w5239;
assign w6478 = ~w5166 & w5208;
assign w6479 = w6457 & w3780;
assign w6480 = (~w5264 & w3939) | (~w5264 & w7065) | (w3939 & w7065);
assign w6481 = ~w3939 & w7066;
assign w6482 = (w5151 & w7067) | (w5151 & w7068) | (w7067 & w7068);
assign w6483 = (~w5281 & w5659) | (~w5281 & w5260) | (w5659 & w5260);
assign w6484 = w5253 & w3829;
assign w6485 = ~w5290 & w3829;
assign w6486 = ~w5290 & w6484;
assign w6487 = ~w5294 & w3829;
assign w6488 = (~w5151 & w7647) | (~w5151 & w7648) | (w7647 & w7648);
assign w6489 = (~w7063 & w7373) | (~w7063 & w7374) | (w7373 & w7374);
assign w6490 = (~w5296 & w5220) | (~w5296 & w7375) | (w5220 & w7375);
assign w6491 = (~w5307 & w5284) | (~w5307 & w7074) | (w5284 & w7074);
assign w6492 = ~w5297 & w5308;
assign w6493 = ~w5284 & w7075;
assign w6494 = w5241 & w5660;
assign w6495 = (~w5243 & w7649) | (~w5243 & w7650) | (w7649 & w7650);
assign w6496 = ~w5297 & w5662;
assign w6497 = ~w5232 & w5333;
assign w6498 = w5351 & ~w3829;
assign w6499 = w5351 & ~w5661;
assign w6500 = (~w5243 & w7651) | (~w5243 & w7652) | (w7651 & w7652);
assign w6501 = (w5385 & w5664) | (w5385 & w5297) | (w5664 & w5297);
assign w6502 = w5312 & w5386;
assign w6503 = w5250 & w5387;
assign w6504 = w5362 & w5384;
assign w6505 = ~w5297 & w5665;
assign w6506 = w919 & w915;
assign w6507 = ~w5411 & ~w5420;
assign w6508 = w45 & w47;
assign w6509 = ~w5392 & ~w5417;
assign w6510 = ~w5428 & ~w5426;
assign w6511 = w5428 & ~w5415;
assign w6512 = w819 & w7078;
assign w6513 = (~w726 & ~w819) | (~w726 & w7079) | (~w819 & w7079);
assign w6514 = w819 & w7080;
assign w6515 = w819 & w7081;
assign w6516 = (~w720 & ~w819) | (~w720 & w7082) | (~w819 & w7082);
assign w6517 = w819 & w7083;
assign w6518 = (~w735 & ~w819) | (~w735 & w7084) | (~w819 & w7084);
assign w6519 = w819 & w7085;
assign w6520 = (~w574 & ~w819) | (~w574 & w7086) | (~w819 & w7086);
assign w6521 = (~w565 & ~w819) | (~w565 & w7087) | (~w819 & w7087);
assign w6522 = w819 & w7088;
assign w6523 = w819 & w7089;
assign w6524 = (~w511 & ~w819) | (~w511 & w7090) | (~w819 & w7090);
assign w6525 = (w847 & ~w828) | (w847 & w7091) | (~w828 & w7091);
assign w6526 = w828 & w7092;
assign w6527 = w819 & w7093;
assign w6528 = (w880 & ~w819) | (w880 & w7094) | (~w819 & w7094);
assign w6529 = w1330 & w7095;
assign w6530 = (~w1695 & ~w1330) | (~w1695 & w7096) | (~w1330 & w7096);
assign w6531 = w819 & w7097;
assign w6532 = (w1022 & ~w819) | (w1022 & w7098) | (~w819 & w7098);
assign w6533 = ~w1991 & ~w1987;
assign w6534 = ~w1974 & ~w1976;
assign w6535 = ~w1976 & ~w1968;
assign w6536 = (w565 & w1962) | (w565 & w5965) | (w1962 & w5965);
assign w6537 = ~w1963 & w5965;
assign w6538 = ~w1710 & w7099;
assign w6539 = ~w2209 & w2205;
assign w6540 = ~w2209 & w1722;
assign w6541 = w2209 & ~w2205;
assign w6542 = w2209 & ~w1722;
assign w6543 = ~w2227 & w2204;
assign w6544 = w2227 & ~w2204;
assign w6545 = (~w726 & w6572) | (~w726 & w7100) | (w6572 & w7100);
assign w6546 = (~w726 & w5672) | (~w726 & w2246) | (w5672 & w2246);
assign w6547 = ~w2246 & w5673;
assign w6548 = ~w2402 & ~w2436;
assign w6549 = w2484 & w5676;
assign w6550 = ~w2546 & ~w1991;
assign w6551 = w2710 & w7793;
assign w6552 = w2710 & w7794;
assign w6553 = w2774 & w7793;
assign w6554 = w2774 & w7794;
assign w6555 = w1710 | w7376;
assign w6556 = (w1715 & w7101) | (w1715 & w7102) | (w7101 & w7102);
assign w6557 = w5687 & w3112;
assign w6558 = (w2852 & w7105) | (w2852 & w7106) | (w7105 & w7106);
assign w6559 = w4033 & w4156;
assign w6560 = w4495 & ~w5036;
assign w6561 = w5107 & w7795;
assign w6562 = (~w6755 & w7377) | (~w6755 & w7378) | (w7377 & w7378);
assign w6563 = (~w6755 & w7379) | (~w6755 & w7380) | (w7379 & w7380);
assign w6564 = (~w6755 & w7381) | (~w6755 & w7382) | (w7381 & w7382);
assign w6565 = (~w6755 & w7383) | (~w6755 & w7384) | (w7383 & w7384);
assign w6566 = (~w6755 & w7385) | (~w6755 & w7386) | (w7385 & w7386);
assign w6567 = (w5284 & w6866) | (w5284 & w7107) | (w6866 & w7107);
assign w6568 = w5232 & w5339;
assign w6569 = (w5828 & w5284) | (w5828 & w7108) | (w5284 & w7108);
assign w6570 = ~w5392 & w5417;
assign w6571 = w1820 & w1963;
assign w6572 = w2393 & ~w726;
assign w6573 = ~w2393 & w726;
assign w6574 = w1959 & ~w726;
assign w6575 = w2393 & w726;
assign w6576 = ~w1959 & w726;
assign w6577 = w1820 & w2436;
assign w6578 = ~w726 & ~w2436;
assign w6579 = w726 & w2436;
assign w6580 = w726 & w5677;
assign w6581 = ~w2393 & ~w726;
assign w6582 = ~w7224 & ~w2903;
assign w6583 = w1820 & w3009;
assign w6584 = w1657 & w7796;
assign w6585 = w1657 & w7797;
assign w6586 = w1502 & w5504;
assign w6587 = w1839 & w2228;
assign w6588 = ~w2045 | w5567;
assign w6589 = (~w2045 & w5567) | (~w2045 & ~w2482) | (w5567 & ~w2482);
assign w6590 = w2482 & w5570;
assign w6591 = w3503 & ~w3722;
assign w6592 = w3595 & ~w3833;
assign w6593 = w5241 & ~w5296;
assign w6594 = w3538 & w3715;
assign w6595 = ~w3854 & ~w3853;
assign w6596 = ~a_8 & a_22;
assign w6597 = ~a_8 & ~w5876;
assign w6598 = a_9 & a_22;
assign w6599 = a_9 & w7798;
assign w6600 = ~w455 & w854;
assign w6601 = ~w455 & w871;
assign w6602 = w871 & ~w1398;
assign w6603 = w428 & w735;
assign w6604 = w735 & ~w1724;
assign w6605 = ~w2395 & w726;
assign w6606 = w2227 & w2204;
assign w6607 = (w2398 & w2410) | (w2398 & w7109) | (w2410 & w7109);
assign w6608 = ~w2410 & w7110;
assign w6609 = (~w726 & w2410) | (~w726 & w7111) | (w2410 & w7111);
assign w6610 = w1959 & ~w565;
assign w6611 = ~w2792 & ~w2229;
assign w6612 = ~w2792 & w5714;
assign w6613 = ~w2812 & w2893;
assign w6614 = ~w2928 & ~w2926;
assign w6615 = w2929 & w2882;
assign w6616 = w2788 & w6904;
assign w6617 = (~w871 & ~w2788) | (~w871 & w6905) | (~w2788 & w6905);
assign w6618 = (w871 & w2410) | (w871 & w7387) | (w2410 & w7387);
assign w6619 = ~w2410 & w7112;
assign w6620 = ~w2484 & w726;
assign w6621 = ~w2482 & w2993;
assign w6622 = w2482 & ~w2993;
assign w6623 = w6555 | w5614;
assign w6624 = (w6555 & w5614) | (w6555 & ~w3024) | (w5614 & ~w3024);
assign w6625 = ~w2812 & w2903;
assign w6626 = ~w2896 & w5620;
assign w6627 = (w2900 & w7113) | (w2900 & w7114) | (w7113 & w7114);
assign w6628 = (~w3161 & w5621) | (~w3161 & w2896) | (w5621 & w2896);
assign w6629 = (~w2878 & ~w6100) | (~w2878 & w7842) | (~w6100 & w7842);
assign w6630 = (~w2878 & ~w6100) | (~w2878 & w7389) | (~w6100 & w7389);
assign w6631 = ~w2812 & w3169;
assign w6632 = w2878 & ~w3216;
assign w6633 = (w2878 & ~w3216) | (w2878 & w7115) | (~w3216 & w7115);
assign w6634 = ~w2812 & w3148;
assign w6635 = w3225 & w7117;
assign w6636 = w2878 & w6103;
assign w6637 = w3243 & w7800;
assign w6638 = w3243 & w7801;
assign w6639 = ~w3250 & w7119;
assign w6640 = ~w3250 & w7391;
assign w6641 = (w2878 & w3311) | (w2878 & w7392) | (w3311 & w7392);
assign w6642 = w2878 & ~w6129;
assign w6643 = w3317 & ~w3309;
assign w6644 = (~w2878 & ~w3323) | (~w2878 & w7393) | (~w3323 & w7393);
assign w6645 = (~w2878 & w6136) | (~w2878 & w2389) | (w6136 & w2389);
assign w6646 = ~w2389 & w6137;
assign w6647 = ~w3358 & w7120;
assign w6648 = w3363 & w7121;
assign w6649 = ~w2812 & w2891;
assign w6650 = w2929 & w2394;
assign w6651 = (~w726 & ~w2788) | (~w726 & w7111) | (~w2788 & w7111);
assign w6652 = w2788 & w7110;
assign w6653 = ~w2896 & w6162;
assign w6654 = (~w3471 & w6163) | (~w3471 & w2896) | (w6163 & w2896);
assign w6655 = (~w2878 & ~w3484) | (~w2878 & w7122) | (~w3484 & w7122);
assign w6656 = (~w2878 & ~w3484) | (~w2878 & w7394) | (~w3484 & w7394);
assign w6657 = ~w2812 & w2411;
assign w6658 = (w3552 & w6176) | (w3552 & w2896) | (w6176 & w2896);
assign w6659 = w3571 & w7123;
assign w6660 = w3571 & w7395;
assign w6661 = ~w3644 & ~w3672;
assign w6662 = w3644 & w3672;
assign w6663 = w3674 & ~w3673;
assign w6664 = ~w3164 & w6904;
assign w6665 = (~w871 & w3164) | (~w871 & w6905) | (w3164 & w6905);
assign w6666 = ~w2812 & w2402;
assign w6667 = w2799 & w1963;
assign w6668 = ~w3863 & ~w3862;
assign w6669 = ~w2812 & w2405;
assign w6670 = (w3472 & w7126) | (w3472 & w7127) | (w7126 & w7127);
assign w6671 = ~w2878 & w7802;
assign w6672 = (~w3472 & w7128) | (~w3472 & w7129) | (w7128 & w7129);
assign w6673 = w2788 & w7398;
assign w6674 = ~w2812 & w1968;
assign w6675 = w4055 & w7130;
assign w6676 = ~w608 & w0;
assign w6677 = (w2878 & w3936) | (w2878 & w7131) | (w3936 & w7131);
assign w6678 = (w3936 & w6976) | (w3936 & w7611) | (w6976 & w7611);
assign w6679 = ~w2812 & w1976;
assign w6680 = ~w2410 & w7132;
assign w6681 = ~w2581 & w4159;
assign w6682 = (w1994 & w2410) | (w1994 & w7133) | (w2410 & w7133);
assign w6683 = w2581 & w4161;
assign w6684 = ~w3164 & w7110;
assign w6685 = (~w726 & w3164) | (~w726 & w7111) | (w3164 & w7111);
assign w6686 = (w6269 & w7399) | (w6269 & w7400) | (w7399 & w7400);
assign w6687 = (~w3555 & w7134) | (~w3555 & w7135) | (w7134 & w7135);
assign w6688 = (~w4207 & w7134) | (~w4207 & w7136) | (w7134 & w7136);
assign w6689 = (w3555 & w7137) | (w3555 & w7138) | (w7137 & w7138);
assign w6690 = (w4207 & w7137) | (w4207 & w7139) | (w7137 & w7139);
assign w6691 = w4145 & ~w4224;
assign w6692 = ~w2799 & w1994;
assign w6693 = ~w2928 & w4269;
assign w6694 = w5765 & w4279;
assign w6695 = (w4279 & w5765) | (w4279 & w4270) | (w5765 & w4270);
assign w6696 = ~w4270 & w5766;
assign w6697 = ~w2812 & w1974;
assign w6698 = (w3472 & w7140) | (w3472 & w7141) | (w7140 & w7141);
assign w6699 = w4318 & ~w6294;
assign w6700 = ~w4130 & w3829;
assign w6701 = ~w4376 & ~w4375;
assign w6702 = ~w2885 & w4385;
assign w6703 = w5770 & ~w4277;
assign w6704 = (~w4277 & w5770) | (~w4277 & w4270) | (w5770 & w4270);
assign w6705 = ~w4270 & w5771;
assign w6706 = ~w4270 & w6310;
assign w6707 = ~w2812 & w1987;
assign w6708 = w4379 & w4466;
assign w6709 = w4472 & ~w4490;
assign w6710 = (~w3555 & w7143) | (~w3555 & w7144) | (w7143 & w7144);
assign w6711 = (~w4207 & w7143) | (~w4207 & w7145) | (w7143 & w7145);
assign w6712 = ~w2812 & w1991;
assign w6713 = ~w3164 & w6849;
assign w6714 = (w565 & w3164) | (w565 & w6850) | (w3164 & w6850);
assign w6715 = (~w4572 & w4563) | (~w4572 & w7403) | (w4563 & w7403);
assign w6716 = (~w726 & w4608) | (~w726 & w7146) | (w4608 & w7146);
assign w6717 = ~w726 & ~w6341;
assign w6718 = w4564 & w4614;
assign w6719 = ~w4563 & w7404;
assign w6720 = ~w4564 & ~w4614;
assign w6721 = ~w2812 & w2546;
assign w6722 = w2812 & ~w1022;
assign w6723 = ~w4749 & w7147;
assign w6724 = ~w726 & w6378;
assign w6725 = ~w4473 & w4805;
assign w6726 = w5653 & ~w4762;
assign w6727 = (~w3555 & w7148) | (~w3555 & w7149) | (w7148 & w7149);
assign w6728 = (~w4207 & w7148) | (~w4207 & w7150) | (w7148 & w7150);
assign w6729 = ~w4824 & w4820;
assign w6730 = w2860 & w7803;
assign w6731 = (~w4516 & w7152) | (~w4516 & w7153) | (w7152 & w7153);
assign w6732 = (w4516 & w7154) | (w4516 & w7155) | (w7154 & w7155);
assign w6733 = ~w4803 & w4866;
assign w6734 = ~w2812 & ~w1022;
assign w6735 = ~w4899 & w4900;
assign w6736 = (~w1022 & ~w4904) | (~w1022 & w7156) | (~w4904 & w7156);
assign w6737 = (~w1022 & ~w4904) | (~w1022 & w7653) | (~w4904 & w7653);
assign w6738 = (~w565 & w4913) | (~w565 & w7157) | (w4913 & w7157);
assign w6739 = ~w565 & ~w6409;
assign w6740 = w5794 & w7804;
assign w6741 = (w4516 & w7158) | (w4516 & w7159) | (w7158 & w7159);
assign w6742 = (w4516 & w7160) | (w4516 & w7161) | (w7160 & w7161);
assign w6743 = (w4516 & w7162) | (w4516 & w7163) | (w7162 & w7163);
assign w6744 = ~w4900 & ~w4893;
assign w6745 = ~w4893 & w7881;
assign w6746 = (w565 & w4982) | (w565 & w7164) | (w4982 & w7164);
assign w6747 = w565 & ~w6425;
assign w6748 = (w4516 & w7165) | (w4516 & w7166) | (w7165 & w7166);
assign w6749 = (w5837 & w4931) | (w5837 & w7167) | (w4931 & w7167);
assign w6750 = (w5837 & w5838) | (w5837 & w7804) | (w5838 & w7804);
assign w6751 = (w4516 & w7168) | (w4516 & w7169) | (w7168 & w7169);
assign w6752 = (w5841 & w4931) | (w5841 & w7170) | (w4931 & w7170);
assign w6753 = (w5841 & w5842) | (w5841 & w7804) | (w5842 & w7804);
assign w6754 = w4963 & w5011;
assign w6755 = ~w5033 & ~w5032;
assign w6756 = (~w6755 & w7405) | (~w6755 & w7406) | (w7405 & w7406);
assign w6757 = (~w3555 & w7171) | (~w3555 & w7172) | (w7171 & w7172);
assign w6758 = (~w4207 & w7171) | (~w4207 & w7173) | (w7171 & w7173);
assign w6759 = w4970 & w7175;
assign w6760 = (w3568 & w7176) | (w3568 & w7177) | (w7176 & w7177);
assign w6761 = w4973 & w7805;
assign w6762 = ~w5021 & ~w5077;
assign w6763 = w5021 & w5077;
assign w6764 = w6444 | w6445;
assign w6765 = (w4973 & w7482) | (w4973 & w7806) | (w7482 & w7806);
assign w6766 = (w3472 & w7178) | (w3472 & w7179) | (w7178 & w7179);
assign w6767 = ~w1022 & w7807;
assign w6768 = (~w3472 & w7180) | (~w3472 & w7181) | (w7180 & w7181);
assign w6769 = (~w5035 & w7407) | (~w5035 & w7408) | (w7407 & w7408);
assign w6770 = (w4674 & w6769) | (w4674 & w7182) | (w6769 & w7182);
assign w6771 = (~w5035 & w7409) | (~w5035 & w7410) | (w7409 & w7410);
assign w6772 = (w4674 & w6771) | (w4674 & w7183) | (w6771 & w7183);
assign w6773 = w5021 & w5134;
assign w6774 = w5139 & ~w5030;
assign w6775 = w5139 & ~w4806;
assign w6776 = w5808 | ~w5142;
assign w6777 = (~w5142 & w5808) | (~w5142 & ~w5021) | (w5808 & ~w5021);
assign w6778 = w6453 & ~w5144;
assign w6779 = (~w5144 & w6453) | (~w5144 & w5145) | (w6453 & w5145);
assign w6780 = ~w5145 & w6454;
assign w6781 = (~w1022 & w5158) | (~w1022 & w7184) | (w5158 & w7184);
assign w6782 = ~w1022 & ~w6460;
assign w6783 = (w7566 & w7185) | (w7566 & w7186) | (w7185 & w7186);
assign w6784 = (w4674 & w7411) | (w4674 & w7412) | (w7411 & w7412);
assign w6785 = (w6869 & w7187) | (w6869 & w7188) | (w7187 & w7188);
assign w6786 = (~w4674 & w7413) | (~w4674 & w7414) | (w7413 & w7414);
assign w6787 = (w7525 & w7189) | (w7525 & w7190) | (w7189 & w7190);
assign w6788 = (w4674 & w7272) | (w4674 & w7273) | (w7272 & w7273);
assign w6789 = (w6872 & w7191) | (w6872 & w7192) | (w7191 & w7192);
assign w6790 = (~w4674 & w7415) | (~w4674 & w7416) | (w7415 & w7416);
assign w6791 = ~w5198 & ~w6454;
assign w6792 = ~w5198 & ~w3829;
assign w6793 = (w3555 & w7193) | (w3555 & w7194) | (w7193 & w7194);
assign w6794 = (w4207 & w7193) | (w4207 & w7195) | (w7193 & w7195);
assign w6795 = w5160 & w6469;
assign w6796 = w6470 & w5204;
assign w6797 = (w5204 & w6470) | (w5204 & ~w5160) | (w6470 & ~w5160);
assign w6798 = (~w5035 & w7417) | (~w5035 & w7418) | (w7417 & w7418);
assign w6799 = (w4674 & w6798) | (w4674 & w7196) | (w6798 & w7196);
assign w6800 = (~w5035 & w7419) | (~w5035 & w7420) | (w7419 & w7420);
assign w6801 = (w4674 & w6800) | (w4674 & w7197) | (w6800 & w7197);
assign w6802 = w5246 & ~w5030;
assign w6803 = w5246 & ~w4806;
assign w6804 = ~w5810 & ~w5249;
assign w6805 = w5254 & w5294;
assign w6806 = ~w5310 & ~w5311;
assign w6807 = (~w5310 & ~w5311) | (~w5310 & w7655) | (~w5311 & w7655);
assign w6808 = w5316 & ~w3829;
assign w6809 = w5316 & ~w6487;
assign w6810 = (w5330 & w6495) | (w5330 & w5311) | (w6495 & w5311);
assign w6811 = (w5311 & w7656) | (w5311 & w7657) | (w7656 & w7657);
assign w6812 = w5335 & ~w5030;
assign w6813 = w5335 & ~w4806;
assign w6814 = w5341 & ~w5030;
assign w6815 = w5341 & ~w4806;
assign w6816 = (~w5243 & w7658) | (~w5243 & w7659) | (w7658 & w7659);
assign w6817 = (w5330 & w5297) | (w5330 & w7660) | (w5297 & w7660);
assign w6818 = w5814 & w5375;
assign w6819 = w5392 & ~w3829;
assign w6820 = (w5392 & w5375) | (w5392 & w6819) | (w5375 & w6819);
assign w6821 = ~w5375 & w5396;
assign w6822 = (w5857 & ~w5297) | (w5857 & w7661) | (~w5297 & w7661);
assign w6823 = (w5400 & w5858) | (w5400 & w5297) | (w5858 & w5297);
assign w6824 = (w5297 & w7662) | (w5297 & w7663) | (w7662 & w7663);
assign w6825 = w5409 & ~w5667;
assign w6826 = (w5821 & w5375) | (w5821 & w7199) | (w5375 & w7199);
assign w6827 = (w5375 & w7200) | (w5375 & w7201) | (w7200 & w7201);
assign w6828 = w3033 & ~w3008;
assign w6829 = ~w4282 & w4266;
assign w6830 = ~w4282 & ~w4173;
assign w6831 = w4282 & ~w4266;
assign w6832 = w4282 & w4173;
assign w6833 = (~w4463 & w5690) | (~w4463 & ~w4379) | (w5690 & ~w4379);
assign w6834 = w5260 & ~w5216;
assign w6835 = (~w6755 & w7421) | (~w6755 & w7422) | (w7421 & w7422);
assign w6836 = (w5151 & w7664) | (w5151 & w7665) | (w7664 & w7665);
assign w6837 = (w7063 & w7423) | (w7063 & w7424) | (w7423 & w7424);
assign w6838 = w871 & ~w3009;
assign w6839 = ~w871 & w3009;
assign w6840 = ~w871 & w5684;
assign w6841 = ~w5057 & w5056;
assign w6842 = w2863 & ~w2900;
assign w6843 = ~w1710 & w7203;
assign w6844 = w2807 & w7204;
assign w6845 = w2807 & w7205;
assign w6846 = ~w2863 & ~w3177;
assign w6847 = w2863 & w3177;
assign w6848 = ~w3206 & ~w3487;
assign w6849 = w1962 & w7206;
assign w6850 = (w565 & ~w1962) | (w565 & w5965) | (~w1962 & w5965);
assign w6851 = ~w6968 & w7425;
assign w6852 = (w3784 & w3562) | (w3784 & w7207) | (w3562 & w7207);
assign w6853 = w4274 & w4279;
assign w6854 = ~w4274 & ~w4279;
assign w6855 = w4307 & w4388;
assign w6856 = ~w4307 & ~w4388;
assign w6857 = w4274 & ~w4277;
assign w6858 = ~w4274 & ~w4407;
assign w6859 = ~w4581 & w4450;
assign w6860 = ~w4581 & ~w5650;
assign w6861 = w4929 & w4940;
assign w6862 = w4948 & ~w4949;
assign w6863 = w4948 & w5796;
assign w6864 = ~w5800 & w5138;
assign w6865 = w1957 & w2436;
assign w6866 = ~w5330 & ~w5307;
assign w6867 = ~w5151 & w7495;
assign w6868 = (w5180 & ~w5691) | (w5180 & w5844) | (~w5691 & w5844);
assign w6869 = (w6755 & w7426) | (w6755 & w7427) | (w7426 & w7427);
assign w6870 = ~w5151 & w7497;
assign w6871 = (w5166 & ~w5691) | (w5166 & w5213) | (~w5691 & w5213);
assign w6872 = w5166 & ~w6564;
assign w6873 = ~w5284 & ~w5232;
assign w6874 = ~w5243 & w6873;
assign w6875 = w5284 & w5232;
assign w6876 = (w5284 & w5243) | (w5284 & w6875) | (w5243 & w6875);
assign w6877 = ~w4929 & ~w4940;
assign w6878 = a_9 & ~a_22;
assign w6879 = ~a_22 & a_12;
assign w6880 = (~w854 & ~w819) | (~w854 & w7208) | (~w819 & w7208);
assign w6881 = ~a_22 & ~a_14;
assign w6882 = a_22 & a_14;
assign w6883 = (~w871 & ~w828) | (~w871 & w7209) | (~w828 & w7209);
assign w6884 = w828 & w7210;
assign w6885 = (w391 & ~w526) | (w391 & w7211) | (~w526 & w7211);
assign w6886 = w693 & w2180;
assign w6887 = ~w1959 & w565;
assign w6888 = ~w2405 & ~w2402;
assign w6889 = ~w1022 & ~w5526;
assign w6890 = ~w1710 & w7213;
assign w6891 = ~w1063 & w7214;
assign w6892 = (w1022 & w1063) | (w1022 & w5963) | (w1063 & w5963);
assign w6893 = ~w2647 & ~w2650;
assign w6894 = ~w2402 & w2398;
assign w6895 = w2402 & w726;
assign w6896 = ~w2402 & ~w726;
assign w6897 = ~w1656 & w2711;
assign w6898 = ~w1656 & w2722;
assign w6899 = w2684 & w2734;
assign w6900 = ~w2684 & ~w2734;
assign w6901 = w2734 & w7215;
assign w6902 = ~w6899 & ~w2844;
assign w6903 = ~w2896 & w2903;
assign w6904 = w2903 & w871;
assign w6905 = ~w2903 & ~w871;
assign w6906 = ~w2884 & w871;
assign w6907 = ~w2891 & ~w2893;
assign w6908 = (w1710 & w6905) | (w1710 & w7216) | (w6905 & w7216);
assign w6909 = (~w871 & w1710) | (~w871 & w7217) | (w1710 & w7217);
assign w6910 = w2893 & w871;
assign w6911 = ~w2893 & ~w871;
assign w6912 = ~w2900 & w7218;
assign w6913 = (w3142 & w2900) | (w3142 & w7219) | (w2900 & w7219);
assign w6914 = ~w2900 & w7220;
assign w6915 = (~w3161 & w2900) | (~w3161 & w7221) | (w2900 & w7221);
assign w6916 = ~w3199 & ~w3200;
assign w6917 = (w2878 & w3164) | (w2878 & w7222) | (w3164 & w7222);
assign w6918 = ~w2896 & w3169;
assign w6919 = ~w3222 & ~w3175;
assign w6920 = w3222 & ~w2878;
assign w6921 = (~w3175 & ~w2788) | (~w3175 & w7223) | (~w2788 & w7223);
assign w6922 = w2788 & w7561;
assign w6923 = (~w3175 & w2410) | (~w3175 & w7505) | (w2410 & w7505);
assign w6924 = ~w871 & ~w5683;
assign w6925 = ~w1710 & w7224;
assign w6926 = ~w1710 & w7225;
assign w6927 = ~w2878 & ~w3175;
assign w6928 = ~w1710 & w7226;
assign w6929 = w3316 & ~w3175;
assign w6930 = w3316 & ~w2878;
assign w6931 = ~w2368 & w3175;
assign w6932 = (w2878 & w2410) | (w2878 & w7222) | (w2410 & w7222);
assign w6933 = ~w2896 & w3173;
assign w6934 = ~w3351 & w2878;
assign w6935 = ~w3351 & w6976;
assign w6936 = ~w2896 & w3148;
assign w6937 = ~w2896 & w2893;
assign w6938 = (w2878 & w3474) | (w2878 & w7222) | (w3474 & w7222);
assign w6939 = ~w2900 & w7227;
assign w6940 = (w3169 & ~w423) | (w3169 & w7228) | (~w423 & w7228);
assign w6941 = ~w3474 & w7229;
assign w6942 = ~w2896 & w2891;
assign w6943 = ~w2896 & w2411;
assign w6944 = ~w1022 & ~w1994;
assign w6945 = ~w1972 & w5965;
assign w6946 = (~w565 & w1972) | (~w565 & w7206) | (w1972 & w7206);
assign w6947 = (~w1976 & w6968) | (~w1976 & w7428) | (w6968 & w7428);
assign w6948 = (w3148 & ~w423) | (w3148 & w7230) | (~w423 & w7230);
assign w6949 = ~w3472 & w7232;
assign w6950 = (w3791 & w7233) | (w3791 & w7234) | (w7233 & w7234);
assign w6951 = (w3791 & w7429) | (w3791 & w7430) | (w7429 & w7430);
assign w6952 = w2788 & w7237;
assign w6953 = (~w565 & ~w2788) | (~w565 & w7238) | (~w2788 & w7238);
assign w6954 = ~w2896 & w2402;
assign w6955 = ~w3904 & ~w726;
assign w6956 = ~w3904 & w6578;
assign w6957 = ~w3474 & w7112;
assign w6958 = (w3173 & ~w423) | (w3173 & w7240) | (~w423 & w7240);
assign w6959 = ~w3944 & ~w6236;
assign w6960 = w2878 & w6237;
assign w6961 = ~w3943 & w7241;
assign w6962 = (~w2878 & w3943) | (~w2878 & w7242) | (w3943 & w7242);
assign w6963 = ~w2896 & w2405;
assign w6964 = (w2903 & ~w423) | (w2903 & w7243) | (~w423 & w7243);
assign w6965 = w4073 & ~w2878;
assign w6966 = ~w2896 & w1968;
assign w6967 = ~w4152 & ~w565;
assign w6968 = (~w565 & w1962) | (~w565 & w6610) | (w1962 & w6610);
assign w6969 = w4152 & w565;
assign w6970 = ~w1962 & w6887;
assign w6971 = w1987 & w4164;
assign w6972 = ~w1987 & ~w4164;
assign w6973 = (w2893 & ~w423) | (w2893 & w7245) | (~w423 & w7245);
assign w6974 = (w3472 & w7246) | (w3472 & w7247) | (w7246 & w7247);
assign w6975 = w4208 & ~w6274;
assign w6976 = ~w3175 & w2878;
assign w6977 = w2878 & ~w6975;
assign w6978 = (w2878 & ~w4208) | (w2878 & w7248) | (~w4208 & w7248);
assign w6979 = ~w2878 & w6975;
assign w6980 = w4208 & w7249;
assign w6981 = ~w1987 & w4264;
assign w6982 = ~w2896 & w1976;
assign w6983 = (~w565 & w4288) | (~w565 & w7250) | (w4288 & w7250);
assign w6984 = ~w4288 & w7251;
assign w6985 = w2411 & ~w726;
assign w6986 = ~w2411 & w726;
assign w6987 = ~w4313 & w7252;
assign w6988 = ~w4313 & w7253;
assign w6989 = (w2891 & ~w423) | (w2891 & w7254) | (~w423 & w7254);
assign w6990 = w4313 & w7255;
assign w6991 = ~w4316 & ~w6296;
assign w6992 = (~w3472 & w7256) | (~w3472 & w7257) | (w7256 & w7257);
assign w6993 = (w3472 & w7609) | (w3472 & w7608) | (w7609 & w7608);
assign w6994 = (w2411 & ~w423) | (w2411 & w7432) | (~w423 & w7432);
assign w6995 = (~w726 & w3472) | (~w726 & w7258) | (w3472 & w7258);
assign w6996 = (w3472 & w6578) | (w3472 & w7259) | (w6578 & w7259);
assign w6997 = ~w4274 & ~w4411;
assign w6998 = w1991 & w1022;
assign w6999 = ~w1991 & ~w1022;
assign w7000 = ~w2896 & w1974;
assign w7001 = (w3009 & ~w3779) | (w3009 & w7260) | (~w3779 & w7260);
assign w7002 = ~w2891 & ~w7001;
assign w7003 = (~w2891 & w6274) | (~w2891 & w6322) | (w6274 & w6322);
assign w7004 = w4399 & ~w4520;
assign w7005 = ~w4399 & w4520;
assign w7006 = ~w2896 & w1987;
assign w7007 = (w2402 & ~w423) | (w2402 & w7261) | (~w423 & w7261);
assign w7008 = (w3472 & w7433) | (w3472 & w7434) | (w7433 & w7434);
assign w7009 = (w2405 & ~w423) | (w2405 & w7435) | (~w423 & w7435);
assign w7010 = ~w4609 & ~w6340;
assign w7011 = ~w4609 & w726;
assign w7012 = ~w2896 & w1991;
assign w7013 = w4517 & ~w4686;
assign w7014 = (w1968 & ~w423) | (w1968 & w7436) | (~w423 & w7436);
assign w7015 = w1976 & ~w565;
assign w7016 = ~w1976 & w565;
assign w7017 = ~w2896 & w2546;
assign w7018 = ~w4732 & ~w1994;
assign w7019 = (w4741 & w4624) | (w4741 & w7437) | (w4624 & w7437);
assign w7020 = w6348 & w4635;
assign w7021 = ~w4750 & ~w2436;
assign w7022 = w4750 & w726;
assign w7023 = (w2436 & ~w3779) | (w2436 & w7438) | (~w3779 & w7438);
assign w7024 = ~w2405 & ~w7023;
assign w7025 = (~w2405 & w6274) | (~w2405 & w6384) | (w6274 & w6384);
assign w7026 = ~w4732 & ~w4728;
assign w7027 = w7018 & ~w4728;
assign w7028 = (w1976 & ~w423) | (w1976 & w7439) | (~w423 & w7439);
assign w7029 = (w3472 & w7440) | (w3472 & w7441) | (w7440 & w7441);
assign w7030 = ~w4753 & ~w4757;
assign w7031 = ~w4664 & ~w4847;
assign w7032 = (w1022 & w3474) | (w1022 & w7443) | (w3474 & w7443);
assign w7033 = (w1974 & ~w423) | (w1974 & w7444) | (~w423 & w7444);
assign w7034 = ~w4914 & ~w6408;
assign w7035 = ~w4914 & w565;
assign w7036 = ~w726 & w4890;
assign w7037 = (w1987 & ~w423) | (w1987 & w7445) | (~w423 & w7445);
assign w7038 = (~w1994 & w3472) | (~w1994 & w7446) | (w3472 & w7446);
assign w7039 = ~w4983 & ~w1963;
assign w7040 = ~w4983 & ~w565;
assign w7041 = (w1963 & ~w3779) | (w1963 & w7447) | (~w3779 & w7447);
assign w7042 = ~w1974 & ~w7041;
assign w7043 = (~w1974 & w6274) | (~w1974 & w6432) | (w6274 & w6432);
assign w7044 = (w1022 & w3472) | (w1022 & w7448) | (w3472 & w7448);
assign w7045 = ~w4969 & ~w5048;
assign w7046 = w4969 & w5048;
assign w7047 = ~w7045 & ~w5085;
assign w7048 = (w2546 & ~w423) | (w2546 & w7449) | (~w423 & w7449);
assign w7049 = ~w5094 & ~w6448;
assign w7050 = w1022 & w6450;
assign w7051 = ~w5095 & w7450;
assign w7052 = (~w1022 & w5095) | (~w1022 & w7451) | (w5095 & w7451);
assign w7053 = (~w1022 & ~w423) | (~w1022 & w7666) | (~w423 & w7666);
assign w7054 = ~w5159 & ~w1994;
assign w7055 = ~w5159 & w1022;
assign w7056 = ~w5157 & w6461;
assign w7057 = ~w5157 & w6462;
assign w7058 = (w1994 & ~w3779) | (w1994 & w7452) | (~w3779 & w7452);
assign w7059 = w1022 & ~w3936;
assign w7060 = ~w3936 & w7453;
assign w7061 = w629 & w5221;
assign w7062 = ~w5206 & ~w5208;
assign w7063 = w4883 & w7454;
assign w7064 = (~w1022 & ~w2545) | (~w1022 & w7455) | (~w2545 & w7455);
assign w7065 = (w1022 & w3472) | (w1022 & w7456) | (w3472 & w7456);
assign w7066 = ~w3472 & w7457;
assign w7067 = w5658 & ~w5208;
assign w7068 = (w5658 & w5166) | (w5658 & w7067) | (w5166 & w7067);
assign w7069 = (w5658 & ~w5260) | (w5658 & w7458) | (~w5260 & w7458);
assign w7070 = w4883 & w7459;
assign w7071 = (~w5277 & w5154) | (~w5277 & w7460) | (w5154 & w7460);
assign w7072 = (w5260 & w7461) | (w5260 & w7462) | (w7461 & w7462);
assign w7073 = (~w4883 & w7463) | (~w4883 & w7464) | (w7463 & w7464);
assign w7074 = ~w5277 & ~w5307;
assign w7075 = w5277 & w5307;
assign w7076 = w5330 & w5307;
assign w7077 = ~w5284 & w7465;
assign w7078 = w818 & w854;
assign w7079 = ~w818 & ~w726;
assign w7080 = w818 & w726;
assign w7081 = w818 & w720;
assign w7082 = ~w818 & ~w720;
assign w7083 = w818 & w735;
assign w7084 = ~w818 & ~w735;
assign w7085 = w818 & w574;
assign w7086 = ~w818 & ~w574;
assign w7087 = ~w818 & ~w565;
assign w7088 = w818 & w565;
assign w7089 = w818 & w511;
assign w7090 = ~w818 & ~w511;
assign w7091 = (w847 & ~w819) | (w847 & w7466) | (~w819 & w7466);
assign w7092 = w819 & w7467;
assign w7093 = w818 & ~w880;
assign w7094 = ~w818 & w880;
assign w7095 = ~w1695 & ~w1256;
assign w7096 = ~w1195 & w7808;
assign w7097 = w818 & ~w1022;
assign w7098 = ~w818 & w1022;
assign w7099 = w1982 & w1963;
assign w7100 = ~w2403 | ~w726;
assign w7101 = (w6555 & w871) | (w6555 & ~w5683) | (w871 & ~w5683);
assign w7102 = (w6555 & w871) | (w6555 & w6925) | (w871 & w6925);
assign w7103 = w5687 & w3111;
assign w7104 = w5687 & w6080;
assign w7105 = (~w3161 & w5688) | (~w3161 & ~w3111) | (w5688 & ~w3111);
assign w7106 = (~w3161 & w5688) | (~w3161 & ~w6080) | (w5688 & ~w6080);
assign w7107 = ~w5330 & w7074;
assign w7108 = ~w5277 & w5828;
assign w7109 = ~w2411 & w2398;
assign w7110 = w2411 & w726;
assign w7111 = ~w2411 & ~w726;
assign w7112 = w2903 & ~w871;
assign w7113 = w5688 | ~w3161;
assign w7114 = (w2852 & w7469) | (w2852 & w7470) | (w7469 & w7470);
assign w7115 = w3175 & w2878;
assign w7116 = (w2655 & w6927) | (w2655 & w7471) | (w6927 & w7471);
assign w7117 = ~w3222 & w2878;
assign w7118 = ~w2410 & w7472;
assign w7119 = ~w3251 & w3253;
assign w7120 = ~w3359 & w3365;
assign w7121 = ~w3175 & w3365;
assign w7122 = ~w3474 & w7561;
assign w7123 = (w2878 & w3474) | (w2878 & w7131) | (w3474 & w7131);
assign w7124 = (w2878 & w3472) | (w2878 & w7473) | (w3472 & w7473);
assign w7125 = (w871 & w3474) | (w871 & w7387) | (w3474 & w7387);
assign w7126 = ~w3175 & w6961;
assign w7127 = w6237 & w6976;
assign w7128 = (~w2878 & w3175) | (~w2878 & w6962) | (w3175 & w6962);
assign w7129 = (~w2878 & ~w6237) | (~w2878 & w7620) | (~w6237 & w7620);
assign w7130 = (w3474 & w7667) | (w3474 & w7668) | (w7667 & w7668);
assign w7131 = ~w3148 & w2878;
assign w7132 = w2659 & w1994;
assign w7133 = ~w2659 & w1994;
assign w7134 = (~w3553 & w7669) | (~w3553 & w7670) | (w7669 & w7670);
assign w7135 = (w6275 & w6276) | (w6275 & w4206) | (w6276 & w4206);
assign w7136 = (w6275 & w6276) | (w6275 & ~w3561) | (w6276 & ~w3561);
assign w7137 = (w3553 & w7474) | (w3553 & w7475) | (w7474 & w7475);
assign w7138 = (w7585 & w6277) | (w7585 & ~w4206) | (w6277 & ~w4206);
assign w7139 = (w7585 & w6277) | (w7585 & w3561) | (w6277 & w3561);
assign w7140 = ~w4314 & w6297;
assign w7141 = ~w4314 & w4317;
assign w7142 = ~w3472 & w7476;
assign w7143 = (w6322 & w7717) | (w6322 & w7810) | (w7717 & w7810);
assign w7144 = (w6322 & w6323) | (w6322 & w4206) | (w6323 & w4206);
assign w7145 = (w6322 & w6323) | (w6322 & ~w3561) | (w6323 & ~w3561);
assign w7146 = w4609 & ~w726;
assign w7147 = ~w4750 & ~w726;
assign w7148 = (w6384 & w7586) | (w6384 & w7811) | (w7586 & w7811);
assign w7149 = (w6384 & w6385) | (w6384 & w4206) | (w6385 & w4206);
assign w7150 = (w6384 & w6385) | (w6384 & ~w3561) | (w6385 & ~w3561);
assign w7151 = (~w1994 & ~w2860) | (~w1994 & w7477) | (~w2860 & w7477);
assign w7152 = w4862 & w4809;
assign w7153 = (w4862 & w4810) | (w4862 & w7152) | (w4810 & w7152);
assign w7154 = ~w4862 & ~w4809;
assign w7155 = ~w4810 & w7154;
assign w7156 = ~w3474 & w7212;
assign w7157 = w4914 & ~w565;
assign w7158 = (w4942 & w5795) | (w4942 & w4883) | (w5795 & w4883);
assign w7159 = (w4942 & w5795) | (w4942 & w5656) | (w5795 & w5656);
assign w7160 = (~w4929 & w5834) | (~w4929 & w4883) | (w5834 & w4883);
assign w7161 = (~w4929 & w5834) | (~w4929 & w5656) | (w5834 & w5656);
assign w7162 = (~w4940 & w5859) | (~w4940 & w4883) | (w5859 & w4883);
assign w7163 = (~w4940 & w5859) | (~w4940 & w5656) | (w5859 & w5656);
assign w7164 = w4983 & w565;
assign w7165 = (w5835 & w5836) | (w5835 & w4883) | (w5836 & w4883);
assign w7166 = (w5835 & w5836) | (w5835 & w5656) | (w5836 & w5656);
assign w7167 = w5837 & w5003;
assign w7168 = (w5839 & w5840) | (w5839 & w4883) | (w5840 & w4883);
assign w7169 = (w5839 & w5840) | (w5839 & w5656) | (w5840 & w5656);
assign w7170 = w5841 & w5008;
assign w7171 = (w6432 & w7587) | (w6432 & w7812) | (w7587 & w7812);
assign w7172 = (w6432 & w6433) | (w6432 & w4206) | (w6433 & w4206);
assign w7173 = (w6432 & w6433) | (w6432 & ~w3561) | (w6433 & ~w3561);
assign w7174 = ~w3472 & w7478;
assign w7175 = w7045 & ~w5048;
assign w7176 = (~w4973 & w7479) | (~w4973 & w7480) | (w7479 & w7480);
assign w7177 = (~w4973 & w7479) | (~w4973 & w7481) | (w7479 & w7481);
assign w7178 = ~w1994 & w7051;
assign w7179 = w6450 & w7477;
assign w7180 = (~w1022 & w1994) | (~w1022 & w7052) | (w1994 & w7052);
assign w7181 = (~w1022 & ~w6450) | (~w1022 & w5775) | (~w6450 & w5775);
assign w7182 = (~w5035 & w7671) | (~w5035 & w7672) | (w7671 & w7672);
assign w7183 = (~w5035 & w7483) | (~w5035 & w7484) | (w7483 & w7484);
assign w7184 = w5159 & ~w1022;
assign w7185 = ~w5151 & w7813;
assign w7186 = (w5843 & ~w4883) | (w5843 & w7485) | (~w4883 & w7485);
assign w7187 = w5844 | w6868;
assign w7188 = (w5844 & w4883) | (w5844 & w7486) | (w4883 & w7486);
assign w7189 = ~w5151 & w7814;
assign w7190 = (w5845 & ~w4883) | (w5845 & w7487) | (~w4883 & w7487);
assign w7191 = w5213 | w6871;
assign w7192 = (w5213 & w4883) | (w5213 & w7488) | (w4883 & w7488);
assign w7193 = (w3553 & w7489) | (w3553 & w7490) | (w7489 & w7490);
assign w7194 = (w1994 & w6465) | (w1994 & ~w4206) | (w6465 & ~w4206);
assign w7195 = (w1994 & w6465) | (w1994 & w3561) | (w6465 & w3561);
assign w7196 = (~w5035 & w7491) | (~w5035 & w7492) | (w7491 & w7492);
assign w7197 = (~w5035 & w7673) | (~w5035 & w7674) | (w7673 & w7674);
assign w7198 = w5330 & ~w6491;
assign w7199 = (w5388 & w7493) | (w5388 & w7494) | (w7493 & w7494);
assign w7200 = w5821 | w5415;
assign w7201 = (w5415 & w5821) | (w5415 & ~w3829) | (w5821 & ~w3829);
assign w7202 = (w5307 & w5267) | (w5307 & w7075) | (w5267 & w7075);
assign w7203 = w2392 & w3009;
assign w7204 = w2895 & ~w3142;
assign w7205 = w2895 & ~w3111;
assign w7206 = ~w1959 & ~w565;
assign w7207 = ~w3555 & w3784;
assign w7208 = ~w818 & ~w854;
assign w7209 = (~w871 & ~w819) | (~w871 & w7498) | (~w819 & w7498);
assign w7210 = w819 & w7499;
assign w7211 = ~w524 & w391;
assign w7212 = ~w1022 & w1987;
assign w7213 = w1991 & ~w1022;
assign w7214 = w565 & ~w1022;
assign w7215 = w2684 & ~w2731;
assign w7216 = ~w871 & w6582;
assign w7217 = ~w2881 & ~w871;
assign w7218 = (~w3142 & ~w2852) | (~w3142 & w7500) | (~w2852 & w7500);
assign w7219 = w2852 & w7501;
assign w7220 = w3161 & w3112;
assign w7221 = (w2852 & w7503) | (w2852 & w7504) | (w7503 & w7504);
assign w7222 = ~w3169 & w2878;
assign w7223 = ~w3169 & ~w3175;
assign w7224 = w2881 & ~w871;
assign w7225 = w2881 & w7882;
assign w7226 = w2881 & w2878;
assign w7227 = w3559 & w3112;
assign w7228 = ~w418 & w3169;
assign w7229 = w3148 & ~w2878;
assign w7230 = ~w418 & w3148;
assign w7231 = (w3550 & w7505) | (w3550 & w7506) | (w7505 & w7506);
assign w7232 = ~w2878 & w7815;
assign w7233 = (w2878 & ~w3804) | (w2878 & w7507) | (~w3804 & w7507);
assign w7234 = (~w3805 & w3472) | (~w3805 & w7508) | (w3472 & w7508);
assign w7235 = w3804 & w7509;
assign w7236 = ~w3472 & w7510;
assign w7237 = w1968 & w565;
assign w7238 = ~w1968 & ~w565;
assign w7239 = ~w2903 & ~w3009;
assign w7240 = ~w418 & w3173;
assign w7241 = ~w3944 & w2878;
assign w7242 = w3944 & ~w2878;
assign w7243 = ~w418 & w2903;
assign w7244 = ~a_0 & ~w3148;
assign w7245 = ~w418 & w2893;
assign w7246 = w871 & ~w4200;
assign w7247 = w871 & w6272;
assign w7248 = w3779 & w7511;
assign w7249 = (~w2878 & ~w3779) | (~w2878 & w7512) | (~w3779 & w7512);
assign w7250 = w1963 & ~w565;
assign w7251 = ~w1963 & w565;
assign w7252 = w3779 & w7513;
assign w7253 = w3009 & w6212;
assign w7254 = ~w418 & w2891;
assign w7255 = w3009 & ~w6212;
assign w7256 = ~w871 & w6990;
assign w7257 = w4313 & w7514;
assign w7258 = (w3550 & w7111) | (w3550 & w7515) | (w7111 & w7515);
assign w7259 = (w3550 & w7676) | (w3550 & w7677) | (w7676 & w7677);
assign w7260 = ~w608 & w3009;
assign w7261 = ~w418 & w2402;
assign w7262 = ~w4588 & ~w4587;
assign w7263 = w5776 & ~w4581;
assign w7264 = (~w4581 & w5776) | (~w4581 & w4495) | (w5776 & w4495);
assign w7265 = ~w4676 & ~w4675;
assign w7266 = w4677 & w4686;
assign w7267 = ~w4690 & ~w4689;
assign w7268 = ~w4701 & w4796;
assign w7269 = w4701 & ~w4796;
assign w7270 = (~w4674 & w7518) | (~w4674 & w7519) | (w7518 & w7519);
assign w7271 = (w4674 & w7522) | (w4674 & w7523) | (w7522 & w7523);
assign w7272 = (~w5035 & w7189) | (~w5035 & w7524) | (w7189 & w7524);
assign w7273 = (~w5035 & w7525) | (~w5035 & w7526) | (w7525 & w7526);
assign w7274 = ~a_10 & a_22;
assign w7275 = ~a_10 & ~w5865;
assign w7276 = ~a_11 & a_22;
assign w7277 = ~a_11 & w7816;
assign w7278 = ~w2666 & w6025;
assign w7279 = (w726 & w6026) | (w726 & w2666) | (w6026 & w2666);
assign w7280 = ~w2666 & w6027;
assign w7281 = ~w2677 & w7527;
assign w7282 = (~w2691 & w2734) | (~w2691 & w7817) | (w2734 & w7817);
assign w7283 = (w2677 & w7678) | (w2677 & w7679) | (w7678 & w7679);
assign w7284 = ~w2677 & w7528;
assign w7285 = (~w2691 & w6044) | (~w2691 & w7818) | (w6044 & w7818);
assign w7286 = w3180 & w2902;
assign w7287 = (w3480 & w6165) | (w3480 & ~w5739) | (w6165 & ~w5739);
assign w7288 = (w3480 & w6165) | (w3480 & w6095) | (w6165 & w6095);
assign w7289 = w3566 & ~w5739;
assign w7290 = w3566 & w6095;
assign w7291 = (w565 & ~w2410) | (w565 & w7529) | (~w2410 & w7529);
assign w7292 = (w565 & w6207) | (w565 & w3740) | (w6207 & w3740);
assign w7293 = ~w3740 & w6208;
assign w7294 = ~w3740 & w6209;
assign w7295 = (~w2878 & ~w3791) | (~w2878 & w7819) | (~w3791 & w7819);
assign w7296 = (~w2878 & ~w3791) | (~w2878 & w7820) | (~w3791 & w7820);
assign w7297 = (w4067 & ~w3786) | (w4067 & w7531) | (~w3786 & w7531);
assign w7298 = (w4069 & w3786) | (w4069 & w7532) | (w3786 & w7532);
assign w7299 = (~w871 & w4201) | (~w871 & w7821) | (w4201 & w7821);
assign w7300 = (~w871 & w4201) | (~w871 & w7822) | (w4201 & w7822);
assign w7301 = (w6689 & w6690) | (w6689 & ~w5739) | (w6690 & ~w5739);
assign w7302 = (w6689 & w6690) | (w6689 & w6095) | (w6690 & w6095);
assign w7303 = ~w4205 & w7823;
assign w7304 = ~w4205 & w7824;
assign w7305 = ~w4287 & ~w4288;
assign w7306 = (w6311 & ~w5770) | (w6311 & w7533) | (~w5770 & w7533);
assign w7307 = ~w4404 & ~w6704;
assign w7308 = w6324 & w7883;
assign w7309 = w6324 & w7826;
assign w7310 = (w726 & w4569) | (w726 & w7827) | (w4569 & w7827);
assign w7311 = (w726 & w4569) | (w726 & w7828) | (w4569 & w7828);
assign w7312 = ~w4623 & ~w4624;
assign w7313 = w3829 & ~w4799;
assign w7314 = ~w3829 & w4799;
assign w7315 = w6386 & w7829;
assign w7316 = w6386 & w7830;
assign w7317 = (w565 & w4836) | (w565 & w7884) | (w4836 & w7884);
assign w7318 = (w565 & w4836) | (w565 & w7885) | (w4836 & w7885);
assign w7319 = ~w726 & w3171;
assign w7320 = ~w4901 & ~w4967;
assign w7321 = w6434 & w7831;
assign w7322 = w6434 & w7832;
assign w7323 = (~w1022 & ~w5041) | (~w1022 & w7886) | (~w5041 & w7886);
assign w7324 = (~w1022 & ~w5041) | (~w1022 & w7887) | (~w5041 & w7887);
assign w7325 = ~w5051 & ~w5046;
assign w7326 = (w6468 & w6467) | (w6468 & w7833) | (w6467 & w7833);
assign w7327 = (w6468 & w6467) | (w6468 & w7834) | (w6467 & w7834);
assign w7328 = ~w5253 & ~w3829;
assign w7329 = ~w5253 & ~w5848;
assign w7330 = w6489 & w6488;
assign w7331 = (w4674 & w7330) | (w4674 & w7534) | (w7330 & w7534);
assign w7332 = (w7535 & w5243) | (w7535 & w7680) | (w5243 & w7680);
assign w7333 = ~w5297 & w7681;
assign w7334 = (~w5243 & w7682) | (~w5243 & w7683) | (w7682 & w7683);
assign w7335 = (w5362 & w5297) | (w5362 & w7684) | (w5297 & w7684);
assign w7336 = (~w5243 & w7685) | (~w5243 & w7686) | (w7685 & w7686);
assign w7337 = (w5297 & w7537) | (w5297 & w7739) | (w7537 & w7739);
assign w7338 = (~w5137 & w7687) | (~w5137 & w7688) | (w7687 & w7688);
assign w7339 = (w5403 & w7539) | (w5403 & w7740) | (w7539 & w7740);
assign w7340 = w6072 & ~w2484;
assign w7341 = w6837 | w6836;
assign w7342 = (w6836 & w6837) | (w6836 & w7835) | (w6837 & w7835);
assign w7343 = ~w5071 & w4883;
assign w7344 = w5071 & ~w4883;
assign w7345 = (~w5137 & w7699) | (~w5137 & w7700) | (w7699 & w7700);
assign w7346 = ~w5071 & ~w4930;
assign w7347 = (w5284 & w7540) | (w5284 & w7541) | (w7540 & w7541);
assign w7348 = (w5400 & ~w5828) | (w5400 & w7836) | (~w5828 & w7836);
assign w7349 = w2607 & ~w2606;
assign w7350 = (w2788 & w7620) | (w2788 & w7542) | (w7620 & w7542);
assign w7351 = (~w2852 & w7543) | (~w2852 & w7544) | (w7543 & w7544);
assign w7352 = (w2852 & w7545) | (w2852 & w7546) | (w7545 & w7546);
assign w7353 = (w3474 & w6976) | (w3474 & w7547) | (w6976 & w7547);
assign w7354 = (w2852 & w7548) | (w2852 & w7549) | (w7548 & w7549);
assign w7355 = ~w2878 & w7837;
assign w7356 = (~w3472 & w7620) | (~w3472 & w7550) | (w7620 & w7550);
assign w7357 = (~w3791 & w7235) | (~w3791 & w7838) | (w7235 & w7838);
assign w7358 = (~w3791 & w7235) | (~w3791 & w7839) | (w7235 & w7839);
assign w7359 = ~w871 & w7888;
assign w7360 = (~w871 & ~w2881) | (~w871 & w7551) | (~w2881 & w7551);
assign w7361 = (~w2885 & w3474) | (~w2885 & w7552) | (w3474 & w7552);
assign w7362 = ~w4152 & w6968;
assign w7363 = (w565 & w6887) | (w565 & w7553) | (w6887 & w7553);
assign w7364 = (w565 & w6970) | (w565 & w4152) | (w6970 & w4152);
assign w7365 = (w3164 & w6578) | (w3164 & w7554) | (w6578 & w7554);
assign w7366 = (w3472 & w7555) | (w3472 & w7556) | (w7555 & w7556);
assign w7367 = w6992 & w3782;
assign w7368 = (w6992 & ~w3786) | (w6992 & w7367) | (~w3786 & w7367);
assign w7369 = (w871 & w6993) | (w871 & ~w3782) | (w6993 & ~w3782);
assign w7370 = (w3786 & w7557) | (w3786 & w7369) | (w7557 & w7369);
assign w7371 = (w3472 & w7689) | (w3472 & w7690) | (w7689 & w7690);
assign w7372 = ~w5093 & w5086;
assign w7373 = (w5260 & w7691) | (w5260 & w7692) | (w7691 & w7692);
assign w7374 = w5278 & w6835;
assign w7375 = (w4496 & w7558) | (w4496 & w7559) | (w7558 & w7559);
assign w7376 = w847 | w871;
assign w7377 = w5107 & w7889;
assign w7378 = w5107 & w7841;
assign w7379 = (~w5111 & w5826) | (~w5111 & w5032) | (w5826 & w5032);
assign w7380 = (~w5111 & w5826) | (~w5111 & w4930) | (w5826 & w4930);
assign w7381 = (~w5151 & w5691) | (~w5151 & w5032) | (w5691 & w5032);
assign w7382 = (~w5151 & w5691) | (~w5151 & w4930) | (w5691 & w4930);
assign w7383 = (w5214 & w5827) | (w5214 & w5032) | (w5827 & w5032);
assign w7384 = (w5214 & w5827) | (w5214 & w4930) | (w5827 & w4930);
assign w7385 = (~w5218 & w5692) | (~w5218 & w5032) | (w5692 & w5032);
assign w7386 = (~w5218 & w5692) | (~w5218 & w4930) | (w5692 & w4930);
assign w7387 = ~w2903 & w871;
assign w7388 = (w3164 & w6976) | (w3164 & w7560) | (w6976 & w7560);
assign w7389 = (w3175 & ~w2878) | (w3175 & w7842) | (~w2878 & w7842);
assign w7390 = w2878 & ~w6923;
assign w7391 = w6923 & w3253;
assign w7392 = ~w3316 & w2878;
assign w7393 = ~w2410 & w7561;
assign w7394 = ~w2878 & w7843;
assign w7395 = (w3474 & w7611) | (w3474 & w6976) | (w7611 & w6976);
assign w7396 = (w3472 & w6976) | (w3472 & w7562) | (w6976 & w7562);
assign w7397 = (w3474 & w6838) | (w3474 & w7693) | (w6838 & w7693);
assign w7398 = w2772 & w1963;
assign w7399 = (~w726 & w2393) | (~w726 & w7563) | (w2393 & w7563);
assign w7400 = (~w2396 & w3164) | (~w2396 & w7564) | (w3164 & w7564);
assign w7401 = (~w3472 & w6579) | (~w3472 & w7694) | (w6579 & w7694);
assign w7402 = w726 & w7844;
assign w7403 = w4425 & ~w4572;
assign w7404 = ~w4425 & w4572;
assign w7405 = ~w5031 & w5032;
assign w7406 = ~w5031 & w4930;
assign w7407 = w5107 & w7846;
assign w7408 = w5108 & w6562;
assign w7409 = w5826 & ~w5111;
assign w7410 = ~w5111 & w6563;
assign w7411 = (~w5035 & w7185) | (~w5035 & w7565) | (w7185 & w7565);
assign w7412 = (~w5035 & w7566) | (~w5035 & w7567) | (w7566 & w7567);
assign w7413 = (w5035 & w7187) | (w5035 & w7695) | (w7187 & w7695);
assign w7414 = (w5035 & w7568) | (w5035 & w7569) | (w7568 & w7569);
assign w7415 = w5846 | w5213;
assign w7416 = (w5213 & w5846) | (w5213 & w5034) | (w5846 & w5034);
assign w7417 = w5827 & w5214;
assign w7418 = w5214 & w6565;
assign w7419 = w5692 & ~w5218;
assign w7420 = ~w5218 & w6566;
assign w7421 = (w5260 & w6834) | (w5260 & w5032) | (w6834 & w5032);
assign w7422 = (w5260 & w6834) | (w5260 & w4930) | (w6834 & w4930);
assign w7423 = (~w5260 & w7696) | (~w5260 & w7697) | (w7696 & w7697);
assign w7424 = (w5307 & w7202) | (w5307 & ~w6835) | (w7202 & ~w6835);
assign w7425 = ~w2563 & ~w1968;
assign w7426 = (w5180 & w5151) | (w5180 & w7847) | (w5151 & w7847);
assign w7427 = (w5180 & w5151) | (w5180 & w7848) | (w5151 & w7848);
assign w7428 = w2563 & ~w1976;
assign w7429 = w7233 & ~w3805;
assign w7430 = (w3472 & w7570) | (w3472 & w7571) | (w7570 & w7571);
assign w7431 = (~w3472 & w7572) | (~w3472 & w7573) | (w7572 & w7573);
assign w7432 = ~w418 & w2411;
assign w7433 = ~w726 & ~w4568;
assign w7434 = ~w726 & w6338;
assign w7435 = ~w418 & w2405;
assign w7436 = ~w418 & w1968;
assign w7437 = w1994 & w4741;
assign w7438 = ~w608 & w2436;
assign w7439 = ~w418 & w1976;
assign w7440 = ~w565 & ~w4835;
assign w7441 = ~w565 & w6395;
assign w7442 = ~w1987 & ~w1994;
assign w7443 = ~w1987 & w1022;
assign w7444 = ~w418 & w1974;
assign w7445 = ~w418 & w1987;
assign w7446 = (w3550 & w7442) | (w3550 & w7574) | (w7442 & w7574);
assign w7447 = ~w608 & w1963;
assign w7448 = (w3550 & w7703) | (w3550 & w7577) | (w7703 & w7577);
assign w7449 = ~w418 & w2546;
assign w7450 = ~w5094 & w1022;
assign w7451 = w5094 & ~w1022;
assign w7452 = ~w608 & w1994;
assign w7453 = w2545 & w7578;
assign w7454 = ~w4927 & w7579;
assign w7455 = w1990 & ~w1022;
assign w7456 = ~w6479 & w1022;
assign w7457 = w6479 & ~w1022;
assign w7458 = w5150 & w7580;
assign w7459 = ~w4927 & w7581;
assign w7460 = ~w3472 & w7582;
assign w7461 = w5659 & ~w5281;
assign w7462 = (~w5281 & w5659) | (~w5281 & w7890) | (w5659 & w7890);
assign w7463 = w5659 | ~w5281;
assign w7464 = (w4927 & w7463) | (w4927 & w7583) | (w7463 & w7583);
assign w7465 = w7075 & w5330;
assign w7466 = ~w818 & w847;
assign w7467 = w818 & ~w847;
assign w7468 = ~w1695 & ~w1197;
assign w7469 = ~w3161 | w7106;
assign w7470 = (~w3161 & w5688) | (~w3161 & ~w7502) | (w5688 & ~w7502);
assign w7471 = ~w3175 & w6101;
assign w7472 = w3148 & w2878;
assign w7473 = (w3550 & w7131) | (w3550 & w7584) | (w7131 & w7584);
assign w7474 = w7585 & w6980;
assign w7475 = w6975 & w7585;
assign w7476 = w726 & w7849;
assign w7477 = w1022 & ~w1994;
assign w7478 = (~w3550 & w7213) | (~w3550 & w7588) | (w7213 & w7588);
assign w7479 = (~w5048 & w4970) | (~w5048 & w7698) | (w4970 & w7698);
assign w7480 = (~w5048 & w6439) | (~w5048 & w6421) | (w6439 & w6421);
assign w7481 = (~w5048 & w6439) | (~w5048 & w4978) | (w6439 & w4978);
assign w7482 = w6445 & w6444;
assign w7483 = (~w5111 & w7409) | (~w5111 & ~w5034) | (w7409 & ~w5034);
assign w7484 = (~w5111 & ~w5034) | (~w5111 & w6563) | (~w5034 & w6563);
assign w7485 = ~w5031 & w5843;
assign w7486 = w5031 | w5844;
assign w7487 = ~w5031 & w5845;
assign w7488 = w5031 | w5213;
assign w7489 = w1994 & w7058;
assign w7490 = ~w6274 & w1994;
assign w7491 = (w5214 & ~w5034) | (w5214 & w7417) | (~w5034 & w7417);
assign w7492 = (w5214 & ~w5034) | (w5214 & w6565) | (~w5034 & w6565);
assign w7493 = (~w5137 & w7699) | (~w5137 & w7700) | (w7699 & w7700);
assign w7494 = (w5403 & w7589) | (w5403 & w7741) | (w7589 & w7741);
assign w7495 = ~w5150 & w5178;
assign w7496 = w5150 & w5180;
assign w7497 = ~w5150 & ~w5166;
assign w7498 = ~w818 & ~w871;
assign w7499 = w818 & w871;
assign w7500 = w2835 & ~w3142;
assign w7501 = ~w2835 & w3142;
assign w7502 = w3161 & w3111;
assign w7503 = ~w3161 & ~w3111;
assign w7504 = ~w3161 & ~w6080;
assign w7505 = (~w3148 & w3168) | (~w3148 & w7244) | (w3168 & w7244);
assign w7506 = ~w3175 & ~w6948;
assign w7507 = (w2878 & ~w2171) | (w2878 & w7590) | (~w2171 & w7590);
assign w7508 = ~w7232 & ~w3805;
assign w7509 = w2171 & w7591;
assign w7510 = w7232 & w3805;
assign w7511 = w608 & w2878;
assign w7512 = ~w608 & ~w2878;
assign w7513 = w608 & w3009;
assign w7514 = w7001 & ~w871;
assign w7515 = ~w726 & ~w6994;
assign w7516 = w6482 | w7069;
assign w7517 = w6482 | ~w6835;
assign w7518 = (w7070 & w7516) | (w7070 & w7517) | (w7516 & w7517);
assign w7519 = (w7070 & w7592) | (w7070 & w7593) | (w7592 & w7593);
assign w7520 = w6483 & w7072;
assign w7521 = w6483 & w6835;
assign w7522 = (w7073 & w7520) | (w7073 & w7521) | (w7520 & w7521);
assign w7523 = (w7073 & w7594) | (w7073 & w7595) | (w7594 & w7595);
assign w7524 = w5845 & w7525;
assign w7525 = (w5845 & w6870) | (w5845 & ~w5034) | (w6870 & ~w5034);
assign w7526 = (w5845 & ~w5034) | (w5845 & w7525) | (~w5034 & w7525);
assign w7527 = w6899 & w2734;
assign w7528 = w2734 & w7850;
assign w7529 = (w565 & w5965) | (w565 & w7596) | (w5965 & w7596);
assign w7530 = ~w3780 & w7851;
assign w7531 = ~w3472 & w7530;
assign w7532 = (w4069 & w3472) | (w4069 & w7597) | (w3472 & w7597);
assign w7533 = ~w4404 | w6311;
assign w7534 = (w6488 & w6489) | (w6488 & ~w5034) | (w6489 & ~w5034);
assign w7535 = (w5284 & w7598) | (w5284 & w7599) | (w7598 & w7599);
assign w7536 = (~w5284 & w7600) | (~w5284 & w7601) | (w7600 & w7601);
assign w7537 = w6504 | w5384;
assign w7538 = ~w5425 & ~w3829;
assign w7539 = (~w5425 & ~w5414) | (~w5425 & w7538) | (~w5414 & w7538);
assign w7540 = ~w5400 & w5828;
assign w7541 = w5828 & w7602;
assign w7542 = ~w2878 & ~w7223;
assign w7543 = w3471 & w7104;
assign w7544 = w5687 & w7604;
assign w7545 = ~w3471 & ~w7104;
assign w7546 = (~w3471 & ~w5687) | (~w3471 & w7605) | (~w5687 & w7605);
assign w7547 = w2878 & w7223;
assign w7548 = w3552 & ~w7104;
assign w7549 = w3552 & ~w7103;
assign w7550 = (~w3550 & w7606) | (~w3550 & w7607) | (w7606 & w7607);
assign w7551 = ~w2884 & ~w871;
assign w7552 = ~w6910 & ~w2885;
assign w7553 = ~w1962 | w565;
assign w7554 = ~w2436 & w7111;
assign w7555 = ~w4200 & w6838;
assign w7556 = w6272 & w6838;
assign w7557 = (w3472 & w7608) | (w3472 & w7609) | (w7608 & w7609);
assign w7558 = (w5231 & ~w6489) | (w5231 & w7610) | (~w6489 & w7610);
assign w7559 = w5231 & ~w7331;
assign w7560 = ~w3175 & w7222;
assign w7561 = w3169 & ~w2878;
assign w7562 = (w3550 & w7611) | (w3550 & w7612) | (w7611 & w7612);
assign w7563 = ~w2395 & ~w726;
assign w7564 = ~w7110 & ~w2396;
assign w7565 = w5843 & w7566;
assign w7566 = (w5843 & w6867) | (w5843 & ~w5034) | (w6867 & ~w5034);
assign w7567 = (w5843 & ~w5034) | (w5843 & w7566) | (~w5034 & w7566);
assign w7568 = (w6755 & w7613) | (w6755 & w7614) | (w7613 & w7614);
assign w7569 = (w5844 & w5034) | (w5844 & w6869) | (w5034 & w6869);
assign w7570 = (~w3805 & w7233) | (~w3805 & ~w3175) | (w7233 & ~w3175);
assign w7571 = (~w3805 & w7233) | (~w3805 & w7231) | (w7233 & w7231);
assign w7572 = w3804 & w7615;
assign w7573 = w7235 & ~w7231;
assign w7574 = ~w1994 & ~w7037;
assign w7575 = ~w1994 & ~w1991;
assign w7576 = (w423 & w7701) | (w423 & w7702) | (w7701 & w7702);
assign w7577 = (w423 & w7703) | (w423 & w7704) | (w7703 & w7704);
assign w7578 = ~w1990 & w1022;
assign w7579 = (~w5206 & w4966) | (~w5206 & w7617) | (w4966 & w7617);
assign w7580 = (w5658 & w5152) | (w5658 & w7618) | (w5152 & w7618);
assign w7581 = (w5658 & w4966) | (w5658 & w7619) | (w4966 & w7619);
assign w7582 = w6457 & ~w5277;
assign w7583 = (~w5281 & w5659) | (~w5281 & w4993) | (w5659 & w4993);
assign w7584 = w2878 & ~w6948;
assign w7585 = ~w3936 & w7620;
assign w7586 = ~w2405 | w6384;
assign w7587 = ~w1974 | w6432;
assign w7588 = (w7213 & ~w423) | (w7213 & w7705) | (~w423 & w7705);
assign w7589 = ~w5414 & ~w3829;
assign w7590 = ~w675 & w2878;
assign w7591 = w675 & ~w2878;
assign w7592 = (w6755 & w7621) | (w6755 & w7622) | (w7621 & w7622);
assign w7593 = (w6482 & w5034) | (w6482 & ~w6835) | (w5034 & ~w6835);
assign w7594 = (w6483 & w7072) | (w6483 & ~w5034) | (w7072 & ~w5034);
assign w7595 = (w6483 & ~w5034) | (w6483 & w6835) | (~w5034 & w6835);
assign w7596 = ~w1972 | w565;
assign w7597 = w3551 & w4069;
assign w7598 = ~w5362 & w6866;
assign w7599 = w7074 & w7623;
assign w7600 = w5362 & ~w6866;
assign w7601 = (w5362 & ~w7074) | (w5362 & w7624) | (~w7074 & w7624);
assign w7602 = ~w5277 & ~w5400;
assign w7603 = w5277 & w5400;
assign w7604 = w3111 & w3471;
assign w7605 = ~w3111 & ~w3471;
assign w7606 = ~w2878 & ~w7505;
assign w7607 = (~w2878 & w6948) | (~w2878 & w7620) | (w6948 & w7620);
assign w7608 = (w871 & ~w4313) | (w871 & w7625) | (~w4313 & w7625);
assign w7609 = ~w6990 & w871;
assign w7610 = (w5151 & w7706) | (w5151 & w7707) | (w7706 & w7707);
assign w7611 = w2878 & w7505;
assign w7612 = ~w6948 & w6976;
assign w7613 = (w5844 & w6868) | (w5844 & ~w5032) | (w6868 & ~w5032);
assign w7614 = (w5844 & w6868) | (w5844 & ~w4930) | (w6868 & ~w4930);
assign w7615 = w7509 & w3175;
assign w7616 = ~w5163 & ~w5206;
assign w7617 = w4992 & ~w5206;
assign w7618 = ~w5163 & w5658;
assign w7619 = w4992 & w5658;
assign w7620 = w3175 & ~w2878;
assign w7621 = (w6482 & w7069) | (w6482 & ~w5032) | (w7069 & ~w5032);
assign w7622 = (w6482 & w7069) | (w6482 & ~w4930) | (w7069 & ~w4930);
assign w7623 = ~w5330 & ~w5362;
assign w7624 = w5330 & w5362;
assign w7625 = ~w7001 & w871;
assign w7626 = (w5231 & w5267) | (w5231 & w7627) | (w5267 & w7627);
assign w7627 = w5277 & w5231;
assign w7628 = w3024 & w5615;
assign w7629 = ~w3261 & w6623;
assign w7630 = ~w3261 & w6624;
assign w7631 = w5163 & ~w6456;
assign w7632 = w5163 & w5099;
assign w7633 = ~w6490 & w6491;
assign w7634 = ~w5284 & w7708;
assign w7635 = (w5307 & w6493) | (w5307 & w6490) | (w6493 & w6490);
assign w7636 = ~w6490 & w6567;
assign w7637 = (w5385 & w7840) | (w5385 & w6490) | (w7840 & w6490);
assign w7638 = ~w6490 & w6569;
assign w7639 = ~w6490 & w7347;
assign w7640 = (~w5828 & w5400) | (~w5828 & w7853) | (w5400 & w7853);
assign w7641 = (w5400 & w7348) | (w5400 & w6490) | (w7348 & w6490);
assign w7642 = w3266 & w6111;
assign w7643 = w3266 & w6110;
assign w7644 = (w3472 & w7709) | (w3472 & w7710) | (w7709 & w7710);
assign w7645 = (w3474 & w7477) | (w3474 & w7711) | (w7477 & w7711);
assign w7646 = (w3472 & w7477) | (w3472 & w7712) | (w7477 & w7712);
assign w7647 = (w5278 & w5208) | (w5278 & w7691) | (w5208 & w7691);
assign w7648 = w5278 & w7854;
assign w7649 = ~w5284 & w7713;
assign w7650 = (w7076 & w7077) | (w7076 & w6490) | (w7077 & w6490);
assign w7651 = w5385 & w7840;
assign w7652 = (w5385 & w7651) | (w5385 & w6490) | (w7651 & w6490);
assign w7653 = ~w1022 & w7855;
assign w7654 = ~w1022 & w7891;
assign w7655 = w5139 & ~w5310;
assign w7656 = w6495 & w5330;
assign w7657 = (w5330 & w6495) | (w5330 & ~w5139) | (w6495 & ~w5139);
assign w7658 = w5330 & w7856;
assign w7659 = (w5330 & w7198) | (w5330 & w6490) | (w7198 & w6490);
assign w7660 = ~w5308 & w5330;
assign w7661 = w5139 & w5857;
assign w7662 = w5858 & w5400;
assign w7663 = (w5400 & w5858) | (w5400 & ~w5139) | (w5858 & ~w5139);
assign w7664 = (~w5208 & w7714) | (~w5208 & w7696) | (w7714 & w7696);
assign w7665 = (w7062 & w7696) | (w7062 & w7715) | (w7696 & w7715);
assign w7666 = ~w418 & ~w1022;
assign w7667 = (~w871 & ~w2881) | (~w871 & w7716) | (~w2881 & w7716);
assign w7668 = ~w2882 & w6911;
assign w7669 = w6275 | w6978;
assign w7670 = (w6275 & ~w6975) | (w6275 & w2878) | (~w6975 & w2878);
assign w7671 = (w5108 & w6561) | (w5108 & ~w5034) | (w6561 & ~w5034);
assign w7672 = (w5108 & ~w5034) | (w5108 & w6562) | (~w5034 & w6562);
assign w7673 = (~w5218 & ~w5034) | (~w5218 & w7419) | (~w5034 & w7419);
assign w7674 = (~w5218 & ~w5034) | (~w5218 & w6566) | (~w5034 & w6566);
assign w7675 = ~w2436 & ~w2411;
assign w7676 = w6578 & ~w2411;
assign w7677 = w6578 & ~w6994;
assign w7678 = w2691 & ~w2734;
assign w7679 = w2691 & w6900;
assign w7680 = ~w6490 & w7535;
assign w7681 = w5662 & ~w5362;
assign w7682 = w5362 & w7857;
assign w7683 = (w5362 & w7536) | (w5362 & w6490) | (w7536 & w6490);
assign w7684 = ~w5662 & w5362;
assign w7685 = (w5384 & w6504) | (w5384 & ~w6567) | (w6504 & ~w6567);
assign w7686 = (w5384 & w6504) | (w5384 & ~w7636) | (w6504 & ~w7636);
assign w7687 = (w7538 & w7539) | (w7538 & w6822) | (w7539 & w6822);
assign w7688 = (~w5297 & w7718) | (~w5297 & w7719) | (w7718 & w7719);
assign w7689 = ~w4568 & w6578;
assign w7690 = w6338 & w6578;
assign w7691 = w5278 & w5206;
assign w7692 = (w5278 & ~w5150) | (w5278 & w7720) | (~w5150 & w7720);
assign w7693 = w871 & w7239;
assign w7694 = (~w3550 & w7721) | (~w3550 & w7722) | (w7721 & w7722);
assign w7695 = w5844 | w6869;
assign w7696 = (w5307 & w7202) | (w5307 & ~w5206) | (w7202 & ~w5206);
assign w7697 = (w5150 & w7714) | (w5150 & w7723) | (w7714 & w7723);
assign w7698 = w7045 | ~w5048;
assign w7699 = w7589 & w6822;
assign w7700 = ~w5297 & w7724;
assign w7701 = w7575 & ~w1994;
assign w7702 = (~w1994 & w7575) | (~w1994 & w418) | (w7575 & w418);
assign w7703 = ~w1991 & w1022;
assign w7704 = (w1022 & w7703) | (w1022 & w418) | (w7703 & w418);
assign w7705 = ~w418 & w7213;
assign w7706 = (~w5208 & w7725) | (~w5208 & w7726) | (w7725 & w7726);
assign w7707 = (w7062 & w7726) | (w7062 & w7727) | (w7726 & w7727);
assign w7708 = w7075 & w5307;
assign w7709 = ~w4835 & w7729;
assign w7710 = w6395 & w7729;
assign w7711 = w1022 & w7442;
assign w7712 = (w3550 & w7730) | (w3550 & w7731) | (w7730 & w7731);
assign w7713 = w5330 & w7708;
assign w7714 = (w5307 & w5267) | (w5307 & w7708) | (w5267 & w7708);
assign w7715 = (w5307 & w7202) | (w5307 & w5166) | (w7202 & w5166);
assign w7716 = ~w2875 & ~w871;
assign w7717 = ~w2891 | w6322;
assign w7718 = ~w5425 & w7858;
assign w7719 = (w7538 & w7539) | (w7538 & w5857) | (w7539 & w5857);
assign w7720 = w5278 & w7859;
assign w7721 = w726 & ~w7675;
assign w7722 = (w726 & w6994) | (w726 & w6579) | (w6994 & w6579);
assign w7723 = (w5152 & w7696) | (w5152 & w7742) | (w7696 & w7742);
assign w7724 = w5857 & w7589;
assign w7725 = (w5231 & w5267) | (w5231 & w7732) | (w5267 & w7732);
assign w7726 = (w5231 & w7626) | (w5231 & ~w5206) | (w7626 & ~w5206);
assign w7727 = (w5231 & w7626) | (w5231 & w5166) | (w7626 & w5166);
assign w7728 = w7603 & w5400;
assign w7729 = ~w1963 & ~w565;
assign w7730 = w1022 & w7575;
assign w7731 = w1022 & w7576;
assign w7732 = w7627 & w5231;
assign w7733 = ~w3288 & ~w3275;
assign w7734 = ~w3326 & ~w3331;
assign w7735 = ~w5414 & w6822;
assign w7736 = ~w5297 & w7743;
assign w7737 = w5414 & ~w6822;
assign w7738 = (w5414 & w5297) | (w5414 & w7744) | (w5297 & w7744);
assign w7739 = (w5384 & w6504) | (w5384 & ~w5662) | (w6504 & ~w5662);
assign w7740 = (~w5425 & w7538) | (~w5425 & w5817) | (w7538 & w5817);
assign w7741 = ~w3829 & w5817;
assign w7742 = (w5307 & w7202) | (w5307 & w7616) | (w7202 & w7616);
assign w7743 = w5857 & ~w5414;
assign w7744 = ~w5857 & w5414;
assign w7745 = w1963 & w565;
assign w7746 = (~a_22 & w5876) | (~a_22 & ~w5) | (w5876 & ~w5);
assign w7747 = (~a_22 & w5878) | (~a_22 & ~w2) | (w5878 & ~w2);
assign w7748 = (w2287 & ~w5553) | (w2287 & ~w2117) | (~w5553 & ~w2117);
assign w7749 = (~w2589 & ~w5587) | (~w2589 & ~w2117) | (~w5587 & ~w2117);
assign w7750 = (w2229 & ~w5714) | (w2229 & ~w5715) | (~w5714 & ~w5715);
assign w7751 = (~w2957 & w2389) | (~w2957 & ~w6063) | (w2389 & ~w6063);
assign w7752 = (w2899 & w2866) | (w2899 & w7286) | (w2866 & w7286);
assign w7753 = (~w3189 & w2803) | (~w3189 & ~w5739) | (w2803 & ~w5739);
assign w7754 = (w6917 & w7388) | (w6917 & ~w3203) | (w7388 & ~w3203);
assign w7755 = (w3218 & w7116) | (w3218 & ~w3078) | (w7116 & ~w3078);
assign w7756 = (w7118 & w7390) | (w7118 & ~w2664) | (w7390 & ~w2664);
assign w7757 = (w2878 & w6976) | (w2878 & ~w3269) | (w6976 & ~w3269);
assign w7758 = (w3351 & ~w2878) | (w3351 & w7861) | (~w2878 & w7861);
assign w7759 = (w3359 & w2878) | (w3359 & w7892) | (w2878 & w7892);
assign w7760 = w6839 & ~w3362;
assign w7761 = (w5739 & ~w6095) | (w5739 & ~w6096) | (~w6095 & ~w6096);
assign w7762 = (w6938 & w7353) | (w6938 & ~w3483) | (w7353 & ~w3483);
assign w7763 = (w5739 & ~w6179) | (w5739 & ~w6180) | (~w6179 & ~w6180);
assign w7764 = (w6941 & w7355) | (w6941 & ~w3568) | (w7355 & ~w3568);
assign w7765 = (w3491 & ~w3386) | (w3491 & ~w5754) | (~w3386 & ~w5754);
assign w7766 = (~w3201 & w2803) | (~w3201 & ~w5740) | (w2803 & ~w5740);
assign w7767 = ~w3789 & ~w3790;
assign w7768 = (w3904 & w726) | (w3904 & w7862) | (w726 & w7862);
assign w7769 = (w7125 & w7397) | (w7125 & ~w3483) | (w7397 & ~w3483);
assign w7770 = (w4072 & ~w6257) | (w4072 & ~w4071) | (~w6257 & ~w4071);
assign w7771 = (w6685 & w7365) | (w6685 & ~w3203) | (w7365 & ~w3203);
assign w7772 = (w7142 & w7401) | (w7142 & ~w3568) | (w7401 & ~w3568);
assign w7773 = (~w4734 & ~w6372) | (~w4734 & ~w3348) | (~w6372 & ~w3348);
assign w7774 = (~w4820 & w7151) | (~w4820 & ~w3203) | (w7151 & ~w3203);
assign w7775 = (w3145 & ~w726) | (w3145 & w7319) | (~w726 & w7319);
assign w7776 = (w7032 & w7645) | (w7032 & ~w3483) | (w7645 & ~w3483);
assign w7777 = (~w4978 & ~w6421) | (~w4978 & ~w3568) | (~w6421 & ~w3568);
assign w7778 = (~w3829 & ~w6441) | (~w3829 & ~w5026) | (~w6441 & ~w5026);
assign w7779 = (w6454 & w3829) | (w6454 & ~w5146) | (w3829 & ~w5146);
assign w7780 = (~w3829 & ~w6484) | (~w3829 & ~w5256) | (~w6484 & ~w5256);
assign w7781 = (w3829 & w6487) | (w3829 & ~w5255) | (w6487 & ~w5255);
assign w7782 = (w3829 & w5661) | (w3829 & ~w5295) | (w5661 & ~w5295);
assign w7783 = w7661 & ~w5137;
assign w7784 = (~w2436 & ~w5677) | (~w2436 & ~w1819) | (~w5677 & ~w1819);
assign w7785 = ~w2712 & w2615;
assign w7786 = (~w3009 & ~w5684) | (~w3009 & ~w1819) | (~w5684 & ~w1819);
assign w7787 = (w4949 & ~w5796) | (w4949 & ~w4807) | (~w5796 & ~w4807);
assign w7788 = (~w5033 & ~w5071) | (~w5033 & w7346) | (~w5071 & w7346);
assign w7789 = (a_10 & a_11) | (a_10 & ~a_22) | (a_11 & ~a_22);
assign w7790 = (~w6111 & ~w6110) | (~w6111 & ~w3269) | (~w6110 & ~w3269);
assign w7791 = (w3144 & w3146) | (w3144 & ~w1022) | (w3146 & ~w1022);
assign w7792 = (~w6461 & ~w6462) | (~w6461 & ~w4071) | (~w6462 & ~w4071);
assign w7793 = (~w2712 & w7785) | (~w2712 & ~w2287) | (w7785 & ~w2287);
assign w7794 = (~w2712 & w7785) | (~w2712 & w5553) | (w7785 & w5553);
assign w7795 = w6841 & ~w5057;
assign w7796 = ~w1695 & w6529;
assign w7797 = (w6529 & ~w1695) | (w6529 & ~w1502) | (~w1695 & ~w1502);
assign w7798 = (a_22 & ~w5877) | (a_22 & ~w5876) | (~w5877 & ~w5876);
assign w7799 = w2903 & ~w2410;
assign w7800 = w6921 | ~w3240;
assign w7801 = (~w3240 & w6921) | (~w3240 & ~w2929) | (w6921 & ~w2929);
assign w7802 = (w6962 & ~w6237) | (w6962 & ~w3472) | (~w6237 & ~w3472);
assign w7803 = (~w1022 & w5775) | (~w1022 & ~w4824) | (w5775 & ~w4824);
assign w7804 = (~w4883 & ~w5656) | (~w4883 & ~w4516) | (~w5656 & ~w4516);
assign w7805 = w6440 & w7777;
assign w7806 = (w6444 & w6445) | (w6444 & w7777) | (w6445 & w7777);
assign w7807 = (w7052 & ~w6450) | (w7052 & ~w3472) | (~w6450 & ~w3472);
assign w7808 = (~w1247 & ~w1695) | (~w1247 & w7468) | (~w1695 & w7468);
assign w7809 = (w4200 & ~w6272) | (w4200 & ~w3472) | (~w6272 & ~w3472);
assign w7810 = (~w7001 & w6274) | (~w7001 & ~w3553) | (w6274 & ~w3553);
assign w7811 = (~w7023 & w6274) | (~w7023 & ~w3553) | (w6274 & ~w3553);
assign w7812 = (~w7041 & w6274) | (~w7041 & ~w3553) | (w6274 & ~w3553);
assign w7813 = w7495 & w5178;
assign w7814 = w7497 & ~w5166;
assign w7815 = (w3148 & w6948) | (w3148 & ~w3550) | (w6948 & ~w3550);
assign w7816 = (a_22 & ~w5866) | (a_22 & ~w5865) | (~w5866 & ~w5865);
assign w7817 = w6899 & ~w2677;
assign w7818 = w6901 & ~w2677;
assign w7819 = w7356 | w6949;
assign w7820 = (w6949 & w7356) | (w6949 & w3789) | (w7356 & w3789);
assign w7821 = (w7809 & ~w871) | (w7809 & w6839) | (~w871 & w6839);
assign w7822 = (w7809 & ~w871) | (w7809 & w7863) | (~w871 & w7863);
assign w7823 = (~w6687 & ~w6688) | (~w6687 & ~w5739) | (~w6688 & ~w5739);
assign w7824 = (~w6687 & ~w6688) | (~w6687 & w6095) | (~w6688 & w6095);
assign w7825 = w3782 | ~w3786;
assign w7826 = (~w6710 & ~w6711) | (~w6710 & w6095) | (~w6711 & w6095);
assign w7827 = (w7844 & w726) | (w7844 & w6579) | (w726 & w6579);
assign w7828 = (w7827 & w7402) | (w7827 & w3789) | (w7402 & w3789);
assign w7829 = (~w6727 & ~w6728) | (~w6727 & ~w5739) | (~w6728 & ~w5739);
assign w7830 = (~w6727 & ~w6728) | (~w6727 & w6095) | (~w6728 & w6095);
assign w7831 = (~w6757 & ~w6758) | (~w6757 & ~w5739) | (~w6758 & ~w5739);
assign w7832 = (~w6757 & ~w6758) | (~w6757 & w6095) | (~w6758 & w6095);
assign w7833 = (w6793 & w6794) | (w6793 & ~w5739) | (w6794 & ~w5739);
assign w7834 = (w6793 & w6794) | (w6793 & w6095) | (w6794 & w6095);
assign w7835 = w5034 | ~w4674;
assign w7836 = w7603 & ~w5284;
assign w7837 = (~w7505 & w3175) | (~w7505 & ~w3474) | (w3175 & ~w3474);
assign w7838 = w7431 | w7236;
assign w7839 = (w7236 & w7431) | (w7236 & w3789) | (w7431 & w3789);
assign w7840 = w5385 & ~w6491;
assign w7841 = (~w5057 & w6841) | (~w5057 & w4930) | (w6841 & w4930);
assign w7842 = w7561 & ~w3164;
assign w7843 = (w3175 & ~w7223) | (w3175 & ~w3474) | (~w7223 & ~w3474);
assign w7844 = (w4568 & ~w6338) | (w4568 & ~w3472) | (~w6338 & ~w3472);
assign w7845 = (w4835 & ~w6395) | (w4835 & ~w3472) | (~w6395 & ~w3472);
assign w7846 = w7795 & ~w5057;
assign w7847 = w7496 & ~w5032;
assign w7848 = w7496 & ~w4930;
assign w7849 = (w2411 & w6994) | (w2411 & ~w3550) | (w6994 & ~w3550);
assign w7850 = ~w2731 & w7215;
assign w7851 = w3936 & ~w3551;
assign w7852 = w5163 & ~w5152;
assign w7853 = w7728 & ~w5284;
assign w7854 = (w5206 & ~w5166) | (w5206 & ~w7062) | (~w5166 & ~w7062);
assign w7855 = (w1994 & ~w7442) | (w1994 & ~w3474) | (~w7442 & ~w3474);
assign w7856 = (w7076 & ~w7074) | (w7076 & ~w5284) | (~w7074 & ~w5284);
assign w7857 = (w7601 & ~w6866) | (w7601 & ~w5284) | (~w6866 & ~w5284);
assign w7858 = (~w3829 & w7538) | (~w3829 & ~w5414) | (w7538 & ~w5414);
assign w7859 = (w5206 & ~w7616) | (w5206 & ~w5152) | (~w7616 & ~w5152);
assign w7860 = (~w7575 & ~w7576) | (~w7575 & ~w3550) | (~w7576 & ~w3550);
assign w7861 = w7620 & ~w3348;
assign w7862 = w6579 & ~w3362;
assign w7863 = w6839 & w3789;
assign w7864 = (a_22 & ~w5867) | (a_22 & ~w506) | (~w5867 & ~w506);
assign w7865 = (~a_22 & w5866) | (~a_22 & w506) | (w5866 & w506);
assign w7866 = (~a_22 & w5877) | (~a_22 & w7746) | (w5877 & w7746);
assign w7867 = w7799 | ~w2956;
assign w7868 = (w6922 & w7350) | (w6922 & w2930) | (w7350 & w2930);
assign w7869 = (w7124 & w7396) | (w7124 & w7767) | (w7396 & w7767);
assign w7870 = (w6974 & w7366) | (w6974 & w7767) | (w7366 & w7767);
assign w7871 = (w3782 & w7825) | (w3782 & ~w3788) | (w7825 & ~w3788);
assign w7872 = (w6710 & w6711) | (w6710 & w7761) | (w6711 & w7761);
assign w7873 = (w7008 & w7371) | (w7008 & w7767) | (w7371 & w7767);
assign w7874 = (w6727 & w6728) | (w6727 & w7761) | (w6728 & w7761);
assign w7875 = (w7029 & w7644) | (w7029 & w7767) | (w7644 & w7767);
assign w7876 = (w6757 & w6758) | (w6757 & w7761) | (w6758 & w7761);
assign w7877 = (w7044 & w7646) | (w7044 & w7767) | (w7646 & w7767);
assign w7878 = w7064 & w7893;
assign w7879 = w7071 & ~w5161;
assign w7880 = (w4972 & w7777) | (w4972 & ~w4971) | (w7777 & ~w4971);
assign w7881 = (~w4900 & ~w4898) | (~w4900 & ~w4893) | (~w4898 & ~w4893);
assign w7882 = w2889 & ~w871;
assign w7883 = (~w6710 & ~w6711) | (~w6710 & ~w5739) | (~w6711 & ~w5739);
assign w7884 = (w7845 & w565) | (w7845 & w7745) | (w565 & w7745);
assign w7885 = (w7845 & w565) | (w7845 & w7894) | (w565 & w7894);
assign w7886 = w7654 | w7174;
assign w7887 = (w7174 & w7654) | (w7174 & w3789) | (w7654 & w3789);
assign w7888 = (w3009 & ~w7239) | (w3009 & ~w3474) | (~w7239 & ~w3474);
assign w7889 = (~w5057 & w6841) | (~w5057 & w5032) | (w6841 & w5032);
assign w7890 = w7852 | ~w5150;
assign w7891 = (w1994 & w7860) | (w1994 & ~w3472) | (w7860 & ~w3472);
assign w7892 = w7115 & ~w3362;
assign w7893 = (~w6793 & ~w6794) | (~w6793 & w7761) | (~w6794 & w7761);
assign w7894 = w7745 & w3789;
assign one = 1;
assign sin_0 = w3826;// level 74
assign sin_1 = ~w3971;// level 77
assign sin_2 = ~w4129;// level 78
assign sin_3 = ~w4257;// level 80
assign sin_4 = ~w4373;// level 81
assign sin_5 = ~w4489;// level 83
assign sin_6 = ~w4605;// level 84
assign sin_7 = ~w4709;// level 85
assign sin_8 = ~w4802;// level 86
assign sin_9 = ~w4882;// level 86
assign sin_10 = ~w4962;// level 87
assign sin_11 = w5029;// level 88
assign sin_12 = w5083;// level 89
assign sin_13 = w5149;// level 89
assign sin_14 = w5201;// level 90
assign sin_15 = w5259;// level 90
assign sin_16 = ~w5293;// level 91
assign sin_17 = w5319;// level 91
assign sin_18 = ~w5354;// level 91
assign sin_19 = w5374;// level 91
assign sin_20 = ~w5395;// level 91
assign sin_21 = w5413;// level 91
assign sin_22 = ~w5423;// level 91
assign sin_23 = ~w5430;// level 91
assign sin_24 = w5432;// level 91
endmodule

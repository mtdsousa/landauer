module bar_best_speed (
        a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, a_64, a_65, a_66, a_67, a_68, a_69, a_70, a_71, a_72, a_73, a_74, a_75, a_76, a_77, a_78, a_79, a_80, a_81, a_82, a_83, a_84, a_85, a_86, a_87, a_88, a_89, a_90, a_91, a_92, a_93, a_94, a_95, a_96, a_97, a_98, a_99, a_100, a_101, a_102, a_103, a_104, a_105, a_106, a_107, a_108, a_109, a_110, a_111, a_112, a_113, a_114, a_115, a_116, a_117, a_118, a_119, a_120, a_121, a_122, a_123, a_124, a_125, a_126, a_127, shift_0, shift_1, shift_2, shift_3, shift_4, shift_5, shift_6, 
        result_0, result_1, result_2, result_3, result_4, result_5, result_6, result_7, result_8, result_9, result_10, result_11, result_12, result_13, result_14, result_15, result_16, result_17, result_18, result_19, result_20, result_21, result_22, result_23, result_24, result_25, result_26, result_27, result_28, result_29, result_30, result_31, result_32, result_33, result_34, result_35, result_36, result_37, result_38, result_39, result_40, result_41, result_42, result_43, result_44, result_45, result_46, result_47, result_48, result_49, result_50, result_51, result_52, result_53, result_54, result_55, result_56, result_57, result_58, result_59, result_60, result_61, result_62, result_63, result_64, result_65, result_66, result_67, result_68, result_69, result_70, result_71, result_72, result_73, result_74, result_75, result_76, result_77, result_78, result_79, result_80, result_81, result_82, result_83, result_84, result_85, result_86, result_87, result_88, result_89, result_90, result_91, result_92, result_93, result_94, result_95, result_96, result_97, result_98, result_99, result_100, result_101, result_102, result_103, result_104, result_105, result_106, result_107, result_108, result_109, result_110, result_111, result_112, result_113, result_114, result_115, result_116, result_117, result_118, result_119, result_120, result_121, result_122, result_123, result_124, result_125, result_126, result_127);
input a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, a_64, a_65, a_66, a_67, a_68, a_69, a_70, a_71, a_72, a_73, a_74, a_75, a_76, a_77, a_78, a_79, a_80, a_81, a_82, a_83, a_84, a_85, a_86, a_87, a_88, a_89, a_90, a_91, a_92, a_93, a_94, a_95, a_96, a_97, a_98, a_99, a_100, a_101, a_102, a_103, a_104, a_105, a_106, a_107, a_108, a_109, a_110, a_111, a_112, a_113, a_114, a_115, a_116, a_117, a_118, a_119, a_120, a_121, a_122, a_123, a_124, a_125, a_126, a_127, shift_0, shift_1, shift_2, shift_3, shift_4, shift_5, shift_6;
output result_0, result_1, result_2, result_3, result_4, result_5, result_6, result_7, result_8, result_9, result_10, result_11, result_12, result_13, result_14, result_15, result_16, result_17, result_18, result_19, result_20, result_21, result_22, result_23, result_24, result_25, result_26, result_27, result_28, result_29, result_30, result_31, result_32, result_33, result_34, result_35, result_36, result_37, result_38, result_39, result_40, result_41, result_42, result_43, result_44, result_45, result_46, result_47, result_48, result_49, result_50, result_51, result_52, result_53, result_54, result_55, result_56, result_57, result_58, result_59, result_60, result_61, result_62, result_63, result_64, result_65, result_66, result_67, result_68, result_69, result_70, result_71, result_72, result_73, result_74, result_75, result_76, result_77, result_78, result_79, result_80, result_81, result_82, result_83, result_84, result_85, result_86, result_87, result_88, result_89, result_90, result_91, result_92, result_93, result_94, result_95, result_96, result_97, result_98, result_99, result_100, result_101, result_102, result_103, result_104, result_105, result_106, result_107, result_108, result_109, result_110, result_111, result_112, result_113, result_114, result_115, result_116, result_117, result_118, result_119, result_120, result_121, result_122, result_123, result_124, result_125, result_126, result_127;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053;
assign w0 = ~a_64 & ~shift_1;
assign w1 = ~a_62 & shift_1;
assign w2 = ~w0 & ~w1;
assign w3 = ~shift_0 & ~w2;
assign w4 = ~a_63 & ~shift_1;
assign w5 = ~a_61 & shift_1;
assign w6 = ~w4 & ~w5;
assign w7 = shift_0 & ~w6;
assign w8 = ~w3 & ~w7;
assign w9 = ~shift_3 & ~w8;
assign w10 = ~a_56 & ~shift_1;
assign w11 = ~a_54 & shift_1;
assign w12 = ~w10 & ~w11;
assign w13 = ~shift_0 & ~w12;
assign w14 = ~a_55 & ~shift_1;
assign w15 = ~a_53 & shift_1;
assign w16 = ~w14 & ~w15;
assign w17 = shift_0 & ~w16;
assign w18 = ~w13 & ~w17;
assign w19 = shift_3 & ~w18;
assign w20 = ~w9 & ~w19;
assign w21 = ~shift_2 & ~w20;
assign w22 = ~a_60 & ~shift_1;
assign w23 = ~a_58 & shift_1;
assign w24 = ~w22 & ~w23;
assign w25 = ~shift_0 & ~w24;
assign w26 = ~a_59 & ~shift_1;
assign w27 = ~a_57 & shift_1;
assign w28 = ~w26 & ~w27;
assign w29 = shift_0 & ~w28;
assign w30 = ~w25 & ~w29;
assign w31 = ~shift_3 & ~w30;
assign w32 = ~a_52 & ~shift_1;
assign w33 = ~a_50 & shift_1;
assign w34 = ~w32 & ~w33;
assign w35 = ~shift_0 & ~w34;
assign w36 = ~a_51 & ~shift_1;
assign w37 = ~a_49 & shift_1;
assign w38 = ~w36 & ~w37;
assign w39 = shift_0 & ~w38;
assign w40 = ~w35 & ~w39;
assign w41 = shift_3 & ~w40;
assign w42 = ~w31 & ~w41;
assign w43 = shift_2 & ~w42;
assign w44 = ~w21 & ~w43;
assign w45 = ~shift_5 & ~w44;
assign w46 = ~a_32 & ~shift_1;
assign w47 = ~a_30 & shift_1;
assign w48 = ~w46 & ~w47;
assign w49 = ~shift_0 & ~w48;
assign w50 = ~a_31 & ~shift_1;
assign w51 = ~a_29 & shift_1;
assign w52 = ~w50 & ~w51;
assign w53 = shift_0 & ~w52;
assign w54 = ~w49 & ~w53;
assign w55 = ~shift_3 & ~w54;
assign w56 = ~a_24 & ~shift_1;
assign w57 = ~a_22 & shift_1;
assign w58 = ~w56 & ~w57;
assign w59 = ~shift_0 & ~w58;
assign w60 = ~a_23 & ~shift_1;
assign w61 = ~a_21 & shift_1;
assign w62 = ~w60 & ~w61;
assign w63 = shift_0 & ~w62;
assign w64 = ~w59 & ~w63;
assign w65 = shift_3 & ~w64;
assign w66 = ~w55 & ~w65;
assign w67 = ~shift_2 & ~w66;
assign w68 = ~a_28 & ~shift_1;
assign w69 = ~a_26 & shift_1;
assign w70 = ~w68 & ~w69;
assign w71 = ~shift_0 & ~w70;
assign w72 = ~a_27 & ~shift_1;
assign w73 = ~a_25 & shift_1;
assign w74 = ~w72 & ~w73;
assign w75 = shift_0 & ~w74;
assign w76 = ~w71 & ~w75;
assign w77 = ~shift_3 & ~w76;
assign w78 = ~a_20 & ~shift_1;
assign w79 = ~a_18 & shift_1;
assign w80 = ~w78 & ~w79;
assign w81 = ~shift_0 & ~w80;
assign w82 = ~a_19 & ~shift_1;
assign w83 = ~a_17 & shift_1;
assign w84 = ~w82 & ~w83;
assign w85 = shift_0 & ~w84;
assign w86 = ~w81 & ~w85;
assign w87 = shift_3 & ~w86;
assign w88 = ~w77 & ~w87;
assign w89 = shift_2 & ~w88;
assign w90 = ~w67 & ~w89;
assign w91 = shift_5 & ~w90;
assign w92 = ~w45 & ~w91;
assign w93 = ~shift_4 & ~w92;
assign w94 = a_38 & shift_1;
assign w95 = a_40 & ~shift_1;
assign w96 = ~w94 & ~w95;
assign w97 = ~shift_0 & ~w96;
assign w98 = a_39 & ~shift_1;
assign w99 = a_37 & shift_1;
assign w100 = ~w98 & ~w99;
assign w101 = shift_0 & ~w100;
assign w102 = ~w97 & ~w101;
assign w103 = shift_3 & w102;
assign w104 = ~a_48 & ~shift_1;
assign w105 = ~a_46 & shift_1;
assign w106 = ~w104 & ~w105;
assign w107 = ~shift_0 & ~w106;
assign w108 = ~a_47 & ~shift_1;
assign w109 = ~a_45 & shift_1;
assign w110 = ~w108 & ~w109;
assign w111 = shift_0 & ~w110;
assign w112 = ~w107 & ~w111;
assign w113 = ~shift_3 & ~w112;
assign w114 = ~w103 & ~w113;
assign w115 = ~shift_2 & ~w114;
assign w116 = ~a_44 & ~shift_1;
assign w117 = ~a_42 & shift_1;
assign w118 = ~w116 & ~w117;
assign w119 = ~shift_0 & ~w118;
assign w120 = ~a_43 & ~shift_1;
assign w121 = ~a_41 & shift_1;
assign w122 = ~w120 & ~w121;
assign w123 = shift_0 & ~w122;
assign w124 = ~w119 & ~w123;
assign w125 = ~shift_3 & ~w124;
assign w126 = ~a_36 & ~shift_1;
assign w127 = ~a_34 & shift_1;
assign w128 = ~w126 & ~w127;
assign w129 = ~shift_0 & ~w128;
assign w130 = ~a_35 & ~shift_1;
assign w131 = ~a_33 & shift_1;
assign w132 = ~w130 & ~w131;
assign w133 = shift_0 & ~w132;
assign w134 = ~w129 & ~w133;
assign w135 = shift_3 & ~w134;
assign w136 = ~w125 & ~w135;
assign w137 = shift_2 & ~w136;
assign w138 = ~w115 & ~w137;
assign w139 = ~shift_5 & ~w138;
assign w140 = ~a_16 & ~shift_1;
assign w141 = ~a_14 & shift_1;
assign w142 = ~w140 & ~w141;
assign w143 = ~shift_0 & ~w142;
assign w144 = ~a_15 & ~shift_1;
assign w145 = ~a_13 & shift_1;
assign w146 = ~w144 & ~w145;
assign w147 = shift_0 & ~w146;
assign w148 = ~w143 & ~w147;
assign w149 = ~shift_3 & ~w148;
assign w150 = ~a_8 & ~shift_1;
assign w151 = ~a_6 & shift_1;
assign w152 = ~w150 & ~w151;
assign w153 = ~shift_0 & ~w152;
assign w154 = ~a_7 & ~shift_1;
assign w155 = ~a_5 & shift_1;
assign w156 = ~w154 & ~w155;
assign w157 = shift_0 & ~w156;
assign w158 = ~w153 & ~w157;
assign w159 = shift_3 & ~w158;
assign w160 = ~w149 & ~w159;
assign w161 = ~shift_2 & ~w160;
assign w162 = ~a_12 & ~shift_1;
assign w163 = ~a_10 & shift_1;
assign w164 = ~w162 & ~w163;
assign w165 = ~shift_0 & ~w164;
assign w166 = ~a_11 & ~shift_1;
assign w167 = ~a_9 & shift_1;
assign w168 = ~w166 & ~w167;
assign w169 = shift_0 & ~w168;
assign w170 = ~w165 & ~w169;
assign w171 = ~shift_3 & ~w170;
assign w172 = ~a_4 & ~shift_1;
assign w173 = ~a_2 & shift_1;
assign w174 = ~w172 & ~w173;
assign w175 = ~shift_0 & ~w174;
assign w176 = ~a_3 & ~shift_1;
assign w177 = ~a_1 & shift_1;
assign w178 = ~w176 & ~w177;
assign w179 = shift_0 & ~w178;
assign w180 = ~w175 & ~w179;
assign w181 = shift_3 & ~w180;
assign w182 = ~w171 & ~w181;
assign w183 = shift_2 & ~w182;
assign w184 = ~w161 & ~w183;
assign w185 = shift_5 & ~w184;
assign w186 = ~w139 & ~w185;
assign w187 = shift_4 & ~w186;
assign w188 = ~w93 & ~w187;
assign w189 = shift_6 & w188;
assign w190 = ~a_0 & ~shift_1;
assign w191 = ~a_126 & shift_1;
assign w192 = ~w190 & ~w191;
assign w193 = ~shift_0 & ~w192;
assign w194 = ~a_127 & ~shift_1;
assign w195 = ~a_125 & shift_1;
assign w196 = ~w194 & ~w195;
assign w197 = shift_0 & ~w196;
assign w198 = ~w193 & ~w197;
assign w199 = ~shift_3 & ~w198;
assign w200 = ~a_120 & ~shift_1;
assign w201 = ~a_118 & shift_1;
assign w202 = ~w200 & ~w201;
assign w203 = ~shift_0 & ~w202;
assign w204 = ~a_119 & ~shift_1;
assign w205 = ~a_117 & shift_1;
assign w206 = ~w204 & ~w205;
assign w207 = shift_0 & ~w206;
assign w208 = ~w203 & ~w207;
assign w209 = shift_3 & ~w208;
assign w210 = ~w199 & ~w209;
assign w211 = ~shift_2 & ~w210;
assign w212 = ~a_124 & ~shift_1;
assign w213 = ~a_122 & shift_1;
assign w214 = ~w212 & ~w213;
assign w215 = ~shift_0 & ~w214;
assign w216 = ~a_123 & ~shift_1;
assign w217 = ~a_121 & shift_1;
assign w218 = ~w216 & ~w217;
assign w219 = shift_0 & ~w218;
assign w220 = ~w215 & ~w219;
assign w221 = ~shift_3 & ~w220;
assign w222 = ~a_116 & ~shift_1;
assign w223 = ~a_114 & shift_1;
assign w224 = ~w222 & ~w223;
assign w225 = ~shift_0 & ~w224;
assign w226 = ~a_115 & ~shift_1;
assign w227 = ~a_113 & shift_1;
assign w228 = ~w226 & ~w227;
assign w229 = shift_0 & ~w228;
assign w230 = ~w225 & ~w229;
assign w231 = shift_3 & ~w230;
assign w232 = ~w221 & ~w231;
assign w233 = shift_2 & ~w232;
assign w234 = ~w211 & ~w233;
assign w235 = ~shift_5 & ~w234;
assign w236 = ~a_96 & ~shift_1;
assign w237 = ~a_94 & shift_1;
assign w238 = ~w236 & ~w237;
assign w239 = ~shift_0 & ~w238;
assign w240 = ~a_95 & ~shift_1;
assign w241 = ~a_93 & shift_1;
assign w242 = ~w240 & ~w241;
assign w243 = shift_0 & ~w242;
assign w244 = ~w239 & ~w243;
assign w245 = ~shift_3 & ~w244;
assign w246 = ~a_88 & ~shift_1;
assign w247 = ~a_86 & shift_1;
assign w248 = ~w246 & ~w247;
assign w249 = ~shift_0 & ~w248;
assign w250 = ~a_87 & ~shift_1;
assign w251 = ~a_85 & shift_1;
assign w252 = ~w250 & ~w251;
assign w253 = shift_0 & ~w252;
assign w254 = ~w249 & ~w253;
assign w255 = shift_3 & ~w254;
assign w256 = ~w245 & ~w255;
assign w257 = ~shift_2 & ~w256;
assign w258 = ~a_92 & ~shift_1;
assign w259 = ~a_90 & shift_1;
assign w260 = ~w258 & ~w259;
assign w261 = ~shift_0 & ~w260;
assign w262 = ~a_91 & ~shift_1;
assign w263 = ~a_89 & shift_1;
assign w264 = ~w262 & ~w263;
assign w265 = shift_0 & ~w264;
assign w266 = ~w261 & ~w265;
assign w267 = ~shift_3 & ~w266;
assign w268 = ~a_84 & ~shift_1;
assign w269 = ~a_82 & shift_1;
assign w270 = ~w268 & ~w269;
assign w271 = ~shift_0 & ~w270;
assign w272 = ~a_83 & ~shift_1;
assign w273 = ~a_81 & shift_1;
assign w274 = ~w272 & ~w273;
assign w275 = shift_0 & ~w274;
assign w276 = ~w271 & ~w275;
assign w277 = shift_3 & ~w276;
assign w278 = ~w267 & ~w277;
assign w279 = shift_2 & ~w278;
assign w280 = ~w257 & ~w279;
assign w281 = shift_5 & ~w280;
assign w282 = ~w235 & ~w281;
assign w283 = ~shift_4 & ~w282;
assign w284 = ~a_112 & ~shift_1;
assign w285 = ~a_110 & shift_1;
assign w286 = ~w284 & ~w285;
assign w287 = ~shift_0 & ~w286;
assign w288 = ~a_111 & ~shift_1;
assign w289 = ~a_109 & shift_1;
assign w290 = ~w288 & ~w289;
assign w291 = shift_0 & ~w290;
assign w292 = ~w287 & ~w291;
assign w293 = ~shift_3 & ~w292;
assign w294 = ~a_104 & ~shift_1;
assign w295 = ~a_102 & shift_1;
assign w296 = ~w294 & ~w295;
assign w297 = ~shift_0 & ~w296;
assign w298 = ~a_103 & ~shift_1;
assign w299 = ~a_101 & shift_1;
assign w300 = ~w298 & ~w299;
assign w301 = shift_0 & ~w300;
assign w302 = ~w297 & ~w301;
assign w303 = shift_3 & ~w302;
assign w304 = ~w293 & ~w303;
assign w305 = ~shift_2 & ~w304;
assign w306 = ~a_108 & ~shift_1;
assign w307 = ~a_106 & shift_1;
assign w308 = ~w306 & ~w307;
assign w309 = ~shift_0 & ~w308;
assign w310 = ~a_107 & ~shift_1;
assign w311 = ~a_105 & shift_1;
assign w312 = ~w310 & ~w311;
assign w313 = shift_0 & ~w312;
assign w314 = ~w309 & ~w313;
assign w315 = ~shift_3 & ~w314;
assign w316 = ~a_100 & ~shift_1;
assign w317 = ~a_98 & shift_1;
assign w318 = ~w316 & ~w317;
assign w319 = ~shift_0 & ~w318;
assign w320 = ~a_99 & ~shift_1;
assign w321 = ~a_97 & shift_1;
assign w322 = ~w320 & ~w321;
assign w323 = shift_0 & ~w322;
assign w324 = ~w319 & ~w323;
assign w325 = shift_3 & ~w324;
assign w326 = ~w315 & ~w325;
assign w327 = shift_2 & ~w326;
assign w328 = ~w305 & ~w327;
assign w329 = ~shift_5 & ~w328;
assign w330 = ~a_80 & ~shift_1;
assign w331 = ~a_78 & shift_1;
assign w332 = ~w330 & ~w331;
assign w333 = ~shift_0 & ~w332;
assign w334 = ~a_79 & ~shift_1;
assign w335 = ~a_77 & shift_1;
assign w336 = ~w334 & ~w335;
assign w337 = shift_0 & ~w336;
assign w338 = ~w333 & ~w337;
assign w339 = ~shift_3 & ~w338;
assign w340 = ~a_72 & ~shift_1;
assign w341 = ~a_70 & shift_1;
assign w342 = ~w340 & ~w341;
assign w343 = ~shift_0 & ~w342;
assign w344 = ~a_71 & ~shift_1;
assign w345 = ~a_69 & shift_1;
assign w346 = ~w344 & ~w345;
assign w347 = shift_0 & ~w346;
assign w348 = ~w343 & ~w347;
assign w349 = shift_3 & ~w348;
assign w350 = ~w339 & ~w349;
assign w351 = ~shift_2 & ~w350;
assign w352 = ~a_76 & ~shift_1;
assign w353 = ~a_74 & shift_1;
assign w354 = ~w352 & ~w353;
assign w355 = ~shift_0 & ~w354;
assign w356 = ~a_75 & ~shift_1;
assign w357 = ~a_73 & shift_1;
assign w358 = ~w356 & ~w357;
assign w359 = shift_0 & ~w358;
assign w360 = ~w355 & ~w359;
assign w361 = ~shift_3 & ~w360;
assign w362 = ~a_68 & ~shift_1;
assign w363 = ~a_66 & shift_1;
assign w364 = ~w362 & ~w363;
assign w365 = ~shift_0 & ~w364;
assign w366 = ~a_67 & ~shift_1;
assign w367 = ~a_65 & shift_1;
assign w368 = ~w366 & ~w367;
assign w369 = shift_0 & ~w368;
assign w370 = ~w365 & ~w369;
assign w371 = shift_3 & ~w370;
assign w372 = ~w361 & ~w371;
assign w373 = shift_2 & ~w372;
assign w374 = ~w351 & ~w373;
assign w375 = shift_5 & ~w374;
assign w376 = ~w329 & ~w375;
assign w377 = shift_4 & ~w376;
assign w378 = ~w283 & ~w377;
assign w379 = ~shift_6 & w378;
assign w380 = ~w189 & ~w379;
assign w381 = a_47 & shift_1;
assign w382 = a_49 & ~shift_1;
assign w383 = ~w381 & ~w382;
assign w384 = ~shift_0 & ~w383;
assign w385 = a_48 & ~shift_1;
assign w386 = a_46 & shift_1;
assign w387 = ~w385 & ~w386;
assign w388 = shift_0 & ~w387;
assign w389 = ~w384 & ~w388;
assign w390 = ~shift_3 & w389;
assign w391 = ~a_41 & ~shift_1;
assign w392 = ~a_39 & shift_1;
assign w393 = ~w391 & ~w392;
assign w394 = ~shift_0 & ~w393;
assign w395 = ~a_40 & ~shift_1;
assign w396 = ~a_38 & shift_1;
assign w397 = ~w395 & ~w396;
assign w398 = shift_0 & ~w397;
assign w399 = ~w394 & ~w398;
assign w400 = shift_3 & ~w399;
assign w401 = ~w390 & ~w400;
assign w402 = ~shift_2 & ~w401;
assign w403 = a_35 & shift_1;
assign w404 = a_37 & ~shift_1;
assign w405 = ~w403 & ~w404;
assign w406 = ~shift_0 & ~w405;
assign w407 = a_36 & ~shift_1;
assign w408 = a_34 & shift_1;
assign w409 = ~w407 & ~w408;
assign w410 = shift_0 & ~w409;
assign w411 = ~w406 & ~w410;
assign w412 = shift_3 & w411;
assign w413 = ~a_45 & ~shift_1;
assign w414 = ~a_43 & shift_1;
assign w415 = ~w413 & ~w414;
assign w416 = ~shift_0 & ~w415;
assign w417 = shift_0 & ~w118;
assign w418 = ~w416 & ~w417;
assign w419 = ~shift_3 & ~w418;
assign w420 = ~w412 & ~w419;
assign w421 = shift_2 & ~w420;
assign w422 = ~w402 & ~w421;
assign w423 = ~shift_5 & ~w422;
assign w424 = a_15 & shift_1;
assign w425 = a_17 & ~shift_1;
assign w426 = ~w424 & ~w425;
assign w427 = ~shift_0 & ~w426;
assign w428 = a_16 & ~shift_1;
assign w429 = a_14 & shift_1;
assign w430 = ~w428 & ~w429;
assign w431 = shift_0 & ~w430;
assign w432 = ~w427 & ~w431;
assign w433 = ~shift_3 & w432;
assign w434 = a_7 & shift_1;
assign w435 = a_9 & ~shift_1;
assign w436 = ~w434 & ~w435;
assign w437 = ~shift_0 & ~w436;
assign w438 = a_8 & ~shift_1;
assign w439 = a_6 & shift_1;
assign w440 = ~w438 & ~w439;
assign w441 = shift_0 & ~w440;
assign w442 = ~w437 & ~w441;
assign w443 = shift_3 & w442;
assign w444 = ~w433 & ~w443;
assign w445 = ~shift_2 & ~w444;
assign w446 = a_11 & shift_1;
assign w447 = a_13 & ~shift_1;
assign w448 = ~w446 & ~w447;
assign w449 = ~shift_0 & ~w448;
assign w450 = a_12 & ~shift_1;
assign w451 = a_10 & shift_1;
assign w452 = ~w450 & ~w451;
assign w453 = shift_0 & ~w452;
assign w454 = ~w449 & ~w453;
assign w455 = ~shift_3 & w454;
assign w456 = a_3 & shift_1;
assign w457 = a_5 & ~shift_1;
assign w458 = ~w456 & ~w457;
assign w459 = ~shift_0 & ~w458;
assign w460 = a_4 & ~shift_1;
assign w461 = a_2 & shift_1;
assign w462 = ~w460 & ~w461;
assign w463 = shift_0 & ~w462;
assign w464 = ~w459 & ~w463;
assign w465 = shift_3 & w464;
assign w466 = ~w455 & ~w465;
assign w467 = shift_2 & ~w466;
assign w468 = ~w445 & ~w467;
assign w469 = shift_5 & ~w468;
assign w470 = ~w423 & ~w469;
assign w471 = shift_4 & ~w470;
assign w472 = a_63 & shift_1;
assign w473 = a_65 & ~shift_1;
assign w474 = ~w472 & ~w473;
assign w475 = ~shift_0 & ~w474;
assign w476 = a_64 & ~shift_1;
assign w477 = a_62 & shift_1;
assign w478 = ~w476 & ~w477;
assign w479 = shift_0 & ~w478;
assign w480 = ~w475 & ~w479;
assign w481 = ~shift_3 & w480;
assign w482 = a_55 & shift_1;
assign w483 = a_57 & ~shift_1;
assign w484 = ~w482 & ~w483;
assign w485 = ~shift_0 & ~w484;
assign w486 = a_56 & ~shift_1;
assign w487 = a_54 & shift_1;
assign w488 = ~w486 & ~w487;
assign w489 = shift_0 & ~w488;
assign w490 = ~w485 & ~w489;
assign w491 = shift_3 & w490;
assign w492 = ~w481 & ~w491;
assign w493 = ~shift_2 & ~w492;
assign w494 = a_59 & shift_1;
assign w495 = a_61 & ~shift_1;
assign w496 = ~w494 & ~w495;
assign w497 = ~shift_0 & ~w496;
assign w498 = a_60 & ~shift_1;
assign w499 = a_58 & shift_1;
assign w500 = ~w498 & ~w499;
assign w501 = shift_0 & ~w500;
assign w502 = ~w497 & ~w501;
assign w503 = ~shift_3 & w502;
assign w504 = a_51 & shift_1;
assign w505 = a_53 & ~shift_1;
assign w506 = ~w504 & ~w505;
assign w507 = ~shift_0 & ~w506;
assign w508 = a_52 & ~shift_1;
assign w509 = a_50 & shift_1;
assign w510 = ~w508 & ~w509;
assign w511 = shift_0 & ~w510;
assign w512 = ~w507 & ~w511;
assign w513 = shift_3 & w512;
assign w514 = ~w503 & ~w513;
assign w515 = shift_2 & ~w514;
assign w516 = ~w493 & ~w515;
assign w517 = ~shift_5 & ~w516;
assign w518 = a_31 & shift_1;
assign w519 = a_33 & ~shift_1;
assign w520 = ~w518 & ~w519;
assign w521 = ~shift_0 & ~w520;
assign w522 = a_32 & ~shift_1;
assign w523 = a_30 & shift_1;
assign w524 = ~w522 & ~w523;
assign w525 = shift_0 & ~w524;
assign w526 = ~w521 & ~w525;
assign w527 = ~shift_3 & w526;
assign w528 = a_23 & shift_1;
assign w529 = a_25 & ~shift_1;
assign w530 = ~w528 & ~w529;
assign w531 = ~shift_0 & ~w530;
assign w532 = a_24 & ~shift_1;
assign w533 = a_22 & shift_1;
assign w534 = ~w532 & ~w533;
assign w535 = shift_0 & ~w534;
assign w536 = ~w531 & ~w535;
assign w537 = shift_3 & w536;
assign w538 = ~w527 & ~w537;
assign w539 = ~shift_2 & ~w538;
assign w540 = a_27 & shift_1;
assign w541 = a_29 & ~shift_1;
assign w542 = ~w540 & ~w541;
assign w543 = ~shift_0 & ~w542;
assign w544 = a_28 & ~shift_1;
assign w545 = a_26 & shift_1;
assign w546 = ~w544 & ~w545;
assign w547 = shift_0 & ~w546;
assign w548 = ~w543 & ~w547;
assign w549 = ~shift_3 & w548;
assign w550 = a_19 & shift_1;
assign w551 = a_21 & ~shift_1;
assign w552 = ~w550 & ~w551;
assign w553 = ~shift_0 & ~w552;
assign w554 = a_20 & ~shift_1;
assign w555 = a_18 & shift_1;
assign w556 = ~w554 & ~w555;
assign w557 = shift_0 & ~w556;
assign w558 = ~w553 & ~w557;
assign w559 = shift_3 & w558;
assign w560 = ~w549 & ~w559;
assign w561 = shift_2 & ~w560;
assign w562 = ~w539 & ~w561;
assign w563 = shift_5 & ~w562;
assign w564 = ~w517 & ~w563;
assign w565 = ~shift_4 & ~w564;
assign w566 = ~w471 & ~w565;
assign w567 = shift_6 & w566;
assign w568 = a_127 & shift_1;
assign w569 = a_1 & ~shift_1;
assign w570 = ~w568 & ~w569;
assign w571 = ~shift_0 & ~w570;
assign w572 = a_0 & ~shift_1;
assign w573 = a_126 & shift_1;
assign w574 = ~w572 & ~w573;
assign w575 = shift_0 & ~w574;
assign w576 = ~w571 & ~w575;
assign w577 = ~shift_3 & w576;
assign w578 = a_119 & shift_1;
assign w579 = a_121 & ~shift_1;
assign w580 = ~w578 & ~w579;
assign w581 = ~shift_0 & ~w580;
assign w582 = a_120 & ~shift_1;
assign w583 = a_118 & shift_1;
assign w584 = ~w582 & ~w583;
assign w585 = shift_0 & ~w584;
assign w586 = ~w581 & ~w585;
assign w587 = shift_3 & w586;
assign w588 = ~w577 & ~w587;
assign w589 = ~shift_2 & ~w588;
assign w590 = a_123 & shift_1;
assign w591 = a_125 & ~shift_1;
assign w592 = ~w590 & ~w591;
assign w593 = ~shift_0 & ~w592;
assign w594 = a_124 & ~shift_1;
assign w595 = a_122 & shift_1;
assign w596 = ~w594 & ~w595;
assign w597 = shift_0 & ~w596;
assign w598 = ~w593 & ~w597;
assign w599 = ~shift_3 & w598;
assign w600 = a_115 & shift_1;
assign w601 = a_117 & ~shift_1;
assign w602 = ~w600 & ~w601;
assign w603 = ~shift_0 & ~w602;
assign w604 = a_116 & ~shift_1;
assign w605 = a_114 & shift_1;
assign w606 = ~w604 & ~w605;
assign w607 = shift_0 & ~w606;
assign w608 = ~w603 & ~w607;
assign w609 = shift_3 & w608;
assign w610 = ~w599 & ~w609;
assign w611 = shift_2 & ~w610;
assign w612 = ~w589 & ~w611;
assign w613 = ~shift_5 & ~w612;
assign w614 = a_95 & shift_1;
assign w615 = a_97 & ~shift_1;
assign w616 = ~w614 & ~w615;
assign w617 = ~shift_0 & ~w616;
assign w618 = a_96 & ~shift_1;
assign w619 = a_94 & shift_1;
assign w620 = ~w618 & ~w619;
assign w621 = shift_0 & ~w620;
assign w622 = ~w617 & ~w621;
assign w623 = ~shift_3 & w622;
assign w624 = a_87 & shift_1;
assign w625 = a_89 & ~shift_1;
assign w626 = ~w624 & ~w625;
assign w627 = ~shift_0 & ~w626;
assign w628 = a_88 & ~shift_1;
assign w629 = a_86 & shift_1;
assign w630 = ~w628 & ~w629;
assign w631 = shift_0 & ~w630;
assign w632 = ~w627 & ~w631;
assign w633 = shift_3 & w632;
assign w634 = ~w623 & ~w633;
assign w635 = ~shift_2 & ~w634;
assign w636 = a_91 & shift_1;
assign w637 = a_93 & ~shift_1;
assign w638 = ~w636 & ~w637;
assign w639 = ~shift_0 & ~w638;
assign w640 = a_92 & ~shift_1;
assign w641 = a_90 & shift_1;
assign w642 = ~w640 & ~w641;
assign w643 = shift_0 & ~w642;
assign w644 = ~w639 & ~w643;
assign w645 = ~shift_3 & w644;
assign w646 = a_83 & shift_1;
assign w647 = a_85 & ~shift_1;
assign w648 = ~w646 & ~w647;
assign w649 = ~shift_0 & ~w648;
assign w650 = a_84 & ~shift_1;
assign w651 = a_82 & shift_1;
assign w652 = ~w650 & ~w651;
assign w653 = shift_0 & ~w652;
assign w654 = ~w649 & ~w653;
assign w655 = shift_3 & w654;
assign w656 = ~w645 & ~w655;
assign w657 = shift_2 & ~w656;
assign w658 = ~w635 & ~w657;
assign w659 = shift_5 & ~w658;
assign w660 = ~w613 & ~w659;
assign w661 = ~shift_4 & ~w660;
assign w662 = a_111 & shift_1;
assign w663 = a_113 & ~shift_1;
assign w664 = ~w662 & ~w663;
assign w665 = ~shift_0 & ~w664;
assign w666 = a_112 & ~shift_1;
assign w667 = a_110 & shift_1;
assign w668 = ~w666 & ~w667;
assign w669 = shift_0 & ~w668;
assign w670 = ~w665 & ~w669;
assign w671 = ~shift_3 & w670;
assign w672 = a_103 & shift_1;
assign w673 = a_105 & ~shift_1;
assign w674 = ~w672 & ~w673;
assign w675 = ~shift_0 & ~w674;
assign w676 = a_104 & ~shift_1;
assign w677 = a_102 & shift_1;
assign w678 = ~w676 & ~w677;
assign w679 = shift_0 & ~w678;
assign w680 = ~w675 & ~w679;
assign w681 = shift_3 & w680;
assign w682 = ~w671 & ~w681;
assign w683 = ~shift_2 & ~w682;
assign w684 = a_107 & shift_1;
assign w685 = a_109 & ~shift_1;
assign w686 = ~w684 & ~w685;
assign w687 = ~shift_0 & ~w686;
assign w688 = a_108 & ~shift_1;
assign w689 = a_106 & shift_1;
assign w690 = ~w688 & ~w689;
assign w691 = shift_0 & ~w690;
assign w692 = ~w687 & ~w691;
assign w693 = ~shift_3 & w692;
assign w694 = a_99 & shift_1;
assign w695 = a_101 & ~shift_1;
assign w696 = ~w694 & ~w695;
assign w697 = ~shift_0 & ~w696;
assign w698 = a_100 & ~shift_1;
assign w699 = a_98 & shift_1;
assign w700 = ~w698 & ~w699;
assign w701 = shift_0 & ~w700;
assign w702 = ~w697 & ~w701;
assign w703 = shift_3 & w702;
assign w704 = ~w693 & ~w703;
assign w705 = shift_2 & ~w704;
assign w706 = ~w683 & ~w705;
assign w707 = ~shift_5 & ~w706;
assign w708 = a_79 & shift_1;
assign w709 = a_81 & ~shift_1;
assign w710 = ~w708 & ~w709;
assign w711 = ~shift_0 & ~w710;
assign w712 = a_80 & ~shift_1;
assign w713 = a_78 & shift_1;
assign w714 = ~w712 & ~w713;
assign w715 = shift_0 & ~w714;
assign w716 = ~w711 & ~w715;
assign w717 = ~shift_3 & w716;
assign w718 = a_71 & shift_1;
assign w719 = a_73 & ~shift_1;
assign w720 = ~w718 & ~w719;
assign w721 = ~shift_0 & ~w720;
assign w722 = a_72 & ~shift_1;
assign w723 = a_70 & shift_1;
assign w724 = ~w722 & ~w723;
assign w725 = shift_0 & ~w724;
assign w726 = ~w721 & ~w725;
assign w727 = shift_3 & w726;
assign w728 = ~w717 & ~w727;
assign w729 = ~shift_2 & ~w728;
assign w730 = a_75 & shift_1;
assign w731 = a_77 & ~shift_1;
assign w732 = ~w730 & ~w731;
assign w733 = ~shift_0 & ~w732;
assign w734 = a_76 & ~shift_1;
assign w735 = a_74 & shift_1;
assign w736 = ~w734 & ~w735;
assign w737 = shift_0 & ~w736;
assign w738 = ~w733 & ~w737;
assign w739 = ~shift_3 & w738;
assign w740 = a_67 & shift_1;
assign w741 = a_69 & ~shift_1;
assign w742 = ~w740 & ~w741;
assign w743 = ~shift_0 & ~w742;
assign w744 = a_68 & ~shift_1;
assign w745 = a_66 & shift_1;
assign w746 = ~w744 & ~w745;
assign w747 = shift_0 & ~w746;
assign w748 = ~w743 & ~w747;
assign w749 = shift_3 & w748;
assign w750 = ~w739 & ~w749;
assign w751 = shift_2 & ~w750;
assign w752 = ~w729 & ~w751;
assign w753 = shift_5 & ~w752;
assign w754 = ~w707 & ~w753;
assign w755 = shift_4 & ~w754;
assign w756 = ~w661 & ~w755;
assign w757 = ~shift_6 & w756;
assign w758 = ~w567 & ~w757;
assign w759 = ~a_50 & ~shift_1;
assign w760 = ~a_48 & shift_1;
assign w761 = ~w759 & ~w760;
assign w762 = ~shift_0 & ~w761;
assign w763 = ~a_49 & ~shift_1;
assign w764 = ~a_47 & shift_1;
assign w765 = ~w763 & ~w764;
assign w766 = shift_0 & ~w765;
assign w767 = ~w762 & ~w766;
assign w768 = ~shift_3 & ~w767;
assign w769 = ~a_42 & ~shift_1;
assign w770 = ~a_40 & shift_1;
assign w771 = ~w769 & ~w770;
assign w772 = ~shift_0 & ~w771;
assign w773 = shift_0 & ~w393;
assign w774 = ~w772 & ~w773;
assign w775 = shift_3 & ~w774;
assign w776 = ~w768 & ~w775;
assign w777 = ~shift_2 & ~w776;
assign w778 = ~a_46 & ~shift_1;
assign w779 = ~a_44 & shift_1;
assign w780 = ~w778 & ~w779;
assign w781 = ~shift_0 & ~w780;
assign w782 = shift_0 & ~w415;
assign w783 = ~w781 & ~w782;
assign w784 = ~shift_3 & ~w783;
assign w785 = ~a_38 & ~shift_1;
assign w786 = ~a_36 & shift_1;
assign w787 = ~w785 & ~w786;
assign w788 = ~shift_0 & ~w787;
assign w789 = ~a_37 & ~shift_1;
assign w790 = ~a_35 & shift_1;
assign w791 = ~w789 & ~w790;
assign w792 = shift_0 & ~w791;
assign w793 = ~w788 & ~w792;
assign w794 = shift_3 & ~w793;
assign w795 = ~w784 & ~w794;
assign w796 = shift_2 & ~w795;
assign w797 = ~w777 & ~w796;
assign w798 = ~shift_5 & ~w797;
assign w799 = ~a_18 & ~shift_1;
assign w800 = ~a_16 & shift_1;
assign w801 = ~w799 & ~w800;
assign w802 = ~shift_0 & ~w801;
assign w803 = ~a_17 & ~shift_1;
assign w804 = ~a_15 & shift_1;
assign w805 = ~w803 & ~w804;
assign w806 = shift_0 & ~w805;
assign w807 = ~w802 & ~w806;
assign w808 = ~shift_3 & ~w807;
assign w809 = ~a_10 & ~shift_1;
assign w810 = ~a_8 & shift_1;
assign w811 = ~w809 & ~w810;
assign w812 = ~shift_0 & ~w811;
assign w813 = ~a_9 & ~shift_1;
assign w814 = ~a_7 & shift_1;
assign w815 = ~w813 & ~w814;
assign w816 = shift_0 & ~w815;
assign w817 = ~w812 & ~w816;
assign w818 = shift_3 & ~w817;
assign w819 = ~w808 & ~w818;
assign w820 = ~shift_2 & ~w819;
assign w821 = ~a_14 & ~shift_1;
assign w822 = ~a_12 & shift_1;
assign w823 = ~w821 & ~w822;
assign w824 = ~shift_0 & ~w823;
assign w825 = ~a_13 & ~shift_1;
assign w826 = ~a_11 & shift_1;
assign w827 = ~w825 & ~w826;
assign w828 = shift_0 & ~w827;
assign w829 = ~w824 & ~w828;
assign w830 = ~shift_3 & ~w829;
assign w831 = ~a_6 & ~shift_1;
assign w832 = ~a_4 & shift_1;
assign w833 = ~w831 & ~w832;
assign w834 = ~shift_0 & ~w833;
assign w835 = ~a_5 & ~shift_1;
assign w836 = ~a_3 & shift_1;
assign w837 = ~w835 & ~w836;
assign w838 = shift_0 & ~w837;
assign w839 = ~w834 & ~w838;
assign w840 = shift_3 & ~w839;
assign w841 = ~w830 & ~w840;
assign w842 = shift_2 & ~w841;
assign w843 = ~w820 & ~w842;
assign w844 = shift_5 & ~w843;
assign w845 = ~w798 & ~w844;
assign w846 = shift_4 & ~w845;
assign w847 = ~a_66 & ~shift_1;
assign w848 = ~a_64 & shift_1;
assign w849 = ~w847 & ~w848;
assign w850 = ~shift_0 & ~w849;
assign w851 = ~a_65 & ~shift_1;
assign w852 = ~a_63 & shift_1;
assign w853 = ~w851 & ~w852;
assign w854 = shift_0 & ~w853;
assign w855 = ~w850 & ~w854;
assign w856 = ~shift_3 & ~w855;
assign w857 = ~a_58 & ~shift_1;
assign w858 = ~a_56 & shift_1;
assign w859 = ~w857 & ~w858;
assign w860 = ~shift_0 & ~w859;
assign w861 = ~a_57 & ~shift_1;
assign w862 = ~a_55 & shift_1;
assign w863 = ~w861 & ~w862;
assign w864 = shift_0 & ~w863;
assign w865 = ~w860 & ~w864;
assign w866 = shift_3 & ~w865;
assign w867 = ~w856 & ~w866;
assign w868 = ~shift_2 & ~w867;
assign w869 = ~a_62 & ~shift_1;
assign w870 = ~a_60 & shift_1;
assign w871 = ~w869 & ~w870;
assign w872 = ~shift_0 & ~w871;
assign w873 = ~a_61 & ~shift_1;
assign w874 = ~a_59 & shift_1;
assign w875 = ~w873 & ~w874;
assign w876 = shift_0 & ~w875;
assign w877 = ~w872 & ~w876;
assign w878 = ~shift_3 & ~w877;
assign w879 = ~a_54 & ~shift_1;
assign w880 = ~a_52 & shift_1;
assign w881 = ~w879 & ~w880;
assign w882 = ~shift_0 & ~w881;
assign w883 = ~a_53 & ~shift_1;
assign w884 = ~a_51 & shift_1;
assign w885 = ~w883 & ~w884;
assign w886 = shift_0 & ~w885;
assign w887 = ~w882 & ~w886;
assign w888 = shift_3 & ~w887;
assign w889 = ~w878 & ~w888;
assign w890 = shift_2 & ~w889;
assign w891 = ~w868 & ~w890;
assign w892 = ~shift_5 & ~w891;
assign w893 = ~a_34 & ~shift_1;
assign w894 = ~a_32 & shift_1;
assign w895 = ~w893 & ~w894;
assign w896 = ~shift_0 & ~w895;
assign w897 = ~a_33 & ~shift_1;
assign w898 = ~a_31 & shift_1;
assign w899 = ~w897 & ~w898;
assign w900 = shift_0 & ~w899;
assign w901 = ~w896 & ~w900;
assign w902 = ~shift_3 & ~w901;
assign w903 = ~a_26 & ~shift_1;
assign w904 = ~a_24 & shift_1;
assign w905 = ~w903 & ~w904;
assign w906 = ~shift_0 & ~w905;
assign w907 = ~a_25 & ~shift_1;
assign w908 = ~a_23 & shift_1;
assign w909 = ~w907 & ~w908;
assign w910 = shift_0 & ~w909;
assign w911 = ~w906 & ~w910;
assign w912 = shift_3 & ~w911;
assign w913 = ~w902 & ~w912;
assign w914 = ~shift_2 & ~w913;
assign w915 = ~a_30 & ~shift_1;
assign w916 = ~a_28 & shift_1;
assign w917 = ~w915 & ~w916;
assign w918 = ~shift_0 & ~w917;
assign w919 = ~a_29 & ~shift_1;
assign w920 = ~a_27 & shift_1;
assign w921 = ~w919 & ~w920;
assign w922 = shift_0 & ~w921;
assign w923 = ~w918 & ~w922;
assign w924 = ~shift_3 & ~w923;
assign w925 = ~a_22 & ~shift_1;
assign w926 = ~a_20 & shift_1;
assign w927 = ~w925 & ~w926;
assign w928 = ~shift_0 & ~w927;
assign w929 = ~a_21 & ~shift_1;
assign w930 = ~a_19 & shift_1;
assign w931 = ~w929 & ~w930;
assign w932 = shift_0 & ~w931;
assign w933 = ~w928 & ~w932;
assign w934 = shift_3 & ~w933;
assign w935 = ~w924 & ~w934;
assign w936 = shift_2 & ~w935;
assign w937 = ~w914 & ~w936;
assign w938 = shift_5 & ~w937;
assign w939 = ~w892 & ~w938;
assign w940 = ~shift_4 & ~w939;
assign w941 = ~w846 & ~w940;
assign w942 = shift_6 & w941;
assign w943 = ~a_2 & ~shift_1;
assign w944 = ~a_0 & shift_1;
assign w945 = ~w943 & ~w944;
assign w946 = ~shift_0 & ~w945;
assign w947 = ~a_1 & ~shift_1;
assign w948 = ~a_127 & shift_1;
assign w949 = ~w947 & ~w948;
assign w950 = shift_0 & ~w949;
assign w951 = ~w946 & ~w950;
assign w952 = ~shift_3 & ~w951;
assign w953 = ~a_122 & ~shift_1;
assign w954 = ~a_120 & shift_1;
assign w955 = ~w953 & ~w954;
assign w956 = ~shift_0 & ~w955;
assign w957 = ~a_121 & ~shift_1;
assign w958 = ~a_119 & shift_1;
assign w959 = ~w957 & ~w958;
assign w960 = shift_0 & ~w959;
assign w961 = ~w956 & ~w960;
assign w962 = shift_3 & ~w961;
assign w963 = ~w952 & ~w962;
assign w964 = ~shift_2 & ~w963;
assign w965 = ~a_126 & ~shift_1;
assign w966 = ~a_124 & shift_1;
assign w967 = ~w965 & ~w966;
assign w968 = ~shift_0 & ~w967;
assign w969 = ~a_125 & ~shift_1;
assign w970 = ~a_123 & shift_1;
assign w971 = ~w969 & ~w970;
assign w972 = shift_0 & ~w971;
assign w973 = ~w968 & ~w972;
assign w974 = ~shift_3 & ~w973;
assign w975 = ~a_118 & ~shift_1;
assign w976 = ~a_116 & shift_1;
assign w977 = ~w975 & ~w976;
assign w978 = ~shift_0 & ~w977;
assign w979 = ~a_117 & ~shift_1;
assign w980 = ~a_115 & shift_1;
assign w981 = ~w979 & ~w980;
assign w982 = shift_0 & ~w981;
assign w983 = ~w978 & ~w982;
assign w984 = shift_3 & ~w983;
assign w985 = ~w974 & ~w984;
assign w986 = shift_2 & ~w985;
assign w987 = ~w964 & ~w986;
assign w988 = ~shift_5 & ~w987;
assign w989 = ~a_98 & ~shift_1;
assign w990 = ~a_96 & shift_1;
assign w991 = ~w989 & ~w990;
assign w992 = ~shift_0 & ~w991;
assign w993 = ~a_97 & ~shift_1;
assign w994 = ~a_95 & shift_1;
assign w995 = ~w993 & ~w994;
assign w996 = shift_0 & ~w995;
assign w997 = ~w992 & ~w996;
assign w998 = ~shift_3 & ~w997;
assign w999 = ~a_90 & ~shift_1;
assign w1000 = ~a_88 & shift_1;
assign w1001 = ~w999 & ~w1000;
assign w1002 = ~shift_0 & ~w1001;
assign w1003 = ~a_89 & ~shift_1;
assign w1004 = ~a_87 & shift_1;
assign w1005 = ~w1003 & ~w1004;
assign w1006 = shift_0 & ~w1005;
assign w1007 = ~w1002 & ~w1006;
assign w1008 = shift_3 & ~w1007;
assign w1009 = ~w998 & ~w1008;
assign w1010 = ~shift_2 & ~w1009;
assign w1011 = ~a_94 & ~shift_1;
assign w1012 = ~a_92 & shift_1;
assign w1013 = ~w1011 & ~w1012;
assign w1014 = ~shift_0 & ~w1013;
assign w1015 = ~a_93 & ~shift_1;
assign w1016 = ~a_91 & shift_1;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = shift_0 & ~w1017;
assign w1019 = ~w1014 & ~w1018;
assign w1020 = ~shift_3 & ~w1019;
assign w1021 = ~a_86 & ~shift_1;
assign w1022 = ~a_84 & shift_1;
assign w1023 = ~w1021 & ~w1022;
assign w1024 = ~shift_0 & ~w1023;
assign w1025 = ~a_85 & ~shift_1;
assign w1026 = ~a_83 & shift_1;
assign w1027 = ~w1025 & ~w1026;
assign w1028 = shift_0 & ~w1027;
assign w1029 = ~w1024 & ~w1028;
assign w1030 = shift_3 & ~w1029;
assign w1031 = ~w1020 & ~w1030;
assign w1032 = shift_2 & ~w1031;
assign w1033 = ~w1010 & ~w1032;
assign w1034 = shift_5 & ~w1033;
assign w1035 = ~w988 & ~w1034;
assign w1036 = ~shift_4 & ~w1035;
assign w1037 = ~a_114 & ~shift_1;
assign w1038 = ~a_112 & shift_1;
assign w1039 = ~w1037 & ~w1038;
assign w1040 = ~shift_0 & ~w1039;
assign w1041 = ~a_113 & ~shift_1;
assign w1042 = ~a_111 & shift_1;
assign w1043 = ~w1041 & ~w1042;
assign w1044 = shift_0 & ~w1043;
assign w1045 = ~w1040 & ~w1044;
assign w1046 = ~shift_3 & ~w1045;
assign w1047 = ~a_106 & ~shift_1;
assign w1048 = ~a_104 & shift_1;
assign w1049 = ~w1047 & ~w1048;
assign w1050 = ~shift_0 & ~w1049;
assign w1051 = ~a_105 & ~shift_1;
assign w1052 = ~a_103 & shift_1;
assign w1053 = ~w1051 & ~w1052;
assign w1054 = shift_0 & ~w1053;
assign w1055 = ~w1050 & ~w1054;
assign w1056 = shift_3 & ~w1055;
assign w1057 = ~w1046 & ~w1056;
assign w1058 = ~shift_2 & ~w1057;
assign w1059 = ~a_110 & ~shift_1;
assign w1060 = ~a_108 & shift_1;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = ~shift_0 & ~w1061;
assign w1063 = ~a_109 & ~shift_1;
assign w1064 = ~a_107 & shift_1;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = shift_0 & ~w1065;
assign w1067 = ~w1062 & ~w1066;
assign w1068 = ~shift_3 & ~w1067;
assign w1069 = ~a_102 & ~shift_1;
assign w1070 = ~a_100 & shift_1;
assign w1071 = ~w1069 & ~w1070;
assign w1072 = ~shift_0 & ~w1071;
assign w1073 = ~a_101 & ~shift_1;
assign w1074 = ~a_99 & shift_1;
assign w1075 = ~w1073 & ~w1074;
assign w1076 = shift_0 & ~w1075;
assign w1077 = ~w1072 & ~w1076;
assign w1078 = shift_3 & ~w1077;
assign w1079 = ~w1068 & ~w1078;
assign w1080 = shift_2 & ~w1079;
assign w1081 = ~w1058 & ~w1080;
assign w1082 = ~shift_5 & ~w1081;
assign w1083 = ~a_82 & ~shift_1;
assign w1084 = ~a_80 & shift_1;
assign w1085 = ~w1083 & ~w1084;
assign w1086 = ~shift_0 & ~w1085;
assign w1087 = ~a_81 & ~shift_1;
assign w1088 = ~a_79 & shift_1;
assign w1089 = ~w1087 & ~w1088;
assign w1090 = shift_0 & ~w1089;
assign w1091 = ~w1086 & ~w1090;
assign w1092 = ~shift_3 & ~w1091;
assign w1093 = ~a_74 & ~shift_1;
assign w1094 = ~a_72 & shift_1;
assign w1095 = ~w1093 & ~w1094;
assign w1096 = ~shift_0 & ~w1095;
assign w1097 = ~a_73 & ~shift_1;
assign w1098 = ~a_71 & shift_1;
assign w1099 = ~w1097 & ~w1098;
assign w1100 = shift_0 & ~w1099;
assign w1101 = ~w1096 & ~w1100;
assign w1102 = shift_3 & ~w1101;
assign w1103 = ~w1092 & ~w1102;
assign w1104 = ~shift_2 & ~w1103;
assign w1105 = ~a_78 & ~shift_1;
assign w1106 = ~a_76 & shift_1;
assign w1107 = ~w1105 & ~w1106;
assign w1108 = ~shift_0 & ~w1107;
assign w1109 = ~a_77 & ~shift_1;
assign w1110 = ~a_75 & shift_1;
assign w1111 = ~w1109 & ~w1110;
assign w1112 = shift_0 & ~w1111;
assign w1113 = ~w1108 & ~w1112;
assign w1114 = ~shift_3 & ~w1113;
assign w1115 = ~a_70 & ~shift_1;
assign w1116 = ~a_68 & shift_1;
assign w1117 = ~w1115 & ~w1116;
assign w1118 = ~shift_0 & ~w1117;
assign w1119 = ~a_69 & ~shift_1;
assign w1120 = ~a_67 & shift_1;
assign w1121 = ~w1119 & ~w1120;
assign w1122 = shift_0 & ~w1121;
assign w1123 = ~w1118 & ~w1122;
assign w1124 = shift_3 & ~w1123;
assign w1125 = ~w1114 & ~w1124;
assign w1126 = shift_2 & ~w1125;
assign w1127 = ~w1104 & ~w1126;
assign w1128 = shift_5 & ~w1127;
assign w1129 = ~w1082 & ~w1128;
assign w1130 = shift_4 & ~w1129;
assign w1131 = ~w1036 & ~w1130;
assign w1132 = ~shift_6 & w1131;
assign w1133 = ~w942 & ~w1132;
assign w1134 = a_65 & shift_1;
assign w1135 = a_67 & ~shift_1;
assign w1136 = ~w1134 & ~w1135;
assign w1137 = ~shift_0 & ~w1136;
assign w1138 = a_66 & ~shift_1;
assign w1139 = a_64 & shift_1;
assign w1140 = ~w1138 & ~w1139;
assign w1141 = shift_0 & ~w1140;
assign w1142 = ~w1137 & ~w1141;
assign w1143 = ~shift_3 & w1142;
assign w1144 = a_57 & shift_1;
assign w1145 = a_59 & ~shift_1;
assign w1146 = ~w1144 & ~w1145;
assign w1147 = ~shift_0 & ~w1146;
assign w1148 = a_58 & ~shift_1;
assign w1149 = a_56 & shift_1;
assign w1150 = ~w1148 & ~w1149;
assign w1151 = shift_0 & ~w1150;
assign w1152 = ~w1147 & ~w1151;
assign w1153 = shift_3 & w1152;
assign w1154 = ~w1143 & ~w1153;
assign w1155 = ~shift_2 & ~w1154;
assign w1156 = a_61 & shift_1;
assign w1157 = a_63 & ~shift_1;
assign w1158 = ~w1156 & ~w1157;
assign w1159 = ~shift_0 & ~w1158;
assign w1160 = a_62 & ~shift_1;
assign w1161 = a_60 & shift_1;
assign w1162 = ~w1160 & ~w1161;
assign w1163 = shift_0 & ~w1162;
assign w1164 = ~w1159 & ~w1163;
assign w1165 = ~shift_3 & w1164;
assign w1166 = a_53 & shift_1;
assign w1167 = a_55 & ~shift_1;
assign w1168 = ~w1166 & ~w1167;
assign w1169 = ~shift_0 & ~w1168;
assign w1170 = a_54 & ~shift_1;
assign w1171 = a_52 & shift_1;
assign w1172 = ~w1170 & ~w1171;
assign w1173 = shift_0 & ~w1172;
assign w1174 = ~w1169 & ~w1173;
assign w1175 = shift_3 & w1174;
assign w1176 = ~w1165 & ~w1175;
assign w1177 = shift_2 & ~w1176;
assign w1178 = ~w1155 & ~w1177;
assign w1179 = ~shift_5 & ~w1178;
assign w1180 = a_33 & shift_1;
assign w1181 = a_35 & ~shift_1;
assign w1182 = ~w1180 & ~w1181;
assign w1183 = ~shift_0 & ~w1182;
assign w1184 = a_34 & ~shift_1;
assign w1185 = a_32 & shift_1;
assign w1186 = ~w1184 & ~w1185;
assign w1187 = shift_0 & ~w1186;
assign w1188 = ~w1183 & ~w1187;
assign w1189 = ~shift_3 & w1188;
assign w1190 = a_25 & shift_1;
assign w1191 = a_27 & ~shift_1;
assign w1192 = ~w1190 & ~w1191;
assign w1193 = ~shift_0 & ~w1192;
assign w1194 = a_26 & ~shift_1;
assign w1195 = a_24 & shift_1;
assign w1196 = ~w1194 & ~w1195;
assign w1197 = shift_0 & ~w1196;
assign w1198 = ~w1193 & ~w1197;
assign w1199 = shift_3 & w1198;
assign w1200 = ~w1189 & ~w1199;
assign w1201 = ~shift_2 & ~w1200;
assign w1202 = a_29 & shift_1;
assign w1203 = a_31 & ~shift_1;
assign w1204 = ~w1202 & ~w1203;
assign w1205 = ~shift_0 & ~w1204;
assign w1206 = a_30 & ~shift_1;
assign w1207 = a_28 & shift_1;
assign w1208 = ~w1206 & ~w1207;
assign w1209 = shift_0 & ~w1208;
assign w1210 = ~w1205 & ~w1209;
assign w1211 = ~shift_3 & w1210;
assign w1212 = a_21 & shift_1;
assign w1213 = a_23 & ~shift_1;
assign w1214 = ~w1212 & ~w1213;
assign w1215 = ~shift_0 & ~w1214;
assign w1216 = a_22 & ~shift_1;
assign w1217 = a_20 & shift_1;
assign w1218 = ~w1216 & ~w1217;
assign w1219 = shift_0 & ~w1218;
assign w1220 = ~w1215 & ~w1219;
assign w1221 = shift_3 & w1220;
assign w1222 = ~w1211 & ~w1221;
assign w1223 = shift_2 & ~w1222;
assign w1224 = ~w1201 & ~w1223;
assign w1225 = shift_5 & ~w1224;
assign w1226 = ~w1179 & ~w1225;
assign w1227 = ~shift_4 & ~w1226;
assign w1228 = ~shift_0 & ~w100;
assign w1229 = a_38 & ~shift_1;
assign w1230 = a_36 & shift_1;
assign w1231 = ~w1229 & ~w1230;
assign w1232 = shift_0 & ~w1231;
assign w1233 = ~w1228 & ~w1232;
assign w1234 = shift_3 & w1233;
assign w1235 = ~shift_0 & ~w110;
assign w1236 = shift_0 & ~w780;
assign w1237 = ~w1235 & ~w1236;
assign w1238 = ~shift_3 & ~w1237;
assign w1239 = ~w1234 & ~w1238;
assign w1240 = shift_2 & ~w1239;
assign w1241 = a_49 & shift_1;
assign w1242 = a_51 & ~shift_1;
assign w1243 = ~w1241 & ~w1242;
assign w1244 = ~shift_0 & ~w1243;
assign w1245 = a_50 & ~shift_1;
assign w1246 = a_48 & shift_1;
assign w1247 = ~w1245 & ~w1246;
assign w1248 = shift_0 & ~w1247;
assign w1249 = ~w1244 & ~w1248;
assign w1250 = ~shift_3 & w1249;
assign w1251 = a_41 & shift_1;
assign w1252 = a_43 & ~shift_1;
assign w1253 = ~w1251 & ~w1252;
assign w1254 = ~shift_0 & ~w1253;
assign w1255 = a_42 & ~shift_1;
assign w1256 = a_40 & shift_1;
assign w1257 = ~w1255 & ~w1256;
assign w1258 = shift_0 & ~w1257;
assign w1259 = ~w1254 & ~w1258;
assign w1260 = shift_3 & w1259;
assign w1261 = ~w1250 & ~w1260;
assign w1262 = ~shift_2 & ~w1261;
assign w1263 = ~w1240 & ~w1262;
assign w1264 = ~shift_5 & ~w1263;
assign w1265 = a_17 & shift_1;
assign w1266 = a_19 & ~shift_1;
assign w1267 = ~w1265 & ~w1266;
assign w1268 = ~shift_0 & ~w1267;
assign w1269 = a_18 & ~shift_1;
assign w1270 = a_16 & shift_1;
assign w1271 = ~w1269 & ~w1270;
assign w1272 = shift_0 & ~w1271;
assign w1273 = ~w1268 & ~w1272;
assign w1274 = ~shift_3 & w1273;
assign w1275 = a_9 & shift_1;
assign w1276 = a_11 & ~shift_1;
assign w1277 = ~w1275 & ~w1276;
assign w1278 = ~shift_0 & ~w1277;
assign w1279 = a_10 & ~shift_1;
assign w1280 = a_8 & shift_1;
assign w1281 = ~w1279 & ~w1280;
assign w1282 = shift_0 & ~w1281;
assign w1283 = ~w1278 & ~w1282;
assign w1284 = shift_3 & w1283;
assign w1285 = ~w1274 & ~w1284;
assign w1286 = ~shift_2 & ~w1285;
assign w1287 = a_13 & shift_1;
assign w1288 = a_15 & ~shift_1;
assign w1289 = ~w1287 & ~w1288;
assign w1290 = ~shift_0 & ~w1289;
assign w1291 = a_14 & ~shift_1;
assign w1292 = a_12 & shift_1;
assign w1293 = ~w1291 & ~w1292;
assign w1294 = shift_0 & ~w1293;
assign w1295 = ~w1290 & ~w1294;
assign w1296 = ~shift_3 & w1295;
assign w1297 = a_5 & shift_1;
assign w1298 = a_7 & ~shift_1;
assign w1299 = ~w1297 & ~w1298;
assign w1300 = ~shift_0 & ~w1299;
assign w1301 = a_6 & ~shift_1;
assign w1302 = a_4 & shift_1;
assign w1303 = ~w1301 & ~w1302;
assign w1304 = shift_0 & ~w1303;
assign w1305 = ~w1300 & ~w1304;
assign w1306 = shift_3 & w1305;
assign w1307 = ~w1296 & ~w1306;
assign w1308 = shift_2 & ~w1307;
assign w1309 = ~w1286 & ~w1308;
assign w1310 = shift_5 & ~w1309;
assign w1311 = ~w1264 & ~w1310;
assign w1312 = shift_4 & ~w1311;
assign w1313 = ~w1227 & ~w1312;
assign w1314 = shift_6 & w1313;
assign w1315 = a_113 & shift_1;
assign w1316 = a_115 & ~shift_1;
assign w1317 = ~w1315 & ~w1316;
assign w1318 = ~shift_0 & ~w1317;
assign w1319 = a_114 & ~shift_1;
assign w1320 = a_112 & shift_1;
assign w1321 = ~w1319 & ~w1320;
assign w1322 = shift_0 & ~w1321;
assign w1323 = ~w1318 & ~w1322;
assign w1324 = ~shift_3 & w1323;
assign w1325 = a_105 & shift_1;
assign w1326 = a_107 & ~shift_1;
assign w1327 = ~w1325 & ~w1326;
assign w1328 = ~shift_0 & ~w1327;
assign w1329 = a_106 & ~shift_1;
assign w1330 = a_104 & shift_1;
assign w1331 = ~w1329 & ~w1330;
assign w1332 = shift_0 & ~w1331;
assign w1333 = ~w1328 & ~w1332;
assign w1334 = shift_3 & w1333;
assign w1335 = ~w1324 & ~w1334;
assign w1336 = ~shift_2 & ~w1335;
assign w1337 = a_109 & shift_1;
assign w1338 = a_111 & ~shift_1;
assign w1339 = ~w1337 & ~w1338;
assign w1340 = ~shift_0 & ~w1339;
assign w1341 = a_110 & ~shift_1;
assign w1342 = a_108 & shift_1;
assign w1343 = ~w1341 & ~w1342;
assign w1344 = shift_0 & ~w1343;
assign w1345 = ~w1340 & ~w1344;
assign w1346 = ~shift_3 & w1345;
assign w1347 = a_101 & shift_1;
assign w1348 = a_103 & ~shift_1;
assign w1349 = ~w1347 & ~w1348;
assign w1350 = ~shift_0 & ~w1349;
assign w1351 = a_102 & ~shift_1;
assign w1352 = a_100 & shift_1;
assign w1353 = ~w1351 & ~w1352;
assign w1354 = shift_0 & ~w1353;
assign w1355 = ~w1350 & ~w1354;
assign w1356 = shift_3 & w1355;
assign w1357 = ~w1346 & ~w1356;
assign w1358 = shift_2 & ~w1357;
assign w1359 = ~w1336 & ~w1358;
assign w1360 = ~shift_5 & ~w1359;
assign w1361 = a_81 & shift_1;
assign w1362 = a_83 & ~shift_1;
assign w1363 = ~w1361 & ~w1362;
assign w1364 = ~shift_0 & ~w1363;
assign w1365 = a_82 & ~shift_1;
assign w1366 = a_80 & shift_1;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = shift_0 & ~w1367;
assign w1369 = ~w1364 & ~w1368;
assign w1370 = ~shift_3 & w1369;
assign w1371 = a_73 & shift_1;
assign w1372 = a_75 & ~shift_1;
assign w1373 = ~w1371 & ~w1372;
assign w1374 = ~shift_0 & ~w1373;
assign w1375 = a_74 & ~shift_1;
assign w1376 = a_72 & shift_1;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = shift_0 & ~w1377;
assign w1379 = ~w1374 & ~w1378;
assign w1380 = shift_3 & w1379;
assign w1381 = ~w1370 & ~w1380;
assign w1382 = ~shift_2 & ~w1381;
assign w1383 = a_77 & shift_1;
assign w1384 = a_79 & ~shift_1;
assign w1385 = ~w1383 & ~w1384;
assign w1386 = ~shift_0 & ~w1385;
assign w1387 = a_78 & ~shift_1;
assign w1388 = a_76 & shift_1;
assign w1389 = ~w1387 & ~w1388;
assign w1390 = shift_0 & ~w1389;
assign w1391 = ~w1386 & ~w1390;
assign w1392 = ~shift_3 & w1391;
assign w1393 = a_69 & shift_1;
assign w1394 = a_71 & ~shift_1;
assign w1395 = ~w1393 & ~w1394;
assign w1396 = ~shift_0 & ~w1395;
assign w1397 = a_70 & ~shift_1;
assign w1398 = a_68 & shift_1;
assign w1399 = ~w1397 & ~w1398;
assign w1400 = shift_0 & ~w1399;
assign w1401 = ~w1396 & ~w1400;
assign w1402 = shift_3 & w1401;
assign w1403 = ~w1392 & ~w1402;
assign w1404 = shift_2 & ~w1403;
assign w1405 = ~w1382 & ~w1404;
assign w1406 = shift_5 & ~w1405;
assign w1407 = ~w1360 & ~w1406;
assign w1408 = shift_4 & ~w1407;
assign w1409 = a_1 & shift_1;
assign w1410 = a_3 & ~shift_1;
assign w1411 = ~w1409 & ~w1410;
assign w1412 = ~shift_0 & ~w1411;
assign w1413 = a_2 & ~shift_1;
assign w1414 = a_0 & shift_1;
assign w1415 = ~w1413 & ~w1414;
assign w1416 = shift_0 & ~w1415;
assign w1417 = ~w1412 & ~w1416;
assign w1418 = ~shift_3 & w1417;
assign w1419 = a_121 & shift_1;
assign w1420 = a_123 & ~shift_1;
assign w1421 = ~w1419 & ~w1420;
assign w1422 = ~shift_0 & ~w1421;
assign w1423 = a_122 & ~shift_1;
assign w1424 = a_120 & shift_1;
assign w1425 = ~w1423 & ~w1424;
assign w1426 = shift_0 & ~w1425;
assign w1427 = ~w1422 & ~w1426;
assign w1428 = shift_3 & w1427;
assign w1429 = ~w1418 & ~w1428;
assign w1430 = ~shift_2 & ~w1429;
assign w1431 = a_125 & shift_1;
assign w1432 = a_127 & ~shift_1;
assign w1433 = ~w1431 & ~w1432;
assign w1434 = ~shift_0 & ~w1433;
assign w1435 = a_126 & ~shift_1;
assign w1436 = a_124 & shift_1;
assign w1437 = ~w1435 & ~w1436;
assign w1438 = shift_0 & ~w1437;
assign w1439 = ~w1434 & ~w1438;
assign w1440 = ~shift_3 & w1439;
assign w1441 = a_117 & shift_1;
assign w1442 = a_119 & ~shift_1;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = ~shift_0 & ~w1443;
assign w1445 = a_118 & ~shift_1;
assign w1446 = a_116 & shift_1;
assign w1447 = ~w1445 & ~w1446;
assign w1448 = shift_0 & ~w1447;
assign w1449 = ~w1444 & ~w1448;
assign w1450 = shift_3 & w1449;
assign w1451 = ~w1440 & ~w1450;
assign w1452 = shift_2 & ~w1451;
assign w1453 = ~w1430 & ~w1452;
assign w1454 = ~shift_5 & ~w1453;
assign w1455 = a_97 & shift_1;
assign w1456 = a_99 & ~shift_1;
assign w1457 = ~w1455 & ~w1456;
assign w1458 = ~shift_0 & ~w1457;
assign w1459 = a_98 & ~shift_1;
assign w1460 = a_96 & shift_1;
assign w1461 = ~w1459 & ~w1460;
assign w1462 = shift_0 & ~w1461;
assign w1463 = ~w1458 & ~w1462;
assign w1464 = ~shift_3 & w1463;
assign w1465 = a_89 & shift_1;
assign w1466 = a_91 & ~shift_1;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = ~shift_0 & ~w1467;
assign w1469 = a_90 & ~shift_1;
assign w1470 = a_88 & shift_1;
assign w1471 = ~w1469 & ~w1470;
assign w1472 = shift_0 & ~w1471;
assign w1473 = ~w1468 & ~w1472;
assign w1474 = shift_3 & w1473;
assign w1475 = ~w1464 & ~w1474;
assign w1476 = ~shift_2 & ~w1475;
assign w1477 = a_93 & shift_1;
assign w1478 = a_95 & ~shift_1;
assign w1479 = ~w1477 & ~w1478;
assign w1480 = ~shift_0 & ~w1479;
assign w1481 = a_94 & ~shift_1;
assign w1482 = a_92 & shift_1;
assign w1483 = ~w1481 & ~w1482;
assign w1484 = shift_0 & ~w1483;
assign w1485 = ~w1480 & ~w1484;
assign w1486 = ~shift_3 & w1485;
assign w1487 = a_85 & shift_1;
assign w1488 = a_87 & ~shift_1;
assign w1489 = ~w1487 & ~w1488;
assign w1490 = ~shift_0 & ~w1489;
assign w1491 = a_86 & ~shift_1;
assign w1492 = a_84 & shift_1;
assign w1493 = ~w1491 & ~w1492;
assign w1494 = shift_0 & ~w1493;
assign w1495 = ~w1490 & ~w1494;
assign w1496 = shift_3 & w1495;
assign w1497 = ~w1486 & ~w1496;
assign w1498 = shift_2 & ~w1497;
assign w1499 = ~w1476 & ~w1498;
assign w1500 = shift_5 & ~w1499;
assign w1501 = ~w1454 & ~w1500;
assign w1502 = ~shift_4 & ~w1501;
assign w1503 = ~w1408 & ~w1502;
assign w1504 = ~shift_6 & w1503;
assign w1505 = ~w1314 & ~w1504;
assign w1506 = shift_2 & ~w20;
assign w1507 = shift_3 & ~w30;
assign w1508 = ~shift_3 & ~w370;
assign w1509 = ~w1507 & ~w1508;
assign w1510 = ~shift_2 & ~w1509;
assign w1511 = ~w1506 & ~w1510;
assign w1512 = ~shift_5 & ~w1511;
assign w1513 = shift_2 & ~w66;
assign w1514 = shift_3 & ~w76;
assign w1515 = ~shift_3 & ~w134;
assign w1516 = ~w1514 & ~w1515;
assign w1517 = ~shift_2 & ~w1516;
assign w1518 = ~w1513 & ~w1517;
assign w1519 = shift_5 & ~w1518;
assign w1520 = ~w1512 & ~w1519;
assign w1521 = ~shift_4 & ~w1520;
assign w1522 = ~shift_3 & ~w40;
assign w1523 = shift_3 & ~w124;
assign w1524 = ~w1522 & ~w1523;
assign w1525 = ~shift_2 & ~w1524;
assign w1526 = shift_2 & ~w114;
assign w1527 = ~w1525 & ~w1526;
assign w1528 = ~shift_5 & ~w1527;
assign w1529 = shift_2 & ~w160;
assign w1530 = shift_3 & ~w170;
assign w1531 = ~shift_3 & ~w86;
assign w1532 = ~w1530 & ~w1531;
assign w1533 = ~shift_2 & ~w1532;
assign w1534 = ~w1529 & ~w1533;
assign w1535 = shift_5 & ~w1534;
assign w1536 = ~w1528 & ~w1535;
assign w1537 = shift_4 & ~w1536;
assign w1538 = ~w1521 & ~w1537;
assign w1539 = shift_6 & w1538;
assign w1540 = shift_2 & ~w210;
assign w1541 = ~shift_3 & ~w180;
assign w1542 = shift_3 & ~w220;
assign w1543 = ~w1541 & ~w1542;
assign w1544 = ~shift_2 & ~w1543;
assign w1545 = ~w1540 & ~w1544;
assign w1546 = ~shift_5 & ~w1545;
assign w1547 = shift_2 & ~w256;
assign w1548 = shift_3 & ~w266;
assign w1549 = ~shift_3 & ~w324;
assign w1550 = ~w1548 & ~w1549;
assign w1551 = ~shift_2 & ~w1550;
assign w1552 = ~w1547 & ~w1551;
assign w1553 = shift_5 & ~w1552;
assign w1554 = ~w1546 & ~w1553;
assign w1555 = ~shift_4 & ~w1554;
assign w1556 = shift_2 & ~w304;
assign w1557 = ~shift_3 & ~w230;
assign w1558 = shift_3 & ~w314;
assign w1559 = ~w1557 & ~w1558;
assign w1560 = ~shift_2 & ~w1559;
assign w1561 = ~w1556 & ~w1560;
assign w1562 = ~shift_5 & ~w1561;
assign w1563 = shift_2 & ~w350;
assign w1564 = shift_3 & ~w360;
assign w1565 = ~shift_3 & ~w276;
assign w1566 = ~w1564 & ~w1565;
assign w1567 = ~shift_2 & ~w1566;
assign w1568 = ~w1563 & ~w1567;
assign w1569 = shift_5 & ~w1568;
assign w1570 = ~w1562 & ~w1569;
assign w1571 = shift_4 & ~w1570;
assign w1572 = ~w1555 & ~w1571;
assign w1573 = ~shift_6 & w1572;
assign w1574 = ~w1539 & ~w1573;
assign w1575 = shift_2 & ~w492;
assign w1576 = ~shift_3 & w748;
assign w1577 = shift_3 & w502;
assign w1578 = ~w1576 & ~w1577;
assign w1579 = ~shift_2 & ~w1578;
assign w1580 = ~w1575 & ~w1579;
assign w1581 = ~shift_5 & ~w1580;
assign w1582 = shift_2 & ~w538;
assign w1583 = ~shift_3 & w411;
assign w1584 = shift_3 & w548;
assign w1585 = ~w1583 & ~w1584;
assign w1586 = ~shift_2 & ~w1585;
assign w1587 = ~w1582 & ~w1586;
assign w1588 = shift_5 & ~w1587;
assign w1589 = ~w1581 & ~w1588;
assign w1590 = ~shift_4 & ~w1589;
assign w1591 = ~shift_3 & w512;
assign w1592 = shift_3 & ~w418;
assign w1593 = ~w1591 & ~w1592;
assign w1594 = ~shift_2 & ~w1593;
assign w1595 = shift_2 & ~w401;
assign w1596 = ~w1594 & ~w1595;
assign w1597 = ~shift_5 & ~w1596;
assign w1598 = shift_2 & ~w444;
assign w1599 = ~shift_3 & w558;
assign w1600 = shift_3 & w454;
assign w1601 = ~w1599 & ~w1600;
assign w1602 = ~shift_2 & ~w1601;
assign w1603 = ~w1598 & ~w1602;
assign w1604 = shift_5 & ~w1603;
assign w1605 = ~w1597 & ~w1604;
assign w1606 = shift_4 & ~w1605;
assign w1607 = ~w1590 & ~w1606;
assign w1608 = shift_6 & w1607;
assign w1609 = shift_2 & ~w588;
assign w1610 = ~shift_3 & w464;
assign w1611 = shift_3 & w598;
assign w1612 = ~w1610 & ~w1611;
assign w1613 = ~shift_2 & ~w1612;
assign w1614 = ~w1609 & ~w1613;
assign w1615 = ~shift_5 & ~w1614;
assign w1616 = shift_2 & ~w634;
assign w1617 = ~shift_3 & w702;
assign w1618 = shift_3 & w644;
assign w1619 = ~w1617 & ~w1618;
assign w1620 = ~shift_2 & ~w1619;
assign w1621 = ~w1616 & ~w1620;
assign w1622 = shift_5 & ~w1621;
assign w1623 = ~w1615 & ~w1622;
assign w1624 = ~shift_4 & ~w1623;
assign w1625 = shift_2 & ~w682;
assign w1626 = ~shift_3 & w608;
assign w1627 = shift_3 & w692;
assign w1628 = ~w1626 & ~w1627;
assign w1629 = ~shift_2 & ~w1628;
assign w1630 = ~w1625 & ~w1629;
assign w1631 = ~shift_5 & ~w1630;
assign w1632 = shift_2 & ~w728;
assign w1633 = ~shift_3 & w654;
assign w1634 = shift_3 & w738;
assign w1635 = ~w1633 & ~w1634;
assign w1636 = ~shift_2 & ~w1635;
assign w1637 = ~w1632 & ~w1636;
assign w1638 = shift_5 & ~w1637;
assign w1639 = ~w1631 & ~w1638;
assign w1640 = shift_4 & ~w1639;
assign w1641 = ~w1624 & ~w1640;
assign w1642 = ~shift_6 & w1641;
assign w1643 = ~w1608 & ~w1642;
assign w1644 = shift_2 & ~w867;
assign w1645 = shift_3 & ~w877;
assign w1646 = ~shift_3 & ~w1123;
assign w1647 = ~w1645 & ~w1646;
assign w1648 = ~shift_2 & ~w1647;
assign w1649 = ~w1644 & ~w1648;
assign w1650 = ~shift_5 & ~w1649;
assign w1651 = shift_2 & ~w913;
assign w1652 = ~shift_3 & ~w793;
assign w1653 = shift_3 & ~w923;
assign w1654 = ~w1652 & ~w1653;
assign w1655 = ~shift_2 & ~w1654;
assign w1656 = ~w1651 & ~w1655;
assign w1657 = shift_5 & ~w1656;
assign w1658 = ~w1650 & ~w1657;
assign w1659 = ~shift_4 & ~w1658;
assign w1660 = shift_2 & ~w776;
assign w1661 = ~shift_3 & ~w887;
assign w1662 = shift_3 & ~w783;
assign w1663 = ~w1661 & ~w1662;
assign w1664 = ~shift_2 & ~w1663;
assign w1665 = ~w1660 & ~w1664;
assign w1666 = ~shift_5 & ~w1665;
assign w1667 = shift_2 & ~w819;
assign w1668 = shift_3 & ~w829;
assign w1669 = ~shift_3 & ~w933;
assign w1670 = ~w1668 & ~w1669;
assign w1671 = ~shift_2 & ~w1670;
assign w1672 = ~w1667 & ~w1671;
assign w1673 = shift_5 & ~w1672;
assign w1674 = ~w1666 & ~w1673;
assign w1675 = shift_4 & ~w1674;
assign w1676 = ~w1659 & ~w1675;
assign w1677 = shift_6 & w1676;
assign w1678 = shift_2 & ~w963;
assign w1679 = ~shift_3 & ~w839;
assign w1680 = shift_3 & ~w973;
assign w1681 = ~w1679 & ~w1680;
assign w1682 = ~shift_2 & ~w1681;
assign w1683 = ~w1678 & ~w1682;
assign w1684 = ~shift_5 & ~w1683;
assign w1685 = shift_2 & ~w1009;
assign w1686 = shift_3 & ~w1019;
assign w1687 = ~shift_3 & ~w1077;
assign w1688 = ~w1686 & ~w1687;
assign w1689 = ~shift_2 & ~w1688;
assign w1690 = ~w1685 & ~w1689;
assign w1691 = shift_5 & ~w1690;
assign w1692 = ~w1684 & ~w1691;
assign w1693 = ~shift_4 & ~w1692;
assign w1694 = shift_2 & ~w1057;
assign w1695 = ~shift_3 & ~w983;
assign w1696 = shift_3 & ~w1067;
assign w1697 = ~w1695 & ~w1696;
assign w1698 = ~shift_2 & ~w1697;
assign w1699 = ~w1694 & ~w1698;
assign w1700 = ~shift_5 & ~w1699;
assign w1701 = shift_2 & ~w1103;
assign w1702 = shift_3 & ~w1113;
assign w1703 = ~shift_3 & ~w1029;
assign w1704 = ~w1702 & ~w1703;
assign w1705 = ~shift_2 & ~w1704;
assign w1706 = ~w1701 & ~w1705;
assign w1707 = shift_5 & ~w1706;
assign w1708 = ~w1700 & ~w1707;
assign w1709 = shift_4 & ~w1708;
assign w1710 = ~w1693 & ~w1709;
assign w1711 = ~shift_6 & w1710;
assign w1712 = ~w1677 & ~w1711;
assign w1713 = shift_2 & ~w1154;
assign w1714 = ~shift_3 & w1401;
assign w1715 = shift_3 & w1164;
assign w1716 = ~w1714 & ~w1715;
assign w1717 = ~shift_2 & ~w1716;
assign w1718 = ~w1713 & ~w1717;
assign w1719 = ~shift_5 & ~w1718;
assign w1720 = shift_2 & ~w1200;
assign w1721 = ~shift_3 & w1233;
assign w1722 = shift_3 & w1210;
assign w1723 = ~w1721 & ~w1722;
assign w1724 = ~shift_2 & ~w1723;
assign w1725 = ~w1720 & ~w1724;
assign w1726 = shift_5 & ~w1725;
assign w1727 = ~w1719 & ~w1726;
assign w1728 = ~shift_4 & ~w1727;
assign w1729 = ~shift_3 & w1174;
assign w1730 = shift_3 & ~w1237;
assign w1731 = ~w1729 & ~w1730;
assign w1732 = ~shift_2 & ~w1731;
assign w1733 = shift_2 & ~w1261;
assign w1734 = ~w1732 & ~w1733;
assign w1735 = ~shift_5 & ~w1734;
assign w1736 = shift_2 & ~w1285;
assign w1737 = ~shift_3 & w1220;
assign w1738 = shift_3 & w1295;
assign w1739 = ~w1737 & ~w1738;
assign w1740 = ~shift_2 & ~w1739;
assign w1741 = ~w1736 & ~w1740;
assign w1742 = shift_5 & ~w1741;
assign w1743 = ~w1735 & ~w1742;
assign w1744 = shift_4 & ~w1743;
assign w1745 = ~w1728 & ~w1744;
assign w1746 = shift_6 & w1745;
assign w1747 = shift_2 & ~w1429;
assign w1748 = ~shift_3 & w1305;
assign w1749 = shift_3 & w1439;
assign w1750 = ~w1748 & ~w1749;
assign w1751 = ~shift_2 & ~w1750;
assign w1752 = ~w1747 & ~w1751;
assign w1753 = ~shift_5 & ~w1752;
assign w1754 = shift_2 & ~w1475;
assign w1755 = ~shift_3 & w1355;
assign w1756 = shift_3 & w1485;
assign w1757 = ~w1755 & ~w1756;
assign w1758 = ~shift_2 & ~w1757;
assign w1759 = ~w1754 & ~w1758;
assign w1760 = shift_5 & ~w1759;
assign w1761 = ~w1753 & ~w1760;
assign w1762 = ~shift_4 & ~w1761;
assign w1763 = shift_2 & ~w1335;
assign w1764 = ~shift_3 & w1449;
assign w1765 = shift_3 & w1345;
assign w1766 = ~w1764 & ~w1765;
assign w1767 = ~shift_2 & ~w1766;
assign w1768 = ~w1763 & ~w1767;
assign w1769 = ~shift_5 & ~w1768;
assign w1770 = shift_2 & ~w1381;
assign w1771 = ~shift_3 & w1495;
assign w1772 = shift_3 & w1391;
assign w1773 = ~w1771 & ~w1772;
assign w1774 = ~shift_2 & ~w1773;
assign w1775 = ~w1770 & ~w1774;
assign w1776 = shift_5 & ~w1775;
assign w1777 = ~w1769 & ~w1776;
assign w1778 = shift_4 & ~w1777;
assign w1779 = ~w1762 & ~w1778;
assign w1780 = ~shift_6 & w1779;
assign w1781 = ~w1746 & ~w1780;
assign w1782 = ~shift_3 & ~w348;
assign w1783 = shift_3 & ~w8;
assign w1784 = ~w1782 & ~w1783;
assign w1785 = ~shift_2 & ~w1784;
assign w1786 = shift_2 & ~w1509;
assign w1787 = ~w1785 & ~w1786;
assign w1788 = ~shift_5 & ~w1787;
assign w1789 = ~shift_3 & w102;
assign w1790 = shift_3 & ~w54;
assign w1791 = ~w1789 & ~w1790;
assign w1792 = ~shift_2 & ~w1791;
assign w1793 = shift_2 & ~w1516;
assign w1794 = ~w1792 & ~w1793;
assign w1795 = shift_5 & ~w1794;
assign w1796 = ~w1788 & ~w1795;
assign w1797 = ~shift_4 & ~w1796;
assign w1798 = ~shift_3 & ~w18;
assign w1799 = shift_3 & ~w112;
assign w1800 = ~w1798 & ~w1799;
assign w1801 = ~shift_2 & ~w1800;
assign w1802 = shift_2 & ~w1524;
assign w1803 = ~w1801 & ~w1802;
assign w1804 = ~shift_5 & ~w1803;
assign w1805 = ~shift_3 & ~w64;
assign w1806 = shift_3 & ~w148;
assign w1807 = ~w1805 & ~w1806;
assign w1808 = ~shift_2 & ~w1807;
assign w1809 = shift_2 & ~w1532;
assign w1810 = ~w1808 & ~w1809;
assign w1811 = shift_5 & ~w1810;
assign w1812 = ~w1804 & ~w1811;
assign w1813 = shift_4 & ~w1812;
assign w1814 = ~w1797 & ~w1813;
assign w1815 = shift_6 & w1814;
assign w1816 = ~shift_3 & ~w158;
assign w1817 = shift_3 & ~w198;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = ~shift_2 & ~w1818;
assign w1820 = shift_2 & ~w1543;
assign w1821 = ~w1819 & ~w1820;
assign w1822 = ~shift_5 & ~w1821;
assign w1823 = ~shift_3 & ~w302;
assign w1824 = shift_3 & ~w244;
assign w1825 = ~w1823 & ~w1824;
assign w1826 = ~shift_2 & ~w1825;
assign w1827 = shift_2 & ~w1550;
assign w1828 = ~w1826 & ~w1827;
assign w1829 = shift_5 & ~w1828;
assign w1830 = ~w1822 & ~w1829;
assign w1831 = ~shift_4 & ~w1830;
assign w1832 = ~shift_3 & ~w208;
assign w1833 = shift_3 & ~w292;
assign w1834 = ~w1832 & ~w1833;
assign w1835 = ~shift_2 & ~w1834;
assign w1836 = shift_2 & ~w1559;
assign w1837 = ~w1835 & ~w1836;
assign w1838 = ~shift_5 & ~w1837;
assign w1839 = ~shift_3 & ~w254;
assign w1840 = shift_3 & ~w338;
assign w1841 = ~w1839 & ~w1840;
assign w1842 = ~shift_2 & ~w1841;
assign w1843 = shift_2 & ~w1566;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = shift_5 & ~w1844;
assign w1846 = ~w1838 & ~w1845;
assign w1847 = shift_4 & ~w1846;
assign w1848 = ~w1831 & ~w1847;
assign w1849 = ~shift_6 & w1848;
assign w1850 = ~w1815 & ~w1849;
assign w1851 = ~shift_3 & w726;
assign w1852 = shift_3 & w480;
assign w1853 = ~w1851 & ~w1852;
assign w1854 = ~shift_2 & ~w1853;
assign w1855 = shift_2 & ~w1578;
assign w1856 = ~w1854 & ~w1855;
assign w1857 = ~shift_5 & ~w1856;
assign w1858 = shift_3 & w526;
assign w1859 = ~shift_3 & ~w399;
assign w1860 = ~w1858 & ~w1859;
assign w1861 = ~shift_2 & ~w1860;
assign w1862 = shift_2 & ~w1585;
assign w1863 = ~w1861 & ~w1862;
assign w1864 = shift_5 & ~w1863;
assign w1865 = ~w1857 & ~w1864;
assign w1866 = ~shift_4 & ~w1865;
assign w1867 = ~shift_3 & w490;
assign w1868 = shift_3 & w389;
assign w1869 = ~w1867 & ~w1868;
assign w1870 = ~shift_2 & ~w1869;
assign w1871 = shift_2 & ~w1593;
assign w1872 = ~w1870 & ~w1871;
assign w1873 = ~shift_5 & ~w1872;
assign w1874 = ~shift_3 & w536;
assign w1875 = shift_3 & w432;
assign w1876 = ~w1874 & ~w1875;
assign w1877 = ~shift_2 & ~w1876;
assign w1878 = shift_2 & ~w1601;
assign w1879 = ~w1877 & ~w1878;
assign w1880 = shift_5 & ~w1879;
assign w1881 = ~w1873 & ~w1880;
assign w1882 = shift_4 & ~w1881;
assign w1883 = ~w1866 & ~w1882;
assign w1884 = shift_6 & w1883;
assign w1885 = shift_2 & ~w1612;
assign w1886 = ~shift_3 & w442;
assign w1887 = shift_3 & w576;
assign w1888 = ~w1886 & ~w1887;
assign w1889 = ~shift_2 & ~w1888;
assign w1890 = ~w1885 & ~w1889;
assign w1891 = ~shift_5 & ~w1890;
assign w1892 = ~shift_3 & w680;
assign w1893 = shift_3 & w622;
assign w1894 = ~w1892 & ~w1893;
assign w1895 = ~shift_2 & ~w1894;
assign w1896 = shift_2 & ~w1619;
assign w1897 = ~w1895 & ~w1896;
assign w1898 = shift_5 & ~w1897;
assign w1899 = ~w1891 & ~w1898;
assign w1900 = ~shift_4 & ~w1899;
assign w1901 = shift_2 & ~w1628;
assign w1902 = ~shift_3 & w586;
assign w1903 = shift_3 & w670;
assign w1904 = ~w1902 & ~w1903;
assign w1905 = ~shift_2 & ~w1904;
assign w1906 = ~w1901 & ~w1905;
assign w1907 = ~shift_5 & ~w1906;
assign w1908 = ~shift_3 & w632;
assign w1909 = shift_3 & w716;
assign w1910 = ~w1908 & ~w1909;
assign w1911 = ~shift_2 & ~w1910;
assign w1912 = shift_2 & ~w1635;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = shift_5 & ~w1913;
assign w1915 = ~w1907 & ~w1914;
assign w1916 = shift_4 & ~w1915;
assign w1917 = ~w1900 & ~w1916;
assign w1918 = ~shift_6 & w1917;
assign w1919 = ~w1884 & ~w1918;
assign w1920 = ~shift_3 & ~w1101;
assign w1921 = shift_3 & ~w855;
assign w1922 = ~w1920 & ~w1921;
assign w1923 = ~shift_2 & ~w1922;
assign w1924 = shift_2 & ~w1647;
assign w1925 = ~w1923 & ~w1924;
assign w1926 = ~shift_5 & ~w1925;
assign w1927 = ~shift_3 & ~w774;
assign w1928 = shift_3 & ~w901;
assign w1929 = ~w1927 & ~w1928;
assign w1930 = ~shift_2 & ~w1929;
assign w1931 = shift_2 & ~w1654;
assign w1932 = ~w1930 & ~w1931;
assign w1933 = shift_5 & ~w1932;
assign w1934 = ~w1926 & ~w1933;
assign w1935 = ~shift_4 & ~w1934;
assign w1936 = ~shift_3 & ~w865;
assign w1937 = shift_3 & ~w767;
assign w1938 = ~w1936 & ~w1937;
assign w1939 = ~shift_2 & ~w1938;
assign w1940 = shift_2 & ~w1663;
assign w1941 = ~w1939 & ~w1940;
assign w1942 = ~shift_5 & ~w1941;
assign w1943 = ~shift_3 & ~w911;
assign w1944 = shift_3 & ~w807;
assign w1945 = ~w1943 & ~w1944;
assign w1946 = ~shift_2 & ~w1945;
assign w1947 = shift_2 & ~w1670;
assign w1948 = ~w1946 & ~w1947;
assign w1949 = shift_5 & ~w1948;
assign w1950 = ~w1942 & ~w1949;
assign w1951 = shift_4 & ~w1950;
assign w1952 = ~w1935 & ~w1951;
assign w1953 = shift_6 & w1952;
assign w1954 = ~shift_3 & ~w817;
assign w1955 = shift_3 & ~w951;
assign w1956 = ~w1954 & ~w1955;
assign w1957 = ~shift_2 & ~w1956;
assign w1958 = shift_2 & ~w1681;
assign w1959 = ~w1957 & ~w1958;
assign w1960 = ~shift_5 & ~w1959;
assign w1961 = ~shift_3 & ~w1055;
assign w1962 = shift_3 & ~w997;
assign w1963 = ~w1961 & ~w1962;
assign w1964 = ~shift_2 & ~w1963;
assign w1965 = shift_2 & ~w1688;
assign w1966 = ~w1964 & ~w1965;
assign w1967 = shift_5 & ~w1966;
assign w1968 = ~w1960 & ~w1967;
assign w1969 = ~shift_4 & ~w1968;
assign w1970 = ~shift_3 & ~w961;
assign w1971 = shift_3 & ~w1045;
assign w1972 = ~w1970 & ~w1971;
assign w1973 = ~shift_2 & ~w1972;
assign w1974 = shift_2 & ~w1697;
assign w1975 = ~w1973 & ~w1974;
assign w1976 = ~shift_5 & ~w1975;
assign w1977 = ~shift_3 & ~w1007;
assign w1978 = shift_3 & ~w1091;
assign w1979 = ~w1977 & ~w1978;
assign w1980 = ~shift_2 & ~w1979;
assign w1981 = shift_2 & ~w1704;
assign w1982 = ~w1980 & ~w1981;
assign w1983 = shift_5 & ~w1982;
assign w1984 = ~w1976 & ~w1983;
assign w1985 = shift_4 & ~w1984;
assign w1986 = ~w1969 & ~w1985;
assign w1987 = ~shift_6 & w1986;
assign w1988 = ~w1953 & ~w1987;
assign w1989 = ~shift_3 & w1379;
assign w1990 = shift_3 & w1142;
assign w1991 = ~w1989 & ~w1990;
assign w1992 = ~shift_2 & ~w1991;
assign w1993 = shift_2 & ~w1716;
assign w1994 = ~w1992 & ~w1993;
assign w1995 = ~shift_5 & ~w1994;
assign w1996 = shift_2 & ~w1723;
assign w1997 = ~shift_3 & w1259;
assign w1998 = shift_3 & w1188;
assign w1999 = ~w1997 & ~w1998;
assign w2000 = ~shift_2 & ~w1999;
assign w2001 = ~w1996 & ~w2000;
assign w2002 = shift_5 & ~w2001;
assign w2003 = ~w1995 & ~w2002;
assign w2004 = ~shift_4 & ~w2003;
assign w2005 = ~shift_3 & w1152;
assign w2006 = shift_3 & w1249;
assign w2007 = ~w2005 & ~w2006;
assign w2008 = ~shift_2 & ~w2007;
assign w2009 = shift_2 & ~w1731;
assign w2010 = ~w2008 & ~w2009;
assign w2011 = ~shift_5 & ~w2010;
assign w2012 = ~shift_3 & w1198;
assign w2013 = shift_3 & w1273;
assign w2014 = ~w2012 & ~w2013;
assign w2015 = ~shift_2 & ~w2014;
assign w2016 = shift_2 & ~w1739;
assign w2017 = ~w2015 & ~w2016;
assign w2018 = shift_5 & ~w2017;
assign w2019 = ~w2011 & ~w2018;
assign w2020 = shift_4 & ~w2019;
assign w2021 = ~w2004 & ~w2020;
assign w2022 = shift_6 & w2021;
assign w2023 = shift_2 & ~w1750;
assign w2024 = ~shift_3 & w1283;
assign w2025 = shift_3 & w1417;
assign w2026 = ~w2024 & ~w2025;
assign w2027 = ~shift_2 & ~w2026;
assign w2028 = ~w2023 & ~w2027;
assign w2029 = ~shift_5 & ~w2028;
assign w2030 = shift_2 & ~w1757;
assign w2031 = ~shift_3 & w1333;
assign w2032 = shift_3 & w1463;
assign w2033 = ~w2031 & ~w2032;
assign w2034 = ~shift_2 & ~w2033;
assign w2035 = ~w2030 & ~w2034;
assign w2036 = shift_5 & ~w2035;
assign w2037 = ~w2029 & ~w2036;
assign w2038 = ~shift_4 & ~w2037;
assign w2039 = ~shift_3 & w1427;
assign w2040 = shift_3 & w1323;
assign w2041 = ~w2039 & ~w2040;
assign w2042 = ~shift_2 & ~w2041;
assign w2043 = shift_2 & ~w1766;
assign w2044 = ~w2042 & ~w2043;
assign w2045 = ~shift_5 & ~w2044;
assign w2046 = shift_2 & ~w1773;
assign w2047 = ~shift_3 & w1473;
assign w2048 = shift_3 & w1369;
assign w2049 = ~w2047 & ~w2048;
assign w2050 = ~shift_2 & ~w2049;
assign w2051 = ~w2046 & ~w2050;
assign w2052 = shift_5 & ~w2051;
assign w2053 = ~w2045 & ~w2052;
assign w2054 = shift_4 & ~w2053;
assign w2055 = ~w2038 & ~w2054;
assign w2056 = ~shift_6 & w2055;
assign w2057 = ~w2022 & ~w2056;
assign w2058 = ~shift_2 & ~w372;
assign w2059 = shift_2 & ~w1784;
assign w2060 = ~w2058 & ~w2059;
assign w2061 = ~shift_5 & ~w2060;
assign w2062 = shift_2 & ~w1791;
assign w2063 = ~shift_2 & ~w136;
assign w2064 = ~w2062 & ~w2063;
assign w2065 = shift_5 & ~w2064;
assign w2066 = ~w2061 & ~w2065;
assign w2067 = ~shift_4 & ~w2066;
assign w2068 = ~shift_2 & ~w42;
assign w2069 = shift_2 & ~w1800;
assign w2070 = ~w2068 & ~w2069;
assign w2071 = ~shift_5 & ~w2070;
assign w2072 = ~shift_2 & ~w88;
assign w2073 = shift_2 & ~w1807;
assign w2074 = ~w2072 & ~w2073;
assign w2075 = shift_5 & ~w2074;
assign w2076 = ~w2071 & ~w2075;
assign w2077 = shift_4 & ~w2076;
assign w2078 = ~w2067 & ~w2077;
assign w2079 = shift_6 & w2078;
assign w2080 = ~shift_2 & ~w182;
assign w2081 = shift_2 & ~w1818;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = ~shift_5 & ~w2082;
assign w2084 = ~shift_2 & ~w326;
assign w2085 = shift_2 & ~w1825;
assign w2086 = ~w2084 & ~w2085;
assign w2087 = shift_5 & ~w2086;
assign w2088 = ~w2083 & ~w2087;
assign w2089 = ~shift_4 & ~w2088;
assign w2090 = ~shift_2 & ~w232;
assign w2091 = shift_2 & ~w1834;
assign w2092 = ~w2090 & ~w2091;
assign w2093 = ~shift_5 & ~w2092;
assign w2094 = ~shift_2 & ~w278;
assign w2095 = shift_2 & ~w1841;
assign w2096 = ~w2094 & ~w2095;
assign w2097 = shift_5 & ~w2096;
assign w2098 = ~w2093 & ~w2097;
assign w2099 = shift_4 & ~w2098;
assign w2100 = ~w2089 & ~w2099;
assign w2101 = ~shift_6 & w2100;
assign w2102 = ~w2079 & ~w2101;
assign w2103 = shift_2 & ~w1853;
assign w2104 = ~shift_2 & ~w750;
assign w2105 = ~w2103 & ~w2104;
assign w2106 = ~shift_5 & ~w2105;
assign w2107 = ~shift_2 & ~w420;
assign w2108 = shift_2 & ~w1860;
assign w2109 = ~w2107 & ~w2108;
assign w2110 = shift_5 & ~w2109;
assign w2111 = ~w2106 & ~w2110;
assign w2112 = ~shift_4 & ~w2111;
assign w2113 = ~shift_2 & ~w514;
assign w2114 = shift_2 & ~w1869;
assign w2115 = ~w2113 & ~w2114;
assign w2116 = ~shift_5 & ~w2115;
assign w2117 = shift_2 & ~w1876;
assign w2118 = ~shift_2 & ~w560;
assign w2119 = ~w2117 & ~w2118;
assign w2120 = shift_5 & ~w2119;
assign w2121 = ~w2116 & ~w2120;
assign w2122 = shift_4 & ~w2121;
assign w2123 = ~w2112 & ~w2122;
assign w2124 = shift_6 & w2123;
assign w2125 = ~shift_2 & ~w466;
assign w2126 = shift_2 & ~w1888;
assign w2127 = ~w2125 & ~w2126;
assign w2128 = ~shift_5 & ~w2127;
assign w2129 = shift_2 & ~w1894;
assign w2130 = ~shift_2 & ~w704;
assign w2131 = ~w2129 & ~w2130;
assign w2132 = shift_5 & ~w2131;
assign w2133 = ~w2128 & ~w2132;
assign w2134 = ~shift_4 & ~w2133;
assign w2135 = ~shift_2 & ~w610;
assign w2136 = shift_2 & ~w1904;
assign w2137 = ~w2135 & ~w2136;
assign w2138 = ~shift_5 & ~w2137;
assign w2139 = shift_2 & ~w1910;
assign w2140 = ~shift_2 & ~w656;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = shift_5 & ~w2141;
assign w2143 = ~w2138 & ~w2142;
assign w2144 = shift_4 & ~w2143;
assign w2145 = ~w2134 & ~w2144;
assign w2146 = ~shift_6 & w2145;
assign w2147 = ~w2124 & ~w2146;
assign w2148 = ~shift_2 & ~w1125;
assign w2149 = shift_2 & ~w1922;
assign w2150 = ~w2148 & ~w2149;
assign w2151 = ~shift_5 & ~w2150;
assign w2152 = ~shift_2 & ~w795;
assign w2153 = shift_2 & ~w1929;
assign w2154 = ~w2152 & ~w2153;
assign w2155 = shift_5 & ~w2154;
assign w2156 = ~w2151 & ~w2155;
assign w2157 = ~shift_4 & ~w2156;
assign w2158 = ~shift_2 & ~w889;
assign w2159 = shift_2 & ~w1938;
assign w2160 = ~w2158 & ~w2159;
assign w2161 = ~shift_5 & ~w2160;
assign w2162 = ~shift_2 & ~w935;
assign w2163 = shift_2 & ~w1945;
assign w2164 = ~w2162 & ~w2163;
assign w2165 = shift_5 & ~w2164;
assign w2166 = ~w2161 & ~w2165;
assign w2167 = shift_4 & ~w2166;
assign w2168 = ~w2157 & ~w2167;
assign w2169 = shift_6 & w2168;
assign w2170 = ~shift_2 & ~w841;
assign w2171 = shift_2 & ~w1956;
assign w2172 = ~w2170 & ~w2171;
assign w2173 = ~shift_5 & ~w2172;
assign w2174 = ~shift_2 & ~w1079;
assign w2175 = shift_2 & ~w1963;
assign w2176 = ~w2174 & ~w2175;
assign w2177 = shift_5 & ~w2176;
assign w2178 = ~w2173 & ~w2177;
assign w2179 = ~shift_4 & ~w2178;
assign w2180 = ~shift_2 & ~w985;
assign w2181 = shift_2 & ~w1972;
assign w2182 = ~w2180 & ~w2181;
assign w2183 = ~shift_5 & ~w2182;
assign w2184 = ~shift_2 & ~w1031;
assign w2185 = shift_2 & ~w1979;
assign w2186 = ~w2184 & ~w2185;
assign w2187 = shift_5 & ~w2186;
assign w2188 = ~w2183 & ~w2187;
assign w2189 = shift_4 & ~w2188;
assign w2190 = ~w2179 & ~w2189;
assign w2191 = ~shift_6 & w2190;
assign w2192 = ~w2169 & ~w2191;
assign w2193 = shift_2 & ~w1991;
assign w2194 = ~shift_2 & ~w1403;
assign w2195 = ~w2193 & ~w2194;
assign w2196 = ~shift_5 & ~w2195;
assign w2197 = ~shift_2 & ~w1239;
assign w2198 = shift_2 & ~w1999;
assign w2199 = ~w2197 & ~w2198;
assign w2200 = shift_5 & ~w2199;
assign w2201 = ~w2196 & ~w2200;
assign w2202 = ~shift_4 & ~w2201;
assign w2203 = ~shift_2 & ~w1176;
assign w2204 = shift_2 & ~w2007;
assign w2205 = ~w2203 & ~w2204;
assign w2206 = ~shift_5 & ~w2205;
assign w2207 = shift_2 & ~w2014;
assign w2208 = ~shift_2 & ~w1222;
assign w2209 = ~w2207 & ~w2208;
assign w2210 = shift_5 & ~w2209;
assign w2211 = ~w2206 & ~w2210;
assign w2212 = shift_4 & ~w2211;
assign w2213 = ~w2202 & ~w2212;
assign w2214 = shift_6 & w2213;
assign w2215 = ~shift_2 & ~w1307;
assign w2216 = shift_2 & ~w2026;
assign w2217 = ~w2215 & ~w2216;
assign w2218 = ~shift_5 & ~w2217;
assign w2219 = ~shift_2 & ~w1357;
assign w2220 = shift_2 & ~w2033;
assign w2221 = ~w2219 & ~w2220;
assign w2222 = shift_5 & ~w2221;
assign w2223 = ~w2218 & ~w2222;
assign w2224 = ~shift_4 & ~w2223;
assign w2225 = shift_2 & ~w2041;
assign w2226 = ~shift_2 & ~w1451;
assign w2227 = ~w2225 & ~w2226;
assign w2228 = ~shift_5 & ~w2227;
assign w2229 = ~shift_2 & ~w1497;
assign w2230 = shift_2 & ~w2049;
assign w2231 = ~w2229 & ~w2230;
assign w2232 = shift_5 & ~w2231;
assign w2233 = ~w2228 & ~w2232;
assign w2234 = shift_4 & ~w2233;
assign w2235 = ~w2224 & ~w2234;
assign w2236 = ~shift_6 & w2235;
assign w2237 = ~w2214 & ~w2236;
assign w2238 = shift_5 & ~w138;
assign w2239 = ~shift_5 & ~w374;
assign w2240 = ~w2238 & ~w2239;
assign w2241 = ~shift_4 & ~w2240;
assign w2242 = shift_4 & ~w92;
assign w2243 = ~w2241 & ~w2242;
assign w2244 = shift_6 & w2243;
assign w2245 = shift_4 & ~w282;
assign w2246 = ~shift_5 & ~w184;
assign w2247 = shift_5 & ~w328;
assign w2248 = ~w2246 & ~w2247;
assign w2249 = ~shift_4 & ~w2248;
assign w2250 = ~w2245 & ~w2249;
assign w2251 = ~shift_6 & w2250;
assign w2252 = ~w2244 & ~w2251;
assign w2253 = shift_4 & ~w564;
assign w2254 = shift_5 & ~w422;
assign w2255 = ~shift_5 & ~w752;
assign w2256 = ~w2254 & ~w2255;
assign w2257 = ~shift_4 & ~w2256;
assign w2258 = ~w2253 & ~w2257;
assign w2259 = shift_6 & w2258;
assign w2260 = shift_4 & ~w660;
assign w2261 = ~shift_5 & ~w468;
assign w2262 = shift_5 & ~w706;
assign w2263 = ~w2261 & ~w2262;
assign w2264 = ~shift_4 & ~w2263;
assign w2265 = ~w2260 & ~w2264;
assign w2266 = ~shift_6 & w2265;
assign w2267 = ~w2259 & ~w2266;
assign w2268 = shift_4 & ~w939;
assign w2269 = shift_5 & ~w797;
assign w2270 = ~shift_5 & ~w1127;
assign w2271 = ~w2269 & ~w2270;
assign w2272 = ~shift_4 & ~w2271;
assign w2273 = ~w2268 & ~w2272;
assign w2274 = shift_6 & w2273;
assign w2275 = shift_4 & ~w1035;
assign w2276 = ~shift_5 & ~w843;
assign w2277 = shift_5 & ~w1081;
assign w2278 = ~w2276 & ~w2277;
assign w2279 = ~shift_4 & ~w2278;
assign w2280 = ~w2275 & ~w2279;
assign w2281 = ~shift_6 & w2280;
assign w2282 = ~w2274 & ~w2281;
assign w2283 = shift_4 & ~w1226;
assign w2284 = shift_5 & ~w1263;
assign w2285 = ~shift_5 & ~w1405;
assign w2286 = ~w2284 & ~w2285;
assign w2287 = ~shift_4 & ~w2286;
assign w2288 = ~w2283 & ~w2287;
assign w2289 = shift_6 & w2288;
assign w2290 = shift_4 & ~w1501;
assign w2291 = ~shift_5 & ~w1309;
assign w2292 = shift_5 & ~w1359;
assign w2293 = ~w2291 & ~w2292;
assign w2294 = ~shift_4 & ~w2293;
assign w2295 = ~w2290 & ~w2294;
assign w2296 = ~shift_6 & w2295;
assign w2297 = ~w2289 & ~w2296;
assign w2298 = ~shift_5 & ~w1568;
assign w2299 = shift_5 & ~w1527;
assign w2300 = ~w2298 & ~w2299;
assign w2301 = ~shift_4 & ~w2300;
assign w2302 = shift_4 & ~w1520;
assign w2303 = ~w2301 & ~w2302;
assign w2304 = shift_6 & w2303;
assign w2305 = shift_4 & ~w1554;
assign w2306 = ~shift_5 & ~w1534;
assign w2307 = shift_5 & ~w1561;
assign w2308 = ~w2306 & ~w2307;
assign w2309 = ~shift_4 & ~w2308;
assign w2310 = ~w2305 & ~w2309;
assign w2311 = ~shift_6 & w2310;
assign w2312 = ~w2304 & ~w2311;
assign w2313 = ~shift_5 & ~w1637;
assign w2314 = shift_5 & ~w1596;
assign w2315 = ~w2313 & ~w2314;
assign w2316 = ~shift_4 & ~w2315;
assign w2317 = shift_4 & ~w1589;
assign w2318 = ~w2316 & ~w2317;
assign w2319 = shift_6 & w2318;
assign w2320 = shift_4 & ~w1623;
assign w2321 = ~shift_5 & ~w1603;
assign w2322 = shift_5 & ~w1630;
assign w2323 = ~w2321 & ~w2322;
assign w2324 = ~shift_4 & ~w2323;
assign w2325 = ~w2320 & ~w2324;
assign w2326 = ~shift_6 & w2325;
assign w2327 = ~w2319 & ~w2326;
assign w2328 = ~shift_5 & ~w1706;
assign w2329 = shift_5 & ~w1665;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = ~shift_4 & ~w2330;
assign w2332 = shift_4 & ~w1658;
assign w2333 = ~w2331 & ~w2332;
assign w2334 = shift_6 & w2333;
assign w2335 = shift_4 & ~w1692;
assign w2336 = ~shift_5 & ~w1672;
assign w2337 = shift_5 & ~w1699;
assign w2338 = ~w2336 & ~w2337;
assign w2339 = ~shift_4 & ~w2338;
assign w2340 = ~w2335 & ~w2339;
assign w2341 = ~shift_6 & w2340;
assign w2342 = ~w2334 & ~w2341;
assign w2343 = ~shift_5 & ~w1775;
assign w2344 = shift_5 & ~w1734;
assign w2345 = ~w2343 & ~w2344;
assign w2346 = ~shift_4 & ~w2345;
assign w2347 = shift_4 & ~w1727;
assign w2348 = ~w2346 & ~w2347;
assign w2349 = shift_6 & w2348;
assign w2350 = shift_4 & ~w1761;
assign w2351 = ~shift_5 & ~w1741;
assign w2352 = shift_5 & ~w1768;
assign w2353 = ~w2351 & ~w2352;
assign w2354 = ~shift_4 & ~w2353;
assign w2355 = ~w2350 & ~w2354;
assign w2356 = ~shift_6 & w2355;
assign w2357 = ~w2349 & ~w2356;
assign w2358 = ~shift_5 & ~w1844;
assign w2359 = shift_5 & ~w1803;
assign w2360 = ~w2358 & ~w2359;
assign w2361 = ~shift_4 & ~w2360;
assign w2362 = shift_4 & ~w1796;
assign w2363 = ~w2361 & ~w2362;
assign w2364 = shift_6 & w2363;
assign w2365 = shift_4 & ~w1830;
assign w2366 = ~shift_5 & ~w1810;
assign w2367 = shift_5 & ~w1837;
assign w2368 = ~w2366 & ~w2367;
assign w2369 = ~shift_4 & ~w2368;
assign w2370 = ~w2365 & ~w2369;
assign w2371 = ~shift_6 & w2370;
assign w2372 = ~w2364 & ~w2371;
assign w2373 = ~shift_5 & ~w1913;
assign w2374 = shift_5 & ~w1872;
assign w2375 = ~w2373 & ~w2374;
assign w2376 = ~shift_4 & ~w2375;
assign w2377 = shift_4 & ~w1865;
assign w2378 = ~w2376 & ~w2377;
assign w2379 = shift_6 & w2378;
assign w2380 = shift_4 & ~w1899;
assign w2381 = ~shift_5 & ~w1879;
assign w2382 = shift_5 & ~w1906;
assign w2383 = ~w2381 & ~w2382;
assign w2384 = ~shift_4 & ~w2383;
assign w2385 = ~w2380 & ~w2384;
assign w2386 = ~shift_6 & w2385;
assign w2387 = ~w2379 & ~w2386;
assign w2388 = ~shift_5 & ~w1982;
assign w2389 = shift_5 & ~w1941;
assign w2390 = ~w2388 & ~w2389;
assign w2391 = ~shift_4 & ~w2390;
assign w2392 = shift_4 & ~w1934;
assign w2393 = ~w2391 & ~w2392;
assign w2394 = shift_6 & w2393;
assign w2395 = shift_4 & ~w1968;
assign w2396 = ~shift_5 & ~w1948;
assign w2397 = shift_5 & ~w1975;
assign w2398 = ~w2396 & ~w2397;
assign w2399 = ~shift_4 & ~w2398;
assign w2400 = ~w2395 & ~w2399;
assign w2401 = ~shift_6 & w2400;
assign w2402 = ~w2394 & ~w2401;
assign w2403 = ~shift_5 & ~w2051;
assign w2404 = shift_5 & ~w2010;
assign w2405 = ~w2403 & ~w2404;
assign w2406 = ~shift_4 & ~w2405;
assign w2407 = shift_4 & ~w2003;
assign w2408 = ~w2406 & ~w2407;
assign w2409 = shift_6 & w2408;
assign w2410 = shift_4 & ~w2037;
assign w2411 = ~shift_5 & ~w2017;
assign w2412 = shift_5 & ~w2044;
assign w2413 = ~w2411 & ~w2412;
assign w2414 = ~shift_4 & ~w2413;
assign w2415 = ~w2410 & ~w2414;
assign w2416 = ~shift_6 & w2415;
assign w2417 = ~w2409 & ~w2416;
assign w2418 = ~shift_5 & ~w2096;
assign w2419 = shift_5 & ~w2070;
assign w2420 = ~w2418 & ~w2419;
assign w2421 = ~shift_4 & ~w2420;
assign w2422 = shift_4 & ~w2066;
assign w2423 = ~w2421 & ~w2422;
assign w2424 = shift_6 & w2423;
assign w2425 = shift_4 & ~w2088;
assign w2426 = ~shift_5 & ~w2074;
assign w2427 = shift_5 & ~w2092;
assign w2428 = ~w2426 & ~w2427;
assign w2429 = ~shift_4 & ~w2428;
assign w2430 = ~w2425 & ~w2429;
assign w2431 = ~shift_6 & w2430;
assign w2432 = ~w2424 & ~w2431;
assign w2433 = ~shift_5 & ~w2141;
assign w2434 = shift_5 & ~w2115;
assign w2435 = ~w2433 & ~w2434;
assign w2436 = ~shift_4 & ~w2435;
assign w2437 = shift_4 & ~w2111;
assign w2438 = ~w2436 & ~w2437;
assign w2439 = shift_6 & w2438;
assign w2440 = shift_4 & ~w2133;
assign w2441 = ~shift_5 & ~w2119;
assign w2442 = shift_5 & ~w2137;
assign w2443 = ~w2441 & ~w2442;
assign w2444 = ~shift_4 & ~w2443;
assign w2445 = ~w2440 & ~w2444;
assign w2446 = ~shift_6 & w2445;
assign w2447 = ~w2439 & ~w2446;
assign w2448 = ~shift_5 & ~w2186;
assign w2449 = shift_5 & ~w2160;
assign w2450 = ~w2448 & ~w2449;
assign w2451 = ~shift_4 & ~w2450;
assign w2452 = shift_4 & ~w2156;
assign w2453 = ~w2451 & ~w2452;
assign w2454 = shift_6 & w2453;
assign w2455 = shift_4 & ~w2178;
assign w2456 = ~shift_5 & ~w2164;
assign w2457 = shift_5 & ~w2182;
assign w2458 = ~w2456 & ~w2457;
assign w2459 = ~shift_4 & ~w2458;
assign w2460 = ~w2455 & ~w2459;
assign w2461 = ~shift_6 & w2460;
assign w2462 = ~w2454 & ~w2461;
assign w2463 = ~shift_5 & ~w2231;
assign w2464 = shift_5 & ~w2205;
assign w2465 = ~w2463 & ~w2464;
assign w2466 = ~shift_4 & ~w2465;
assign w2467 = shift_4 & ~w2201;
assign w2468 = ~w2466 & ~w2467;
assign w2469 = shift_6 & w2468;
assign w2470 = shift_4 & ~w2223;
assign w2471 = ~shift_5 & ~w2209;
assign w2472 = shift_5 & ~w2227;
assign w2473 = ~w2471 & ~w2472;
assign w2474 = ~shift_4 & ~w2473;
assign w2475 = ~w2470 & ~w2474;
assign w2476 = ~shift_6 & w2475;
assign w2477 = ~w2469 & ~w2476;
assign w2478 = ~shift_5 & ~w280;
assign w2479 = shift_5 & ~w44;
assign w2480 = ~w2478 & ~w2479;
assign w2481 = ~shift_4 & ~w2480;
assign w2482 = shift_4 & ~w2240;
assign w2483 = ~w2481 & ~w2482;
assign w2484 = shift_6 & w2483;
assign w2485 = ~shift_5 & ~w90;
assign w2486 = shift_5 & ~w234;
assign w2487 = ~w2485 & ~w2486;
assign w2488 = ~shift_4 & ~w2487;
assign w2489 = shift_4 & ~w2248;
assign w2490 = ~w2488 & ~w2489;
assign w2491 = ~shift_6 & w2490;
assign w2492 = ~w2484 & ~w2491;
assign w2493 = ~shift_5 & ~w658;
assign w2494 = shift_5 & ~w516;
assign w2495 = ~w2493 & ~w2494;
assign w2496 = ~shift_4 & ~w2495;
assign w2497 = shift_4 & ~w2256;
assign w2498 = ~w2496 & ~w2497;
assign w2499 = shift_6 & w2498;
assign w2500 = ~shift_5 & ~w562;
assign w2501 = shift_5 & ~w612;
assign w2502 = ~w2500 & ~w2501;
assign w2503 = ~shift_4 & ~w2502;
assign w2504 = shift_4 & ~w2263;
assign w2505 = ~w2503 & ~w2504;
assign w2506 = ~shift_6 & w2505;
assign w2507 = ~w2499 & ~w2506;
assign w2508 = ~shift_5 & ~w1033;
assign w2509 = shift_5 & ~w891;
assign w2510 = ~w2508 & ~w2509;
assign w2511 = ~shift_4 & ~w2510;
assign w2512 = shift_4 & ~w2271;
assign w2513 = ~w2511 & ~w2512;
assign w2514 = shift_6 & w2513;
assign w2515 = ~shift_5 & ~w937;
assign w2516 = shift_5 & ~w987;
assign w2517 = ~w2515 & ~w2516;
assign w2518 = ~shift_4 & ~w2517;
assign w2519 = shift_4 & ~w2278;
assign w2520 = ~w2518 & ~w2519;
assign w2521 = ~shift_6 & w2520;
assign w2522 = ~w2514 & ~w2521;
assign w2523 = ~shift_5 & ~w1499;
assign w2524 = shift_5 & ~w1178;
assign w2525 = ~w2523 & ~w2524;
assign w2526 = ~shift_4 & ~w2525;
assign w2527 = shift_4 & ~w2286;
assign w2528 = ~w2526 & ~w2527;
assign w2529 = shift_6 & w2528;
assign w2530 = shift_5 & ~w1453;
assign w2531 = ~shift_5 & ~w1224;
assign w2532 = ~w2530 & ~w2531;
assign w2533 = ~shift_4 & ~w2532;
assign w2534 = shift_4 & ~w2293;
assign w2535 = ~w2533 & ~w2534;
assign w2536 = ~shift_6 & w2535;
assign w2537 = ~w2529 & ~w2536;
assign w2538 = shift_5 & ~w1511;
assign w2539 = ~shift_5 & ~w1552;
assign w2540 = ~w2538 & ~w2539;
assign w2541 = ~shift_4 & ~w2540;
assign w2542 = shift_4 & ~w2300;
assign w2543 = ~w2541 & ~w2542;
assign w2544 = shift_6 & w2543;
assign w2545 = shift_4 & ~w2308;
assign w2546 = ~shift_5 & ~w1518;
assign w2547 = shift_5 & ~w1545;
assign w2548 = ~w2546 & ~w2547;
assign w2549 = ~shift_4 & ~w2548;
assign w2550 = ~w2545 & ~w2549;
assign w2551 = ~shift_6 & w2550;
assign w2552 = ~w2544 & ~w2551;
assign w2553 = shift_5 & ~w1580;
assign w2554 = ~shift_5 & ~w1621;
assign w2555 = ~w2553 & ~w2554;
assign w2556 = ~shift_4 & ~w2555;
assign w2557 = shift_4 & ~w2315;
assign w2558 = ~w2556 & ~w2557;
assign w2559 = shift_6 & w2558;
assign w2560 = shift_4 & ~w2323;
assign w2561 = ~shift_5 & ~w1587;
assign w2562 = shift_5 & ~w1614;
assign w2563 = ~w2561 & ~w2562;
assign w2564 = ~shift_4 & ~w2563;
assign w2565 = ~w2560 & ~w2564;
assign w2566 = ~shift_6 & w2565;
assign w2567 = ~w2559 & ~w2566;
assign w2568 = shift_5 & ~w1649;
assign w2569 = ~shift_5 & ~w1690;
assign w2570 = ~w2568 & ~w2569;
assign w2571 = ~shift_4 & ~w2570;
assign w2572 = shift_4 & ~w2330;
assign w2573 = ~w2571 & ~w2572;
assign w2574 = shift_6 & w2573;
assign w2575 = shift_4 & ~w2338;
assign w2576 = ~shift_5 & ~w1656;
assign w2577 = shift_5 & ~w1683;
assign w2578 = ~w2576 & ~w2577;
assign w2579 = ~shift_4 & ~w2578;
assign w2580 = ~w2575 & ~w2579;
assign w2581 = ~shift_6 & w2580;
assign w2582 = ~w2574 & ~w2581;
assign w2583 = shift_5 & ~w1718;
assign w2584 = ~shift_5 & ~w1759;
assign w2585 = ~w2583 & ~w2584;
assign w2586 = ~shift_4 & ~w2585;
assign w2587 = shift_4 & ~w2345;
assign w2588 = ~w2586 & ~w2587;
assign w2589 = shift_6 & w2588;
assign w2590 = shift_4 & ~w2353;
assign w2591 = ~shift_5 & ~w1725;
assign w2592 = shift_5 & ~w1752;
assign w2593 = ~w2591 & ~w2592;
assign w2594 = ~shift_4 & ~w2593;
assign w2595 = ~w2590 & ~w2594;
assign w2596 = ~shift_6 & w2595;
assign w2597 = ~w2589 & ~w2596;
assign w2598 = shift_5 & ~w1787;
assign w2599 = ~shift_5 & ~w1828;
assign w2600 = ~w2598 & ~w2599;
assign w2601 = ~shift_4 & ~w2600;
assign w2602 = shift_4 & ~w2360;
assign w2603 = ~w2601 & ~w2602;
assign w2604 = shift_6 & w2603;
assign w2605 = shift_4 & ~w2368;
assign w2606 = ~shift_5 & ~w1794;
assign w2607 = shift_5 & ~w1821;
assign w2608 = ~w2606 & ~w2607;
assign w2609 = ~shift_4 & ~w2608;
assign w2610 = ~w2605 & ~w2609;
assign w2611 = ~shift_6 & w2610;
assign w2612 = ~w2604 & ~w2611;
assign w2613 = shift_5 & ~w1856;
assign w2614 = ~shift_5 & ~w1897;
assign w2615 = ~w2613 & ~w2614;
assign w2616 = ~shift_4 & ~w2615;
assign w2617 = shift_4 & ~w2375;
assign w2618 = ~w2616 & ~w2617;
assign w2619 = shift_6 & w2618;
assign w2620 = shift_4 & ~w2383;
assign w2621 = ~shift_5 & ~w1863;
assign w2622 = shift_5 & ~w1890;
assign w2623 = ~w2621 & ~w2622;
assign w2624 = ~shift_4 & ~w2623;
assign w2625 = ~w2620 & ~w2624;
assign w2626 = ~shift_6 & w2625;
assign w2627 = ~w2619 & ~w2626;
assign w2628 = shift_5 & ~w1925;
assign w2629 = ~shift_5 & ~w1966;
assign w2630 = ~w2628 & ~w2629;
assign w2631 = ~shift_4 & ~w2630;
assign w2632 = shift_4 & ~w2390;
assign w2633 = ~w2631 & ~w2632;
assign w2634 = shift_6 & w2633;
assign w2635 = shift_4 & ~w2398;
assign w2636 = ~shift_5 & ~w1932;
assign w2637 = shift_5 & ~w1959;
assign w2638 = ~w2636 & ~w2637;
assign w2639 = ~shift_4 & ~w2638;
assign w2640 = ~w2635 & ~w2639;
assign w2641 = ~shift_6 & w2640;
assign w2642 = ~w2634 & ~w2641;
assign w2643 = shift_5 & ~w1994;
assign w2644 = ~shift_5 & ~w2035;
assign w2645 = ~w2643 & ~w2644;
assign w2646 = ~shift_4 & ~w2645;
assign w2647 = shift_4 & ~w2405;
assign w2648 = ~w2646 & ~w2647;
assign w2649 = shift_6 & w2648;
assign w2650 = shift_4 & ~w2413;
assign w2651 = ~shift_5 & ~w2001;
assign w2652 = shift_5 & ~w2028;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = ~shift_4 & ~w2653;
assign w2655 = ~w2650 & ~w2654;
assign w2656 = ~shift_6 & w2655;
assign w2657 = ~w2649 & ~w2656;
assign w2658 = shift_5 & ~w2060;
assign w2659 = ~shift_5 & ~w2086;
assign w2660 = ~w2658 & ~w2659;
assign w2661 = ~shift_4 & ~w2660;
assign w2662 = shift_4 & ~w2420;
assign w2663 = ~w2661 & ~w2662;
assign w2664 = shift_6 & w2663;
assign w2665 = shift_4 & ~w2428;
assign w2666 = ~shift_5 & ~w2064;
assign w2667 = shift_5 & ~w2082;
assign w2668 = ~w2666 & ~w2667;
assign w2669 = ~shift_4 & ~w2668;
assign w2670 = ~w2665 & ~w2669;
assign w2671 = ~shift_6 & w2670;
assign w2672 = ~w2664 & ~w2671;
assign w2673 = shift_5 & ~w2105;
assign w2674 = ~shift_5 & ~w2131;
assign w2675 = ~w2673 & ~w2674;
assign w2676 = ~shift_4 & ~w2675;
assign w2677 = shift_4 & ~w2435;
assign w2678 = ~w2676 & ~w2677;
assign w2679 = shift_6 & w2678;
assign w2680 = shift_4 & ~w2443;
assign w2681 = ~shift_5 & ~w2109;
assign w2682 = shift_5 & ~w2127;
assign w2683 = ~w2681 & ~w2682;
assign w2684 = ~shift_4 & ~w2683;
assign w2685 = ~w2680 & ~w2684;
assign w2686 = ~shift_6 & w2685;
assign w2687 = ~w2679 & ~w2686;
assign w2688 = shift_5 & ~w2150;
assign w2689 = ~shift_5 & ~w2176;
assign w2690 = ~w2688 & ~w2689;
assign w2691 = ~shift_4 & ~w2690;
assign w2692 = shift_4 & ~w2450;
assign w2693 = ~w2691 & ~w2692;
assign w2694 = shift_6 & w2693;
assign w2695 = shift_4 & ~w2458;
assign w2696 = ~shift_5 & ~w2154;
assign w2697 = shift_5 & ~w2172;
assign w2698 = ~w2696 & ~w2697;
assign w2699 = ~shift_4 & ~w2698;
assign w2700 = ~w2695 & ~w2699;
assign w2701 = ~shift_6 & w2700;
assign w2702 = ~w2694 & ~w2701;
assign w2703 = shift_5 & ~w2195;
assign w2704 = ~shift_5 & ~w2221;
assign w2705 = ~w2703 & ~w2704;
assign w2706 = ~shift_4 & ~w2705;
assign w2707 = shift_4 & ~w2465;
assign w2708 = ~w2706 & ~w2707;
assign w2709 = shift_6 & w2708;
assign w2710 = shift_4 & ~w2473;
assign w2711 = ~shift_5 & ~w2199;
assign w2712 = shift_5 & ~w2217;
assign w2713 = ~w2711 & ~w2712;
assign w2714 = ~shift_4 & ~w2713;
assign w2715 = ~w2710 & ~w2714;
assign w2716 = ~shift_6 & w2715;
assign w2717 = ~w2709 & ~w2716;
assign w2718 = ~shift_4 & ~w376;
assign w2719 = shift_4 & ~w2480;
assign w2720 = ~w2718 & ~w2719;
assign w2721 = shift_6 & w2720;
assign w2722 = ~shift_4 & ~w186;
assign w2723 = shift_4 & ~w2487;
assign w2724 = ~w2722 & ~w2723;
assign w2725 = ~shift_6 & w2724;
assign w2726 = ~w2721 & ~w2725;
assign w2727 = ~shift_4 & ~w754;
assign w2728 = shift_4 & ~w2495;
assign w2729 = ~w2727 & ~w2728;
assign w2730 = shift_6 & w2729;
assign w2731 = ~shift_4 & ~w470;
assign w2732 = shift_4 & ~w2502;
assign w2733 = ~w2731 & ~w2732;
assign w2734 = ~shift_6 & w2733;
assign w2735 = ~w2730 & ~w2734;
assign w2736 = ~shift_4 & ~w1129;
assign w2737 = shift_4 & ~w2510;
assign w2738 = ~w2736 & ~w2737;
assign w2739 = shift_6 & w2738;
assign w2740 = ~shift_4 & ~w845;
assign w2741 = shift_4 & ~w2517;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = ~shift_6 & w2742;
assign w2744 = ~w2739 & ~w2743;
assign w2745 = ~shift_4 & ~w1407;
assign w2746 = shift_4 & ~w2525;
assign w2747 = ~w2745 & ~w2746;
assign w2748 = shift_6 & w2747;
assign w2749 = ~shift_4 & ~w1311;
assign w2750 = shift_4 & ~w2532;
assign w2751 = ~w2749 & ~w2750;
assign w2752 = ~shift_6 & w2751;
assign w2753 = ~w2748 & ~w2752;
assign w2754 = ~shift_4 & ~w1570;
assign w2755 = shift_4 & ~w2540;
assign w2756 = ~w2754 & ~w2755;
assign w2757 = shift_6 & w2756;
assign w2758 = shift_4 & ~w2548;
assign w2759 = ~shift_4 & ~w1536;
assign w2760 = ~w2758 & ~w2759;
assign w2761 = ~shift_6 & w2760;
assign w2762 = ~w2757 & ~w2761;
assign w2763 = ~shift_4 & ~w1639;
assign w2764 = shift_4 & ~w2555;
assign w2765 = ~w2763 & ~w2764;
assign w2766 = shift_6 & w2765;
assign w2767 = shift_4 & ~w2563;
assign w2768 = ~shift_4 & ~w1605;
assign w2769 = ~w2767 & ~w2768;
assign w2770 = ~shift_6 & w2769;
assign w2771 = ~w2766 & ~w2770;
assign w2772 = ~shift_4 & ~w1708;
assign w2773 = shift_4 & ~w2570;
assign w2774 = ~w2772 & ~w2773;
assign w2775 = shift_6 & w2774;
assign w2776 = shift_4 & ~w2578;
assign w2777 = ~shift_4 & ~w1674;
assign w2778 = ~w2776 & ~w2777;
assign w2779 = ~shift_6 & w2778;
assign w2780 = ~w2775 & ~w2779;
assign w2781 = ~shift_4 & ~w1777;
assign w2782 = shift_4 & ~w2585;
assign w2783 = ~w2781 & ~w2782;
assign w2784 = shift_6 & w2783;
assign w2785 = shift_4 & ~w2593;
assign w2786 = ~shift_4 & ~w1743;
assign w2787 = ~w2785 & ~w2786;
assign w2788 = ~shift_6 & w2787;
assign w2789 = ~w2784 & ~w2788;
assign w2790 = ~shift_4 & ~w1846;
assign w2791 = shift_4 & ~w2600;
assign w2792 = ~w2790 & ~w2791;
assign w2793 = shift_6 & w2792;
assign w2794 = shift_4 & ~w2608;
assign w2795 = ~shift_4 & ~w1812;
assign w2796 = ~w2794 & ~w2795;
assign w2797 = ~shift_6 & w2796;
assign w2798 = ~w2793 & ~w2797;
assign w2799 = ~shift_4 & ~w1915;
assign w2800 = shift_4 & ~w2615;
assign w2801 = ~w2799 & ~w2800;
assign w2802 = shift_6 & w2801;
assign w2803 = shift_4 & ~w2623;
assign w2804 = ~shift_4 & ~w1881;
assign w2805 = ~w2803 & ~w2804;
assign w2806 = ~shift_6 & w2805;
assign w2807 = ~w2802 & ~w2806;
assign w2808 = ~shift_4 & ~w1984;
assign w2809 = shift_4 & ~w2630;
assign w2810 = ~w2808 & ~w2809;
assign w2811 = shift_6 & w2810;
assign w2812 = shift_4 & ~w2638;
assign w2813 = ~shift_4 & ~w1950;
assign w2814 = ~w2812 & ~w2813;
assign w2815 = ~shift_6 & w2814;
assign w2816 = ~w2811 & ~w2815;
assign w2817 = ~shift_4 & ~w2053;
assign w2818 = shift_4 & ~w2645;
assign w2819 = ~w2817 & ~w2818;
assign w2820 = shift_6 & w2819;
assign w2821 = shift_4 & ~w2653;
assign w2822 = ~shift_4 & ~w2019;
assign w2823 = ~w2821 & ~w2822;
assign w2824 = ~shift_6 & w2823;
assign w2825 = ~w2820 & ~w2824;
assign w2826 = ~shift_4 & ~w2098;
assign w2827 = shift_4 & ~w2660;
assign w2828 = ~w2826 & ~w2827;
assign w2829 = shift_6 & w2828;
assign w2830 = shift_4 & ~w2668;
assign w2831 = ~shift_4 & ~w2076;
assign w2832 = ~w2830 & ~w2831;
assign w2833 = ~shift_6 & w2832;
assign w2834 = ~w2829 & ~w2833;
assign w2835 = ~shift_4 & ~w2143;
assign w2836 = shift_4 & ~w2675;
assign w2837 = ~w2835 & ~w2836;
assign w2838 = shift_6 & w2837;
assign w2839 = shift_4 & ~w2683;
assign w2840 = ~shift_4 & ~w2121;
assign w2841 = ~w2839 & ~w2840;
assign w2842 = ~shift_6 & w2841;
assign w2843 = ~w2838 & ~w2842;
assign w2844 = ~shift_4 & ~w2188;
assign w2845 = shift_4 & ~w2690;
assign w2846 = ~w2844 & ~w2845;
assign w2847 = shift_6 & w2846;
assign w2848 = shift_4 & ~w2698;
assign w2849 = ~shift_4 & ~w2166;
assign w2850 = ~w2848 & ~w2849;
assign w2851 = ~shift_6 & w2850;
assign w2852 = ~w2847 & ~w2851;
assign w2853 = ~shift_4 & ~w2233;
assign w2854 = shift_4 & ~w2705;
assign w2855 = ~w2853 & ~w2854;
assign w2856 = shift_6 & w2855;
assign w2857 = shift_4 & ~w2713;
assign w2858 = ~shift_4 & ~w2211;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = ~shift_6 & w2859;
assign w2861 = ~w2856 & ~w2860;
assign w2862 = shift_6 & w378;
assign w2863 = ~shift_6 & w188;
assign w2864 = ~w2862 & ~w2863;
assign w2865 = shift_6 & w756;
assign w2866 = ~shift_6 & w566;
assign w2867 = ~w2865 & ~w2866;
assign w2868 = shift_6 & w1131;
assign w2869 = ~shift_6 & w941;
assign w2870 = ~w2868 & ~w2869;
assign w2871 = shift_6 & w1503;
assign w2872 = ~shift_6 & w1313;
assign w2873 = ~w2871 & ~w2872;
assign w2874 = shift_6 & w1572;
assign w2875 = ~shift_6 & w1538;
assign w2876 = ~w2874 & ~w2875;
assign w2877 = shift_6 & w1641;
assign w2878 = ~shift_6 & w1607;
assign w2879 = ~w2877 & ~w2878;
assign w2880 = shift_6 & w1710;
assign w2881 = ~shift_6 & w1676;
assign w2882 = ~w2880 & ~w2881;
assign w2883 = shift_6 & w1779;
assign w2884 = ~shift_6 & w1745;
assign w2885 = ~w2883 & ~w2884;
assign w2886 = shift_6 & w1848;
assign w2887 = ~shift_6 & w1814;
assign w2888 = ~w2886 & ~w2887;
assign w2889 = shift_6 & w1917;
assign w2890 = ~shift_6 & w1883;
assign w2891 = ~w2889 & ~w2890;
assign w2892 = shift_6 & w1986;
assign w2893 = ~shift_6 & w1952;
assign w2894 = ~w2892 & ~w2893;
assign w2895 = shift_6 & w2055;
assign w2896 = ~shift_6 & w2021;
assign w2897 = ~w2895 & ~w2896;
assign w2898 = shift_6 & w2100;
assign w2899 = ~shift_6 & w2078;
assign w2900 = ~w2898 & ~w2899;
assign w2901 = shift_6 & w2145;
assign w2902 = ~shift_6 & w2123;
assign w2903 = ~w2901 & ~w2902;
assign w2904 = shift_6 & w2190;
assign w2905 = ~shift_6 & w2168;
assign w2906 = ~w2904 & ~w2905;
assign w2907 = shift_6 & w2235;
assign w2908 = ~shift_6 & w2213;
assign w2909 = ~w2907 & ~w2908;
assign w2910 = shift_6 & w2250;
assign w2911 = ~shift_6 & w2243;
assign w2912 = ~w2910 & ~w2911;
assign w2913 = shift_6 & w2265;
assign w2914 = ~shift_6 & w2258;
assign w2915 = ~w2913 & ~w2914;
assign w2916 = shift_6 & w2280;
assign w2917 = ~shift_6 & w2273;
assign w2918 = ~w2916 & ~w2917;
assign w2919 = shift_6 & w2295;
assign w2920 = ~shift_6 & w2288;
assign w2921 = ~w2919 & ~w2920;
assign w2922 = shift_6 & w2310;
assign w2923 = ~shift_6 & w2303;
assign w2924 = ~w2922 & ~w2923;
assign w2925 = shift_6 & w2325;
assign w2926 = ~shift_6 & w2318;
assign w2927 = ~w2925 & ~w2926;
assign w2928 = shift_6 & w2340;
assign w2929 = ~shift_6 & w2333;
assign w2930 = ~w2928 & ~w2929;
assign w2931 = shift_6 & w2355;
assign w2932 = ~shift_6 & w2348;
assign w2933 = ~w2931 & ~w2932;
assign w2934 = shift_6 & w2370;
assign w2935 = ~shift_6 & w2363;
assign w2936 = ~w2934 & ~w2935;
assign w2937 = shift_6 & w2385;
assign w2938 = ~shift_6 & w2378;
assign w2939 = ~w2937 & ~w2938;
assign w2940 = shift_6 & w2400;
assign w2941 = ~shift_6 & w2393;
assign w2942 = ~w2940 & ~w2941;
assign w2943 = shift_6 & w2415;
assign w2944 = ~shift_6 & w2408;
assign w2945 = ~w2943 & ~w2944;
assign w2946 = shift_6 & w2430;
assign w2947 = ~shift_6 & w2423;
assign w2948 = ~w2946 & ~w2947;
assign w2949 = shift_6 & w2445;
assign w2950 = ~shift_6 & w2438;
assign w2951 = ~w2949 & ~w2950;
assign w2952 = shift_6 & w2460;
assign w2953 = ~shift_6 & w2453;
assign w2954 = ~w2952 & ~w2953;
assign w2955 = shift_6 & w2475;
assign w2956 = ~shift_6 & w2468;
assign w2957 = ~w2955 & ~w2956;
assign w2958 = shift_6 & w2490;
assign w2959 = ~shift_6 & w2483;
assign w2960 = ~w2958 & ~w2959;
assign w2961 = shift_6 & w2505;
assign w2962 = ~shift_6 & w2498;
assign w2963 = ~w2961 & ~w2962;
assign w2964 = shift_6 & w2520;
assign w2965 = ~shift_6 & w2513;
assign w2966 = ~w2964 & ~w2965;
assign w2967 = shift_6 & w2535;
assign w2968 = ~shift_6 & w2528;
assign w2969 = ~w2967 & ~w2968;
assign w2970 = shift_6 & w2550;
assign w2971 = ~shift_6 & w2543;
assign w2972 = ~w2970 & ~w2971;
assign w2973 = shift_6 & w2565;
assign w2974 = ~shift_6 & w2558;
assign w2975 = ~w2973 & ~w2974;
assign w2976 = shift_6 & w2580;
assign w2977 = ~shift_6 & w2573;
assign w2978 = ~w2976 & ~w2977;
assign w2979 = shift_6 & w2595;
assign w2980 = ~shift_6 & w2588;
assign w2981 = ~w2979 & ~w2980;
assign w2982 = shift_6 & w2610;
assign w2983 = ~shift_6 & w2603;
assign w2984 = ~w2982 & ~w2983;
assign w2985 = shift_6 & w2625;
assign w2986 = ~shift_6 & w2618;
assign w2987 = ~w2985 & ~w2986;
assign w2988 = shift_6 & w2640;
assign w2989 = ~shift_6 & w2633;
assign w2990 = ~w2988 & ~w2989;
assign w2991 = shift_6 & w2655;
assign w2992 = ~shift_6 & w2648;
assign w2993 = ~w2991 & ~w2992;
assign w2994 = shift_6 & w2670;
assign w2995 = ~shift_6 & w2663;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = shift_6 & w2685;
assign w2998 = ~shift_6 & w2678;
assign w2999 = ~w2997 & ~w2998;
assign w3000 = shift_6 & w2700;
assign w3001 = ~shift_6 & w2693;
assign w3002 = ~w3000 & ~w3001;
assign w3003 = shift_6 & w2715;
assign w3004 = ~shift_6 & w2708;
assign w3005 = ~w3003 & ~w3004;
assign w3006 = shift_6 & w2724;
assign w3007 = ~shift_6 & w2720;
assign w3008 = ~w3006 & ~w3007;
assign w3009 = shift_6 & w2733;
assign w3010 = ~shift_6 & w2729;
assign w3011 = ~w3009 & ~w3010;
assign w3012 = shift_6 & w2742;
assign w3013 = ~shift_6 & w2738;
assign w3014 = ~w3012 & ~w3013;
assign w3015 = shift_6 & w2751;
assign w3016 = ~shift_6 & w2747;
assign w3017 = ~w3015 & ~w3016;
assign w3018 = shift_6 & w2760;
assign w3019 = ~shift_6 & w2756;
assign w3020 = ~w3018 & ~w3019;
assign w3021 = shift_6 & w2769;
assign w3022 = ~shift_6 & w2765;
assign w3023 = ~w3021 & ~w3022;
assign w3024 = shift_6 & w2778;
assign w3025 = ~shift_6 & w2774;
assign w3026 = ~w3024 & ~w3025;
assign w3027 = shift_6 & w2787;
assign w3028 = ~shift_6 & w2783;
assign w3029 = ~w3027 & ~w3028;
assign w3030 = shift_6 & w2796;
assign w3031 = ~shift_6 & w2792;
assign w3032 = ~w3030 & ~w3031;
assign w3033 = shift_6 & w2805;
assign w3034 = ~shift_6 & w2801;
assign w3035 = ~w3033 & ~w3034;
assign w3036 = shift_6 & w2814;
assign w3037 = ~shift_6 & w2810;
assign w3038 = ~w3036 & ~w3037;
assign w3039 = shift_6 & w2823;
assign w3040 = ~shift_6 & w2819;
assign w3041 = ~w3039 & ~w3040;
assign w3042 = shift_6 & w2832;
assign w3043 = ~shift_6 & w2828;
assign w3044 = ~w3042 & ~w3043;
assign w3045 = shift_6 & w2841;
assign w3046 = ~shift_6 & w2837;
assign w3047 = ~w3045 & ~w3046;
assign w3048 = shift_6 & w2850;
assign w3049 = ~shift_6 & w2846;
assign w3050 = ~w3048 & ~w3049;
assign w3051 = shift_6 & w2859;
assign w3052 = ~shift_6 & w2855;
assign w3053 = ~w3051 & ~w3052;
assign one = 1;
assign result_0 = ~w380;
assign result_1 = ~w758;
assign result_2 = ~w1133;
assign result_3 = ~w1505;
assign result_4 = ~w1574;
assign result_5 = ~w1643;
assign result_6 = ~w1712;
assign result_7 = ~w1781;
assign result_8 = ~w1850;
assign result_9 = ~w1919;
assign result_10 = ~w1988;
assign result_11 = ~w2057;
assign result_12 = ~w2102;
assign result_13 = ~w2147;
assign result_14 = ~w2192;
assign result_15 = ~w2237;
assign result_16 = ~w2252;
assign result_17 = ~w2267;
assign result_18 = ~w2282;
assign result_19 = ~w2297;
assign result_20 = ~w2312;
assign result_21 = ~w2327;
assign result_22 = ~w2342;
assign result_23 = ~w2357;
assign result_24 = ~w2372;
assign result_25 = ~w2387;
assign result_26 = ~w2402;
assign result_27 = ~w2417;
assign result_28 = ~w2432;
assign result_29 = ~w2447;
assign result_30 = ~w2462;
assign result_31 = ~w2477;
assign result_32 = ~w2492;
assign result_33 = ~w2507;
assign result_34 = ~w2522;
assign result_35 = ~w2537;
assign result_36 = ~w2552;
assign result_37 = ~w2567;
assign result_38 = ~w2582;
assign result_39 = ~w2597;
assign result_40 = ~w2612;
assign result_41 = ~w2627;
assign result_42 = ~w2642;
assign result_43 = ~w2657;
assign result_44 = ~w2672;
assign result_45 = ~w2687;
assign result_46 = ~w2702;
assign result_47 = ~w2717;
assign result_48 = ~w2726;
assign result_49 = ~w2735;
assign result_50 = ~w2744;
assign result_51 = ~w2753;
assign result_52 = ~w2762;
assign result_53 = ~w2771;
assign result_54 = ~w2780;
assign result_55 = ~w2789;
assign result_56 = ~w2798;
assign result_57 = ~w2807;
assign result_58 = ~w2816;
assign result_59 = ~w2825;
assign result_60 = ~w2834;
assign result_61 = ~w2843;
assign result_62 = ~w2852;
assign result_63 = ~w2861;
assign result_64 = ~w2864;
assign result_65 = ~w2867;
assign result_66 = ~w2870;
assign result_67 = ~w2873;
assign result_68 = ~w2876;
assign result_69 = ~w2879;
assign result_70 = ~w2882;
assign result_71 = ~w2885;
assign result_72 = ~w2888;
assign result_73 = ~w2891;
assign result_74 = ~w2894;
assign result_75 = ~w2897;
assign result_76 = ~w2900;
assign result_77 = ~w2903;
assign result_78 = ~w2906;
assign result_79 = ~w2909;
assign result_80 = ~w2912;
assign result_81 = ~w2915;
assign result_82 = ~w2918;
assign result_83 = ~w2921;
assign result_84 = ~w2924;
assign result_85 = ~w2927;
assign result_86 = ~w2930;
assign result_87 = ~w2933;
assign result_88 = ~w2936;
assign result_89 = ~w2939;
assign result_90 = ~w2942;
assign result_91 = ~w2945;
assign result_92 = ~w2948;
assign result_93 = ~w2951;
assign result_94 = ~w2954;
assign result_95 = ~w2957;
assign result_96 = ~w2960;
assign result_97 = ~w2963;
assign result_98 = ~w2966;
assign result_99 = ~w2969;
assign result_100 = ~w2972;
assign result_101 = ~w2975;
assign result_102 = ~w2978;
assign result_103 = ~w2981;
assign result_104 = ~w2984;
assign result_105 = ~w2987;
assign result_106 = ~w2990;
assign result_107 = ~w2993;
assign result_108 = ~w2996;
assign result_109 = ~w2999;
assign result_110 = ~w3002;
assign result_111 = ~w3005;
assign result_112 = ~w3008;
assign result_113 = ~w3011;
assign result_114 = ~w3014;
assign result_115 = ~w3017;
assign result_116 = ~w3020;
assign result_117 = ~w3023;
assign result_118 = ~w3026;
assign result_119 = ~w3029;
assign result_120 = ~w3032;
assign result_121 = ~w3035;
assign result_122 = ~w3038;
assign result_123 = ~w3041;
assign result_124 = ~w3044;
assign result_125 = ~w3047;
assign result_126 = ~w3050;
assign result_127 = ~w3053;
endmodule

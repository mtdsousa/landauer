module mem_ctrl_best_speed (
        pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, 
        po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361;
assign w0 = ~pi0039 & ~pi0087;
assign w1 = ~pi0092 & w0;
assign w2 = ~pi0038 & ~pi0054;
assign w3 = ~pi0074 & ~pi0075;
assign w4 = w2 & w3;
assign w5 = ~pi0100 & w4;
assign w6 = w1 & w5;
assign w7 = pi0095 & ~pi0479;
assign w8 = pi0234 & w7;
assign w9 = pi0105 & pi0228;
assign w10 = ~pi0215 & ~pi0216;
assign w11 = ~pi0221 & pi0299;
assign w12 = w10 & w11;
assign w13 = w9 & w12;
assign w14 = ~pi0222 & ~pi0223;
assign w15 = ~pi0224 & ~pi0299;
assign w16 = w14 & w15;
assign w17 = ~w8 & w16;
assign w18 = (~w8 & w13) | (~w8 & w17) | (w13 & w17);
assign w19 = ~pi0216 & pi0833;
assign w20 = ~pi0215 & ~pi0221;
assign w21 = (~pi0215 & w19) | (~pi0215 & w20) | (w19 & w20);
assign w22 = ~pi0221 & pi0265;
assign w23 = pi0221 & pi0929;
assign w24 = ~pi0216 & ~w23;
assign w25 = ~w22 & ~w24;
assign w26 = w21 & ~w25;
assign w27 = ~pi1144 & ~w21;
assign w28 = pi0299 & w27;
assign w29 = (pi0299 & w26) | (pi0299 & w28) | (w26 & w28);
assign w30 = ~pi0153 & ~pi0215;
assign w31 = (~pi0215 & w9) | (~pi0215 & w30) | (w9 & w30);
assign w32 = ~pi0216 & ~pi0221;
assign w33 = w31 & w32;
assign w34 = ~w18 & w33;
assign w35 = (~w18 & ~w29) | (~w18 & w34) | (~w29 & w34);
assign w36 = ~pi0161 & ~pi0166;
assign w37 = ~pi0146 & pi0152;
assign w38 = (~pi0146 & ~w36) | (~pi0146 & w37) | (~w36 & w37);
assign w39 = pi0100 & pi0252;
assign w40 = ~w38 & w39;
assign w41 = ~pi0228 & w4;
assign w42 = ~w40 & w41;
assign w43 = pi0092 & ~pi0100;
assign w44 = ~pi0092 & pi0100;
assign w45 = ~w43 & ~w44;
assign w46 = ~pi0087 & ~w45;
assign w47 = pi0039 & ~pi0087;
assign w48 = ~pi0092 & ~pi0100;
assign w49 = w47 & w48;
assign w50 = pi0039 & ~w49;
assign w51 = ~pi0039 & pi0087;
assign w52 = w48 & w51;
assign w53 = ~w49 & ~w52;
assign w54 = (~w46 & w50) | (~w46 & w53) | (w50 & w53);
assign w55 = w42 & ~w54;
assign w56 = ~w13 & ~w16;
assign w57 = ~pi0036 & ~pi0045;
assign w58 = ~pi0049 & ~pi0089;
assign w59 = w57 & w58;
assign w60 = ~pi0104 & w59;
assign w61 = ~pi0048 & ~pi0061;
assign w62 = ~pi0076 & ~pi0085;
assign w63 = w61 & w62;
assign w64 = ~pi0106 & w63;
assign w65 = w60 & w64;
assign w66 = ~pi0081 & ~pi0088;
assign w67 = ~pi0098 & w66;
assign w68 = ~pi0066 & ~pi0069;
assign w69 = ~pi0082 & ~pi0083;
assign w70 = w68 & w69;
assign w71 = ~pi0103 & ~pi0111;
assign w72 = w70 & w71;
assign w73 = w67 & w72;
assign w74 = w65 & w73;
assign w75 = ~pi0063 & ~pi0064;
assign w76 = ~pi0065 & ~pi0102;
assign w77 = w75 & w76;
assign w78 = ~pi0107 & w77;
assign w79 = ~pi0067 & ~pi0068;
assign w80 = ~pi0071 & ~pi0073;
assign w81 = w79 & w80;
assign w82 = ~pi0084 & w81;
assign w83 = w78 & w82;
assign w84 = w56 & ~w83;
assign w85 = (w56 & ~w74) | (w56 & w84) | (~w74 & w84);
assign w86 = w55 & ~w85;
assign w87 = ~pi0046 & ~pi0047;
assign w88 = ~pi0058 & ~pi0091;
assign w89 = w87 & w88;
assign w90 = ~pi0109 & ~pi0110;
assign w91 = w89 & w90;
assign w92 = ~pi0050 & ~pi0053;
assign w93 = ~pi0060 & ~pi0077;
assign w94 = w92 & w93;
assign w95 = ~pi0097 & ~pi0108;
assign w96 = ~pi0086 & ~pi0094;
assign w97 = w95 & w96;
assign w98 = w94 & w97;
assign w99 = w91 & w98;
assign w100 = ~pi0032 & ~pi0035;
assign w101 = ~pi0040 & ~pi0090;
assign w102 = w100 & w101;
assign w103 = ~pi0093 & ~pi0095;
assign w104 = w102 & w103;
assign w105 = ~pi0072 & ~pi0096;
assign w106 = ~pi0051 & ~pi0070;
assign w107 = w105 & w106;
assign w108 = w104 & w107;
assign w109 = w99 & w108;
assign w110 = w35 & ~w109;
assign w111 = (w35 & ~w86) | (w35 & w110) | (~w86 & w110);
assign w112 = w74 & w83;
assign w113 = w109 & w112;
assign w114 = ~pi0221 & w10;
assign w115 = w55 & w114;
assign w116 = w113 & w115;
assign w117 = ~pi0038 & ~pi0039;
assign w118 = ~pi0087 & w117;
assign w119 = w113 & w118;
assign w120 = w29 & ~w33;
assign w121 = w118 & ~w120;
assign w122 = w113 & w121;
assign w123 = (w116 & w119) | (w116 & w122) | (w119 & w122);
assign w124 = ~pi0210 & ~w38;
assign w125 = ~pi0137 & ~w124;
assign w126 = w29 & w125;
assign w127 = ~pi0174 & ~pi0189;
assign w128 = ~pi0142 & pi0144;
assign w129 = (~pi0142 & ~w127) | (~pi0142 & w128) | (~w127 & w128);
assign w130 = ~pi0137 & pi0198;
assign w131 = (~pi0137 & w129) | (~pi0137 & w130) | (w129 & w130);
assign w132 = w16 & w131;
assign w133 = pi0075 & ~pi0100;
assign w134 = ~pi0075 & pi0100;
assign w135 = ~w133 & ~w134;
assign w136 = ~pi0074 & ~pi0092;
assign w137 = ~pi0054 & w136;
assign w138 = ~w135 & w137;
assign w139 = ~w132 & w138;
assign w140 = ~pi0074 & pi0092;
assign w141 = pi0074 & ~pi0092;
assign w142 = ~w140 & ~w141;
assign w143 = ~pi0054 & ~w142;
assign w144 = pi0054 & w136;
assign w145 = pi0137 & w144;
assign w146 = (pi0137 & w143) | (pi0137 & w145) | (w143 & w145);
assign w147 = ~pi0075 & ~pi0100;
assign w148 = w146 & w147;
assign w149 = ~w139 & ~w148;
assign w150 = ~w126 & ~w149;
assign w151 = ~w111 & ~w150;
assign w152 = (~w111 & ~w123) | (~w111 & w151) | (~w123 & w151);
assign w153 = ~w16 & ~w29;
assign w154 = ~pi0105 & pi0228;
assign w155 = w114 & ~w154;
assign w156 = pi0137 & w155;
assign w157 = (pi0137 & ~w29) | (pi0137 & w156) | (~w29 & w156);
assign w158 = ~w153 & ~w157;
assign w159 = pi0087 & ~pi0092;
assign w160 = ~pi0087 & pi0092;
assign w161 = ~w159 & ~w160;
assign w162 = ~pi0039 & ~w161;
assign w163 = w5 & w162;
assign w164 = pi0039 & ~w5;
assign w165 = ~pi0039 & w33;
assign w166 = ~w5 & ~w165;
assign w167 = (w29 & w164) | (w29 & w166) | (w164 & w166);
assign w168 = ~pi0054 & ~pi0074;
assign w169 = ~pi0075 & ~pi0087;
assign w170 = w168 & w169;
assign w171 = w48 & w170;
assign w172 = ~w163 & ~w171;
assign w173 = (~w163 & w167) | (~w163 & w172) | (w167 & w172);
assign w174 = ~w158 & ~w173;
assign w175 = w113 & w174;
assign w176 = ~w6 & w175;
assign w177 = (~w6 & ~w152) | (~w6 & w176) | (~w152 & w176);
assign w178 = ~pi0055 & ~pi0056;
assign w179 = ~pi0057 & ~pi0059;
assign w180 = w178 & w179;
assign w181 = ~pi0062 & ~pi0332;
assign w182 = w180 & w181;
assign w183 = ~w177 & w182;
assign w184 = ~pi0035 & ~pi0051;
assign w185 = ~pi0070 & ~pi0090;
assign w186 = w184 & w185;
assign w187 = ~pi0093 & w105;
assign w188 = w186 & w187;
assign w189 = w95 & w188;
assign w190 = w94 & w96;
assign w191 = w91 & w190;
assign w192 = w189 & w191;
assign w193 = w67 & w78;
assign w194 = w192 & w193;
assign w195 = w72 & w82;
assign w196 = w65 & w195;
assign w197 = ~pi0040 & ~pi0095;
assign w198 = pi0032 & w197;
assign w199 = pi0040 & ~pi0095;
assign w200 = ~pi0040 & pi0095;
assign w201 = ~w199 & ~w200;
assign w202 = ~pi0032 & ~w201;
assign w203 = ~w198 & ~w202;
assign w204 = w196 & w203;
assign w205 = w194 & w204;
assign w206 = ~pi0228 & ~w205;
assign w207 = pi0102 & ~pi0107;
assign w208 = ~pi0102 & pi0107;
assign w209 = ~w207 & ~w208;
assign w210 = ~pi0098 & ~w209;
assign w211 = ~pi0102 & ~pi0107;
assign w212 = ~pi0088 & pi0098;
assign w213 = w211 & w212;
assign w214 = (~pi0088 & w210) | (~pi0088 & w213) | (w210 & w213);
assign w215 = ~pi0098 & w211;
assign w216 = pi0081 & ~pi0088;
assign w217 = pi0081 & ~w216;
assign w218 = (pi0081 & ~w215) | (pi0081 & w217) | (~w215 & w217);
assign w219 = w215 & w216;
assign w220 = pi0088 & ~pi0098;
assign w221 = w211 & w220;
assign w222 = ~pi0081 & w221;
assign w223 = ~w219 & ~w222;
assign w224 = (~w214 & w218) | (~w214 & w223) | (w218 & w223);
assign w225 = ~pi0065 & w75;
assign w226 = ~w224 & w225;
assign w227 = pi0064 & pi0065;
assign w228 = ~pi0063 & ~w227;
assign w229 = ~pi0064 & ~pi0065;
assign w230 = ~pi0102 & w229;
assign w231 = (~pi0102 & w228) | (~pi0102 & w230) | (w228 & w230);
assign w232 = w67 & w231;
assign w233 = w224 & w232;
assign w234 = ~w226 & ~w233;
assign w235 = pi0060 & pi0077;
assign w236 = ~pi0053 & ~w235;
assign w237 = ~pi0050 & w93;
assign w238 = (~pi0050 & w236) | (~pi0050 & w237) | (w236 & w237);
assign w239 = ~pi0046 & ~pi0109;
assign w240 = ~pi0053 & ~pi0109;
assign w241 = w93 & w240;
assign w242 = ~pi0046 & w241;
assign w243 = (w238 & w239) | (w238 & w242) | (w239 & w242);
assign w244 = w196 & w243;
assign w245 = pi0097 & pi0108;
assign w246 = w96 & ~w245;
assign w247 = ~w95 & ~w246;
assign w248 = ~w94 & ~w97;
assign w249 = (~w97 & w247) | (~w97 & w248) | (w247 & w248);
assign w250 = w193 & ~w249;
assign w251 = w244 & w250;
assign w252 = ~w98 & ~w250;
assign w253 = w244 & ~w252;
assign w254 = (~w234 & w251) | (~w234 & w253) | (w251 & w253);
assign w255 = pi0048 & pi0076;
assign w256 = ~pi0085 & ~pi0106;
assign w257 = ~w255 & w256;
assign w258 = ~pi0061 & w257;
assign w259 = pi0085 & ~pi0106;
assign w260 = ~pi0085 & pi0106;
assign w261 = ~w259 & ~w260;
assign w262 = ~pi0061 & ~w261;
assign w263 = pi0061 & ~pi0076;
assign w264 = w256 & w263;
assign w265 = (~pi0076 & w262) | (~pi0076 & w264) | (w262 & w264);
assign w266 = pi0048 & pi0061;
assign w267 = (pi0048 & ~w257) | (pi0048 & w266) | (~w257 & w266);
assign w268 = (~w258 & ~w265) | (~w258 & w267) | (~w265 & w267);
assign w269 = pi0089 & pi0104;
assign w270 = ~pi0049 & ~w269;
assign w271 = ~pi0089 & ~pi0104;
assign w272 = ~w270 & ~w271;
assign w273 = w64 & ~w272;
assign w274 = ~pi0049 & w271;
assign w275 = ~w273 & ~w274;
assign w276 = ~w268 & ~w275;
assign w277 = ~pi0066 & ~pi0068;
assign w278 = ~pi0073 & ~pi0084;
assign w279 = w277 & w278;
assign w280 = ~pi0048 & ~pi0049;
assign w281 = ~pi0076 & ~pi0089;
assign w282 = w280 & w281;
assign w283 = ~pi0061 & ~pi0104;
assign w284 = w256 & w283;
assign w285 = w282 & w284;
assign w286 = ~pi0045 & w279;
assign w287 = (w279 & w285) | (w279 & w286) | (w285 & w286);
assign w288 = w276 & w287;
assign w289 = pi0073 & ~pi0084;
assign w290 = ~pi0073 & pi0084;
assign w291 = ~w289 & ~w290;
assign w292 = ~pi0068 & ~w291;
assign w293 = ~pi0066 & pi0068;
assign w294 = w278 & w293;
assign w295 = (~pi0066 & w292) | (~pi0066 & w294) | (w292 & w294);
assign w296 = ~pi0045 & ~pi0049;
assign w297 = w271 & w296;
assign w298 = w64 & w297;
assign w299 = pi0066 & ~pi0068;
assign w300 = w278 & w299;
assign w301 = w297 & w300;
assign w302 = w64 & w301;
assign w303 = (w295 & w298) | (w295 & w302) | (w298 & w302);
assign w304 = ~pi0048 & ~pi0076;
assign w305 = ~pi0048 & w264;
assign w306 = (w262 & w304) | (w262 & w305) | (w304 & w305);
assign w307 = ~w275 & w306;
assign w308 = w258 & ~w287;
assign w309 = w303 & w308;
assign w310 = (w303 & w307) | (w303 & w309) | (w307 & w309);
assign w311 = ~w288 & ~w310;
assign w312 = w98 & w193;
assign w313 = w243 & w312;
assign w314 = ~w311 & w313;
assign w315 = pi0083 & ~pi0103;
assign w316 = ~pi0083 & pi0103;
assign w317 = ~w315 & ~w316;
assign w318 = ~pi0069 & ~w317;
assign w319 = ~pi0083 & ~pi0103;
assign w320 = pi0069 & ~pi0071;
assign w321 = w319 & w320;
assign w322 = (~pi0071 & w318) | (~pi0071 & w321) | (w318 & w321);
assign w323 = w279 & w297;
assign w324 = w64 & w323;
assign w325 = ~pi0036 & ~pi0067;
assign w326 = ~pi0082 & ~pi0111;
assign w327 = w325 & w326;
assign w328 = w324 & w327;
assign w329 = w322 & w328;
assign w330 = pi0071 & ~w327;
assign w331 = (pi0071 & ~w324) | (pi0071 & w330) | (~w324 & w330);
assign w332 = ~w324 & ~w327;
assign w333 = ~pi0069 & ~pi0083;
assign w334 = ~pi0103 & w333;
assign w335 = pi0082 & pi0111;
assign w336 = ~pi0067 & ~w335;
assign w337 = ~pi0036 & w326;
assign w338 = (~pi0036 & w336) | (~pi0036 & w337) | (w336 & w337);
assign w339 = ~pi0067 & w326;
assign w340 = w334 & w339;
assign w341 = (w334 & w338) | (w334 & w340) | (w338 & w340);
assign w342 = ~w332 & w341;
assign w343 = ~w331 & w342;
assign w344 = ~w329 & ~w343;
assign w345 = ~w254 & w344;
assign w346 = (~w254 & ~w314) | (~w254 & w345) | (~w314 & w345);
assign w347 = ~pi0032 & ~pi0040;
assign w348 = ~pi0095 & w347;
assign w349 = w107 & w348;
assign w350 = pi0086 & pi0094;
assign w351 = ~pi0047 & ~pi0058;
assign w352 = ~pi0090 & ~pi0091;
assign w353 = w351 & w352;
assign w354 = ~pi0093 & ~pi0110;
assign w355 = ~pi0035 & ~pi0093;
assign w356 = w354 & w355;
assign w357 = w353 & w356;
assign w358 = ~w350 & w357;
assign w359 = w98 & w355;
assign w360 = (~w350 & w358) | (~w350 & w359) | (w358 & w359);
assign w361 = w358 & w360;
assign w362 = pi0091 & pi0110;
assign w363 = ~pi0090 & ~w362;
assign w364 = ~pi0091 & ~pi0110;
assign w365 = ~pi0058 & w364;
assign w366 = (~pi0058 & w363) | (~pi0058 & w365) | (w363 & w365);
assign w367 = ~pi0058 & ~pi0090;
assign w368 = w364 & w367;
assign w369 = pi0047 & ~w368;
assign w370 = ~pi0047 & ~pi0090;
assign w371 = w364 & w370;
assign w372 = ~w368 & ~w371;
assign w373 = (~w366 & w369) | (~w366 & w372) | (w369 & w372);
assign w374 = w243 & ~w373;
assign w375 = (w358 & w360) | (w358 & w374) | (w360 & w374);
assign w376 = (w112 & w361) | (w112 & w375) | (w361 & w375);
assign w377 = w349 & w376;
assign w378 = ~w346 & w377;
assign w379 = ~pi0046 & w354;
assign w380 = w353 & w379;
assign w381 = ~w374 & w380;
assign w382 = w353 & w354;
assign w383 = w374 & ~w382;
assign w384 = ~w381 & ~w383;
assign w385 = w83 & w359;
assign w386 = w74 & w385;
assign w387 = ~w384 & w386;
assign w388 = ~pi0070 & w105;
assign w389 = pi0072 & pi0096;
assign w390 = ~pi0070 & ~w389;
assign w391 = ~pi0051 & w105;
assign w392 = (~pi0051 & w390) | (~pi0051 & w391) | (w390 & w391);
assign w393 = ~w388 & ~w392;
assign w394 = ~w104 & ~w188;
assign w395 = (~w188 & w393) | (~w188 & w394) | (w393 & w394);
assign w396 = w99 & ~w395;
assign w397 = w112 & w396;
assign w398 = ~w349 & ~w397;
assign w399 = pi0035 & ~pi0093;
assign w400 = ~pi0035 & pi0093;
assign w401 = ~w399 & ~w400;
assign w402 = ~pi0090 & ~w401;
assign w403 = w349 & w402;
assign w404 = w99 & w403;
assign w405 = w112 & w404;
assign w406 = ~w397 & ~w405;
assign w407 = (~w387 & w398) | (~w387 & w406) | (w398 & w406);
assign w408 = w206 & ~w407;
assign w409 = (w206 & w378) | (w206 & w408) | (w378 & w408);
assign w410 = ~w205 & w397;
assign w411 = pi0210 & pi0299;
assign w412 = pi0198 & ~pi0299;
assign w413 = ~w411 & ~w412;
assign w414 = pi0032 & pi0225;
assign w415 = pi0225 & pi0841;
assign w416 = pi0032 & w415;
assign w417 = (~w413 & w414) | (~w413 & w416) | (w414 & w416);
assign w418 = pi0070 & pi0332;
assign w419 = ~w417 & ~w418;
assign w420 = w410 & ~w419;
assign w421 = ~w153 & ~w420;
assign w422 = w9 & w29;
assign w423 = ~w16 & ~w422;
assign w424 = ~w420 & ~w423;
assign w425 = (w409 & w421) | (w409 & w424) | (w421 & w424);
assign w426 = ~pi0070 & ~pi0072;
assign w427 = w184 & w426;
assign w428 = ~pi0090 & ~pi0093;
assign w429 = w427 & w428;
assign w430 = w348 & w429;
assign w431 = w99 & w430;
assign w432 = pi0096 & w431;
assign w433 = w112 & w432;
assign w434 = (pi0234 & w8) | (pi0234 & w433) | (w8 & w433);
assign w435 = ~w7 & ~w433;
assign w436 = w104 & ~w393;
assign w437 = w188 & ~w203;
assign w438 = ~w436 & ~w437;
assign w439 = w112 & ~w438;
assign w440 = ~w99 & ~w349;
assign w441 = (~w349 & ~w439) | (~w349 & w440) | (~w439 & w440);
assign w442 = w435 & ~w441;
assign w443 = ~pi0053 & ~pi0060;
assign w444 = ~pi0035 & ~pi0137;
assign w445 = w443 & w444;
assign w446 = pi0299 & ~w38;
assign w447 = ~pi0299 & ~w129;
assign w448 = ~w446 & ~w447;
assign w449 = ~pi0833 & pi0957;
assign w450 = ~pi1091 & pi1093;
assign w451 = (pi1093 & w449) | (pi1093 & w450) | (w449 & w450);
assign w452 = pi0829 & pi0950;
assign w453 = pi1092 & w452;
assign w454 = ~w451 & w453;
assign w455 = w413 & w454;
assign w456 = ~w448 & w455;
assign w457 = pi0097 & pi1093;
assign w458 = pi0096 & ~pi0841;
assign w459 = ~w457 & ~w458;
assign w460 = w445 & w459;
assign w461 = (w445 & ~w456) | (w445 & w460) | (~w456 & w460);
assign w462 = ~w434 & w461;
assign w463 = (~w434 & ~w442) | (~w434 & w462) | (~w442 & w462);
assign w464 = w83 & w98;
assign w465 = w74 & w464;
assign w466 = pi0046 & ~pi0047;
assign w467 = w90 & w466;
assign w468 = w367 & ~w467;
assign w469 = pi0109 & ~pi0110;
assign w470 = ~pi0109 & pi0110;
assign w471 = ~w469 & ~w470;
assign w472 = ~pi0047 & ~w471;
assign w473 = ~pi0046 & pi0047;
assign w474 = w90 & w473;
assign w475 = (~pi0046 & w472) | (~pi0046 & w474) | (w472 & w474);
assign w476 = w468 & ~w475;
assign w477 = w465 & ~w476;
assign w478 = ~w254 & w313;
assign w479 = w67 & w95;
assign w480 = w78 & w479;
assign w481 = ~pi0094 & w480;
assign w482 = w254 & ~w481;
assign w483 = ~w478 & ~w482;
assign w484 = ~w311 & ~w344;
assign w485 = ~w477 & ~w484;
assign w486 = (~w477 & w483) | (~w477 & w485) | (w483 & w485);
assign w487 = ~w98 & w254;
assign w488 = w376 & w387;
assign w489 = (w376 & w487) | (w376 & w488) | (w487 & w488);
assign w490 = (w376 & ~w486) | (w376 & w489) | (~w486 & w489);
assign w491 = w83 & w99;
assign w492 = w74 & w491;
assign w493 = w105 & w355;
assign w494 = ~pi0040 & ~pi0051;
assign w495 = w493 & w494;
assign w496 = ~pi0093 & pi0225;
assign w497 = pi0035 & ~w496;
assign w498 = ~w495 & ~w497;
assign w499 = ~pi0090 & w498;
assign w500 = ~pi0095 & ~w499;
assign w501 = (~pi0095 & ~w492) | (~pi0095 & w500) | (~w492 & w500);
assign w502 = ~w463 & ~w501;
assign w503 = (~w463 & w490) | (~w463 & w502) | (w490 & w502);
assign w504 = w425 & ~w503;
assign w505 = ~pi0221 & ~pi0228;
assign w506 = w10 & w505;
assign w507 = ~w407 & w506;
assign w508 = (w378 & w506) | (w378 & w507) | (w506 & w507);
assign w509 = w6 & ~w120;
assign w510 = w120 & w205;
assign w511 = w6 & ~w510;
assign w512 = (w508 & w509) | (w508 & w511) | (w509 & w511);
assign w513 = w183 & ~w512;
assign w514 = (w183 & w504) | (w183 & w513) | (w504 & w513);
assign w515 = ~pi0224 & pi0833;
assign w516 = (~pi0223 & w14) | (~pi0223 & w515) | (w14 & w515);
assign w517 = ~pi0299 & ~w516;
assign w518 = ~pi0224 & pi0929;
assign w519 = pi0224 & pi0265;
assign w520 = ~pi0222 & ~w519;
assign w521 = ~w518 & ~w520;
assign w522 = ~w517 & ~w521;
assign w523 = ~pi0299 & pi1144;
assign w524 = ~w516 & w523;
assign w525 = ~pi0062 & ~pi0299;
assign w526 = w180 & w525;
assign w527 = ~w524 & w526;
assign w528 = ~w522 & w527;
assign w529 = ~pi0062 & w180;
assign w530 = w27 & ~w529;
assign w531 = (w26 & ~w529) | (w26 & w530) | (~w529 & w530);
assign w532 = ~pi0063 & ~pi0107;
assign w533 = ~pi0100 & w532;
assign w534 = w4 & w533;
assign w535 = w1 & w179;
assign w536 = w534 & w535;
assign w537 = pi0056 & ~pi0062;
assign w538 = ~pi0056 & pi0062;
assign w539 = ~w537 & ~w538;
assign w540 = ~pi0040 & ~pi0055;
assign w541 = ~w539 & w540;
assign w542 = w536 & w541;
assign w543 = w109 & ~w542;
assign w544 = pi0056 & pi0062;
assign w545 = ~pi0055 & ~w544;
assign w546 = ~pi0056 & ~pi0062;
assign w547 = w179 & w546;
assign w548 = (w179 & w545) | (w179 & w547) | (w545 & w547);
assign w549 = w1 & w548;
assign w550 = w5 & w549;
assign w551 = w112 & w550;
assign w552 = w543 & w551;
assign w553 = w109 & w550;
assign w554 = w112 & w553;
assign w555 = pi0234 & w9;
assign w556 = w7 & w555;
assign w557 = ~pi0153 & ~w9;
assign w558 = ~w556 & ~w557;
assign w559 = ~w554 & ~w558;
assign w560 = ~w552 & ~w559;
assign w561 = pi0153 & pi0228;
assign w562 = ~pi0105 & w561;
assign w563 = w114 & ~w562;
assign w564 = w531 & ~w563;
assign w565 = (w531 & w560) | (w531 & w564) | (w560 & w564);
assign w566 = w6 & w109;
assign w567 = w112 & w566;
assign w568 = w1 & w114;
assign w569 = w5 & w568;
assign w570 = w542 & w569;
assign w571 = pi0057 & ~pi0059;
assign w572 = ~pi0057 & pi0059;
assign w573 = ~w571 & ~w572;
assign w574 = ~pi0055 & ~w573;
assign w575 = pi0055 & w179;
assign w576 = w546 & w575;
assign w577 = (w546 & w574) | (w546 & w576) | (w574 & w576);
assign w578 = ~w542 & ~w577;
assign w579 = w569 & ~w578;
assign w580 = (w567 & w570) | (w567 & w579) | (w570 & w579);
assign w581 = ~pi0228 & w179;
assign w582 = pi0137 & w9;
assign w583 = (pi0137 & w581) | (pi0137 & w582) | (w581 & w582);
assign w584 = pi0137 & ~pi0153;
assign w585 = (~pi0153 & w154) | (~pi0153 & w584) | (w154 & w584);
assign w586 = ~w583 & ~w585;
assign w587 = w113 & ~w586;
assign w588 = w580 & w587;
assign w589 = ~w528 & w588;
assign w590 = (~w528 & ~w565) | (~w528 & w589) | (~w565 & w589);
assign w591 = ~pi0332 & ~w590;
assign w592 = ~w514 & ~w591;
assign w593 = w6 & w529;
assign w594 = ~w205 & w593;
assign w595 = w205 & ~w593;
assign w596 = w377 & w595;
assign w597 = ~w594 & ~w596;
assign w598 = (w346 & ~w594) | (w346 & w597) | (~w594 & w597);
assign w599 = ~w407 & ~w598;
assign w600 = w377 & w594;
assign w601 = ~w346 & w600;
assign w602 = w550 & w601;
assign w603 = (w550 & w599) | (w550 & w602) | (w599 & w602);
assign w604 = pi0239 & w9;
assign w605 = w7 & w604;
assign w606 = ~pi0154 & ~w9;
assign w607 = w114 & w606;
assign w608 = (w114 & w605) | (w114 & w607) | (w605 & w607);
assign w609 = pi0221 & pi0833;
assign w610 = w10 & w609;
assign w611 = pi0939 & w610;
assign w612 = ~pi0215 & pi0216;
assign w613 = ~pi0221 & pi0276;
assign w614 = w612 & w613;
assign w615 = ~w611 & ~w614;
assign w616 = pi1146 & ~w21;
assign w617 = w615 & ~w616;
assign w618 = ~w608 & w617;
assign w619 = ~w506 & ~w526;
assign w620 = ~w618 & w619;
assign w621 = w55 & w109;
assign w622 = w112 & w621;
assign w623 = ~w526 & ~w529;
assign w624 = (~w526 & ~w622) | (~w526 & w623) | (~w622 & w623);
assign w625 = ~w619 & ~w624;
assign w626 = ~w618 & ~w625;
assign w627 = (~w603 & w620) | (~w603 & w626) | (w620 & w626);
assign w628 = w7 & w16;
assign w629 = (w7 & w13) | (w7 & w628) | (w13 & w628);
assign w630 = ~w1 & ~w7;
assign w631 = (~w5 & ~w7) | (~w5 & w630) | (~w7 & w630);
assign w632 = ~w56 & ~w631;
assign w633 = (w433 & w629) | (w433 & w632) | (w629 & w632);
assign w634 = w1 & w506;
assign w635 = w5 & w634;
assign w636 = pi0299 & w635;
assign w637 = ~w395 & w636;
assign w638 = w7 & w347;
assign w639 = ~pi0096 & ~w638;
assign w640 = w637 & ~w639;
assign w641 = w492 & w640;
assign w642 = ~w633 & ~w641;
assign w643 = pi0222 & ~pi0223;
assign w644 = w15 & w643;
assign w645 = pi0833 & pi0939;
assign w646 = w644 & w645;
assign w647 = pi0224 & ~pi0299;
assign w648 = w14 & w647;
assign w649 = pi0276 & w648;
assign w650 = ~w646 & ~w649;
assign w651 = ~pi0299 & pi1146;
assign w652 = ~w516 & w651;
assign w653 = w650 & ~w652;
assign w654 = w529 & ~w653;
assign w655 = ~pi0239 & w653;
assign w656 = w529 & ~w655;
assign w657 = (~w642 & w654) | (~w642 & w656) | (w654 & w656);
assign w658 = ~w627 & ~w657;
assign w659 = (w603 & ~w619) | (w603 & w625) | (~w619 & w625);
assign w660 = w9 & w114;
assign w661 = pi0235 & w7;
assign w662 = w660 & w661;
assign w663 = ~pi0151 & ~w9;
assign w664 = w114 & ~w663;
assign w665 = ~pi0927 & w610;
assign w666 = ~pi0221 & w612;
assign w667 = pi0274 & w666;
assign w668 = ~w665 & ~w667;
assign w669 = ~pi1145 & ~w21;
assign w670 = w668 & ~w669;
assign w671 = ~w664 & w670;
assign w672 = ~w662 & ~w671;
assign w673 = ~w659 & ~w672;
assign w674 = pi0235 & ~w642;
assign w675 = pi0833 & w644;
assign w676 = pi0927 & w675;
assign w677 = ~pi0274 & w648;
assign w678 = ~w676 & ~w677;
assign w679 = pi1145 & w517;
assign w680 = w678 & ~w679;
assign w681 = ~w674 & w680;
assign w682 = w529 & ~w681;
assign w683 = ~w673 & ~w682;
assign w684 = pi0228 & ~w9;
assign w685 = (~w9 & w205) | (~w9 & w684) | (w205 & w684);
assign w686 = w569 & ~w685;
assign w687 = (~w9 & w407) | (~w9 & w685) | (w407 & w685);
assign w688 = w569 & ~w687;
assign w689 = (w378 & w686) | (w378 & w688) | (w686 & w688);
assign w690 = ~pi0284 & w9;
assign w691 = ~w7 & w690;
assign w692 = pi0146 & ~w9;
assign w693 = w114 & w692;
assign w694 = (w114 & w691) | (w114 & w693) | (w691 & w693);
assign w695 = pi0944 & w610;
assign w696 = ~pi0221 & ~pi0264;
assign w697 = w612 & w696;
assign w698 = ~w695 & ~w697;
assign w699 = pi1143 & ~w21;
assign w700 = w698 & ~w699;
assign w701 = ~w694 & w700;
assign w702 = ~w115 & w701;
assign w703 = (~w113 & w701) | (~w113 & w702) | (w701 & w702);
assign w704 = ~pi0095 & w703;
assign w705 = ~w115 & ~w701;
assign w706 = (~w113 & ~w701) | (~w113 & w705) | (~w701 & w705);
assign w707 = ~pi0228 & ~pi0284;
assign w708 = w348 & w707;
assign w709 = w7 & w9;
assign w710 = w114 & w709;
assign w711 = (w114 & w708) | (w114 & w710) | (w708 & w710);
assign w712 = ~w706 & ~w711;
assign w713 = ~w704 & ~w712;
assign w714 = ~w689 & ~w713;
assign w715 = ~w7 & w569;
assign w716 = pi0284 & w715;
assign w717 = ~w433 & w716;
assign w718 = ~w685 & w717;
assign w719 = ~w687 & w717;
assign w720 = (w378 & w718) | (w378 & w719) | (w718 & w719);
assign w721 = pi0299 & w720;
assign w722 = (pi0299 & w714) | (pi0299 & w721) | (w714 & w721);
assign w723 = ~pi0299 & ~pi1143;
assign w724 = ~w516 & w723;
assign w725 = pi0833 & ~pi0944;
assign w726 = w644 & w725;
assign w727 = ~w724 & ~w726;
assign w728 = pi0264 & w648;
assign w729 = w529 & ~w728;
assign w730 = w727 & w729;
assign w731 = pi0238 & ~w642;
assign w732 = pi0284 & w16;
assign w733 = ~w492 & ~w732;
assign w734 = (~w640 & ~w732) | (~w640 & w733) | (~w732 & w733);
assign w735 = ~w633 & w734;
assign w736 = w730 & w735;
assign w737 = (w730 & w731) | (w730 & w736) | (w731 & w736);
assign w738 = ~w722 & w737;
assign w739 = pi0228 & pi0238;
assign w740 = w711 & w739;
assign w741 = ~w506 & ~w739;
assign w742 = w711 & ~w741;
assign w743 = (w554 & w740) | (w554 & w742) | (w740 & w742);
assign w744 = ~w506 & ~w701;
assign w745 = (~w554 & ~w701) | (~w554 & w744) | (~w701 & w744);
assign w746 = ~w743 & ~w745;
assign w747 = ~w529 & ~w746;
assign w748 = ~w738 & ~w747;
assign w749 = ~pi0249 & ~w435;
assign w750 = ~w9 & ~w622;
assign w751 = ~pi0228 & w6;
assign w752 = ~w205 & w751;
assign w753 = w750 & ~w752;
assign w754 = w6 & w206;
assign w755 = ~w407 & w754;
assign w756 = w750 & ~w755;
assign w757 = (~w378 & w753) | (~w378 & w756) | (w753 & w756);
assign w758 = w749 & ~w757;
assign w759 = (~w378 & w685) | (~w378 & w687) | (w685 & w687);
assign w760 = pi0262 & w435;
assign w761 = ~w759 & w760;
assign w762 = pi0172 & w759;
assign w763 = ~w761 & ~w762;
assign w764 = ~w758 & w763;
assign w765 = w12 & w593;
assign w766 = ~w764 & w765;
assign w767 = pi0215 & ~pi1142;
assign w768 = pi0216 & ~pi0221;
assign w769 = ~pi0277 & w768;
assign w770 = pi0932 & w19;
assign w771 = pi1142 & ~w19;
assign w772 = ~w770 & ~w771;
assign w773 = pi0221 & ~w772;
assign w774 = ~w769 & ~w773;
assign w775 = ~pi0215 & w774;
assign w776 = ~w767 & ~w775;
assign w777 = ~pi0228 & w83;
assign w778 = w74 & w777;
assign w779 = w553 & w778;
assign w780 = ~w9 & ~w779;
assign w781 = ~pi0172 & w780;
assign w782 = ~w709 & ~w781;
assign w783 = w529 & w622;
assign w784 = w780 & ~w783;
assign w785 = ~pi0262 & ~w784;
assign w786 = w782 & ~w785;
assign w787 = w114 & ~w786;
assign w788 = ~w776 & ~w787;
assign w789 = pi0262 & w116;
assign w790 = pi0299 & ~w789;
assign w791 = w529 & ~w790;
assign w792 = ~pi0249 & w710;
assign w793 = ~w791 & ~w792;
assign w794 = ~w788 & w793;
assign w795 = (~w7 & ~w433) | (~w7 & w631) | (~w433 & w631);
assign w796 = ~pi0262 & w795;
assign w797 = pi0249 & ~w795;
assign w798 = ~w796 & ~w797;
assign w799 = w16 & ~w798;
assign w800 = w6 & w12;
assign w801 = pi0932 & w675;
assign w802 = ~pi0277 & w648;
assign w803 = ~w801 & ~w802;
assign w804 = pi1142 & w517;
assign w805 = w803 & ~w804;
assign w806 = ~w800 & w805;
assign w807 = ~w799 & w806;
assign w808 = w529 & ~w807;
assign w809 = ~w794 & ~w808;
assign w810 = ~w766 & ~w809;
assign w811 = ~pi0299 & ~pi0861;
assign w812 = (~pi0299 & w7) | (~pi0299 & w811) | (w7 & w811);
assign w813 = ~w1 & ~w812;
assign w814 = (~w5 & ~w812) | (~w5 & w813) | (~w812 & w813);
assign w815 = ~w529 & ~w710;
assign w816 = pi0241 & ~w815;
assign w817 = w83 & w506;
assign w818 = w74 & w817;
assign w819 = w550 & w818;
assign w820 = pi0861 & w109;
assign w821 = w819 & w820;
assign w822 = ~w7 & w9;
assign w823 = pi0861 & w822;
assign w824 = ~pi0171 & ~w9;
assign w825 = w114 & ~w824;
assign w826 = ~w823 & w825;
assign w827 = ~pi1141 & ~w21;
assign w828 = ~w826 & ~w827;
assign w829 = pi0270 & w768;
assign w830 = ~pi0216 & pi0221;
assign w831 = pi0833 & ~pi0935;
assign w832 = w830 & w831;
assign w833 = ~w829 & ~w832;
assign w834 = ~pi0215 & ~w833;
assign w835 = w828 & ~w834;
assign w836 = w553 & w818;
assign w837 = w835 & ~w836;
assign w838 = ~w821 & ~w837;
assign w839 = w529 & ~w816;
assign w840 = (~w816 & w838) | (~w816 & w839) | (w838 & w839);
assign w841 = w529 & ~w629;
assign w842 = w529 & ~w632;
assign w843 = (~w433 & w841) | (~w433 & w842) | (w841 & w842);
assign w844 = ~w641 & w843;
assign w845 = ~w814 & w844;
assign w846 = (~w814 & w840) | (~w814 & w845) | (w840 & w845);
assign w847 = ~w7 & w114;
assign w848 = pi0861 & w847;
assign w849 = ~w433 & w848;
assign w850 = ~w685 & w849;
assign w851 = ~w687 & w849;
assign w852 = (w378 & w850) | (w378 & w851) | (w850 & w851);
assign w853 = pi0299 & ~w852;
assign w854 = w114 & ~w685;
assign w855 = w114 & ~w687;
assign w856 = (w378 & w854) | (w378 & w855) | (w854 & w855);
assign w857 = w835 & ~w856;
assign w858 = w853 & ~w857;
assign w859 = pi0861 & ~w7;
assign w860 = w16 & ~w859;
assign w861 = (w16 & w433) | (w16 & w860) | (w433 & w860);
assign w862 = w846 & w861;
assign w863 = (w846 & w858) | (w846 & w862) | (w858 & w862);
assign w864 = ~w840 & ~w844;
assign w865 = ~pi0861 & w115;
assign w866 = w113 & w865;
assign w867 = ~w115 & ~w835;
assign w868 = (~w113 & ~w835) | (~w113 & w867) | (~w835 & w867);
assign w869 = ~w866 & ~w868;
assign w870 = ~pi0299 & ~pi1141;
assign w871 = ~w516 & w870;
assign w872 = w644 & w831;
assign w873 = pi0270 & w648;
assign w874 = ~w872 & ~w873;
assign w875 = w529 & w874;
assign w876 = ~w871 & w875;
assign w877 = pi0299 & ~w6;
assign w878 = w875 & ~w877;
assign w879 = ~w871 & w878;
assign w880 = (w869 & w876) | (w869 & w879) | (w876 & w879);
assign w881 = ~w864 & ~w880;
assign w882 = ~w863 & ~w881;
assign w883 = pi1140 & ~w21;
assign w884 = ~pi0221 & ~pi0282;
assign w885 = pi0221 & ~pi0921;
assign w886 = ~pi0216 & ~w885;
assign w887 = ~w884 & ~w886;
assign w888 = w21 & ~w887;
assign w889 = ~w883 & ~w888;
assign w890 = w529 & ~w889;
assign w891 = pi0299 & w890;
assign w892 = w642 & w891;
assign w893 = (w378 & w752) | (w378 & w755) | (w752 & w755);
assign w894 = ~pi0869 & ~w750;
assign w895 = (~pi0869 & w893) | (~pi0869 & w894) | (w893 & w894);
assign w896 = pi0170 & w750;
assign w897 = ~w893 & w896;
assign w898 = ~w895 & ~w897;
assign w899 = ~w114 & w892;
assign w900 = (w892 & w898) | (w892 & w899) | (w898 & w899);
assign w901 = pi0248 & ~w815;
assign w902 = w629 & ~w901;
assign w903 = w632 & ~w901;
assign w904 = (w433 & w902) | (w433 & w903) | (w902 & w903);
assign w905 = pi0869 & w16;
assign w906 = ~pi0282 & w648;
assign w907 = ~w905 & ~w906;
assign w908 = ~pi0299 & pi1140;
assign w909 = ~w516 & w908;
assign w910 = pi0833 & pi0921;
assign w911 = w644 & w910;
assign w912 = ~w909 & ~w911;
assign w913 = w907 & w912;
assign w914 = w529 & ~w913;
assign w915 = ~w904 & w914;
assign w916 = ~w901 & ~w914;
assign w917 = ~w904 & ~w916;
assign w918 = (~w844 & w915) | (~w844 & w917) | (w915 & w917);
assign w919 = ~pi0170 & ~w9;
assign w920 = ~w779 & w919;
assign w921 = pi0869 & ~w7;
assign w922 = w9 & w921;
assign w923 = (w779 & w921) | (w779 & w922) | (w921 & w922);
assign w924 = ~w920 & ~w923;
assign w925 = ~w529 & ~w889;
assign w926 = ~w114 & ~w889;
assign w927 = ~w529 & w926;
assign w928 = (~w924 & w925) | (~w924 & w927) | (w925 & w927);
assign w929 = ~w918 & ~w928;
assign w930 = ~w900 & w929;
assign w931 = pi0862 & w435;
assign w932 = pi0247 & ~w435;
assign w933 = ~w931 & ~w932;
assign w934 = ~w759 & w933;
assign w935 = pi0148 & w759;
assign w936 = ~w934 & ~w935;
assign w937 = w569 & ~w936;
assign w938 = pi0862 & w116;
assign w939 = ~pi0247 & w7;
assign w940 = ~pi0862 & ~w7;
assign w941 = ~w939 & ~w940;
assign w942 = w9 & ~w941;
assign w943 = pi0148 & ~w9;
assign w944 = ~w942 & ~w943;
assign w945 = w114 & ~w944;
assign w946 = ~pi1139 & ~w21;
assign w947 = ~w945 & ~w946;
assign w948 = ~pi0920 & w610;
assign w949 = pi0281 & w666;
assign w950 = ~w948 & ~w949;
assign w951 = w947 & w950;
assign w952 = ~w569 & ~w951;
assign w953 = ~w116 & ~w952;
assign w954 = ~w938 & ~w953;
assign w955 = pi0247 & ~w795;
assign w956 = pi0862 & w795;
assign w957 = ~w955 & ~w956;
assign w958 = w16 & w957;
assign w959 = ~pi1139 & w517;
assign w960 = ~pi0920 & w675;
assign w961 = ~w959 & ~w960;
assign w962 = pi0281 & w648;
assign w963 = w529 & ~w962;
assign w964 = w961 & w963;
assign w965 = ~w958 & w964;
assign w966 = ~w954 & w965;
assign w967 = ~w937 & w966;
assign w968 = w506 & w554;
assign w969 = pi0862 & w968;
assign w970 = w951 & ~w968;
assign w971 = ~w969 & ~w970;
assign w972 = ~w529 & ~w971;
assign w973 = ~pi0299 & w965;
assign w974 = ~w972 & ~w973;
assign w975 = ~w967 & w974;
assign w976 = ~pi0877 & w435;
assign w977 = ~pi0246 & ~w435;
assign w978 = ~w976 & ~w977;
assign w979 = ~w759 & ~w978;
assign w980 = pi0169 & w759;
assign w981 = ~w979 & ~w980;
assign w982 = w569 & ~w981;
assign w983 = pi1138 & w517;
assign w984 = ~w633 & ~w983;
assign w985 = pi0940 & w675;
assign w986 = ~pi0269 & w648;
assign w987 = ~w985 & ~w986;
assign w988 = pi0877 & w16;
assign w989 = w987 & ~w988;
assign w990 = w984 & w989;
assign w991 = ~pi0246 & w633;
assign w992 = ~w990 & ~w991;
assign w993 = w529 & ~w992;
assign w994 = w982 & w993;
assign w995 = pi0246 & w710;
assign w996 = ~pi0169 & w780;
assign w997 = ~pi0228 & w109;
assign w998 = ~w822 & ~w997;
assign w999 = (~w551 & ~w822) | (~w551 & w998) | (~w822 & w998);
assign w1000 = pi0877 & ~w999;
assign w1001 = ~w996 & ~w1000;
assign w1002 = w114 & w1001;
assign w1003 = ~pi0940 & w610;
assign w1004 = pi0269 & w666;
assign w1005 = ~w1003 & ~w1004;
assign w1006 = ~pi1138 & ~w21;
assign w1007 = w1005 & ~w1006;
assign w1008 = ~w1002 & w1007;
assign w1009 = ~w995 & ~w1008;
assign w1010 = ~w529 & w1009;
assign w1011 = ~pi0169 & w750;
assign w1012 = pi0877 & ~w7;
assign w1013 = ~w750 & w1012;
assign w1014 = ~w1011 & ~w1013;
assign w1015 = ~w6 & w114;
assign w1016 = w1014 & w1015;
assign w1017 = pi0299 & ~w1016;
assign w1018 = w1007 & w1017;
assign w1019 = w993 & ~w1018;
assign w1020 = ~w1010 & ~w1019;
assign w1021 = ~w994 & w1020;
assign w1022 = ~pi0168 & w685;
assign w1023 = ~pi0168 & w687;
assign w1024 = (~w378 & w1022) | (~w378 & w1023) | (w1022 & w1023);
assign w1025 = pi0878 & ~w7;
assign w1026 = ~w433 & w1025;
assign w1027 = pi0240 & w7;
assign w1028 = (pi0240 & w433) | (pi0240 & w1027) | (w433 & w1027);
assign w1029 = ~w1026 & ~w1028;
assign w1030 = ~w685 & ~w1029;
assign w1031 = ~w687 & ~w1029;
assign w1032 = (w378 & w1030) | (w378 & w1031) | (w1030 & w1031);
assign w1033 = ~w1024 & ~w1032;
assign w1034 = ~pi0299 & ~pi1137;
assign w1035 = ~w516 & w1034;
assign w1036 = pi0833 & ~pi0933;
assign w1037 = w644 & w1036;
assign w1038 = ~w1035 & ~w1037;
assign w1039 = w529 & w1038;
assign w1040 = w16 & ~w1025;
assign w1041 = pi0280 & w648;
assign w1042 = ~w1040 & ~w1041;
assign w1043 = w1039 & w1042;
assign w1044 = ~w12 & ~w629;
assign w1045 = w6 & ~w1044;
assign w1046 = ~w12 & ~w632;
assign w1047 = w6 & ~w1046;
assign w1048 = (w433 & w1045) | (w433 & w1047) | (w1045 & w1047);
assign w1049 = ~pi0878 & w115;
assign w1050 = w113 & w1049;
assign w1051 = pi0878 & w9;
assign w1052 = ~w7 & w1051;
assign w1053 = ~pi0168 & ~w9;
assign w1054 = w114 & w1053;
assign w1055 = (w114 & w1052) | (w114 & w1054) | (w1052 & w1054);
assign w1056 = ~pi0221 & ~pi0280;
assign w1057 = w612 & w1056;
assign w1058 = ~w1055 & ~w1057;
assign w1059 = ~w115 & w1058;
assign w1060 = (~w113 & w1058) | (~w113 & w1059) | (w1058 & w1059);
assign w1061 = ~w1050 & ~w1060;
assign w1062 = pi1137 & ~w21;
assign w1063 = pi0933 & w610;
assign w1064 = ~w1062 & ~w1063;
assign w1065 = pi0299 & w1064;
assign w1066 = ~w1048 & ~w1065;
assign w1067 = (~w1048 & w1061) | (~w1048 & w1066) | (w1061 & w1066);
assign w1068 = w1043 & w1067;
assign w1069 = ~w1 & ~w709;
assign w1070 = (~w5 & ~w709) | (~w5 & w1069) | (~w709 & w1069);
assign w1071 = w12 & ~w1070;
assign w1072 = ~w1067 & ~w1071;
assign w1073 = w1043 & ~w1072;
assign w1074 = (~w1033 & w1068) | (~w1033 & w1073) | (w1068 & w1073);
assign w1075 = ~pi0062 & pi0240;
assign w1076 = w180 & w1075;
assign w1077 = w628 & w1076;
assign w1078 = w16 & ~w631;
assign w1079 = w1076 & w1078;
assign w1080 = (w433 & w1077) | (w433 & w1079) | (w1077 & w1079);
assign w1081 = ~pi0878 & w506;
assign w1082 = w554 & w1081;
assign w1083 = pi0240 & w710;
assign w1084 = ~w506 & ~w1083;
assign w1085 = w1058 & w1084;
assign w1086 = w1064 & w1085;
assign w1087 = w1058 & ~w1083;
assign w1088 = w1064 & w1087;
assign w1089 = (~w554 & w1086) | (~w554 & w1088) | (w1086 & w1088);
assign w1090 = ~w1082 & ~w1089;
assign w1091 = w529 & ~w1080;
assign w1092 = (~w1080 & ~w1090) | (~w1080 & w1091) | (~w1090 & w1091);
assign w1093 = ~w1074 & w1092;
assign w1094 = pi0928 & w610;
assign w1095 = ~pi0221 & pi0266;
assign w1096 = w612 & w1095;
assign w1097 = ~w1094 & ~w1096;
assign w1098 = pi1136 & ~w21;
assign w1099 = ~w526 & ~w1098;
assign w1100 = w1097 & w1099;
assign w1101 = w9 & ~w529;
assign w1102 = (~w529 & w779) | (~w529 & w1101) | (w779 & w1101);
assign w1103 = w9 & w529;
assign w1104 = (w529 & w622) | (w529 & w1103) | (w622 & w1103);
assign w1105 = ~w1102 & ~w1104;
assign w1106 = pi0875 & ~w1105;
assign w1107 = ~w9 & ~w529;
assign w1108 = ~w779 & w1107;
assign w1109 = ~w9 & w529;
assign w1110 = ~w622 & w1109;
assign w1111 = ~w1108 & ~w1110;
assign w1112 = pi0166 & ~w1111;
assign w1113 = ~w1106 & ~w1112;
assign w1114 = w759 & ~w1113;
assign w1115 = ~pi0875 & ~w7;
assign w1116 = ~w433 & w1115;
assign w1117 = ~pi0245 & w7;
assign w1118 = (~pi0245 & w433) | (~pi0245 & w1117) | (w433 & w1117);
assign w1119 = ~w1116 & ~w1118;
assign w1120 = ~w7 & ~w593;
assign w1121 = ~w593 & ~w709;
assign w1122 = (~w622 & w1120) | (~w622 & w1121) | (w1120 & w1121);
assign w1123 = ~w1119 & ~w1122;
assign w1124 = ~w1122 & ~w1123;
assign w1125 = (~w1113 & ~w1123) | (~w1113 & w1124) | (~w1123 & w1124);
assign w1126 = ~w759 & w1125;
assign w1127 = ~w1114 & ~w1126;
assign w1128 = ~w114 & w1100;
assign w1129 = (w1100 & w1127) | (w1100 & w1128) | (w1127 & w1128);
assign w1130 = ~pi0875 & w631;
assign w1131 = (~w433 & w1115) | (~w433 & w1130) | (w1115 & w1130);
assign w1132 = ~pi0245 & ~w631;
assign w1133 = (w433 & w1117) | (w433 & w1132) | (w1117 & w1132);
assign w1134 = ~w1131 & ~w1133;
assign w1135 = pi0833 & ~pi0928;
assign w1136 = w644 & w1135;
assign w1137 = ~pi0266 & w648;
assign w1138 = ~w1136 & ~w1137;
assign w1139 = ~pi0299 & ~pi1136;
assign w1140 = ~w516 & w1139;
assign w1141 = w1138 & ~w1140;
assign w1142 = w529 & ~w1141;
assign w1143 = ~w16 & w1141;
assign w1144 = w529 & ~w1143;
assign w1145 = (~w1134 & w1142) | (~w1134 & w1144) | (w1142 & w1144);
assign w1146 = ~w1129 & ~w1145;
assign w1147 = pi0244 & ~w642;
assign w1148 = ~w12 & ~w16;
assign w1149 = pi0879 & ~w1148;
assign w1150 = pi0879 & ~w56;
assign w1151 = (w622 & w1149) | (w622 & w1150) | (w1149 & w1150);
assign w1152 = w795 & w1151;
assign w1153 = pi0938 & w610;
assign w1154 = ~pi0221 & pi0279;
assign w1155 = w612 & w1154;
assign w1156 = ~w1153 & ~w1155;
assign w1157 = pi1135 & ~w21;
assign w1158 = pi0299 & w1157;
assign w1159 = (pi0299 & ~w1156) | (pi0299 & w1158) | (~w1156 & w1158);
assign w1160 = ~pi0299 & pi1135;
assign w1161 = ~w516 & w1160;
assign w1162 = ~w1159 & ~w1161;
assign w1163 = pi0833 & pi0938;
assign w1164 = w644 & w1163;
assign w1165 = pi0279 & w648;
assign w1166 = ~w1164 & ~w1165;
assign w1167 = w529 & w1166;
assign w1168 = w1162 & w1167;
assign w1169 = ~w1152 & w1168;
assign w1170 = ~w1147 & w1169;
assign w1171 = pi0161 & w757;
assign w1172 = pi0879 & ~w7;
assign w1173 = ~w433 & w1172;
assign w1174 = ~w757 & w1173;
assign w1175 = ~w1171 & ~w1174;
assign w1176 = ~w12 & w1170;
assign w1177 = (w1170 & w1175) | (w1170 & w1176) | (w1175 & w1176);
assign w1178 = pi0879 & ~w999;
assign w1179 = pi0244 & w709;
assign w1180 = pi0161 & ~w9;
assign w1181 = ~w1179 & ~w1180;
assign w1182 = (w779 & ~w1179) | (w779 & w1181) | (~w1179 & w1181);
assign w1183 = w114 & ~w1182;
assign w1184 = (w114 & w1178) | (w114 & w1183) | (w1178 & w1183);
assign w1185 = w1156 & ~w1157;
assign w1186 = ~w529 & w1185;
assign w1187 = ~w1184 & w1186;
assign w1188 = ~w1177 & ~w1187;
assign w1189 = ~pi0152 & w757;
assign w1190 = w636 & ~w639;
assign w1191 = ~w633 & ~w1190;
assign w1192 = pi0846 & w1191;
assign w1193 = pi0242 & ~w1191;
assign w1194 = ~w1192 & ~w1193;
assign w1195 = ~w757 & w1194;
assign w1196 = ~w1189 & ~w1195;
assign w1197 = ~pi0846 & ~w7;
assign w1198 = ~pi0242 & w7;
assign w1199 = ~w1197 & ~w1198;
assign w1200 = ~w780 & w1199;
assign w1201 = pi0152 & w780;
assign w1202 = ~w1200 & ~w1201;
assign w1203 = w114 & w1202;
assign w1204 = ~pi0930 & w610;
assign w1205 = ~pi0278 & w666;
assign w1206 = ~w1204 & ~w1205;
assign w1207 = ~w1203 & w1206;
assign w1208 = ~w529 & w1207;
assign w1209 = ~w1196 & ~w1208;
assign w1210 = w12 & w1209;
assign w1211 = pi0242 & ~w795;
assign w1212 = pi0846 & w795;
assign w1213 = ~w1211 & ~w1212;
assign w1214 = w16 & w1213;
assign w1215 = ~pi0930 & w675;
assign w1216 = ~pi0278 & w648;
assign w1217 = ~w1215 & ~w1216;
assign w1218 = w529 & w1217;
assign w1219 = pi0299 & ~w1206;
assign w1220 = w1218 & ~w1219;
assign w1221 = ~w1214 & w1220;
assign w1222 = ~w1208 & ~w1221;
assign w1223 = ~w517 & w526;
assign w1224 = w21 & ~w526;
assign w1225 = ~w1223 & ~w1224;
assign w1226 = ~pi1134 & w1225;
assign w1227 = ~w1222 & ~w1226;
assign w1228 = ~w1210 & w1227;
assign w1229 = ~pi0252 & ~pi1001;
assign w1230 = ~pi0287 & ~pi0984;
assign w1231 = ~w1229 & w1230;
assign w1232 = pi0835 & ~pi0979;
assign w1233 = w1231 & w1232;
assign w1234 = pi1091 & pi1093;
assign w1235 = ~w449 & w1234;
assign w1236 = w453 & w1235;
assign w1237 = w1233 & w1236;
assign w1238 = ~pi0907 & ~pi0947;
assign w1239 = ~pi0960 & ~pi0963;
assign w1240 = w1238 & w1239;
assign w1241 = ~pi0332 & ~pi0468;
assign w1242 = w1240 & w1241;
assign w1243 = ~pi0970 & ~pi0972;
assign w1244 = ~pi0975 & ~pi0978;
assign w1245 = w1243 & w1244;
assign w1246 = w1242 & w1245;
assign w1247 = pi0603 & ~pi0614;
assign w1248 = ~pi0616 & ~pi0642;
assign w1249 = w1247 & w1248;
assign w1250 = ~w1241 & ~w1249;
assign w1251 = ~pi0661 & ~pi0662;
assign w1252 = pi0680 & ~pi0681;
assign w1253 = w1251 & w1252;
assign w1254 = w1250 & ~w1253;
assign w1255 = ~w1246 & ~w1254;
assign w1256 = pi0221 & pi0299;
assign w1257 = w612 & w1256;
assign w1258 = w1255 & w1257;
assign w1259 = w643 & w647;
assign w1260 = ~pi0587 & ~pi0602;
assign w1261 = ~pi0961 & ~pi0967;
assign w1262 = w1260 & w1261;
assign w1263 = w1241 & w1262;
assign w1264 = ~pi0969 & ~pi0971;
assign w1265 = ~pi0974 & ~pi0977;
assign w1266 = w1264 & w1265;
assign w1267 = w1263 & w1266;
assign w1268 = ~w1254 & ~w1267;
assign w1269 = w1259 & w1268;
assign w1270 = ~w1258 & ~w1269;
assign w1271 = w1237 & ~w1270;
assign w1272 = w5 & ~w1271;
assign w1273 = ~pi0299 & w1241;
assign w1274 = w1262 & w1266;
assign w1275 = w1273 & w1274;
assign w1276 = ~w1241 & ~w1253;
assign w1277 = ~w1249 & w1276;
assign w1278 = ~w1275 & ~w1277;
assign w1279 = w449 & w1234;
assign w1280 = pi0950 & pi1092;
assign w1281 = ~w1279 & w1280;
assign w1282 = ~pi0824 & ~pi0829;
assign w1283 = (~pi0824 & w450) | (~pi0824 & w1282) | (w450 & w1282);
assign w1284 = w1281 & ~w1283;
assign w1285 = w1278 & w1284;
assign w1286 = w1241 & w1245;
assign w1287 = w1240 & w1286;
assign w1288 = pi0215 & ~w1287;
assign w1289 = pi0299 & ~w1288;
assign w1290 = ~pi0223 & ~pi0299;
assign w1291 = ~w1289 & ~w1290;
assign w1292 = w1285 & w1291;
assign w1293 = w1233 & w1292;
assign w1294 = w1272 & ~w1293;
assign w1295 = pi0039 & ~w1294;
assign w1296 = w109 & w529;
assign w1297 = w112 & w1296;
assign w1298 = ~w1295 & w1297;
assign w1299 = ~pi0092 & w147;
assign w1300 = w118 & w1299;
assign w1301 = ~pi0054 & w1300;
assign w1302 = ~pi0092 & w168;
assign w1303 = ~pi0075 & w1302;
assign w1304 = ~w1301 & ~w1303;
assign w1305 = w1298 & ~w1304;
assign w1306 = ~pi0087 & ~pi0100;
assign w1307 = ~w117 & w1306;
assign w1308 = ~pi0074 & ~w1307;
assign w1309 = ~pi0087 & pi0100;
assign w1310 = ~pi0042 & ~pi0043;
assign w1311 = ~pi0114 & ~pi0115;
assign w1312 = w1310 & w1311;
assign w1313 = ~pi0052 & ~pi0116;
assign w1314 = w1312 & w1313;
assign w1315 = ~pi0041 & ~pi0044;
assign w1316 = ~pi0099 & ~pi0101;
assign w1317 = w1315 & w1316;
assign w1318 = ~pi0113 & w1317;
assign w1319 = w1314 & w1318;
assign w1320 = w448 & ~w1319;
assign w1321 = pi1092 & ~pi1093;
assign w1322 = ~w1282 & w1321;
assign w1323 = pi0129 & pi0250;
assign w1324 = pi0250 & ~w1323;
assign w1325 = ~pi0250 & ~pi0950;
assign w1326 = ~w1323 & ~w1325;
assign w1327 = (w1322 & w1324) | (w1322 & w1326) | (w1324 & w1326);
assign w1328 = pi0683 & ~w1327;
assign w1329 = w1320 & w1328;
assign w1330 = pi0252 & ~w448;
assign w1331 = ~w1329 & ~w1330;
assign w1332 = w1309 & w1331;
assign w1333 = pi0087 & ~pi0100;
assign w1334 = ~w1332 & ~w1333;
assign w1335 = w117 & ~w1334;
assign w1336 = w1308 & ~w1335;
assign w1337 = w1305 & ~w1336;
assign w1338 = w546 & w567;
assign w1339 = ~pi0055 & w1338;
assign w1340 = w571 & w1339;
assign w1341 = ~pi0032 & ~pi0095;
assign w1342 = w188 & w1341;
assign w1343 = w542 & w1342;
assign w1344 = ~pi0071 & ~pi0084;
assign w1345 = w79 & w1344;
assign w1346 = w64 & w1345;
assign w1347 = w60 & w72;
assign w1348 = w1346 & w1347;
assign w1349 = w66 & w229;
assign w1350 = ~pi0098 & ~pi0102;
assign w1351 = w1349 & w1350;
assign w1352 = w1348 & w1351;
assign w1353 = w1343 & w1352;
assign w1354 = ~pi0073 & w99;
assign w1355 = w1353 & w1354;
assign w1356 = ~w1340 & ~w1355;
assign w1357 = pi0095 & w347;
assign w1358 = w194 & w196;
assign w1359 = w593 & w1358;
assign w1360 = w1357 & w1359;
assign w1361 = w1356 & ~w1360;
assign w1362 = ~w1337 & w1361;
assign w1363 = ~pi0841 & w413;
assign w1364 = pi0032 & ~w1363;
assign w1365 = ~pi0841 & w400;
assign w1366 = w105 & ~w399;
assign w1367 = ~w1365 & w1366;
assign w1368 = w494 & w1367;
assign w1369 = ~w1364 & w1368;
assign w1370 = w486 & w1369;
assign w1371 = w83 & w402;
assign w1372 = w74 & w1371;
assign w1373 = ~w99 & w349;
assign w1374 = (w349 & ~w1372) | (w349 & w1373) | (~w1372 & w1373);
assign w1375 = ~w376 & w1374;
assign w1376 = ~w489 & w1374;
assign w1377 = (w486 & w1375) | (w486 & w1376) | (w1375 & w1376);
assign w1378 = ~w441 & w593;
assign w1379 = ~w1377 & w1378;
assign w1380 = ~w1370 & w1379;
assign w1381 = w1362 & ~w1380;
assign w1382 = ~w387 & w1374;
assign w1383 = ~w487 & w1382;
assign w1384 = ~pi0228 & ~w1383;
assign w1385 = (~pi0228 & ~w486) | (~pi0228 & w1384) | (~w486 & w1384);
assign w1386 = ~pi0032 & w7;
assign w1387 = w188 & w1386;
assign w1388 = w1354 & w1387;
assign w1389 = w1352 & w1388;
assign w1390 = pi0032 & ~pi0040;
assign w1391 = ~pi0095 & w1390;
assign w1392 = w413 & w1391;
assign w1393 = ~pi0841 & w1392;
assign w1394 = w196 & w1393;
assign w1395 = w194 & w1394;
assign w1396 = ~w1389 & ~w1395;
assign w1397 = w349 & w593;
assign w1398 = ~w104 & ~w349;
assign w1399 = (~w349 & w393) | (~w349 & w1398) | (w393 & w1398);
assign w1400 = w593 & ~w1399;
assign w1401 = (w492 & w1397) | (w492 & w1400) | (w1397 & w1400);
assign w1402 = (w593 & ~w1396) | (w593 & w1401) | (~w1396 & w1401);
assign w1403 = ~w1375 & w1402;
assign w1404 = pi0103 & ~pi0314;
assign w1405 = ~pi0072 & ~w1404;
assign w1406 = ~pi0081 & w196;
assign w1407 = ~w481 & w1406;
assign w1408 = ~pi0066 & pi0084;
assign w1409 = pi0066 & ~pi0084;
assign w1410 = ~w1408 & ~w1409;
assign w1411 = ~pi0073 & ~w1410;
assign w1412 = ~pi0066 & ~pi0084;
assign w1413 = ~pi0068 & pi0073;
assign w1414 = w1412 & w1413;
assign w1415 = (~pi0068 & w1411) | (~pi0068 & w1414) | (w1411 & w1414);
assign w1416 = pi0068 & ~pi0073;
assign w1417 = w1412 & w1416;
assign w1418 = ~pi0082 & ~pi0085;
assign w1419 = ~w1417 & w1418;
assign w1420 = ~w1415 & w1419;
assign w1421 = ~pi0085 & ~w1417;
assign w1422 = ~w1415 & w1421;
assign w1423 = ~pi0067 & w333;
assign w1424 = pi0069 & pi0083;
assign w1425 = ~w1423 & ~w1424;
assign w1426 = ~pi0071 & ~pi0082;
assign w1427 = pi0067 & ~pi0071;
assign w1428 = ~w333 & w1427;
assign w1429 = ~pi0082 & w1428;
assign w1430 = (~w1425 & w1426) | (~w1425 & w1429) | (w1426 & w1429);
assign w1431 = ~w196 & w1430;
assign w1432 = w1422 & w1431;
assign w1433 = (w1407 & w1420) | (w1407 & w1432) | (w1420 & w1432);
assign w1434 = ~pi0058 & ~pi0110;
assign w1435 = ~pi0047 & w1434;
assign w1436 = w494 & w1435;
assign w1437 = w1367 & w1436;
assign w1438 = w1405 & ~w1437;
assign w1439 = (w1405 & w1433) | (w1405 & w1438) | (w1433 & w1438);
assign w1440 = w1403 & ~w1439;
assign w1441 = w1385 & w1440;
assign w1442 = pi0252 & w134;
assign w1443 = ~w448 & w1442;
assign w1444 = (w134 & w1329) | (w134 & w1443) | (w1329 & w1443);
assign w1445 = ~pi0030 & pi0228;
assign w1446 = ~pi0062 & ~w1445;
assign w1447 = w180 & w1446;
assign w1448 = pi0075 & ~pi0092;
assign w1449 = ~pi0075 & pi0092;
assign w1450 = ~w1448 & ~w1449;
assign w1451 = ~pi0074 & ~w1450;
assign w1452 = ~pi0075 & ~pi0092;
assign w1453 = ~pi0054 & pi0074;
assign w1454 = w1452 & w1453;
assign w1455 = (~pi0054 & w1451) | (~pi0054 & w1454) | (w1451 & w1454);
assign w1456 = w117 & w1306;
assign w1457 = pi0054 & ~pi0074;
assign w1458 = w1452 & w1457;
assign w1459 = ~pi0100 & w1458;
assign w1460 = w118 & w1459;
assign w1461 = (w1455 & w1456) | (w1455 & w1460) | (w1456 & w1460);
assign w1462 = w1447 & w1461;
assign w1463 = w4 & ~w54;
assign w1464 = ~w1461 & ~w1463;
assign w1465 = w1447 & ~w1464;
assign w1466 = (w1444 & w1462) | (w1444 & w1465) | (w1462 & w1465);
assign w1467 = ~pi0215 & pi0221;
assign w1468 = ~pi0216 & pi0299;
assign w1469 = w1467 & w1468;
assign w1470 = ~w644 & ~w1469;
assign w1471 = w1237 & w1470;
assign w1472 = pi0829 & pi1091;
assign w1473 = (pi1091 & w449) | (pi1091 & w1472) | (w449 & w1472);
assign w1474 = pi0824 & pi0950;
assign w1475 = pi1092 & pi1093;
assign w1476 = w1474 & w1475;
assign w1477 = ~w1473 & w1476;
assign w1478 = w1233 & w1477;
assign w1479 = ~pi0038 & w1478;
assign w1480 = (~pi0038 & w1471) | (~pi0038 & w1479) | (w1471 & w1479);
assign w1481 = w171 & w529;
assign w1482 = pi0038 & ~pi0039;
assign w1483 = ~pi0228 & w1482;
assign w1484 = w1481 & w1483;
assign w1485 = ~pi0228 & w1481;
assign w1486 = ~pi0299 & w643;
assign w1487 = pi0299 & w1467;
assign w1488 = ~w1486 & ~w1487;
assign w1489 = ~pi0039 & ~w1482;
assign w1490 = (~w1482 & w1488) | (~w1482 & w1489) | (w1488 & w1489);
assign w1491 = w1485 & ~w1490;
assign w1492 = (w1480 & w1484) | (w1480 & w1491) | (w1484 & w1491);
assign w1493 = w113 & w1492;
assign w1494 = (w113 & w1466) | (w113 & w1493) | (w1466 & w1493);
assign w1495 = pi0228 & w1447;
assign w1496 = ~w1494 & ~w1495;
assign w1497 = ~w1241 & w1253;
assign w1498 = pi0158 & pi0159;
assign w1499 = pi0160 & pi0197;
assign w1500 = w1498 & w1499;
assign w1501 = pi0109 & pi0232;
assign w1502 = ~pi0228 & w1501;
assign w1503 = w1500 & w1502;
assign w1504 = ~w526 & ~w1503;
assign w1505 = pi0907 & w1241;
assign w1506 = ~w1497 & ~w1505;
assign w1507 = (~w1497 & ~w1504) | (~w1497 & w1506) | (~w1504 & w1506);
assign w1508 = pi0232 & w1500;
assign w1509 = pi0109 & pi0299;
assign w1510 = pi0109 & pi0145;
assign w1511 = pi0180 & pi0181;
assign w1512 = w1510 & w1511;
assign w1513 = pi0182 & pi0232;
assign w1514 = ~w1509 & ~w1513;
assign w1515 = (~w1509 & ~w1512) | (~w1509 & w1514) | (~w1512 & w1514);
assign w1516 = w1508 & ~w1515;
assign w1517 = ~pi0299 & w1513;
assign w1518 = w1512 & w1517;
assign w1519 = w1241 & w1518;
assign w1520 = (w1241 & w1516) | (w1241 & w1519) | (w1516 & w1519);
assign w1521 = w1507 & w1520;
assign w1522 = w1496 & w1521;
assign w1523 = pi0030 & pi0228;
assign w1524 = pi0062 & w1523;
assign w1525 = (~w180 & w1523) | (~w180 & w1524) | (w1523 & w1524);
assign w1526 = ~w529 & w1523;
assign w1527 = pi0228 & ~w1523;
assign w1528 = ~w529 & ~w1527;
assign w1529 = (w577 & w1526) | (w577 & w1528) | (w1526 & w1528);
assign w1530 = (w567 & w1525) | (w567 & w1529) | (w1525 & w1529);
assign w1531 = ~w1507 & w1530;
assign w1532 = ~w1521 & w1531;
assign w1533 = w1496 & ~w1532;
assign w1534 = (~w1441 & w1522) | (~w1441 & w1533) | (w1522 & w1533);
assign w1535 = ~pi0299 & pi0602;
assign w1536 = w1241 & w1535;
assign w1537 = w1507 & ~w1536;
assign w1538 = ~w1534 & ~w1537;
assign w1539 = ~pi0228 & ~w1520;
assign w1540 = ~w1383 & w1539;
assign w1541 = (~w486 & w1539) | (~w486 & w1540) | (w1539 & w1540);
assign w1542 = ~w1440 & w1496;
assign w1543 = (w1496 & ~w1541) | (w1496 & w1542) | (~w1541 & w1542);
assign w1544 = pi0299 & ~pi0947;
assign w1545 = ~pi0299 & ~pi0587;
assign w1546 = ~w1544 & ~w1545;
assign w1547 = w1241 & ~w1546;
assign w1548 = ~w1250 & ~w1547;
assign w1549 = ~w1543 & w1548;
assign w1550 = pi0947 & w1241;
assign w1551 = ~w1241 & w1249;
assign w1552 = ~w1550 & ~w1551;
assign w1553 = w1525 & ~w1552;
assign w1554 = w1529 & ~w1552;
assign w1555 = (w567 & w1553) | (w567 & w1554) | (w1553 & w1554);
assign w1556 = ~w1549 & ~w1555;
assign w1557 = w1440 & w1541;
assign w1558 = w1241 & w1504;
assign w1559 = pi0970 & w1558;
assign w1560 = w1530 & w1559;
assign w1561 = w1496 & ~w1560;
assign w1562 = ~w1557 & w1561;
assign w1563 = pi0967 & w1273;
assign w1564 = ~w1559 & ~w1563;
assign w1565 = ~w1562 & ~w1564;
assign w1566 = w1500 & w1501;
assign w1567 = pi0299 & pi0972;
assign w1568 = ~w1566 & w1567;
assign w1569 = w1512 & w1513;
assign w1570 = ~pi0299 & pi0961;
assign w1571 = ~w1569 & w1570;
assign w1572 = ~w1568 & ~w1571;
assign w1573 = w1441 & ~w1572;
assign w1574 = ~w1567 & ~w1570;
assign w1575 = ~w1496 & ~w1574;
assign w1576 = pi0972 & w1530;
assign w1577 = ~w1575 & ~w1576;
assign w1578 = ~w1573 & w1577;
assign w1579 = w1241 & ~w1578;
assign w1580 = pi0960 & w1558;
assign w1581 = w1530 & w1580;
assign w1582 = w1496 & ~w1581;
assign w1583 = ~w1557 & w1582;
assign w1584 = pi0977 & w1273;
assign w1585 = ~w1580 & ~w1584;
assign w1586 = ~w1583 & ~w1585;
assign w1587 = pi0963 & w1558;
assign w1588 = w1530 & w1587;
assign w1589 = w1496 & ~w1588;
assign w1590 = ~w1557 & w1589;
assign w1591 = pi0969 & w1273;
assign w1592 = ~w1587 & ~w1591;
assign w1593 = ~w1590 & ~w1592;
assign w1594 = pi0975 & w1558;
assign w1595 = w1530 & w1594;
assign w1596 = w1496 & ~w1595;
assign w1597 = ~w1557 & w1596;
assign w1598 = pi0971 & w1273;
assign w1599 = ~w1594 & ~w1598;
assign w1600 = ~w1597 & ~w1599;
assign w1601 = pi0978 & w1558;
assign w1602 = w1530 & w1601;
assign w1603 = w1496 & ~w1602;
assign w1604 = ~w1557 & w1603;
assign w1605 = pi0974 & w1273;
assign w1606 = ~w1601 & ~w1605;
assign w1607 = ~w1604 & ~w1606;
assign w1608 = ~w1383 & ~w1520;
assign w1609 = (~w486 & ~w1520) | (~w486 & w1608) | (~w1520 & w1608);
assign w1610 = ~pi0954 & ~w1440;
assign w1611 = (~pi0954 & ~w1609) | (~pi0954 & w1610) | (~w1609 & w1610);
assign w1612 = w567 & w577;
assign w1613 = w109 & w1481;
assign w1614 = w112 & w1613;
assign w1615 = w1482 & w1614;
assign w1616 = ~w1612 & ~w1615;
assign w1617 = w109 & w1461;
assign w1618 = w112 & w1617;
assign w1619 = w529 & w1618;
assign w1620 = w1616 & ~w1619;
assign w1621 = w118 & w1302;
assign w1622 = w1297 & w1621;
assign w1623 = w1444 & w1622;
assign w1624 = w529 & w1486;
assign w1625 = w1268 & w1624;
assign w1626 = ~pi0215 & ~w526;
assign w1627 = pi0221 & w1626;
assign w1628 = w1255 & w1627;
assign w1629 = ~w1625 & ~w1628;
assign w1630 = w1478 & ~w1629;
assign w1631 = ~w1271 & ~w1630;
assign w1632 = w65 & w193;
assign w1633 = w1354 & w1632;
assign w1634 = ~pi0051 & ~pi0087;
assign w1635 = w1345 & w1634;
assign w1636 = w1633 & w1635;
assign w1637 = ~pi0035 & ~pi0070;
assign w1638 = w428 & w1637;
assign w1639 = w72 & w1638;
assign w1640 = ~pi0095 & ~pi0096;
assign w1641 = w347 & w1640;
assign w1642 = w5 & w1641;
assign w1643 = w1639 & w1642;
assign w1644 = ~pi0062 & ~pi0092;
assign w1645 = pi0039 & ~pi0072;
assign w1646 = w1644 & w1645;
assign w1647 = w180 & w1646;
assign w1648 = w1643 & w1647;
assign w1649 = w1636 & w1648;
assign w1650 = ~w1631 & w1649;
assign w1651 = ~w1623 & ~w1650;
assign w1652 = w1620 & w1651;
assign w1653 = w1611 & w1652;
assign w1654 = pi0024 & pi0954;
assign w1655 = ~w1653 & ~w1654;
assign w1656 = ~pi0228 & ~w603;
assign w1657 = pi0087 & pi0092;
assign w1658 = ~pi0087 & ~pi0092;
assign w1659 = ~w1657 & ~w1658;
assign w1660 = ~pi0039 & ~w1659;
assign w1661 = w1330 & w1660;
assign w1662 = w109 & w1463;
assign w1663 = w112 & w1662;
assign w1664 = w529 & w1663;
assign w1665 = ~w1661 & w1664;
assign w1666 = w1656 & ~w1665;
assign w1667 = ~w154 & ~w1666;
assign w1668 = ~pi0119 & ~pi0228;
assign w1669 = pi0252 & w1668;
assign w1670 = pi0119 & ~pi1056;
assign w1671 = ~w1669 & ~w1670;
assign w1672 = ~pi0468 & ~w1671;
assign w1673 = pi0119 & ~pi1077;
assign w1674 = ~w1669 & ~w1673;
assign w1675 = ~pi0468 & ~w1674;
assign w1676 = pi0119 & ~pi1073;
assign w1677 = ~w1669 & ~w1676;
assign w1678 = ~pi0468 & ~w1677;
assign w1679 = pi0119 & ~pi1041;
assign w1680 = ~w1669 & ~w1679;
assign w1681 = ~pi0468 & ~w1680;
assign w1682 = ~pi0378 & pi0379;
assign w1683 = pi0378 & ~pi0379;
assign w1684 = ~w1682 & ~w1683;
assign w1685 = ~pi0381 & ~pi0382;
assign w1686 = pi0381 & pi0382;
assign w1687 = ~w1685 & ~w1686;
assign w1688 = ~w1684 & ~w1687;
assign w1689 = pi0381 & ~pi0382;
assign w1690 = ~pi0381 & pi0382;
assign w1691 = ~w1689 & ~w1690;
assign w1692 = pi0378 & pi0379;
assign w1693 = ~pi0378 & ~pi0379;
assign w1694 = ~w1692 & ~w1693;
assign w1695 = ~w1691 & ~w1694;
assign w1696 = ~w1688 & ~w1695;
assign w1697 = pi0385 & pi0439;
assign w1698 = ~pi0385 & ~pi0439;
assign w1699 = ~w1697 & ~w1698;
assign w1700 = ~w1696 & ~w1699;
assign w1701 = ~w1684 & ~w1691;
assign w1702 = ~w1687 & ~w1694;
assign w1703 = ~w1701 & ~w1702;
assign w1704 = pi0385 & ~pi0439;
assign w1705 = ~pi0385 & pi0439;
assign w1706 = ~w1704 & ~w1705;
assign w1707 = ~w1703 & ~w1706;
assign w1708 = ~w1700 & ~w1707;
assign w1709 = pi0317 & w1708;
assign w1710 = ~pi0317 & ~w1708;
assign w1711 = ~w1709 & ~w1710;
assign w1712 = ~pi0376 & ~pi0377;
assign w1713 = pi0376 & pi0377;
assign w1714 = ~w1712 & ~w1713;
assign w1715 = ~w1711 & ~w1714;
assign w1716 = pi0317 & ~w1708;
assign w1717 = ~pi0317 & w1708;
assign w1718 = ~w1716 & ~w1717;
assign w1719 = pi0376 & ~pi0377;
assign w1720 = ~pi0376 & pi0377;
assign w1721 = ~w1719 & ~w1720;
assign w1722 = ~w1718 & ~w1721;
assign w1723 = ~w1715 & ~w1722;
assign w1724 = pi1199 & ~w1723;
assign w1725 = ~pi0363 & pi0372;
assign w1726 = pi0363 & ~pi0372;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = ~pi0380 & ~pi0386;
assign w1729 = pi0380 & pi0386;
assign w1730 = ~w1728 & ~w1729;
assign w1731 = ~w1727 & ~w1730;
assign w1732 = pi0380 & ~pi0386;
assign w1733 = ~pi0380 & pi0386;
assign w1734 = ~w1732 & ~w1733;
assign w1735 = pi0363 & pi0372;
assign w1736 = ~pi0363 & ~pi0372;
assign w1737 = ~w1735 & ~w1736;
assign w1738 = ~w1734 & ~w1737;
assign w1739 = ~w1731 & ~w1738;
assign w1740 = pi0387 & pi0388;
assign w1741 = ~pi0387 & ~pi0388;
assign w1742 = ~w1740 & ~w1741;
assign w1743 = ~w1739 & ~w1742;
assign w1744 = ~w1727 & ~w1734;
assign w1745 = ~w1730 & ~w1737;
assign w1746 = ~w1744 & ~w1745;
assign w1747 = pi0387 & ~pi0388;
assign w1748 = ~pi0387 & pi0388;
assign w1749 = ~w1747 & ~w1748;
assign w1750 = ~w1746 & ~w1749;
assign w1751 = ~w1743 & ~w1750;
assign w1752 = pi0337 & w1751;
assign w1753 = ~pi0337 & ~w1751;
assign w1754 = ~w1752 & ~w1753;
assign w1755 = ~pi0338 & ~pi0339;
assign w1756 = pi0338 & pi0339;
assign w1757 = ~w1755 & ~w1756;
assign w1758 = ~w1754 & ~w1757;
assign w1759 = pi0337 & ~w1751;
assign w1760 = ~pi0337 & w1751;
assign w1761 = ~w1759 & ~w1760;
assign w1762 = pi0338 & ~pi0339;
assign w1763 = ~pi0338 & pi0339;
assign w1764 = ~w1762 & ~w1763;
assign w1765 = ~w1761 & ~w1764;
assign w1766 = ~w1758 & ~w1765;
assign w1767 = pi1196 & ~w1766;
assign w1768 = ~w1724 & ~w1767;
assign w1769 = ~pi0366 & pi0367;
assign w1770 = pi0366 & ~pi0367;
assign w1771 = ~w1769 & ~w1770;
assign w1772 = ~pi0368 & ~pi0383;
assign w1773 = pi0368 & pi0383;
assign w1774 = ~w1772 & ~w1773;
assign w1775 = ~w1771 & ~w1774;
assign w1776 = pi0368 & ~pi0383;
assign w1777 = ~pi0368 & pi0383;
assign w1778 = ~w1776 & ~w1777;
assign w1779 = pi0366 & pi0367;
assign w1780 = ~pi0366 & ~pi0367;
assign w1781 = ~w1779 & ~w1780;
assign w1782 = ~w1778 & ~w1781;
assign w1783 = ~w1775 & ~w1782;
assign w1784 = pi0389 & pi0447;
assign w1785 = ~pi0389 & ~pi0447;
assign w1786 = ~w1784 & ~w1785;
assign w1787 = ~w1783 & ~w1786;
assign w1788 = ~w1771 & ~w1778;
assign w1789 = ~w1774 & ~w1781;
assign w1790 = ~w1788 & ~w1789;
assign w1791 = pi0389 & ~pi0447;
assign w1792 = ~pi0389 & pi0447;
assign w1793 = ~w1791 & ~w1792;
assign w1794 = ~w1790 & ~w1793;
assign w1795 = ~w1787 & ~w1794;
assign w1796 = pi0336 & w1795;
assign w1797 = ~pi0336 & ~w1795;
assign w1798 = ~w1796 & ~w1797;
assign w1799 = ~pi0364 & ~pi0365;
assign w1800 = pi0364 & pi0365;
assign w1801 = ~w1799 & ~w1800;
assign w1802 = ~w1798 & ~w1801;
assign w1803 = pi0336 & ~w1795;
assign w1804 = ~pi0336 & w1795;
assign w1805 = ~w1803 & ~w1804;
assign w1806 = pi0364 & ~pi0365;
assign w1807 = ~pi0364 & pi0365;
assign w1808 = ~w1806 & ~w1807;
assign w1809 = ~w1805 & ~w1808;
assign w1810 = ~w1802 & ~w1809;
assign w1811 = pi1197 & ~w1810;
assign w1812 = ~pi0373 & pi0374;
assign w1813 = pi0373 & ~pi0374;
assign w1814 = ~w1812 & ~w1813;
assign w1815 = ~pi0375 & ~pi0384;
assign w1816 = pi0375 & pi0384;
assign w1817 = ~w1815 & ~w1816;
assign w1818 = ~w1814 & ~w1817;
assign w1819 = pi0375 & ~pi0384;
assign w1820 = ~pi0375 & pi0384;
assign w1821 = ~w1819 & ~w1820;
assign w1822 = pi0373 & pi0374;
assign w1823 = ~pi0373 & ~pi0374;
assign w1824 = ~w1822 & ~w1823;
assign w1825 = ~w1821 & ~w1824;
assign w1826 = ~w1818 & ~w1825;
assign w1827 = pi0440 & pi0442;
assign w1828 = ~pi0440 & ~pi0442;
assign w1829 = ~w1827 & ~w1828;
assign w1830 = ~w1826 & ~w1829;
assign w1831 = ~w1814 & ~w1821;
assign w1832 = ~w1817 & ~w1824;
assign w1833 = ~w1831 & ~w1832;
assign w1834 = pi0440 & ~pi0442;
assign w1835 = ~pi0440 & pi0442;
assign w1836 = ~w1834 & ~w1835;
assign w1837 = ~w1833 & ~w1836;
assign w1838 = ~w1830 & ~w1837;
assign w1839 = pi0369 & w1838;
assign w1840 = ~pi0369 & ~w1838;
assign w1841 = ~w1839 & ~w1840;
assign w1842 = ~pi0370 & ~pi0371;
assign w1843 = pi0370 & pi0371;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = ~w1841 & ~w1844;
assign w1846 = pi0369 & ~w1838;
assign w1847 = ~pi0369 & w1838;
assign w1848 = ~w1846 & ~w1847;
assign w1849 = pi0370 & ~pi0371;
assign w1850 = ~pi0370 & pi0371;
assign w1851 = ~w1849 & ~w1850;
assign w1852 = ~w1848 & ~w1851;
assign w1853 = ~w1845 & ~w1852;
assign w1854 = pi1198 & ~w1853;
assign w1855 = ~w1811 & ~w1854;
assign w1856 = w1768 & w1855;
assign w1857 = ~pi0590 & pi0591;
assign w1858 = ~pi0591 & ~pi0592;
assign w1859 = ~pi0590 & ~w1858;
assign w1860 = (~w1856 & w1857) | (~w1856 & w1859) | (w1857 & w1859);
assign w1861 = ~pi0344 & pi0345;
assign w1862 = pi0344 & ~pi0345;
assign w1863 = ~w1861 & ~w1862;
assign w1864 = ~pi0346 & ~pi0358;
assign w1865 = pi0346 & pi0358;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = ~w1863 & ~w1866;
assign w1868 = pi0346 & ~pi0358;
assign w1869 = ~pi0346 & pi0358;
assign w1870 = ~w1868 & ~w1869;
assign w1871 = pi0344 & pi0345;
assign w1872 = ~pi0344 & ~pi0345;
assign w1873 = ~w1871 & ~w1872;
assign w1874 = ~w1870 & ~w1873;
assign w1875 = ~w1867 & ~w1874;
assign w1876 = pi0362 & pi0450;
assign w1877 = ~pi0362 & ~pi0450;
assign w1878 = ~w1876 & ~w1877;
assign w1879 = ~w1875 & ~w1878;
assign w1880 = ~w1863 & ~w1870;
assign w1881 = ~w1866 & ~w1873;
assign w1882 = ~w1880 & ~w1881;
assign w1883 = pi0362 & ~pi0450;
assign w1884 = ~pi0362 & pi0450;
assign w1885 = ~w1883 & ~w1884;
assign w1886 = ~w1882 & ~w1885;
assign w1887 = ~w1879 & ~w1886;
assign w1888 = ~pi0323 & ~w1887;
assign w1889 = pi0323 & w1887;
assign w1890 = ~w1888 & ~w1889;
assign w1891 = pi0327 & ~pi0343;
assign w1892 = ~pi0327 & pi0343;
assign w1893 = ~w1891 & ~w1892;
assign w1894 = pi1197 & w1893;
assign w1895 = (pi1197 & w1890) | (pi1197 & w1894) | (w1890 & w1894);
assign w1896 = pi0323 & ~w1887;
assign w1897 = ~pi0323 & w1887;
assign w1898 = ~w1896 & ~w1897;
assign w1899 = pi0327 & pi0343;
assign w1900 = ~pi0327 & ~pi0343;
assign w1901 = ~w1899 & ~w1900;
assign w1902 = ~w1898 & ~w1901;
assign w1903 = w1895 & ~w1902;
assign w1904 = ~pi0354 & pi0356;
assign w1905 = pi0354 & ~pi0356;
assign w1906 = ~w1904 & ~w1905;
assign w1907 = ~pi0357 & ~pi0360;
assign w1908 = pi0357 & pi0360;
assign w1909 = ~w1907 & ~w1908;
assign w1910 = ~w1906 & ~w1909;
assign w1911 = pi0357 & ~pi0360;
assign w1912 = ~pi0357 & pi0360;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = pi0354 & pi0356;
assign w1915 = ~pi0354 & ~pi0356;
assign w1916 = ~w1914 & ~w1915;
assign w1917 = ~w1913 & ~w1916;
assign w1918 = ~w1910 & ~w1917;
assign w1919 = pi0461 & pi0462;
assign w1920 = ~pi0461 & ~pi0462;
assign w1921 = ~w1919 & ~w1920;
assign w1922 = ~w1918 & ~w1921;
assign w1923 = ~w1906 & ~w1913;
assign w1924 = ~w1909 & ~w1916;
assign w1925 = ~w1923 & ~w1924;
assign w1926 = pi0461 & ~pi0462;
assign w1927 = ~pi0461 & pi0462;
assign w1928 = ~w1926 & ~w1927;
assign w1929 = ~w1925 & ~w1928;
assign w1930 = ~w1922 & ~w1929;
assign w1931 = pi0351 & w1930;
assign w1932 = ~pi0351 & ~w1930;
assign w1933 = ~w1931 & ~w1932;
assign w1934 = ~pi0352 & ~pi0353;
assign w1935 = pi0352 & pi0353;
assign w1936 = ~w1934 & ~w1935;
assign w1937 = ~w1933 & ~w1936;
assign w1938 = pi0351 & ~w1930;
assign w1939 = ~pi0351 & w1930;
assign w1940 = ~w1938 & ~w1939;
assign w1941 = pi0352 & ~pi0353;
assign w1942 = ~pi0352 & pi0353;
assign w1943 = ~w1941 & ~w1942;
assign w1944 = ~w1940 & ~w1943;
assign w1945 = ~w1937 & ~w1944;
assign w1946 = pi1199 & ~w1945;
assign w1947 = ~w1903 & ~w1946;
assign w1948 = ~pi0361 & pi0441;
assign w1949 = pi0361 & ~pi0441;
assign w1950 = ~w1948 & ~w1949;
assign w1951 = ~pi0452 & ~pi0455;
assign w1952 = pi0452 & pi0455;
assign w1953 = ~w1951 & ~w1952;
assign w1954 = ~w1950 & ~w1953;
assign w1955 = pi0452 & ~pi0455;
assign w1956 = ~pi0452 & pi0455;
assign w1957 = ~w1955 & ~w1956;
assign w1958 = pi0361 & pi0441;
assign w1959 = ~pi0361 & ~pi0441;
assign w1960 = ~w1958 & ~w1959;
assign w1961 = ~w1957 & ~w1960;
assign w1962 = ~w1954 & ~w1961;
assign w1963 = pi0458 & pi0460;
assign w1964 = ~pi0458 & ~pi0460;
assign w1965 = ~w1963 & ~w1964;
assign w1966 = ~w1962 & ~w1965;
assign w1967 = ~w1950 & ~w1957;
assign w1968 = ~w1953 & ~w1960;
assign w1969 = ~w1967 & ~w1968;
assign w1970 = pi0458 & ~pi0460;
assign w1971 = ~pi0458 & pi0460;
assign w1972 = ~w1970 & ~w1971;
assign w1973 = ~w1969 & ~w1972;
assign w1974 = ~w1966 & ~w1973;
assign w1975 = ~pi0320 & ~w1974;
assign w1976 = pi0320 & w1974;
assign w1977 = ~w1975 & ~w1976;
assign w1978 = pi0342 & ~pi0355;
assign w1979 = ~pi0342 & pi0355;
assign w1980 = ~w1978 & ~w1979;
assign w1981 = pi1196 & w1980;
assign w1982 = (pi1196 & w1977) | (pi1196 & w1981) | (w1977 & w1981);
assign w1983 = pi0320 & ~w1974;
assign w1984 = ~pi0320 & w1974;
assign w1985 = ~w1983 & ~w1984;
assign w1986 = pi0342 & pi0355;
assign w1987 = ~pi0342 & ~pi0355;
assign w1988 = ~w1986 & ~w1987;
assign w1989 = ~w1985 & ~w1988;
assign w1990 = w1982 & ~w1989;
assign w1991 = ~pi0322 & pi0347;
assign w1992 = pi0322 & ~pi0347;
assign w1993 = ~w1991 & ~w1992;
assign w1994 = ~pi0348 & ~pi0349;
assign w1995 = pi0348 & pi0349;
assign w1996 = ~w1994 & ~w1995;
assign w1997 = ~w1993 & ~w1996;
assign w1998 = pi0348 & ~pi0349;
assign w1999 = ~pi0348 & pi0349;
assign w2000 = ~w1998 & ~w1999;
assign w2001 = pi0322 & pi0347;
assign w2002 = ~pi0322 & ~pi0347;
assign w2003 = ~w2001 & ~w2002;
assign w2004 = ~w2000 & ~w2003;
assign w2005 = ~w1997 & ~w2004;
assign w2006 = pi0350 & pi0359;
assign w2007 = ~pi0350 & ~pi0359;
assign w2008 = ~w2006 & ~w2007;
assign w2009 = ~w2005 & ~w2008;
assign w2010 = ~w1993 & ~w2000;
assign w2011 = ~w1996 & ~w2003;
assign w2012 = ~w2010 & ~w2011;
assign w2013 = pi0350 & ~pi0359;
assign w2014 = ~pi0350 & pi0359;
assign w2015 = ~w2013 & ~w2014;
assign w2016 = ~w2012 & ~w2015;
assign w2017 = ~w2009 & ~w2016;
assign w2018 = pi0315 & w2017;
assign w2019 = ~pi0315 & ~w2017;
assign w2020 = ~w2018 & ~w2019;
assign w2021 = ~pi0316 & ~pi0321;
assign w2022 = pi0316 & pi0321;
assign w2023 = ~w2021 & ~w2022;
assign w2024 = ~w2020 & ~w2023;
assign w2025 = pi0315 & ~w2017;
assign w2026 = ~pi0315 & w2017;
assign w2027 = ~w2025 & ~w2026;
assign w2028 = pi0316 & ~pi0321;
assign w2029 = ~pi0316 & pi0321;
assign w2030 = ~w2028 & ~w2029;
assign w2031 = ~w2027 & ~w2030;
assign w2032 = ~w2024 & ~w2031;
assign w2033 = pi1198 & ~w2032;
assign w2034 = ~w1990 & ~w2033;
assign w2035 = w1947 & w2034;
assign w2036 = pi0590 & w1858;
assign w2037 = ~w2035 & w2036;
assign w2038 = ~w1860 & ~w2037;
assign w2039 = ~pi0122 & ~pi1091;
assign w2040 = w1476 & w2039;
assign w2041 = ~pi0285 & ~pi0286;
assign w2042 = ~pi0288 & ~pi0289;
assign w2043 = w2041 & w2042;
assign w2044 = ~pi1161 & ~pi1162;
assign w2045 = ~pi1163 & w2044;
assign w2046 = ~w2043 & w2045;
assign w2047 = w2040 & w2046;
assign w2048 = ~pi0098 & pi0567;
assign w2049 = w2047 & w2048;
assign w2050 = ~pi0397 & pi0404;
assign w2051 = pi0397 & ~pi0404;
assign w2052 = ~w2050 & ~w2051;
assign w2053 = ~pi0410 & ~pi0411;
assign w2054 = pi0410 & pi0411;
assign w2055 = ~w2053 & ~w2054;
assign w2056 = ~w2052 & ~w2055;
assign w2057 = pi0410 & ~pi0411;
assign w2058 = ~pi0410 & pi0411;
assign w2059 = ~w2057 & ~w2058;
assign w2060 = pi0397 & pi0404;
assign w2061 = ~pi0397 & ~pi0404;
assign w2062 = ~w2060 & ~w2061;
assign w2063 = ~w2059 & ~w2062;
assign w2064 = ~w2056 & ~w2063;
assign w2065 = pi0412 & pi0456;
assign w2066 = ~pi0412 & ~pi0456;
assign w2067 = ~w2065 & ~w2066;
assign w2068 = ~w2064 & ~w2067;
assign w2069 = ~w2052 & ~w2059;
assign w2070 = ~w2055 & ~w2062;
assign w2071 = ~w2069 & ~w2070;
assign w2072 = pi0412 & ~pi0456;
assign w2073 = ~pi0412 & pi0456;
assign w2074 = ~w2072 & ~w2073;
assign w2075 = ~w2071 & ~w2074;
assign w2076 = ~w2068 & ~w2075;
assign w2077 = pi0319 & w2076;
assign w2078 = ~pi0319 & ~w2076;
assign w2079 = ~w2077 & ~w2078;
assign w2080 = ~pi0324 & ~pi0390;
assign w2081 = pi0324 & pi0390;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = ~w2079 & ~w2082;
assign w2084 = pi0319 & ~w2076;
assign w2085 = ~pi0319 & w2076;
assign w2086 = ~w2084 & ~w2085;
assign w2087 = pi0324 & ~pi0390;
assign w2088 = ~pi0324 & pi0390;
assign w2089 = ~w2087 & ~w2088;
assign w2090 = ~w2086 & ~w2089;
assign w2091 = ~w2083 & ~w2090;
assign w2092 = pi1196 & ~w2091;
assign w2093 = ~pi0401 & pi0402;
assign w2094 = pi0401 & ~pi0402;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = ~pi0403 & ~pi0405;
assign w2097 = pi0403 & pi0405;
assign w2098 = ~w2096 & ~w2097;
assign w2099 = ~w2095 & ~w2098;
assign w2100 = pi0403 & ~pi0405;
assign w2101 = ~pi0403 & pi0405;
assign w2102 = ~w2100 & ~w2101;
assign w2103 = pi0401 & pi0402;
assign w2104 = ~pi0401 & ~pi0402;
assign w2105 = ~w2103 & ~w2104;
assign w2106 = ~w2102 & ~w2105;
assign w2107 = ~w2099 & ~w2106;
assign w2108 = pi0406 & pi0409;
assign w2109 = ~pi0406 & ~pi0409;
assign w2110 = ~w2108 & ~w2109;
assign w2111 = ~w2107 & ~w2110;
assign w2112 = ~w2095 & ~w2102;
assign w2113 = ~w2098 & ~w2105;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = pi0406 & ~pi0409;
assign w2116 = ~pi0406 & pi0409;
assign w2117 = ~w2115 & ~w2116;
assign w2118 = ~w2114 & ~w2117;
assign w2119 = ~w2111 & ~w2118;
assign w2120 = pi0318 & w2119;
assign w2121 = ~pi0318 & ~w2119;
assign w2122 = ~w2120 & ~w2121;
assign w2123 = ~pi0325 & ~pi0326;
assign w2124 = pi0325 & pi0326;
assign w2125 = ~w2123 & ~w2124;
assign w2126 = ~w2122 & ~w2125;
assign w2127 = pi0318 & ~w2119;
assign w2128 = ~pi0318 & w2119;
assign w2129 = ~w2127 & ~w2128;
assign w2130 = pi0325 & ~pi0326;
assign w2131 = ~pi0325 & pi0326;
assign w2132 = ~w2130 & ~w2131;
assign w2133 = ~w2129 & ~w2132;
assign w2134 = ~w2126 & ~w2133;
assign w2135 = pi1199 & ~w2134;
assign w2136 = ~w2092 & ~w2135;
assign w2137 = ~pi0391 & pi0392;
assign w2138 = pi0391 & ~pi0392;
assign w2139 = ~w2137 & ~w2138;
assign w2140 = ~pi0393 & ~pi0407;
assign w2141 = pi0393 & pi0407;
assign w2142 = ~w2140 & ~w2141;
assign w2143 = ~w2139 & ~w2142;
assign w2144 = pi0393 & ~pi0407;
assign w2145 = ~pi0393 & pi0407;
assign w2146 = ~w2144 & ~w2145;
assign w2147 = pi0391 & pi0392;
assign w2148 = ~pi0391 & ~pi0392;
assign w2149 = ~w2147 & ~w2148;
assign w2150 = ~w2146 & ~w2149;
assign w2151 = ~w2143 & ~w2150;
assign w2152 = pi0413 & pi0463;
assign w2153 = ~pi0413 & ~pi0463;
assign w2154 = ~w2152 & ~w2153;
assign w2155 = ~w2151 & ~w2154;
assign w2156 = ~w2139 & ~w2146;
assign w2157 = ~w2142 & ~w2149;
assign w2158 = ~w2156 & ~w2157;
assign w2159 = pi0413 & ~pi0463;
assign w2160 = ~pi0413 & pi0463;
assign w2161 = ~w2159 & ~w2160;
assign w2162 = ~w2158 & ~w2161;
assign w2163 = ~w2155 & ~w2162;
assign w2164 = pi0333 & w2163;
assign w2165 = ~pi0333 & ~w2163;
assign w2166 = ~w2164 & ~w2165;
assign w2167 = ~pi0334 & ~pi0335;
assign w2168 = pi0334 & pi0335;
assign w2169 = ~w2167 & ~w2168;
assign w2170 = ~w2166 & ~w2169;
assign w2171 = pi0333 & ~w2163;
assign w2172 = ~pi0333 & w2163;
assign w2173 = ~w2171 & ~w2172;
assign w2174 = pi0334 & ~pi0335;
assign w2175 = ~pi0334 & pi0335;
assign w2176 = ~w2174 & ~w2175;
assign w2177 = ~w2173 & ~w2176;
assign w2178 = ~w2170 & ~w2177;
assign w2179 = pi1197 & ~w2178;
assign w2180 = ~pi0395 & pi0396;
assign w2181 = pi0395 & ~pi0396;
assign w2182 = ~w2180 & ~w2181;
assign w2183 = ~pi0398 & ~pi0399;
assign w2184 = pi0398 & pi0399;
assign w2185 = ~w2183 & ~w2184;
assign w2186 = ~w2182 & ~w2185;
assign w2187 = pi0398 & ~pi0399;
assign w2188 = ~pi0398 & pi0399;
assign w2189 = ~w2187 & ~w2188;
assign w2190 = pi0395 & pi0396;
assign w2191 = ~pi0395 & ~pi0396;
assign w2192 = ~w2190 & ~w2191;
assign w2193 = ~w2189 & ~w2192;
assign w2194 = ~w2186 & ~w2193;
assign w2195 = pi0400 & pi0408;
assign w2196 = ~pi0400 & ~pi0408;
assign w2197 = ~w2195 & ~w2196;
assign w2198 = ~w2194 & ~w2197;
assign w2199 = ~w2182 & ~w2189;
assign w2200 = ~w2185 & ~w2192;
assign w2201 = ~w2199 & ~w2200;
assign w2202 = pi0400 & ~pi0408;
assign w2203 = ~pi0400 & pi0408;
assign w2204 = ~w2202 & ~w2203;
assign w2205 = ~w2201 & ~w2204;
assign w2206 = ~w2198 & ~w2205;
assign w2207 = pi0328 & w2206;
assign w2208 = ~pi0328 & ~w2206;
assign w2209 = ~w2207 & ~w2208;
assign w2210 = ~pi0329 & ~pi0394;
assign w2211 = pi0329 & pi0394;
assign w2212 = ~w2210 & ~w2211;
assign w2213 = ~w2209 & ~w2212;
assign w2214 = pi0328 & ~w2206;
assign w2215 = ~pi0328 & w2206;
assign w2216 = ~w2214 & ~w2215;
assign w2217 = pi0329 & ~pi0394;
assign w2218 = ~pi0329 & pi0394;
assign w2219 = ~w2217 & ~w2218;
assign w2220 = ~w2216 & ~w2219;
assign w2221 = ~w2213 & ~w2220;
assign w2222 = pi1198 & ~w2221;
assign w2223 = ~w2179 & ~w2222;
assign w2224 = w2136 & w2223;
assign w2225 = ~pi0217 & ~pi0591;
assign w2226 = w2048 & ~w2225;
assign w2227 = w2047 & w2226;
assign w2228 = pi0591 & pi0592;
assign w2229 = ~pi0217 & ~w2228;
assign w2230 = w2048 & ~w2229;
assign w2231 = w2047 & w2230;
assign w2232 = (w2224 & w2227) | (w2224 & w2231) | (w2227 & w2231);
assign w2233 = ~pi0418 & pi0431;
assign w2234 = pi0418 & ~pi0431;
assign w2235 = ~w2233 & ~w2234;
assign w2236 = ~pi0437 & ~pi0438;
assign w2237 = pi0437 & pi0438;
assign w2238 = ~w2236 & ~w2237;
assign w2239 = ~w2235 & ~w2238;
assign w2240 = pi0437 & ~pi0438;
assign w2241 = ~pi0437 & pi0438;
assign w2242 = ~w2240 & ~w2241;
assign w2243 = pi0418 & pi0431;
assign w2244 = ~pi0418 & ~pi0431;
assign w2245 = ~w2243 & ~w2244;
assign w2246 = ~w2242 & ~w2245;
assign w2247 = ~w2239 & ~w2246;
assign w2248 = pi0453 & pi0464;
assign w2249 = ~pi0453 & ~pi0464;
assign w2250 = ~w2248 & ~w2249;
assign w2251 = ~w2247 & ~w2250;
assign w2252 = ~w2235 & ~w2242;
assign w2253 = ~w2238 & ~w2245;
assign w2254 = ~w2252 & ~w2253;
assign w2255 = pi0453 & ~pi0464;
assign w2256 = ~pi0453 & pi0464;
assign w2257 = ~w2255 & ~w2256;
assign w2258 = ~w2254 & ~w2257;
assign w2259 = ~w2251 & ~w2258;
assign w2260 = pi0415 & w2259;
assign w2261 = ~pi0415 & ~w2259;
assign w2262 = ~w2260 & ~w2261;
assign w2263 = ~pi0416 & ~pi0417;
assign w2264 = pi0416 & pi0417;
assign w2265 = ~w2263 & ~w2264;
assign w2266 = ~w2262 & ~w2265;
assign w2267 = pi0415 & ~w2259;
assign w2268 = ~pi0415 & w2259;
assign w2269 = ~w2267 & ~w2268;
assign w2270 = pi0416 & ~pi0417;
assign w2271 = ~pi0416 & pi0417;
assign w2272 = ~w2270 & ~w2271;
assign w2273 = ~w2269 & ~w2272;
assign w2274 = ~w2266 & ~w2273;
assign w2275 = pi1197 & ~w2274;
assign w2276 = ~pi0423 & pi0424;
assign w2277 = pi0423 & ~pi0424;
assign w2278 = ~w2276 & ~w2277;
assign w2279 = ~pi0425 & ~pi0432;
assign w2280 = pi0425 & pi0432;
assign w2281 = ~w2279 & ~w2280;
assign w2282 = ~w2278 & ~w2281;
assign w2283 = pi0425 & ~pi0432;
assign w2284 = ~pi0425 & pi0432;
assign w2285 = ~w2283 & ~w2284;
assign w2286 = pi0423 & pi0424;
assign w2287 = ~pi0423 & ~pi0424;
assign w2288 = ~w2286 & ~w2287;
assign w2289 = ~w2285 & ~w2288;
assign w2290 = ~w2282 & ~w2289;
assign w2291 = pi0454 & pi0459;
assign w2292 = ~pi0454 & ~pi0459;
assign w2293 = ~w2291 & ~w2292;
assign w2294 = ~w2290 & ~w2293;
assign w2295 = ~w2278 & ~w2285;
assign w2296 = ~w2281 & ~w2288;
assign w2297 = ~w2295 & ~w2296;
assign w2298 = pi0454 & ~pi0459;
assign w2299 = ~pi0454 & pi0459;
assign w2300 = ~w2298 & ~w2299;
assign w2301 = ~w2297 & ~w2300;
assign w2302 = ~w2294 & ~w2301;
assign w2303 = pi0419 & w2302;
assign w2304 = ~pi0419 & ~w2302;
assign w2305 = ~w2303 & ~w2304;
assign w2306 = ~pi0420 & ~pi0421;
assign w2307 = pi0420 & pi0421;
assign w2308 = ~w2306 & ~w2307;
assign w2309 = ~w2305 & ~w2308;
assign w2310 = pi0419 & ~w2302;
assign w2311 = ~pi0419 & w2302;
assign w2312 = ~w2310 & ~w2311;
assign w2313 = pi0420 & ~pi0421;
assign w2314 = ~pi0420 & pi0421;
assign w2315 = ~w2313 & ~w2314;
assign w2316 = ~w2312 & ~w2315;
assign w2317 = ~w2309 & ~w2316;
assign w2318 = pi1198 & ~w2317;
assign w2319 = ~w2275 & ~w2318;
assign w2320 = ~pi0434 & pi0435;
assign w2321 = pi0434 & ~pi0435;
assign w2322 = ~w2320 & ~w2321;
assign w2323 = ~pi0436 & ~pi0443;
assign w2324 = pi0436 & pi0443;
assign w2325 = ~w2323 & ~w2324;
assign w2326 = ~w2322 & ~w2325;
assign w2327 = pi0436 & ~pi0443;
assign w2328 = ~pi0436 & pi0443;
assign w2329 = ~w2327 & ~w2328;
assign w2330 = pi0434 & pi0435;
assign w2331 = ~pi0434 & ~pi0435;
assign w2332 = ~w2330 & ~w2331;
assign w2333 = ~w2329 & ~w2332;
assign w2334 = ~w2326 & ~w2333;
assign w2335 = pi0444 & pi0446;
assign w2336 = ~pi0444 & ~pi0446;
assign w2337 = ~w2335 & ~w2336;
assign w2338 = ~w2334 & ~w2337;
assign w2339 = ~w2322 & ~w2329;
assign w2340 = ~w2325 & ~w2332;
assign w2341 = ~w2339 & ~w2340;
assign w2342 = pi0444 & ~pi0446;
assign w2343 = ~pi0444 & pi0446;
assign w2344 = ~w2342 & ~w2343;
assign w2345 = ~w2341 & ~w2344;
assign w2346 = ~w2338 & ~w2345;
assign w2347 = pi0414 & w2346;
assign w2348 = ~pi0414 & ~w2346;
assign w2349 = ~w2347 & ~w2348;
assign w2350 = ~pi0422 & ~pi0429;
assign w2351 = pi0422 & pi0429;
assign w2352 = ~w2350 & ~w2351;
assign w2353 = ~w2349 & ~w2352;
assign w2354 = pi0414 & ~w2346;
assign w2355 = ~pi0414 & w2346;
assign w2356 = ~w2354 & ~w2355;
assign w2357 = pi0422 & ~pi0429;
assign w2358 = ~pi0422 & pi0429;
assign w2359 = ~w2357 & ~w2358;
assign w2360 = ~w2356 & ~w2359;
assign w2361 = ~w2353 & ~w2360;
assign w2362 = pi1196 & ~w2361;
assign w2363 = ~pi0430 & pi0433;
assign w2364 = pi0430 & ~pi0433;
assign w2365 = ~w2363 & ~w2364;
assign w2366 = ~pi0445 & ~pi0448;
assign w2367 = pi0445 & pi0448;
assign w2368 = ~w2366 & ~w2367;
assign w2369 = ~w2365 & ~w2368;
assign w2370 = pi0445 & ~pi0448;
assign w2371 = ~pi0445 & pi0448;
assign w2372 = ~w2370 & ~w2371;
assign w2373 = pi0430 & pi0433;
assign w2374 = ~pi0430 & ~pi0433;
assign w2375 = ~w2373 & ~w2374;
assign w2376 = ~w2372 & ~w2375;
assign w2377 = ~w2369 & ~w2376;
assign w2378 = pi0449 & pi0451;
assign w2379 = ~pi0449 & ~pi0451;
assign w2380 = ~w2378 & ~w2379;
assign w2381 = ~w2377 & ~w2380;
assign w2382 = ~w2365 & ~w2372;
assign w2383 = ~w2368 & ~w2375;
assign w2384 = ~w2382 & ~w2383;
assign w2385 = pi0449 & ~pi0451;
assign w2386 = ~pi0449 & pi0451;
assign w2387 = ~w2385 & ~w2386;
assign w2388 = ~w2384 & ~w2387;
assign w2389 = ~w2381 & ~w2388;
assign w2390 = pi0426 & w2389;
assign w2391 = ~pi0426 & ~w2389;
assign w2392 = ~w2390 & ~w2391;
assign w2393 = ~pi0427 & ~pi0428;
assign w2394 = pi0427 & pi0428;
assign w2395 = ~w2393 & ~w2394;
assign w2396 = ~w2392 & ~w2395;
assign w2397 = pi0426 & ~w2389;
assign w2398 = ~pi0426 & w2389;
assign w2399 = ~w2397 & ~w2398;
assign w2400 = pi0427 & ~pi0428;
assign w2401 = ~pi0427 & pi0428;
assign w2402 = ~w2400 & ~w2401;
assign w2403 = ~w2399 & ~w2402;
assign w2404 = ~w2396 & ~w2403;
assign w2405 = pi1199 & ~w2404;
assign w2406 = ~w2362 & ~w2405;
assign w2407 = w2319 & w2406;
assign w2408 = ~pi0590 & ~pi0591;
assign w2409 = pi0588 & ~pi0592;
assign w2410 = w2408 & w2409;
assign w2411 = pi0588 & ~w2410;
assign w2412 = (pi0588 & w2407) | (pi0588 & w2411) | (w2407 & w2411);
assign w2413 = (w2049 & w2232) | (w2049 & w2412) | (w2232 & w2412);
assign w2414 = ~w2407 & w2410;
assign w2415 = (w2049 & w2232) | (w2049 & ~w2414) | (w2232 & ~w2414);
assign w2416 = (w2038 & w2413) | (w2038 & w2415) | (w2413 & w2415);
assign w2417 = ~pi0031 & pi1161;
assign w2418 = w1475 & w2417;
assign w2419 = pi1162 & ~pi1163;
assign w2420 = w2418 & w2419;
assign w2421 = ~w2416 & ~w2420;
assign w2422 = w450 & w2225;
assign w2423 = w450 & w2229;
assign w2424 = (~w2224 & w2422) | (~w2224 & w2423) | (w2422 & w2423);
assign w2425 = ~w2412 & w2424;
assign w2426 = w2414 & w2424;
assign w2427 = (~w2038 & w2425) | (~w2038 & w2426) | (w2425 & w2426);
assign w2428 = ~pi1091 & w1475;
assign w2429 = pi0098 & w106;
assign w2430 = w382 & w2429;
assign w2431 = w359 & w2430;
assign w2432 = w244 & w2431;
assign w2433 = ~w234 & w2432;
assign w2434 = pi0090 & ~pi0093;
assign w2435 = ~pi0090 & pi0093;
assign w2436 = ~w2434 & ~w2435;
assign w2437 = ~pi0051 & ~pi0841;
assign w2438 = ~w2436 & w2437;
assign w2439 = ~pi0035 & pi0051;
assign w2440 = w428 & w2439;
assign w2441 = ~pi0070 & w2440;
assign w2442 = (w1637 & w2438) | (w1637 & w2441) | (w2438 & w2441);
assign w2443 = w99 & w2442;
assign w2444 = ~pi0096 & ~w2443;
assign w2445 = (~pi0096 & ~w112) | (~pi0096 & w2444) | (~w112 & w2444);
assign w2446 = ~w2428 & ~w2445;
assign w2447 = (~w2428 & w2433) | (~w2428 & w2446) | (w2433 & w2446);
assign w2448 = ~pi0072 & ~w1283;
assign w2449 = w1281 & w2448;
assign w2450 = w2447 & w2449;
assign w2451 = ~pi0122 & w1236;
assign w2452 = pi0097 & w354;
assign w2453 = w353 & w2452;
assign w2454 = w429 & w2453;
assign w2455 = w2451 & w2454;
assign w2456 = w429 & w2451;
assign w2457 = (~pi0109 & w238) | (~pi0109 & w241) | (w238 & w241);
assign w2458 = ~pi0024 & ~pi0046;
assign w2459 = w351 & w2458;
assign w2460 = pi0091 & ~pi0110;
assign w2461 = w2459 & w2460;
assign w2462 = ~w2453 & ~w2461;
assign w2463 = (~w2453 & ~w2457) | (~w2453 & w2462) | (~w2457 & w2462);
assign w2464 = w2456 & ~w2463;
assign w2465 = (w465 & w2455) | (w465 & w2464) | (w2455 & w2464);
assign w2466 = w2457 & w2461;
assign w2467 = w2456 & w2466;
assign w2468 = w465 & w2467;
assign w2469 = (w254 & w2465) | (w254 & w2468) | (w2465 & w2468);
assign w2470 = ~w2450 & ~w2469;
assign w2471 = ~pi0116 & w1312;
assign w2472 = ~pi0052 & ~pi0113;
assign w2473 = w1317 & w2472;
assign w2474 = w2471 & w2473;
assign w2475 = ~pi0152 & ~pi0161;
assign w2476 = ~pi0166 & pi0299;
assign w2477 = w2475 & w2476;
assign w2478 = ~pi0144 & ~pi0174;
assign w2479 = ~pi0189 & ~pi0299;
assign w2480 = w2478 & w2479;
assign w2481 = ~w2477 & ~w2480;
assign w2482 = pi0232 & ~pi0332;
assign w2483 = ~pi0468 & w2482;
assign w2484 = ~w2481 & w2483;
assign w2485 = ~w2474 & ~w2484;
assign w2486 = ~pi0087 & pi0252;
assign w2487 = ~pi0024 & ~pi0100;
assign w2488 = w2486 & w2487;
assign w2489 = ~pi0122 & w2488;
assign w2490 = w1236 & w2489;
assign w2491 = ~w147 & ~w2490;
assign w2492 = (~w147 & ~w2485) | (~w147 & w2491) | (~w2485 & w2491);
assign w2493 = w1284 & ~w2492;
assign w2494 = w113 & w2493;
assign w2495 = w117 & ~w169;
assign w2496 = w1302 & w2495;
assign w2497 = w2494 & w2496;
assign w2498 = w4 & w109;
assign w2499 = w112 & w2498;
assign w2500 = ~pi0100 & w1658;
assign w2501 = ~w1 & ~w2500;
assign w2502 = (~w5 & ~w2500) | (~w5 & w2501) | (~w2500 & w2501);
assign w2503 = ~pi0122 & pi0228;
assign w2504 = pi0100 & ~w2503;
assign w2505 = w1658 & ~w2504;
assign w2506 = (w1236 & w2500) | (w1236 & w2505) | (w2500 & w2505);
assign w2507 = ~w6 & ~w2506;
assign w2508 = (~w2485 & w2502) | (~w2485 & w2507) | (w2502 & w2507);
assign w2509 = (~w6 & ~w2499) | (~w6 & w2508) | (~w2499 & w2508);
assign w2510 = ~pi0222 & ~pi0224;
assign w2511 = w1290 & ~w2510;
assign w2512 = w1268 & w2511;
assign w2513 = w1255 & ~w2511;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = pi0039 & w1470;
assign w2516 = (pi0039 & ~w1237) | (pi0039 & w2515) | (~w1237 & w2515);
assign w2517 = (pi0039 & w2514) | (pi0039 & w2516) | (w2514 & w2516);
assign w2518 = ~w2509 & ~w2517;
assign w2519 = pi0039 & pi0100;
assign w2520 = pi0087 & ~w1283;
assign w2521 = w1281 & w2520;
assign w2522 = ~pi0039 & ~pi0100;
assign w2523 = ~w2519 & ~w2522;
assign w2524 = (~w2519 & w2521) | (~w2519 & w2523) | (w2521 & w2523);
assign w2525 = ~pi0039 & ~pi0072;
assign w2526 = ~pi1091 & w2525;
assign w2527 = w1476 & w2526;
assign w2528 = w1641 & w2527;
assign w2529 = w2442 & w2528;
assign w2530 = ~w2524 & ~w2529;
assign w2531 = (~w492 & ~w2524) | (~w492 & w2530) | (~w2524 & w2530);
assign w2532 = ~pi0093 & w186;
assign w2533 = ~pi0095 & ~pi0122;
assign w2534 = w347 & w2533;
assign w2535 = pi0829 & ~pi0841;
assign w2536 = w2534 & w2535;
assign w2537 = w2532 & w2536;
assign w2538 = ~w1641 & ~w2537;
assign w2539 = (~w492 & ~w1641) | (~w492 & w2538) | (~w1641 & w2538);
assign w2540 = w2531 & w2539;
assign w2541 = w2518 & ~w2540;
assign w2542 = ~w2497 & ~w2541;
assign w2543 = w2518 & ~w2531;
assign w2544 = ~w2497 & ~w2543;
assign w2545 = (w2470 & w2542) | (w2470 & w2544) | (w2542 & w2544);
assign w2546 = w1475 & ~w2048;
assign w2547 = w2045 & ~w2546;
assign w2548 = w529 & w2547;
assign w2549 = ~w2545 & w2548;
assign w2550 = ~w2427 & w2549;
assign w2551 = w2421 & ~w2550;
assign w2552 = ~w377 & w407;
assign w2553 = (w346 & w407) | (w346 & w2552) | (w407 & w2552);
assign w2554 = w594 & ~w2553;
assign w2555 = ~pi0024 & pi0050;
assign w2556 = ~w454 & ~w2043;
assign w2557 = ~pi0137 & ~w2556;
assign w2558 = pi0076 & w2557;
assign w2559 = w413 & w2558;
assign w2560 = ~pi0050 & w2559;
assign w2561 = ~w2555 & ~w2560;
assign w2562 = pi0024 & w413;
assign w2563 = ~pi0841 & ~w2562;
assign w2564 = pi0032 & ~w2563;
assign w2565 = w2561 & ~w2564;
assign w2566 = w2554 & ~w2565;
assign w2567 = w134 & ~w2485;
assign w2568 = pi0950 & w1322;
assign w2569 = ~pi0299 & w129;
assign w2570 = pi0299 & w38;
assign w2571 = ~w2569 & ~w2570;
assign w2572 = ~pi0250 & ~w2571;
assign w2573 = ~w2568 & w2572;
assign w2574 = pi0250 & ~w2571;
assign w2575 = pi0252 & w2571;
assign w2576 = ~w2574 & ~w2575;
assign w2577 = pi0129 & ~w2576;
assign w2578 = ~w2573 & ~w2577;
assign w2579 = w2567 & ~w2578;
assign w2580 = pi0252 & ~w2485;
assign w2581 = w2487 & ~w2580;
assign w2582 = pi0075 & w2581;
assign w2583 = ~w454 & w2582;
assign w2584 = ~w1320 & w2583;
assign w2585 = ~w2579 & ~w2584;
assign w2586 = ~pi0137 & ~w2585;
assign w2587 = w1622 & w2586;
assign w2588 = ~w2566 & ~w2587;
assign w2589 = pi0073 & pi0299;
assign w2590 = ~pi0152 & w2589;
assign w2591 = ~pi0210 & ~pi0841;
assign w2592 = pi0032 & w2591;
assign w2593 = ~pi0050 & ~pi0070;
assign w2594 = w443 & w2593;
assign w2595 = ~w2592 & w2594;
assign w2596 = ~pi0073 & pi0149;
assign w2597 = pi0299 & w2596;
assign w2598 = ~w2590 & ~w2597;
assign w2599 = (~w2590 & w2595) | (~w2590 & w2598) | (w2595 & w2598);
assign w2600 = ~pi0198 & ~pi0841;
assign w2601 = pi0032 & w2600;
assign w2602 = w2594 & ~w2601;
assign w2603 = pi0183 & ~pi0299;
assign w2604 = ~w2602 & w2603;
assign w2605 = w2599 & ~w2604;
assign w2606 = w594 & ~w2605;
assign w2607 = ~w2553 & w2606;
assign w2608 = pi0073 & w377;
assign w2609 = ~pi0174 & ~pi0299;
assign w2610 = w2608 & w2609;
assign w2611 = ~w346 & w2610;
assign w2612 = pi0193 & ~pi0299;
assign w2613 = pi0172 & pi0299;
assign w2614 = ~w2612 & ~w2613;
assign w2615 = ~pi0058 & pi0090;
assign w2616 = ~pi0841 & w2615;
assign w2617 = pi0058 & ~pi0090;
assign w2618 = ~w2616 & ~w2617;
assign w2619 = ~pi0095 & w107;
assign w2620 = ~w2618 & w2619;
assign w2621 = ~pi0032 & w2620;
assign w2622 = w374 & w2621;
assign w2623 = w386 & w2622;
assign w2624 = ~w2614 & w2623;
assign w2625 = pi0180 & ~pi0299;
assign w2626 = pi0158 & pi0299;
assign w2627 = ~w2625 & ~w2626;
assign w2628 = w7 & ~w2627;
assign w2629 = w196 & w2628;
assign w2630 = w194 & w2629;
assign w2631 = ~pi0040 & w2630;
assign w2632 = (~pi0040 & w2624) | (~pi0040 & w2631) | (w2624 & w2631);
assign w2633 = pi0032 & ~pi0039;
assign w2634 = (~pi0039 & ~w2632) | (~pi0039 & w2633) | (~w2632 & w2633);
assign w2635 = ~w2611 & w2634;
assign w2636 = ~w2607 & w2635;
assign w2637 = w1240 & w1245;
assign w2638 = ~pi0152 & w1257;
assign w2639 = ~w2637 & w2638;
assign w2640 = ~pi0174 & w1259;
assign w2641 = ~w1274 & w2640;
assign w2642 = ~w2639 & ~w2641;
assign w2643 = w1478 & ~w2642;
assign w2644 = pi0154 & w1257;
assign w2645 = ~w2637 & w2644;
assign w2646 = pi0176 & w1259;
assign w2647 = ~w1274 & w2646;
assign w2648 = ~w2645 & ~w2647;
assign w2649 = w1237 & ~w2648;
assign w2650 = ~w2643 & ~w2649;
assign w2651 = w113 & ~w2650;
assign w2652 = ~pi0038 & w171;
assign w2653 = w2483 & w2652;
assign w2654 = ~pi0039 & w171;
assign w2655 = ~pi0038 & w2654;
assign w2656 = w2483 & w2655;
assign w2657 = (w2651 & w2653) | (w2651 & w2656) | (w2653 & w2656);
assign w2658 = ~w2636 & w2657;
assign w2659 = w254 & w377;
assign w2660 = ~pi0164 & pi0299;
assign w2661 = ~pi0186 & ~pi0299;
assign w2662 = ~w2660 & ~w2661;
assign w2663 = w2483 & w2662;
assign w2664 = ~pi0074 & w2;
assign w2665 = (~pi0074 & w2663) | (~pi0074 & w2664) | (w2663 & w2664);
assign w2666 = pi0033 & pi0954;
assign w2667 = ~pi0033 & ~pi0954;
assign w2668 = ~w2666 & ~w2667;
assign w2669 = ~pi0138 & ~pi0139;
assign w2670 = ~pi0195 & ~pi0196;
assign w2671 = w2669 & w2670;
assign w2672 = ~pi0079 & ~pi0118;
assign w2673 = ~pi0033 & w2672;
assign w2674 = w2671 & w2673;
assign w2675 = pi0034 & ~w2668;
assign w2676 = (~w2668 & ~w2674) | (~w2668 & w2675) | (~w2674 & w2675);
assign w2677 = w2665 & ~w2676;
assign w2678 = ~pi0040 & w532;
assign w2679 = w1300 & w2678;
assign w2680 = w2677 & w2679;
assign w2681 = w2594 & w2680;
assign w2682 = w104 & ~w2594;
assign w2683 = ~w393 & w2682;
assign w2684 = w492 & w2683;
assign w2685 = w2680 & ~w2684;
assign w2686 = (~w2659 & w2681) | (~w2659 & w2685) | (w2681 & w2685);
assign w2687 = ~w357 & ~w359;
assign w2688 = (~w357 & ~w374) | (~w357 & w2687) | (~w374 & w2687);
assign w2689 = (~w112 & ~w357) | (~w112 & w2688) | (~w357 & w2688);
assign w2690 = ~w1389 & ~w2621;
assign w2691 = w1395 & ~w2689;
assign w2692 = (~w2689 & ~w2690) | (~w2689 & w2691) | (~w2690 & w2691);
assign w2693 = w99 & w1342;
assign w2694 = pi0073 & w2693;
assign w2695 = w1352 & w2694;
assign w2696 = ~w2692 & ~w2695;
assign w2697 = w2686 & w2696;
assign w2698 = ~w1237 & ~w1478;
assign w2699 = ~w1270 & ~w2698;
assign w2700 = w1342 & w1351;
assign w2701 = w1348 & w2700;
assign w2702 = w1354 & w1658;
assign w2703 = w2701 & w2702;
assign w2704 = w2699 & w2703;
assign w2705 = w2 & w2678;
assign w2706 = (w2663 & w2678) | (w2663 & w2705) | (w2678 & w2705);
assign w2707 = ~pi0074 & w147;
assign w2708 = w2706 & w2707;
assign w2709 = ~w2704 & w2708;
assign w2710 = ~pi0034 & w2672;
assign w2711 = w2671 & w2710;
assign w2712 = ~pi0033 & pi0954;
assign w2713 = pi0033 & ~pi0954;
assign w2714 = ~w2712 & ~w2713;
assign w2715 = ~w0 & ~w2714;
assign w2716 = pi0954 & ~w2712;
assign w2717 = ~w0 & ~w2716;
assign w2718 = (w2711 & w2715) | (w2711 & w2717) | (w2715 & w2717);
assign w2719 = w1342 & w1354;
assign w2720 = w1352 & w2719;
assign w2721 = pi0092 & ~w2714;
assign w2722 = pi0092 & ~w2716;
assign w2723 = (w2711 & w2721) | (w2711 & w2722) | (w2721 & w2722);
assign w2724 = ~w2720 & ~w2723;
assign w2725 = pi0154 & pi0299;
assign w2726 = pi0176 & ~pi0299;
assign w2727 = ~w2725 & ~w2726;
assign w2728 = w2483 & ~w2727;
assign w2729 = pi0092 & w0;
assign w2730 = w2728 & w2729;
assign w2731 = w1351 & ~w2730;
assign w2732 = w1348 & w2731;
assign w2733 = w2719 & w2732;
assign w2734 = ~w2718 & w2733;
assign w2735 = (~w2718 & w2724) | (~w2718 & w2734) | (w2724 & w2734);
assign w2736 = w2709 & ~w2735;
assign w2737 = ~w2697 & ~w2736;
assign w2738 = w83 & w2532;
assign w2739 = w74 & w2738;
assign w2740 = w1658 & w2525;
assign w2741 = w1641 & w2740;
assign w2742 = ~pi0054 & w2741;
assign w2743 = w99 & w2742;
assign w2744 = ~w2 & ~w2743;
assign w2745 = (~w2 & ~w2739) | (~w2 & w2744) | (~w2739 & w2744);
assign w2746 = ~pi0149 & pi0157;
assign w2747 = pi0149 & ~pi0157;
assign w2748 = ~w2746 & ~w2747;
assign w2749 = pi0299 & ~w2748;
assign w2750 = pi0178 & ~pi0183;
assign w2751 = ~pi0178 & pi0183;
assign w2752 = ~w2750 & ~w2751;
assign w2753 = ~pi0299 & ~w2752;
assign w2754 = ~w2749 & ~w2753;
assign w2755 = ~w147 & w2483;
assign w2756 = ~w2754 & w2755;
assign w2757 = pi0191 & ~pi0299;
assign w2758 = pi0169 & pi0299;
assign w2759 = ~w2757 & ~w2758;
assign w2760 = w2483 & ~w2759;
assign w2761 = pi0074 & w2760;
assign w2762 = w147 & ~w2761;
assign w2763 = ~w2756 & ~w2762;
assign w2764 = w147 & ~w2665;
assign w2765 = ~w2761 & w2764;
assign w2766 = ~w2756 & ~w2765;
assign w2767 = (w2745 & w2763) | (w2745 & w2766) | (w2763 & w2766);
assign w2768 = w529 & ~w2767;
assign w2769 = w2737 & w2768;
assign w2770 = ~w2658 & w2769;
assign w2771 = pi0074 & pi0169;
assign w2772 = w2 & w179;
assign w2773 = ~pi0074 & pi0164;
assign w2774 = ~w2771 & ~w2773;
assign w2775 = (~w2771 & w2772) | (~w2771 & w2774) | (w2772 & w2774);
assign w2776 = w147 & ~w2483;
assign w2777 = (w147 & w2775) | (w147 & w2776) | (w2775 & w2776);
assign w2778 = ~w147 & ~w2748;
assign w2779 = w2483 & w2778;
assign w2780 = ~w2777 & ~w2779;
assign w2781 = ~w529 & ~w2780;
assign w2782 = pi0149 & w546;
assign w2783 = w2483 & w2782;
assign w2784 = w567 & w2783;
assign w2785 = ~w546 & ~w2676;
assign w2786 = (~w567 & ~w2676) | (~w567 & w2785) | (~w2676 & w2785);
assign w2787 = ~w2784 & ~w2786;
assign w2788 = ~pi0040 & w179;
assign w2789 = w534 & w2788;
assign w2790 = w2781 & ~w2789;
assign w2791 = (w2781 & w2787) | (w2781 & w2790) | (w2787 & w2790);
assign w2792 = ~w2770 & ~w2791;
assign w2793 = pi0162 & pi0299;
assign w2794 = ~w2595 & w2793;
assign w2795 = pi0140 & ~pi0299;
assign w2796 = ~w2602 & w2795;
assign w2797 = ~w2794 & ~w2796;
assign w2798 = ~pi0159 & pi0299;
assign w2799 = ~pi0181 & ~pi0299;
assign w2800 = ~w2798 & ~w2799;
assign w2801 = w7 & w2800;
assign w2802 = ~pi0161 & pi0299;
assign w2803 = ~pi0144 & ~pi0299;
assign w2804 = ~w2802 & ~w2803;
assign w2805 = pi0073 & ~w2804;
assign w2806 = ~w2801 & ~w2805;
assign w2807 = w2797 & w2806;
assign w2808 = ~pi0146 & pi0299;
assign w2809 = ~pi0142 & ~pi0299;
assign w2810 = ~w2808 & ~w2809;
assign w2811 = w2807 & w2810;
assign w2812 = (~w2623 & w2807) | (~w2623 & w2811) | (w2807 & w2811);
assign w2813 = w2483 & ~w2812;
assign w2814 = w594 & w2813;
assign w2815 = ~w2553 & w2814;
assign w2816 = ~pi0073 & w1;
assign w2817 = w99 & w2816;
assign w2818 = w546 & w2817;
assign w2819 = w2701 & w2818;
assign w2820 = pi0055 & pi0162;
assign w2821 = w2789 & w2820;
assign w2822 = w2819 & w2821;
assign w2823 = w1354 & w2701;
assign w2824 = ~pi0055 & w546;
assign w2825 = ~w1 & w2824;
assign w2826 = (~w5 & w2824) | (~w5 & w2825) | (w2824 & w2825);
assign w2827 = w2789 & w2826;
assign w2828 = w2823 & w2827;
assign w2829 = w2699 & w2828;
assign w2830 = ~pi0161 & ~w1472;
assign w2831 = (~w1257 & ~w1472) | (~w1257 & w2830) | (~w1472 & w2830);
assign w2832 = pi0144 & ~w1257;
assign w2833 = w2831 & ~w2832;
assign w2834 = ~pi0155 & w1257;
assign w2835 = ~w2637 & w2834;
assign w2836 = ~pi0177 & ~w1257;
assign w2837 = (~pi0177 & w2637) | (~pi0177 & w2836) | (w2637 & w2836);
assign w2838 = ~w2835 & ~w2837;
assign w2839 = ~w1236 & ~w2833;
assign w2840 = (~w2833 & ~w2838) | (~w2833 & w2839) | (~w2838 & w2839);
assign w2841 = w1658 & ~w2840;
assign w2842 = ~w2822 & ~w2841;
assign w2843 = (~w2822 & ~w2829) | (~w2822 & w2842) | (~w2829 & w2842);
assign w2844 = ~pi0162 & ~pi0197;
assign w2845 = pi0162 & pi0197;
assign w2846 = ~w2844 & ~w2845;
assign w2847 = ~pi0149 & ~pi0157;
assign w2848 = ~w2846 & w2847;
assign w2849 = pi0162 & ~pi0197;
assign w2850 = ~pi0162 & pi0197;
assign w2851 = ~w2849 & ~w2850;
assign w2852 = ~w2847 & ~w2851;
assign w2853 = ~w2848 & ~w2852;
assign w2854 = ~w147 & w2853;
assign w2855 = pi0074 & pi0148;
assign w2856 = ~pi0074 & pi0167;
assign w2857 = ~w2855 & ~w2856;
assign w2858 = (w2772 & ~w2855) | (w2772 & w2857) | (~w2855 & w2857);
assign w2859 = w147 & ~w2858;
assign w2860 = ~w529 & ~w2859;
assign w2861 = ~w2854 & w2860;
assign w2862 = pi0188 & ~pi0299;
assign w2863 = pi0167 & pi0299;
assign w2864 = ~w2862 & ~w2863;
assign w2865 = w2707 & ~w2864;
assign w2866 = w2745 & w2865;
assign w2867 = pi0140 & pi0145;
assign w2868 = ~pi0140 & ~pi0145;
assign w2869 = ~w2867 & ~w2868;
assign w2870 = ~pi0178 & ~pi0183;
assign w2871 = ~w2869 & w2870;
assign w2872 = pi0140 & ~pi0145;
assign w2873 = ~pi0140 & pi0145;
assign w2874 = ~w2872 & ~w2873;
assign w2875 = ~w2870 & ~w2874;
assign w2876 = ~w2871 & ~w2875;
assign w2877 = ~pi0299 & ~w2876;
assign w2878 = pi0299 & ~w2853;
assign w2879 = ~w2877 & ~w2878;
assign w2880 = pi0148 & pi0299;
assign w2881 = pi0141 & ~pi0299;
assign w2882 = ~w2880 & ~w2881;
assign w2883 = pi0074 & w147;
assign w2884 = ~w2882 & w2883;
assign w2885 = w529 & ~w2884;
assign w2886 = w147 & ~w2884;
assign w2887 = w529 & w2886;
assign w2888 = (~w2879 & w2885) | (~w2879 & w2887) | (w2885 & w2887);
assign w2889 = ~w2861 & ~w2888;
assign w2890 = (~w2861 & w2866) | (~w2861 & w2889) | (w2866 & w2889);
assign w2891 = w2483 & w2890;
assign w2892 = (w2483 & ~w2843) | (w2483 & w2891) | (~w2843 & w2891);
assign w2893 = ~w2815 & ~w2892;
assign w2894 = w593 & w2594;
assign w2895 = w593 & ~w2684;
assign w2896 = (~w2659 & w2894) | (~w2659 & w2895) | (w2894 & w2895);
assign w2897 = w2696 & w2896;
assign w2898 = pi0034 & ~w2667;
assign w2899 = ~pi0034 & ~pi0954;
assign w2900 = ~pi0033 & pi0034;
assign w2901 = w2899 & w2900;
assign w2902 = ~w2898 & ~w2901;
assign w2903 = ~pi0033 & w2899;
assign w2904 = ~w2898 & ~w2903;
assign w2905 = (w2674 & w2902) | (w2674 & w2904) | (w2902 & w2904);
assign w2906 = w2789 & w2905;
assign w2907 = pi0055 & ~w2817;
assign w2908 = (pi0055 & ~w2701) | (pi0055 & w2907) | (~w2701 & w2907);
assign w2909 = w546 & ~w2908;
assign w2910 = w2789 & ~w2909;
assign w2911 = w2905 & w2910;
assign w2912 = (w2897 & w2906) | (w2897 & w2911) | (w2906 & w2911);
assign w2913 = w2893 & ~w2912;
assign w2914 = ~pi0032 & w0;
assign w2915 = ~pi0095 & w2914;
assign w2916 = w188 & w2915;
assign w2917 = w1354 & w2916;
assign w2918 = w1352 & w2917;
assign w2919 = pi0177 & ~pi0299;
assign w2920 = pi0155 & pi0299;
assign w2921 = ~w2919 & ~w2920;
assign w2922 = w2483 & ~w2921;
assign w2923 = w2918 & w2922;
assign w2924 = w2905 & ~w2918;
assign w2925 = ~w2923 & ~w2924;
assign w2926 = ~w2704 & ~w2925;
assign w2927 = w2827 & w2926;
assign w2928 = w2913 & ~w2927;
assign w2929 = ~pi0024 & ~pi0054;
assign w2930 = pi0059 & ~w2929;
assign w2931 = ~pi0057 & w546;
assign w2932 = ~pi0074 & w2931;
assign w2933 = ~w2930 & w2932;
assign w2934 = ~pi0055 & w2933;
assign w2935 = ~pi0074 & ~w2772;
assign w2936 = w348 & w1358;
assign w2937 = w1 & w2936;
assign w2938 = w2935 & ~w2937;
assign w2939 = w2934 & ~w2938;
assign w2940 = w1300 & w2939;
assign w2941 = ~pi0054 & ~w1395;
assign w2942 = ~pi0024 & ~w2941;
assign w2943 = ~pi0059 & ~w2942;
assign w2944 = ~w2940 & w2943;
assign w2945 = w2934 & w2944;
assign w2946 = w2 & w134;
assign w2947 = pi1091 & w449;
assign w2948 = pi1093 & w2947;
assign w2949 = pi0824 & ~w2948;
assign w2950 = w1280 & w2949;
assign w2951 = pi0683 & w2950;
assign w2952 = w2485 & ~w2951;
assign w2953 = ~pi0137 & ~w2485;
assign w2954 = ~w2952 & ~w2953;
assign w2955 = pi0252 & ~w2954;
assign w2956 = ~w1323 & ~w2573;
assign w2957 = pi0137 & ~w2956;
assign w2958 = w1318 & w2471;
assign w2959 = ~pi0052 & w2958;
assign w2960 = w2957 & w2959;
assign w2961 = pi0129 & w2571;
assign w2962 = ~w2960 & ~w2961;
assign w2963 = ~w2955 & ~w2962;
assign w2964 = w2946 & w2963;
assign w2965 = ~pi0038 & pi0075;
assign w2966 = pi0137 & ~w1320;
assign w2967 = ~w454 & w2966;
assign w2968 = ~w2580 & ~w2967;
assign w2969 = w2965 & ~w2968;
assign w2970 = pi0038 & ~pi0075;
assign w2971 = ~w2969 & ~w2970;
assign w2972 = w2487 & ~w2971;
assign w2973 = ~w2964 & ~w2972;
assign w2974 = w2937 & ~w2973;
assign w2975 = w2945 & w2974;
assign w2976 = w378 & w407;
assign w2977 = ~w205 & ~w407;
assign w2978 = ~w2976 & ~w2977;
assign w2979 = ~pi0035 & pi0841;
assign w2980 = ~pi0093 & ~pi0841;
assign w2981 = ~w2979 & ~w2980;
assign w2982 = ~w1236 & ~w2043;
assign w2983 = ~pi0122 & ~w2568;
assign w2984 = ~w2982 & w2983;
assign w2985 = ~pi0137 & w413;
assign w2986 = pi0076 & ~w2985;
assign w2987 = w2984 & w2986;
assign w2988 = ~pi0058 & ~w2987;
assign w2989 = ~w2981 & w2988;
assign w2990 = pi0040 & pi1082;
assign w2991 = w2989 & ~w2990;
assign w2992 = pi0035 & ~pi0841;
assign w2993 = ~w2991 & ~w2992;
assign w2994 = ~w2978 & w2993;
assign w2995 = w2943 & ~w2994;
assign w2996 = w2940 & ~w2995;
assign w2997 = ~w2975 & ~w2996;
assign w2998 = w465 & w2466;
assign w2999 = pi0036 & w99;
assign w3000 = w193 & w484;
assign w3001 = w2999 & w3000;
assign w3002 = ~w2998 & ~w3001;
assign w3003 = w104 & w529;
assign w3004 = w6 & w3003;
assign w3005 = w107 & w3004;
assign w3006 = ~w3002 & w3005;
assign w3007 = w2568 & w3006;
assign w3008 = w1440 & w1609;
assign w3009 = ~w1650 & ~w3008;
assign w3010 = ~w1623 & w3009;
assign w3011 = w1620 & w3010;
assign w3012 = w99 & w3005;
assign w3013 = w484 & w3012;
assign w3014 = w193 & w3013;
assign w3015 = pi0089 & pi0332;
assign w3016 = w3014 & w3015;
assign w3017 = w196 & w3012;
assign w3018 = ~w234 & w3017;
assign w3019 = pi0064 & w3018;
assign w3020 = ~w3016 & ~w3019;
assign w3021 = ~pi0841 & ~w3020;
assign w3022 = pi0024 & w1615;
assign w3023 = ~w3021 & ~w3022;
assign w3024 = pi0835 & pi0984;
assign w3025 = ~w1229 & ~w3024;
assign w3026 = ~pi0979 & w3025;
assign w3027 = ~pi1093 & ~w1293;
assign w3028 = pi0299 & w1240;
assign w3029 = w1286 & w3028;
assign w3030 = w1278 & ~w3029;
assign w3031 = w1284 & w3030;
assign w3032 = ~w3027 & w3031;
assign w3033 = pi0835 & w3032;
assign w3034 = pi0835 & w3031;
assign w3035 = ~pi1082 & ~w3034;
assign w3036 = pi0786 & w3035;
assign w3037 = ~w3033 & ~w3036;
assign w3038 = w3026 & w3037;
assign w3039 = ~pi0287 & w1648;
assign w3040 = w1636 & w3039;
assign w3041 = w3038 & w3040;
assign w3042 = w349 & w380;
assign w3043 = w359 & w3042;
assign w3044 = w99 & w348;
assign w3045 = w355 & w388;
assign w3046 = (w355 & w392) | (w355 & w3045) | (w392 & w3045);
assign w3047 = w107 & ~w401;
assign w3048 = ~pi0090 & w3047;
assign w3049 = (~pi0090 & w3046) | (~pi0090 & w3048) | (w3046 & w3048);
assign w3050 = w3044 & w3049;
assign w3051 = ~w3043 & ~w3050;
assign w3052 = w112 & ~w3051;
assign w3053 = ~w254 & ~w313;
assign w3054 = (~w254 & ~w484) | (~w254 & w3053) | (~w484 & w3053);
assign w3055 = ~w377 & ~w3052;
assign w3056 = (~w3052 & w3054) | (~w3052 & w3055) | (w3054 & w3055);
assign w3057 = ~pi0035 & ~pi0048;
assign w3058 = pi0841 & ~w3057;
assign w3059 = ~pi0986 & ~w2568;
assign w3060 = pi0252 & ~w3059;
assign w3061 = pi0314 & ~w3060;
assign w3062 = pi0108 & w3061;
assign w3063 = ~pi0048 & ~w3062;
assign w3064 = ~pi0035 & w3063;
assign w3065 = ~pi0047 & w3064;
assign w3066 = ~w3058 & ~w3065;
assign w3067 = ~w3056 & w3066;
assign w3068 = pi0032 & ~w413;
assign w3069 = ~pi0040 & w3068;
assign w3070 = ~pi0095 & w3069;
assign w3071 = ~pi0841 & w3070;
assign w3072 = w1358 & w3071;
assign w3073 = ~w3067 & ~w3072;
assign w3074 = w593 & ~w3073;
assign w3075 = ~w3041 & ~w3074;
assign w3076 = pi0040 & ~pi1082;
assign w3077 = ~pi0040 & pi0102;
assign w3078 = ~w3076 & ~w3077;
assign w3079 = w2554 & ~w3078;
assign w3080 = w180 & w1644;
assign w3081 = w1643 & w3080;
assign w3082 = w1633 & w3081;
assign w3083 = ~pi0189 & w525;
assign w3084 = w180 & w3083;
assign w3085 = pi0144 & ~pi0174;
assign w3086 = w3084 & w3085;
assign w3087 = ~pi0152 & pi0161;
assign w3088 = ~pi0166 & w3087;
assign w3089 = ~w526 & w3088;
assign w3090 = ~w3086 & ~w3089;
assign w3091 = pi0287 & w1634;
assign w3092 = w1345 & w3091;
assign w3093 = w2483 & ~w3092;
assign w3094 = ~w3090 & w3093;
assign w3095 = pi0039 & ~w3094;
assign w3096 = w2483 & ~w3090;
assign w3097 = pi0039 & ~w3096;
assign w3098 = (w3082 & w3095) | (w3082 & w3097) | (w3095 & w3097);
assign w3099 = ~w2433 & w2445;
assign w3100 = w429 & w2461;
assign w3101 = w2457 & w3100;
assign w3102 = w2451 & w3101;
assign w3103 = w465 & w3102;
assign w3104 = pi0096 & ~w454;
assign w3105 = ~w3103 & w3104;
assign w3106 = (w3099 & ~w3103) | (w3099 & w3105) | (~w3103 & w3105);
assign w3107 = pi0228 & w169;
assign w3108 = pi0100 & ~pi0122;
assign w3109 = w3107 & ~w3108;
assign w3110 = (~w1236 & w3107) | (~w1236 & w3109) | (w3107 & w3109);
assign w3111 = (~w2485 & w3107) | (~w2485 & w3110) | (w3107 & w3110);
assign w3112 = w429 & w453;
assign w3113 = w382 & w1235;
assign w3114 = w3112 & w3113;
assign w3115 = pi0097 & ~pi0122;
assign w3116 = w3114 & w3115;
assign w3117 = w3111 & ~w3116;
assign w3118 = (~w251 & w3111) | (~w251 & w3117) | (w3111 & w3117);
assign w3119 = ~w2539 & ~w3118;
assign w3120 = (~w2539 & ~w3106) | (~w2539 & w3119) | (~w3106 & w3119);
assign w3121 = ~pi0094 & pi0110;
assign w3122 = ~pi0480 & pi0949;
assign w3123 = w3121 & w3122;
assign w3124 = pi0094 & ~pi0110;
assign w3125 = ~pi0250 & pi0252;
assign w3126 = pi0901 & ~pi0959;
assign w3127 = w3125 & w3126;
assign w3128 = w3124 & w3127;
assign w3129 = ~w3123 & ~w3128;
assign w3130 = w254 & ~w3129;
assign w3131 = w112 & w374;
assign w3132 = ~pi0070 & ~w350;
assign w3133 = ~pi0051 & w3132;
assign w3134 = w357 & w3133;
assign w3135 = ~pi0228 & ~w3134;
assign w3136 = w106 & w360;
assign w3137 = ~pi0228 & ~w3136;
assign w3138 = (~w3131 & w3135) | (~w3131 & w3137) | (w3135 & w3137);
assign w3139 = (~pi0228 & ~w3130) | (~pi0228 & w3138) | (~w3130 & w3138);
assign w3140 = w3120 & ~w3139;
assign w3141 = w147 & w169;
assign w3142 = w169 & w3141;
assign w3143 = (w169 & w2490) | (w169 & w3141) | (w2490 & w3141);
assign w3144 = (w2485 & w3142) | (w2485 & w3143) | (w3142 & w3143);
assign w3145 = ~w147 & ~w169;
assign w3146 = ~w2490 & w3145;
assign w3147 = (~w2485 & w3145) | (~w2485 & w3146) | (w3145 & w3146);
assign w3148 = ~w3144 & w3147;
assign w3149 = (~w113 & ~w3144) | (~w113 & w3148) | (~w3144 & w3148);
assign w3150 = ~pi0038 & ~pi0092;
assign w3151 = w168 & w3150;
assign w3152 = w529 & w3151;
assign w3153 = ~w3149 & w3152;
assign w3154 = ~pi0044 & ~pi0101;
assign w3155 = w3153 & w3154;
assign w3156 = ~pi0041 & ~w3155;
assign w3157 = (~pi0041 & ~w3140) | (~pi0041 & w3156) | (~w3140 & w3156);
assign w3158 = pi0041 & w3154;
assign w3159 = w3153 & w3158;
assign w3160 = w3140 & w3159;
assign w3161 = ~w3157 & ~w3160;
assign w3162 = pi0039 & ~w3098;
assign w3163 = (~w3098 & w3161) | (~w3098 & w3162) | (w3161 & w3162);
assign w3164 = ~pi0072 & ~w3163;
assign w3165 = ~w3139 & w3153;
assign w3166 = w3120 & w3165;
assign w3167 = ~pi0042 & ~pi0116;
assign w3168 = w1311 & w3167;
assign w3169 = w1318 & w3168;
assign w3170 = w3166 & w3169;
assign w3171 = ~pi0116 & w1311;
assign w3172 = w1318 & w3171;
assign w3173 = pi0042 & ~w3172;
assign w3174 = (pi0042 & ~w3166) | (pi0042 & w3173) | (~w3166 & w3173);
assign w3175 = ~w3170 & ~w3174;
assign w3176 = w2525 & ~w3175;
assign w3177 = pi0207 & pi0208;
assign w3178 = ~pi0199 & ~pi0200;
assign w3179 = (~pi0199 & ~w3177) | (~pi0199 & w3178) | (~w3177 & w3178);
assign w3180 = w526 & w3179;
assign w3181 = pi0211 & pi0214;
assign w3182 = ~pi0212 & ~pi0219;
assign w3183 = (~pi0219 & ~w3181) | (~pi0219 & w3182) | (~w3181 & w3182);
assign w3184 = ~w526 & w3183;
assign w3185 = ~w3180 & ~w3184;
assign w3186 = pi0166 & ~w525;
assign w3187 = (pi0166 & ~w180) | (pi0166 & w3186) | (~w180 & w3186);
assign w3188 = pi0189 & w525;
assign w3189 = w180 & w3188;
assign w3190 = ~w3187 & ~w3189;
assign w3191 = w1645 & ~w2483;
assign w3192 = (w1645 & ~w3190) | (w1645 & w3191) | (~w3190 & w3191);
assign w3193 = w3185 & w3192;
assign w3194 = w3093 & w3190;
assign w3195 = w1645 & ~w3194;
assign w3196 = w3185 & w3195;
assign w3197 = (w3082 & w3193) | (w3082 & w3196) | (w3193 & w3196);
assign w3198 = ~w3176 & ~w3197;
assign w3199 = w3166 & w3172;
assign w3200 = w1310 & w3199;
assign w3201 = pi0043 & ~w3170;
assign w3202 = ~w3200 & ~w3201;
assign w3203 = w2525 & ~w3202;
assign w3204 = (w3082 & w3192) | (w3082 & w3195) | (w3192 & w3195);
assign w3205 = ~pi0200 & w3177;
assign w3206 = ~pi0199 & w3205;
assign w3207 = pi0200 & ~w3177;
assign w3208 = ~w3206 & ~w3207;
assign w3209 = w526 & ~w3208;
assign w3210 = ~pi0211 & pi0214;
assign w3211 = pi0212 & ~pi0219;
assign w3212 = w3210 & w3211;
assign w3213 = pi0212 & pi0214;
assign w3214 = pi0211 & ~w3213;
assign w3215 = ~w3212 & ~w3214;
assign w3216 = ~w526 & ~w3215;
assign w3217 = ~w3209 & ~w3216;
assign w3218 = w3204 & ~w3217;
assign w3219 = ~w3203 & ~w3218;
assign w3220 = ~pi0044 & w3166;
assign w3221 = pi0044 & ~w3166;
assign w3222 = ~w3220 & ~w3221;
assign w3223 = ~pi0039 & ~w3222;
assign w3224 = (w2483 & ~w3082) | (w2483 & w3093) | (~w3082 & w3093);
assign w3225 = ~pi0189 & w2478;
assign w3226 = w526 & w3225;
assign w3227 = ~pi0166 & w2475;
assign w3228 = ~w526 & w3227;
assign w3229 = ~w3226 & ~w3228;
assign w3230 = pi0039 & ~w3229;
assign w3231 = w3224 & w3230;
assign w3232 = ~w3223 & ~w3231;
assign w3233 = ~pi0072 & ~w3232;
assign w3234 = pi0979 & w3040;
assign w3235 = pi0061 & ~pi0841;
assign w3236 = w3014 & w3235;
assign w3237 = w477 & ~w2689;
assign w3238 = w349 & w3237;
assign w3239 = w593 & w3238;
assign w3240 = pi0046 & w3239;
assign w3241 = pi0024 & w3240;
assign w3242 = ~w3236 & ~w3241;
assign w3243 = pi0104 & w3014;
assign w3244 = pi0088 & w3018;
assign w3245 = ~w3243 & ~w3244;
assign w3246 = ~w2950 & ~w3245;
assign w3247 = pi0824 & ~pi1093;
assign w3248 = w1280 & w3247;
assign w3249 = ~w454 & ~w3248;
assign w3250 = w3006 & w3249;
assign w3251 = ~w3246 & ~w3250;
assign w3252 = pi0048 & w3014;
assign w3253 = pi0841 & w3252;
assign w3254 = pi0049 & pi0841;
assign w3255 = w3014 & w3254;
assign w3256 = ~pi0092 & w2929;
assign w3257 = ~pi0100 & w3256;
assign w3258 = w118 & w3257;
assign w3259 = pi0074 & w3258;
assign w3260 = ~pi0075 & w3259;
assign w3261 = w1297 & w3260;
assign w3262 = ~w3255 & ~w3261;
assign w3263 = pi0050 & w443;
assign w3264 = ~pi0077 & w97;
assign w3265 = ~pi0109 & w89;
assign w3266 = w112 & w3005;
assign w3267 = w3265 & w3266;
assign w3268 = w3264 & w3267;
assign w3269 = pi0024 & w3268;
assign w3270 = ~pi0110 & w3269;
assign w3271 = w3263 & w3270;
assign w3272 = w95 & w3267;
assign w3273 = w94 & w3272;
assign w3274 = ~pi0086 & w3273;
assign w3275 = pi0094 & w3274;
assign w3276 = ~pi0110 & w3275;
assign w3277 = ~pi0252 & w2485;
assign w3278 = pi0252 & w454;
assign w3279 = ~w3277 & ~w3278;
assign w3280 = w3276 & ~w3279;
assign w3281 = ~w3271 & ~w3280;
assign w3282 = pi0075 & w2487;
assign w3283 = ~w454 & w3282;
assign w3284 = ~w1444 & ~w3283;
assign w3285 = w1320 & ~w3284;
assign w3286 = w1622 & w3285;
assign w3287 = w3281 & ~w3286;
assign w3288 = w193 & w3012;
assign w3289 = w65 & w279;
assign w3290 = ~pi0067 & w3289;
assign w3291 = ~pi0071 & w3290;
assign w3292 = w3288 & w3291;
assign w3293 = w334 & w3292;
assign w3294 = pi0082 & w3293;
assign w3295 = ~pi0111 & w3294;
assign w3296 = w1319 & w3166;
assign w3297 = pi0052 & ~w2958;
assign w3298 = (pi0052 & ~w3166) | (pi0052 & w3297) | (~w3166 & w3297);
assign w3299 = ~w3296 & ~w3298;
assign w3300 = w2525 & ~w3299;
assign w3301 = ~w3177 & w3178;
assign w3302 = pi0199 & pi0200;
assign w3303 = ~w3301 & ~w3302;
assign w3304 = w526 & ~w3303;
assign w3305 = ~pi0211 & ~pi0219;
assign w3306 = ~w3213 & w3305;
assign w3307 = pi0211 & pi0219;
assign w3308 = ~w3306 & ~w3307;
assign w3309 = ~w526 & ~w3308;
assign w3310 = ~w3304 & ~w3309;
assign w3311 = ~w3185 & ~w3310;
assign w3312 = w3192 & w3311;
assign w3313 = w3195 & w3311;
assign w3314 = (w3082 & w3312) | (w3082 & w3313) | (w3312 & w3313);
assign w3315 = ~w3300 & ~w3314;
assign w3316 = ~pi0050 & w3268;
assign w3317 = pi0053 & w3316;
assign w3318 = ~pi0060 & w3317;
assign w3319 = ~pi0110 & w3318;
assign w3320 = pi0024 & w3319;
assign w3321 = ~pi0979 & w3024;
assign w3322 = w3040 & w3321;
assign w3323 = ~w3320 & ~w3322;
assign w3324 = pi0024 & ~pi0074;
assign w3325 = w1300 & w1619;
assign w3326 = w3324 & w3325;
assign w3327 = w193 & w3005;
assign w3328 = w99 & w3327;
assign w3329 = w342 & w3328;
assign w3330 = ~pi0071 & w3329;
assign w3331 = w484 & w3330;
assign w3332 = pi0106 & w3331;
assign w3333 = ~pi0841 & w3332;
assign w3334 = ~w3326 & ~w3333;
assign w3335 = w2819 & ~w3014;
assign w3336 = pi0024 & w2789;
assign w3337 = w3335 & w3336;
assign w3338 = pi0045 & w3014;
assign w3339 = ~w3337 & ~w3338;
assign w3340 = ~pi0055 & pi0056;
assign w3341 = pi0841 & w3340;
assign w3342 = pi0055 & ~pi0056;
assign w3343 = ~pi0024 & w3342;
assign w3344 = ~w3341 & ~w3343;
assign w3345 = w2789 & ~w3344;
assign w3346 = ~pi0062 & w3345;
assign w3347 = w2823 & w3346;
assign w3348 = w1 & w3347;
assign w3349 = ~pi0056 & pi0924;
assign w3350 = w1355 & ~w3349;
assign w3351 = ~pi0841 & w3350;
assign w3352 = pi0024 & w1338;
assign w3353 = ~pi0055 & w3352;
assign w3354 = pi0057 & w3353;
assign w3355 = ~pi0059 & w3354;
assign w3356 = ~w3351 & ~w3355;
assign w3357 = w349 & w492;
assign w3358 = w593 & w3357;
assign w3359 = w355 & w3358;
assign w3360 = pi0090 & w3359;
assign w3361 = ~pi0841 & w3360;
assign w3362 = ~pi0841 & pi0924;
assign w3363 = pi0062 & w1355;
assign w3364 = w3362 & w3363;
assign w3365 = w567 & w2824;
assign w3366 = pi0024 & w3365;
assign w3367 = ~pi0057 & w3366;
assign w3368 = pi0059 & w3367;
assign w3369 = ~w3364 & ~w3368;
assign w3370 = ~pi0053 & pi0060;
assign w3371 = ~pi0050 & w3270;
assign w3372 = w3370 & w3371;
assign w3373 = ~w3024 & w3040;
assign w3374 = ~pi0252 & w3373;
assign w3375 = ~pi0979 & w3374;
assign w3376 = ~pi1001 & w3375;
assign w3377 = ~w3372 & ~w3376;
assign w3378 = pi0061 & pi0841;
assign w3379 = w3014 & w3378;
assign w3380 = ~pi0024 & ~pi0050;
assign w3381 = ~pi0053 & w3380;
assign w3382 = pi0060 & w3381;
assign w3383 = w3268 & w3382;
assign w3384 = ~pi0110 & w3383;
assign w3385 = ~w3379 & ~w3384;
assign w3386 = ~pi0057 & pi0062;
assign w3387 = pi0841 & w3386;
assign w3388 = pi0057 & ~pi0062;
assign w3389 = ~pi0024 & w3388;
assign w3390 = ~w3387 & ~w3389;
assign w3391 = ~w1355 & ~w1619;
assign w3392 = w1616 & w3391;
assign w3393 = ~w1664 & w3392;
assign w3394 = ~w3390 & ~w3393;
assign w3395 = ~pi0024 & w3240;
assign w3396 = w1352 & w1354;
assign w3397 = w3005 & w3396;
assign w3398 = pi0063 & w3397;
assign w3399 = ~pi0107 & w3398;
assign w3400 = pi0999 & w3399;
assign w3401 = ~w3395 & ~w3400;
assign w3402 = pi0064 & pi0841;
assign w3403 = ~pi0107 & ~w3402;
assign w3404 = w3018 & ~w3403;
assign w3405 = w3035 & w3040;
assign w3406 = pi0786 & w3405;
assign w3407 = w3026 & w3406;
assign w3408 = pi0199 & ~pi0299;
assign w3409 = pi0219 & pi0299;
assign w3410 = ~w3408 & ~w3409;
assign w3411 = pi0081 & w78;
assign w3412 = ~pi0088 & w3411;
assign w3413 = ~pi0098 & w3412;
assign w3414 = pi0314 & w3413;
assign w3415 = w3017 & w3414;
assign w3416 = ~w3410 & w3415;
assign w3417 = ~pi0069 & w3292;
assign w3418 = ~pi0082 & w3417;
assign w3419 = ~pi0111 & w3418;
assign w3420 = pi0083 & w3419;
assign w3421 = ~pi0103 & w3420;
assign w3422 = pi0314 & w3421;
assign w3423 = pi0299 & w666;
assign w3424 = w1255 & w3423;
assign w3425 = w648 & w1268;
assign w3426 = ~w3424 & ~w3425;
assign w3427 = w1649 & ~w3426;
assign w3428 = w1478 & w3427;
assign w3429 = ~pi0314 & w320;
assign w3430 = ~pi0069 & pi0071;
assign w3431 = ~w3429 & ~w3430;
assign w3432 = w3014 & ~w3431;
assign w3433 = pi0024 & pi0070;
assign w3434 = w593 & w3052;
assign w3435 = w593 & ~w3055;
assign w3436 = (~w3054 & w3434) | (~w3054 & w3435) | (w3434 & w3435);
assign w3437 = w3433 & w3436;
assign w3438 = pi0210 & w1255;
assign w3439 = w12 & w3438;
assign w3440 = w16 & w1268;
assign w3441 = pi0198 & w3440;
assign w3442 = ~w3439 & ~w3441;
assign w3443 = pi0589 & ~w3442;
assign w3444 = ~pi0593 & w3443;
assign w3445 = ~w2698 & w3444;
assign w3446 = ~pi0287 & ~w3445;
assign w3447 = w1649 & ~w3446;
assign w3448 = ~w3437 & ~w3447;
assign w3449 = ~pi0076 & w61;
assign w3450 = pi0085 & w3449;
assign w3451 = ~pi0106 & w3450;
assign w3452 = w323 & w3451;
assign w3453 = pi0314 & w3452;
assign w3454 = w3330 & w3453;
assign w3455 = pi0200 & ~pi0299;
assign w3456 = ~pi0199 & w3455;
assign w3457 = ~pi0219 & pi0299;
assign w3458 = pi0211 & w3457;
assign w3459 = ~w3456 & ~w3458;
assign w3460 = w3415 & ~w3459;
assign w3461 = ~w3454 & ~w3460;
assign w3462 = pi0024 & w1641;
assign w3463 = pi0072 & w3462;
assign w3464 = w492 & w2532;
assign w3465 = w3463 & w3464;
assign w3466 = w1476 & ~w2947;
assign w3467 = pi0088 & w3466;
assign w3468 = w378 & w3467;
assign w3469 = ~w3465 & ~w3468;
assign w3470 = w593 & ~w3469;
assign w3471 = pi0299 & ~w32;
assign w3472 = ~pi0215 & w3471;
assign w3473 = w1255 & w3472;
assign w3474 = ~w2512 & ~w3473;
assign w3475 = w1649 & ~w3474;
assign w3476 = w1478 & w3475;
assign w3477 = ~w1470 & w3476;
assign w3478 = ~w3470 & ~w3477;
assign w3479 = ~pi0314 & pi1050;
assign w3480 = ~pi0039 & ~w3479;
assign w3481 = ~w1270 & w1478;
assign w3482 = w1649 & w3481;
assign w3483 = pi0073 & w529;
assign w3484 = w6 & w3483;
assign w3485 = ~w3482 & ~w3484;
assign w3486 = w378 & ~w3485;
assign w3487 = ~w3480 & w3486;
assign w3488 = pi0024 & pi0074;
assign w3489 = w1619 & w3488;
assign w3490 = pi0096 & ~pi0479;
assign w3491 = ~pi0841 & w3490;
assign w3492 = pi0479 & ~w413;
assign w3493 = ~pi0096 & ~w3492;
assign w3494 = ~w2568 & w3493;
assign w3495 = ~w3491 & ~w3494;
assign w3496 = ~w454 & ~w3495;
assign w3497 = ~pi0035 & w349;
assign w3498 = w254 & w382;
assign w3499 = pi0097 & w3498;
assign w3500 = w3497 & w3499;
assign w3501 = ~w433 & ~w3500;
assign w3502 = w593 & ~w3501;
assign w3503 = w3496 & w3502;
assign w3504 = ~w3489 & ~w3503;
assign w3505 = pi0024 & pi0075;
assign w3506 = w1619 & w3505;
assign w3507 = pi1093 & ~w432;
assign w3508 = ~w458 & ~w3507;
assign w3509 = w3502 & ~w3508;
assign w3510 = w454 & w3509;
assign w3511 = ~w3506 & ~w3510;
assign w3512 = ~pi0076 & pi0094;
assign w3513 = ~w2485 & w3512;
assign w3514 = ~pi0137 & w2043;
assign w3515 = w413 & w3514;
assign w3516 = ~w2984 & ~w3515;
assign w3517 = pi0076 & w3516;
assign w3518 = ~w3513 & ~w3517;
assign w3519 = ~pi0094 & w413;
assign w3520 = ~pi0137 & w3519;
assign w3521 = pi0094 & pi0252;
assign w3522 = ~w3520 & ~w3521;
assign w3523 = w454 & ~w3522;
assign w3524 = ~w3518 & ~w3523;
assign w3525 = w2554 & w3524;
assign w3526 = pi0077 & ~pi0314;
assign w3527 = ~pi0077 & pi0086;
assign w3528 = ~w3526 & ~w3527;
assign w3529 = w3436 & ~w3528;
assign w3530 = pi0119 & pi0232;
assign w3531 = ~pi0468 & w3530;
assign w3532 = (~w2594 & w2659) | (~w2594 & w2684) | (w2659 & w2684);
assign w3533 = w2696 & ~w3532;
assign w3534 = w6 & ~w3533;
assign w3535 = ~pi0034 & w2667;
assign w3536 = pi0079 & ~w3535;
assign w3537 = ~pi0118 & w2671;
assign w3538 = ~pi0079 & ~w3537;
assign w3539 = ~pi0954 & w3538;
assign w3540 = ~pi0033 & w3539;
assign w3541 = ~pi0034 & w3540;
assign w3542 = ~w3536 & ~w3541;
assign w3543 = ~w3534 & ~w3542;
assign w3544 = pi0189 & ~pi0299;
assign w3545 = pi0166 & pi0299;
assign w3546 = ~w3544 & ~w3545;
assign w3547 = w2695 & ~w3546;
assign w3548 = ~pi0175 & ~pi0299;
assign w3549 = pi0058 & pi0090;
assign w3550 = ~w367 & ~w3549;
assign w3551 = pi0153 & w3550;
assign w3552 = pi0299 & ~w3551;
assign w3553 = ~pi0095 & w3552;
assign w3554 = ~w3548 & ~w3553;
assign w3555 = w2623 & ~w3554;
assign w3556 = ~w3547 & ~w3555;
assign w3557 = pi0182 & ~pi0299;
assign w3558 = pi0160 & pi0299;
assign w3559 = ~w3557 & ~w3558;
assign w3560 = w1387 & w3559;
assign w3561 = pi0032 & ~pi0299;
assign w3562 = (~pi0299 & ~w2594) | (~pi0299 & w3561) | (~w2594 & w3561);
assign w3563 = ~pi0184 & w3562;
assign w3564 = ~w3560 & ~w3563;
assign w3565 = ~pi0073 & ~pi0163;
assign w3566 = w3553 & w3565;
assign w3567 = w2483 & ~w3566;
assign w3568 = w3564 & w3567;
assign w3569 = w3556 & w3568;
assign w3570 = w3534 & ~w3569;
assign w3571 = ~w3543 & ~w3570;
assign w3572 = ~pi0039 & ~w3571;
assign w3573 = w1257 & ~w2637;
assign w3574 = ~pi0166 & w3573;
assign w3575 = w1259 & ~w1274;
assign w3576 = ~pi0189 & w3575;
assign w3577 = ~w3574 & ~w3576;
assign w3578 = w1478 & ~w3577;
assign w3579 = pi0156 & w3573;
assign w3580 = pi0179 & w3575;
assign w3581 = ~w3579 & ~w3580;
assign w3582 = w1237 & ~w3581;
assign w3583 = ~w3578 & ~w3582;
assign w3584 = w2483 & ~w3583;
assign w3585 = w2823 & w3584;
assign w3586 = pi0039 & ~w3585;
assign w3587 = w2699 & w2823;
assign w3588 = w3542 & ~w3587;
assign w3589 = w3586 & ~w3588;
assign w3590 = ~w2845 & w2847;
assign w3591 = ~w2844 & ~w3590;
assign w3592 = pi0163 & ~w3591;
assign w3593 = ~w2844 & ~w2847;
assign w3594 = ~w2845 & ~w3593;
assign w3595 = ~pi0163 & ~w3594;
assign w3596 = ~w3592 & ~w3595;
assign w3597 = pi0299 & ~w3596;
assign w3598 = ~pi0183 & ~w2867;
assign w3599 = ~pi0178 & w3598;
assign w3600 = ~w2868 & ~w3599;
assign w3601 = pi0184 & ~w3600;
assign w3602 = ~w2868 & ~w2870;
assign w3603 = ~w2867 & ~w3602;
assign w3604 = ~pi0184 & ~w3603;
assign w3605 = ~w3601 & ~w3604;
assign w3606 = ~pi0299 & ~w3605;
assign w3607 = ~w3597 & ~w3606;
assign w3608 = ~pi0468 & ~w147;
assign w3609 = ~pi0332 & w3608;
assign w3610 = pi0232 & w3609;
assign w3611 = ~w3607 & w3610;
assign w3612 = pi0187 & ~pi0299;
assign w3613 = pi0147 & pi0299;
assign w3614 = ~w3612 & ~w3613;
assign w3615 = ~pi0468 & ~w3614;
assign w3616 = ~pi0332 & w3615;
assign w3617 = pi0232 & w3616;
assign w3618 = ~pi0100 & ~w2;
assign w3619 = ~pi0075 & w3618;
assign w3620 = ~pi0074 & w3619;
assign w3621 = ~w3617 & w3620;
assign w3622 = ~w3611 & ~w3621;
assign w3623 = w532 & w3622;
assign w3624 = w1658 & w3623;
assign w3625 = w529 & w3624;
assign w3626 = ~pi0038 & w3625;
assign w3627 = ~w3589 & w3626;
assign w3628 = ~w3572 & w3627;
assign w3629 = ~pi0040 & w5;
assign w3630 = ~w2824 & w3629;
assign w3631 = pi0163 & w2819;
assign w3632 = w2483 & w3631;
assign w3633 = ~w2819 & w3542;
assign w3634 = ~w3632 & ~w3633;
assign w3635 = w532 & ~w3634;
assign w3636 = w3630 & ~w3635;
assign w3637 = pi0179 & ~pi0299;
assign w3638 = pi0156 & pi0299;
assign w3639 = ~w3637 & ~w3638;
assign w3640 = w2483 & ~w3639;
assign w3641 = w2918 & ~w3640;
assign w3642 = ~w171 & w532;
assign w3643 = ~w3641 & w3642;
assign w3644 = ~w2745 & ~w3643;
assign w3645 = ~w5 & ~w171;
assign w3646 = ~pi0040 & ~w3645;
assign w3647 = w3644 & w3646;
assign w3648 = ~w2918 & ~w3542;
assign w3649 = w3629 & w3648;
assign w3650 = w3622 & ~w3649;
assign w3651 = ~w3647 & w3650;
assign w3652 = w2824 & ~w3651;
assign w3653 = ~w3636 & ~w3652;
assign w3654 = w179 & ~w3653;
assign w3655 = ~w5 & ~w2824;
assign w3656 = w179 & ~w3655;
assign w3657 = pi0147 & w2483;
assign w3658 = ~pi0100 & ~w3657;
assign w3659 = ~pi0075 & w3658;
assign w3660 = ~pi0074 & w3659;
assign w3661 = w2755 & ~w3596;
assign w3662 = ~w3660 & ~w3661;
assign w3663 = ~w3656 & ~w3662;
assign w3664 = ~w3654 & ~w3663;
assign w3665 = ~w3628 & ~w3664;
assign w3666 = (~w2224 & w2225) | (~w2224 & w2229) | (w2225 & w2229);
assign w3667 = ~w2412 & w3666;
assign w3668 = w2414 & w3666;
assign w3669 = (~w2038 & w3667) | (~w2038 & w3668) | (w3667 & w3668);
assign w3670 = ~pi0080 & w2546;
assign w3671 = ~pi0087 & w2442;
assign w3672 = w492 & w3671;
assign w3673 = pi0087 & w196;
assign w3674 = w194 & w3673;
assign w3675 = ~w3672 & ~w3674;
assign w3676 = w2043 & ~w2546;
assign w3677 = (~w2040 & ~w2546) | (~w2040 & w3676) | (~w2546 & w3676);
assign w3678 = ~pi0080 & ~w3677;
assign w3679 = w5 & w529;
assign w3680 = ~pi0092 & w2525;
assign w3681 = w1641 & w3680;
assign w3682 = ~pi1091 & w1476;
assign w3683 = w3681 & w3682;
assign w3684 = w3679 & w3683;
assign w3685 = (~pi0080 & w3678) | (~pi0080 & w3684) | (w3678 & w3684);
assign w3686 = (~w3675 & w3678) | (~w3675 & w3685) | (w3678 & w3685);
assign w3687 = (w3669 & w3670) | (w3669 & w3686) | (w3670 & w3686);
assign w3688 = w2045 & w3687;
assign w3689 = pi0081 & ~pi0314;
assign w3690 = ~pi0068 & ~w3689;
assign w3691 = ~w3014 & ~w3018;
assign w3692 = ~w3690 & ~w3691;
assign w3693 = pi0069 & pi0314;
assign w3694 = pi0066 & ~pi0069;
assign w3695 = ~w3693 & ~w3694;
assign w3696 = w3014 & ~w3695;
assign w3697 = ~pi0103 & ~pi0314;
assign w3698 = w3420 & w3697;
assign w3699 = ~pi0073 & w78;
assign w3700 = w74 & w3699;
assign w3701 = w3012 & w3700;
assign w3702 = ~pi0067 & w3701;
assign w3703 = ~pi0068 & w3702;
assign w3704 = ~pi0071 & w3703;
assign w3705 = pi0084 & w3704;
assign w3706 = ~w3698 & ~w3705;
assign w3707 = ~pi0200 & ~pi0299;
assign w3708 = ~pi0199 & w3707;
assign w3709 = ~pi0211 & w3457;
assign w3710 = ~w3708 & ~w3709;
assign w3711 = w3415 & ~w3710;
assign w3712 = ~pi0314 & w3452;
assign w3713 = ~pi0067 & ~w3712;
assign w3714 = w3330 & ~w3713;
assign w3715 = w1237 & w3427;
assign w3716 = ~pi0083 & w3419;
assign w3717 = pi0103 & w3716;
assign w3718 = pi0314 & w3717;
assign w3719 = pi0104 & w2043;
assign w3720 = w2950 & w3014;
assign w3721 = w3719 & w3720;
assign w3722 = w1280 & w3018;
assign w3723 = pi0088 & w3722;
assign w3724 = pi0824 & w3723;
assign w3725 = ~pi1093 & w3724;
assign w3726 = ~w3721 & ~w3725;
assign w3727 = ~pi0070 & pi0841;
assign w3728 = pi0089 & w3727;
assign w3729 = ~pi0024 & pi0070;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = w3436 & ~w3730;
assign w3732 = ~pi1050 & w3436;
assign w3733 = pi0073 & w3732;
assign w3734 = pi0841 & w3360;
assign w3735 = ~w3733 & ~w3734;
assign w3736 = pi0024 & ~pi0036;
assign w3737 = ~w1236 & ~w3736;
assign w3738 = ~pi0036 & ~pi0091;
assign w3739 = w1379 & ~w3738;
assign w3740 = w1237 & w3475;
assign w3741 = ~w1470 & w3740;
assign w3742 = ~w3739 & ~w3741;
assign w3743 = ~w3737 & ~w3742;
assign w3744 = ~pi0039 & pi0092;
assign w3745 = w3479 & w3744;
assign w3746 = pi0039 & ~pi0092;
assign w3747 = w1271 & w3746;
assign w3748 = ~w3745 & ~w3747;
assign w3749 = w1297 & ~w3748;
assign w3750 = w5 & w3749;
assign w3751 = ~pi0087 & w3750;
assign w3752 = pi0841 & w3436;
assign w3753 = pi0093 & w3752;
assign w3754 = w5 & w1297;
assign w3755 = w118 & w3754;
assign w3756 = pi0092 & w3755;
assign w3757 = ~pi1050 & w3756;
assign w3758 = ~w3753 & ~w3757;
assign w3759 = pi0049 & ~pi0841;
assign w3760 = w3014 & w3759;
assign w3761 = pi0252 & w2485;
assign w3762 = ~w454 & w3761;
assign w3763 = w3276 & w3762;
assign w3764 = ~w3760 & ~w3763;
assign w3765 = ~pi0332 & ~pi0841;
assign w3766 = pi0089 & w3014;
assign w3767 = w3765 & w3766;
assign w3768 = w12 & w1255;
assign w3769 = ~w3440 & ~w3768;
assign w3770 = ~w2698 & ~w3769;
assign w3771 = w1649 & w3770;
assign w3772 = ~w3443 & w3771;
assign w3773 = pi0024 & w1360;
assign w3774 = ~w3772 & ~w3773;
assign w3775 = ~w3767 & w3774;
assign w3776 = pi0479 & ~w454;
assign w3777 = ~pi0841 & ~w3776;
assign w3778 = pi0096 & ~w3777;
assign w3779 = ~pi0095 & w3778;
assign w3780 = pi0095 & ~pi0096;
assign w3781 = ~pi0024 & w3780;
assign w3782 = ~w3779 & ~w3781;
assign w3783 = w3464 & ~w3782;
assign w3784 = w593 & w3783;
assign w3785 = ~pi0032 & w3784;
assign w3786 = ~pi0040 & w3785;
assign w3787 = ~pi0072 & w3786;
assign w3788 = pi0593 & ~w2698;
assign w3789 = w1649 & w3443;
assign w3790 = w3788 & w3789;
assign w3791 = ~w2568 & ~w3492;
assign w3792 = ~w1236 & ~w3791;
assign w3793 = w3005 & w3792;
assign w3794 = w3499 & w3793;
assign w3795 = ~w3790 & ~w3794;
assign w3796 = w378 & w3484;
assign w3797 = ~w3756 & ~w3796;
assign w3798 = pi1050 & ~w3797;
assign w3799 = pi0314 & w3798;
assign w3800 = w3140 & w3155;
assign w3801 = ~pi0041 & ~pi0099;
assign w3802 = w3800 & w3801;
assign w3803 = ~pi0041 & w3154;
assign w3804 = w3166 & w3803;
assign w3805 = pi0099 & ~w3804;
assign w3806 = ~w3802 & ~w3805;
assign w3807 = w2525 & ~w3806;
assign w3808 = pi0174 & w526;
assign w3809 = ~pi0189 & w3808;
assign w3810 = pi0144 & w3809;
assign w3811 = pi0152 & ~w526;
assign w3812 = ~pi0166 & w3811;
assign w3813 = pi0161 & w3812;
assign w3814 = ~w3810 & ~w3813;
assign w3815 = w1645 & ~w3814;
assign w3816 = w3224 & w3815;
assign w3817 = ~w3807 & ~w3816;
assign w3818 = pi0129 & ~w2572;
assign w3819 = ~w2573 & ~w3818;
assign w3820 = w2571 & ~w2950;
assign w3821 = pi0683 & ~w3820;
assign w3822 = pi0252 & ~w3821;
assign w3823 = ~pi0683 & ~w2571;
assign w3824 = ~w3822 & ~w3823;
assign w3825 = w2485 & ~w3824;
assign w3826 = ~w3819 & ~w3825;
assign w3827 = w134 & ~w3826;
assign w3828 = w454 & w2582;
assign w3829 = ~w3827 & ~w3828;
assign w3830 = w1622 & ~w3829;
assign w3831 = pi0101 & ~w3220;
assign w3832 = ~w3800 & ~w3831;
assign w3833 = w2525 & ~w3832;
assign w3834 = ~pi0144 & w3809;
assign w3835 = ~pi0161 & w3812;
assign w3836 = ~w3834 & ~w3835;
assign w3837 = w1645 & ~w3836;
assign w3838 = w3224 & w3837;
assign w3839 = ~w3833 & ~w3838;
assign w3840 = pi0065 & w3018;
assign w3841 = ~pi0109 & ~w1404;
assign w3842 = w3436 & ~w3841;
assign w3843 = pi0104 & w2950;
assign w3844 = ~w2043 & w3014;
assign w3845 = w3843 & w3844;
assign w3846 = w2485 & w2950;
assign w3847 = w98 & w3267;
assign w3848 = pi0110 & w3847;
assign w3849 = ~w3846 & w3848;
assign w3850 = ~w3845 & ~w3849;
assign w3851 = ~pi0024 & w3319;
assign w3852 = pi0841 & w3332;
assign w3853 = ~w3851 & ~w3852;
assign w3854 = ~pi0999 & w3399;
assign w3855 = pi0108 & ~w3061;
assign w3856 = ~pi0098 & ~w3855;
assign w3857 = w254 & w376;
assign w3858 = w3005 & w3857;
assign w3859 = ~w3856 & w3858;
assign w3860 = pi0051 & ~pi0087;
assign w3861 = ~pi0051 & pi0087;
assign w3862 = ~w3860 & ~w3861;
assign w3863 = w2525 & ~w3862;
assign w3864 = w1345 & w3863;
assign w3865 = w3082 & w3864;
assign w3866 = ~w3859 & ~w3865;
assign w3867 = pi0077 & w1379;
assign w3868 = pi0314 & w3867;
assign w3869 = w2950 & w3848;
assign w3870 = w2485 & w3869;
assign w3871 = ~pi0082 & w3293;
assign w3872 = pi0111 & w3871;
assign w3873 = pi0314 & w3872;
assign w3874 = ~w3870 & ~w3873;
assign w3875 = ~pi0024 & w1641;
assign w3876 = pi0072 & w3875;
assign w3877 = w593 & w3876;
assign w3878 = w3464 & w3877;
assign w3879 = ~pi0314 & w3872;
assign w3880 = ~w3878 & ~w3879;
assign w3881 = pi0124 & ~pi0468;
assign w3882 = ~pi0099 & ~pi0113;
assign w3883 = ~pi0041 & w3882;
assign w3884 = w3800 & w3883;
assign w3885 = pi0113 & ~w3802;
assign w3886 = ~w3884 & ~w3885;
assign w3887 = w2525 & ~w3886;
assign w3888 = ~pi0114 & ~pi0116;
assign w3889 = w1318 & w3166;
assign w3890 = ~pi0115 & w3889;
assign w3891 = w3888 & w3890;
assign w3892 = ~pi0115 & ~pi0116;
assign w3893 = w3889 & w3892;
assign w3894 = pi0114 & ~w3893;
assign w3895 = ~w3891 & ~w3894;
assign w3896 = w2525 & ~w3895;
assign w3897 = ~pi0116 & w3889;
assign w3898 = pi0115 & ~w3897;
assign w3899 = ~w3893 & ~w3898;
assign w3900 = w2525 & ~w3899;
assign w3901 = pi0116 & ~w3889;
assign w3902 = ~w3897 & ~w3901;
assign w3903 = w2525 & ~w3902;
assign w3904 = ~w603 & ~w1665;
assign w3905 = ~w526 & w2824;
assign w3906 = pi0165 & ~pi0468;
assign w3907 = w2482 & w3906;
assign w3908 = w147 & ~w3907;
assign w3909 = w2935 & w3908;
assign w3910 = pi0150 & w2844;
assign w3911 = (pi0150 & w3590) | (pi0150 & w3910) | (w3590 & w3910);
assign w3912 = ~pi0163 & w3911;
assign w3913 = ~pi0163 & ~w2845;
assign w3914 = ~w3593 & w3913;
assign w3915 = ~pi0150 & ~w3914;
assign w3916 = ~w3912 & ~w3915;
assign w3917 = ~w2755 & ~w3909;
assign w3918 = (~w3909 & w3916) | (~w3909 & w3917) | (w3916 & w3917);
assign w3919 = w3905 & w3918;
assign w3920 = pi0143 & ~pi0468;
assign w3921 = w2482 & w3920;
assign w3922 = w147 & ~w3921;
assign w3923 = w2935 & w3922;
assign w3924 = (~pi0140 & w2868) | (~pi0140 & w2870) | (w2868 & w2870);
assign w3925 = ~pi0145 & w2870;
assign w3926 = ~w3924 & ~w3925;
assign w3927 = pi0184 & ~pi0185;
assign w3928 = (~pi0185 & w3926) | (~pi0185 & w3927) | (w3926 & w3927);
assign w3929 = ~pi0184 & pi0185;
assign w3930 = ~w3926 & w3929;
assign w3931 = ~w3928 & ~w3930;
assign w3932 = ~w2755 & ~w3923;
assign w3933 = (~w3923 & w3931) | (~w3923 & w3932) | (w3931 & w3932);
assign w3934 = w526 & w3933;
assign w3935 = ~w3919 & ~w3934;
assign w3936 = ~pi0150 & pi0299;
assign w3937 = ~w2595 & w3936;
assign w3938 = ~pi0168 & pi0299;
assign w3939 = ~pi0190 & ~pi0299;
assign w3940 = ~w3938 & ~w3939;
assign w3941 = pi0073 & ~w3940;
assign w3942 = ~pi0185 & ~pi0299;
assign w3943 = ~pi0185 & w3561;
assign w3944 = (~w2594 & w3942) | (~w2594 & w3943) | (w3942 & w3943);
assign w3945 = ~w3941 & ~w3944;
assign w3946 = ~w3937 & w3945;
assign w3947 = ~pi0173 & ~pi0299;
assign w3948 = ~pi0151 & pi0299;
assign w3949 = ~w3947 & ~w3948;
assign w3950 = w2483 & w3949;
assign w3951 = ~w1387 & ~w3950;
assign w3952 = w3946 & ~w3951;
assign w3953 = ~w1387 & ~w2483;
assign w3954 = w3946 & ~w3953;
assign w3955 = (~w2623 & w3952) | (~w2623 & w3954) | (w3952 & w3954);
assign w3956 = w6 & ~w3955;
assign w3957 = ~w3533 & w3956;
assign w3958 = ~w2698 & w3746;
assign w3959 = ~w3744 & ~w3958;
assign w3960 = (w1270 & ~w3744) | (w1270 & w3959) | (~w3744 & w3959);
assign w3961 = ~pi0039 & ~pi0092;
assign w3962 = pi0038 & w3961;
assign w3963 = ~pi0087 & w3962;
assign w3964 = w113 & w3963;
assign w3965 = pi0038 & ~w3962;
assign w3966 = ~pi0087 & ~w3965;
assign w3967 = w113 & w3966;
assign w3968 = (~w3960 & w3964) | (~w3960 & w3967) | (w3964 & w3967);
assign w3969 = w147 & w168;
assign w3970 = ~pi0118 & ~pi0954;
assign w3971 = ~pi0079 & w3970;
assign w3972 = ~pi0033 & ~pi0034;
assign w3973 = ~w2671 & w3972;
assign w3974 = w3971 & w3973;
assign w3975 = ~pi0079 & ~pi0954;
assign w3976 = w3972 & w3975;
assign w3977 = pi0118 & ~w3976;
assign w3978 = ~pi0038 & w3977;
assign w3979 = (~pi0038 & w3974) | (~pi0038 & w3978) | (w3974 & w3978);
assign w3980 = ~pi0074 & w3979;
assign w3981 = ~pi0054 & w3980;
assign w3982 = w147 & w3981;
assign w3983 = (w3968 & w3969) | (w3968 & w3982) | (w3969 & w3982);
assign w3984 = ~w6 & w3983;
assign w3985 = (w3533 & w3983) | (w3533 & w3984) | (w3983 & w3984);
assign w3986 = ~w3957 & ~w3985;
assign w3987 = ~pi0178 & ~pi0299;
assign w3988 = ~pi0157 & pi0299;
assign w3989 = ~w3987 & ~w3988;
assign w3990 = w3744 & w3989;
assign w3991 = pi0157 & w1237;
assign w3992 = pi0168 & w1478;
assign w3993 = ~w3991 & ~w3992;
assign w3994 = w3573 & ~w3993;
assign w3995 = pi0178 & w1237;
assign w3996 = pi0190 & w1478;
assign w3997 = ~w3995 & ~w3996;
assign w3998 = w3575 & ~w3997;
assign w3999 = ~w3994 & ~w3998;
assign w4000 = ~w3746 & ~w3990;
assign w4001 = (~w3990 & w3999) | (~w3990 & w4000) | (w3999 & w4000);
assign w4002 = w1354 & w2483;
assign w4003 = w2701 & w4002;
assign w4004 = ~pi0087 & w4003;
assign w4005 = w2678 & ~w4004;
assign w4006 = (w2678 & w4001) | (w2678 & w4005) | (w4001 & w4005);
assign w4007 = ~w3935 & ~w4006;
assign w4008 = (~w3935 & w3986) | (~w3935 & w4007) | (w3986 & w4007);
assign w4009 = ~w3974 & ~w3977;
assign w4010 = ~w546 & w4009;
assign w4011 = (~w567 & w4009) | (~w567 & w4010) | (w4009 & w4010);
assign w4012 = pi0150 & ~pi0468;
assign w4013 = w2482 & w4012;
assign w4014 = w546 & w4013;
assign w4015 = w567 & w4014;
assign w4016 = ~w4011 & ~w4015;
assign w4017 = ~w529 & w3918;
assign w4018 = ~w529 & ~w2789;
assign w4019 = w3918 & w4018;
assign w4020 = (~w4016 & w4017) | (~w4016 & w4019) | (w4017 & w4019);
assign w4021 = ~w4008 & ~w4020;
assign w4022 = ~pi0228 & ~w3756;
assign w4023 = ~w135 & w1622;
assign w4024 = w1237 & ~w3474;
assign w4025 = w1649 & w4024;
assign w4026 = ~w4023 & ~w4025;
assign w4027 = ~pi0086 & ~pi0109;
assign w4028 = ~pi0077 & w4027;
assign w4029 = ~w1520 & ~w4028;
assign w4030 = pi0036 & pi0097;
assign w4031 = ~pi0036 & ~pi0097;
assign w4032 = ~w4030 & ~w4031;
assign w4033 = w1236 & w4032;
assign w4034 = ~pi0091 & ~w4033;
assign w4035 = ~pi0093 & w4034;
assign w4036 = ~w4029 & w4035;
assign w4037 = w593 & ~w4036;
assign w4038 = ~w2553 & w4037;
assign w4039 = w4026 & ~w4038;
assign w4040 = w4022 & w4039;
assign w4041 = ~pi0128 & pi0228;
assign w4042 = ~w4040 & ~w4041;
assign w4043 = w2040 & ~w2043;
assign w4044 = ~w2470 & ~w2539;
assign w4045 = w112 & w2443;
assign w4046 = ~w2433 & ~w4045;
assign w4047 = w2525 & ~w4046;
assign w4048 = w1284 & w1641;
assign w4049 = w4047 & w4048;
assign w4050 = ~pi0075 & ~w4049;
assign w4051 = ~w2524 & w4050;
assign w4052 = ~w4044 & w4051;
assign w4053 = w113 & ~w2492;
assign w4054 = w117 & w1302;
assign w4055 = w4053 & w4054;
assign w4056 = ~w2518 & ~w4055;
assign w4057 = w529 & ~w4056;
assign w4058 = ~w4052 & w4057;
assign w4059 = pi0818 & pi1093;
assign w4060 = ~pi0031 & ~pi0080;
assign w4061 = w4059 & w4060;
assign w4062 = ~pi0120 & ~w4061;
assign w4063 = w1475 & w2045;
assign w4064 = pi0951 & w4063;
assign w4065 = pi0982 & w4064;
assign w4066 = w4062 & ~w4065;
assign w4067 = ~w4058 & ~w4066;
assign w4068 = ~w4043 & w4067;
assign w4069 = pi0051 & ~pi0146;
assign w4070 = ~pi0051 & ~pi0161;
assign w4071 = ~w4069 & ~w4070;
assign w4072 = ~w526 & ~w4071;
assign w4073 = ~pi0051 & ~pi0144;
assign w4074 = pi0051 & ~pi0142;
assign w4075 = ~w4073 & ~w4074;
assign w4076 = w526 & ~w4075;
assign w4077 = ~w4072 & ~w4076;
assign w4078 = ~pi0087 & ~w4077;
assign w4079 = pi0163 & ~w525;
assign w4080 = (pi0163 & ~w180) | (pi0163 & w4079) | (~w180 & w4079);
assign w4081 = pi0184 & w525;
assign w4082 = w180 & w4081;
assign w4083 = ~w4080 & ~w4082;
assign w4084 = pi0087 & ~w4083;
assign w4085 = ~w1635 & w4084;
assign w4086 = (~w1635 & w4078) | (~w1635 & w4085) | (w4078 & w4085);
assign w4087 = pi0159 & w1257;
assign w4088 = pi0181 & w1259;
assign w4089 = ~w4087 & ~w4088;
assign w4090 = ~w4086 & w4089;
assign w4091 = (~w3040 & ~w4086) | (~w3040 & w4090) | (~w4086 & w4090);
assign w4092 = w2483 & ~w4091;
assign w4093 = pi0077 & pi0314;
assign w4094 = ~pi0024 & w4093;
assign w4095 = ~w2627 & w4094;
assign w4096 = w4091 & ~w4095;
assign w4097 = w2483 & ~w4096;
assign w4098 = (w3436 & w4092) | (w3436 & w4097) | (w4092 & w4097);
assign w4099 = w254 & ~w1433;
assign w4100 = ~pi0092 & w3679;
assign w4101 = w3497 & w4100;
assign w4102 = ~pi0024 & ~pi0314;
assign w4103 = ~pi0077 & ~pi0086;
assign w4104 = (~pi0086 & w4102) | (~pi0086 & w4103) | (w4102 & w4103);
assign w4105 = ~pi0039 & ~w4104;
assign w4106 = w4101 & w4105;
assign w4107 = w382 & w4106;
assign w4108 = ~pi0024 & pi0077;
assign w4109 = w4107 & ~w4108;
assign w4110 = w4099 & w4109;
assign w4111 = w3640 & w4110;
assign w4112 = ~pi0125 & ~pi0133;
assign w4113 = pi0121 & ~w4112;
assign w4114 = ~pi0134 & ~pi0135;
assign w4115 = ~pi0126 & ~pi0130;
assign w4116 = w4114 & w4115;
assign w4117 = ~pi0132 & ~pi0136;
assign w4118 = ~pi0125 & ~w4117;
assign w4119 = (~pi0125 & ~w4116) | (~pi0125 & w4118) | (~w4116 & w4118);
assign w4120 = ~pi0121 & ~pi0133;
assign w4121 = ~w4113 & ~w4120;
assign w4122 = (~w4113 & ~w4119) | (~w4113 & w4121) | (~w4119 & w4121);
assign w4123 = pi0039 & pi0072;
assign w4124 = pi0072 & ~w4123;
assign w4125 = ~w2525 & ~w4123;
assign w4126 = (~w1488 & w4124) | (~w1488 & w4125) | (w4124 & w4125);
assign w4127 = w4122 & ~w4126;
assign w4128 = (~w3082 & w4122) | (~w3082 & w4127) | (w4122 & w4127);
assign w4129 = ~w4107 & w4128;
assign w4130 = (~w4099 & w4128) | (~w4099 & w4129) | (w4128 & w4129);
assign w4131 = w1635 & w4130;
assign w4132 = (w1635 & w4111) | (w1635 & w4131) | (w4111 & w4131);
assign w4133 = ~w4098 & ~w4132;
assign w4134 = ~w4043 & ~w4058;
assign w4135 = ~pi0039 & pi0110;
assign w4136 = w2483 & ~w3229;
assign w4137 = w2950 & ~w4136;
assign w4138 = ~w2959 & w4137;
assign w4139 = w4135 & w4138;
assign w4140 = pi0039 & ~pi0110;
assign w4141 = w1630 & w4140;
assign w4142 = ~w4139 & ~w4141;
assign w4143 = (~pi0071 & ~w1425) | (~pi0071 & w1428) | (~w1425 & w1428);
assign w4144 = w1422 & w4143;
assign w4145 = ~pi0072 & w4144;
assign w4146 = ~pi0081 & w4145;
assign w4147 = ~pi0090 & w4146;
assign w4148 = ~pi0111 & w4147;
assign w4149 = w3436 & ~w4148;
assign w4150 = w4142 & ~w4149;
assign w4151 = ~w2793 & ~w2795;
assign w4152 = pi0087 & ~w4151;
assign w4153 = w2483 & w4152;
assign w4154 = w529 & ~w4153;
assign w4155 = w99 & w3699;
assign w4156 = w74 & w4155;
assign w4157 = w1638 & w1641;
assign w4158 = ~pi0072 & w4157;
assign w4159 = ~w1257 & ~w1259;
assign w4160 = w4158 & ~w4159;
assign w4161 = w5 & w4160;
assign w4162 = w4156 & w4161;
assign w4163 = w3746 & w4162;
assign w4164 = pi0051 & pi0193;
assign w4165 = ~pi0051 & ~pi0174;
assign w4166 = ~w4164 & ~w4165;
assign w4167 = (w1345 & ~w4164) | (w1345 & w4166) | (~w4164 & w4166);
assign w4168 = ~pi0299 & ~w4167;
assign w4169 = pi0051 & pi0172;
assign w4170 = ~pi0051 & ~pi0152;
assign w4171 = ~w4169 & ~w4170;
assign w4172 = (w1345 & ~w4169) | (w1345 & w4171) | (~w4169 & w4171);
assign w4173 = pi0299 & ~w4172;
assign w4174 = ~w4168 & ~w4173;
assign w4175 = w2483 & ~w4174;
assign w4176 = ~pi0121 & w4117;
assign w4177 = w4116 & w4176;
assign w4178 = ~pi0125 & pi0133;
assign w4179 = pi0133 & ~w4178;
assign w4180 = pi0125 & ~pi0133;
assign w4181 = ~w4178 & ~w4180;
assign w4182 = (~w4177 & w4179) | (~w4177 & w4181) | (w4179 & w4181);
assign w4183 = w1635 & ~w4182;
assign w4184 = ~pi0087 & w4183;
assign w4185 = (~pi0087 & w4175) | (~pi0087 & w4184) | (w4175 & w4184);
assign w4186 = w4154 & ~w4185;
assign w4187 = (w4154 & w4163) | (w4154 & w4186) | (w4163 & w4186);
assign w4188 = ~pi0174 & w1241;
assign w4189 = ~w1345 & w4188;
assign w4190 = pi0180 & ~pi0287;
assign w4191 = w1241 & w4190;
assign w4192 = ~pi0223 & ~pi0224;
assign w4193 = pi0222 & w4192;
assign w4194 = (w643 & w4191) | (w643 & w4193) | (w4191 & w4193);
assign w4195 = w1345 & w4194;
assign w4196 = w4158 & w4195;
assign w4197 = ~w4189 & ~w4196;
assign w4198 = (~w4156 & ~w4189) | (~w4156 & w4197) | (~w4189 & w4197);
assign w4199 = pi0051 & ~pi0193;
assign w4200 = (pi0051 & ~w1241) | (pi0051 & w4199) | (~w1241 & w4199);
assign w4201 = ~pi0299 & w4200;
assign w4202 = pi0051 & ~w4200;
assign w4203 = ~pi0299 & ~w4202;
assign w4204 = (w4198 & w4201) | (w4198 & w4203) | (w4201 & w4203);
assign w4205 = pi0232 & ~pi0299;
assign w4206 = pi0299 & ~w1241;
assign w4207 = pi0232 & ~w4206;
assign w4208 = (~w4172 & w4205) | (~w4172 & w4207) | (w4205 & w4207);
assign w4209 = pi0158 & ~pi0215;
assign w4210 = w1241 & w4209;
assign w4211 = pi0221 & pi0232;
assign w4212 = ~pi0287 & w4211;
assign w4213 = w4210 & w4212;
assign w4214 = w1470 & ~w4213;
assign w4215 = w109 & ~w4214;
assign w4216 = w112 & w4215;
assign w4217 = ~w4208 & ~w4216;
assign w4218 = ~w4204 & ~w4217;
assign w4219 = pi0039 & ~w4218;
assign w4220 = ~pi0072 & w4104;
assign w4221 = w3052 & ~w4220;
assign w4222 = ~w3055 & ~w4220;
assign w4223 = (~w3054 & w4221) | (~w3054 & w4222) | (w4221 & w4222);
assign w4224 = pi0039 & ~w4219;
assign w4225 = (~w4219 & w4223) | (~w4219 & w4224) | (w4223 & w4224);
assign w4226 = w5 & w171;
assign w4227 = w4187 & ~w4226;
assign w4228 = (w4187 & ~w4225) | (w4187 & w4227) | (~w4225 & w4227);
assign w4229 = pi0087 & pi0162;
assign w4230 = w2483 & w4229;
assign w4231 = pi0087 & ~w4229;
assign w4232 = w2483 & ~w4231;
assign w4233 = (~w4172 & w4230) | (~w4172 & w4232) | (w4230 & w4232);
assign w4234 = ~w529 & ~w4233;
assign w4235 = ~w4183 & w4234;
assign w4236 = ~pi0092 & w349;
assign w4237 = w3679 & w4236;
assign w4238 = w382 & ~w4104;
assign w4239 = ~pi0035 & w4238;
assign w4240 = w4237 & w4239;
assign w4241 = w254 & w4240;
assign w4242 = ~w1433 & w4241;
assign w4243 = ~pi0024 & ~pi0086;
assign w4244 = ~w2921 & ~w4243;
assign w4245 = pi0145 & ~pi0299;
assign w4246 = pi0197 & pi0299;
assign w4247 = ~w4245 & ~w4246;
assign w4248 = w4243 & ~w4247;
assign w4249 = ~w4244 & ~w4248;
assign w4250 = w2483 & ~w4249;
assign w4251 = w6 & ~w4250;
assign w4252 = ~w4235 & ~w4251;
assign w4253 = (~w4235 & ~w4242) | (~w4235 & w4252) | (~w4242 & w4252);
assign w4254 = ~w4228 & w4253;
assign w4255 = w6 & w4242;
assign w4256 = w4116 & w4117;
assign w4257 = ~pi0121 & w4112;
assign w4258 = pi0126 & ~w4257;
assign w4259 = ~pi0126 & ~pi0133;
assign w4260 = ~pi0121 & ~pi0125;
assign w4261 = w4259 & w4260;
assign w4262 = ~w4258 & ~w4261;
assign w4263 = ~w4256 & ~w4262;
assign w4264 = w1635 & w4263;
assign w4265 = ~w4255 & ~w4264;
assign w4266 = (~pi0072 & w1488) | (~pi0072 & w2525) | (w1488 & w2525);
assign w4267 = w3082 & ~w4266;
assign w4268 = ~w4265 & ~w4267;
assign w4269 = ~pi0182 & w1259;
assign w4270 = ~pi0287 & w2483;
assign w4271 = ~w4269 & w4270;
assign w4272 = pi0160 & w4271;
assign w4273 = pi0182 & w4270;
assign w4274 = w1259 & ~w4273;
assign w4275 = ~w1257 & ~w4274;
assign w4276 = ~w4272 & ~w4275;
assign w4277 = ~pi0072 & w4276;
assign w4278 = pi0072 & w4263;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = pi0039 & ~w4279;
assign w4281 = w3082 & w4280;
assign w4282 = ~w4268 & ~w4281;
assign w4283 = ~pi0051 & ~pi0166;
assign w4284 = pi0051 & pi0153;
assign w4285 = ~w4283 & ~w4284;
assign w4286 = w2483 & ~w4285;
assign w4287 = ~w529 & w4286;
assign w4288 = ~pi0087 & w4287;
assign w4289 = ~w1635 & ~w4288;
assign w4290 = w4282 & ~w4289;
assign w4291 = ~w2800 & w4243;
assign w4292 = ~w3989 & ~w4243;
assign w4293 = ~w4291 & ~w4292;
assign w4294 = w4255 & w4293;
assign w4295 = ~pi0087 & w529;
assign w4296 = ~pi0051 & ~w1345;
assign w4297 = w3546 & w4296;
assign w4298 = pi0175 & ~pi0299;
assign w4299 = pi0153 & pi0299;
assign w4300 = ~w4298 & ~w4299;
assign w4301 = pi0051 & ~w4300;
assign w4302 = ~w4297 & ~w4301;
assign w4303 = w4295 & ~w4302;
assign w4304 = pi0185 & w526;
assign w4305 = pi0150 & ~w526;
assign w4306 = ~w4304 & ~w4305;
assign w4307 = pi0087 & ~w4306;
assign w4308 = ~w4303 & ~w4307;
assign w4309 = ~w4294 & w4308;
assign w4310 = w2483 & ~w4309;
assign w4311 = ~w4290 & ~w4310;
assign w4312 = ~pi0063 & w1378;
assign w4313 = w3393 & ~w4312;
assign w4314 = (w1377 & w3393) | (w1377 & w4313) | (w3393 & w4313);
assign w4315 = pi0129 & ~w4314;
assign w4316 = pi0250 & pi0252;
assign w4317 = ~pi0127 & ~w4316;
assign w4318 = (~pi0127 & ~w2485) | (~pi0127 & w4317) | (~w2485 & w4317);
assign w4319 = w2568 & w4316;
assign w4320 = w2485 & w4319;
assign w4321 = ~w4318 & ~w4320;
assign w4322 = pi0094 & ~w4321;
assign w4323 = w4315 & ~w4322;
assign w4324 = pi0129 & ~w3761;
assign w4325 = pi0075 & ~w4324;
assign w4326 = ~pi0100 & ~w4325;
assign w4327 = ~pi0100 & ~w3761;
assign w4328 = ~pi0250 & ~w4327;
assign w4329 = ~w2568 & w4328;
assign w4330 = ~w4326 & ~w4329;
assign w4331 = ~w1323 & w4330;
assign w4332 = ~w3393 & ~w4331;
assign w4333 = ~w2554 & ~w4332;
assign w4334 = ~pi0092 & w5;
assign w4335 = ~pi0039 & ~w4223;
assign w4336 = pi0140 & w1486;
assign w4337 = pi0162 & w1487;
assign w4338 = ~w4336 & ~w4337;
assign w4339 = w4270 & ~w4338;
assign w4340 = w1470 & ~w4339;
assign w4341 = w113 & ~w4340;
assign w4342 = pi0039 & ~w4341;
assign w4343 = ~w4335 & ~w4342;
assign w4344 = w4334 & w4343;
assign w4345 = pi0130 & ~pi0132;
assign w4346 = ~pi0126 & w4260;
assign w4347 = ~pi0133 & w4346;
assign w4348 = w4345 & w4347;
assign w4349 = ~pi0132 & w4347;
assign w4350 = ~pi0136 & w4114;
assign w4351 = w4349 & ~w4350;
assign w4352 = ~pi0130 & ~w4351;
assign w4353 = ~w4348 & ~w4352;
assign w4354 = w1345 & ~w4353;
assign w4355 = ~w4163 & w4354;
assign w4356 = ~w1345 & w2760;
assign w4357 = ~w4355 & ~w4356;
assign w4358 = w1634 & w4357;
assign w4359 = w529 & w4358;
assign w4360 = ~w4344 & w4359;
assign w4361 = pi0169 & ~w1345;
assign w4362 = ~pi0087 & ~w4361;
assign w4363 = w2483 & ~w4362;
assign w4364 = ~pi0051 & ~w4363;
assign w4365 = ~w4354 & w4364;
assign w4366 = ~w529 & w4365;
assign w4367 = ~pi0188 & w526;
assign w4368 = ~pi0167 & ~w526;
assign w4369 = ~w4367 & ~w4368;
assign w4370 = w2483 & w4369;
assign w4371 = pi0087 & ~w4370;
assign w4372 = ~w4366 & ~w4371;
assign w4373 = ~w4360 & w4372;
assign w4374 = ~w3756 & ~w4038;
assign w4375 = w4026 & w4374;
assign w4376 = w4099 & w4107;
assign w4377 = w6 & ~w4108;
assign w4378 = w4376 & ~w4377;
assign w4379 = ~pi0039 & pi0072;
assign w4380 = ~w1645 & ~w4379;
assign w4381 = w3082 & ~w4380;
assign w4382 = ~pi0072 & w1470;
assign w4383 = w4381 & ~w4382;
assign w4384 = ~w4256 & w4349;
assign w4385 = pi0132 & ~w4347;
assign w4386 = ~w4384 & ~w4385;
assign w4387 = ~w4383 & ~w4386;
assign w4388 = w3082 & ~w4159;
assign w4389 = w1645 & w4388;
assign w4390 = ~w4387 & ~w4389;
assign w4391 = ~w4381 & ~w4386;
assign w4392 = pi0183 & w1486;
assign w4393 = pi0149 & w1487;
assign w4394 = ~w4392 & ~w4393;
assign w4395 = w4270 & ~w4394;
assign w4396 = ~w4391 & w4395;
assign w4397 = ~w4390 & ~w4396;
assign w4398 = w1635 & ~w4397;
assign w4399 = ~w4376 & ~w4398;
assign w4400 = ~w4378 & ~w4399;
assign w4401 = w1635 & ~w3559;
assign w4402 = w4376 & w4401;
assign w4403 = pi0164 & ~w526;
assign w4404 = pi0186 & w526;
assign w4405 = ~w4403 & ~w4404;
assign w4406 = pi0087 & ~w4405;
assign w4407 = ~pi0051 & ~pi0168;
assign w4408 = pi0051 & ~pi0151;
assign w4409 = ~w4407 & ~w4408;
assign w4410 = ~w526 & ~w4409;
assign w4411 = pi0051 & ~pi0173;
assign w4412 = ~pi0051 & ~pi0190;
assign w4413 = ~w4411 & ~w4412;
assign w4414 = w526 & ~w4413;
assign w4415 = ~w4410 & ~w4414;
assign w4416 = ~pi0087 & w4415;
assign w4417 = ~w4406 & ~w4416;
assign w4418 = ~w1635 & ~w4417;
assign w4419 = ~w4402 & ~w4418;
assign w4420 = w2483 & ~w4419;
assign w4421 = ~w4400 & ~w4420;
assign w4422 = ~pi0154 & pi0299;
assign w4423 = ~pi0176 & ~pi0299;
assign w4424 = ~w4422 & ~w4423;
assign w4425 = w2483 & w4424;
assign w4426 = ~w4243 & ~w4425;
assign w4427 = w4255 & ~w4426;
assign w4428 = pi0145 & w1486;
assign w4429 = pi0197 & w1487;
assign w4430 = ~w4428 & ~w4429;
assign w4431 = w4270 & ~w4430;
assign w4432 = w4382 & ~w4431;
assign w4433 = w1635 & ~w4432;
assign w4434 = w4381 & w4433;
assign w4435 = ~w4427 & ~w4434;
assign w4436 = ~pi0125 & w4256;
assign w4437 = ~pi0121 & w4436;
assign w4438 = ~pi0133 & ~w4437;
assign w4439 = w1645 & ~w4159;
assign w4440 = w3082 & w4439;
assign w4441 = w1635 & ~w4440;
assign w4442 = ~w4438 & w4441;
assign w4443 = pi0149 & ~w526;
assign w4444 = pi0183 & w526;
assign w4445 = ~w4443 & ~w4444;
assign w4446 = w2483 & ~w4445;
assign w4447 = pi0087 & w4446;
assign w4448 = ~w4442 & ~w4447;
assign w4449 = ~w4255 & ~w4448;
assign w4450 = w4435 & ~w4449;
assign w4451 = w3082 & ~w4123;
assign w4452 = ~pi0135 & ~pi0136;
assign w4453 = w4347 & w4452;
assign w4454 = ~pi0130 & ~pi0132;
assign w4455 = w4453 & w4454;
assign w4456 = pi0134 & ~w4455;
assign w4457 = ~w4451 & w4456;
assign w4458 = pi0039 & ~w1488;
assign w4459 = w3082 & w4458;
assign w4460 = ~w4456 & ~w4459;
assign w4461 = pi0186 & w1486;
assign w4462 = pi0164 & w1487;
assign w4463 = ~w4461 & ~w4462;
assign w4464 = w4270 & ~w4463;
assign w4465 = w1470 & ~w4464;
assign w4466 = ~w4460 & w4465;
assign w4467 = ~pi0039 & w4456;
assign w4468 = ~w4466 & ~w4467;
assign w4469 = ~pi0072 & ~w4468;
assign w4470 = ~w4457 & ~w4469;
assign w4471 = w1345 & ~w4470;
assign w4472 = pi0192 & w526;
assign w4473 = pi0171 & ~w526;
assign w4474 = ~w4472 & ~w4473;
assign w4475 = w2483 & ~w4474;
assign w4476 = ~w1345 & ~w4475;
assign w4477 = ~w4471 & ~w4476;
assign w4478 = w1634 & ~w4477;
assign w4479 = ~w4376 & w4478;
assign w4480 = ~w4159 & w4381;
assign w4481 = pi0134 & w4454;
assign w4482 = w4453 & w4481;
assign w4483 = ~pi0136 & w4347;
assign w4484 = w4454 & w4483;
assign w4485 = pi0135 & ~w4484;
assign w4486 = ~w4482 & ~w4485;
assign w4487 = ~w4480 & w4486;
assign w4488 = pi0185 & w1486;
assign w4489 = pi0150 & w1487;
assign w4490 = ~w4488 & ~w4489;
assign w4491 = w4270 & ~w4490;
assign w4492 = ~w4487 & ~w4491;
assign w4493 = w4382 & w4492;
assign w4494 = ~w4381 & ~w4486;
assign w4495 = ~w4493 & ~w4494;
assign w4496 = w1345 & ~w4495;
assign w4497 = pi0194 & w526;
assign w4498 = pi0170 & ~w526;
assign w4499 = ~w4497 & ~w4498;
assign w4500 = w2483 & ~w4499;
assign w4501 = ~w1345 & ~w4500;
assign w4502 = ~w4496 & ~w4501;
assign w4503 = w1634 & ~w4502;
assign w4504 = ~w4376 & w4503;
assign w4505 = w4100 & ~w4335;
assign w4506 = w2483 & ~w2882;
assign w4507 = ~w1345 & w4506;
assign w4508 = w4156 & w4158;
assign w4509 = pi0184 & w1486;
assign w4510 = pi0163 & w1487;
assign w4511 = ~w4509 & ~w4510;
assign w4512 = w4270 & ~w4511;
assign w4513 = w1470 & ~w4512;
assign w4514 = w4508 & ~w4513;
assign w4515 = pi0039 & ~w4514;
assign w4516 = w1345 & ~w4515;
assign w4517 = ~w4507 & ~w4516;
assign w4518 = w4505 & ~w4517;
assign w4519 = pi0148 & ~w526;
assign w4520 = pi0141 & w526;
assign w4521 = ~w4519 & ~w4520;
assign w4522 = ~w1345 & ~w4521;
assign w4523 = w2483 & w4522;
assign w4524 = ~pi0130 & w4117;
assign w4525 = ~w4114 & w4347;
assign w4526 = w4524 & w4525;
assign w4527 = w4347 & w4454;
assign w4528 = pi0136 & ~w4527;
assign w4529 = ~w4526 & ~w4528;
assign w4530 = w1345 & w4529;
assign w4531 = ~w4523 & ~w4530;
assign w4532 = ~w4389 & ~w4531;
assign w4533 = ~w4518 & ~w4532;
assign w4534 = w1634 & w4533;
assign w4535 = ~pi0039 & pi0137;
assign w4536 = pi0039 & ~w3204;
assign w4537 = ~pi0198 & w526;
assign w4538 = w3225 & w4537;
assign w4539 = ~pi0210 & ~w526;
assign w4540 = w3227 & w4539;
assign w4541 = ~w4538 & ~w4540;
assign w4542 = w2483 & ~w4541;
assign w4543 = w4536 & w4542;
assign w4544 = ~w4535 & ~w4543;
assign w4545 = w3486 & w4506;
assign w4546 = ~w2594 & w3052;
assign w4547 = ~w2594 & ~w3055;
assign w4548 = (~w3054 & w4546) | (~w3054 & w4547) | (w4546 & w4547);
assign w4549 = pi0039 & w1237;
assign w4550 = ~w1270 & w4549;
assign w4551 = w2823 & w4550;
assign w4552 = pi0039 & ~w4551;
assign w4553 = w2621 & ~w2689;
assign w4554 = (~w1396 & ~w2689) | (~w1396 & w4553) | (~w2689 & w4553);
assign w4555 = ~pi0039 & w4554;
assign w4556 = ~w4551 & ~w4555;
assign w4557 = (~w4548 & w4552) | (~w4548 & w4556) | (w4552 & w4556);
assign w4558 = ~w4545 & w4557;
assign w4559 = w1481 & ~w4558;
assign w4560 = w2701 & w2817;
assign w4561 = pi0055 & w546;
assign w4562 = w4560 & w4561;
assign w4563 = ~w1619 & ~w4562;
assign w4564 = w2789 & w4563;
assign w4565 = ~pi0138 & ~w2670;
assign w4566 = ~pi0034 & w2673;
assign w4567 = ~pi0139 & w4566;
assign w4568 = ~pi0954 & w4567;
assign w4569 = w4565 & w4568;
assign w4570 = pi0138 & ~w4568;
assign w4571 = ~w4569 & ~w4570;
assign w4572 = w4564 & ~w4571;
assign w4573 = ~w3486 & ~w4572;
assign w4574 = ~w4559 & ~w4573;
assign w4575 = pi0139 & ~w2899;
assign w4576 = (pi0139 & ~w2673) | (pi0139 & w4575) | (~w2673 & w4575);
assign w4577 = ~pi0139 & ~pi0954;
assign w4578 = ~pi0034 & w4577;
assign w4579 = w2673 & w4578;
assign w4580 = ~w4576 & ~w4579;
assign w4581 = ~w2671 & ~w4580;
assign w4582 = w2789 & w4581;
assign w4583 = w4563 & w4582;
assign w4584 = w1658 & w2824;
assign w4585 = w4583 & ~w4584;
assign w4586 = (w4557 & w4583) | (w4557 & w4585) | (w4583 & w4585);
assign w4587 = ~w3486 & ~w4586;
assign w4588 = w2760 & ~w3485;
assign w4589 = w378 & w4588;
assign w4590 = ~w4587 & ~w4589;
assign w4591 = pi0665 & pi1091;
assign w4592 = pi0628 & pi1156;
assign w4593 = ~pi0628 & ~pi1156;
assign w4594 = ~w4592 & ~w4593;
assign w4595 = pi0792 & w4594;
assign w4596 = ~pi0715 & pi1160;
assign w4597 = pi0715 & ~pi1160;
assign w4598 = ~w4596 & ~w4597;
assign w4599 = pi0790 & ~w4598;
assign w4600 = ~pi0648 & pi1159;
assign w4601 = pi0648 & ~pi1159;
assign w4602 = ~w4600 & ~w4601;
assign w4603 = pi0789 & ~w4602;
assign w4604 = ~w4599 & ~w4603;
assign w4605 = ~w4595 & w4604;
assign w4606 = pi0625 & pi1153;
assign w4607 = ~pi0625 & ~pi1153;
assign w4608 = ~w4606 & ~w4607;
assign w4609 = pi0778 & w4608;
assign w4610 = ~pi0641 & pi1158;
assign w4611 = pi0641 & ~pi1158;
assign w4612 = ~w4610 & ~w4611;
assign w4613 = pi0788 & ~w4612;
assign w4614 = pi0647 & ~pi1157;
assign w4615 = ~pi0647 & pi1157;
assign w4616 = ~w4614 & ~w4615;
assign w4617 = pi0787 & ~w4616;
assign w4618 = ~w4613 & ~w4617;
assign w4619 = ~w4609 & w4618;
assign w4620 = ~pi0660 & pi1155;
assign w4621 = pi0660 & ~pi1155;
assign w4622 = ~w4620 & ~w4621;
assign w4623 = pi0785 & ~w4622;
assign w4624 = ~pi0627 & pi1154;
assign w4625 = pi0627 & ~pi1154;
assign w4626 = ~w4624 & ~w4625;
assign w4627 = pi0781 & ~w4626;
assign w4628 = ~w4623 & ~w4627;
assign w4629 = w4619 & w4628;
assign w4630 = pi0680 & w4629;
assign w4631 = w4605 & w4630;
assign w4632 = ~w4591 & w4631;
assign w4633 = pi0621 & pi1091;
assign w4634 = pi0629 & pi1156;
assign w4635 = ~pi0629 & ~pi1156;
assign w4636 = ~w4634 & ~w4635;
assign w4637 = pi0792 & w4636;
assign w4638 = ~pi0644 & pi1160;
assign w4639 = pi0644 & ~pi1160;
assign w4640 = ~w4638 & ~w4639;
assign w4641 = pi0790 & ~w4640;
assign w4642 = ~pi0619 & pi1159;
assign w4643 = pi0619 & ~pi1159;
assign w4644 = ~w4642 & ~w4643;
assign w4645 = pi0789 & ~w4644;
assign w4646 = ~w4641 & ~w4645;
assign w4647 = ~w4637 & w4646;
assign w4648 = pi0630 & pi1157;
assign w4649 = ~pi0630 & ~pi1157;
assign w4650 = ~w4648 & ~w4649;
assign w4651 = pi0787 & w4650;
assign w4652 = pi0603 & ~w4651;
assign w4653 = ~pi0618 & pi1154;
assign w4654 = pi0618 & ~pi1154;
assign w4655 = ~w4653 & ~w4654;
assign w4656 = pi0781 & ~w4655;
assign w4657 = ~pi0608 & pi1153;
assign w4658 = pi0608 & ~pi1153;
assign w4659 = ~w4657 & ~w4658;
assign w4660 = pi0778 & ~w4659;
assign w4661 = ~w4656 & ~w4660;
assign w4662 = w4652 & w4661;
assign w4663 = ~pi0626 & pi1158;
assign w4664 = pi0626 & ~pi1158;
assign w4665 = ~w4663 & ~w4664;
assign w4666 = pi0788 & ~w4665;
assign w4667 = ~pi0609 & pi1155;
assign w4668 = pi0609 & ~pi1155;
assign w4669 = ~w4667 & ~w4668;
assign w4670 = pi0785 & ~w4669;
assign w4671 = ~w4666 & ~w4670;
assign w4672 = w4662 & w4671;
assign w4673 = w4647 & w4672;
assign w4674 = ~w4633 & w4673;
assign w4675 = w4632 & ~w4674;
assign w4676 = ~pi0738 & w4675;
assign w4677 = ~pi0761 & w4674;
assign w4678 = ~w4676 & ~w4677;
assign w4679 = pi0108 & pi0314;
assign w4680 = ~pi0102 & ~w4679;
assign w4681 = ~pi0045 & w4680;
assign w4682 = pi0040 & w4681;
assign w4683 = ~pi0252 & ~w4682;
assign w4684 = w3700 & w4683;
assign w4685 = ~pi0040 & ~w2992;
assign w4686 = ~pi0047 & w4685;
assign w4687 = w4681 & w4686;
assign w4688 = ~w4684 & ~w4687;
assign w4689 = ~w3467 & ~w4688;
assign w4690 = ~w205 & ~w4689;
assign w4691 = ~w2553 & w4690;
assign w4692 = ~w1649 & ~w4691;
assign w4693 = w193 & w3071;
assign w4694 = w1284 & w4693;
assign w4695 = w192 & w196;
assign w4696 = w4694 & w4695;
assign w4697 = ~pi0038 & ~w4696;
assign w4698 = ~pi0832 & w4697;
assign w4699 = w4692 & w4698;
assign w4700 = ~w2698 & ~w3474;
assign w4701 = w1233 & w1284;
assign w4702 = w1278 & w1291;
assign w4703 = w4701 & w4702;
assign w4704 = ~pi0287 & ~w3026;
assign w4705 = ~pi0120 & ~w4704;
assign w4706 = ~w4703 & ~w4705;
assign w4707 = ~w4700 & ~w4706;
assign w4708 = w1649 & ~w4707;
assign w4709 = pi0038 & ~w113;
assign w4710 = ~pi0039 & w1481;
assign w4711 = ~w4709 & w4710;
assign w4712 = ~pi0832 & ~w4711;
assign w4713 = ~w4708 & w4712;
assign w4714 = w1475 & ~w4713;
assign w4715 = ~w4699 & w4714;
assign w4716 = ~w4678 & w4715;
assign w4717 = ~pi0140 & ~w4715;
assign w4718 = ~w4716 & ~w4717;
assign w4719 = pi0706 & w4675;
assign w4720 = pi0749 & w4674;
assign w4721 = ~w4719 & ~w4720;
assign w4722 = w4715 & ~w4721;
assign w4723 = ~pi0141 & ~w4715;
assign w4724 = ~w4722 & ~w4723;
assign w4725 = pi0735 & w4675;
assign w4726 = pi0743 & w4674;
assign w4727 = ~w4725 & ~w4726;
assign w4728 = w4715 & ~w4727;
assign w4729 = pi0142 & ~w4715;
assign w4730 = ~w4728 & ~w4729;
assign w4731 = pi0687 & w4675;
assign w4732 = ~pi0774 & w4674;
assign w4733 = ~w4731 & ~w4732;
assign w4734 = w4715 & ~w4733;
assign w4735 = ~pi0143 & ~w4715;
assign w4736 = ~w4734 & ~w4735;
assign w4737 = pi0736 & w4675;
assign w4738 = pi0758 & w4674;
assign w4739 = ~w4737 & ~w4738;
assign w4740 = w4715 & ~w4739;
assign w4741 = pi0144 & ~w4715;
assign w4742 = ~w4740 & ~w4741;
assign w4743 = ~pi0698 & w4675;
assign w4744 = ~pi0767 & w4674;
assign w4745 = ~w4743 & ~w4744;
assign w4746 = w4715 & ~w4745;
assign w4747 = ~pi0145 & ~w4715;
assign w4748 = ~w4746 & ~w4747;
assign w4749 = pi0743 & pi0947;
assign w4750 = pi0907 & ~pi0947;
assign w4751 = pi0735 & w4750;
assign w4752 = ~w4749 & ~w4751;
assign w4753 = w4715 & ~w4752;
assign w4754 = pi0146 & ~w4715;
assign w4755 = ~w4753 & ~w4754;
assign w4756 = ~pi0770 & pi0947;
assign w4757 = pi0726 & w4750;
assign w4758 = ~w4756 & ~w4757;
assign w4759 = w4715 & ~w4758;
assign w4760 = ~pi0147 & ~w4715;
assign w4761 = ~w4759 & ~w4760;
assign w4762 = pi0749 & pi0947;
assign w4763 = pi0706 & w4750;
assign w4764 = ~w4762 & ~w4763;
assign w4765 = w4715 & ~w4764;
assign w4766 = ~pi0148 & ~w4715;
assign w4767 = ~w4765 & ~w4766;
assign w4768 = ~pi0725 & w4750;
assign w4769 = ~pi0755 & pi0947;
assign w4770 = ~w4768 & ~w4769;
assign w4771 = w4715 & ~w4770;
assign w4772 = ~pi0149 & ~w4715;
assign w4773 = ~w4771 & ~w4772;
assign w4774 = ~pi0701 & w4750;
assign w4775 = ~pi0751 & pi0947;
assign w4776 = ~w4774 & ~w4775;
assign w4777 = w4715 & ~w4776;
assign w4778 = ~pi0150 & ~w4715;
assign w4779 = ~w4777 & ~w4778;
assign w4780 = ~pi0723 & w4750;
assign w4781 = ~pi0745 & pi0947;
assign w4782 = ~w4780 & ~w4781;
assign w4783 = w4715 & ~w4782;
assign w4784 = ~pi0151 & ~w4715;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = pi0759 & pi0947;
assign w4787 = pi0696 & w4750;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = w4715 & ~w4788;
assign w4790 = pi0152 & ~w4715;
assign w4791 = ~w4789 & ~w4790;
assign w4792 = pi0766 & pi0947;
assign w4793 = pi0700 & w4750;
assign w4794 = ~w4792 & ~w4793;
assign w4795 = w4715 & ~w4794;
assign w4796 = ~pi0153 & ~w4715;
assign w4797 = ~w4795 & ~w4796;
assign w4798 = ~pi0704 & w4750;
assign w4799 = ~pi0742 & pi0947;
assign w4800 = ~w4798 & ~w4799;
assign w4801 = w4715 & ~w4800;
assign w4802 = ~pi0154 & ~w4715;
assign w4803 = ~w4801 & ~w4802;
assign w4804 = ~pi0686 & w4750;
assign w4805 = ~pi0757 & pi0947;
assign w4806 = ~w4804 & ~w4805;
assign w4807 = w4715 & ~w4806;
assign w4808 = ~pi0155 & ~w4715;
assign w4809 = ~w4807 & ~w4808;
assign w4810 = ~pi0724 & w4750;
assign w4811 = ~pi0741 & pi0947;
assign w4812 = ~w4810 & ~w4811;
assign w4813 = w4715 & ~w4812;
assign w4814 = ~pi0156 & ~w4715;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = ~pi0688 & w4750;
assign w4817 = ~pi0760 & pi0947;
assign w4818 = ~w4816 & ~w4817;
assign w4819 = w4715 & ~w4818;
assign w4820 = ~pi0157 & ~w4715;
assign w4821 = ~w4819 & ~w4820;
assign w4822 = ~pi0702 & w4750;
assign w4823 = ~pi0753 & pi0947;
assign w4824 = ~w4822 & ~w4823;
assign w4825 = w4715 & ~w4824;
assign w4826 = ~pi0158 & ~w4715;
assign w4827 = ~w4825 & ~w4826;
assign w4828 = ~pi0709 & w4750;
assign w4829 = ~pi0754 & pi0947;
assign w4830 = ~w4828 & ~w4829;
assign w4831 = w4715 & ~w4830;
assign w4832 = ~pi0159 & ~w4715;
assign w4833 = ~w4831 & ~w4832;
assign w4834 = ~pi0734 & w4750;
assign w4835 = ~pi0756 & pi0947;
assign w4836 = ~w4834 & ~w4835;
assign w4837 = w4715 & ~w4836;
assign w4838 = ~pi0160 & ~w4715;
assign w4839 = ~w4837 & ~w4838;
assign w4840 = pi0758 & pi0947;
assign w4841 = pi0736 & w4750;
assign w4842 = ~w4840 & ~w4841;
assign w4843 = w4715 & ~w4842;
assign w4844 = pi0161 & ~w4715;
assign w4845 = ~w4843 & ~w4844;
assign w4846 = ~pi0738 & w4750;
assign w4847 = ~pi0761 & pi0947;
assign w4848 = ~w4846 & ~w4847;
assign w4849 = w4715 & ~w4848;
assign w4850 = ~pi0162 & ~w4715;
assign w4851 = ~w4849 & ~w4850;
assign w4852 = ~pi0737 & w4750;
assign w4853 = ~pi0777 & pi0947;
assign w4854 = ~w4852 & ~w4853;
assign w4855 = w4715 & ~w4854;
assign w4856 = ~pi0163 & ~w4715;
assign w4857 = ~w4855 & ~w4856;
assign w4858 = ~pi0752 & pi0947;
assign w4859 = pi0703 & w4750;
assign w4860 = ~w4858 & ~w4859;
assign w4861 = w4715 & ~w4860;
assign w4862 = ~pi0164 & ~w4715;
assign w4863 = ~w4861 & ~w4862;
assign w4864 = ~pi0774 & pi0947;
assign w4865 = pi0687 & w4750;
assign w4866 = ~w4864 & ~w4865;
assign w4867 = w4715 & ~w4866;
assign w4868 = ~pi0165 & ~w4715;
assign w4869 = ~w4867 & ~w4868;
assign w4870 = pi0772 & pi0947;
assign w4871 = pi0727 & w4750;
assign w4872 = ~w4870 & ~w4871;
assign w4873 = w4715 & ~w4872;
assign w4874 = pi0166 & ~w4715;
assign w4875 = ~w4873 & ~w4874;
assign w4876 = ~pi0768 & pi0947;
assign w4877 = pi0705 & w4750;
assign w4878 = ~w4876 & ~w4877;
assign w4879 = w4715 & ~w4878;
assign w4880 = ~pi0167 & ~w4715;
assign w4881 = ~w4879 & ~w4880;
assign w4882 = pi0763 & pi0947;
assign w4883 = pi0699 & w4750;
assign w4884 = ~w4882 & ~w4883;
assign w4885 = w4715 & ~w4884;
assign w4886 = ~pi0168 & ~w4715;
assign w4887 = ~w4885 & ~w4886;
assign w4888 = pi0746 & pi0947;
assign w4889 = pi0729 & w4750;
assign w4890 = ~w4888 & ~w4889;
assign w4891 = w4715 & ~w4890;
assign w4892 = ~pi0169 & ~w4715;
assign w4893 = ~w4891 & ~w4892;
assign w4894 = pi0748 & pi0947;
assign w4895 = pi0730 & w4750;
assign w4896 = ~w4894 & ~w4895;
assign w4897 = w4715 & ~w4896;
assign w4898 = ~pi0170 & ~w4715;
assign w4899 = ~w4897 & ~w4898;
assign w4900 = pi0764 & pi0947;
assign w4901 = pi0691 & w4750;
assign w4902 = ~w4900 & ~w4901;
assign w4903 = w4715 & ~w4902;
assign w4904 = ~pi0171 & ~w4715;
assign w4905 = ~w4903 & ~w4904;
assign w4906 = pi0739 & pi0947;
assign w4907 = pi0690 & w4750;
assign w4908 = ~w4906 & ~w4907;
assign w4909 = w4715 & ~w4908;
assign w4910 = ~pi0172 & ~w4715;
assign w4911 = ~w4909 & ~w4910;
assign w4912 = ~pi0723 & w4675;
assign w4913 = ~pi0745 & w4674;
assign w4914 = ~w4912 & ~w4913;
assign w4915 = w4715 & ~w4914;
assign w4916 = ~pi0173 & ~w4715;
assign w4917 = ~w4915 & ~w4916;
assign w4918 = pi0696 & w4675;
assign w4919 = pi0759 & w4674;
assign w4920 = ~w4918 & ~w4919;
assign w4921 = w4715 & ~w4920;
assign w4922 = pi0174 & ~w4715;
assign w4923 = ~w4921 & ~w4922;
assign w4924 = pi0700 & w4675;
assign w4925 = pi0766 & w4674;
assign w4926 = ~w4924 & ~w4925;
assign w4927 = w4715 & ~w4926;
assign w4928 = ~pi0175 & ~w4715;
assign w4929 = ~w4927 & ~w4928;
assign w4930 = ~pi0704 & w4675;
assign w4931 = ~pi0742 & w4674;
assign w4932 = ~w4930 & ~w4931;
assign w4933 = w4715 & ~w4932;
assign w4934 = ~pi0176 & ~w4715;
assign w4935 = ~w4933 & ~w4934;
assign w4936 = ~pi0686 & w4675;
assign w4937 = ~pi0757 & w4674;
assign w4938 = ~w4936 & ~w4937;
assign w4939 = w4715 & ~w4938;
assign w4940 = ~pi0177 & ~w4715;
assign w4941 = ~w4939 & ~w4940;
assign w4942 = ~pi0688 & w4675;
assign w4943 = ~pi0760 & w4674;
assign w4944 = ~w4942 & ~w4943;
assign w4945 = w4715 & ~w4944;
assign w4946 = ~pi0178 & ~w4715;
assign w4947 = ~w4945 & ~w4946;
assign w4948 = ~pi0724 & w4675;
assign w4949 = ~pi0741 & w4674;
assign w4950 = ~w4948 & ~w4949;
assign w4951 = w4715 & ~w4950;
assign w4952 = ~pi0179 & ~w4715;
assign w4953 = ~w4951 & ~w4952;
assign w4954 = ~pi0702 & w4675;
assign w4955 = ~pi0753 & w4674;
assign w4956 = ~w4954 & ~w4955;
assign w4957 = w4715 & ~w4956;
assign w4958 = ~pi0180 & ~w4715;
assign w4959 = ~w4957 & ~w4958;
assign w4960 = ~pi0709 & w4675;
assign w4961 = ~pi0754 & w4674;
assign w4962 = ~w4960 & ~w4961;
assign w4963 = w4715 & ~w4962;
assign w4964 = ~pi0181 & ~w4715;
assign w4965 = ~w4963 & ~w4964;
assign w4966 = ~pi0734 & w4675;
assign w4967 = ~pi0756 & w4674;
assign w4968 = ~w4966 & ~w4967;
assign w4969 = w4715 & ~w4968;
assign w4970 = ~pi0182 & ~w4715;
assign w4971 = ~w4969 & ~w4970;
assign w4972 = ~pi0725 & w4675;
assign w4973 = ~pi0755 & w4674;
assign w4974 = ~w4972 & ~w4973;
assign w4975 = w4715 & ~w4974;
assign w4976 = ~pi0183 & ~w4715;
assign w4977 = ~w4975 & ~w4976;
assign w4978 = ~pi0737 & w4675;
assign w4979 = ~pi0777 & w4674;
assign w4980 = ~w4978 & ~w4979;
assign w4981 = w4715 & ~w4980;
assign w4982 = ~pi0184 & ~w4715;
assign w4983 = ~w4981 & ~w4982;
assign w4984 = ~pi0701 & w4675;
assign w4985 = ~pi0751 & w4674;
assign w4986 = ~w4984 & ~w4985;
assign w4987 = w4715 & ~w4986;
assign w4988 = ~pi0185 & ~w4715;
assign w4989 = ~w4987 & ~w4988;
assign w4990 = pi0703 & w4675;
assign w4991 = ~pi0752 & w4674;
assign w4992 = ~w4990 & ~w4991;
assign w4993 = w4715 & ~w4992;
assign w4994 = ~pi0186 & ~w4715;
assign w4995 = ~w4993 & ~w4994;
assign w4996 = pi0726 & w4675;
assign w4997 = ~pi0770 & w4674;
assign w4998 = ~w4996 & ~w4997;
assign w4999 = w4715 & ~w4998;
assign w5000 = ~pi0187 & ~w4715;
assign w5001 = ~w4999 & ~w5000;
assign w5002 = pi0705 & w4675;
assign w5003 = ~pi0768 & w4674;
assign w5004 = ~w5002 & ~w5003;
assign w5005 = w4715 & ~w5004;
assign w5006 = ~pi0188 & ~w4715;
assign w5007 = ~w5005 & ~w5006;
assign w5008 = pi0727 & w4675;
assign w5009 = pi0772 & w4674;
assign w5010 = ~w5008 & ~w5009;
assign w5011 = w4715 & ~w5010;
assign w5012 = pi0189 & ~w4715;
assign w5013 = ~w5011 & ~w5012;
assign w5014 = pi0699 & w4675;
assign w5015 = pi0763 & w4674;
assign w5016 = ~w5014 & ~w5015;
assign w5017 = w4715 & ~w5016;
assign w5018 = ~pi0190 & ~w4715;
assign w5019 = ~w5017 & ~w5018;
assign w5020 = pi0729 & w4675;
assign w5021 = pi0746 & w4674;
assign w5022 = ~w5020 & ~w5021;
assign w5023 = w4715 & ~w5022;
assign w5024 = ~pi0191 & ~w4715;
assign w5025 = ~w5023 & ~w5024;
assign w5026 = pi0691 & w4675;
assign w5027 = pi0764 & w4674;
assign w5028 = ~w5026 & ~w5027;
assign w5029 = w4715 & ~w5028;
assign w5030 = ~pi0192 & ~w4715;
assign w5031 = ~w5029 & ~w5030;
assign w5032 = pi0690 & w4675;
assign w5033 = pi0739 & w4674;
assign w5034 = ~w5032 & ~w5033;
assign w5035 = w4715 & ~w5034;
assign w5036 = ~pi0193 & ~w4715;
assign w5037 = ~w5035 & ~w5036;
assign w5038 = pi0730 & w4675;
assign w5039 = pi0748 & w4674;
assign w5040 = ~w5038 & ~w5039;
assign w5041 = w4715 & ~w5040;
assign w5042 = ~pi0194 & ~w4715;
assign w5043 = ~w5041 & ~w5042;
assign w5044 = ~pi0196 & w4568;
assign w5045 = ~pi0138 & w5044;
assign w5046 = pi0195 & ~w5045;
assign w5047 = w4564 & w5046;
assign w5048 = w1658 & w5047;
assign w5049 = w2824 & ~w4557;
assign w5050 = w5048 & w5049;
assign w5051 = ~w3486 & ~w5047;
assign w5052 = ~w5050 & ~w5051;
assign w5053 = pi0171 & pi0299;
assign w5054 = pi0192 & ~pi0299;
assign w5055 = ~w5053 & ~w5054;
assign w5056 = ~w3485 & ~w5055;
assign w5057 = w378 & w5056;
assign w5058 = w2483 & w5057;
assign w5059 = w5052 & ~w5058;
assign w5060 = pi0194 & ~pi0299;
assign w5061 = pi0170 & pi0299;
assign w5062 = ~w5060 & ~w5061;
assign w5063 = w2483 & ~w5062;
assign w5064 = w3486 & w5063;
assign w5065 = w4557 & ~w5064;
assign w5066 = w1481 & ~w5065;
assign w5067 = ~pi0138 & pi0195;
assign w5068 = w5044 & w5067;
assign w5069 = ~pi0138 & w4568;
assign w5070 = pi0196 & ~w5069;
assign w5071 = ~w5068 & ~w5070;
assign w5072 = w4564 & ~w5071;
assign w5073 = ~w3486 & ~w5072;
assign w5074 = ~w5066 & ~w5073;
assign w5075 = ~pi0698 & w4750;
assign w5076 = ~pi0767 & pi0947;
assign w5077 = ~w5075 & ~w5076;
assign w5078 = w4715 & ~w5077;
assign w5079 = ~pi0197 & ~w4715;
assign w5080 = ~w5078 & ~w5079;
assign w5081 = pi0634 & w4675;
assign w5082 = pi0633 & w4674;
assign w5083 = ~w5081 & ~w5082;
assign w5084 = ~w4691 & w4697;
assign w5085 = ~w1649 & w5084;
assign w5086 = ~w4708 & ~w4711;
assign w5087 = w1475 & ~w5086;
assign w5088 = ~w5085 & w5087;
assign w5089 = ~w5083 & w5088;
assign w5090 = pi0198 & ~w5088;
assign w5091 = ~w5089 & ~w5090;
assign w5092 = pi0637 & w4675;
assign w5093 = pi0617 & w4674;
assign w5094 = ~w5092 & ~w5093;
assign w5095 = w5088 & ~w5094;
assign w5096 = pi0199 & ~w5088;
assign w5097 = ~w5095 & ~w5096;
assign w5098 = pi0643 & w4675;
assign w5099 = pi0606 & w4674;
assign w5100 = ~w5098 & ~w5099;
assign w5101 = w5088 & ~w5100;
assign w5102 = pi0200 & ~w5088;
assign w5103 = ~w5101 & ~w5102;
assign w5104 = pi0233 & pi0237;
assign w5105 = ~w4537 & ~w4539;
assign w5106 = ~pi0070 & ~w5105;
assign w5107 = pi0032 & w5106;
assign w5108 = ~pi0841 & w5107;
assign w5109 = ~pi0032 & pi0070;
assign w5110 = ~w5108 & ~w5109;
assign w5111 = w5104 & ~w5110;
assign w5112 = ~w443 & w3858;
assign w5113 = ~pi0055 & ~pi0059;
assign w5114 = pi0054 & w5113;
assign w5115 = pi0055 & ~pi0059;
assign w5116 = ~pi0055 & pi0059;
assign w5117 = ~w5115 & ~w5116;
assign w5118 = ~pi0054 & ~w5117;
assign w5119 = ~w5114 & ~w5118;
assign w5120 = w2932 & ~w5119;
assign w5121 = w1300 & w5120;
assign w5122 = w113 & w5121;
assign w5123 = ~w5112 & ~w5122;
assign w5124 = ~pi0332 & w5123;
assign w5125 = ~w5111 & w5124;
assign w5126 = ~pi0587 & w526;
assign w5127 = ~pi0947 & ~w526;
assign w5128 = ~w5126 & ~w5127;
assign w5129 = ~pi0468 & ~w5128;
assign w5130 = pi0468 & ~w1249;
assign w5131 = ~w5129 & ~w5130;
assign w5132 = ~pi0332 & ~w5131;
assign w5133 = ~w5125 & ~w5132;
assign w5134 = ~pi0201 & ~w5133;
assign w5135 = pi0210 & ~w526;
assign w5136 = pi0198 & w526;
assign w5137 = ~w5135 & ~w5136;
assign w5138 = pi0947 & ~w526;
assign w5139 = pi0587 & w526;
assign w5140 = ~w5138 & ~w5139;
assign w5141 = w1241 & ~w5140;
assign w5142 = ~w1551 & ~w5141;
assign w5143 = ~w5137 & ~w5142;
assign w5144 = pi0096 & w5143;
assign w5145 = w5104 & w5144;
assign w5146 = ~w5134 & ~w5145;
assign w5147 = ~pi0233 & pi0237;
assign w5148 = ~w5110 & w5147;
assign w5149 = w5124 & ~w5148;
assign w5150 = ~w5132 & ~w5149;
assign w5151 = ~pi0202 & ~w5150;
assign w5152 = w5144 & w5147;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = ~pi0233 & ~pi0237;
assign w5155 = ~w5110 & w5154;
assign w5156 = w5124 & ~w5155;
assign w5157 = ~w5132 & ~w5156;
assign w5158 = ~pi0203 & ~w5157;
assign w5159 = w5144 & w5154;
assign w5160 = ~w5158 & ~w5159;
assign w5161 = ~pi0602 & w526;
assign w5162 = ~pi0907 & ~w526;
assign w5163 = ~w5161 & ~w5162;
assign w5164 = ~pi0468 & ~w5163;
assign w5165 = pi0468 & ~w1253;
assign w5166 = ~w5164 & ~w5165;
assign w5167 = ~pi0332 & ~w5166;
assign w5168 = ~w5125 & ~w5167;
assign w5169 = ~pi0204 & ~w5168;
assign w5170 = pi0907 & ~w526;
assign w5171 = pi0602 & w526;
assign w5172 = ~w5170 & ~w5171;
assign w5173 = w1241 & ~w5172;
assign w5174 = ~w1497 & ~w5173;
assign w5175 = ~w5137 & ~w5174;
assign w5176 = pi0096 & w5175;
assign w5177 = w5104 & w5176;
assign w5178 = ~w5169 & ~w5177;
assign w5179 = ~w5149 & ~w5167;
assign w5180 = ~pi0205 & ~w5179;
assign w5181 = w5147 & w5176;
assign w5182 = ~w5180 & ~w5181;
assign w5183 = pi0233 & ~pi0237;
assign w5184 = ~w5110 & w5183;
assign w5185 = w5124 & ~w5184;
assign w5186 = ~w5167 & ~w5185;
assign w5187 = ~pi0206 & ~w5186;
assign w5188 = w5176 & w5183;
assign w5189 = ~w5187 & ~w5188;
assign w5190 = pi0710 & w4675;
assign w5191 = pi0623 & w4674;
assign w5192 = ~w5190 & ~w5191;
assign w5193 = w5088 & ~w5192;
assign w5194 = ~pi0207 & ~w5088;
assign w5195 = ~w5193 & ~w5194;
assign w5196 = pi0638 & w4675;
assign w5197 = pi0607 & w4674;
assign w5198 = ~w5196 & ~w5197;
assign w5199 = w5088 & ~w5198;
assign w5200 = ~pi0208 & ~w5088;
assign w5201 = ~w5199 & ~w5200;
assign w5202 = pi0639 & w4675;
assign w5203 = pi0622 & w4674;
assign w5204 = ~w5202 & ~w5203;
assign w5205 = w5088 & ~w5204;
assign w5206 = ~pi0209 & ~w5088;
assign w5207 = ~w5205 & ~w5206;
assign w5208 = pi0634 & w4750;
assign w5209 = pi0633 & pi0947;
assign w5210 = ~w5208 & ~w5209;
assign w5211 = w5088 & ~w5210;
assign w5212 = pi0210 & ~w5088;
assign w5213 = ~w5211 & ~w5212;
assign w5214 = pi0643 & w4750;
assign w5215 = pi0606 & pi0947;
assign w5216 = ~w5214 & ~w5215;
assign w5217 = w5088 & ~w5216;
assign w5218 = pi0211 & ~w5088;
assign w5219 = ~w5217 & ~w5218;
assign w5220 = pi0638 & w4750;
assign w5221 = pi0607 & pi0947;
assign w5222 = ~w5220 & ~w5221;
assign w5223 = w5088 & ~w5222;
assign w5224 = ~pi0212 & ~w5088;
assign w5225 = ~w5223 & ~w5224;
assign w5226 = pi0639 & w4750;
assign w5227 = pi0622 & pi0947;
assign w5228 = ~w5226 & ~w5227;
assign w5229 = w5088 & ~w5228;
assign w5230 = ~pi0213 & ~w5088;
assign w5231 = ~w5229 & ~w5230;
assign w5232 = pi0710 & w4750;
assign w5233 = pi0623 & pi0947;
assign w5234 = ~w5232 & ~w5233;
assign w5235 = w5088 & ~w5234;
assign w5236 = ~pi0214 & ~w5088;
assign w5237 = ~w5235 & ~w5236;
assign w5238 = pi0681 & w4750;
assign w5239 = pi0642 & pi0947;
assign w5240 = ~w5238 & ~w5239;
assign w5241 = w5088 & ~w5240;
assign w5242 = pi0215 & ~w5088;
assign w5243 = ~w5241 & ~w5242;
assign w5244 = pi0662 & w4750;
assign w5245 = pi0614 & pi0947;
assign w5246 = ~w5244 & ~w5245;
assign w5247 = w5088 & ~w5246;
assign w5248 = pi0216 & ~w5088;
assign w5249 = ~w5247 & ~w5248;
assign w5250 = ~pi0695 & w4675;
assign w5251 = pi0612 & w4674;
assign w5252 = ~w5250 & ~w5251;
assign w5253 = w5088 & ~w5252;
assign w5254 = ~pi0217 & ~w5088;
assign w5255 = ~w5253 & ~w5254;
assign w5256 = ~w5156 & ~w5167;
assign w5257 = ~pi0218 & ~w5256;
assign w5258 = w5154 & w5176;
assign w5259 = ~w5257 & ~w5258;
assign w5260 = pi0637 & w4750;
assign w5261 = pi0617 & pi0947;
assign w5262 = ~w5260 & ~w5261;
assign w5263 = w5088 & ~w5262;
assign w5264 = pi0219 & ~w5088;
assign w5265 = ~w5263 & ~w5264;
assign w5266 = ~w5132 & ~w5185;
assign w5267 = ~pi0220 & ~w5266;
assign w5268 = w5144 & w5183;
assign w5269 = ~w5267 & ~w5268;
assign w5270 = pi0661 & w4750;
assign w5271 = pi0616 & pi0947;
assign w5272 = ~w5270 & ~w5271;
assign w5273 = w5088 & ~w5272;
assign w5274 = pi0221 & ~w5088;
assign w5275 = ~w5273 & ~w5274;
assign w5276 = pi0661 & w4675;
assign w5277 = pi0616 & w4674;
assign w5278 = ~w5276 & ~w5277;
assign w5279 = w5088 & ~w5278;
assign w5280 = pi0222 & ~w5088;
assign w5281 = ~w5279 & ~w5280;
assign w5282 = pi0681 & w4675;
assign w5283 = pi0642 & w4674;
assign w5284 = ~w5282 & ~w5283;
assign w5285 = w5088 & ~w5284;
assign w5286 = pi0223 & ~w5088;
assign w5287 = ~w5285 & ~w5286;
assign w5288 = pi0662 & w4675;
assign w5289 = pi0614 & w4674;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = w5088 & ~w5290;
assign w5292 = pi0224 & ~w5088;
assign w5293 = ~w5291 & ~w5292;
assign w5294 = w413 & ~w448;
assign w5295 = ~w147 & w5294;
assign w5296 = ~pi0055 & ~w5295;
assign w5297 = ~pi0137 & w5296;
assign w5298 = ~w3393 & ~w5297;
assign w5299 = ~w490 & w501;
assign w5300 = ~w441 & ~w461;
assign w5301 = ~w5299 & w5300;
assign w5302 = ~w420 & ~w5301;
assign w5303 = w593 & ~w5302;
assign w5304 = ~w5298 & ~w5303;
assign w5305 = pi0228 & pi0231;
assign w5306 = ~pi0032 & w443;
assign w5307 = ~pi0070 & ~pi0095;
assign w5308 = w5306 & w5307;
assign w5309 = ~w1364 & ~w5308;
assign w5310 = ~w2553 & ~w5309;
assign w5311 = w593 & w5310;
assign w5312 = ~w205 & w5311;
assign w5313 = ~pi0054 & w1619;
assign w5314 = ~w1360 & ~w5313;
assign w5315 = ~w1355 & w5314;
assign w5316 = ~w1664 & w5315;
assign w5317 = ~pi0479 & w1360;
assign w5318 = ~w5316 & ~w5317;
assign w5319 = ~w5312 & ~w5318;
assign w5320 = ~pi0228 & ~w5319;
assign w5321 = ~w5305 & ~w5320;
assign w5322 = ~pi0036 & ~pi0104;
assign w5323 = ~pi0088 & w5322;
assign w5324 = ~w2950 & ~w5323;
assign w5325 = pi0036 & pi1093;
assign w5326 = ~pi0047 & ~w5325;
assign w5327 = ~pi0091 & w5326;
assign w5328 = ~pi0072 & w5327;
assign w5329 = ~w5324 & w5328;
assign w5330 = pi0036 & w454;
assign w5331 = ~w5329 & ~w5330;
assign w5332 = w2554 & w5331;
assign w5333 = ~w3477 & ~w5332;
assign w5334 = ~pi0039 & w3502;
assign w5335 = ~w3771 & ~w5334;
assign w5336 = ~pi1093 & ~w453;
assign w5337 = ~w450 & ~w5336;
assign w5338 = ~w5335 & w5337;
assign w5339 = ~pi0039 & ~w3771;
assign w5340 = pi0228 & w5339;
assign w5341 = ~w5338 & ~w5340;
assign w5342 = ~pi0047 & w2568;
assign w5343 = w112 & ~w2823;
assign w5344 = w5342 & w5343;
assign w5345 = ~w2553 & ~w4689;
assign w5346 = ~w205 & w5345;
assign w5347 = w4697 & ~w5346;
assign w5348 = w4711 & ~w5347;
assign w5349 = ~w4708 & ~w5348;
assign w5350 = ~w5344 & ~w5349;
assign w5351 = pi0065 & ~pi0102;
assign w5352 = ~pi0065 & pi0102;
assign w5353 = ~w5351 & ~w5352;
assign w5354 = w67 & ~w5353;
assign w5355 = ~pi0064 & w532;
assign w5356 = w5354 & w5355;
assign w5357 = ~w2990 & ~w5356;
assign w5358 = w1379 & w5357;
assign w5359 = ~w3393 & ~w3407;
assign w5360 = ~w5358 & ~w5359;
assign w5361 = ~pi0212 & ~pi0214;
assign w5362 = pi0219 & ~w5361;
assign w5363 = pi1142 & w5362;
assign w5364 = ~pi0211 & w5363;
assign w5365 = ~pi0211 & pi1143;
assign w5366 = pi0211 & pi1142;
assign w5367 = ~w5365 & ~w5366;
assign w5368 = pi0212 & ~w5367;
assign w5369 = pi0214 & w5368;
assign w5370 = ~pi0211 & pi1144;
assign w5371 = pi0211 & pi1143;
assign w5372 = ~w5370 & ~w5371;
assign w5373 = ~pi0212 & pi0214;
assign w5374 = pi0212 & ~pi0214;
assign w5375 = ~w5373 & ~w5374;
assign w5376 = ~w5372 & ~w5375;
assign w5377 = ~w5369 & ~w5376;
assign w5378 = ~pi0219 & ~w5377;
assign w5379 = ~w5364 & ~w5378;
assign w5380 = pi0213 & ~w5379;
assign w5381 = pi0211 & ~pi0219;
assign w5382 = pi1156 & w5381;
assign w5383 = pi0219 & pi1155;
assign w5384 = ~pi0219 & pi1157;
assign w5385 = ~w5383 & ~w5384;
assign w5386 = ~pi0211 & ~w5385;
assign w5387 = ~w5382 & ~w5386;
assign w5388 = pi0214 & ~w5387;
assign w5389 = ~pi0212 & w5388;
assign w5390 = ~pi0214 & pi1154;
assign w5391 = pi0214 & pi1153;
assign w5392 = ~w5390 & ~w5391;
assign w5393 = pi0219 & ~w5392;
assign w5394 = ~pi0211 & w5393;
assign w5395 = ~pi1154 & w3181;
assign w5396 = ~pi0211 & ~pi0214;
assign w5397 = ~pi1156 & w5396;
assign w5398 = ~w5395 & ~w5397;
assign w5399 = pi0211 & ~pi0214;
assign w5400 = ~w3210 & ~w5399;
assign w5401 = ~pi1155 & ~w5400;
assign w5402 = w5398 & ~w5401;
assign w5403 = ~pi0219 & w5402;
assign w5404 = ~w5394 & ~w5403;
assign w5405 = pi0212 & ~w5404;
assign w5406 = ~w5389 & ~w5405;
assign w5407 = ~pi0213 & ~w5406;
assign w5408 = ~w5380 & ~w5407;
assign w5409 = ~w526 & ~w5408;
assign w5410 = pi0230 & ~w5409;
assign w5411 = ~pi0207 & ~pi0208;
assign w5412 = pi0199 & ~w5411;
assign w5413 = pi1142 & w5412;
assign w5414 = ~pi0200 & w5413;
assign w5415 = ~pi0200 & pi1143;
assign w5416 = pi0200 & pi1142;
assign w5417 = ~w5415 & ~w5416;
assign w5418 = pi0207 & ~w5417;
assign w5419 = pi0208 & w5418;
assign w5420 = ~pi0200 & pi1144;
assign w5421 = pi0200 & pi1143;
assign w5422 = ~w5420 & ~w5421;
assign w5423 = pi0207 & ~pi0208;
assign w5424 = ~pi0207 & pi0208;
assign w5425 = ~w5423 & ~w5424;
assign w5426 = ~w5422 & ~w5425;
assign w5427 = ~w5419 & ~w5426;
assign w5428 = ~pi0199 & ~w5427;
assign w5429 = ~w5414 & ~w5428;
assign w5430 = pi0209 & ~w5429;
assign w5431 = ~pi0199 & pi0200;
assign w5432 = pi1155 & w5431;
assign w5433 = pi0199 & pi1154;
assign w5434 = ~pi0199 & pi1156;
assign w5435 = ~w5433 & ~w5434;
assign w5436 = ~pi0200 & ~w5435;
assign w5437 = ~w5432 & ~w5436;
assign w5438 = w5424 & ~w5437;
assign w5439 = pi1156 & w5431;
assign w5440 = pi0199 & pi1155;
assign w5441 = ~pi0199 & pi1157;
assign w5442 = ~w5440 & ~w5441;
assign w5443 = ~pi0200 & ~w5442;
assign w5444 = ~w5439 & ~w5443;
assign w5445 = ~pi0208 & ~w5444;
assign w5446 = pi1154 & w5431;
assign w5447 = pi0199 & pi1153;
assign w5448 = ~pi0199 & pi1155;
assign w5449 = ~w5447 & ~w5448;
assign w5450 = ~pi0200 & ~w5449;
assign w5451 = ~w5446 & ~w5450;
assign w5452 = pi0208 & ~w5451;
assign w5453 = ~w5445 & ~w5452;
assign w5454 = pi0207 & ~w5453;
assign w5455 = ~w5438 & ~w5454;
assign w5456 = ~pi0209 & ~w5455;
assign w5457 = ~w5430 & ~w5456;
assign w5458 = w526 & ~w5457;
assign w5459 = w5410 & ~w5458;
assign w5460 = ~pi0230 & pi0233;
assign w5461 = ~w5459 & ~w5460;
assign w5462 = ~pi0230 & pi0234;
assign w5463 = ~pi0208 & w526;
assign w5464 = ~pi0207 & w5463;
assign w5465 = ~pi0214 & ~w526;
assign w5466 = ~pi0212 & w5465;
assign w5467 = ~w5464 & ~w5466;
assign w5468 = pi1154 & w5467;
assign w5469 = w3185 & w3310;
assign w5470 = w5468 & w5469;
assign w5471 = pi0213 & ~w526;
assign w5472 = ~pi0211 & pi0212;
assign w5473 = pi0214 & pi1155;
assign w5474 = w5472 & w5473;
assign w5475 = pi0211 & pi1155;
assign w5476 = ~pi0211 & pi1156;
assign w5477 = ~w5475 & ~w5476;
assign w5478 = ~w5375 & ~w5477;
assign w5479 = ~w5474 & ~w5478;
assign w5480 = ~pi0219 & ~w5479;
assign w5481 = w5471 & ~w5480;
assign w5482 = ~pi0200 & pi1156;
assign w5483 = pi0200 & pi1155;
assign w5484 = ~w5482 & ~w5483;
assign w5485 = ~w5425 & ~w5484;
assign w5486 = ~pi0200 & pi0207;
assign w5487 = pi0208 & pi1155;
assign w5488 = w5486 & w5487;
assign w5489 = ~w5485 & ~w5488;
assign w5490 = ~pi0199 & ~w5489;
assign w5491 = w526 & ~w5490;
assign w5492 = pi0209 & w5491;
assign w5493 = ~w5481 & ~w5492;
assign w5494 = ~w5470 & ~w5493;
assign w5495 = pi0209 & w526;
assign w5496 = ~w5471 & ~w5495;
assign w5497 = pi1152 & w5469;
assign w5498 = pi1154 & ~w3310;
assign w5499 = pi1153 & w3310;
assign w5500 = ~w5498 & ~w5499;
assign w5501 = ~w3185 & ~w5500;
assign w5502 = ~w5497 & ~w5501;
assign w5503 = w5467 & ~w5502;
assign w5504 = w5496 & ~w5503;
assign w5505 = ~w5494 & ~w5504;
assign w5506 = pi0230 & w5505;
assign w5507 = ~w5462 & ~w5506;
assign w5508 = ~pi0213 & pi1154;
assign w5509 = pi0213 & pi1156;
assign w5510 = ~w5508 & ~w5509;
assign w5511 = ~pi0211 & ~w5510;
assign w5512 = ~pi0213 & pi1153;
assign w5513 = pi0213 & pi1155;
assign w5514 = ~w5512 & ~w5513;
assign w5515 = pi0211 & ~w5514;
assign w5516 = ~w5511 & ~w5515;
assign w5517 = ~pi0219 & ~w5516;
assign w5518 = w3213 & w5517;
assign w5519 = pi0211 & ~w5510;
assign w5520 = ~pi0219 & w5519;
assign w5521 = pi0213 & ~pi0219;
assign w5522 = pi1157 & w5521;
assign w5523 = ~pi0213 & pi0219;
assign w5524 = pi1153 & w5523;
assign w5525 = ~w5522 & ~w5524;
assign w5526 = pi0213 & pi0219;
assign w5527 = ~pi0213 & ~pi0219;
assign w5528 = ~w5526 & ~w5527;
assign w5529 = pi1155 & ~w5528;
assign w5530 = w5525 & ~w5529;
assign w5531 = ~pi0211 & ~w5530;
assign w5532 = ~w5520 & ~w5531;
assign w5533 = ~w5375 & ~w5532;
assign w5534 = ~w5518 & ~w5533;
assign w5535 = ~w526 & ~w5534;
assign w5536 = ~pi0209 & pi1154;
assign w5537 = pi0209 & pi1156;
assign w5538 = ~w5536 & ~w5537;
assign w5539 = ~pi0200 & ~w5538;
assign w5540 = ~pi0209 & pi1153;
assign w5541 = pi0209 & pi1155;
assign w5542 = ~w5540 & ~w5541;
assign w5543 = pi0200 & ~w5542;
assign w5544 = ~w5539 & ~w5543;
assign w5545 = ~pi0199 & ~w5544;
assign w5546 = w3177 & w5545;
assign w5547 = pi0209 & w5444;
assign w5548 = ~pi0209 & w5451;
assign w5549 = ~w5547 & ~w5548;
assign w5550 = ~w5425 & w5549;
assign w5551 = ~w5546 & ~w5550;
assign w5552 = w526 & ~w5551;
assign w5553 = ~w5535 & ~w5552;
assign w5554 = pi0230 & ~w5553;
assign w5555 = ~pi0230 & pi0235;
assign w5556 = ~w5554 & ~w5555;
assign w5557 = ~pi0230 & ~pi0237;
assign w5558 = pi0208 & ~w5437;
assign w5559 = pi1157 & w5431;
assign w5560 = pi0199 & pi1156;
assign w5561 = ~pi0199 & pi1158;
assign w5562 = ~w5560 & ~w5561;
assign w5563 = ~pi0200 & ~w5562;
assign w5564 = ~w5559 & ~w5563;
assign w5565 = ~pi0208 & ~w5564;
assign w5566 = ~w5558 & ~w5565;
assign w5567 = pi0207 & ~w5566;
assign w5568 = w5424 & ~w5444;
assign w5569 = ~w5567 & ~w5568;
assign w5570 = ~pi0209 & w5569;
assign w5571 = pi1143 & w5412;
assign w5572 = ~pi0200 & w5571;
assign w5573 = pi0207 & ~w5422;
assign w5574 = pi0208 & w5573;
assign w5575 = ~pi0200 & pi1145;
assign w5576 = pi0200 & pi1144;
assign w5577 = ~w5575 & ~w5576;
assign w5578 = ~w5425 & ~w5577;
assign w5579 = ~w5574 & ~w5578;
assign w5580 = ~pi0199 & ~w5579;
assign w5581 = ~w5572 & ~w5580;
assign w5582 = pi0209 & w5581;
assign w5583 = ~w5570 & ~w5582;
assign w5584 = w526 & ~w5583;
assign w5585 = ~pi0211 & pi1158;
assign w5586 = pi0211 & pi1157;
assign w5587 = ~w5585 & ~w5586;
assign w5588 = ~pi0219 & ~w5587;
assign w5589 = ~pi0211 & pi0219;
assign w5590 = pi1156 & w5589;
assign w5591 = ~w5588 & ~w5590;
assign w5592 = w5373 & ~w5591;
assign w5593 = ~pi0214 & pi1155;
assign w5594 = pi0214 & pi1154;
assign w5595 = ~w5593 & ~w5594;
assign w5596 = pi0219 & ~w5595;
assign w5597 = ~pi0211 & w5596;
assign w5598 = pi1155 & w3181;
assign w5599 = pi1157 & w5396;
assign w5600 = ~w5598 & ~w5599;
assign w5601 = pi1156 & ~w5400;
assign w5602 = w5600 & ~w5601;
assign w5603 = ~pi0219 & ~w5602;
assign w5604 = ~w5597 & ~w5603;
assign w5605 = pi0212 & ~w5604;
assign w5606 = ~w5592 & ~w5605;
assign w5607 = ~pi0213 & ~w5606;
assign w5608 = pi1143 & w5362;
assign w5609 = ~pi0211 & w5608;
assign w5610 = pi0212 & ~w5372;
assign w5611 = pi0214 & w5610;
assign w5612 = ~pi0211 & pi1145;
assign w5613 = pi0211 & pi1144;
assign w5614 = ~w5612 & ~w5613;
assign w5615 = ~w5375 & ~w5614;
assign w5616 = ~w5611 & ~w5615;
assign w5617 = ~pi0219 & ~w5616;
assign w5618 = ~w5609 & ~w5617;
assign w5619 = pi0213 & ~w5618;
assign w5620 = ~w5607 & ~w5619;
assign w5621 = ~w526 & w5620;
assign w5622 = ~w5584 & ~w5621;
assign w5623 = pi0230 & w5622;
assign w5624 = ~w5557 & ~w5623;
assign w5625 = pi1151 & w5469;
assign w5626 = pi1153 & ~w3310;
assign w5627 = pi1152 & w3310;
assign w5628 = ~w5626 & ~w5627;
assign w5629 = ~w3185 & ~w5628;
assign w5630 = ~w5625 & ~w5629;
assign w5631 = w5467 & ~w5630;
assign w5632 = w5496 & ~w5631;
assign w5633 = pi0230 & ~w5632;
assign w5634 = pi0214 & w5589;
assign w5635 = pi0214 & w5381;
assign w5636 = ~w5589 & ~w5635;
assign w5637 = pi0212 & ~w5636;
assign w5638 = ~w5634 & ~w5637;
assign w5639 = pi1153 & ~w5638;
assign w5640 = ~pi0211 & pi1155;
assign w5641 = pi0211 & pi1154;
assign w5642 = ~w5640 & ~w5641;
assign w5643 = ~w5375 & ~w5642;
assign w5644 = w5472 & w5594;
assign w5645 = ~w5643 & ~w5644;
assign w5646 = ~pi0219 & ~w5645;
assign w5647 = ~w5639 & ~w5646;
assign w5648 = w5471 & w5647;
assign w5649 = pi0199 & ~pi0200;
assign w5650 = pi1153 & w5649;
assign w5651 = ~pi0200 & ~w3177;
assign w5652 = pi1155 & w5651;
assign w5653 = ~w3205 & ~w3207;
assign w5654 = pi1154 & ~w5653;
assign w5655 = ~w5652 & ~w5654;
assign w5656 = ~pi0199 & ~w5655;
assign w5657 = ~w5650 & ~w5656;
assign w5658 = pi0208 & ~w5657;
assign w5659 = ~pi0207 & ~w5658;
assign w5660 = pi1153 & w5431;
assign w5661 = pi0208 & w5660;
assign w5662 = w5657 & ~w5661;
assign w5663 = ~w5659 & ~w5662;
assign w5664 = pi0209 & ~w5663;
assign w5665 = w526 & w5664;
assign w5666 = ~w5648 & ~w5665;
assign w5667 = w5633 & w5666;
assign w5668 = ~pi0230 & pi0238;
assign w5669 = ~w5667 & ~w5668;
assign w5670 = pi0209 & ~w5564;
assign w5671 = ~pi0209 & ~w5437;
assign w5672 = ~w5670 & ~w5671;
assign w5673 = ~pi0208 & ~w5672;
assign w5674 = pi0207 & w5673;
assign w5675 = w526 & w5674;
assign w5676 = pi0213 & ~w5591;
assign w5677 = ~pi0213 & ~w5604;
assign w5678 = ~w5676 & ~w5677;
assign w5679 = pi0214 & ~w5678;
assign w5680 = ~pi0212 & w5679;
assign w5681 = ~w526 & w5680;
assign w5682 = ~w5675 & ~w5681;
assign w5683 = pi0230 & ~w5682;
assign w5684 = ~pi0230 & pi0239;
assign w5685 = ~w5683 & ~w5684;
assign w5686 = pi1147 & w5469;
assign w5687 = pi1149 & ~w3310;
assign w5688 = pi1148 & w3310;
assign w5689 = ~w5687 & ~w5688;
assign w5690 = ~w3185 & ~w5689;
assign w5691 = ~w5686 & ~w5690;
assign w5692 = w5467 & ~w5691;
assign w5693 = ~w5496 & w5692;
assign w5694 = pi1145 & w5469;
assign w5695 = pi1147 & ~w3310;
assign w5696 = pi1146 & w3310;
assign w5697 = ~w5695 & ~w5696;
assign w5698 = ~w3185 & ~w5697;
assign w5699 = ~w5694 & ~w5698;
assign w5700 = w5467 & ~w5699;
assign w5701 = w5496 & w5700;
assign w5702 = ~w5693 & ~w5701;
assign w5703 = pi0230 & ~w5702;
assign w5704 = ~pi0230 & pi0240;
assign w5705 = ~w5703 & ~w5704;
assign w5706 = pi1149 & w5469;
assign w5707 = pi1151 & ~w3310;
assign w5708 = pi1150 & w3310;
assign w5709 = ~w5707 & ~w5708;
assign w5710 = ~w3185 & ~w5709;
assign w5711 = ~w5706 & ~w5710;
assign w5712 = w5467 & ~w5711;
assign w5713 = w5496 & w5712;
assign w5714 = ~w5496 & w5631;
assign w5715 = ~w5713 & ~w5714;
assign w5716 = pi0230 & ~w5715;
assign w5717 = ~pi0230 & pi0241;
assign w5718 = ~w5716 & ~w5717;
assign w5719 = ~pi0230 & pi0242;
assign w5720 = ~pi0213 & ~w526;
assign w5721 = w5379 & w5720;
assign w5722 = ~pi0209 & w526;
assign w5723 = w5429 & w5722;
assign w5724 = ~w5721 & ~w5723;
assign w5725 = pi1144 & w5469;
assign w5726 = pi1146 & ~w3310;
assign w5727 = pi1145 & w3310;
assign w5728 = ~w5726 & ~w5727;
assign w5729 = ~w3185 & ~w5728;
assign w5730 = ~w5725 & ~w5729;
assign w5731 = w5467 & ~w5730;
assign w5732 = ~w5496 & ~w5731;
assign w5733 = w5724 & ~w5732;
assign w5734 = pi0230 & w5733;
assign w5735 = ~w5719 & ~w5734;
assign w5736 = pi0199 & w525;
assign w5737 = w180 & w5736;
assign w5738 = pi0219 & ~w525;
assign w5739 = (pi0219 & ~w180) | (pi0219 & w5738) | (~w180 & w5738);
assign w5740 = ~w5737 & ~w5739;
assign w5741 = ~pi0083 & ~pi0085;
assign w5742 = pi0314 & ~w5741;
assign w5743 = pi0271 & w5742;
assign w5744 = ~pi0081 & ~pi0083;
assign w5745 = ~pi0085 & w5744;
assign w5746 = pi0314 & ~w5745;
assign w5747 = pi0271 & w5746;
assign w5748 = (w5740 & w5743) | (w5740 & w5747) | (w5743 & w5747);
assign w5749 = pi0273 & pi0276;
assign w5750 = pi0283 & w5749;
assign w5751 = pi0802 & w5750;
assign w5752 = pi0253 & w5751;
assign w5753 = pi0268 & w5752;
assign w5754 = w5748 & w5753;
assign w5755 = pi0272 & pi0275;
assign w5756 = pi0254 & ~pi0263;
assign w5757 = pi0267 & w5756;
assign w5758 = w5755 & w5757;
assign w5759 = ~pi0243 & ~w5758;
assign w5760 = (~pi0243 & ~w5754) | (~pi0243 & w5759) | (~w5754 & w5759);
assign w5761 = pi0243 & pi0267;
assign w5762 = w5756 & w5761;
assign w5763 = w5755 & w5762;
assign w5764 = w5754 & w5763;
assign w5765 = ~w5760 & ~w5764;
assign w5766 = ~pi0230 & ~pi1091;
assign w5767 = ~w5765 & w5766;
assign w5768 = ~pi0200 & w525;
assign w5769 = w180 & w5768;
assign w5770 = ~pi0199 & w5769;
assign w5771 = ~pi0219 & ~w525;
assign w5772 = (~pi0219 & ~w180) | (~pi0219 & w5771) | (~w180 & w5771);
assign w5773 = ~pi0211 & w5772;
assign w5774 = ~w5770 & ~w5773;
assign w5775 = pi1155 & ~w5774;
assign w5776 = pi0199 & w5769;
assign w5777 = ~pi0211 & w5739;
assign w5778 = ~w5776 & ~w5777;
assign w5779 = pi1157 & ~w5778;
assign w5780 = ~w5775 & ~w5779;
assign w5781 = pi0211 & w5772;
assign w5782 = pi0200 & w525;
assign w5783 = w180 & w5782;
assign w5784 = ~pi0199 & w5783;
assign w5785 = ~w5781 & ~w5784;
assign w5786 = pi1156 & ~w5785;
assign w5787 = ~w5766 & w5786;
assign w5788 = (~w5766 & ~w5780) | (~w5766 & w5787) | (~w5780 & w5787);
assign w5789 = ~w5767 & ~w5788;
assign w5790 = ~pi0230 & pi0244;
assign w5791 = w5618 & w5720;
assign w5792 = w5581 & w5722;
assign w5793 = ~w5791 & ~w5792;
assign w5794 = ~w5496 & ~w5700;
assign w5795 = w5793 & ~w5794;
assign w5796 = pi0230 & w5795;
assign w5797 = ~w5790 & ~w5796;
assign w5798 = pi1146 & w5469;
assign w5799 = pi1148 & ~w3310;
assign w5800 = pi1147 & w3310;
assign w5801 = ~w5799 & ~w5800;
assign w5802 = ~w3185 & ~w5801;
assign w5803 = ~w5798 & ~w5802;
assign w5804 = w5467 & ~w5803;
assign w5805 = ~w5496 & w5804;
assign w5806 = w5496 & w5731;
assign w5807 = ~w5805 & ~w5806;
assign w5808 = pi0230 & ~w5807;
assign w5809 = ~pi0230 & pi0245;
assign w5810 = ~w5808 & ~w5809;
assign w5811 = pi1148 & w5469;
assign w5812 = pi1150 & ~w3310;
assign w5813 = pi1149 & w3310;
assign w5814 = ~w5812 & ~w5813;
assign w5815 = ~w3185 & ~w5814;
assign w5816 = ~w5811 & ~w5815;
assign w5817 = w5467 & ~w5816;
assign w5818 = ~w5496 & w5817;
assign w5819 = w5496 & w5804;
assign w5820 = ~w5818 & ~w5819;
assign w5821 = pi0230 & ~w5820;
assign w5822 = ~pi0230 & pi0246;
assign w5823 = ~w5821 & ~w5822;
assign w5824 = ~w5496 & w5712;
assign w5825 = w5496 & w5692;
assign w5826 = ~w5824 & ~w5825;
assign w5827 = pi0230 & ~w5826;
assign w5828 = ~pi0230 & pi0247;
assign w5829 = ~w5827 & ~w5828;
assign w5830 = pi1150 & w5469;
assign w5831 = pi1152 & ~w3310;
assign w5832 = pi1151 & w3310;
assign w5833 = ~w5831 & ~w5832;
assign w5834 = ~w3185 & ~w5833;
assign w5835 = ~w5830 & ~w5834;
assign w5836 = w5467 & ~w5835;
assign w5837 = ~w5496 & w5836;
assign w5838 = w5496 & w5817;
assign w5839 = ~w5837 & ~w5838;
assign w5840 = pi0230 & ~w5839;
assign w5841 = ~pi0230 & pi0248;
assign w5842 = ~w5840 & ~w5841;
assign w5843 = w5496 & w5836;
assign w5844 = ~w5496 & w5503;
assign w5845 = ~w5843 & ~w5844;
assign w5846 = pi0230 & ~w5845;
assign w5847 = ~pi0230 & pi0249;
assign w5848 = ~w5846 & ~w5847;
assign w5849 = ~w3276 & ~w4023;
assign w5850 = ~pi0250 & ~w5849;
assign w5851 = ~pi0200 & pi1053;
assign w5852 = pi0200 & pi1039;
assign w5853 = ~w5851 & ~w5852;
assign w5854 = ~pi0200 & pi0897;
assign w5855 = pi0200 & ~pi0476;
assign w5856 = ~w5854 & ~w5855;
assign w5857 = ~pi0199 & ~w5856;
assign w5858 = ~w5853 & w5857;
assign w5859 = pi0251 & ~w5857;
assign w5860 = ~w5858 & ~w5859;
assign w5861 = w1233 & w1649;
assign w5862 = w3031 & w5861;
assign w5863 = pi1093 & ~w2045;
assign w5864 = pi0252 & ~w5863;
assign w5865 = pi1092 & w5864;
assign w5866 = ~w5862 & ~w5865;
assign w5867 = pi1151 & ~w5774;
assign w5868 = pi1153 & ~w5778;
assign w5869 = ~w5867 & ~w5868;
assign w5870 = pi1152 & ~w5785;
assign w5871 = w5869 & ~w5870;
assign w5872 = ~w5766 & ~w5871;
assign w5873 = w5748 & w5751;
assign w5874 = pi0268 & w5873;
assign w5875 = w5755 & w5874;
assign w5876 = ~pi0253 & ~w5875;
assign w5877 = pi0253 & pi0275;
assign w5878 = pi0272 & w5877;
assign w5879 = w5874 & w5878;
assign w5880 = ~w5876 & ~w5879;
assign w5881 = w5766 & w5880;
assign w5882 = ~w5872 & ~w5881;
assign w5883 = w5754 & w5755;
assign w5884 = ~pi0254 & w5883;
assign w5885 = pi0254 & ~w5883;
assign w5886 = ~w5884 & ~w5885;
assign w5887 = w5766 & ~w5886;
assign w5888 = pi1152 & ~w5774;
assign w5889 = pi1154 & ~w5778;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = pi1153 & ~w5785;
assign w5892 = w5890 & ~w5891;
assign w5893 = ~w5766 & ~w5892;
assign w5894 = ~w5887 & ~w5893;
assign w5895 = ~pi0200 & pi1049;
assign w5896 = pi0200 & pi1036;
assign w5897 = ~w5895 & ~w5896;
assign w5898 = w5857 & ~w5897;
assign w5899 = pi0255 & ~w5857;
assign w5900 = ~w5898 & ~w5899;
assign w5901 = ~pi0200 & pi1048;
assign w5902 = pi0200 & pi1070;
assign w5903 = ~w5901 & ~w5902;
assign w5904 = w5857 & ~w5903;
assign w5905 = pi0256 & ~w5857;
assign w5906 = ~w5904 & ~w5905;
assign w5907 = ~pi0200 & pi1084;
assign w5908 = pi0200 & pi1065;
assign w5909 = ~w5907 & ~w5908;
assign w5910 = w5857 & ~w5909;
assign w5911 = pi0257 & ~w5857;
assign w5912 = ~w5910 & ~w5911;
assign w5913 = ~pi0200 & pi1072;
assign w5914 = pi0200 & pi1062;
assign w5915 = ~w5913 & ~w5914;
assign w5916 = w5857 & ~w5915;
assign w5917 = pi0258 & ~w5857;
assign w5918 = ~w5916 & ~w5917;
assign w5919 = ~pi0200 & pi1059;
assign w5920 = pi0200 & pi1069;
assign w5921 = ~w5919 & ~w5920;
assign w5922 = w5857 & ~w5921;
assign w5923 = pi0259 & ~w5857;
assign w5924 = ~w5922 & ~w5923;
assign w5925 = ~pi0200 & pi1044;
assign w5926 = pi0200 & pi1067;
assign w5927 = ~w5925 & ~w5926;
assign w5928 = w5857 & ~w5927;
assign w5929 = pi0260 & ~w5857;
assign w5930 = ~w5928 & ~w5929;
assign w5931 = ~pi0200 & pi1037;
assign w5932 = pi0200 & pi1040;
assign w5933 = ~w5931 & ~w5932;
assign w5934 = w5857 & ~w5933;
assign w5935 = pi0261 & ~w5857;
assign w5936 = ~w5934 & ~w5935;
assign w5937 = ~pi0228 & pi1093;
assign w5938 = ~pi0123 & pi0228;
assign w5939 = ~w5937 & ~w5938;
assign w5940 = pi1142 & ~w5939;
assign w5941 = ~w3185 & w5467;
assign w5942 = w5940 & w5941;
assign w5943 = ~pi0262 & w5939;
assign w5944 = ~w5942 & ~w5943;
assign w5945 = pi0263 & pi0267;
assign w5946 = pi0254 & w5883;
assign w5947 = w5945 & w5946;
assign w5948 = pi0254 & pi0267;
assign w5949 = w5883 & w5948;
assign w5950 = ~pi0263 & ~w5949;
assign w5951 = ~w5947 & ~w5950;
assign w5952 = w5766 & ~w5951;
assign w5953 = pi1154 & ~w5774;
assign w5954 = pi1156 & ~w5778;
assign w5955 = ~w5953 & ~w5954;
assign w5956 = pi1155 & ~w5785;
assign w5957 = w5955 & ~w5956;
assign w5958 = ~w5766 & ~w5957;
assign w5959 = ~w5952 & ~w5958;
assign w5960 = (w5740 & w5742) | (w5740 & w5746) | (w5742 & w5746);
assign w5961 = ~pi0264 & ~w5960;
assign w5962 = pi0796 & w5960;
assign w5963 = ~w5961 & ~w5962;
assign w5964 = w5766 & ~w5963;
assign w5965 = pi1141 & ~w5774;
assign w5966 = pi1143 & ~w5778;
assign w5967 = ~w5965 & ~w5966;
assign w5968 = pi1142 & ~w5785;
assign w5969 = w5967 & ~w5968;
assign w5970 = ~w5766 & ~w5969;
assign w5971 = ~w5964 & ~w5970;
assign w5972 = ~pi0265 & ~w5960;
assign w5973 = pi0819 & w5960;
assign w5974 = ~w5972 & ~w5973;
assign w5975 = w5766 & ~w5974;
assign w5976 = pi1142 & ~w5774;
assign w5977 = pi1144 & ~w5778;
assign w5978 = ~w5976 & ~w5977;
assign w5979 = pi1143 & ~w5785;
assign w5980 = w5978 & ~w5979;
assign w5981 = ~w5766 & ~w5980;
assign w5982 = ~w5975 & ~w5981;
assign w5983 = pi0266 & ~w5960;
assign w5984 = pi0948 & w5960;
assign w5985 = ~w5983 & ~w5984;
assign w5986 = w5766 & ~w5985;
assign w5987 = pi1134 & ~w5774;
assign w5988 = pi1136 & ~w5778;
assign w5989 = ~w5987 & ~w5988;
assign w5990 = pi1135 & ~w5785;
assign w5991 = w5989 & ~w5990;
assign w5992 = ~w5766 & ~w5991;
assign w5993 = ~w5986 & ~w5992;
assign w5994 = pi0254 & ~pi0267;
assign w5995 = w5883 & w5994;
assign w5996 = pi0267 & ~w5946;
assign w5997 = ~w5995 & ~w5996;
assign w5998 = w5766 & ~w5997;
assign w5999 = pi1153 & ~w5774;
assign w6000 = pi1155 & ~w5778;
assign w6001 = ~w5999 & ~w6000;
assign w6002 = pi1154 & ~w5785;
assign w6003 = w6001 & ~w6002;
assign w6004 = ~w5766 & ~w6003;
assign w6005 = ~w5998 & ~w6004;
assign w6006 = w5755 & w5873;
assign w6007 = pi0268 & ~w6006;
assign w6008 = ~pi0268 & pi0275;
assign w6009 = pi0272 & w5873;
assign w6010 = w6008 & w6009;
assign w6011 = ~w6007 & ~w6010;
assign w6012 = w5766 & ~w6011;
assign w6013 = pi1150 & ~w5774;
assign w6014 = pi1152 & ~w5778;
assign w6015 = ~w6013 & ~w6014;
assign w6016 = pi1151 & ~w5785;
assign w6017 = w6015 & ~w6016;
assign w6018 = ~w5766 & ~w6017;
assign w6019 = ~w6012 & ~w6018;
assign w6020 = ~pi0269 & ~w5960;
assign w6021 = pi0817 & w5960;
assign w6022 = ~w6020 & ~w6021;
assign w6023 = w5766 & ~w6022;
assign w6024 = pi1136 & ~w5774;
assign w6025 = pi1138 & ~w5778;
assign w6026 = ~w6024 & ~w6025;
assign w6027 = pi1137 & ~w5785;
assign w6028 = w6026 & ~w6027;
assign w6029 = ~w5766 & ~w6028;
assign w6030 = ~w6023 & ~w6029;
assign w6031 = ~pi0270 & ~w5960;
assign w6032 = pi0805 & w5960;
assign w6033 = ~w6031 & ~w6032;
assign w6034 = w5766 & ~w6033;
assign w6035 = pi1139 & ~w5774;
assign w6036 = pi1141 & ~w5778;
assign w6037 = ~w6035 & ~w6036;
assign w6038 = pi1140 & ~w5785;
assign w6039 = w6037 & ~w6038;
assign w6040 = ~w5766 & ~w6039;
assign w6041 = ~w6034 & ~w6040;
assign w6042 = pi0276 & pi0802;
assign w6043 = w5960 & w6042;
assign w6044 = pi0271 & ~w6043;
assign w6045 = ~pi0271 & pi0802;
assign w6046 = pi0276 & w5960;
assign w6047 = w6045 & w6046;
assign w6048 = ~w6044 & ~w6047;
assign w6049 = w5766 & ~w6048;
assign w6050 = pi1145 & ~w5774;
assign w6051 = pi1147 & ~w5778;
assign w6052 = ~w6050 & ~w6051;
assign w6053 = pi1146 & ~w5785;
assign w6054 = w6052 & ~w6053;
assign w6055 = ~w5766 & ~w6054;
assign w6056 = ~w6049 & ~w6055;
assign w6057 = ~pi0272 & w5873;
assign w6058 = pi0272 & ~w5873;
assign w6059 = ~w6057 & ~w6058;
assign w6060 = w5766 & ~w6059;
assign w6061 = pi1148 & ~w5774;
assign w6062 = pi1150 & ~w5778;
assign w6063 = ~w6061 & ~w6062;
assign w6064 = pi1149 & ~w5785;
assign w6065 = w6063 & ~w6064;
assign w6066 = ~w5766 & ~w6065;
assign w6067 = ~w6060 & ~w6066;
assign w6068 = pi1146 & ~w5774;
assign w6069 = pi1148 & ~w5778;
assign w6070 = ~w6068 & ~w6069;
assign w6071 = pi1147 & ~w5785;
assign w6072 = w6070 & ~w6071;
assign w6073 = ~w5766 & ~w6072;
assign w6074 = w5748 & w6042;
assign w6075 = ~pi0273 & ~w6074;
assign w6076 = pi0273 & pi0802;
assign w6077 = pi0276 & w6076;
assign w6078 = w5748 & w6077;
assign w6079 = ~w6075 & ~w6078;
assign w6080 = w5766 & w6079;
assign w6081 = ~w6073 & ~w6080;
assign w6082 = ~pi0274 & ~w5960;
assign w6083 = pi0659 & w5960;
assign w6084 = ~w6082 & ~w6083;
assign w6085 = w5766 & ~w6084;
assign w6086 = pi1143 & ~w5774;
assign w6087 = pi1145 & ~w5778;
assign w6088 = ~w6086 & ~w6087;
assign w6089 = pi1144 & ~w5785;
assign w6090 = w6088 & ~w6089;
assign w6091 = ~w5766 & ~w6090;
assign w6092 = ~w6085 & ~w6091;
assign w6093 = pi0272 & ~pi0275;
assign w6094 = w5873 & w6093;
assign w6095 = pi0275 & ~w6009;
assign w6096 = ~w6094 & ~w6095;
assign w6097 = w5766 & ~w6096;
assign w6098 = pi1149 & ~w5774;
assign w6099 = pi1151 & ~w5778;
assign w6100 = ~w6098 & ~w6099;
assign w6101 = pi1150 & ~w5785;
assign w6102 = w6100 & ~w6101;
assign w6103 = ~w5766 & ~w6102;
assign w6104 = ~w6097 & ~w6103;
assign w6105 = ~pi0276 & pi0802;
assign w6106 = w5960 & w6105;
assign w6107 = pi0802 & w5960;
assign w6108 = pi0276 & ~w6107;
assign w6109 = ~w6106 & ~w6108;
assign w6110 = w5766 & ~w6109;
assign w6111 = pi1144 & ~w5774;
assign w6112 = pi1146 & ~w5778;
assign w6113 = ~w6111 & ~w6112;
assign w6114 = pi1145 & ~w5785;
assign w6115 = w6113 & ~w6114;
assign w6116 = ~w5766 & ~w6115;
assign w6117 = ~w6110 & ~w6116;
assign w6118 = ~pi0277 & ~w5960;
assign w6119 = pi0820 & w5960;
assign w6120 = ~w6118 & ~w6119;
assign w6121 = w5766 & ~w6120;
assign w6122 = pi1140 & ~w5774;
assign w6123 = pi1142 & ~w5778;
assign w6124 = ~w6122 & ~w6123;
assign w6125 = pi1141 & ~w5785;
assign w6126 = w6124 & ~w6125;
assign w6127 = ~w5766 & ~w6126;
assign w6128 = ~w6121 & ~w6127;
assign w6129 = pi0278 & ~w5960;
assign w6130 = pi0976 & w5960;
assign w6131 = ~w6129 & ~w6130;
assign w6132 = w5766 & ~w6131;
assign w6133 = pi1132 & ~w5774;
assign w6134 = pi1134 & ~w5778;
assign w6135 = ~w6133 & ~w6134;
assign w6136 = pi1133 & ~w5785;
assign w6137 = w6135 & ~w6136;
assign w6138 = ~w5766 & ~w6137;
assign w6139 = ~w6132 & ~w6138;
assign w6140 = pi0279 & ~w5960;
assign w6141 = pi0958 & w5960;
assign w6142 = ~w6140 & ~w6141;
assign w6143 = w5766 & ~w6142;
assign w6144 = pi1133 & ~w5774;
assign w6145 = pi1135 & ~w5778;
assign w6146 = ~w6144 & ~w6145;
assign w6147 = pi1134 & ~w5785;
assign w6148 = w6146 & ~w6147;
assign w6149 = ~w5766 & ~w6148;
assign w6150 = ~w6143 & ~w6149;
assign w6151 = ~pi0280 & ~w5960;
assign w6152 = pi0914 & w5960;
assign w6153 = ~w6151 & ~w6152;
assign w6154 = w5766 & ~w6153;
assign w6155 = pi1135 & ~w5774;
assign w6156 = pi1137 & ~w5778;
assign w6157 = ~w6155 & ~w6156;
assign w6158 = pi1136 & ~w5785;
assign w6159 = w6157 & ~w6158;
assign w6160 = ~w5766 & ~w6159;
assign w6161 = ~w6154 & ~w6160;
assign w6162 = ~pi0281 & ~w5960;
assign w6163 = pi0830 & w5960;
assign w6164 = ~w6162 & ~w6163;
assign w6165 = w5766 & ~w6164;
assign w6166 = pi1137 & ~w5774;
assign w6167 = pi1139 & ~w5778;
assign w6168 = ~w6166 & ~w6167;
assign w6169 = pi1138 & ~w5785;
assign w6170 = w6168 & ~w6169;
assign w6171 = ~w5766 & ~w6170;
assign w6172 = ~w6165 & ~w6171;
assign w6173 = ~pi0282 & ~w5960;
assign w6174 = pi0836 & w5960;
assign w6175 = ~w6173 & ~w6174;
assign w6176 = w5766 & ~w6175;
assign w6177 = pi1138 & ~w5774;
assign w6178 = pi1140 & ~w5778;
assign w6179 = ~w6177 & ~w6178;
assign w6180 = pi1139 & ~w5785;
assign w6181 = w6179 & ~w6180;
assign w6182 = ~w5766 & ~w6181;
assign w6183 = ~w6176 & ~w6182;
assign w6184 = pi1147 & ~w5774;
assign w6185 = pi1149 & ~w5778;
assign w6186 = ~w6184 & ~w6185;
assign w6187 = pi1148 & ~w5785;
assign w6188 = w6186 & ~w6187;
assign w6189 = ~w5766 & ~w6188;
assign w6190 = pi0271 & pi0273;
assign w6191 = w5960 & w6190;
assign w6192 = pi0283 & pi0802;
assign w6193 = pi0276 & w6192;
assign w6194 = w6191 & w6193;
assign w6195 = pi0273 & w6042;
assign w6196 = w5748 & w6195;
assign w6197 = ~pi0283 & ~w6196;
assign w6198 = ~w6194 & ~w6197;
assign w6199 = w5766 & w6198;
assign w6200 = ~w6189 & ~w6199;
assign w6201 = pi1143 & ~w5939;
assign w6202 = w3311 & w5467;
assign w6203 = w6201 & w6202;
assign w6204 = ~pi0284 & w5939;
assign w6205 = ~w6203 & ~w6204;
assign w6206 = w94 & w3123;
assign w6207 = (w94 & w3128) | (w94 & w6206) | (w3128 & w6206);
assign w6208 = ~pi0086 & w6207;
assign w6209 = w3005 & w6208;
assign w6210 = w95 & w112;
assign w6211 = w6209 & w6210;
assign w6212 = ~pi0288 & pi0289;
assign w6213 = ~w2040 & w6212;
assign w6214 = pi0286 & w3265;
assign w6215 = pi0288 & ~pi0289;
assign w6216 = w6214 & w6215;
assign w6217 = ~w6212 & ~w6216;
assign w6218 = ~w2040 & ~w6217;
assign w6219 = (w6211 & w6213) | (w6211 & w6218) | (w6213 & w6218);
assign w6220 = pi0286 & ~pi0288;
assign w6221 = ~pi0286 & ~w3265;
assign w6222 = ~pi0288 & ~w6221;
assign w6223 = (w6211 & w6220) | (w6211 & w6222) | (w6220 & w6222);
assign w6224 = pi0288 & ~w6214;
assign w6225 = (pi0288 & ~w6211) | (pi0288 & w6224) | (~w6211 & w6224);
assign w6226 = ~w6223 & ~w6225;
assign w6227 = ~pi0289 & ~w6219;
assign w6228 = (~w6219 & w6226) | (~w6219 & w6227) | (w6226 & w6227);
assign w6229 = pi0288 & pi0289;
assign w6230 = ~pi0286 & w2042;
assign w6231 = pi0285 & w6230;
assign w6232 = ~w6229 & ~w6231;
assign w6233 = w2040 & ~w6232;
assign w6234 = pi0285 & ~w3265;
assign w6235 = w6230 & w6234;
assign w6236 = ~w6229 & ~w6235;
assign w6237 = w2040 & ~w6236;
assign w6238 = (~w6211 & w6233) | (~w6211 & w6237) | (w6233 & w6237);
assign w6239 = pi0286 & pi0289;
assign w6240 = ~w6238 & ~w6239;
assign w6241 = w6228 & w6240;
assign w6242 = pi0289 & w6238;
assign w6243 = (pi0289 & ~w6228) | (pi0289 & w6242) | (~w6228 & w6242);
assign w6244 = ~w6241 & ~w6243;
assign w6245 = pi0285 & ~w6244;
assign w6246 = ~pi0285 & ~w6238;
assign w6247 = pi0289 & w6246;
assign w6248 = w6228 & w6247;
assign w6249 = pi0285 & w6238;
assign w6250 = (pi0285 & ~w6228) | (pi0285 & w6249) | (~w6228 & w6249);
assign w6251 = ~w6248 & ~w6250;
assign w6252 = pi0286 & ~w6251;
assign w6253 = ~w6245 & ~w6252;
assign w6254 = ~pi0793 & ~w6253;
assign w6255 = ~pi0288 & ~w4043;
assign w6256 = pi0288 & w4043;
assign w6257 = ~w6255 & ~w6256;
assign w6258 = pi0286 & ~w6257;
assign w6259 = w3265 & w6211;
assign w6260 = ~pi0286 & ~pi0288;
assign w6261 = w4043 & w6260;
assign w6262 = pi0286 & pi0288;
assign w6263 = ~w6261 & ~w6262;
assign w6264 = ~w6259 & ~w6263;
assign w6265 = ~w6258 & ~w6264;
assign w6266 = ~pi0286 & pi0288;
assign w6267 = ~w4043 & w6266;
assign w6268 = ~w6220 & ~w6267;
assign w6269 = w6259 & ~w6268;
assign w6270 = w6265 & ~w6269;
assign w6271 = ~pi0793 & ~w6270;
assign w6272 = ~pi0287 & pi0457;
assign w6273 = ~pi0332 & ~w6272;
assign w6274 = ~pi0288 & w6259;
assign w6275 = w2043 & w6274;
assign w6276 = pi0288 & ~w6259;
assign w6277 = ~w6274 & ~w6276;
assign w6278 = ~w2040 & ~w6277;
assign w6279 = ~w6275 & ~w6278;
assign w6280 = ~pi0288 & ~w6259;
assign w6281 = ~w2043 & w6280;
assign w6282 = pi0288 & w6259;
assign w6283 = ~w6281 & ~w6282;
assign w6284 = w2040 & ~w6283;
assign w6285 = w6279 & ~w6284;
assign w6286 = ~pi0793 & ~w6285;
assign w6287 = w6228 & ~w6238;
assign w6288 = ~pi0793 & ~w6287;
assign w6289 = ~pi0476 & pi1048;
assign w6290 = pi0290 & pi0476;
assign w6291 = ~w6289 & ~w6290;
assign w6292 = ~pi0476 & pi1049;
assign w6293 = pi0291 & pi0476;
assign w6294 = ~w6292 & ~w6293;
assign w6295 = ~pi0476 & pi1084;
assign w6296 = pi0292 & pi0476;
assign w6297 = ~w6295 & ~w6296;
assign w6298 = ~pi0476 & pi1059;
assign w6299 = pi0293 & pi0476;
assign w6300 = ~w6298 & ~w6299;
assign w6301 = ~pi0476 & pi1072;
assign w6302 = pi0294 & pi0476;
assign w6303 = ~w6301 & ~w6302;
assign w6304 = ~pi0476 & pi1053;
assign w6305 = pi0295 & pi0476;
assign w6306 = ~w6304 & ~w6305;
assign w6307 = ~pi0476 & pi1037;
assign w6308 = pi0296 & pi0476;
assign w6309 = ~w6307 & ~w6308;
assign w6310 = ~pi0476 & pi1044;
assign w6311 = pi0297 & pi0476;
assign w6312 = ~w6310 & ~w6311;
assign w6313 = ~pi0478 & pi1044;
assign w6314 = pi0298 & pi0478;
assign w6315 = ~w6313 & ~w6314;
assign w6316 = w529 & w5122;
assign w6317 = ~w3319 & ~w6316;
assign w6318 = pi0039 & w3024;
assign w6319 = ~pi0287 & w6318;
assign w6320 = ~pi0979 & w6319;
assign w6321 = w6317 & ~w6320;
assign w6322 = ~w3332 & w6321;
assign w6323 = ~pi0024 & w1338;
assign w6324 = pi0057 & w6323;
assign w6325 = ~pi0059 & w6324;
assign w6326 = ~pi0312 & w6325;
assign w6327 = pi0300 & w6326;
assign w6328 = ~pi0300 & ~w6326;
assign w6329 = ~w6327 & ~w6328;
assign w6330 = ~pi0055 & ~w6329;
assign w6331 = ~pi0300 & pi0301;
assign w6332 = w6326 & w6331;
assign w6333 = ~pi0300 & w6326;
assign w6334 = ~pi0301 & ~w6333;
assign w6335 = ~w6332 & ~w6334;
assign w6336 = ~pi0055 & ~w6335;
assign w6337 = pi1148 & w1225;
assign w6338 = ~w526 & w666;
assign w6339 = w526 & w648;
assign w6340 = ~w6338 & ~w6339;
assign w6341 = pi0273 & ~w6340;
assign w6342 = ~w6337 & ~w6341;
assign w6343 = w114 & ~w526;
assign w6344 = w16 & w526;
assign w6345 = ~w6343 & ~w6344;
assign w6346 = ~pi0237 & ~w6345;
assign w6347 = ~w526 & w610;
assign w6348 = w526 & w675;
assign w6349 = ~w6347 & ~w6348;
assign w6350 = pi0937 & ~w6349;
assign w6351 = ~w6346 & ~w6350;
assign w6352 = w6342 & w6351;
assign w6353 = ~pi0478 & pi1049;
assign w6354 = pi0303 & pi0478;
assign w6355 = ~w6353 & ~w6354;
assign w6356 = ~pi0478 & pi1048;
assign w6357 = pi0304 & pi0478;
assign w6358 = ~w6356 & ~w6357;
assign w6359 = ~pi0478 & pi1084;
assign w6360 = pi0305 & pi0478;
assign w6361 = ~w6359 & ~w6360;
assign w6362 = ~pi0478 & pi1059;
assign w6363 = pi0306 & pi0478;
assign w6364 = ~w6362 & ~w6363;
assign w6365 = ~pi0478 & pi1053;
assign w6366 = pi0307 & pi0478;
assign w6367 = ~w6365 & ~w6366;
assign w6368 = ~pi0478 & pi1037;
assign w6369 = pi0308 & pi0478;
assign w6370 = ~w6368 & ~w6369;
assign w6371 = ~pi0478 & pi1072;
assign w6372 = pi0309 & pi0478;
assign w6373 = ~w6371 & ~w6372;
assign w6374 = pi1147 & w1225;
assign w6375 = pi0271 & ~w6340;
assign w6376 = ~w6374 & ~w6375;
assign w6377 = ~pi0233 & ~w6345;
assign w6378 = pi0934 & ~w6349;
assign w6379 = ~w6377 & ~w6378;
assign w6380 = w6376 & w6379;
assign w6381 = pi0301 & pi0311;
assign w6382 = w6333 & w6381;
assign w6383 = ~pi0311 & ~w6332;
assign w6384 = ~w6382 & ~w6383;
assign w6385 = ~pi0055 & ~w6384;
assign w6386 = ~pi0059 & ~pi0312;
assign w6387 = pi0057 & w6386;
assign w6388 = w6323 & w6387;
assign w6389 = w571 & w6323;
assign w6390 = pi0312 & ~w6389;
assign w6391 = ~w6388 & ~w6390;
assign w6392 = ~pi0055 & ~w6391;
assign w6393 = pi0314 & w2568;
assign w6394 = w3872 & ~w6393;
assign w6395 = ~w2568 & w3848;
assign w6396 = ~w6394 & ~w6395;
assign w6397 = ~pi0954 & ~w6396;
assign w6398 = ~pi0313 & pi0954;
assign w6399 = ~w6397 & ~w6398;
assign w6400 = ~w4376 & w4441;
assign w6401 = w4256 & w6400;
assign w6402 = ~pi0121 & w6401;
assign w6403 = ~pi0125 & w6402;
assign w6404 = ~pi0133 & w6403;
assign w6405 = ~pi0340 & w6259;
assign w6406 = pi1080 & w6405;
assign w6407 = pi0315 & ~w6405;
assign w6408 = ~w6406 & ~w6407;
assign w6409 = pi1047 & w6405;
assign w6410 = pi0316 & ~w6405;
assign w6411 = ~w6409 & ~w6410;
assign w6412 = ~pi0330 & w6259;
assign w6413 = pi1078 & w6412;
assign w6414 = pi0317 & ~w6412;
assign w6415 = ~w6413 & ~w6414;
assign w6416 = ~pi0341 & w6259;
assign w6417 = pi1074 & w6416;
assign w6418 = pi0318 & ~w6416;
assign w6419 = ~w6417 & ~w6418;
assign w6420 = pi1072 & w6416;
assign w6421 = pi0319 & ~w6416;
assign w6422 = ~w6420 & ~w6421;
assign w6423 = pi1048 & w6405;
assign w6424 = pi0320 & ~w6405;
assign w6425 = ~w6423 & ~w6424;
assign w6426 = pi1058 & w6405;
assign w6427 = pi0321 & ~w6405;
assign w6428 = ~w6426 & ~w6427;
assign w6429 = pi1051 & w6405;
assign w6430 = pi0322 & ~w6405;
assign w6431 = ~w6429 & ~w6430;
assign w6432 = pi1065 & w6405;
assign w6433 = pi0323 & ~w6405;
assign w6434 = ~w6432 & ~w6433;
assign w6435 = pi1086 & w6416;
assign w6436 = pi0324 & ~w6416;
assign w6437 = ~w6435 & ~w6436;
assign w6438 = pi1063 & w6416;
assign w6439 = pi0325 & ~w6416;
assign w6440 = ~w6438 & ~w6439;
assign w6441 = pi1057 & w6416;
assign w6442 = pi0326 & ~w6416;
assign w6443 = ~w6441 & ~w6442;
assign w6444 = pi1040 & w6405;
assign w6445 = pi0327 & ~w6405;
assign w6446 = ~w6444 & ~w6445;
assign w6447 = pi1058 & w6416;
assign w6448 = pi0328 & ~w6416;
assign w6449 = ~w6447 & ~w6448;
assign w6450 = pi1043 & w6416;
assign w6451 = pi0329 & ~w6416;
assign w6452 = ~w6450 & ~w6451;
assign w6453 = ~pi0330 & ~w6259;
assign w6454 = ~w6405 & ~w6453;
assign w6455 = ~w1234 & ~w6454;
assign w6456 = pi1092 & w6455;
assign w6457 = ~pi0331 & ~w6259;
assign w6458 = ~w6416 & ~w6457;
assign w6459 = ~w1234 & ~w6458;
assign w6460 = pi1092 & w6459;
assign w6461 = ~pi0070 & ~pi0089;
assign w6462 = w2554 & ~w6461;
assign w6463 = pi0332 & w6462;
assign w6464 = pi0287 & w1649;
assign w6465 = ~w3240 & ~w6464;
assign w6466 = ~w6463 & w6465;
assign w6467 = ~w1615 & w6466;
assign w6468 = pi1040 & w6416;
assign w6469 = pi0333 & ~w6416;
assign w6470 = ~w6468 & ~w6469;
assign w6471 = pi1065 & w6416;
assign w6472 = pi0334 & ~w6416;
assign w6473 = ~w6471 & ~w6472;
assign w6474 = pi1069 & w6416;
assign w6475 = pi0335 & ~w6416;
assign w6476 = ~w6474 & ~w6475;
assign w6477 = pi1070 & w6412;
assign w6478 = pi0336 & ~w6412;
assign w6479 = ~w6477 & ~w6478;
assign w6480 = pi1044 & w6412;
assign w6481 = pi0337 & ~w6412;
assign w6482 = ~w6480 & ~w6481;
assign w6483 = pi1072 & w6412;
assign w6484 = pi0338 & ~w6412;
assign w6485 = ~w6483 & ~w6484;
assign w6486 = pi1086 & w6412;
assign w6487 = pi0339 & ~w6412;
assign w6488 = ~w6486 & ~w6487;
assign w6489 = ~pi0331 & w6259;
assign w6490 = ~w1234 & ~w6489;
assign w6491 = ~pi0340 & ~w6259;
assign w6492 = pi1092 & ~w6491;
assign w6493 = w6490 & w6492;
assign w6494 = ~pi0341 & ~w6259;
assign w6495 = ~w6412 & ~w6494;
assign w6496 = ~w1234 & ~w6495;
assign w6497 = pi1092 & w6496;
assign w6498 = pi1049 & w6405;
assign w6499 = pi0342 & ~w6405;
assign w6500 = ~w6498 & ~w6499;
assign w6501 = pi1062 & w6405;
assign w6502 = pi0343 & ~w6405;
assign w6503 = ~w6501 & ~w6502;
assign w6504 = pi1069 & w6405;
assign w6505 = pi0344 & ~w6405;
assign w6506 = ~w6504 & ~w6505;
assign w6507 = pi1039 & w6405;
assign w6508 = pi0345 & ~w6405;
assign w6509 = ~w6507 & ~w6508;
assign w6510 = pi1067 & w6405;
assign w6511 = pi0346 & ~w6405;
assign w6512 = ~w6510 & ~w6511;
assign w6513 = pi1055 & w6405;
assign w6514 = pi0347 & ~w6405;
assign w6515 = ~w6513 & ~w6514;
assign w6516 = pi1087 & w6405;
assign w6517 = pi0348 & ~w6405;
assign w6518 = ~w6516 & ~w6517;
assign w6519 = pi1043 & w6405;
assign w6520 = pi0349 & ~w6405;
assign w6521 = ~w6519 & ~w6520;
assign w6522 = pi1035 & w6405;
assign w6523 = pi0350 & ~w6405;
assign w6524 = ~w6522 & ~w6523;
assign w6525 = pi1079 & w6405;
assign w6526 = pi0351 & ~w6405;
assign w6527 = ~w6525 & ~w6526;
assign w6528 = pi1078 & w6405;
assign w6529 = pi0352 & ~w6405;
assign w6530 = ~w6528 & ~w6529;
assign w6531 = pi1063 & w6405;
assign w6532 = pi0353 & ~w6405;
assign w6533 = ~w6531 & ~w6532;
assign w6534 = pi1045 & w6405;
assign w6535 = pi0354 & ~w6405;
assign w6536 = ~w6534 & ~w6535;
assign w6537 = pi1084 & w6405;
assign w6538 = pi0355 & ~w6405;
assign w6539 = ~w6537 & ~w6538;
assign w6540 = pi1081 & w6405;
assign w6541 = pi0356 & ~w6405;
assign w6542 = ~w6540 & ~w6541;
assign w6543 = pi1076 & w6405;
assign w6544 = pi0357 & ~w6405;
assign w6545 = ~w6543 & ~w6544;
assign w6546 = pi1071 & w6405;
assign w6547 = pi0358 & ~w6405;
assign w6548 = ~w6546 & ~w6547;
assign w6549 = pi1068 & w6405;
assign w6550 = pi0359 & ~w6405;
assign w6551 = ~w6549 & ~w6550;
assign w6552 = pi1042 & w6405;
assign w6553 = pi0360 & ~w6405;
assign w6554 = ~w6552 & ~w6553;
assign w6555 = pi1059 & w6405;
assign w6556 = pi0361 & ~w6405;
assign w6557 = ~w6555 & ~w6556;
assign w6558 = pi1070 & w6405;
assign w6559 = pi0362 & ~w6405;
assign w6560 = ~w6558 & ~w6559;
assign w6561 = pi1049 & w6412;
assign w6562 = pi0363 & ~w6412;
assign w6563 = ~w6561 & ~w6562;
assign w6564 = pi1062 & w6412;
assign w6565 = pi0364 & ~w6412;
assign w6566 = ~w6564 & ~w6565;
assign w6567 = pi1065 & w6412;
assign w6568 = pi0365 & ~w6412;
assign w6569 = ~w6567 & ~w6568;
assign w6570 = pi1069 & w6412;
assign w6571 = pi0366 & ~w6412;
assign w6572 = ~w6570 & ~w6571;
assign w6573 = pi1039 & w6412;
assign w6574 = pi0367 & ~w6412;
assign w6575 = ~w6573 & ~w6574;
assign w6576 = pi1067 & w6412;
assign w6577 = pi0368 & ~w6412;
assign w6578 = ~w6576 & ~w6577;
assign w6579 = pi1080 & w6412;
assign w6580 = pi0369 & ~w6412;
assign w6581 = ~w6579 & ~w6580;
assign w6582 = pi1055 & w6412;
assign w6583 = pi0370 & ~w6412;
assign w6584 = ~w6582 & ~w6583;
assign w6585 = pi1051 & w6412;
assign w6586 = pi0371 & ~w6412;
assign w6587 = ~w6585 & ~w6586;
assign w6588 = pi1048 & w6412;
assign w6589 = pi0372 & ~w6412;
assign w6590 = ~w6588 & ~w6589;
assign w6591 = pi1087 & w6412;
assign w6592 = pi0373 & ~w6412;
assign w6593 = ~w6591 & ~w6592;
assign w6594 = pi1035 & w6412;
assign w6595 = pi0374 & ~w6412;
assign w6596 = ~w6594 & ~w6595;
assign w6597 = pi1047 & w6412;
assign w6598 = pi0375 & ~w6412;
assign w6599 = ~w6597 & ~w6598;
assign w6600 = pi1079 & w6412;
assign w6601 = pi0376 & ~w6412;
assign w6602 = ~w6600 & ~w6601;
assign w6603 = pi1074 & w6412;
assign w6604 = pi0377 & ~w6412;
assign w6605 = ~w6603 & ~w6604;
assign w6606 = pi1063 & w6412;
assign w6607 = pi0378 & ~w6412;
assign w6608 = ~w6606 & ~w6607;
assign w6609 = pi1045 & w6412;
assign w6610 = pi0379 & ~w6412;
assign w6611 = ~w6609 & ~w6610;
assign w6612 = pi1084 & w6412;
assign w6613 = pi0380 & ~w6412;
assign w6614 = ~w6612 & ~w6613;
assign w6615 = pi1081 & w6412;
assign w6616 = pi0381 & ~w6412;
assign w6617 = ~w6615 & ~w6616;
assign w6618 = pi1076 & w6412;
assign w6619 = pi0382 & ~w6412;
assign w6620 = ~w6618 & ~w6619;
assign w6621 = pi1071 & w6412;
assign w6622 = pi0383 & ~w6412;
assign w6623 = ~w6621 & ~w6622;
assign w6624 = pi1068 & w6412;
assign w6625 = pi0384 & ~w6412;
assign w6626 = ~w6624 & ~w6625;
assign w6627 = pi1042 & w6412;
assign w6628 = pi0385 & ~w6412;
assign w6629 = ~w6627 & ~w6628;
assign w6630 = pi1059 & w6412;
assign w6631 = pi0386 & ~w6412;
assign w6632 = ~w6630 & ~w6631;
assign w6633 = pi1053 & w6412;
assign w6634 = pi0387 & ~w6412;
assign w6635 = ~w6633 & ~w6634;
assign w6636 = pi1037 & w6412;
assign w6637 = pi0388 & ~w6412;
assign w6638 = ~w6636 & ~w6637;
assign w6639 = pi1036 & w6412;
assign w6640 = pi0389 & ~w6412;
assign w6641 = ~w6639 & ~w6640;
assign w6642 = pi1049 & w6416;
assign w6643 = pi0390 & ~w6416;
assign w6644 = ~w6642 & ~w6643;
assign w6645 = pi1062 & w6416;
assign w6646 = pi0391 & ~w6416;
assign w6647 = ~w6645 & ~w6646;
assign w6648 = pi1039 & w6416;
assign w6649 = pi0392 & ~w6416;
assign w6650 = ~w6648 & ~w6649;
assign w6651 = pi1067 & w6416;
assign w6652 = pi0393 & ~w6416;
assign w6653 = ~w6651 & ~w6652;
assign w6654 = pi1080 & w6416;
assign w6655 = pi0394 & ~w6416;
assign w6656 = ~w6654 & ~w6655;
assign w6657 = pi1055 & w6416;
assign w6658 = pi0395 & ~w6416;
assign w6659 = ~w6657 & ~w6658;
assign w6660 = pi1051 & w6416;
assign w6661 = pi0396 & ~w6416;
assign w6662 = ~w6660 & ~w6661;
assign w6663 = pi1048 & w6416;
assign w6664 = pi0397 & ~w6416;
assign w6665 = ~w6663 & ~w6664;
assign w6666 = pi1087 & w6416;
assign w6667 = pi0398 & ~w6416;
assign w6668 = ~w6666 & ~w6667;
assign w6669 = pi1047 & w6416;
assign w6670 = pi0399 & ~w6416;
assign w6671 = ~w6669 & ~w6670;
assign w6672 = pi1035 & w6416;
assign w6673 = pi0400 & ~w6416;
assign w6674 = ~w6672 & ~w6673;
assign w6675 = pi1079 & w6416;
assign w6676 = pi0401 & ~w6416;
assign w6677 = ~w6675 & ~w6676;
assign w6678 = pi1078 & w6416;
assign w6679 = pi0402 & ~w6416;
assign w6680 = ~w6678 & ~w6679;
assign w6681 = pi1045 & w6416;
assign w6682 = pi0403 & ~w6416;
assign w6683 = ~w6681 & ~w6682;
assign w6684 = pi1084 & w6416;
assign w6685 = pi0404 & ~w6416;
assign w6686 = ~w6684 & ~w6685;
assign w6687 = pi1081 & w6416;
assign w6688 = pi0405 & ~w6416;
assign w6689 = ~w6687 & ~w6688;
assign w6690 = pi1076 & w6416;
assign w6691 = pi0406 & ~w6416;
assign w6692 = ~w6690 & ~w6691;
assign w6693 = pi1071 & w6416;
assign w6694 = pi0407 & ~w6416;
assign w6695 = ~w6693 & ~w6694;
assign w6696 = pi1068 & w6416;
assign w6697 = pi0408 & ~w6416;
assign w6698 = ~w6696 & ~w6697;
assign w6699 = pi1042 & w6416;
assign w6700 = pi0409 & ~w6416;
assign w6701 = ~w6699 & ~w6700;
assign w6702 = pi1059 & w6416;
assign w6703 = pi0410 & ~w6416;
assign w6704 = ~w6702 & ~w6703;
assign w6705 = pi1053 & w6416;
assign w6706 = pi0411 & ~w6416;
assign w6707 = ~w6705 & ~w6706;
assign w6708 = pi1037 & w6416;
assign w6709 = pi0412 & ~w6416;
assign w6710 = ~w6708 & ~w6709;
assign w6711 = pi1036 & w6416;
assign w6712 = pi0413 & ~w6416;
assign w6713 = ~w6711 & ~w6712;
assign w6714 = pi1049 & w6489;
assign w6715 = pi0414 & ~w6489;
assign w6716 = ~w6714 & ~w6715;
assign w6717 = pi1062 & w6489;
assign w6718 = pi0415 & ~w6489;
assign w6719 = ~w6717 & ~w6718;
assign w6720 = pi1069 & w6489;
assign w6721 = pi0416 & ~w6489;
assign w6722 = ~w6720 & ~w6721;
assign w6723 = pi1039 & w6489;
assign w6724 = pi0417 & ~w6489;
assign w6725 = ~w6723 & ~w6724;
assign w6726 = pi1067 & w6489;
assign w6727 = pi0418 & ~w6489;
assign w6728 = ~w6726 & ~w6727;
assign w6729 = pi1080 & w6489;
assign w6730 = pi0419 & ~w6489;
assign w6731 = ~w6729 & ~w6730;
assign w6732 = pi1055 & w6489;
assign w6733 = pi0420 & ~w6489;
assign w6734 = ~w6732 & ~w6733;
assign w6735 = pi1051 & w6489;
assign w6736 = pi0421 & ~w6489;
assign w6737 = ~w6735 & ~w6736;
assign w6738 = pi1048 & w6489;
assign w6739 = pi0422 & ~w6489;
assign w6740 = ~w6738 & ~w6739;
assign w6741 = pi1087 & w6489;
assign w6742 = pi0423 & ~w6489;
assign w6743 = ~w6741 & ~w6742;
assign w6744 = pi1047 & w6489;
assign w6745 = pi0424 & ~w6489;
assign w6746 = ~w6744 & ~w6745;
assign w6747 = pi1035 & w6489;
assign w6748 = pi0425 & ~w6489;
assign w6749 = ~w6747 & ~w6748;
assign w6750 = pi1079 & w6489;
assign w6751 = pi0426 & ~w6489;
assign w6752 = ~w6750 & ~w6751;
assign w6753 = pi1078 & w6489;
assign w6754 = pi0427 & ~w6489;
assign w6755 = ~w6753 & ~w6754;
assign w6756 = pi1045 & w6489;
assign w6757 = pi0428 & ~w6489;
assign w6758 = ~w6756 & ~w6757;
assign w6759 = pi1084 & w6489;
assign w6760 = pi0429 & ~w6489;
assign w6761 = ~w6759 & ~w6760;
assign w6762 = pi1076 & w6489;
assign w6763 = pi0430 & ~w6489;
assign w6764 = ~w6762 & ~w6763;
assign w6765 = pi1071 & w6489;
assign w6766 = pi0431 & ~w6489;
assign w6767 = ~w6765 & ~w6766;
assign w6768 = pi1068 & w6489;
assign w6769 = pi0432 & ~w6489;
assign w6770 = ~w6768 & ~w6769;
assign w6771 = pi1042 & w6489;
assign w6772 = pi0433 & ~w6489;
assign w6773 = ~w6771 & ~w6772;
assign w6774 = pi1059 & w6489;
assign w6775 = pi0434 & ~w6489;
assign w6776 = ~w6774 & ~w6775;
assign w6777 = pi1053 & w6489;
assign w6778 = pi0435 & ~w6489;
assign w6779 = ~w6777 & ~w6778;
assign w6780 = pi1037 & w6489;
assign w6781 = pi0436 & ~w6489;
assign w6782 = ~w6780 & ~w6781;
assign w6783 = pi1070 & w6489;
assign w6784 = pi0437 & ~w6489;
assign w6785 = ~w6783 & ~w6784;
assign w6786 = pi1036 & w6489;
assign w6787 = pi0438 & ~w6489;
assign w6788 = ~w6786 & ~w6787;
assign w6789 = pi1057 & w6412;
assign w6790 = pi0439 & ~w6412;
assign w6791 = ~w6789 & ~w6790;
assign w6792 = pi1043 & w6412;
assign w6793 = pi0440 & ~w6412;
assign w6794 = ~w6792 & ~w6793;
assign w6795 = pi1044 & w6405;
assign w6796 = pi0441 & ~w6405;
assign w6797 = ~w6795 & ~w6796;
assign w6798 = pi1058 & w6412;
assign w6799 = pi0442 & ~w6412;
assign w6800 = ~w6798 & ~w6799;
assign w6801 = pi1044 & w6489;
assign w6802 = pi0443 & ~w6489;
assign w6803 = ~w6801 & ~w6802;
assign w6804 = pi1072 & w6489;
assign w6805 = pi0444 & ~w6489;
assign w6806 = ~w6804 & ~w6805;
assign w6807 = pi1081 & w6489;
assign w6808 = pi0445 & ~w6489;
assign w6809 = ~w6807 & ~w6808;
assign w6810 = pi1086 & w6489;
assign w6811 = pi0446 & ~w6489;
assign w6812 = ~w6810 & ~w6811;
assign w6813 = pi1040 & w6412;
assign w6814 = pi0447 & ~w6412;
assign w6815 = ~w6813 & ~w6814;
assign w6816 = pi1074 & w6489;
assign w6817 = pi0448 & ~w6489;
assign w6818 = ~w6816 & ~w6817;
assign w6819 = pi1057 & w6489;
assign w6820 = pi0449 & ~w6489;
assign w6821 = ~w6819 & ~w6820;
assign w6822 = pi1036 & w6405;
assign w6823 = pi0450 & ~w6405;
assign w6824 = ~w6822 & ~w6823;
assign w6825 = pi1063 & w6489;
assign w6826 = pi0451 & ~w6489;
assign w6827 = ~w6825 & ~w6826;
assign w6828 = pi1053 & w6405;
assign w6829 = pi0452 & ~w6405;
assign w6830 = ~w6828 & ~w6829;
assign w6831 = pi1040 & w6489;
assign w6832 = pi0453 & ~w6489;
assign w6833 = ~w6831 & ~w6832;
assign w6834 = pi1043 & w6489;
assign w6835 = pi0454 & ~w6489;
assign w6836 = ~w6834 & ~w6835;
assign w6837 = pi1037 & w6405;
assign w6838 = pi0455 & ~w6405;
assign w6839 = ~w6837 & ~w6838;
assign w6840 = pi1044 & w6416;
assign w6841 = pi0456 & ~w6416;
assign w6842 = ~w6840 & ~w6841;
assign w6843 = pi0600 & ~pi0810;
assign w6844 = pi0804 & ~w6843;
assign w6845 = pi0601 & ~w6844;
assign w6846 = ~pi0804 & ~pi0810;
assign w6847 = ~w6845 & ~w6846;
assign w6848 = ~pi0815 & ~w6847;
assign w6849 = pi0599 & pi0815;
assign w6850 = pi0810 & ~w6849;
assign w6851 = pi0596 & ~w6850;
assign w6852 = pi0804 & ~w6851;
assign w6853 = pi0595 & ~w6852;
assign w6854 = ~w6846 & ~w6853;
assign w6855 = pi0594 & pi0597;
assign w6856 = pi0600 & w6855;
assign w6857 = pi0601 & w6856;
assign w6858 = ~w6854 & w6857;
assign w6859 = ~w6848 & ~w6858;
assign w6860 = pi0605 & ~w6859;
assign w6861 = pi0594 & pi0600;
assign w6862 = pi0804 & w6861;
assign w6863 = pi0810 & w6862;
assign w6864 = ~pi0815 & w6863;
assign w6865 = pi0990 & w6864;
assign w6866 = ~w6860 & ~w6865;
assign w6867 = pi0821 & ~w6866;
assign w6868 = pi1072 & w6405;
assign w6869 = pi0458 & ~w6405;
assign w6870 = ~w6868 & ~w6869;
assign w6871 = pi1058 & w6489;
assign w6872 = pi0459 & ~w6489;
assign w6873 = ~w6871 & ~w6872;
assign w6874 = pi1086 & w6405;
assign w6875 = pi0460 & ~w6405;
assign w6876 = ~w6874 & ~w6875;
assign w6877 = pi1057 & w6405;
assign w6878 = pi0461 & ~w6405;
assign w6879 = ~w6877 & ~w6878;
assign w6880 = pi1074 & w6405;
assign w6881 = pi0462 & ~w6405;
assign w6882 = ~w6880 & ~w6881;
assign w6883 = pi1070 & w6416;
assign w6884 = pi0463 & ~w6416;
assign w6885 = ~w6883 & ~w6884;
assign w6886 = pi1065 & w6489;
assign w6887 = pi0464 & ~w6489;
assign w6888 = ~w6886 & ~w6887;
assign w6889 = pi0926 & ~w6349;
assign w6890 = ~pi0243 & ~w6340;
assign w6891 = ~w6889 & ~w6890;
assign w6892 = pi1157 & w1225;
assign w6893 = w6891 & ~w6892;
assign w6894 = pi0943 & ~w6349;
assign w6895 = pi0275 & ~w6340;
assign w6896 = ~w6894 & ~w6895;
assign w6897 = pi1151 & w1225;
assign w6898 = w6896 & ~w6897;
assign w6899 = w3017 & w5356;
assign w6900 = pi0040 & ~w1284;
assign w6901 = ~pi0287 & w6900;
assign w6902 = ~pi0979 & w6901;
assign w6903 = ~pi0984 & w6902;
assign w6904 = pi1001 & w6903;
assign w6905 = ~w6899 & ~w6904;
assign w6906 = ~pi0024 & w1615;
assign w6907 = pi0468 & ~w6906;
assign w6908 = ~w3376 & ~w6907;
assign w6909 = pi0942 & ~w6349;
assign w6910 = ~pi0263 & ~w6340;
assign w6911 = ~w6909 & ~w6910;
assign w6912 = pi1156 & w1225;
assign w6913 = w6911 & ~w6912;
assign w6914 = pi0925 & ~w6349;
assign w6915 = pi0267 & ~w6340;
assign w6916 = ~w6914 & ~w6915;
assign w6917 = pi1155 & w1225;
assign w6918 = w6916 & ~w6917;
assign w6919 = pi0941 & ~w6349;
assign w6920 = pi0253 & ~w6340;
assign w6921 = ~w6919 & ~w6920;
assign w6922 = pi1153 & w1225;
assign w6923 = w6921 & ~w6922;
assign w6924 = pi0923 & ~w6349;
assign w6925 = pi0254 & ~w6340;
assign w6926 = ~w6924 & ~w6925;
assign w6927 = pi1154 & w1225;
assign w6928 = w6926 & ~w6927;
assign w6929 = pi0922 & ~w6349;
assign w6930 = pi0268 & ~w6340;
assign w6931 = ~w6929 & ~w6930;
assign w6932 = pi1152 & w1225;
assign w6933 = w6931 & ~w6932;
assign w6934 = pi0931 & ~w6349;
assign w6935 = pi0272 & ~w6340;
assign w6936 = ~w6934 & ~w6935;
assign w6937 = pi1150 & w1225;
assign w6938 = w6936 & ~w6937;
assign w6939 = pi0936 & ~w6349;
assign w6940 = pi0283 & ~w6340;
assign w6941 = ~w6939 & ~w6940;
assign w6942 = pi1149 & w1225;
assign w6943 = w6941 & ~w6942;
assign w6944 = pi0071 & ~w5785;
assign w6945 = ~w3705 & ~w6944;
assign w6946 = w2568 & ~w3879;
assign w6947 = ~w3848 & ~w3872;
assign w6948 = ~w6946 & ~w6947;
assign w6949 = pi0071 & ~w5774;
assign w6950 = pi0481 & ~w5145;
assign w6951 = pi0248 & w5145;
assign w6952 = ~w6950 & ~w6951;
assign w6953 = pi0482 & ~w5159;
assign w6954 = pi0249 & w5159;
assign w6955 = ~w6953 & ~w6954;
assign w6956 = pi0483 & ~w5188;
assign w6957 = pi0242 & w5188;
assign w6958 = ~w6956 & ~w6957;
assign w6959 = pi0484 & ~w5188;
assign w6960 = pi0249 & w5188;
assign w6961 = ~w6959 & ~w6960;
assign w6962 = pi0485 & ~w5258;
assign w6963 = pi0234 & w5258;
assign w6964 = ~w6962 & ~w6963;
assign w6965 = pi0486 & ~w5258;
assign w6966 = pi0244 & w5258;
assign w6967 = ~w6965 & ~w6966;
assign w6968 = pi0487 & ~w5145;
assign w6969 = pi0246 & w5145;
assign w6970 = ~w6968 & ~w6969;
assign w6971 = ~pi0488 & ~w5145;
assign w6972 = pi0239 & w5145;
assign w6973 = ~w6971 & ~w6972;
assign w6974 = pi0489 & ~w5258;
assign w6975 = pi0242 & w5258;
assign w6976 = ~w6974 & ~w6975;
assign w6977 = pi0490 & ~w5188;
assign w6978 = pi0241 & w5188;
assign w6979 = ~w6977 & ~w6978;
assign w6980 = pi0491 & ~w5188;
assign w6981 = pi0238 & w5188;
assign w6982 = ~w6980 & ~w6981;
assign w6983 = pi0492 & ~w5188;
assign w6984 = pi0240 & w5188;
assign w6985 = ~w6983 & ~w6984;
assign w6986 = pi0493 & ~w5188;
assign w6987 = pi0244 & w5188;
assign w6988 = ~w6986 & ~w6987;
assign w6989 = ~pi0494 & ~w5188;
assign w6990 = pi0239 & w5188;
assign w6991 = ~w6989 & ~w6990;
assign w6992 = pi0495 & ~w5188;
assign w6993 = pi0235 & w5188;
assign w6994 = ~w6992 & ~w6993;
assign w6995 = pi0496 & ~w5181;
assign w6996 = pi0249 & w5181;
assign w6997 = ~w6995 & ~w6996;
assign w6998 = ~pi0497 & ~w5181;
assign w6999 = pi0239 & w5181;
assign w7000 = ~w6998 & ~w6999;
assign w7001 = pi0498 & ~w5159;
assign w7002 = pi0238 & w5159;
assign w7003 = ~w7001 & ~w7002;
assign w7004 = pi0499 & ~w5181;
assign w7005 = pi0246 & w5181;
assign w7006 = ~w7004 & ~w7005;
assign w7007 = pi0500 & ~w5181;
assign w7008 = pi0241 & w5181;
assign w7009 = ~w7007 & ~w7008;
assign w7010 = pi0501 & ~w5181;
assign w7011 = pi0248 & w5181;
assign w7012 = ~w7010 & ~w7011;
assign w7013 = pi0502 & ~w5181;
assign w7014 = pi0247 & w5181;
assign w7015 = ~w7013 & ~w7014;
assign w7016 = pi0503 & ~w5181;
assign w7017 = pi0245 & w5181;
assign w7018 = ~w7016 & ~w7017;
assign w7019 = pi0504 & ~w5177;
assign w7020 = pi0242 & w5177;
assign w7021 = ~w7019 & ~w7020;
assign w7022 = pi0505 & ~w5181;
assign w7023 = pi0234 & w5181;
assign w7024 = ~w7022 & ~w7023;
assign w7025 = pi0506 & ~w5177;
assign w7026 = pi0241 & w5177;
assign w7027 = ~w7025 & ~w7026;
assign w7028 = pi0507 & ~w5177;
assign w7029 = pi0238 & w5177;
assign w7030 = ~w7028 & ~w7029;
assign w7031 = pi0508 & ~w5177;
assign w7032 = pi0247 & w5177;
assign w7033 = ~w7031 & ~w7032;
assign w7034 = pi0509 & ~w5177;
assign w7035 = pi0245 & w5177;
assign w7036 = ~w7034 & ~w7035;
assign w7037 = pi0510 & ~w5145;
assign w7038 = pi0242 & w5145;
assign w7039 = ~w7037 & ~w7038;
assign w7040 = pi0511 & ~w5145;
assign w7041 = pi0234 & w5145;
assign w7042 = ~w7040 & ~w7041;
assign w7043 = pi0512 & ~w5145;
assign w7044 = pi0235 & w5145;
assign w7045 = ~w7043 & ~w7044;
assign w7046 = pi0513 & ~w5145;
assign w7047 = pi0244 & w5145;
assign w7048 = ~w7046 & ~w7047;
assign w7049 = pi0514 & ~w5145;
assign w7050 = pi0245 & w5145;
assign w7051 = ~w7049 & ~w7050;
assign w7052 = pi0515 & ~w5145;
assign w7053 = pi0240 & w5145;
assign w7054 = ~w7052 & ~w7053;
assign w7055 = pi0516 & ~w5145;
assign w7056 = pi0247 & w5145;
assign w7057 = ~w7055 & ~w7056;
assign w7058 = pi0517 & ~w5145;
assign w7059 = pi0238 & w5145;
assign w7060 = ~w7058 & ~w7059;
assign w7061 = pi0518 & ~w5152;
assign w7062 = pi0234 & w5152;
assign w7063 = ~w7061 & ~w7062;
assign w7064 = ~pi0519 & ~w5152;
assign w7065 = pi0239 & w5152;
assign w7066 = ~w7064 & ~w7065;
assign w7067 = pi0520 & ~w5152;
assign w7068 = pi0246 & w5152;
assign w7069 = ~w7067 & ~w7068;
assign w7070 = pi0521 & ~w5152;
assign w7071 = pi0248 & w5152;
assign w7072 = ~w7070 & ~w7071;
assign w7073 = pi0522 & ~w5152;
assign w7074 = pi0238 & w5152;
assign w7075 = ~w7073 & ~w7074;
assign w7076 = pi0523 & ~w5268;
assign w7077 = pi0234 & w5268;
assign w7078 = ~w7076 & ~w7077;
assign w7079 = ~pi0524 & ~w5268;
assign w7080 = pi0239 & w5268;
assign w7081 = ~w7079 & ~w7080;
assign w7082 = pi0525 & ~w5268;
assign w7083 = pi0245 & w5268;
assign w7084 = ~w7082 & ~w7083;
assign w7085 = pi0526 & ~w5268;
assign w7086 = pi0246 & w5268;
assign w7087 = ~w7085 & ~w7086;
assign w7088 = pi0527 & ~w5268;
assign w7089 = pi0247 & w5268;
assign w7090 = ~w7088 & ~w7089;
assign w7091 = pi0528 & ~w5268;
assign w7092 = pi0249 & w5268;
assign w7093 = ~w7091 & ~w7092;
assign w7094 = pi0529 & ~w5268;
assign w7095 = pi0238 & w5268;
assign w7096 = ~w7094 & ~w7095;
assign w7097 = pi0530 & ~w5268;
assign w7098 = pi0240 & w5268;
assign w7099 = ~w7097 & ~w7098;
assign w7100 = pi0531 & ~w5159;
assign w7101 = pi0235 & w5159;
assign w7102 = ~w7100 & ~w7101;
assign w7103 = pi0532 & ~w5159;
assign w7104 = pi0247 & w5159;
assign w7105 = ~w7103 & ~w7104;
assign w7106 = pi0533 & ~w5177;
assign w7107 = pi0235 & w5177;
assign w7108 = ~w7106 & ~w7107;
assign w7109 = ~pi0534 & ~w5177;
assign w7110 = pi0239 & w5177;
assign w7111 = ~w7109 & ~w7110;
assign w7112 = pi0535 & ~w5177;
assign w7113 = pi0240 & w5177;
assign w7114 = ~w7112 & ~w7113;
assign w7115 = pi0536 & ~w5177;
assign w7116 = pi0246 & w5177;
assign w7117 = ~w7115 & ~w7116;
assign w7118 = pi0537 & ~w5177;
assign w7119 = pi0248 & w5177;
assign w7120 = ~w7118 & ~w7119;
assign w7121 = pi0538 & ~w5177;
assign w7122 = pi0249 & w5177;
assign w7123 = ~w7121 & ~w7122;
assign w7124 = pi0539 & ~w5181;
assign w7125 = pi0242 & w5181;
assign w7126 = ~w7124 & ~w7125;
assign w7127 = pi0540 & ~w5181;
assign w7128 = pi0235 & w5181;
assign w7129 = ~w7127 & ~w7128;
assign w7130 = pi0541 & ~w5181;
assign w7131 = pi0244 & w5181;
assign w7132 = ~w7130 & ~w7131;
assign w7133 = pi0542 & ~w5181;
assign w7134 = pi0240 & w5181;
assign w7135 = ~w7133 & ~w7134;
assign w7136 = pi0543 & ~w5181;
assign w7137 = pi0238 & w5181;
assign w7138 = ~w7136 & ~w7137;
assign w7139 = pi0544 & ~w5188;
assign w7140 = pi0234 & w5188;
assign w7141 = ~w7139 & ~w7140;
assign w7142 = pi0545 & ~w5188;
assign w7143 = pi0245 & w5188;
assign w7144 = ~w7142 & ~w7143;
assign w7145 = pi0546 & ~w5188;
assign w7146 = pi0246 & w5188;
assign w7147 = ~w7145 & ~w7146;
assign w7148 = pi0547 & ~w5188;
assign w7149 = pi0247 & w5188;
assign w7150 = ~w7148 & ~w7149;
assign w7151 = pi0548 & ~w5188;
assign w7152 = pi0248 & w5188;
assign w7153 = ~w7151 & ~w7152;
assign w7154 = pi0549 & ~w5258;
assign w7155 = pi0235 & w5258;
assign w7156 = ~w7154 & ~w7155;
assign w7157 = ~pi0550 & ~w5258;
assign w7158 = pi0239 & w5258;
assign w7159 = ~w7157 & ~w7158;
assign w7160 = pi0551 & ~w5258;
assign w7161 = pi0240 & w5258;
assign w7162 = ~w7160 & ~w7161;
assign w7163 = pi0552 & ~w5258;
assign w7164 = pi0247 & w5258;
assign w7165 = ~w7163 & ~w7164;
assign w7166 = pi0553 & ~w5258;
assign w7167 = pi0241 & w5258;
assign w7168 = ~w7166 & ~w7167;
assign w7169 = pi0554 & ~w5258;
assign w7170 = pi0248 & w5258;
assign w7171 = ~w7169 & ~w7170;
assign w7172 = pi0555 & ~w5258;
assign w7173 = pi0249 & w5258;
assign w7174 = ~w7172 & ~w7173;
assign w7175 = pi0556 & ~w5159;
assign w7176 = pi0242 & w5159;
assign w7177 = ~w7175 & ~w7176;
assign w7178 = pi0557 & ~w5177;
assign w7179 = pi0234 & w5177;
assign w7180 = ~w7178 & ~w7179;
assign w7181 = pi0558 & ~w5177;
assign w7182 = pi0244 & w5177;
assign w7183 = ~w7181 & ~w7182;
assign w7184 = pi0559 & ~w5145;
assign w7185 = pi0241 & w5145;
assign w7186 = ~w7184 & ~w7185;
assign w7187 = pi0560 & ~w5159;
assign w7188 = pi0240 & w5159;
assign w7189 = ~w7187 & ~w7188;
assign w7190 = pi0561 & ~w5152;
assign w7191 = pi0247 & w5152;
assign w7192 = ~w7190 & ~w7191;
assign w7193 = pi0562 & ~w5159;
assign w7194 = pi0241 & w5159;
assign w7195 = ~w7193 & ~w7194;
assign w7196 = pi0563 & ~w5258;
assign w7197 = pi0246 & w5258;
assign w7198 = ~w7196 & ~w7197;
assign w7199 = pi0564 & ~w5159;
assign w7200 = pi0246 & w5159;
assign w7201 = ~w7199 & ~w7200;
assign w7202 = pi0565 & ~w5159;
assign w7203 = pi0248 & w5159;
assign w7204 = ~w7202 & ~w7203;
assign w7205 = pi0566 & ~w5159;
assign w7206 = pi0244 & w5159;
assign w7207 = ~w7205 & ~w7206;
assign w7208 = pi0621 & w4673;
assign w7209 = pi0665 & w4631;
assign w7210 = ~w7208 & ~w7209;
assign w7211 = pi1091 & ~w7210;
assign w7212 = pi0230 & pi1093;
assign w7213 = w7211 & w7212;
assign w7214 = ~pi0567 & ~w7212;
assign w7215 = ~w7213 & ~w7214;
assign w7216 = pi1092 & ~w7215;
assign w7217 = pi0568 & ~w5159;
assign w7218 = pi0245 & w5159;
assign w7219 = ~w7217 & ~w7218;
assign w7220 = ~pi0569 & ~w5159;
assign w7221 = pi0239 & w5159;
assign w7222 = ~w7220 & ~w7221;
assign w7223 = pi0570 & ~w5159;
assign w7224 = pi0234 & w5159;
assign w7225 = ~w7223 & ~w7224;
assign w7226 = pi0571 & ~w5268;
assign w7227 = pi0241 & w5268;
assign w7228 = ~w7226 & ~w7227;
assign w7229 = pi0572 & ~w5268;
assign w7230 = pi0244 & w5268;
assign w7231 = ~w7229 & ~w7230;
assign w7232 = pi0573 & ~w5268;
assign w7233 = pi0242 & w5268;
assign w7234 = ~w7232 & ~w7233;
assign w7235 = pi0574 & ~w5152;
assign w7236 = pi0241 & w5152;
assign w7237 = ~w7235 & ~w7236;
assign w7238 = pi0575 & ~w5268;
assign w7239 = pi0235 & w5268;
assign w7240 = ~w7238 & ~w7239;
assign w7241 = pi0576 & ~w5268;
assign w7242 = pi0248 & w5268;
assign w7243 = ~w7241 & ~w7242;
assign w7244 = pi0577 & ~w5258;
assign w7245 = pi0238 & w5258;
assign w7246 = ~w7244 & ~w7245;
assign w7247 = pi0578 & ~w5152;
assign w7248 = pi0249 & w5152;
assign w7249 = ~w7247 & ~w7248;
assign w7250 = pi0579 & ~w5145;
assign w7251 = pi0249 & w5145;
assign w7252 = ~w7250 & ~w7251;
assign w7253 = pi0580 & ~w5258;
assign w7254 = pi0245 & w5258;
assign w7255 = ~w7253 & ~w7254;
assign w7256 = pi0581 & ~w5152;
assign w7257 = pi0235 & w5152;
assign w7258 = ~w7256 & ~w7257;
assign w7259 = pi0582 & ~w5152;
assign w7260 = pi0240 & w5152;
assign w7261 = ~w7259 & ~w7260;
assign w7262 = pi0584 & ~w5152;
assign w7263 = pi0245 & w5152;
assign w7264 = ~w7262 & ~w7263;
assign w7265 = pi0585 & ~w5152;
assign w7266 = pi0244 & w5152;
assign w7267 = ~w7265 & ~w7266;
assign w7268 = pi0586 & ~w5152;
assign w7269 = pi0242 & w5152;
assign w7270 = ~w7268 & ~w7269;
assign w7271 = ~pi0230 & pi0587;
assign w7272 = pi0230 & w4674;
assign w7273 = ~w7271 & ~w7272;
assign w7274 = ~pi0123 & pi0824;
assign w7275 = pi0950 & w7274;
assign w7276 = pi0591 & w7275;
assign w7277 = pi0588 & ~w7275;
assign w7278 = ~w7276 & ~w7277;
assign w7279 = ~w1234 & ~w7278;
assign w7280 = pi1092 & w7279;
assign w7281 = ~pi0203 & ~pi0237;
assign w7282 = ~pi0202 & pi0237;
assign w7283 = ~w7281 & ~w7282;
assign w7284 = ~pi0233 & ~w7283;
assign w7285 = ~pi0201 & pi0237;
assign w7286 = ~pi0220 & ~pi0237;
assign w7287 = ~w7285 & ~w7286;
assign w7288 = pi0233 & ~w7287;
assign w7289 = ~w7284 & ~w7288;
assign w7290 = ~w5142 & ~w7289;
assign w7291 = ~pi0205 & pi0237;
assign w7292 = ~pi0218 & ~pi0237;
assign w7293 = ~w7291 & ~w7292;
assign w7294 = ~pi0233 & ~w7293;
assign w7295 = ~pi0206 & ~pi0237;
assign w7296 = ~pi0204 & pi0237;
assign w7297 = ~w7295 & ~w7296;
assign w7298 = pi0233 & ~w7297;
assign w7299 = ~w7294 & ~w7298;
assign w7300 = ~w5174 & ~w7299;
assign w7301 = ~w7290 & ~w7300;
assign w7302 = pi0588 & w7275;
assign w7303 = ~w1234 & ~w7302;
assign w7304 = pi0590 & ~w7275;
assign w7305 = pi1092 & ~w7304;
assign w7306 = w7303 & w7305;
assign w7307 = pi0592 & w7275;
assign w7308 = pi0591 & ~w7275;
assign w7309 = ~w7307 & ~w7308;
assign w7310 = ~w1234 & ~w7309;
assign w7311 = pi1092 & w7310;
assign w7312 = pi0592 & ~w7275;
assign w7313 = pi0590 & w7275;
assign w7314 = ~w7312 & ~w7313;
assign w7315 = ~w1234 & ~w7314;
assign w7316 = pi1092 & w7315;
assign w7317 = pi0234 & pi0485;
assign w7318 = ~pi0234 & ~pi0485;
assign w7319 = ~w7317 & ~w7318;
assign w7320 = ~pi0233 & ~w7319;
assign w7321 = ~pi0249 & ~pi0555;
assign w7322 = pi0249 & pi0555;
assign w7323 = ~w7321 & ~w7322;
assign w7324 = ~pi0248 & ~pi0554;
assign w7325 = pi0248 & pi0554;
assign w7326 = ~w7324 & ~w7325;
assign w7327 = ~w7323 & ~w7326;
assign w7328 = pi0241 & pi0553;
assign w7329 = ~pi0241 & ~pi0553;
assign w7330 = ~w7328 & ~w7329;
assign w7331 = pi0242 & pi0489;
assign w7332 = ~pi0242 & ~pi0489;
assign w7333 = ~w7331 & ~w7332;
assign w7334 = ~w7330 & ~w7333;
assign w7335 = w7327 & w7334;
assign w7336 = w7320 & w7335;
assign w7337 = ~pi0245 & ~pi0580;
assign w7338 = pi0245 & pi0580;
assign w7339 = ~w7337 & ~w7338;
assign w7340 = pi0247 & pi0552;
assign w7341 = ~pi0247 & ~pi0552;
assign w7342 = ~w7340 & ~w7341;
assign w7343 = ~w7339 & ~w7342;
assign w7344 = pi0238 & pi0577;
assign w7345 = ~pi0238 & ~pi0577;
assign w7346 = ~w7344 & ~w7345;
assign w7347 = pi0246 & pi0563;
assign w7348 = ~pi0246 & ~pi0563;
assign w7349 = ~w7347 & ~w7348;
assign w7350 = ~w7346 & ~w7349;
assign w7351 = w7343 & w7350;
assign w7352 = pi0239 & ~pi0550;
assign w7353 = ~pi0239 & pi0550;
assign w7354 = ~w7352 & ~w7353;
assign w7355 = ~pi0244 & ~pi0486;
assign w7356 = pi0244 & pi0486;
assign w7357 = ~w7355 & ~w7356;
assign w7358 = ~w7354 & ~w7357;
assign w7359 = pi0235 & pi0549;
assign w7360 = ~pi0235 & ~pi0549;
assign w7361 = ~w7359 & ~w7360;
assign w7362 = ~pi0240 & ~pi0551;
assign w7363 = pi0240 & pi0551;
assign w7364 = ~w7362 & ~w7363;
assign w7365 = ~w7361 & ~w7364;
assign w7366 = w7358 & w7365;
assign w7367 = w7351 & w7366;
assign w7368 = w7336 & w7367;
assign w7369 = pi0238 & pi0491;
assign w7370 = ~pi0238 & ~pi0491;
assign w7371 = ~w7369 & ~w7370;
assign w7372 = pi0233 & ~w7371;
assign w7373 = ~pi0246 & ~pi0546;
assign w7374 = pi0246 & pi0546;
assign w7375 = ~w7373 & ~w7374;
assign w7376 = ~pi0239 & pi0494;
assign w7377 = pi0239 & ~pi0494;
assign w7378 = ~w7376 & ~w7377;
assign w7379 = ~w7375 & ~w7378;
assign w7380 = pi0244 & pi0493;
assign w7381 = ~pi0244 & ~pi0493;
assign w7382 = ~w7380 & ~w7381;
assign w7383 = pi0249 & pi0484;
assign w7384 = ~pi0249 & ~pi0484;
assign w7385 = ~w7383 & ~w7384;
assign w7386 = ~w7382 & ~w7385;
assign w7387 = w7379 & w7386;
assign w7388 = w7372 & w7387;
assign w7389 = pi0245 & pi0545;
assign w7390 = ~pi0245 & ~pi0545;
assign w7391 = ~w7389 & ~w7390;
assign w7392 = ~pi0234 & ~pi0544;
assign w7393 = pi0234 & pi0544;
assign w7394 = ~w7392 & ~w7393;
assign w7395 = ~w7391 & ~w7394;
assign w7396 = pi0247 & pi0547;
assign w7397 = ~pi0247 & ~pi0547;
assign w7398 = ~w7396 & ~w7397;
assign w7399 = ~pi0248 & ~pi0548;
assign w7400 = pi0248 & pi0548;
assign w7401 = ~w7399 & ~w7400;
assign w7402 = ~w7398 & ~w7401;
assign w7403 = w7395 & w7402;
assign w7404 = ~pi0235 & ~pi0495;
assign w7405 = pi0235 & pi0495;
assign w7406 = ~w7404 & ~w7405;
assign w7407 = ~pi0242 & ~pi0483;
assign w7408 = pi0242 & pi0483;
assign w7409 = ~w7407 & ~w7408;
assign w7410 = ~w7406 & ~w7409;
assign w7411 = pi0240 & pi0492;
assign w7412 = ~pi0240 & ~pi0492;
assign w7413 = ~w7411 & ~w7412;
assign w7414 = pi0241 & pi0490;
assign w7415 = ~pi0241 & ~pi0490;
assign w7416 = ~w7414 & ~w7415;
assign w7417 = ~w7413 & ~w7416;
assign w7418 = w7410 & w7417;
assign w7419 = w7403 & w7418;
assign w7420 = w7388 & w7419;
assign w7421 = ~w7368 & ~w7420;
assign w7422 = ~pi0237 & ~w7421;
assign w7423 = pi0245 & pi0509;
assign w7424 = ~pi0245 & ~pi0509;
assign w7425 = ~w7423 & ~w7424;
assign w7426 = pi0233 & ~w7425;
assign w7427 = ~pi0248 & ~pi0537;
assign w7428 = pi0248 & pi0537;
assign w7429 = ~w7427 & ~w7428;
assign w7430 = ~pi0239 & pi0534;
assign w7431 = pi0239 & ~pi0534;
assign w7432 = ~w7430 & ~w7431;
assign w7433 = ~w7429 & ~w7432;
assign w7434 = pi0238 & pi0507;
assign w7435 = ~pi0238 & ~pi0507;
assign w7436 = ~w7434 & ~w7435;
assign w7437 = ~pi0246 & ~pi0536;
assign w7438 = pi0246 & pi0536;
assign w7439 = ~w7437 & ~w7438;
assign w7440 = ~w7436 & ~w7439;
assign w7441 = w7433 & w7440;
assign w7442 = w7426 & w7441;
assign w7443 = pi0249 & pi0538;
assign w7444 = ~pi0249 & ~pi0538;
assign w7445 = ~w7443 & ~w7444;
assign w7446 = ~pi0247 & ~pi0508;
assign w7447 = pi0247 & pi0508;
assign w7448 = ~w7446 & ~w7447;
assign w7449 = ~w7445 & ~w7448;
assign w7450 = pi0234 & pi0557;
assign w7451 = ~pi0234 & ~pi0557;
assign w7452 = ~w7450 & ~w7451;
assign w7453 = ~pi0244 & ~pi0558;
assign w7454 = pi0244 & pi0558;
assign w7455 = ~w7453 & ~w7454;
assign w7456 = ~w7452 & ~w7455;
assign w7457 = w7449 & w7456;
assign w7458 = ~pi0240 & ~pi0535;
assign w7459 = pi0240 & pi0535;
assign w7460 = ~w7458 & ~w7459;
assign w7461 = ~pi0241 & ~pi0506;
assign w7462 = pi0241 & pi0506;
assign w7463 = ~w7461 & ~w7462;
assign w7464 = ~w7460 & ~w7463;
assign w7465 = pi0235 & pi0533;
assign w7466 = ~pi0235 & ~pi0533;
assign w7467 = ~w7465 & ~w7466;
assign w7468 = pi0242 & pi0504;
assign w7469 = ~pi0242 & ~pi0504;
assign w7470 = ~w7468 & ~w7469;
assign w7471 = ~w7467 & ~w7470;
assign w7472 = w7464 & w7471;
assign w7473 = w7457 & w7472;
assign w7474 = w7442 & w7473;
assign w7475 = pi0247 & pi0502;
assign w7476 = ~pi0247 & ~pi0502;
assign w7477 = ~w7475 & ~w7476;
assign w7478 = ~pi0233 & ~w7477;
assign w7479 = ~pi0235 & ~pi0540;
assign w7480 = pi0235 & pi0540;
assign w7481 = ~w7479 & ~w7480;
assign w7482 = ~pi0245 & ~pi0503;
assign w7483 = pi0245 & pi0503;
assign w7484 = ~w7482 & ~w7483;
assign w7485 = ~w7481 & ~w7484;
assign w7486 = pi0238 & pi0543;
assign w7487 = ~pi0238 & ~pi0543;
assign w7488 = ~w7486 & ~w7487;
assign w7489 = pi0249 & pi0496;
assign w7490 = ~pi0249 & ~pi0496;
assign w7491 = ~w7489 & ~w7490;
assign w7492 = ~w7488 & ~w7491;
assign w7493 = w7485 & w7492;
assign w7494 = w7478 & w7493;
assign w7495 = ~pi0244 & ~pi0541;
assign w7496 = pi0244 & pi0541;
assign w7497 = ~w7495 & ~w7496;
assign w7498 = pi0248 & pi0501;
assign w7499 = ~pi0248 & ~pi0501;
assign w7500 = ~w7498 & ~w7499;
assign w7501 = ~w7497 & ~w7500;
assign w7502 = pi0240 & pi0542;
assign w7503 = ~pi0240 & ~pi0542;
assign w7504 = ~w7502 & ~w7503;
assign w7505 = pi0242 & pi0539;
assign w7506 = ~pi0242 & ~pi0539;
assign w7507 = ~w7505 & ~w7506;
assign w7508 = ~w7504 & ~w7507;
assign w7509 = w7501 & w7508;
assign w7510 = ~pi0246 & ~pi0499;
assign w7511 = pi0246 & pi0499;
assign w7512 = ~w7510 & ~w7511;
assign w7513 = ~pi0239 & pi0497;
assign w7514 = pi0239 & ~pi0497;
assign w7515 = ~w7513 & ~w7514;
assign w7516 = ~w7512 & ~w7515;
assign w7517 = pi0234 & pi0505;
assign w7518 = ~pi0234 & ~pi0505;
assign w7519 = ~w7517 & ~w7518;
assign w7520 = pi0241 & pi0500;
assign w7521 = ~pi0241 & ~pi0500;
assign w7522 = ~w7520 & ~w7521;
assign w7523 = ~w7519 & ~w7522;
assign w7524 = w7516 & w7523;
assign w7525 = w7509 & w7524;
assign w7526 = w7494 & w7525;
assign w7527 = ~w7474 & ~w7526;
assign w7528 = pi0237 & ~w7527;
assign w7529 = ~w7422 & ~w7528;
assign w7530 = ~w5174 & ~w7529;
assign w7531 = pi0246 & pi0526;
assign w7532 = ~pi0246 & ~pi0526;
assign w7533 = ~w7531 & ~w7532;
assign w7534 = pi0233 & ~w7533;
assign w7535 = ~pi0235 & ~pi0575;
assign w7536 = pi0235 & pi0575;
assign w7537 = ~w7535 & ~w7536;
assign w7538 = ~pi0240 & ~pi0530;
assign w7539 = pi0240 & pi0530;
assign w7540 = ~w7538 & ~w7539;
assign w7541 = ~w7537 & ~w7540;
assign w7542 = pi0247 & pi0527;
assign w7543 = ~pi0247 & ~pi0527;
assign w7544 = ~w7542 & ~w7543;
assign w7545 = ~pi0249 & ~pi0528;
assign w7546 = pi0249 & pi0528;
assign w7547 = ~w7545 & ~w7546;
assign w7548 = ~w7544 & ~w7547;
assign w7549 = w7541 & w7548;
assign w7550 = w7534 & w7549;
assign w7551 = pi0242 & pi0573;
assign w7552 = ~pi0242 & ~pi0573;
assign w7553 = ~w7551 & ~w7552;
assign w7554 = ~pi0241 & ~pi0571;
assign w7555 = pi0241 & pi0571;
assign w7556 = ~w7554 & ~w7555;
assign w7557 = ~w7553 & ~w7556;
assign w7558 = pi0244 & pi0572;
assign w7559 = ~pi0244 & ~pi0572;
assign w7560 = ~w7558 & ~w7559;
assign w7561 = ~pi0248 & ~pi0576;
assign w7562 = pi0248 & pi0576;
assign w7563 = ~w7561 & ~w7562;
assign w7564 = ~w7560 & ~w7563;
assign w7565 = w7557 & w7564;
assign w7566 = ~pi0234 & ~pi0523;
assign w7567 = pi0234 & pi0523;
assign w7568 = ~w7566 & ~w7567;
assign w7569 = pi0239 & ~pi0524;
assign w7570 = ~pi0239 & pi0524;
assign w7571 = ~w7569 & ~w7570;
assign w7572 = ~w7568 & ~w7571;
assign w7573 = pi0238 & pi0529;
assign w7574 = ~pi0238 & ~pi0529;
assign w7575 = ~w7573 & ~w7574;
assign w7576 = pi0245 & pi0525;
assign w7577 = ~pi0245 & ~pi0525;
assign w7578 = ~w7576 & ~w7577;
assign w7579 = ~w7575 & ~w7578;
assign w7580 = w7572 & w7579;
assign w7581 = w7565 & w7580;
assign w7582 = w7550 & w7581;
assign w7583 = ~pi0237 & ~w7582;
assign w7584 = pi0249 & pi0482;
assign w7585 = ~pi0249 & ~pi0482;
assign w7586 = ~w7584 & ~w7585;
assign w7587 = ~pi0233 & ~w7586;
assign w7588 = pi0239 & ~pi0569;
assign w7589 = ~pi0239 & pi0569;
assign w7590 = ~w7588 & ~w7589;
assign w7591 = ~pi0241 & ~pi0562;
assign w7592 = pi0241 & pi0562;
assign w7593 = ~w7591 & ~w7592;
assign w7594 = ~w7590 & ~w7593;
assign w7595 = pi0240 & pi0560;
assign w7596 = ~pi0240 & ~pi0560;
assign w7597 = ~w7595 & ~w7596;
assign w7598 = pi0242 & pi0556;
assign w7599 = ~pi0242 & ~pi0556;
assign w7600 = ~w7598 & ~w7599;
assign w7601 = ~w7597 & ~w7600;
assign w7602 = w7594 & w7601;
assign w7603 = w7587 & w7602;
assign w7604 = ~pi0245 & ~pi0568;
assign w7605 = pi0245 & pi0568;
assign w7606 = ~w7604 & ~w7605;
assign w7607 = pi0246 & pi0564;
assign w7608 = ~pi0246 & ~pi0564;
assign w7609 = ~w7607 & ~w7608;
assign w7610 = ~w7606 & ~w7609;
assign w7611 = pi0234 & pi0570;
assign w7612 = ~pi0234 & ~pi0570;
assign w7613 = ~w7611 & ~w7612;
assign w7614 = pi0248 & pi0565;
assign w7615 = ~pi0248 & ~pi0565;
assign w7616 = ~w7614 & ~w7615;
assign w7617 = ~w7613 & ~w7616;
assign w7618 = w7610 & w7617;
assign w7619 = ~pi0244 & ~pi0566;
assign w7620 = pi0244 & pi0566;
assign w7621 = ~w7619 & ~w7620;
assign w7622 = ~pi0238 & ~pi0498;
assign w7623 = pi0238 & pi0498;
assign w7624 = ~w7622 & ~w7623;
assign w7625 = ~w7621 & ~w7624;
assign w7626 = pi0235 & pi0531;
assign w7627 = ~pi0235 & ~pi0531;
assign w7628 = ~w7626 & ~w7627;
assign w7629 = ~pi0247 & ~pi0532;
assign w7630 = pi0247 & pi0532;
assign w7631 = ~w7629 & ~w7630;
assign w7632 = ~w7628 & ~w7631;
assign w7633 = w7625 & w7632;
assign w7634 = w7618 & w7633;
assign w7635 = w7603 & w7634;
assign w7636 = w7583 & ~w7635;
assign w7637 = pi0246 & pi0520;
assign w7638 = ~pi0246 & ~pi0520;
assign w7639 = ~w7637 & ~w7638;
assign w7640 = ~pi0233 & ~w7639;
assign w7641 = ~pi0244 & ~pi0585;
assign w7642 = pi0244 & pi0585;
assign w7643 = ~w7641 & ~w7642;
assign w7644 = ~pi0240 & ~pi0582;
assign w7645 = pi0240 & pi0582;
assign w7646 = ~w7644 & ~w7645;
assign w7647 = ~w7643 & ~w7646;
assign w7648 = ~pi0247 & ~pi0561;
assign w7649 = pi0247 & pi0561;
assign w7650 = ~w7648 & ~w7649;
assign w7651 = pi0239 & ~pi0519;
assign w7652 = ~pi0239 & pi0519;
assign w7653 = ~w7651 & ~w7652;
assign w7654 = ~w7650 & ~w7653;
assign w7655 = w7647 & w7654;
assign w7656 = w7640 & w7655;
assign w7657 = ~pi0245 & ~pi0584;
assign w7658 = pi0245 & pi0584;
assign w7659 = ~w7657 & ~w7658;
assign w7660 = pi0249 & pi0578;
assign w7661 = ~pi0249 & ~pi0578;
assign w7662 = ~w7660 & ~w7661;
assign w7663 = ~w7659 & ~w7662;
assign w7664 = pi0235 & pi0581;
assign w7665 = ~pi0235 & ~pi0581;
assign w7666 = ~w7664 & ~w7665;
assign w7667 = ~pi0242 & ~pi0586;
assign w7668 = pi0242 & pi0586;
assign w7669 = ~w7667 & ~w7668;
assign w7670 = ~w7666 & ~w7669;
assign w7671 = w7663 & w7670;
assign w7672 = ~pi0238 & ~pi0522;
assign w7673 = pi0238 & pi0522;
assign w7674 = ~w7672 & ~w7673;
assign w7675 = ~pi0234 & ~pi0518;
assign w7676 = pi0234 & pi0518;
assign w7677 = ~w7675 & ~w7676;
assign w7678 = ~w7674 & ~w7677;
assign w7679 = pi0241 & pi0574;
assign w7680 = ~pi0241 & ~pi0574;
assign w7681 = ~w7679 & ~w7680;
assign w7682 = pi0248 & pi0521;
assign w7683 = ~pi0248 & ~pi0521;
assign w7684 = ~w7682 & ~w7683;
assign w7685 = ~w7681 & ~w7684;
assign w7686 = w7678 & w7685;
assign w7687 = w7671 & w7686;
assign w7688 = w7656 & w7687;
assign w7689 = pi0237 & ~w7688;
assign w7690 = pi0242 & pi0510;
assign w7691 = ~pi0242 & ~pi0510;
assign w7692 = ~w7690 & ~w7691;
assign w7693 = pi0233 & ~w7692;
assign w7694 = ~pi0241 & ~pi0559;
assign w7695 = pi0241 & pi0559;
assign w7696 = ~w7694 & ~w7695;
assign w7697 = ~pi0235 & ~pi0512;
assign w7698 = pi0235 & pi0512;
assign w7699 = ~w7697 & ~w7698;
assign w7700 = ~w7696 & ~w7699;
assign w7701 = pi0246 & pi0487;
assign w7702 = ~pi0246 & ~pi0487;
assign w7703 = ~w7701 & ~w7702;
assign w7704 = ~pi0247 & ~pi0516;
assign w7705 = pi0247 & pi0516;
assign w7706 = ~w7704 & ~w7705;
assign w7707 = ~w7703 & ~w7706;
assign w7708 = w7700 & w7707;
assign w7709 = w7693 & w7708;
assign w7710 = ~pi0238 & ~pi0517;
assign w7711 = pi0238 & pi0517;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = pi0245 & pi0514;
assign w7714 = ~pi0245 & ~pi0514;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = ~w7712 & ~w7715;
assign w7717 = pi0240 & pi0515;
assign w7718 = ~pi0240 & ~pi0515;
assign w7719 = ~w7717 & ~w7718;
assign w7720 = ~pi0249 & ~pi0579;
assign w7721 = pi0249 & pi0579;
assign w7722 = ~w7720 & ~w7721;
assign w7723 = ~w7719 & ~w7722;
assign w7724 = w7716 & w7723;
assign w7725 = ~pi0244 & ~pi0513;
assign w7726 = pi0244 & pi0513;
assign w7727 = ~w7725 & ~w7726;
assign w7728 = ~pi0248 & ~pi0481;
assign w7729 = pi0248 & pi0481;
assign w7730 = ~w7728 & ~w7729;
assign w7731 = ~w7727 & ~w7730;
assign w7732 = pi0234 & pi0511;
assign w7733 = ~pi0234 & ~pi0511;
assign w7734 = ~w7732 & ~w7733;
assign w7735 = pi0239 & ~pi0488;
assign w7736 = ~pi0239 & pi0488;
assign w7737 = ~w7735 & ~w7736;
assign w7738 = ~w7734 & ~w7737;
assign w7739 = w7731 & w7738;
assign w7740 = w7724 & w7739;
assign w7741 = w7709 & w7740;
assign w7742 = w7689 & ~w7741;
assign w7743 = ~w7636 & ~w7742;
assign w7744 = ~w5142 & w7743;
assign w7745 = ~w7530 & ~w7744;
assign w7746 = ~pi0806 & pi0990;
assign w7747 = pi0600 & w7746;
assign w7748 = pi0594 & ~w7747;
assign w7749 = ~pi0594 & pi0990;
assign w7750 = pi0600 & ~pi0806;
assign w7751 = w7749 & w7750;
assign w7752 = ~w7748 & ~w7751;
assign w7753 = ~pi0332 & ~w7752;
assign w7754 = ~pi0595 & ~pi0806;
assign w7755 = pi0605 & w6857;
assign w7756 = w7754 & w7755;
assign w7757 = pi0605 & ~pi0806;
assign w7758 = w6857 & w7757;
assign w7759 = pi0595 & ~w7758;
assign w7760 = ~w7756 & ~w7759;
assign w7761 = ~pi0332 & ~w7760;
assign w7762 = pi0594 & pi0595;
assign w7763 = pi0597 & w7762;
assign w7764 = pi0600 & w7763;
assign w7765 = ~pi0806 & w7764;
assign w7766 = pi0990 & w7765;
assign w7767 = ~pi0596 & w7766;
assign w7768 = pi0596 & ~w7766;
assign w7769 = ~w7767 & ~w7768;
assign w7770 = ~pi0332 & ~w7769;
assign w7771 = ~pi0597 & pi0990;
assign w7772 = ~pi0806 & w7771;
assign w7773 = w6861 & w7772;
assign w7774 = w6861 & w7746;
assign w7775 = pi0597 & ~w7774;
assign w7776 = ~w7773 & ~w7775;
assign w7777 = ~pi0332 & ~w7776;
assign w7778 = ~pi0882 & w529;
assign w7779 = pi0947 & w7778;
assign w7780 = pi0598 & ~w7779;
assign w7781 = pi0740 & pi0780;
assign w7782 = w1249 & w7781;
assign w7783 = ~w7780 & ~w7782;
assign w7784 = pi0596 & ~pi0599;
assign w7785 = w7766 & w7784;
assign w7786 = pi0596 & w7766;
assign w7787 = pi0599 & ~w7786;
assign w7788 = ~w7785 & ~w7787;
assign w7789 = ~pi0332 & ~w7788;
assign w7790 = ~pi0600 & pi0990;
assign w7791 = ~pi0806 & w7790;
assign w7792 = pi0600 & ~w7746;
assign w7793 = ~w7791 & ~w7792;
assign w7794 = ~pi0332 & ~w7793;
assign w7795 = ~pi0806 & pi0989;
assign w7796 = pi0601 & pi0806;
assign w7797 = ~w7795 & ~w7796;
assign w7798 = ~pi0332 & ~w7797;
assign w7799 = ~pi0230 & pi0602;
assign w7800 = pi0230 & w4632;
assign w7801 = ~w7799 & ~w7800;
assign w7802 = ~pi0872 & pi0966;
assign w7803 = ~pi0871 & w7802;
assign w7804 = pi0832 & pi0952;
assign w7805 = ~pi0980 & w7804;
assign w7806 = pi1038 & w7805;
assign w7807 = pi1060 & w7806;
assign w7808 = ~pi1061 & w7807;
assign w7809 = ~pi1100 & w7808;
assign w7810 = ~pi0603 & ~w7808;
assign w7811 = ~w7809 & ~w7810;
assign w7812 = ~pi0966 & ~w7811;
assign w7813 = ~w7803 & ~w7812;
assign w7814 = pi0907 & pi0983;
assign w7815 = ~pi0299 & w7814;
assign w7816 = pi0604 & ~w7815;
assign w7817 = ~pi0681 & w1251;
assign w7818 = pi0823 & w7817;
assign w7819 = ~w7816 & ~w7818;
assign w7820 = pi0779 & w7818;
assign w7821 = ~w7819 & ~w7820;
assign w7822 = pi0605 & pi0806;
assign w7823 = ~pi0605 & ~pi0806;
assign w7824 = ~w7822 & ~w7823;
assign w7825 = ~pi0332 & ~w7824;
assign w7826 = pi0606 & ~w7808;
assign w7827 = pi1104 & w7808;
assign w7828 = ~w7826 & ~w7827;
assign w7829 = ~pi0966 & ~w7828;
assign w7830 = pi0837 & pi0966;
assign w7831 = ~w7829 & ~w7830;
assign w7832 = pi0607 & ~w7808;
assign w7833 = pi1107 & w7808;
assign w7834 = ~w7832 & ~w7833;
assign w7835 = ~pi0966 & ~w7834;
assign w7836 = pi0608 & ~w7808;
assign w7837 = pi1116 & w7808;
assign w7838 = ~w7836 & ~w7837;
assign w7839 = ~pi0966 & ~w7838;
assign w7840 = pi0609 & ~w7808;
assign w7841 = pi1118 & w7808;
assign w7842 = ~w7840 & ~w7841;
assign w7843 = ~pi0966 & ~w7842;
assign w7844 = pi0610 & ~w7808;
assign w7845 = pi1113 & w7808;
assign w7846 = ~w7844 & ~w7845;
assign w7847 = ~pi0966 & ~w7846;
assign w7848 = pi0611 & ~w7808;
assign w7849 = pi1114 & w7808;
assign w7850 = ~w7848 & ~w7849;
assign w7851 = ~pi0966 & ~w7850;
assign w7852 = pi0612 & ~w7808;
assign w7853 = pi1111 & w7808;
assign w7854 = ~w7852 & ~w7853;
assign w7855 = ~pi0966 & ~w7854;
assign w7856 = pi0613 & ~w7808;
assign w7857 = pi1115 & w7808;
assign w7858 = ~w7856 & ~w7857;
assign w7859 = ~pi0966 & ~w7858;
assign w7860 = pi0614 & ~w7808;
assign w7861 = pi1102 & w7808;
assign w7862 = ~w7860 & ~w7861;
assign w7863 = ~pi0966 & ~w7862;
assign w7864 = pi0871 & pi0966;
assign w7865 = ~w7863 & ~w7864;
assign w7866 = pi0907 & w7778;
assign w7867 = ~pi0615 & ~w7866;
assign w7868 = pi0779 & pi0797;
assign w7869 = w1253 & w7868;
assign w7870 = ~w7867 & ~w7869;
assign w7871 = pi0616 & ~w7808;
assign w7872 = pi1101 & w7808;
assign w7873 = ~w7871 & ~w7872;
assign w7874 = ~pi0966 & ~w7873;
assign w7875 = pi0872 & pi0966;
assign w7876 = ~w7874 & ~w7875;
assign w7877 = pi0617 & ~w7808;
assign w7878 = pi1105 & w7808;
assign w7879 = ~w7877 & ~w7878;
assign w7880 = ~pi0966 & ~w7879;
assign w7881 = pi0850 & pi0966;
assign w7882 = ~w7880 & ~w7881;
assign w7883 = pi0618 & ~w7808;
assign w7884 = pi1117 & w7808;
assign w7885 = ~w7883 & ~w7884;
assign w7886 = ~pi0966 & ~w7885;
assign w7887 = pi0619 & ~w7808;
assign w7888 = pi1122 & w7808;
assign w7889 = ~w7887 & ~w7888;
assign w7890 = ~pi0966 & ~w7889;
assign w7891 = pi0620 & ~w7808;
assign w7892 = pi1112 & w7808;
assign w7893 = ~w7891 & ~w7892;
assign w7894 = ~pi0966 & ~w7893;
assign w7895 = pi0621 & ~w7808;
assign w7896 = pi1108 & w7808;
assign w7897 = ~w7895 & ~w7896;
assign w7898 = ~pi0966 & ~w7897;
assign w7899 = pi0622 & ~w7808;
assign w7900 = pi1109 & w7808;
assign w7901 = ~w7899 & ~w7900;
assign w7902 = ~pi0966 & ~w7901;
assign w7903 = pi0623 & ~w7808;
assign w7904 = pi1106 & w7808;
assign w7905 = ~w7903 & ~w7904;
assign w7906 = ~pi0966 & ~w7905;
assign w7907 = pi0947 & pi0983;
assign w7908 = ~pi0299 & w7907;
assign w7909 = pi0624 & ~w7908;
assign w7910 = ~pi0614 & ~pi0616;
assign w7911 = ~pi0642 & w7910;
assign w7912 = pi0831 & w7911;
assign w7913 = ~w7909 & ~w7912;
assign w7914 = pi0780 & w7912;
assign w7915 = ~w7913 & ~w7914;
assign w7916 = pi0832 & ~pi0953;
assign w7917 = ~pi0973 & w7916;
assign w7918 = ~pi1054 & w7917;
assign w7919 = pi1066 & w7918;
assign w7920 = pi1088 & w7919;
assign w7921 = pi0625 & ~w7920;
assign w7922 = pi1116 & w7920;
assign w7923 = ~w7921 & ~w7922;
assign w7924 = ~pi0962 & ~w7923;
assign w7925 = pi0626 & ~w7808;
assign w7926 = pi1121 & w7808;
assign w7927 = ~w7925 & ~w7926;
assign w7928 = ~pi0966 & ~w7927;
assign w7929 = pi0627 & ~w7920;
assign w7930 = pi1117 & w7920;
assign w7931 = ~w7929 & ~w7930;
assign w7932 = ~pi0962 & ~w7931;
assign w7933 = pi0628 & ~w7920;
assign w7934 = pi1119 & w7920;
assign w7935 = ~w7933 & ~w7934;
assign w7936 = ~pi0962 & ~w7935;
assign w7937 = pi0629 & ~w7808;
assign w7938 = pi1119 & w7808;
assign w7939 = ~w7937 & ~w7938;
assign w7940 = ~pi0966 & ~w7939;
assign w7941 = pi0630 & ~w7808;
assign w7942 = pi1120 & w7808;
assign w7943 = ~w7941 & ~w7942;
assign w7944 = ~pi0966 & ~w7943;
assign w7945 = ~pi0631 & ~w7920;
assign w7946 = pi1113 & w7920;
assign w7947 = ~w7945 & ~w7946;
assign w7948 = ~pi0962 & ~w7947;
assign w7949 = ~pi0632 & ~w7920;
assign w7950 = pi1115 & w7920;
assign w7951 = ~w7949 & ~w7950;
assign w7952 = ~pi0962 & ~w7951;
assign w7953 = pi0633 & ~w7808;
assign w7954 = pi1110 & w7808;
assign w7955 = ~w7953 & ~w7954;
assign w7956 = ~pi0966 & ~w7955;
assign w7957 = pi0634 & ~w7920;
assign w7958 = pi1110 & w7920;
assign w7959 = ~w7957 & ~w7958;
assign w7960 = ~pi0962 & ~w7959;
assign w7961 = ~pi0635 & ~w7920;
assign w7962 = pi1112 & w7920;
assign w7963 = ~w7961 & ~w7962;
assign w7964 = ~pi0962 & ~w7963;
assign w7965 = pi0636 & ~w7808;
assign w7966 = pi1127 & w7808;
assign w7967 = ~w7965 & ~w7966;
assign w7968 = ~pi0966 & ~w7967;
assign w7969 = pi0637 & ~w7920;
assign w7970 = pi1105 & w7920;
assign w7971 = ~w7969 & ~w7970;
assign w7972 = ~pi0962 & ~w7971;
assign w7973 = pi0638 & ~w7920;
assign w7974 = pi1107 & w7920;
assign w7975 = ~w7973 & ~w7974;
assign w7976 = ~pi0962 & ~w7975;
assign w7977 = pi0639 & ~w7920;
assign w7978 = pi1109 & w7920;
assign w7979 = ~w7977 & ~w7978;
assign w7980 = ~pi0962 & ~w7979;
assign w7981 = pi0640 & ~w7808;
assign w7982 = pi1128 & w7808;
assign w7983 = ~w7981 & ~w7982;
assign w7984 = ~pi0966 & ~w7983;
assign w7985 = pi0641 & ~w7920;
assign w7986 = pi1121 & w7920;
assign w7987 = ~w7985 & ~w7986;
assign w7988 = ~pi0962 & ~w7987;
assign w7989 = pi0642 & ~w7808;
assign w7990 = pi1103 & w7808;
assign w7991 = ~w7989 & ~w7990;
assign w7992 = ~pi0966 & ~w7991;
assign w7993 = pi0643 & ~w7920;
assign w7994 = pi1104 & w7920;
assign w7995 = ~w7993 & ~w7994;
assign w7996 = ~pi0962 & ~w7995;
assign w7997 = pi0644 & ~w7808;
assign w7998 = pi1123 & w7808;
assign w7999 = ~w7997 & ~w7998;
assign w8000 = ~pi0966 & ~w7999;
assign w8001 = pi0645 & ~w7808;
assign w8002 = pi1125 & w7808;
assign w8003 = ~w8001 & ~w8002;
assign w8004 = ~pi0966 & ~w8003;
assign w8005 = ~pi0646 & ~w7920;
assign w8006 = pi1114 & w7920;
assign w8007 = ~w8005 & ~w8006;
assign w8008 = ~pi0962 & ~w8007;
assign w8009 = pi0647 & ~w7920;
assign w8010 = pi1120 & w7920;
assign w8011 = ~w8009 & ~w8010;
assign w8012 = ~pi0962 & ~w8011;
assign w8013 = pi0648 & ~w7920;
assign w8014 = pi1122 & w7920;
assign w8015 = ~w8013 & ~w8014;
assign w8016 = ~pi0962 & ~w8015;
assign w8017 = ~pi0649 & ~w7920;
assign w8018 = pi1126 & w7920;
assign w8019 = ~w8017 & ~w8018;
assign w8020 = ~pi0962 & ~w8019;
assign w8021 = ~pi0650 & ~w7920;
assign w8022 = pi1127 & w7920;
assign w8023 = ~w8021 & ~w8022;
assign w8024 = ~pi0962 & ~w8023;
assign w8025 = pi0651 & ~w7808;
assign w8026 = pi1130 & w7808;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = ~pi0966 & ~w8027;
assign w8029 = pi0652 & ~w7808;
assign w8030 = pi1131 & w7808;
assign w8031 = ~w8029 & ~w8030;
assign w8032 = ~pi0966 & ~w8031;
assign w8033 = pi0653 & ~w7808;
assign w8034 = pi1129 & w7808;
assign w8035 = ~w8033 & ~w8034;
assign w8036 = ~pi0966 & ~w8035;
assign w8037 = ~pi0654 & ~w7920;
assign w8038 = pi1130 & w7920;
assign w8039 = ~w8037 & ~w8038;
assign w8040 = ~pi0962 & ~w8039;
assign w8041 = ~pi0655 & ~w7920;
assign w8042 = pi1124 & w7920;
assign w8043 = ~w8041 & ~w8042;
assign w8044 = ~pi0962 & ~w8043;
assign w8045 = pi0656 & ~w7808;
assign w8046 = pi1126 & w7808;
assign w8047 = ~w8045 & ~w8046;
assign w8048 = ~pi0966 & ~w8047;
assign w8049 = ~pi0657 & ~w7920;
assign w8050 = pi1131 & w7920;
assign w8051 = ~w8049 & ~w8050;
assign w8052 = ~pi0962 & ~w8051;
assign w8053 = pi0658 & ~w7808;
assign w8054 = pi1124 & w7808;
assign w8055 = ~w8053 & ~w8054;
assign w8056 = ~pi0966 & ~w8055;
assign w8057 = pi0274 & ~pi0277;
assign w8058 = ~pi0270 & w8057;
assign w8059 = ~pi0264 & ~pi0265;
assign w8060 = pi0266 & ~pi0269;
assign w8061 = ~pi0280 & w8060;
assign w8062 = ~pi0281 & w8061;
assign w8063 = ~pi0282 & w8062;
assign w8064 = pi0992 & w8063;
assign w8065 = w8059 & w8064;
assign w8066 = w8058 & w8065;
assign w8067 = ~pi0270 & ~pi0277;
assign w8068 = ~pi0265 & w8067;
assign w8069 = ~pi0264 & w8064;
assign w8070 = w8068 & w8069;
assign w8071 = ~pi0274 & ~w8070;
assign w8072 = ~w8066 & ~w8071;
assign w8073 = pi0660 & ~w7920;
assign w8074 = pi1118 & w7920;
assign w8075 = ~w8073 & ~w8074;
assign w8076 = ~pi0962 & ~w8075;
assign w8077 = pi0661 & ~w7920;
assign w8078 = pi1101 & w7920;
assign w8079 = ~w8077 & ~w8078;
assign w8080 = ~pi0962 & ~w8079;
assign w8081 = pi0662 & ~w7920;
assign w8082 = pi1102 & w7920;
assign w8083 = ~w8081 & ~w8082;
assign w8084 = ~pi0962 & ~w8083;
assign w8085 = ~pi0815 & ~pi1136;
assign w8086 = ~pi0633 & pi1136;
assign w8087 = ~w8085 & ~w8086;
assign w8088 = ~pi1134 & ~w8087;
assign w8089 = ~pi0766 & pi1136;
assign w8090 = ~pi0855 & ~pi1136;
assign w8091 = ~w8089 & ~w8090;
assign w8092 = pi1134 & ~w8091;
assign w8093 = ~w8088 & ~w8092;
assign w8094 = ~pi1135 & w8093;
assign w8095 = pi1134 & pi1136;
assign w8096 = pi0700 & w8095;
assign w8097 = pi0634 & pi1136;
assign w8098 = pi0784 & ~pi1136;
assign w8099 = ~w8097 & ~w8098;
assign w8100 = ~pi1134 & ~w8099;
assign w8101 = ~w8096 & ~w8100;
assign w8102 = pi1135 & ~w8101;
assign w8103 = ~w8094 & ~w8102;
assign w8104 = ~pi1137 & ~w2045;
assign w8105 = ~pi1138 & w8104;
assign w8106 = ~w8103 & w8105;
assign w8107 = ~pi0199 & pi0257;
assign w8108 = pi0199 & pi1065;
assign w8109 = ~w8107 & ~w8108;
assign w8110 = ~w4192 & ~w8109;
assign w8111 = ~pi0591 & w2409;
assign w8112 = pi0464 & ~pi0590;
assign w8113 = w8111 & w8112;
assign w8114 = pi0323 & pi0590;
assign w8115 = w1858 & w8114;
assign w8116 = ~pi0591 & pi0592;
assign w8117 = pi0365 & w8116;
assign w8118 = pi0591 & ~pi0592;
assign w8119 = pi0334 & w8118;
assign w8120 = ~w8117 & ~w8119;
assign w8121 = ~pi0590 & ~w8120;
assign w8122 = ~w8115 & ~w8121;
assign w8123 = ~pi0588 & ~w8122;
assign w8124 = ~w8113 & ~w8123;
assign w8125 = w4192 & ~w8124;
assign w8126 = ~w8110 & ~w8125;
assign w8127 = w2045 & ~w8126;
assign w8128 = ~w8106 & ~w8127;
assign w8129 = ~pi0811 & ~pi1136;
assign w8130 = ~pi0614 & pi1136;
assign w8131 = ~w8129 & ~w8130;
assign w8132 = ~pi1134 & ~w8131;
assign w8133 = ~pi0772 & pi1136;
assign w8134 = ~pi0872 & ~pi1136;
assign w8135 = ~w8133 & ~w8134;
assign w8136 = pi1134 & ~w8135;
assign w8137 = ~w8132 & ~w8136;
assign w8138 = ~pi1135 & w8137;
assign w8139 = pi0727 & w8095;
assign w8140 = pi0662 & pi1136;
assign w8141 = pi0785 & ~pi1136;
assign w8142 = ~w8140 & ~w8141;
assign w8143 = ~pi1134 & ~w8142;
assign w8144 = ~w8139 & ~w8143;
assign w8145 = pi1135 & ~w8144;
assign w8146 = ~w8138 & ~w8145;
assign w8147 = w8105 & ~w8146;
assign w8148 = ~pi0199 & pi0292;
assign w8149 = pi0199 & pi1084;
assign w8150 = ~w8148 & ~w8149;
assign w8151 = ~w4192 & ~w8150;
assign w8152 = pi0429 & ~pi0590;
assign w8153 = w8111 & w8152;
assign w8154 = pi0404 & w8118;
assign w8155 = pi0380 & w8116;
assign w8156 = ~w8154 & ~w8155;
assign w8157 = ~pi0590 & ~w8156;
assign w8158 = pi0355 & pi0590;
assign w8159 = w1858 & w8158;
assign w8160 = ~w8157 & ~w8159;
assign w8161 = ~pi0588 & ~w8160;
assign w8162 = ~w8153 & ~w8161;
assign w8163 = w4192 & ~w8162;
assign w8164 = ~w8151 & ~w8163;
assign w8165 = w2045 & ~w8164;
assign w8166 = ~w8147 & ~w8165;
assign w8167 = pi0665 & ~w7920;
assign w8168 = pi1108 & w7920;
assign w8169 = ~w8167 & ~w8168;
assign w8170 = ~pi0962 & ~w8169;
assign w8171 = ~pi0799 & ~pi1136;
assign w8172 = pi0607 & pi1136;
assign w8173 = ~w8171 & ~w8172;
assign w8174 = ~pi1134 & ~w8173;
assign w8175 = pi0764 & pi1136;
assign w8176 = pi0873 & ~pi1136;
assign w8177 = ~w8175 & ~w8176;
assign w8178 = pi1134 & ~w8177;
assign w8179 = ~w8174 & ~w8178;
assign w8180 = ~pi1135 & ~w8179;
assign w8181 = pi0691 & w8095;
assign w8182 = pi0638 & pi1136;
assign w8183 = pi0790 & ~pi1136;
assign w8184 = ~w8182 & ~w8183;
assign w8185 = ~pi1134 & ~w8184;
assign w8186 = ~w8181 & ~w8185;
assign w8187 = pi1135 & ~w8186;
assign w8188 = ~w8180 & ~w8187;
assign w8189 = w8105 & ~w8188;
assign w8190 = ~pi0199 & pi0297;
assign w8191 = pi0199 & pi1044;
assign w8192 = ~w8190 & ~w8191;
assign w8193 = ~w4192 & ~w8192;
assign w8194 = pi0443 & ~pi0590;
assign w8195 = w8111 & w8194;
assign w8196 = pi0441 & pi0590;
assign w8197 = w1858 & w8196;
assign w8198 = pi0337 & w8116;
assign w8199 = pi0456 & w8118;
assign w8200 = ~w8198 & ~w8199;
assign w8201 = ~pi0590 & ~w8200;
assign w8202 = ~w8197 & ~w8201;
assign w8203 = ~pi0588 & ~w8202;
assign w8204 = ~w8195 & ~w8203;
assign w8205 = w4192 & ~w8204;
assign w8206 = ~w8193 & ~w8205;
assign w8207 = w2045 & ~w8206;
assign w8208 = ~w8189 & ~w8207;
assign w8209 = ~pi0809 & ~pi1136;
assign w8210 = pi0642 & pi1136;
assign w8211 = ~w8209 & ~w8210;
assign w8212 = ~pi1134 & ~w8211;
assign w8213 = pi0763 & pi1136;
assign w8214 = pi0871 & ~pi1136;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = pi1134 & ~w8215;
assign w8217 = ~w8212 & ~w8216;
assign w8218 = ~pi1135 & ~w8217;
assign w8219 = pi0699 & w8095;
assign w8220 = pi0681 & pi1136;
assign w8221 = pi0792 & ~pi1136;
assign w8222 = ~w8220 & ~w8221;
assign w8223 = ~pi1134 & ~w8222;
assign w8224 = ~w8219 & ~w8223;
assign w8225 = pi1135 & ~w8224;
assign w8226 = ~w8218 & ~w8225;
assign w8227 = w8105 & ~w8226;
assign w8228 = ~pi0199 & pi0294;
assign w8229 = pi0199 & pi1072;
assign w8230 = ~w8228 & ~w8229;
assign w8231 = ~w4192 & ~w8230;
assign w8232 = pi0444 & ~pi0590;
assign w8233 = w8111 & w8232;
assign w8234 = pi0458 & pi0590;
assign w8235 = w1858 & w8234;
assign w8236 = pi0338 & w8116;
assign w8237 = pi0319 & w8118;
assign w8238 = ~w8236 & ~w8237;
assign w8239 = ~pi0590 & ~w8238;
assign w8240 = ~w8235 & ~w8239;
assign w8241 = ~pi0588 & ~w8240;
assign w8242 = ~w8233 & ~w8241;
assign w8243 = w4192 & ~w8242;
assign w8244 = ~w8231 & ~w8243;
assign w8245 = w2045 & ~w8244;
assign w8246 = ~w8227 & ~w8245;
assign w8247 = ~pi0603 & pi1136;
assign w8248 = ~pi0981 & ~pi1136;
assign w8249 = ~w8247 & ~w8248;
assign w8250 = ~pi1134 & ~w8249;
assign w8251 = ~pi0837 & ~pi1136;
assign w8252 = ~pi0759 & pi1136;
assign w8253 = ~w8251 & ~w8252;
assign w8254 = pi1134 & ~w8253;
assign w8255 = ~w8250 & ~w8254;
assign w8256 = ~pi1135 & w8255;
assign w8257 = pi0696 & w8095;
assign w8258 = pi0680 & pi1136;
assign w8259 = pi0778 & ~pi1136;
assign w8260 = ~w8258 & ~w8259;
assign w8261 = ~pi1134 & ~w8260;
assign w8262 = ~w8257 & ~w8261;
assign w8263 = pi1135 & ~w8262;
assign w8264 = ~w8256 & ~w8263;
assign w8265 = w8105 & ~w8264;
assign w8266 = ~pi0199 & pi0291;
assign w8267 = pi0199 & pi1049;
assign w8268 = ~w8266 & ~w8267;
assign w8269 = ~w4192 & ~w8268;
assign w8270 = pi0414 & ~pi0590;
assign w8271 = w8111 & w8270;
assign w8272 = pi0390 & w8118;
assign w8273 = pi0363 & w8116;
assign w8274 = ~w8272 & ~w8273;
assign w8275 = ~pi0590 & ~w8274;
assign w8276 = pi0342 & pi0590;
assign w8277 = w1858 & w8276;
assign w8278 = ~w8275 & ~w8277;
assign w8279 = ~pi0588 & ~w8278;
assign w8280 = ~w8271 & ~w8279;
assign w8281 = w4192 & ~w8280;
assign w8282 = ~w8269 & ~w8281;
assign w8283 = w2045 & ~w8282;
assign w8284 = ~w8265 & ~w8283;
assign w8285 = ~pi0669 & ~w7920;
assign w8286 = pi1125 & w7920;
assign w8287 = ~w8285 & ~w8286;
assign w8288 = ~pi0962 & ~w8287;
assign w8289 = pi0612 & ~pi1135;
assign w8290 = ~pi0695 & pi1135;
assign w8291 = ~w8289 & ~w8290;
assign w8292 = ~pi1134 & ~w8291;
assign w8293 = ~pi0723 & pi1135;
assign w8294 = ~pi0745 & ~pi1135;
assign w8295 = ~w8293 & ~w8294;
assign w8296 = pi1134 & ~w8295;
assign w8297 = ~w8292 & ~w8296;
assign w8298 = pi1136 & ~w8297;
assign w8299 = pi1134 & ~pi1135;
assign w8300 = ~pi1136 & w8299;
assign w8301 = pi0852 & w8300;
assign w8302 = ~w8298 & ~w8301;
assign w8303 = w8105 & ~w8302;
assign w8304 = ~pi0199 & pi0258;
assign w8305 = pi0199 & pi1062;
assign w8306 = ~w8304 & ~w8305;
assign w8307 = ~w4192 & ~w8306;
assign w8308 = pi0415 & ~pi0590;
assign w8309 = w8111 & w8308;
assign w8310 = pi0391 & w8118;
assign w8311 = pi0364 & w8116;
assign w8312 = ~w8310 & ~w8311;
assign w8313 = ~pi0590 & ~w8312;
assign w8314 = pi0343 & pi0590;
assign w8315 = w1858 & w8314;
assign w8316 = ~w8313 & ~w8315;
assign w8317 = ~pi0588 & ~w8316;
assign w8318 = ~w8309 & ~w8317;
assign w8319 = w4192 & ~w8318;
assign w8320 = ~w8307 & ~w8319;
assign w8321 = w2045 & ~w8320;
assign w8322 = ~w8303 & ~w8321;
assign w8323 = pi0865 & w8300;
assign w8324 = pi0611 & ~pi1135;
assign w8325 = ~pi0646 & pi1135;
assign w8326 = ~w8324 & ~w8325;
assign w8327 = ~pi1134 & ~w8326;
assign w8328 = ~pi0724 & pi1135;
assign w8329 = ~pi0741 & ~pi1135;
assign w8330 = ~w8328 & ~w8329;
assign w8331 = pi1134 & ~w8330;
assign w8332 = ~w8327 & ~w8331;
assign w8333 = pi1136 & ~w8332;
assign w8334 = ~w8323 & ~w8333;
assign w8335 = w8105 & ~w8334;
assign w8336 = ~pi0199 & pi0261;
assign w8337 = pi0199 & pi1040;
assign w8338 = ~w8336 & ~w8337;
assign w8339 = ~w4192 & ~w8338;
assign w8340 = pi0453 & ~pi0590;
assign w8341 = w8111 & w8340;
assign w8342 = pi0327 & pi0590;
assign w8343 = w1858 & w8342;
assign w8344 = pi0447 & w8116;
assign w8345 = pi0333 & w8118;
assign w8346 = ~w8344 & ~w8345;
assign w8347 = ~pi0590 & ~w8346;
assign w8348 = ~w8343 & ~w8347;
assign w8349 = ~pi0588 & ~w8348;
assign w8350 = ~w8341 & ~w8349;
assign w8351 = w4192 & ~w8350;
assign w8352 = ~w8339 & ~w8351;
assign w8353 = w2045 & ~w8352;
assign w8354 = ~w8335 & ~w8353;
assign w8355 = ~pi0808 & ~pi1136;
assign w8356 = ~pi0616 & pi1136;
assign w8357 = ~w8355 & ~w8356;
assign w8358 = ~pi1134 & ~w8357;
assign w8359 = ~pi0758 & pi1136;
assign w8360 = ~pi0850 & ~pi1136;
assign w8361 = ~w8359 & ~w8360;
assign w8362 = pi1134 & ~w8361;
assign w8363 = ~w8358 & ~w8362;
assign w8364 = ~pi1135 & w8363;
assign w8365 = pi0736 & w8095;
assign w8366 = pi0661 & pi1136;
assign w8367 = pi0781 & ~pi1136;
assign w8368 = ~w8366 & ~w8367;
assign w8369 = ~pi1134 & ~w8368;
assign w8370 = ~w8365 & ~w8369;
assign w8371 = pi1135 & ~w8370;
assign w8372 = ~w8364 & ~w8371;
assign w8373 = w8105 & ~w8372;
assign w8374 = ~pi0199 & pi0290;
assign w8375 = pi0199 & pi1048;
assign w8376 = ~w8374 & ~w8375;
assign w8377 = ~w4192 & ~w8376;
assign w8378 = pi0422 & ~pi0590;
assign w8379 = w8111 & w8378;
assign w8380 = pi0397 & w8118;
assign w8381 = pi0372 & w8116;
assign w8382 = ~w8380 & ~w8381;
assign w8383 = ~pi0590 & ~w8382;
assign w8384 = pi0320 & pi0590;
assign w8385 = w1858 & w8384;
assign w8386 = ~w8383 & ~w8385;
assign w8387 = ~pi0588 & ~w8386;
assign w8388 = ~w8379 & ~w8387;
assign w8389 = w4192 & ~w8388;
assign w8390 = ~w8377 & ~w8389;
assign w8391 = w2045 & ~w8390;
assign w8392 = ~w8373 & ~w8391;
assign w8393 = ~pi0814 & ~pi1136;
assign w8394 = pi0617 & pi1136;
assign w8395 = ~w8393 & ~w8394;
assign w8396 = ~pi1134 & ~w8395;
assign w8397 = pi0749 & pi1136;
assign w8398 = pi0866 & ~pi1136;
assign w8399 = ~w8397 & ~w8398;
assign w8400 = pi1134 & ~w8399;
assign w8401 = ~w8396 & ~w8400;
assign w8402 = ~pi1135 & ~w8401;
assign w8403 = pi0706 & w8095;
assign w8404 = pi0637 & pi1136;
assign w8405 = pi0788 & ~pi1136;
assign w8406 = ~w8404 & ~w8405;
assign w8407 = ~pi1134 & ~w8406;
assign w8408 = ~w8403 & ~w8407;
assign w8409 = pi1135 & ~w8408;
assign w8410 = ~w8402 & ~w8409;
assign w8411 = w8105 & ~w8410;
assign w8412 = ~pi0199 & pi0295;
assign w8413 = pi0199 & pi1053;
assign w8414 = ~w8412 & ~w8413;
assign w8415 = ~w4192 & ~w8414;
assign w8416 = pi0435 & ~pi0590;
assign w8417 = w8111 & w8416;
assign w8418 = pi0387 & w8116;
assign w8419 = pi0411 & w8118;
assign w8420 = ~w8418 & ~w8419;
assign w8421 = ~pi0590 & ~w8420;
assign w8422 = pi0452 & pi0590;
assign w8423 = w1858 & w8422;
assign w8424 = ~w8421 & ~w8423;
assign w8425 = ~pi0588 & ~w8424;
assign w8426 = ~w8417 & ~w8425;
assign w8427 = w4192 & ~w8426;
assign w8428 = ~w8415 & ~w8427;
assign w8429 = w2045 & ~w8428;
assign w8430 = ~w8411 & ~w8429;
assign w8431 = ~pi0804 & ~pi1136;
assign w8432 = ~pi0622 & pi1136;
assign w8433 = ~w8431 & ~w8432;
assign w8434 = ~pi1134 & ~w8433;
assign w8435 = ~pi0743 & pi1136;
assign w8436 = ~pi0859 & ~pi1136;
assign w8437 = ~w8435 & ~w8436;
assign w8438 = pi1134 & ~w8437;
assign w8439 = ~w8434 & ~w8438;
assign w8440 = ~pi1135 & w8439;
assign w8441 = pi0735 & w8095;
assign w8442 = pi0639 & pi1136;
assign w8443 = pi0783 & ~pi1136;
assign w8444 = ~w8442 & ~w8443;
assign w8445 = ~pi1134 & ~w8444;
assign w8446 = ~w8441 & ~w8445;
assign w8447 = pi1135 & ~w8446;
assign w8448 = ~w8440 & ~w8447;
assign w8449 = w8105 & ~w8448;
assign w8450 = ~pi0199 & pi0256;
assign w8451 = pi0199 & pi1070;
assign w8452 = ~w8450 & ~w8451;
assign w8453 = ~w4192 & ~w8452;
assign w8454 = pi0437 & ~pi0590;
assign w8455 = w8111 & w8454;
assign w8456 = pi0362 & pi0590;
assign w8457 = w1858 & w8456;
assign w8458 = pi0336 & w8116;
assign w8459 = pi0463 & w8118;
assign w8460 = ~w8458 & ~w8459;
assign w8461 = ~pi0590 & ~w8460;
assign w8462 = ~w8457 & ~w8461;
assign w8463 = ~pi0588 & ~w8462;
assign w8464 = ~w8455 & ~w8463;
assign w8465 = w4192 & ~w8464;
assign w8466 = ~w8453 & ~w8465;
assign w8467 = w2045 & ~w8466;
assign w8468 = ~w8449 & ~w8467;
assign w8469 = ~pi0803 & ~pi1136;
assign w8470 = pi0623 & pi1136;
assign w8471 = ~w8469 & ~w8470;
assign w8472 = ~pi1134 & ~w8471;
assign w8473 = pi0748 & pi1136;
assign w8474 = pi0876 & ~pi1136;
assign w8475 = ~w8473 & ~w8474;
assign w8476 = pi1134 & ~w8475;
assign w8477 = ~w8472 & ~w8476;
assign w8478 = ~pi1135 & ~w8477;
assign w8479 = pi0730 & w8095;
assign w8480 = pi0710 & pi1136;
assign w8481 = pi0789 & ~pi1136;
assign w8482 = ~w8480 & ~w8481;
assign w8483 = ~pi1134 & ~w8482;
assign w8484 = ~w8479 & ~w8483;
assign w8485 = pi1135 & ~w8484;
assign w8486 = ~w8478 & ~w8485;
assign w8487 = w8105 & ~w8486;
assign w8488 = ~pi0199 & pi0296;
assign w8489 = pi0199 & pi1037;
assign w8490 = ~w8488 & ~w8489;
assign w8491 = ~w4192 & ~w8490;
assign w8492 = pi0436 & ~pi0590;
assign w8493 = w8111 & w8492;
assign w8494 = pi0388 & w8116;
assign w8495 = pi0412 & w8118;
assign w8496 = ~w8494 & ~w8495;
assign w8497 = ~pi0590 & ~w8496;
assign w8498 = pi0455 & pi0590;
assign w8499 = w1858 & w8498;
assign w8500 = ~w8497 & ~w8499;
assign w8501 = ~pi0588 & ~w8500;
assign w8502 = ~w8493 & ~w8501;
assign w8503 = w4192 & ~w8502;
assign w8504 = ~w8491 & ~w8503;
assign w8505 = w2045 & ~w8504;
assign w8506 = ~w8487 & ~w8505;
assign w8507 = ~pi0812 & ~pi1136;
assign w8508 = pi0606 & pi1136;
assign w8509 = ~w8507 & ~w8508;
assign w8510 = ~pi1134 & ~w8509;
assign w8511 = pi0746 & pi1136;
assign w8512 = pi0881 & ~pi1136;
assign w8513 = ~w8511 & ~w8512;
assign w8514 = pi1134 & ~w8513;
assign w8515 = ~w8510 & ~w8514;
assign w8516 = ~pi1135 & ~w8515;
assign w8517 = pi0729 & w8095;
assign w8518 = pi0643 & pi1136;
assign w8519 = pi0787 & ~pi1136;
assign w8520 = ~w8518 & ~w8519;
assign w8521 = ~pi1134 & ~w8520;
assign w8522 = ~w8517 & ~w8521;
assign w8523 = pi1135 & ~w8522;
assign w8524 = ~w8516 & ~w8523;
assign w8525 = w8105 & ~w8524;
assign w8526 = ~pi0199 & pi0293;
assign w8527 = pi0199 & pi1059;
assign w8528 = ~w8526 & ~w8527;
assign w8529 = ~w4192 & ~w8528;
assign w8530 = pi0434 & ~pi0590;
assign w8531 = w8111 & w8530;
assign w8532 = pi0410 & w8118;
assign w8533 = pi0386 & w8116;
assign w8534 = ~w8532 & ~w8533;
assign w8535 = ~pi0590 & ~w8534;
assign w8536 = pi0361 & pi0590;
assign w8537 = w1858 & w8536;
assign w8538 = ~w8535 & ~w8537;
assign w8539 = ~pi0588 & ~w8538;
assign w8540 = ~w8531 & ~w8539;
assign w8541 = w4192 & ~w8540;
assign w8542 = ~w8529 & ~w8541;
assign w8543 = w2045 & ~w8542;
assign w8544 = ~w8525 & ~w8543;
assign w8545 = pi0870 & w8300;
assign w8546 = pi0620 & ~pi1135;
assign w8547 = ~pi0635 & pi1135;
assign w8548 = ~w8546 & ~w8547;
assign w8549 = ~pi1134 & ~w8548;
assign w8550 = ~pi0704 & pi1135;
assign w8551 = ~pi0742 & ~pi1135;
assign w8552 = ~w8550 & ~w8551;
assign w8553 = pi1134 & ~w8552;
assign w8554 = ~w8549 & ~w8553;
assign w8555 = pi1136 & ~w8554;
assign w8556 = ~w8545 & ~w8555;
assign w8557 = w8105 & ~w8556;
assign w8558 = ~pi0199 & pi0259;
assign w8559 = pi0199 & pi1069;
assign w8560 = ~w8558 & ~w8559;
assign w8561 = ~w4192 & ~w8560;
assign w8562 = pi0416 & ~pi0590;
assign w8563 = w8111 & w8562;
assign w8564 = pi0366 & w8116;
assign w8565 = pi0335 & w8118;
assign w8566 = ~w8564 & ~w8565;
assign w8567 = ~pi0590 & ~w8566;
assign w8568 = pi0344 & pi0590;
assign w8569 = w1858 & w8568;
assign w8570 = ~w8567 & ~w8569;
assign w8571 = ~pi0588 & ~w8570;
assign w8572 = ~w8563 & ~w8571;
assign w8573 = w4192 & ~w8572;
assign w8574 = ~w8561 & ~w8573;
assign w8575 = w2045 & ~w8574;
assign w8576 = ~w8557 & ~w8575;
assign w8577 = pi0856 & w8300;
assign w8578 = pi0613 & ~pi1135;
assign w8579 = ~pi0632 & pi1135;
assign w8580 = ~w8578 & ~w8579;
assign w8581 = ~pi1134 & ~w8580;
assign w8582 = ~pi0688 & pi1135;
assign w8583 = ~pi0760 & ~pi1135;
assign w8584 = ~w8582 & ~w8583;
assign w8585 = pi1134 & ~w8584;
assign w8586 = ~w8581 & ~w8585;
assign w8587 = pi1136 & ~w8586;
assign w8588 = ~w8577 & ~w8587;
assign w8589 = w8105 & ~w8588;
assign w8590 = ~pi0199 & pi0260;
assign w8591 = pi0199 & pi1067;
assign w8592 = ~w8590 & ~w8591;
assign w8593 = ~w4192 & ~w8592;
assign w8594 = pi0418 & ~pi0590;
assign w8595 = w8111 & w8594;
assign w8596 = pi0393 & w8118;
assign w8597 = pi0368 & w8116;
assign w8598 = ~w8596 & ~w8597;
assign w8599 = ~pi0590 & ~w8598;
assign w8600 = pi0346 & pi0590;
assign w8601 = w1858 & w8600;
assign w8602 = ~w8599 & ~w8601;
assign w8603 = ~pi0588 & ~w8602;
assign w8604 = ~w8595 & ~w8603;
assign w8605 = w4192 & ~w8604;
assign w8606 = ~w8593 & ~w8605;
assign w8607 = w2045 & ~w8606;
assign w8608 = ~w8589 & ~w8607;
assign w8609 = ~pi0810 & ~pi1136;
assign w8610 = ~pi0621 & pi1136;
assign w8611 = ~w8609 & ~w8610;
assign w8612 = ~pi1134 & ~w8611;
assign w8613 = ~pi0739 & pi1136;
assign w8614 = ~pi0874 & ~pi1136;
assign w8615 = ~w8613 & ~w8614;
assign w8616 = pi1134 & ~w8615;
assign w8617 = ~w8612 & ~w8616;
assign w8618 = ~pi1135 & w8617;
assign w8619 = pi0690 & w8095;
assign w8620 = pi0665 & pi1136;
assign w8621 = pi0791 & ~pi1136;
assign w8622 = ~w8620 & ~w8621;
assign w8623 = ~pi1134 & ~w8622;
assign w8624 = ~w8619 & ~w8623;
assign w8625 = pi1135 & ~w8624;
assign w8626 = ~w8618 & ~w8625;
assign w8627 = w8105 & ~w8626;
assign w8628 = ~pi0199 & pi0255;
assign w8629 = pi0199 & pi1036;
assign w8630 = ~w8628 & ~w8629;
assign w8631 = ~w4192 & ~w8630;
assign w8632 = pi0438 & ~pi0590;
assign w8633 = w8111 & w8632;
assign w8634 = pi0389 & w8116;
assign w8635 = pi0413 & w8118;
assign w8636 = ~w8634 & ~w8635;
assign w8637 = ~pi0590 & ~w8636;
assign w8638 = pi0450 & pi0590;
assign w8639 = w1858 & w8638;
assign w8640 = ~w8637 & ~w8639;
assign w8641 = ~pi0588 & ~w8640;
assign w8642 = ~w8633 & ~w8641;
assign w8643 = w4192 & ~w8642;
assign w8644 = ~w8631 & ~w8643;
assign w8645 = w2045 & ~w8644;
assign w8646 = ~w8627 & ~w8645;
assign w8647 = pi0680 & ~w7920;
assign w8648 = pi1100 & w7920;
assign w8649 = ~w8647 & ~w8648;
assign w8650 = ~pi0962 & ~w8649;
assign w8651 = pi0681 & ~w7920;
assign w8652 = pi1103 & w7920;
assign w8653 = ~w8651 & ~w8652;
assign w8654 = ~pi0962 & ~w8653;
assign w8655 = pi0848 & w8300;
assign w8656 = pi0610 & ~pi1135;
assign w8657 = ~pi0631 & pi1135;
assign w8658 = ~w8656 & ~w8657;
assign w8659 = ~pi1134 & ~w8658;
assign w8660 = ~pi0686 & pi1135;
assign w8661 = ~pi0757 & ~pi1135;
assign w8662 = ~w8660 & ~w8661;
assign w8663 = pi1134 & ~w8662;
assign w8664 = ~w8659 & ~w8663;
assign w8665 = pi1136 & ~w8664;
assign w8666 = ~w8655 & ~w8665;
assign w8667 = w8105 & ~w8666;
assign w8668 = ~pi0199 & pi0251;
assign w8669 = pi0199 & pi1039;
assign w8670 = ~w8668 & ~w8669;
assign w8671 = ~w4192 & ~w8670;
assign w8672 = pi0417 & ~pi0590;
assign w8673 = w8111 & w8672;
assign w8674 = pi0392 & w8118;
assign w8675 = pi0367 & w8116;
assign w8676 = ~w8674 & ~w8675;
assign w8677 = ~pi0590 & ~w8676;
assign w8678 = pi0345 & pi0590;
assign w8679 = w1858 & w8678;
assign w8680 = ~w8677 & ~w8679;
assign w8681 = ~pi0588 & ~w8680;
assign w8682 = ~w8673 & ~w8681;
assign w8683 = w4192 & ~w8682;
assign w8684 = ~w8671 & ~w8683;
assign w8685 = w2045 & ~w8684;
assign w8686 = ~w8667 & ~w8685;
assign w8687 = pi0832 & pi0953;
assign w8688 = ~pi0973 & w8687;
assign w8689 = ~pi1054 & w8688;
assign w8690 = pi1066 & w8689;
assign w8691 = pi1088 & w8690;
assign w8692 = ~pi0684 & ~w8691;
assign w8693 = pi1130 & w8691;
assign w8694 = ~w8692 & ~w8693;
assign w8695 = ~pi0962 & ~w8694;
assign w8696 = ~pi0199 & ~w5927;
assign w8697 = pi0199 & pi1076;
assign w8698 = ~w8696 & ~w8697;
assign w8699 = ~w4192 & ~w8698;
assign w8700 = pi0430 & ~pi0590;
assign w8701 = w8111 & w8700;
assign w8702 = pi0406 & w8118;
assign w8703 = pi0382 & w8116;
assign w8704 = ~w8702 & ~w8703;
assign w8705 = ~pi0590 & ~w8704;
assign w8706 = pi0357 & pi0590;
assign w8707 = w1858 & w8706;
assign w8708 = ~w8705 & ~w8707;
assign w8709 = ~pi0588 & ~w8708;
assign w8710 = ~w8701 & ~w8709;
assign w8711 = w4192 & ~w8710;
assign w8712 = ~w8699 & ~w8711;
assign w8713 = w2045 & ~w8712;
assign w8714 = pi0813 & ~pi1134;
assign w8715 = pi0860 & pi1134;
assign w8716 = ~w8714 & ~w8715;
assign w8717 = ~pi1136 & ~w8716;
assign w8718 = ~pi1135 & w8717;
assign w8719 = pi0652 & ~pi1135;
assign w8720 = ~pi0657 & pi1135;
assign w8721 = ~w8719 & ~w8720;
assign w8722 = ~pi1134 & ~w8721;
assign w8723 = ~pi0728 & pi1135;
assign w8724 = ~pi0744 & ~pi1135;
assign w8725 = ~w8723 & ~w8724;
assign w8726 = pi1134 & ~w8725;
assign w8727 = ~w8722 & ~w8726;
assign w8728 = pi1136 & ~w8727;
assign w8729 = ~w8718 & ~w8728;
assign w8730 = w8105 & ~w8729;
assign w8731 = ~w8713 & ~w8730;
assign w8732 = ~pi0686 & ~w8691;
assign w8733 = pi1113 & w8691;
assign w8734 = ~w8732 & ~w8733;
assign w8735 = ~pi0962 & ~w8734;
assign w8736 = pi0687 & ~w8691;
assign w8737 = pi1127 & w8691;
assign w8738 = ~w8736 & ~w8737;
assign w8739 = ~pi0962 & ~w8738;
assign w8740 = ~pi0688 & ~w8691;
assign w8741 = pi1115 & w8691;
assign w8742 = ~w8740 & ~w8741;
assign w8743 = ~pi0962 & ~w8742;
assign w8744 = ~pi0199 & ~w5897;
assign w8745 = pi0199 & pi1079;
assign w8746 = ~w8744 & ~w8745;
assign w8747 = ~w4192 & ~w8746;
assign w8748 = pi0426 & ~pi0590;
assign w8749 = w8111 & w8748;
assign w8750 = pi0401 & w8118;
assign w8751 = pi0376 & w8116;
assign w8752 = ~w8750 & ~w8751;
assign w8753 = ~pi0590 & ~w8752;
assign w8754 = pi0351 & pi0590;
assign w8755 = w1858 & w8754;
assign w8756 = ~w8753 & ~w8755;
assign w8757 = ~pi0588 & ~w8756;
assign w8758 = ~w8749 & ~w8757;
assign w8759 = w4192 & ~w8758;
assign w8760 = ~w8747 & ~w8759;
assign w8761 = w2045 & ~w8760;
assign w8762 = pi0798 & ~pi1134;
assign w8763 = pi0843 & pi1134;
assign w8764 = ~w8762 & ~w8763;
assign w8765 = ~pi1136 & ~w8764;
assign w8766 = ~pi1135 & w8765;
assign w8767 = pi0655 & pi1135;
assign w8768 = ~pi0658 & ~pi1135;
assign w8769 = ~w8767 & ~w8768;
assign w8770 = ~pi1134 & ~w8769;
assign w8771 = ~pi0703 & pi1135;
assign w8772 = pi0752 & ~pi1135;
assign w8773 = ~w8771 & ~w8772;
assign w8774 = pi1134 & ~w8773;
assign w8775 = ~w8770 & ~w8774;
assign w8776 = pi1136 & w8775;
assign w8777 = ~w8766 & ~w8776;
assign w8778 = w8105 & ~w8777;
assign w8779 = ~w8761 & ~w8778;
assign w8780 = pi0690 & ~w8691;
assign w8781 = pi1108 & w8691;
assign w8782 = ~w8780 & ~w8781;
assign w8783 = ~pi0962 & ~w8782;
assign w8784 = pi0691 & ~w8691;
assign w8785 = pi1107 & w8691;
assign w8786 = ~w8784 & ~w8785;
assign w8787 = ~pi0962 & ~w8786;
assign w8788 = ~pi0199 & ~w5909;
assign w8789 = pi0199 & pi1078;
assign w8790 = ~w8788 & ~w8789;
assign w8791 = ~w4192 & ~w8790;
assign w8792 = pi0427 & ~pi0590;
assign w8793 = w8111 & w8792;
assign w8794 = pi0352 & pi0590;
assign w8795 = w1858 & w8794;
assign w8796 = pi0317 & w8116;
assign w8797 = pi0402 & w8118;
assign w8798 = ~w8796 & ~w8797;
assign w8799 = ~pi0590 & ~w8798;
assign w8800 = ~w8795 & ~w8799;
assign w8801 = ~pi0588 & ~w8800;
assign w8802 = ~w8793 & ~w8801;
assign w8803 = w4192 & ~w8802;
assign w8804 = ~w8791 & ~w8803;
assign w8805 = w2045 & ~w8804;
assign w8806 = pi0801 & ~pi1134;
assign w8807 = pi0844 & pi1134;
assign w8808 = ~w8806 & ~w8807;
assign w8809 = ~pi1136 & ~w8808;
assign w8810 = ~pi1135 & w8809;
assign w8811 = pi0649 & pi1135;
assign w8812 = ~pi0656 & ~pi1135;
assign w8813 = ~w8811 & ~w8812;
assign w8814 = ~pi1134 & ~w8813;
assign w8815 = ~pi0726 & pi1135;
assign w8816 = pi0770 & ~pi1135;
assign w8817 = ~w8815 & ~w8816;
assign w8818 = pi1134 & ~w8817;
assign w8819 = ~w8814 & ~w8818;
assign w8820 = pi1136 & w8819;
assign w8821 = ~w8810 & ~w8820;
assign w8822 = w8105 & ~w8821;
assign w8823 = ~w8805 & ~w8822;
assign w8824 = ~pi0693 & ~w7920;
assign w8825 = pi1129 & w7920;
assign w8826 = ~w8824 & ~w8825;
assign w8827 = ~pi0962 & ~w8826;
assign w8828 = ~pi0694 & ~w8691;
assign w8829 = pi1128 & w8691;
assign w8830 = ~w8828 & ~w8829;
assign w8831 = ~pi0962 & ~w8830;
assign w8832 = ~pi0695 & ~w7920;
assign w8833 = pi1111 & w7920;
assign w8834 = ~w8832 & ~w8833;
assign w8835 = ~pi0962 & ~w8834;
assign w8836 = pi0696 & ~w8691;
assign w8837 = pi1100 & w8691;
assign w8838 = ~w8836 & ~w8837;
assign w8839 = ~pi0962 & ~w8838;
assign w8840 = ~pi0697 & ~w8691;
assign w8841 = pi1129 & w8691;
assign w8842 = ~w8840 & ~w8841;
assign w8843 = ~pi0962 & ~w8842;
assign w8844 = ~pi0698 & ~w8691;
assign w8845 = pi1116 & w8691;
assign w8846 = ~w8844 & ~w8845;
assign w8847 = ~pi0962 & ~w8846;
assign w8848 = pi0699 & ~w8691;
assign w8849 = pi1103 & w8691;
assign w8850 = ~w8848 & ~w8849;
assign w8851 = ~pi0962 & ~w8850;
assign w8852 = pi0700 & ~w8691;
assign w8853 = pi1110 & w8691;
assign w8854 = ~w8852 & ~w8853;
assign w8855 = ~pi0962 & ~w8854;
assign w8856 = ~pi0701 & ~w8691;
assign w8857 = pi1123 & w8691;
assign w8858 = ~w8856 & ~w8857;
assign w8859 = ~pi0962 & ~w8858;
assign w8860 = ~pi0702 & ~w8691;
assign w8861 = pi1117 & w8691;
assign w8862 = ~w8860 & ~w8861;
assign w8863 = ~pi0962 & ~w8862;
assign w8864 = pi0703 & ~w8691;
assign w8865 = pi1124 & w8691;
assign w8866 = ~w8864 & ~w8865;
assign w8867 = ~pi0962 & ~w8866;
assign w8868 = ~pi0704 & ~w8691;
assign w8869 = pi1112 & w8691;
assign w8870 = ~w8868 & ~w8869;
assign w8871 = ~pi0962 & ~w8870;
assign w8872 = pi0705 & ~w8691;
assign w8873 = pi1125 & w8691;
assign w8874 = ~w8872 & ~w8873;
assign w8875 = ~pi0962 & ~w8874;
assign w8876 = pi0706 & ~w8691;
assign w8877 = pi1105 & w8691;
assign w8878 = ~w8876 & ~w8877;
assign w8879 = ~pi0962 & ~w8878;
assign w8880 = pi0200 & pi1048;
assign w8881 = ~pi0200 & pi0304;
assign w8882 = ~w8880 & ~w8881;
assign w8883 = ~pi0199 & ~w8882;
assign w8884 = pi0199 & pi1055;
assign w8885 = ~w8883 & ~w8884;
assign w8886 = ~w4192 & ~w8885;
assign w8887 = pi0420 & ~pi0590;
assign w8888 = w8111 & w8887;
assign w8889 = pi0395 & w8118;
assign w8890 = pi0370 & w8116;
assign w8891 = ~w8889 & ~w8890;
assign w8892 = ~pi0590 & ~w8891;
assign w8893 = pi0347 & pi0590;
assign w8894 = w1858 & w8893;
assign w8895 = ~w8892 & ~w8894;
assign w8896 = ~pi0588 & ~w8895;
assign w8897 = ~w8888 & ~w8896;
assign w8898 = w4192 & ~w8897;
assign w8899 = ~w8886 & ~w8898;
assign w8900 = w2045 & ~w8899;
assign w8901 = pi0847 & w8300;
assign w8902 = pi0627 & pi1135;
assign w8903 = pi0618 & ~pi1135;
assign w8904 = ~w8902 & ~w8903;
assign w8905 = ~pi1134 & ~w8904;
assign w8906 = ~pi0702 & pi1135;
assign w8907 = ~pi0753 & ~pi1135;
assign w8908 = ~w8906 & ~w8907;
assign w8909 = pi1134 & ~w8908;
assign w8910 = ~w8905 & ~w8909;
assign w8911 = pi1136 & ~w8910;
assign w8912 = ~w8901 & ~w8911;
assign w8913 = w8105 & ~w8912;
assign w8914 = ~w8900 & ~w8913;
assign w8915 = ~pi0200 & pi0305;
assign w8916 = pi0200 & pi1084;
assign w8917 = ~w8915 & ~w8916;
assign w8918 = ~pi0199 & ~w8917;
assign w8919 = pi0199 & pi1058;
assign w8920 = ~w8918 & ~w8919;
assign w8921 = ~w4192 & ~w8920;
assign w8922 = pi0459 & ~pi0590;
assign w8923 = w8111 & w8922;
assign w8924 = pi0321 & pi0590;
assign w8925 = w1858 & w8924;
assign w8926 = pi0442 & w8116;
assign w8927 = pi0328 & w8118;
assign w8928 = ~w8926 & ~w8927;
assign w8929 = ~pi0590 & ~w8928;
assign w8930 = ~w8925 & ~w8929;
assign w8931 = ~pi0588 & ~w8930;
assign w8932 = ~w8923 & ~w8931;
assign w8933 = w4192 & ~w8932;
assign w8934 = ~w8921 & ~w8933;
assign w8935 = w2045 & ~w8934;
assign w8936 = pi0857 & w8300;
assign w8937 = pi0660 & pi1135;
assign w8938 = pi0609 & ~pi1135;
assign w8939 = ~w8937 & ~w8938;
assign w8940 = ~pi1134 & ~w8939;
assign w8941 = ~pi0709 & pi1135;
assign w8942 = ~pi0754 & ~pi1135;
assign w8943 = ~w8941 & ~w8942;
assign w8944 = pi1134 & ~w8943;
assign w8945 = ~w8940 & ~w8944;
assign w8946 = pi1136 & ~w8945;
assign w8947 = ~w8936 & ~w8946;
assign w8948 = w8105 & ~w8947;
assign w8949 = ~w8935 & ~w8948;
assign w8950 = ~pi0709 & ~w8691;
assign w8951 = pi1118 & w8691;
assign w8952 = ~w8950 & ~w8951;
assign w8953 = ~pi0962 & ~w8952;
assign w8954 = pi0710 & ~w7920;
assign w8955 = pi1106 & w7920;
assign w8956 = ~w8954 & ~w8955;
assign w8957 = ~pi0962 & ~w8956;
assign w8958 = pi0200 & pi1059;
assign w8959 = ~pi0200 & pi0306;
assign w8960 = ~w8958 & ~w8959;
assign w8961 = ~pi0199 & ~w8960;
assign w8962 = pi0199 & pi1087;
assign w8963 = ~w8961 & ~w8962;
assign w8964 = ~w4192 & ~w8963;
assign w8965 = pi0423 & ~pi0590;
assign w8966 = w8111 & w8965;
assign w8967 = pi0398 & w8118;
assign w8968 = pi0373 & w8116;
assign w8969 = ~w8967 & ~w8968;
assign w8970 = ~pi0590 & ~w8969;
assign w8971 = pi0348 & pi0590;
assign w8972 = w1858 & w8971;
assign w8973 = ~w8970 & ~w8972;
assign w8974 = ~pi0588 & ~w8973;
assign w8975 = ~w8966 & ~w8974;
assign w8976 = w4192 & ~w8975;
assign w8977 = ~w8964 & ~w8976;
assign w8978 = w2045 & ~w8977;
assign w8979 = pi0858 & w8300;
assign w8980 = pi0647 & pi1135;
assign w8981 = pi0630 & ~pi1135;
assign w8982 = ~w8980 & ~w8981;
assign w8983 = ~pi1134 & ~w8982;
assign w8984 = ~pi0725 & pi1135;
assign w8985 = ~pi0755 & ~pi1135;
assign w8986 = ~w8984 & ~w8985;
assign w8987 = pi1134 & ~w8986;
assign w8988 = ~w8983 & ~w8987;
assign w8989 = pi1136 & ~w8988;
assign w8990 = ~w8979 & ~w8989;
assign w8991 = w8105 & ~w8990;
assign w8992 = ~w8978 & ~w8991;
assign w8993 = ~pi0200 & pi0298;
assign w8994 = pi0200 & pi1044;
assign w8995 = ~w8993 & ~w8994;
assign w8996 = ~pi0199 & ~w8995;
assign w8997 = pi0199 & pi1035;
assign w8998 = ~w8996 & ~w8997;
assign w8999 = ~w4192 & ~w8998;
assign w9000 = pi0425 & ~pi0590;
assign w9001 = w8111 & w9000;
assign w9002 = pi0400 & w8118;
assign w9003 = pi0374 & w8116;
assign w9004 = ~w9002 & ~w9003;
assign w9005 = ~pi0590 & ~w9004;
assign w9006 = pi0350 & pi0590;
assign w9007 = w1858 & w9006;
assign w9008 = ~w9005 & ~w9007;
assign w9009 = ~pi0588 & ~w9008;
assign w9010 = ~w9001 & ~w9009;
assign w9011 = w4192 & ~w9010;
assign w9012 = ~w8999 & ~w9011;
assign w9013 = w2045 & ~w9012;
assign w9014 = pi0842 & w8300;
assign w9015 = pi0644 & ~pi1135;
assign w9016 = pi0715 & pi1135;
assign w9017 = ~w9015 & ~w9016;
assign w9018 = ~pi1134 & ~w9017;
assign w9019 = ~pi0701 & pi1135;
assign w9020 = ~pi0751 & ~pi1135;
assign w9021 = ~w9019 & ~w9020;
assign w9022 = pi1134 & ~w9021;
assign w9023 = ~w9018 & ~w9022;
assign w9024 = pi1136 & ~w9023;
assign w9025 = ~w9014 & ~w9024;
assign w9026 = w8105 & ~w9025;
assign w9027 = ~w9013 & ~w9026;
assign w9028 = ~pi0200 & pi0309;
assign w9029 = pi0200 & pi1072;
assign w9030 = ~w9028 & ~w9029;
assign w9031 = ~pi0199 & ~w9030;
assign w9032 = pi0199 & pi1051;
assign w9033 = ~w9031 & ~w9032;
assign w9034 = ~w4192 & ~w9033;
assign w9035 = pi0421 & ~pi0590;
assign w9036 = w8111 & w9035;
assign w9037 = pi0396 & w8118;
assign w9038 = pi0371 & w8116;
assign w9039 = ~w9037 & ~w9038;
assign w9040 = ~pi0590 & ~w9039;
assign w9041 = pi0322 & pi0590;
assign w9042 = w1858 & w9041;
assign w9043 = ~w9040 & ~w9042;
assign w9044 = ~pi0588 & ~w9043;
assign w9045 = ~w9036 & ~w9044;
assign w9046 = w4192 & ~w9045;
assign w9047 = ~w9034 & ~w9046;
assign w9048 = w2045 & ~w9047;
assign w9049 = pi0854 & w8300;
assign w9050 = pi0628 & pi1135;
assign w9051 = pi0629 & ~pi1135;
assign w9052 = ~w9050 & ~w9051;
assign w9053 = ~pi1134 & ~w9052;
assign w9054 = ~pi0734 & pi1135;
assign w9055 = ~pi0756 & ~pi1135;
assign w9056 = ~w9054 & ~w9055;
assign w9057 = pi1134 & ~w9056;
assign w9058 = ~w9053 & ~w9057;
assign w9059 = pi1136 & ~w9058;
assign w9060 = ~w9049 & ~w9059;
assign w9061 = w8105 & ~w9060;
assign w9062 = ~w9048 & ~w9061;
assign w9063 = ~pi0199 & ~w5853;
assign w9064 = pi0199 & pi1057;
assign w9065 = ~w9063 & ~w9064;
assign w9066 = ~w4192 & ~w9065;
assign w9067 = pi0449 & ~pi0590;
assign w9068 = w8111 & w9067;
assign w9069 = pi0461 & pi0590;
assign w9070 = w1858 & w9069;
assign w9071 = pi0439 & w8116;
assign w9072 = pi0326 & w8118;
assign w9073 = ~w9071 & ~w9072;
assign w9074 = ~pi0590 & ~w9073;
assign w9075 = ~w9070 & ~w9074;
assign w9076 = ~pi0588 & ~w9075;
assign w9077 = ~w9068 & ~w9076;
assign w9078 = w4192 & ~w9077;
assign w9079 = ~w9066 & ~w9078;
assign w9080 = w2045 & ~w9079;
assign w9081 = pi0816 & ~pi1134;
assign w9082 = pi0867 & pi1134;
assign w9083 = ~w9081 & ~w9082;
assign w9084 = ~pi1136 & ~w9083;
assign w9085 = ~pi1135 & w9084;
assign w9086 = pi0653 & ~pi1135;
assign w9087 = ~pi0693 & pi1135;
assign w9088 = ~w9086 & ~w9087;
assign w9089 = ~pi1134 & ~w9088;
assign w9090 = ~pi0697 & pi1135;
assign w9091 = ~pi0762 & ~pi1135;
assign w9092 = ~w9090 & ~w9091;
assign w9093 = pi1134 & ~w9092;
assign w9094 = ~w9089 & ~w9093;
assign w9095 = pi1136 & ~w9094;
assign w9096 = ~w9085 & ~w9095;
assign w9097 = w8105 & ~w9096;
assign w9098 = ~w9080 & ~w9097;
assign w9099 = pi0715 & ~w7920;
assign w9100 = pi1123 & w7920;
assign w9101 = ~w9099 & ~w9100;
assign w9102 = ~pi0962 & ~w9101;
assign w9103 = ~pi0200 & pi0307;
assign w9104 = pi0200 & pi1053;
assign w9105 = ~w9103 & ~w9104;
assign w9106 = ~pi0199 & ~w9105;
assign w9107 = pi0199 & pi1043;
assign w9108 = ~w9106 & ~w9107;
assign w9109 = ~w4192 & ~w9108;
assign w9110 = pi0454 & ~pi0590;
assign w9111 = w8111 & w9110;
assign w9112 = pi0440 & w8116;
assign w9113 = pi0329 & w8118;
assign w9114 = ~w9112 & ~w9113;
assign w9115 = ~pi0590 & ~w9114;
assign w9116 = pi0349 & pi0590;
assign w9117 = w1858 & w9116;
assign w9118 = ~w9115 & ~w9117;
assign w9119 = ~pi0588 & ~w9118;
assign w9120 = ~w9111 & ~w9119;
assign w9121 = w4192 & ~w9120;
assign w9122 = ~w9109 & ~w9121;
assign w9123 = w2045 & ~w9122;
assign w9124 = pi0845 & w8300;
assign w9125 = pi0641 & pi1135;
assign w9126 = pi0626 & ~pi1135;
assign w9127 = ~w9125 & ~w9126;
assign w9128 = ~pi1134 & ~w9127;
assign w9129 = ~pi0738 & pi1135;
assign w9130 = ~pi0761 & ~pi1135;
assign w9131 = ~w9129 & ~w9130;
assign w9132 = pi1134 & ~w9131;
assign w9133 = ~w9128 & ~w9132;
assign w9134 = pi1136 & ~w9133;
assign w9135 = ~w9124 & ~w9134;
assign w9136 = w8105 & ~w9135;
assign w9137 = ~w9123 & ~w9136;
assign w9138 = ~pi0199 & ~w5903;
assign w9139 = pi0199 & pi1074;
assign w9140 = ~w9138 & ~w9139;
assign w9141 = ~w4192 & ~w9140;
assign w9142 = pi0448 & ~pi0590;
assign w9143 = w8111 & w9142;
assign w9144 = pi0462 & pi0590;
assign w9145 = w1858 & w9144;
assign w9146 = pi0377 & w8116;
assign w9147 = pi0318 & w8118;
assign w9148 = ~w9146 & ~w9147;
assign w9149 = ~pi0590 & ~w9148;
assign w9150 = ~w9145 & ~w9149;
assign w9151 = ~pi0588 & ~w9150;
assign w9152 = ~w9143 & ~w9151;
assign w9153 = w4192 & ~w9152;
assign w9154 = ~w9141 & ~w9153;
assign w9155 = w2045 & ~w9154;
assign w9156 = pi0800 & ~pi1134;
assign w9157 = pi0839 & pi1134;
assign w9158 = ~w9156 & ~w9157;
assign w9159 = ~pi1136 & ~w9158;
assign w9160 = ~pi1135 & w9159;
assign w9161 = pi0705 & pi1135;
assign w9162 = ~pi0768 & ~pi1135;
assign w9163 = ~w9161 & ~w9162;
assign w9164 = pi1134 & ~w9163;
assign w9165 = pi0645 & ~pi1135;
assign w9166 = ~pi0669 & pi1135;
assign w9167 = ~w9165 & ~w9166;
assign w9168 = ~pi1134 & ~w9167;
assign w9169 = ~w9164 & ~w9168;
assign w9170 = pi1136 & ~w9169;
assign w9171 = ~w9160 & ~w9170;
assign w9172 = w8105 & ~w9171;
assign w9173 = ~w9155 & ~w9172;
assign w9174 = pi0200 & pi1049;
assign w9175 = ~pi0200 & pi0303;
assign w9176 = ~w9174 & ~w9175;
assign w9177 = ~pi0199 & ~w9176;
assign w9178 = pi0199 & pi1080;
assign w9179 = ~w9177 & ~w9178;
assign w9180 = ~w4192 & ~w9179;
assign w9181 = pi0419 & ~pi0590;
assign w9182 = w8111 & w9181;
assign w9183 = pi0394 & w8118;
assign w9184 = pi0369 & w8116;
assign w9185 = ~w9183 & ~w9184;
assign w9186 = ~pi0590 & ~w9185;
assign w9187 = pi0315 & pi0590;
assign w9188 = w1858 & w9187;
assign w9189 = ~w9186 & ~w9188;
assign w9190 = ~pi0588 & ~w9189;
assign w9191 = ~w9182 & ~w9190;
assign w9192 = w4192 & ~w9191;
assign w9193 = ~w9180 & ~w9192;
assign w9194 = w2045 & ~w9193;
assign w9195 = pi0853 & w8300;
assign w9196 = pi0625 & pi1135;
assign w9197 = pi0608 & ~pi1135;
assign w9198 = ~w9196 & ~w9197;
assign w9199 = ~pi1134 & ~w9198;
assign w9200 = ~pi0698 & pi1135;
assign w9201 = ~pi0767 & ~pi1135;
assign w9202 = ~w9200 & ~w9201;
assign w9203 = pi1134 & ~w9202;
assign w9204 = ~w9199 & ~w9203;
assign w9205 = pi1136 & ~w9204;
assign w9206 = ~w9195 & ~w9205;
assign w9207 = w8105 & ~w9206;
assign w9208 = ~w9194 & ~w9207;
assign w9209 = ~pi0199 & ~w5915;
assign w9210 = pi0199 & pi1063;
assign w9211 = ~w9209 & ~w9210;
assign w9212 = ~w4192 & ~w9211;
assign w9213 = pi0451 & ~pi0590;
assign w9214 = w8111 & w9213;
assign w9215 = pi0378 & w8116;
assign w9216 = pi0325 & w8118;
assign w9217 = ~w9215 & ~w9216;
assign w9218 = ~pi0590 & ~w9217;
assign w9219 = pi0353 & pi0590;
assign w9220 = w1858 & w9219;
assign w9221 = ~w9218 & ~w9220;
assign w9222 = ~pi0588 & ~w9221;
assign w9223 = ~w9214 & ~w9222;
assign w9224 = w4192 & ~w9223;
assign w9225 = ~w9212 & ~w9224;
assign w9226 = w2045 & ~w9225;
assign w9227 = pi0807 & ~pi1134;
assign w9228 = pi0868 & pi1134;
assign w9229 = ~w9227 & ~w9228;
assign w9230 = ~pi1136 & ~w9229;
assign w9231 = ~pi1135 & w9230;
assign w9232 = pi0687 & pi1135;
assign w9233 = ~pi0774 & ~pi1135;
assign w9234 = ~w9232 & ~w9233;
assign w9235 = pi1134 & ~w9234;
assign w9236 = pi0636 & ~pi1135;
assign w9237 = ~pi0650 & pi1135;
assign w9238 = ~w9236 & ~w9237;
assign w9239 = ~pi1134 & ~w9238;
assign w9240 = ~w9235 & ~w9239;
assign w9241 = pi1136 & ~w9240;
assign w9242 = ~w9231 & ~w9241;
assign w9243 = w8105 & ~w9242;
assign w9244 = ~w9226 & ~w9243;
assign w9245 = ~pi0199 & ~w5933;
assign w9246 = pi0199 & pi1081;
assign w9247 = ~w9245 & ~w9246;
assign w9248 = ~w4192 & ~w9247;
assign w9249 = pi0445 & ~pi0590;
assign w9250 = w8111 & w9249;
assign w9251 = pi0405 & w8118;
assign w9252 = pi0381 & w8116;
assign w9253 = ~w9251 & ~w9252;
assign w9254 = ~pi0590 & ~w9253;
assign w9255 = pi0356 & pi0590;
assign w9256 = w1858 & w9255;
assign w9257 = ~w9254 & ~w9256;
assign w9258 = ~pi0588 & ~w9257;
assign w9259 = ~w9250 & ~w9258;
assign w9260 = w4192 & ~w9259;
assign w9261 = ~w9248 & ~w9260;
assign w9262 = w2045 & ~w9261;
assign w9263 = pi0794 & ~pi1134;
assign w9264 = pi0880 & pi1134;
assign w9265 = ~w9263 & ~w9264;
assign w9266 = ~pi1136 & ~w9265;
assign w9267 = ~pi1135 & w9266;
assign w9268 = pi0651 & ~pi1135;
assign w9269 = ~pi0654 & pi1135;
assign w9270 = ~w9268 & ~w9269;
assign w9271 = ~pi1134 & ~w9270;
assign w9272 = ~pi0684 & pi1135;
assign w9273 = ~pi0750 & ~pi1135;
assign w9274 = ~w9272 & ~w9273;
assign w9275 = pi1134 & ~w9274;
assign w9276 = ~w9271 & ~w9275;
assign w9277 = pi1136 & ~w9276;
assign w9278 = ~w9267 & ~w9277;
assign w9279 = w8105 & ~w9278;
assign w9280 = ~w9262 & ~w9279;
assign w9281 = pi0731 & pi0747;
assign w9282 = pi0773 & w9281;
assign w9283 = pi0775 & w9282;
assign w9284 = ~pi0945 & w9283;
assign w9285 = pi0988 & w9284;
assign w9286 = pi0769 & w9285;
assign w9287 = pi0721 & ~w9286;
assign w9288 = ~pi0721 & pi0769;
assign w9289 = w9285 & w9288;
assign w9290 = ~w9287 & ~w9289;
assign w9291 = pi0775 & pi0816;
assign w9292 = ~pi0775 & ~pi0816;
assign w9293 = ~w9291 & ~w9292;
assign w9294 = ~pi0731 & ~pi0795;
assign w9295 = pi0731 & pi0795;
assign w9296 = ~w9294 & ~w9295;
assign w9297 = ~w9293 & ~w9296;
assign w9298 = pi0747 & pi0807;
assign w9299 = ~pi0747 & ~pi0807;
assign w9300 = ~w9298 & ~w9299;
assign w9301 = pi0773 & pi0801;
assign w9302 = ~pi0773 & ~pi0801;
assign w9303 = ~w9301 & ~w9302;
assign w9304 = ~w9300 & ~w9303;
assign w9305 = w9297 & w9304;
assign w9306 = ~pi0771 & ~pi0800;
assign w9307 = pi0771 & pi0800;
assign w9308 = ~w9306 & ~w9307;
assign w9309 = ~pi0769 & ~pi0794;
assign w9310 = pi0769 & pi0794;
assign w9311 = ~w9309 & ~w9310;
assign w9312 = ~w9308 & ~w9311;
assign w9313 = pi0721 & pi0813;
assign w9314 = ~pi0721 & ~pi0813;
assign w9315 = ~w9313 & ~w9314;
assign w9316 = pi0765 & pi0798;
assign w9317 = ~pi0765 & ~pi0798;
assign w9318 = ~w9316 & ~w9317;
assign w9319 = ~w9315 & ~w9318;
assign w9320 = w9312 & w9319;
assign w9321 = w9305 & w9320;
assign w9322 = ~w9290 & ~w9321;
assign w9323 = ~pi0199 & ~w5921;
assign w9324 = pi0199 & pi1045;
assign w9325 = ~w9323 & ~w9324;
assign w9326 = ~w4192 & ~w9325;
assign w9327 = pi0428 & ~pi0590;
assign w9328 = w8111 & w9327;
assign w9329 = pi0403 & w8118;
assign w9330 = pi0379 & w8116;
assign w9331 = ~w9329 & ~w9330;
assign w9332 = ~pi0590 & ~w9331;
assign w9333 = pi0354 & pi0590;
assign w9334 = w1858 & w9333;
assign w9335 = ~w9332 & ~w9334;
assign w9336 = ~pi0588 & ~w9335;
assign w9337 = ~w9328 & ~w9336;
assign w9338 = w4192 & ~w9337;
assign w9339 = ~w9326 & ~w9338;
assign w9340 = w2045 & ~w9339;
assign w9341 = pi0795 & ~pi1134;
assign w9342 = pi0851 & pi1134;
assign w9343 = ~w9341 & ~w9342;
assign w9344 = ~pi1136 & ~w9343;
assign w9345 = ~pi1135 & w9344;
assign w9346 = ~pi0732 & pi1135;
assign w9347 = pi0640 & ~pi1135;
assign w9348 = ~w9346 & ~w9347;
assign w9349 = ~pi1134 & ~w9348;
assign w9350 = ~pi0694 & pi1135;
assign w9351 = ~pi0776 & ~pi1135;
assign w9352 = ~w9350 & ~w9351;
assign w9353 = pi1134 & ~w9352;
assign w9354 = ~w9349 & ~w9353;
assign w9355 = pi1136 & ~w9354;
assign w9356 = ~w9345 & ~w9355;
assign w9357 = w8105 & ~w9356;
assign w9358 = ~w9340 & ~w9357;
assign w9359 = ~pi0723 & ~w8691;
assign w9360 = pi1111 & w8691;
assign w9361 = ~w9359 & ~w9360;
assign w9362 = ~pi0962 & ~w9361;
assign w9363 = ~pi0724 & ~w8691;
assign w9364 = pi1114 & w8691;
assign w9365 = ~w9363 & ~w9364;
assign w9366 = ~pi0962 & ~w9365;
assign w9367 = ~pi0725 & ~w8691;
assign w9368 = pi1120 & w8691;
assign w9369 = ~w9367 & ~w9368;
assign w9370 = ~pi0962 & ~w9369;
assign w9371 = pi0726 & ~w8691;
assign w9372 = pi1126 & w8691;
assign w9373 = ~w9371 & ~w9372;
assign w9374 = ~pi0962 & ~w9373;
assign w9375 = pi0727 & ~w8691;
assign w9376 = pi1102 & w8691;
assign w9377 = ~w9375 & ~w9376;
assign w9378 = ~pi0962 & ~w9377;
assign w9379 = ~pi0728 & ~w8691;
assign w9380 = pi1131 & w8691;
assign w9381 = ~w9379 & ~w9380;
assign w9382 = ~pi0962 & ~w9381;
assign w9383 = pi0729 & ~w8691;
assign w9384 = pi1104 & w8691;
assign w9385 = ~w9383 & ~w9384;
assign w9386 = ~pi0962 & ~w9385;
assign w9387 = pi0730 & ~w8691;
assign w9388 = pi1106 & w8691;
assign w9389 = ~w9387 & ~w9388;
assign w9390 = ~pi0962 & ~w9389;
assign w9391 = ~pi0731 & pi0988;
assign w9392 = ~pi0945 & w9391;
assign w9393 = pi0747 & pi0773;
assign w9394 = w9392 & w9393;
assign w9395 = ~pi0945 & pi0988;
assign w9396 = w9393 & w9395;
assign w9397 = pi0731 & ~w9396;
assign w9398 = ~w9394 & ~w9397;
assign w9399 = ~w9321 & ~w9398;
assign w9400 = ~pi0732 & ~w7920;
assign w9401 = pi1128 & w7920;
assign w9402 = ~w9400 & ~w9401;
assign w9403 = ~pi0962 & ~w9402;
assign w9404 = pi0200 & pi1037;
assign w9405 = ~pi0200 & pi0308;
assign w9406 = ~w9404 & ~w9405;
assign w9407 = ~pi0199 & ~w9406;
assign w9408 = pi0199 & pi1047;
assign w9409 = ~w9407 & ~w9408;
assign w9410 = ~w4192 & ~w9409;
assign w9411 = pi0424 & ~pi0590;
assign w9412 = w8111 & w9411;
assign w9413 = pi0399 & w8118;
assign w9414 = pi0375 & w8116;
assign w9415 = ~w9413 & ~w9414;
assign w9416 = ~pi0590 & ~w9415;
assign w9417 = pi0316 & pi0590;
assign w9418 = w1858 & w9417;
assign w9419 = ~w9416 & ~w9418;
assign w9420 = ~pi0588 & ~w9419;
assign w9421 = ~w9412 & ~w9420;
assign w9422 = w4192 & ~w9421;
assign w9423 = ~w9410 & ~w9422;
assign w9424 = w2045 & ~w9423;
assign w9425 = pi0838 & w8300;
assign w9426 = pi0648 & pi1135;
assign w9427 = pi0619 & ~pi1135;
assign w9428 = ~w9426 & ~w9427;
assign w9429 = ~pi1134 & ~w9428;
assign w9430 = ~pi0737 & pi1135;
assign w9431 = ~pi0777 & ~pi1135;
assign w9432 = ~w9430 & ~w9431;
assign w9433 = pi1134 & ~w9432;
assign w9434 = ~w9429 & ~w9433;
assign w9435 = pi1136 & ~w9434;
assign w9436 = ~w9425 & ~w9435;
assign w9437 = w8105 & ~w9436;
assign w9438 = ~w9424 & ~w9437;
assign w9439 = ~pi0734 & ~w8691;
assign w9440 = pi1119 & w8691;
assign w9441 = ~w9439 & ~w9440;
assign w9442 = ~pi0962 & ~w9441;
assign w9443 = pi0735 & ~w8691;
assign w9444 = pi1109 & w8691;
assign w9445 = ~w9443 & ~w9444;
assign w9446 = ~pi0962 & ~w9445;
assign w9447 = pi0736 & ~w8691;
assign w9448 = pi1101 & w8691;
assign w9449 = ~w9447 & ~w9448;
assign w9450 = ~pi0962 & ~w9449;
assign w9451 = ~pi0737 & ~w8691;
assign w9452 = pi1122 & w8691;
assign w9453 = ~w9451 & ~w9452;
assign w9454 = ~pi0962 & ~w9453;
assign w9455 = ~pi0738 & ~w8691;
assign w9456 = pi1121 & w8691;
assign w9457 = ~w9455 & ~w9456;
assign w9458 = ~pi0962 & ~w9457;
assign w9459 = pi0832 & ~pi0952;
assign w9460 = ~pi0980 & w9459;
assign w9461 = pi1038 & w9460;
assign w9462 = pi1060 & w9461;
assign w9463 = ~pi1061 & w9462;
assign w9464 = ~pi1108 & w9463;
assign w9465 = ~pi0739 & ~w9463;
assign w9466 = ~w9464 & ~w9465;
assign w9467 = ~pi0966 & ~w9466;
assign w9468 = ~pi1114 & w9463;
assign w9469 = pi0741 & ~w9463;
assign w9470 = ~w9468 & ~w9469;
assign w9471 = ~pi0966 & ~w9470;
assign w9472 = ~pi1112 & w9463;
assign w9473 = pi0742 & ~w9463;
assign w9474 = ~w9472 & ~w9473;
assign w9475 = ~pi0966 & ~w9474;
assign w9476 = ~pi1109 & w9463;
assign w9477 = ~pi0743 & ~w9463;
assign w9478 = ~w9476 & ~w9477;
assign w9479 = ~pi0966 & ~w9478;
assign w9480 = ~pi1131 & w9463;
assign w9481 = pi0744 & ~w9463;
assign w9482 = ~w9480 & ~w9481;
assign w9483 = ~pi0966 & ~w9482;
assign w9484 = ~pi1111 & w9463;
assign w9485 = pi0745 & ~w9463;
assign w9486 = ~w9484 & ~w9485;
assign w9487 = ~pi0966 & ~w9486;
assign w9488 = ~pi1104 & w9463;
assign w9489 = ~pi0746 & ~w9463;
assign w9490 = ~w9488 & ~w9489;
assign w9491 = ~pi0966 & ~w9490;
assign w9492 = pi0773 & w9395;
assign w9493 = pi0747 & ~w9492;
assign w9494 = ~pi0747 & pi0988;
assign w9495 = pi0773 & ~pi0945;
assign w9496 = w9494 & w9495;
assign w9497 = ~w9493 & ~w9496;
assign w9498 = ~w9321 & ~w9497;
assign w9499 = ~pi1106 & w9463;
assign w9500 = ~pi0748 & ~w9463;
assign w9501 = ~w9499 & ~w9500;
assign w9502 = ~pi0966 & ~w9501;
assign w9503 = ~pi1105 & w9463;
assign w9504 = ~pi0749 & ~w9463;
assign w9505 = ~w9503 & ~w9504;
assign w9506 = ~pi0966 & ~w9505;
assign w9507 = ~pi1130 & w9463;
assign w9508 = pi0750 & ~w9463;
assign w9509 = ~w9507 & ~w9508;
assign w9510 = ~pi0966 & ~w9509;
assign w9511 = ~pi1123 & w9463;
assign w9512 = pi0751 & ~w9463;
assign w9513 = ~w9511 & ~w9512;
assign w9514 = ~pi0966 & ~w9513;
assign w9515 = ~pi1124 & w9463;
assign w9516 = pi0752 & ~w9463;
assign w9517 = ~w9515 & ~w9516;
assign w9518 = ~pi0966 & ~w9517;
assign w9519 = ~pi1117 & w9463;
assign w9520 = pi0753 & ~w9463;
assign w9521 = ~w9519 & ~w9520;
assign w9522 = ~pi0966 & ~w9521;
assign w9523 = ~pi1118 & w9463;
assign w9524 = pi0754 & ~w9463;
assign w9525 = ~w9523 & ~w9524;
assign w9526 = ~pi0966 & ~w9525;
assign w9527 = ~pi1120 & w9463;
assign w9528 = pi0755 & ~w9463;
assign w9529 = ~w9527 & ~w9528;
assign w9530 = ~pi0966 & ~w9529;
assign w9531 = ~pi1119 & w9463;
assign w9532 = pi0756 & ~w9463;
assign w9533 = ~w9531 & ~w9532;
assign w9534 = ~pi0966 & ~w9533;
assign w9535 = ~pi1113 & w9463;
assign w9536 = pi0757 & ~w9463;
assign w9537 = ~w9535 & ~w9536;
assign w9538 = ~pi0966 & ~w9537;
assign w9539 = ~pi1101 & w9463;
assign w9540 = ~pi0758 & ~w9463;
assign w9541 = ~w9539 & ~w9540;
assign w9542 = ~pi0966 & ~w9541;
assign w9543 = ~pi1100 & w9463;
assign w9544 = ~pi0759 & ~w9463;
assign w9545 = ~w9543 & ~w9544;
assign w9546 = ~pi0966 & ~w9545;
assign w9547 = ~pi1115 & w9463;
assign w9548 = pi0760 & ~w9463;
assign w9549 = ~w9547 & ~w9548;
assign w9550 = ~pi0966 & ~w9549;
assign w9551 = ~pi1121 & w9463;
assign w9552 = pi0761 & ~w9463;
assign w9553 = ~w9551 & ~w9552;
assign w9554 = ~pi0966 & ~w9553;
assign w9555 = ~pi1129 & w9463;
assign w9556 = pi0762 & ~w9463;
assign w9557 = ~w9555 & ~w9556;
assign w9558 = ~pi0966 & ~w9557;
assign w9559 = ~pi1103 & w9463;
assign w9560 = ~pi0763 & ~w9463;
assign w9561 = ~w9559 & ~w9560;
assign w9562 = ~pi0966 & ~w9561;
assign w9563 = ~pi1107 & w9463;
assign w9564 = ~pi0764 & ~w9463;
assign w9565 = ~w9563 & ~w9564;
assign w9566 = ~pi0966 & ~w9565;
assign w9567 = pi0765 & pi0945;
assign w9568 = ~pi0765 & ~pi0945;
assign w9569 = ~w9567 & ~w9568;
assign w9570 = ~pi0795 & ~pi0816;
assign w9571 = ~pi0794 & w9570;
assign w9572 = ~pi0721 & ~pi0747;
assign w9573 = ~pi0765 & w9572;
assign w9574 = ~pi0771 & w9573;
assign w9575 = ~pi0773 & w9574;
assign w9576 = w9571 & w9575;
assign w9577 = w9321 & ~w9576;
assign w9578 = ~w9569 & ~w9577;
assign w9579 = ~pi1110 & w9463;
assign w9580 = ~pi0766 & ~w9463;
assign w9581 = ~w9579 & ~w9580;
assign w9582 = ~pi0966 & ~w9581;
assign w9583 = ~pi1116 & w9463;
assign w9584 = pi0767 & ~w9463;
assign w9585 = ~w9583 & ~w9584;
assign w9586 = ~pi0966 & ~w9585;
assign w9587 = ~pi1125 & w9463;
assign w9588 = pi0768 & ~w9463;
assign w9589 = ~w9587 & ~w9588;
assign w9590 = ~pi0966 & ~w9589;
assign w9591 = ~pi0769 & w9285;
assign w9592 = pi0769 & ~w9285;
assign w9593 = ~w9591 & ~w9592;
assign w9594 = ~w9321 & ~w9593;
assign w9595 = ~pi1126 & w9463;
assign w9596 = pi0770 & ~w9463;
assign w9597 = ~w9595 & ~w9596;
assign w9598 = ~pi0966 & ~w9597;
assign w9599 = ~pi0945 & pi0987;
assign w9600 = pi0771 & pi0945;
assign w9601 = ~w9599 & ~w9600;
assign w9602 = ~w9577 & ~w9601;
assign w9603 = ~pi1102 & w9463;
assign w9604 = ~pi0772 & ~w9463;
assign w9605 = ~w9603 & ~w9604;
assign w9606 = ~pi0966 & ~w9605;
assign w9607 = ~pi0773 & pi0988;
assign w9608 = ~pi0945 & w9607;
assign w9609 = pi0773 & ~w9395;
assign w9610 = ~w9608 & ~w9609;
assign w9611 = ~w9577 & ~w9610;
assign w9612 = ~pi1127 & w9463;
assign w9613 = pi0774 & ~w9463;
assign w9614 = ~w9612 & ~w9613;
assign w9615 = ~pi0966 & ~w9614;
assign w9616 = pi0765 & w9281;
assign w9617 = pi0771 & w9616;
assign w9618 = pi0773 & w9617;
assign w9619 = ~pi0945 & w9618;
assign w9620 = ~pi0775 & w9619;
assign w9621 = pi0775 & ~w9619;
assign w9622 = ~w9620 & ~w9621;
assign w9623 = ~w9321 & ~w9622;
assign w9624 = ~pi1128 & w9463;
assign w9625 = pi0776 & ~w9463;
assign w9626 = ~w9624 & ~w9625;
assign w9627 = ~pi0966 & ~w9626;
assign w9628 = ~pi1122 & w9463;
assign w9629 = pi0777 & ~w9463;
assign w9630 = ~w9628 & ~w9629;
assign w9631 = ~pi0966 & ~w9630;
assign w9632 = pi0832 & pi0956;
assign w9633 = ~pi0968 & w9632;
assign w9634 = ~pi1046 & w9633;
assign w9635 = ~pi1083 & w9634;
assign w9636 = pi1085 & w9635;
assign w9637 = pi1100 & w9636;
assign w9638 = pi0778 & ~w9636;
assign w9639 = ~w9637 & ~w9638;
assign w9640 = pi0779 & ~w7866;
assign w9641 = pi0780 & ~w7779;
assign w9642 = pi1101 & w9636;
assign w9643 = pi0781 & ~w9636;
assign w9644 = ~w9642 & ~w9643;
assign w9645 = ~pi0299 & pi0983;
assign w9646 = ~pi0979 & ~pi0984;
assign w9647 = ~w9645 & ~w9646;
assign w9648 = ~w7778 & w9647;
assign w9649 = pi1109 & w9636;
assign w9650 = pi0783 & ~w9636;
assign w9651 = ~w9649 & ~w9650;
assign w9652 = pi1110 & w9636;
assign w9653 = pi0784 & ~w9636;
assign w9654 = ~w9652 & ~w9653;
assign w9655 = pi1102 & w9636;
assign w9656 = pi0785 & ~w9636;
assign w9657 = ~w9655 & ~w9656;
assign w9658 = ~pi0786 & pi0954;
assign w9659 = ~pi0024 & ~pi0954;
assign w9660 = ~w9658 & ~w9659;
assign w9661 = pi1104 & w9636;
assign w9662 = pi0787 & ~w9636;
assign w9663 = ~w9661 & ~w9662;
assign w9664 = pi1105 & w9636;
assign w9665 = pi0788 & ~w9636;
assign w9666 = ~w9664 & ~w9665;
assign w9667 = pi1106 & w9636;
assign w9668 = pi0789 & ~w9636;
assign w9669 = ~w9667 & ~w9668;
assign w9670 = pi1107 & w9636;
assign w9671 = pi0790 & ~w9636;
assign w9672 = ~w9670 & ~w9671;
assign w9673 = pi1108 & w9636;
assign w9674 = pi0791 & ~w9636;
assign w9675 = ~w9673 & ~w9674;
assign w9676 = pi1103 & w9636;
assign w9677 = pi0792 & ~w9636;
assign w9678 = ~w9676 & ~w9677;
assign w9679 = pi0968 & w9632;
assign w9680 = ~pi1046 & w9679;
assign w9681 = ~pi1083 & w9680;
assign w9682 = pi1085 & w9681;
assign w9683 = pi1130 & w9682;
assign w9684 = pi0794 & ~w9682;
assign w9685 = ~w9683 & ~w9684;
assign w9686 = pi1128 & w9682;
assign w9687 = pi0795 & ~w9682;
assign w9688 = ~w9686 & ~w9687;
assign w9689 = pi0264 & pi0279;
assign w9690 = pi0278 & w9689;
assign w9691 = w8063 & w8067;
assign w9692 = w9690 & w9691;
assign w9693 = pi0278 & pi0279;
assign w9694 = ~pi0277 & w9693;
assign w9695 = ~pi0270 & w8063;
assign w9696 = w9694 & w9695;
assign w9697 = ~pi0264 & ~w9696;
assign w9698 = ~w9692 & ~w9697;
assign w9699 = pi1124 & w9682;
assign w9700 = pi0798 & ~w9682;
assign w9701 = ~w9699 & ~w9700;
assign w9702 = pi1107 & w9682;
assign w9703 = ~pi0799 & ~w9682;
assign w9704 = ~w9702 & ~w9703;
assign w9705 = pi1125 & w9682;
assign w9706 = pi0800 & ~w9682;
assign w9707 = ~w9705 & ~w9706;
assign w9708 = pi1126 & w9682;
assign w9709 = pi0801 & ~w9682;
assign w9710 = ~w9708 & ~w9709;
assign w9711 = ~pi0265 & w8069;
assign w9712 = ~pi0270 & w9711;
assign w9713 = ~pi0274 & w9712;
assign w9714 = ~pi0277 & w9713;
assign w9715 = pi1106 & w9682;
assign w9716 = ~pi0803 & ~w9682;
assign w9717 = ~w9715 & ~w9716;
assign w9718 = pi1109 & w9682;
assign w9719 = pi0804 & ~w9682;
assign w9720 = ~w9718 & ~w9719;
assign w9721 = pi0270 & w8064;
assign w9722 = ~pi0270 & ~w8064;
assign w9723 = ~w9721 & ~w9722;
assign w9724 = pi1127 & w9682;
assign w9725 = pi0807 & ~w9682;
assign w9726 = ~w9724 & ~w9725;
assign w9727 = pi1101 & w9682;
assign w9728 = pi0808 & ~w9682;
assign w9729 = ~w9727 & ~w9728;
assign w9730 = pi1103 & w9682;
assign w9731 = ~pi0809 & ~w9682;
assign w9732 = ~w9730 & ~w9731;
assign w9733 = pi1108 & w9682;
assign w9734 = pi0810 & ~w9682;
assign w9735 = ~w9733 & ~w9734;
assign w9736 = pi1102 & w9682;
assign w9737 = pi0811 & ~w9682;
assign w9738 = ~w9736 & ~w9737;
assign w9739 = pi1104 & w9682;
assign w9740 = ~pi0812 & ~w9682;
assign w9741 = ~w9739 & ~w9740;
assign w9742 = pi1131 & w9682;
assign w9743 = pi0813 & ~w9682;
assign w9744 = ~w9742 & ~w9743;
assign w9745 = pi1105 & w9682;
assign w9746 = ~pi0814 & ~w9682;
assign w9747 = ~w9745 & ~w9746;
assign w9748 = pi1110 & w9682;
assign w9749 = pi0815 & ~w9682;
assign w9750 = ~w9748 & ~w9749;
assign w9751 = pi1129 & w9682;
assign w9752 = pi0816 & ~w9682;
assign w9753 = ~w9751 & ~w9752;
assign w9754 = pi0269 & pi0992;
assign w9755 = pi0266 & ~pi0280;
assign w9756 = w9754 & w9755;
assign w9757 = ~pi0280 & pi0992;
assign w9758 = pi0266 & w9757;
assign w9759 = ~pi0269 & ~w9758;
assign w9760 = ~w9756 & ~w9759;
assign w9761 = ~pi0080 & pi0818;
assign w9762 = ~pi0031 & w9761;
assign w9763 = ~w4065 & ~w9762;
assign w9764 = pi0265 & ~pi0277;
assign w9765 = ~pi0270 & w9764;
assign w9766 = w8069 & w9765;
assign w9767 = w8067 & w8069;
assign w9768 = ~pi0265 & ~w9767;
assign w9769 = ~w9766 & ~w9768;
assign w9770 = ~pi0270 & pi0277;
assign w9771 = w8064 & w9770;
assign w9772 = ~pi0270 & w8064;
assign w9773 = ~pi0277 & ~w9772;
assign w9774 = ~w9771 & ~w9773;
assign w9775 = ~pi0811 & ~pi0893;
assign w9776 = pi1093 & w2045;
assign w9777 = pi0982 & ~w9776;
assign w9778 = ~pi1091 & ~w9777;
assign w9779 = pi1093 & w449;
assign w9780 = ~pi0982 & ~w9779;
assign w9781 = ~w9778 & ~w9780;
assign w9782 = w1280 & ~w9781;
assign w9783 = pi0123 & ~pi0222;
assign w9784 = w4192 & w9783;
assign w9785 = pi1128 & ~pi1129;
assign w9786 = ~pi1128 & pi1129;
assign w9787 = ~w9785 & ~w9786;
assign w9788 = ~pi1124 & pi1125;
assign w9789 = pi1124 & ~pi1125;
assign w9790 = ~w9788 & ~w9789;
assign w9791 = ~pi1126 & ~pi1127;
assign w9792 = pi1126 & pi1127;
assign w9793 = ~w9791 & ~w9792;
assign w9794 = ~w9790 & ~w9793;
assign w9795 = pi1124 & pi1125;
assign w9796 = ~pi1124 & ~pi1125;
assign w9797 = ~w9795 & ~w9796;
assign w9798 = pi1126 & ~pi1127;
assign w9799 = ~pi1126 & pi1127;
assign w9800 = ~w9798 & ~w9799;
assign w9801 = ~w9797 & ~w9800;
assign w9802 = ~w9794 & ~w9801;
assign w9803 = ~w9787 & ~w9802;
assign w9804 = pi1128 & pi1129;
assign w9805 = ~pi1128 & ~pi1129;
assign w9806 = ~w9804 & ~w9805;
assign w9807 = w9802 & ~w9806;
assign w9808 = ~w9803 & ~w9807;
assign w9809 = pi1130 & pi1131;
assign w9810 = ~pi1130 & ~pi1131;
assign w9811 = ~w9809 & ~w9810;
assign w9812 = ~w9808 & ~w9811;
assign w9813 = ~w9802 & ~w9806;
assign w9814 = ~w9787 & w9802;
assign w9815 = ~w9813 & ~w9814;
assign w9816 = pi1130 & ~pi1131;
assign w9817 = ~pi1130 & pi1131;
assign w9818 = ~w9816 & ~w9817;
assign w9819 = ~w9815 & ~w9818;
assign w9820 = ~w9812 & ~w9819;
assign w9821 = ~w9784 & w9820;
assign w9822 = ~pi0825 & w4192;
assign w9823 = w9783 & w9822;
assign w9824 = ~w9821 & ~w9823;
assign w9825 = pi1120 & ~pi1121;
assign w9826 = ~pi1120 & pi1121;
assign w9827 = ~w9825 & ~w9826;
assign w9828 = ~pi1116 & pi1117;
assign w9829 = pi1116 & ~pi1117;
assign w9830 = ~w9828 & ~w9829;
assign w9831 = ~pi1118 & ~pi1119;
assign w9832 = pi1118 & pi1119;
assign w9833 = ~w9831 & ~w9832;
assign w9834 = ~w9830 & ~w9833;
assign w9835 = pi1116 & pi1117;
assign w9836 = ~pi1116 & ~pi1117;
assign w9837 = ~w9835 & ~w9836;
assign w9838 = pi1118 & ~pi1119;
assign w9839 = ~pi1118 & pi1119;
assign w9840 = ~w9838 & ~w9839;
assign w9841 = ~w9837 & ~w9840;
assign w9842 = ~w9834 & ~w9841;
assign w9843 = ~w9827 & ~w9842;
assign w9844 = pi1120 & pi1121;
assign w9845 = ~pi1120 & ~pi1121;
assign w9846 = ~w9844 & ~w9845;
assign w9847 = w9842 & ~w9846;
assign w9848 = ~w9843 & ~w9847;
assign w9849 = pi1122 & pi1123;
assign w9850 = ~pi1122 & ~pi1123;
assign w9851 = ~w9849 & ~w9850;
assign w9852 = ~w9848 & ~w9851;
assign w9853 = ~w9842 & ~w9846;
assign w9854 = ~w9827 & w9842;
assign w9855 = ~w9853 & ~w9854;
assign w9856 = pi1122 & ~pi1123;
assign w9857 = ~pi1122 & pi1123;
assign w9858 = ~w9856 & ~w9857;
assign w9859 = ~w9855 & ~w9858;
assign w9860 = ~w9852 & ~w9859;
assign w9861 = ~w9784 & w9860;
assign w9862 = ~pi0826 & w4192;
assign w9863 = w9783 & w9862;
assign w9864 = ~w9861 & ~w9863;
assign w9865 = pi1104 & ~pi1105;
assign w9866 = ~pi1104 & pi1105;
assign w9867 = ~w9865 & ~w9866;
assign w9868 = ~pi1100 & pi1101;
assign w9869 = pi1100 & ~pi1101;
assign w9870 = ~w9868 & ~w9869;
assign w9871 = ~pi1102 & ~pi1103;
assign w9872 = pi1102 & pi1103;
assign w9873 = ~w9871 & ~w9872;
assign w9874 = ~w9870 & ~w9873;
assign w9875 = pi1100 & pi1101;
assign w9876 = ~pi1100 & ~pi1101;
assign w9877 = ~w9875 & ~w9876;
assign w9878 = pi1102 & ~pi1103;
assign w9879 = ~pi1102 & pi1103;
assign w9880 = ~w9878 & ~w9879;
assign w9881 = ~w9877 & ~w9880;
assign w9882 = ~w9874 & ~w9881;
assign w9883 = ~w9867 & ~w9882;
assign w9884 = pi1104 & pi1105;
assign w9885 = ~pi1104 & ~pi1105;
assign w9886 = ~w9884 & ~w9885;
assign w9887 = w9882 & ~w9886;
assign w9888 = ~w9883 & ~w9887;
assign w9889 = pi1106 & pi1107;
assign w9890 = ~pi1106 & ~pi1107;
assign w9891 = ~w9889 & ~w9890;
assign w9892 = ~w9888 & ~w9891;
assign w9893 = ~w9882 & ~w9886;
assign w9894 = ~w9867 & w9882;
assign w9895 = ~w9893 & ~w9894;
assign w9896 = pi1106 & ~pi1107;
assign w9897 = ~pi1106 & pi1107;
assign w9898 = ~w9896 & ~w9897;
assign w9899 = ~w9895 & ~w9898;
assign w9900 = ~w9892 & ~w9899;
assign w9901 = ~w9784 & w9900;
assign w9902 = ~pi0827 & w4192;
assign w9903 = w9783 & w9902;
assign w9904 = ~w9901 & ~w9903;
assign w9905 = pi1112 & ~pi1113;
assign w9906 = ~pi1112 & pi1113;
assign w9907 = ~w9905 & ~w9906;
assign w9908 = ~pi1108 & pi1109;
assign w9909 = pi1108 & ~pi1109;
assign w9910 = ~w9908 & ~w9909;
assign w9911 = ~pi1110 & ~pi1111;
assign w9912 = pi1110 & pi1111;
assign w9913 = ~w9911 & ~w9912;
assign w9914 = ~w9910 & ~w9913;
assign w9915 = pi1108 & pi1109;
assign w9916 = ~pi1108 & ~pi1109;
assign w9917 = ~w9915 & ~w9916;
assign w9918 = pi1110 & ~pi1111;
assign w9919 = ~pi1110 & pi1111;
assign w9920 = ~w9918 & ~w9919;
assign w9921 = ~w9917 & ~w9920;
assign w9922 = ~w9914 & ~w9921;
assign w9923 = ~w9907 & ~w9922;
assign w9924 = pi1112 & pi1113;
assign w9925 = ~pi1112 & ~pi1113;
assign w9926 = ~w9924 & ~w9925;
assign w9927 = w9922 & ~w9926;
assign w9928 = ~w9923 & ~w9927;
assign w9929 = pi1114 & pi1115;
assign w9930 = ~pi1114 & ~pi1115;
assign w9931 = ~w9929 & ~w9930;
assign w9932 = ~w9928 & ~w9931;
assign w9933 = ~w9922 & ~w9926;
assign w9934 = ~w9907 & w9922;
assign w9935 = ~w9933 & ~w9934;
assign w9936 = pi1114 & ~pi1115;
assign w9937 = ~pi1114 & pi1115;
assign w9938 = ~w9936 & ~w9937;
assign w9939 = ~w9935 & ~w9938;
assign w9940 = ~w9932 & ~w9939;
assign w9941 = ~w9784 & w9940;
assign w9942 = ~pi0828 & w4192;
assign w9943 = w9783 & w9942;
assign w9944 = ~w9941 & ~w9943;
assign w9945 = w1234 & w2045;
assign w9946 = pi0951 & ~w9945;
assign w9947 = pi1092 & ~w9946;
assign w9948 = ~pi0280 & pi0281;
assign w9949 = pi0279 & w9948;
assign w9950 = ~pi0269 & pi0278;
assign w9951 = pi0266 & w9950;
assign w9952 = w9949 & w9951;
assign w9953 = pi0279 & ~pi0280;
assign w9954 = pi0278 & w9953;
assign w9955 = w8060 & w9954;
assign w9956 = ~pi0281 & ~w9955;
assign w9957 = ~w9952 & ~w9956;
assign w9958 = ~pi0832 & w1475;
assign w9959 = pi1091 & w9958;
assign w9960 = pi1161 & w9959;
assign w9961 = pi1162 & w9960;
assign w9962 = ~pi1163 & w9961;
assign w9963 = pi1091 & w1475;
assign w9964 = pi0833 & ~w1475;
assign w9965 = ~w9963 & ~w9964;
assign w9966 = pi0946 & w1475;
assign w9967 = pi0282 & pi0992;
assign w9968 = ~pi0281 & w9967;
assign w9969 = ~pi0269 & ~pi0280;
assign w9970 = pi0266 & w9969;
assign w9971 = w9968 & w9970;
assign w9972 = ~pi0281 & pi0992;
assign w9973 = ~pi0280 & w9972;
assign w9974 = w8060 & w9973;
assign w9975 = ~pi0282 & ~w9974;
assign w9976 = ~w9971 & ~w9975;
assign w9977 = ~pi0955 & pi1049;
assign w9978 = pi0837 & pi0955;
assign w9979 = ~w9977 & ~w9978;
assign w9980 = ~pi0955 & pi1047;
assign w9981 = pi0838 & pi0955;
assign w9982 = ~w9980 & ~w9981;
assign w9983 = ~pi0955 & pi1074;
assign w9984 = pi0839 & pi0955;
assign w9985 = ~w9983 & ~w9984;
assign w9986 = pi1196 & w1475;
assign w9987 = pi0840 & ~w1475;
assign w9988 = ~w9986 & ~w9987;
assign w9989 = ~pi0034 & w2674;
assign w9990 = ~pi0955 & pi1035;
assign w9991 = pi0842 & pi0955;
assign w9992 = ~w9990 & ~w9991;
assign w9993 = ~pi0955 & pi1079;
assign w9994 = pi0843 & pi0955;
assign w9995 = ~w9993 & ~w9994;
assign w9996 = ~pi0955 & pi1078;
assign w9997 = pi0844 & pi0955;
assign w9998 = ~w9996 & ~w9997;
assign w9999 = ~pi0955 & pi1043;
assign w10000 = pi0845 & pi0955;
assign w10001 = ~w9999 & ~w10000;
assign w10002 = pi1134 & ~w5939;
assign w10003 = pi0846 & w5939;
assign w10004 = ~w10002 & ~w10003;
assign w10005 = ~pi0955 & pi1055;
assign w10006 = pi0847 & pi0955;
assign w10007 = ~w10005 & ~w10006;
assign w10008 = ~pi0955 & pi1039;
assign w10009 = pi0848 & pi0955;
assign w10010 = ~w10008 & ~w10009;
assign w10011 = pi1198 & w1475;
assign w10012 = pi0849 & ~w1475;
assign w10013 = ~w10011 & ~w10012;
assign w10014 = ~pi0955 & pi1048;
assign w10015 = pi0850 & pi0955;
assign w10016 = ~w10014 & ~w10015;
assign w10017 = ~pi0955 & pi1045;
assign w10018 = pi0851 & pi0955;
assign w10019 = ~w10017 & ~w10018;
assign w10020 = ~pi0955 & pi1062;
assign w10021 = pi0852 & pi0955;
assign w10022 = ~w10020 & ~w10021;
assign w10023 = ~pi0955 & pi1080;
assign w10024 = pi0853 & pi0955;
assign w10025 = ~w10023 & ~w10024;
assign w10026 = ~pi0955 & pi1051;
assign w10027 = pi0854 & pi0955;
assign w10028 = ~w10026 & ~w10027;
assign w10029 = ~pi0955 & pi1065;
assign w10030 = pi0855 & pi0955;
assign w10031 = ~w10029 & ~w10030;
assign w10032 = ~pi0955 & pi1067;
assign w10033 = pi0856 & pi0955;
assign w10034 = ~w10032 & ~w10033;
assign w10035 = ~pi0955 & pi1058;
assign w10036 = pi0857 & pi0955;
assign w10037 = ~w10035 & ~w10036;
assign w10038 = ~pi0955 & pi1087;
assign w10039 = pi0858 & pi0955;
assign w10040 = ~w10038 & ~w10039;
assign w10041 = ~pi0955 & pi1070;
assign w10042 = pi0859 & pi0955;
assign w10043 = ~w10041 & ~w10042;
assign w10044 = ~pi0955 & pi1076;
assign w10045 = pi0860 & pi0955;
assign w10046 = ~w10044 & ~w10045;
assign w10047 = pi1141 & ~w5939;
assign w10048 = pi0861 & w5939;
assign w10049 = ~w10047 & ~w10048;
assign w10050 = pi1139 & ~w5939;
assign w10051 = pi0862 & w5939;
assign w10052 = ~w10050 & ~w10051;
assign w10053 = pi1199 & w1475;
assign w10054 = pi0863 & ~w1475;
assign w10055 = ~w10053 & ~w10054;
assign w10056 = pi1197 & w1475;
assign w10057 = pi0864 & ~w1475;
assign w10058 = ~w10056 & ~w10057;
assign w10059 = ~pi0955 & pi1040;
assign w10060 = pi0865 & pi0955;
assign w10061 = ~w10059 & ~w10060;
assign w10062 = ~pi0955 & pi1053;
assign w10063 = pi0866 & pi0955;
assign w10064 = ~w10062 & ~w10063;
assign w10065 = ~pi0955 & pi1057;
assign w10066 = pi0867 & pi0955;
assign w10067 = ~w10065 & ~w10066;
assign w10068 = ~pi0955 & pi1063;
assign w10069 = pi0868 & pi0955;
assign w10070 = ~w10068 & ~w10069;
assign w10071 = pi1140 & ~w5939;
assign w10072 = pi0869 & w5939;
assign w10073 = ~w10071 & ~w10072;
assign w10074 = ~pi0955 & pi1069;
assign w10075 = pi0870 & pi0955;
assign w10076 = ~w10074 & ~w10075;
assign w10077 = ~pi0955 & pi1072;
assign w10078 = pi0871 & pi0955;
assign w10079 = ~w10077 & ~w10078;
assign w10080 = ~pi0955 & pi1084;
assign w10081 = pi0872 & pi0955;
assign w10082 = ~w10080 & ~w10081;
assign w10083 = ~pi0955 & pi1044;
assign w10084 = pi0873 & pi0955;
assign w10085 = ~w10083 & ~w10084;
assign w10086 = ~pi0955 & pi1036;
assign w10087 = pi0874 & pi0955;
assign w10088 = ~w10086 & ~w10087;
assign w10089 = pi1136 & ~w5939;
assign w10090 = pi0875 & w5939;
assign w10091 = ~w10089 & ~w10090;
assign w10092 = ~pi0955 & pi1037;
assign w10093 = pi0876 & pi0955;
assign w10094 = ~w10092 & ~w10093;
assign w10095 = pi1138 & ~w5939;
assign w10096 = pi0877 & w5939;
assign w10097 = ~w10095 & ~w10096;
assign w10098 = pi1137 & ~w5939;
assign w10099 = pi0878 & w5939;
assign w10100 = ~w10098 & ~w10099;
assign w10101 = pi1135 & ~w5939;
assign w10102 = pi0879 & w5939;
assign w10103 = ~w10101 & ~w10102;
assign w10104 = ~pi0955 & pi1081;
assign w10105 = pi0880 & pi0955;
assign w10106 = ~w10104 & ~w10105;
assign w10107 = ~pi0955 & pi1059;
assign w10108 = pi0881 & pi0955;
assign w10109 = ~w10107 & ~w10108;
assign w10110 = pi0123 & ~pi0883;
assign w10111 = ~pi0222 & w4192;
assign w10112 = w10110 & w10111;
assign w10113 = pi0123 & w10111;
assign w10114 = pi1107 & ~w10113;
assign w10115 = ~w10112 & ~w10114;
assign w10116 = pi0123 & ~pi0884;
assign w10117 = w10111 & w10116;
assign w10118 = pi1124 & ~w10113;
assign w10119 = ~w10117 & ~w10118;
assign w10120 = pi0123 & ~pi0885;
assign w10121 = w10111 & w10120;
assign w10122 = pi1125 & ~w10113;
assign w10123 = ~w10121 & ~w10122;
assign w10124 = pi0123 & ~pi0886;
assign w10125 = w10111 & w10124;
assign w10126 = pi1109 & ~w10113;
assign w10127 = ~w10125 & ~w10126;
assign w10128 = pi0123 & ~pi0887;
assign w10129 = w10111 & w10128;
assign w10130 = pi1100 & ~w10113;
assign w10131 = ~w10129 & ~w10130;
assign w10132 = pi0123 & ~pi0888;
assign w10133 = w10111 & w10132;
assign w10134 = pi1120 & ~w10113;
assign w10135 = ~w10133 & ~w10134;
assign w10136 = pi0123 & ~pi0889;
assign w10137 = w10111 & w10136;
assign w10138 = pi1103 & ~w10113;
assign w10139 = ~w10137 & ~w10138;
assign w10140 = pi0123 & ~pi0890;
assign w10141 = w10111 & w10140;
assign w10142 = pi1126 & ~w10113;
assign w10143 = ~w10141 & ~w10142;
assign w10144 = pi0123 & ~pi0891;
assign w10145 = w10111 & w10144;
assign w10146 = pi1116 & ~w10113;
assign w10147 = ~w10145 & ~w10146;
assign w10148 = pi0123 & ~pi0892;
assign w10149 = w10111 & w10148;
assign w10150 = pi1101 & ~w10113;
assign w10151 = ~w10149 & ~w10150;
assign w10152 = pi0123 & ~pi0894;
assign w10153 = w10111 & w10152;
assign w10154 = pi1119 & ~w10113;
assign w10155 = ~w10153 & ~w10154;
assign w10156 = pi0123 & ~pi0895;
assign w10157 = w10111 & w10156;
assign w10158 = pi1113 & ~w10113;
assign w10159 = ~w10157 & ~w10158;
assign w10160 = pi0123 & ~pi0896;
assign w10161 = w10111 & w10160;
assign w10162 = pi1118 & ~w10113;
assign w10163 = ~w10161 & ~w10162;
assign w10164 = pi0123 & ~pi0898;
assign w10165 = w10111 & w10164;
assign w10166 = pi1129 & ~w10113;
assign w10167 = ~w10165 & ~w10166;
assign w10168 = pi0123 & ~pi0899;
assign w10169 = w10111 & w10168;
assign w10170 = pi1115 & ~w10113;
assign w10171 = ~w10169 & ~w10170;
assign w10172 = pi0123 & ~pi0900;
assign w10173 = w10111 & w10172;
assign w10174 = pi1110 & ~w10113;
assign w10175 = ~w10173 & ~w10174;
assign w10176 = pi0123 & ~pi0902;
assign w10177 = w10111 & w10176;
assign w10178 = pi1111 & ~w10113;
assign w10179 = ~w10177 & ~w10178;
assign w10180 = pi0123 & ~pi0903;
assign w10181 = w10111 & w10180;
assign w10182 = pi1121 & ~w10113;
assign w10183 = ~w10181 & ~w10182;
assign w10184 = pi0123 & ~pi0904;
assign w10185 = w10111 & w10184;
assign w10186 = pi1127 & ~w10113;
assign w10187 = ~w10185 & ~w10186;
assign w10188 = pi0123 & ~pi0905;
assign w10189 = w10111 & w10188;
assign w10190 = pi1131 & ~w10113;
assign w10191 = ~w10189 & ~w10190;
assign w10192 = pi0123 & ~pi0906;
assign w10193 = w10111 & w10192;
assign w10194 = pi1128 & ~w10113;
assign w10195 = ~w10193 & ~w10194;
assign w10196 = ~pi0782 & pi0907;
assign w10197 = ~pi0598 & pi0979;
assign w10198 = ~pi0615 & w10197;
assign w10199 = ~pi0624 & ~pi0979;
assign w10200 = pi0604 & w10199;
assign w10201 = ~w10198 & ~w10200;
assign w10202 = pi0782 & ~w10201;
assign w10203 = ~w10196 & ~w10202;
assign w10204 = pi0123 & ~pi0908;
assign w10205 = w10111 & w10204;
assign w10206 = pi1122 & ~w10113;
assign w10207 = ~w10205 & ~w10206;
assign w10208 = pi0123 & ~pi0909;
assign w10209 = w10111 & w10208;
assign w10210 = pi1105 & ~w10113;
assign w10211 = ~w10209 & ~w10210;
assign w10212 = pi0123 & ~pi0910;
assign w10213 = w10111 & w10212;
assign w10214 = pi1117 & ~w10113;
assign w10215 = ~w10213 & ~w10214;
assign w10216 = pi0123 & ~pi0911;
assign w10217 = w10111 & w10216;
assign w10218 = pi1130 & ~w10113;
assign w10219 = ~w10217 & ~w10218;
assign w10220 = pi0123 & ~pi0912;
assign w10221 = w10111 & w10220;
assign w10222 = pi1114 & ~w10113;
assign w10223 = ~w10221 & ~w10222;
assign w10224 = pi0123 & ~pi0913;
assign w10225 = w10111 & w10224;
assign w10226 = pi1106 & ~w10113;
assign w10227 = ~w10225 & ~w10226;
assign w10228 = pi0280 & pi0992;
assign w10229 = pi0266 & w10228;
assign w10230 = pi0266 & pi0992;
assign w10231 = ~pi0280 & ~w10230;
assign w10232 = ~w10229 & ~w10231;
assign w10233 = pi0123 & ~pi0915;
assign w10234 = w10111 & w10233;
assign w10235 = pi1108 & ~w10113;
assign w10236 = ~w10234 & ~w10235;
assign w10237 = pi0123 & ~pi0916;
assign w10238 = w10111 & w10237;
assign w10239 = pi1123 & ~w10113;
assign w10240 = ~w10238 & ~w10239;
assign w10241 = pi0123 & ~pi0917;
assign w10242 = w10111 & w10241;
assign w10243 = pi1112 & ~w10113;
assign w10244 = ~w10242 & ~w10243;
assign w10245 = pi0123 & ~pi0918;
assign w10246 = w10111 & w10245;
assign w10247 = pi1104 & ~w10113;
assign w10248 = ~w10246 & ~w10247;
assign w10249 = pi0123 & ~pi0919;
assign w10250 = w10111 & w10249;
assign w10251 = pi1102 & ~w10113;
assign w10252 = ~w10250 & ~w10251;
assign w10253 = pi1093 & pi1139;
assign w10254 = pi0920 & ~pi1093;
assign w10255 = ~w10253 & ~w10254;
assign w10256 = pi1093 & pi1140;
assign w10257 = pi0921 & ~pi1093;
assign w10258 = ~w10256 & ~w10257;
assign w10259 = pi1093 & pi1152;
assign w10260 = pi0922 & ~pi1093;
assign w10261 = ~w10259 & ~w10260;
assign w10262 = pi1093 & pi1154;
assign w10263 = pi0923 & ~pi1093;
assign w10264 = ~w10262 & ~w10263;
assign w10265 = pi0311 & w6331;
assign w10266 = ~pi0312 & w10265;
assign w10267 = pi1093 & pi1155;
assign w10268 = pi0925 & ~pi1093;
assign w10269 = ~w10267 & ~w10268;
assign w10270 = pi1093 & pi1157;
assign w10271 = pi0926 & ~pi1093;
assign w10272 = ~w10270 & ~w10271;
assign w10273 = pi1093 & pi1145;
assign w10274 = pi0927 & ~pi1093;
assign w10275 = ~w10273 & ~w10274;
assign w10276 = pi1093 & pi1136;
assign w10277 = pi0928 & ~pi1093;
assign w10278 = ~w10276 & ~w10277;
assign w10279 = pi1093 & pi1144;
assign w10280 = pi0929 & ~pi1093;
assign w10281 = ~w10279 & ~w10280;
assign w10282 = pi1093 & pi1134;
assign w10283 = pi0930 & ~pi1093;
assign w10284 = ~w10282 & ~w10283;
assign w10285 = pi1093 & pi1150;
assign w10286 = pi0931 & ~pi1093;
assign w10287 = ~w10285 & ~w10286;
assign w10288 = pi1093 & pi1142;
assign w10289 = pi0932 & ~pi1093;
assign w10290 = ~w10288 & ~w10289;
assign w10291 = pi1093 & pi1137;
assign w10292 = pi0933 & ~pi1093;
assign w10293 = ~w10291 & ~w10292;
assign w10294 = pi1093 & pi1147;
assign w10295 = pi0934 & ~pi1093;
assign w10296 = ~w10294 & ~w10295;
assign w10297 = pi1093 & pi1141;
assign w10298 = pi0935 & ~pi1093;
assign w10299 = ~w10297 & ~w10298;
assign w10300 = pi1093 & pi1149;
assign w10301 = pi0936 & ~pi1093;
assign w10302 = ~w10300 & ~w10301;
assign w10303 = pi1093 & pi1148;
assign w10304 = pi0937 & ~pi1093;
assign w10305 = ~w10303 & ~w10304;
assign w10306 = pi1093 & pi1135;
assign w10307 = pi0938 & ~pi1093;
assign w10308 = ~w10306 & ~w10307;
assign w10309 = pi1093 & pi1146;
assign w10310 = pi0939 & ~pi1093;
assign w10311 = ~w10309 & ~w10310;
assign w10312 = pi1093 & pi1138;
assign w10313 = pi0940 & ~pi1093;
assign w10314 = ~w10312 & ~w10313;
assign w10315 = pi1093 & pi1153;
assign w10316 = pi0941 & ~pi1093;
assign w10317 = ~w10315 & ~w10316;
assign w10318 = pi1093 & pi1156;
assign w10319 = pi0942 & ~pi1093;
assign w10320 = ~w10318 & ~w10319;
assign w10321 = pi1093 & pi1151;
assign w10322 = pi0943 & ~pi1093;
assign w10323 = ~w10321 & ~w10322;
assign w10324 = pi1093 & pi1143;
assign w10325 = pi0944 & ~pi1093;
assign w10326 = ~w10324 & ~w10325;
assign w10327 = ~w1249 & ~w1253;
assign w10328 = pi0230 & w1475;
assign w10329 = pi0624 & ~pi0979;
assign w10330 = pi0598 & pi0979;
assign w10331 = ~w10329 & ~w10330;
assign w10332 = pi0782 & ~w10331;
assign w10333 = ~pi0782 & pi0947;
assign w10334 = ~w10332 & ~w10333;
assign w10335 = ~pi0266 & pi0992;
assign w10336 = pi0266 & ~pi0992;
assign w10337 = ~w10335 & ~w10336;
assign w10338 = pi0949 & pi0954;
assign w10339 = ~pi0313 & ~pi0954;
assign w10340 = ~w10338 & ~w10339;
assign w10341 = w449 & w1475;
assign w10342 = pi1091 & w10341;
assign w10343 = pi0829 & ~w450;
assign w10344 = pi1092 & w10343;
assign w10345 = pi0957 & pi1092;
assign w10346 = ~pi0031 & ~w10345;
assign w10347 = ~pi0782 & pi0960;
assign w10348 = ~pi0230 & pi0961;
assign w10349 = ~pi0782 & pi0963;
assign w10350 = ~pi0230 & pi0967;
assign w10351 = ~pi0230 & pi0969;
assign w10352 = ~pi0782 & pi0970;
assign w10353 = ~pi0230 & pi0971;
assign w10354 = ~pi0782 & pi0972;
assign w10355 = ~pi0230 & pi0974;
assign w10356 = ~pi0782 & pi0975;
assign w10357 = ~pi0230 & pi0977;
assign w10358 = ~pi0782 & pi0978;
assign w10359 = ~pi0598 & pi0615;
assign w10360 = pi0824 & pi1092;
assign w10361 = ~pi0604 & ~pi0624;
assign one = 1;
assign po0000 = pi0668;
assign po0001 = pi0672;
assign po0002 = pi0664;
assign po0003 = pi0667;
assign po0004 = pi0676;
assign po0005 = pi0673;
assign po0006 = pi0675;
assign po0007 = pi0666;
assign po0008 = pi0679;
assign po0009 = pi0674;
assign po0010 = pi0663;
assign po0011 = pi0670;
assign po0012 = pi0677;
assign po0013 = pi0682;
assign po0014 = pi0671;
assign po0015 = pi0678;
assign po0016 = pi0718;
assign po0017 = pi0707;
assign po0018 = pi0708;
assign po0019 = pi0713;
assign po0020 = pi0711;
assign po0021 = pi0716;
assign po0022 = pi0733;
assign po0023 = pi0712;
assign po0024 = pi0689;
assign po0025 = pi0717;
assign po0026 = pi0692;
assign po0027 = pi0719;
assign po0028 = pi0722;
assign po0029 = pi0714;
assign po0030 = pi0720;
assign po0031 = pi0685;
assign po0032 = pi0837;
assign po0033 = pi0850;
assign po0034 = pi0872;
assign po0035 = pi0871;
assign po0036 = pi0881;
assign po0037 = pi0866;
assign po0038 = pi0876;
assign po0039 = pi0873;
assign po0040 = pi0874;
assign po0041 = pi0859;
assign po0042 = pi0855;
assign po0043 = pi0852;
assign po0044 = pi0870;
assign po0045 = pi0848;
assign po0046 = pi0865;
assign po0047 = pi0856;
assign po0048 = pi0853;
assign po0049 = pi0847;
assign po0050 = pi0857;
assign po0051 = pi0854;
assign po0052 = pi0858;
assign po0053 = pi0845;
assign po0054 = pi0838;
assign po0055 = pi0842;
assign po0056 = pi0843;
assign po0057 = pi0839;
assign po0058 = pi0844;
assign po0059 = pi0868;
assign po0060 = pi0851;
assign po0061 = pi0867;
assign po0062 = pi0880;
assign po0063 = pi0860;
assign po0064 = pi1030;
assign po0065 = pi1034;
assign po0066 = pi1015;
assign po0067 = pi1020;
assign po0068 = pi1025;
assign po0069 = pi1005;
assign po0070 = pi0996;
assign po0071 = pi1012;
assign po0072 = pi0993;
assign po0073 = pi1016;
assign po0074 = pi1021;
assign po0075 = pi1010;
assign po0076 = pi1027;
assign po0077 = pi1018;
assign po0078 = pi1017;
assign po0079 = pi1024;
assign po0080 = pi1009;
assign po0081 = pi1032;
assign po0082 = pi1003;
assign po0083 = pi0997;
assign po0084 = pi1013;
assign po0085 = pi1011;
assign po0086 = pi1008;
assign po0087 = pi1019;
assign po0088 = pi1031;
assign po0089 = pi1022;
assign po0090 = pi1000;
assign po0091 = pi1023;
assign po0092 = pi1002;
assign po0093 = pi1026;
assign po0094 = pi1006;
assign po0095 = pi0998;
assign po0096 = pi0031;
assign po0097 = pi0080;
assign po0098 = pi0893;
assign po0099 = pi0467;
assign po0100 = pi0078;
assign po0101 = pi0112;
assign po0102 = pi0013;
assign po0103 = pi0025;
assign po0104 = pi0226;
assign po0105 = pi0127;
assign po0106 = pi0822;
assign po0107 = pi0808;
assign po0108 = pi0227;
assign po0109 = pi0477;
assign po0110 = pi0834;
assign po0111 = pi0229;
assign po0112 = pi0012;
assign po0113 = pi0011;
assign po0114 = pi0010;
assign po0115 = pi0009;
assign po0116 = pi0008;
assign po0117 = pi0007;
assign po0118 = pi0006;
assign po0119 = pi0005;
assign po0120 = pi0004;
assign po0121 = pi0003;
assign po0122 = pi0000;
assign po0123 = pi0002;
assign po0124 = pi0001;
assign po0125 = pi0310;
assign po0126 = pi0302;
assign po0127 = pi0475;
assign po0128 = pi0474;
assign po0129 = pi0466;
assign po0130 = pi0473;
assign po0131 = pi0471;
assign po0132 = pi0472;
assign po0133 = pi0470;
assign po0134 = pi0469;
assign po0135 = pi0465;
assign po0136 = pi1028;
assign po0137 = pi1033;
assign po0138 = pi0995;
assign po0139 = pi0994;
assign po0140 = pi0028;
assign po0141 = pi0027;
assign po0142 = pi0026;
assign po0143 = pi0029;
assign po0144 = pi0015;
assign po0145 = pi0014;
assign po0146 = pi0021;
assign po0147 = pi0020;
assign po0148 = pi0019;
assign po0149 = pi0018;
assign po0150 = pi0017;
assign po0151 = pi0016;
assign po0152 = pi1096;
assign po0153 = w592;
assign po0154 = ~w658;
assign po0155 = ~w683;
assign po0156 = ~w748;
assign po0157 = w810;
assign po0158 = w882;
assign po0159 = ~w930;
assign po0160 = ~w975;
assign po0161 = w1021;
assign po0162 = ~w1093;
assign po0163 = w1146;
assign po0164 = w1188;
assign po0165 = w1228;
assign po0166 = one;
assign po0167 = ~w1381;
assign po0168 = pi0228;
assign po0169 = pi0022;
assign po0170 = ~pi1090;
assign po0171 = ~w1538;
assign po0172 = w1556;
assign po0173 = ~w1565;
assign po0174 = ~w1579;
assign po0175 = ~w1586;
assign po0176 = ~w1593;
assign po0177 = ~w1600;
assign po0178 = ~w1607;
assign po0179 = pi1089;
assign po0180 = pi0023;
assign po0181 = ~w1381;
assign po0182 = w1655;
assign po0183 = w1667;
assign po0184 = ~w1672;
assign po0185 = ~w1675;
assign po0186 = ~w1678;
assign po0187 = ~w1681;
assign po0188 = pi0037;
assign po0189 = ~w2551;
assign po0190 = ~w2588;
assign po0191 = ~w2792;
assign po0192 = w2928;
assign po0193 = ~w2997;
assign po0194 = w3007;
assign po0195 = ~w3011;
assign po0196 = ~w3023;
assign po0197 = ~w3075;
assign po0198 = w3079;
assign po0199 = ~w3164;
assign po0200 = ~w3198;
assign po0201 = ~w3219;
assign po0202 = w3233;
assign po0203 = w3234;
assign po0204 = ~w3242;
assign po0205 = ~w3251;
assign po0206 = w3253;
assign po0207 = ~w3262;
assign po0208 = ~w3287;
assign po0209 = w3295;
assign po0210 = ~w3315;
assign po0211 = ~w3323;
assign po0212 = ~w3334;
assign po0213 = ~w3339;
assign po0214 = w3348;
assign po0215 = ~w3356;
assign po0216 = w3361;
assign po0217 = ~w3369;
assign po0218 = ~w3377;
assign po0219 = ~w3385;
assign po0220 = w3394;
assign po0221 = ~w3401;
assign po0222 = w3404;
assign po0223 = w3407;
assign po0224 = w3416;
assign po0225 = w3422;
assign po0226 = w3428;
assign po0227 = w3432;
assign po0228 = ~w3448;
assign po0229 = ~w3461;
assign po0230 = ~w3478;
assign po0231 = w3487;
assign po0232 = ~w3504;
assign po0233 = ~w3511;
assign po0234 = w3525;
assign po0235 = w3529;
assign po0236 = w3531;
assign po0237 = w3665;
assign po0238 = w3688;
assign po0239 = w3692;
assign po0240 = w3696;
assign po0241 = ~w3706;
assign po0242 = w3711;
assign po0243 = w3714;
assign po0244 = w3715;
assign po0245 = w3718;
assign po0246 = ~w3726;
assign po0247 = w3731;
assign po0248 = ~w3735;
assign po0249 = w3743;
assign po0250 = w3751;
assign po0251 = ~w3758;
assign po0252 = ~w3764;
assign po0253 = ~w3775;
assign po0254 = w3787;
assign po0255 = ~w3795;
assign po0256 = w3799;
assign po0257 = ~w3817;
assign po0258 = w3830;
assign po0259 = ~w3839;
assign po0260 = w3840;
assign po0261 = w3842;
assign po0262 = ~w3850;
assign po0263 = pi0117;
assign po0264 = ~w3853;
assign po0265 = w3854;
assign po0266 = ~w3866;
assign po0267 = w3868;
assign po0268 = ~w3874;
assign po0269 = ~w3880;
assign po0270 = ~w3881;
assign po0271 = w3887;
assign po0272 = w3896;
assign po0273 = w3900;
assign po0274 = w3903;
assign po0275 = ~w3904;
assign po0276 = w4021;
assign po0277 = w4042;
assign po0278 = w4068;
assign po0279 = w4133;
assign po0280 = ~w4134;
assign po0281 = w4150;
assign po0282 = ~w4254;
assign po0283 = w4311;
assign po0284 = w4323;
assign po0285 = pi0131;
assign po0286 = ~w4333;
assign po0287 = ~w4373;
assign po0288 = ~w4375;
assign po0289 = w4421;
assign po0290 = w4450;
assign po0291 = w4479;
assign po0292 = w4504;
assign po0293 = w4534;
assign po0294 = ~w4544;
assign po0295 = w4574;
assign po0296 = w4590;
assign po0297 = ~w4718;
assign po0298 = ~w4724;
assign po0299 = ~w4730;
assign po0300 = ~w4736;
assign po0301 = ~w4742;
assign po0302 = ~w4748;
assign po0303 = ~w4755;
assign po0304 = ~w4761;
assign po0305 = ~w4767;
assign po0306 = ~w4773;
assign po0307 = ~w4779;
assign po0308 = ~w4785;
assign po0309 = ~w4791;
assign po0310 = ~w4797;
assign po0311 = ~w4803;
assign po0312 = ~w4809;
assign po0313 = ~w4815;
assign po0314 = ~w4821;
assign po0315 = ~w4827;
assign po0316 = ~w4833;
assign po0317 = ~w4839;
assign po0318 = ~w4845;
assign po0319 = ~w4851;
assign po0320 = ~w4857;
assign po0321 = ~w4863;
assign po0322 = ~w4869;
assign po0323 = ~w4875;
assign po0324 = ~w4881;
assign po0325 = ~w4887;
assign po0326 = ~w4893;
assign po0327 = ~w4899;
assign po0328 = ~w4905;
assign po0329 = ~w4911;
assign po0330 = ~w4917;
assign po0331 = ~w4923;
assign po0332 = ~w4929;
assign po0333 = ~w4935;
assign po0334 = ~w4941;
assign po0335 = ~w4947;
assign po0336 = ~w4953;
assign po0337 = ~w4959;
assign po0338 = ~w4965;
assign po0339 = ~w4971;
assign po0340 = ~w4977;
assign po0341 = ~w4983;
assign po0342 = ~w4989;
assign po0343 = ~w4995;
assign po0344 = ~w5001;
assign po0345 = ~w5007;
assign po0346 = ~w5013;
assign po0347 = ~w5019;
assign po0348 = ~w5025;
assign po0349 = ~w5031;
assign po0350 = ~w5037;
assign po0351 = ~w5043;
assign po0352 = w5059;
assign po0353 = w5074;
assign po0354 = ~w5080;
assign po0355 = ~w5091;
assign po0356 = ~w5097;
assign po0357 = ~w5103;
assign po0358 = ~w5146;
assign po0359 = ~w5153;
assign po0360 = ~w5160;
assign po0361 = ~w5178;
assign po0362 = ~w5182;
assign po0363 = ~w5189;
assign po0364 = ~w5195;
assign po0365 = ~w5201;
assign po0366 = ~w5207;
assign po0367 = ~w5213;
assign po0368 = ~w5219;
assign po0369 = ~w5225;
assign po0370 = ~w5231;
assign po0371 = ~w5237;
assign po0372 = ~w5243;
assign po0373 = ~w5249;
assign po0374 = ~w5255;
assign po0375 = ~w5259;
assign po0376 = ~w5265;
assign po0377 = ~w5269;
assign po0378 = ~w5275;
assign po0379 = ~w5281;
assign po0380 = ~w5287;
assign po0381 = ~w5293;
assign po0382 = ~w5304;
assign po0383 = ~w5321;
assign po0384 = w5333;
assign po0385 = ~w5341;
assign po0386 = pi0232;
assign po0387 = w5350;
assign po0388 = pi0236;
assign po0389 = ~w5360;
assign po0390 = w5461;
assign po0391 = ~w5507;
assign po0392 = ~w5556;
assign po0393 = ~w5319;
assign po0394 = ~w5624;
assign po0395 = ~w5669;
assign po0396 = ~w5685;
assign po0397 = ~w5705;
assign po0398 = ~w5718;
assign po0399 = ~w5735;
assign po0400 = ~w5789;
assign po0401 = ~w5797;
assign po0402 = ~w5810;
assign po0403 = ~w5823;
assign po0404 = ~w5829;
assign po0405 = ~w5842;
assign po0406 = ~w5848;
assign po0407 = w5850;
assign po0408 = ~w5860;
assign po0409 = ~w5866;
assign po0410 = ~w5882;
assign po0411 = ~w5894;
assign po0412 = ~w5900;
assign po0413 = ~w5906;
assign po0414 = ~w5912;
assign po0415 = ~w5918;
assign po0416 = ~w5924;
assign po0417 = ~w5930;
assign po0418 = ~w5936;
assign po0419 = ~w5944;
assign po0420 = ~w5959;
assign po0421 = ~w5971;
assign po0422 = ~w5982;
assign po0423 = ~w5993;
assign po0424 = ~w6005;
assign po0425 = ~w6019;
assign po0426 = ~w6030;
assign po0427 = ~w6041;
assign po0428 = ~w6056;
assign po0429 = ~w6067;
assign po0430 = ~w6081;
assign po0431 = ~w6092;
assign po0432 = ~w6104;
assign po0433 = ~w6117;
assign po0434 = ~w6128;
assign po0435 = ~w6139;
assign po0436 = ~w6150;
assign po0437 = ~w6161;
assign po0438 = ~w6172;
assign po0439 = ~w6183;
assign po0440 = ~w6200;
assign po0441 = ~w6205;
assign po0442 = w6254;
assign po0443 = w6271;
assign po0444 = w6273;
assign po0445 = w6286;
assign po0446 = w6288;
assign po0447 = ~w6291;
assign po0448 = ~w6294;
assign po0449 = ~w6297;
assign po0450 = ~w6300;
assign po0451 = ~w6303;
assign po0452 = ~w6306;
assign po0453 = ~w6309;
assign po0454 = ~w6312;
assign po0455 = ~w6315;
assign po0456 = ~w6322;
assign po0457 = ~w6330;
assign po0458 = w6336;
assign po0459 = ~w6352;
assign po0460 = ~w6355;
assign po0461 = ~w6358;
assign po0462 = ~w6361;
assign po0463 = ~w6364;
assign po0464 = ~w6367;
assign po0465 = ~w6370;
assign po0466 = ~w6373;
assign po0467 = ~w6380;
assign po0468 = w6385;
assign po0469 = w6392;
assign po0470 = ~w6399;
assign po0471 = w6404;
assign po0472 = ~w6408;
assign po0473 = ~w6411;
assign po0474 = ~w6415;
assign po0475 = ~w6419;
assign po0476 = ~w6422;
assign po0477 = ~w6425;
assign po0478 = ~w6428;
assign po0479 = ~w6431;
assign po0480 = ~w6434;
assign po0481 = ~w6437;
assign po0482 = ~w6440;
assign po0483 = ~w6443;
assign po0484 = ~w6446;
assign po0485 = ~w6449;
assign po0486 = ~w6452;
assign po0487 = w6456;
assign po0488 = w6460;
assign po0489 = ~w6467;
assign po0490 = ~w6470;
assign po0491 = ~w6473;
assign po0492 = ~w6476;
assign po0493 = ~w6479;
assign po0494 = ~w6482;
assign po0495 = ~w6485;
assign po0496 = ~w6488;
assign po0497 = ~w6493;
assign po0498 = w6497;
assign po0499 = ~w6500;
assign po0500 = ~w6503;
assign po0501 = ~w6506;
assign po0502 = ~w6509;
assign po0503 = ~w6512;
assign po0504 = ~w6515;
assign po0505 = ~w6518;
assign po0506 = ~w6521;
assign po0507 = ~w6524;
assign po0508 = ~w6527;
assign po0509 = ~w6530;
assign po0510 = ~w6533;
assign po0511 = ~w6536;
assign po0512 = ~w6539;
assign po0513 = ~w6542;
assign po0514 = ~w6545;
assign po0515 = ~w6548;
assign po0516 = ~w6551;
assign po0517 = ~w6554;
assign po0518 = ~w6557;
assign po0519 = ~w6560;
assign po0520 = ~w6563;
assign po0521 = ~w6566;
assign po0522 = ~w6569;
assign po0523 = ~w6572;
assign po0524 = ~w6575;
assign po0525 = ~w6578;
assign po0526 = ~w6581;
assign po0527 = ~w6584;
assign po0528 = ~w6587;
assign po0529 = ~w6590;
assign po0530 = ~w6593;
assign po0531 = ~w6596;
assign po0532 = ~w6599;
assign po0533 = ~w6602;
assign po0534 = ~w6605;
assign po0535 = ~w6608;
assign po0536 = ~w6611;
assign po0537 = ~w6614;
assign po0538 = ~w6617;
assign po0539 = ~w6620;
assign po0540 = ~w6623;
assign po0541 = ~w6626;
assign po0542 = ~w6629;
assign po0543 = ~w6632;
assign po0544 = ~w6635;
assign po0545 = ~w6638;
assign po0546 = ~w6641;
assign po0547 = ~w6644;
assign po0548 = ~w6647;
assign po0549 = ~w6650;
assign po0550 = ~w6653;
assign po0551 = ~w6656;
assign po0552 = ~w6659;
assign po0553 = ~w6662;
assign po0554 = ~w6665;
assign po0555 = ~w6668;
assign po0556 = ~w6671;
assign po0557 = ~w6674;
assign po0558 = ~w6677;
assign po0559 = ~w6680;
assign po0560 = ~w6683;
assign po0561 = ~w6686;
assign po0562 = ~w6689;
assign po0563 = ~w6692;
assign po0564 = ~w6695;
assign po0565 = ~w6698;
assign po0566 = ~w6701;
assign po0567 = ~w6704;
assign po0568 = ~w6707;
assign po0569 = ~w6710;
assign po0570 = ~w6713;
assign po0571 = ~w6716;
assign po0572 = ~w6719;
assign po0573 = ~w6722;
assign po0574 = ~w6725;
assign po0575 = ~w6728;
assign po0576 = ~w6731;
assign po0577 = ~w6734;
assign po0578 = ~w6737;
assign po0579 = ~w6740;
assign po0580 = ~w6743;
assign po0581 = ~w6746;
assign po0582 = ~w6749;
assign po0583 = ~w6752;
assign po0584 = ~w6755;
assign po0585 = ~w6758;
assign po0586 = ~w6761;
assign po0587 = ~w6764;
assign po0588 = ~w6767;
assign po0589 = ~w6770;
assign po0590 = ~w6773;
assign po0591 = ~w6776;
assign po0592 = ~w6779;
assign po0593 = ~w6782;
assign po0594 = ~w6785;
assign po0595 = ~w6788;
assign po0596 = ~w6791;
assign po0597 = ~w6794;
assign po0598 = ~w6797;
assign po0599 = ~w6800;
assign po0600 = ~w6803;
assign po0601 = ~w6806;
assign po0602 = ~w6809;
assign po0603 = ~w6812;
assign po0604 = ~w6815;
assign po0605 = ~w6818;
assign po0606 = ~w6821;
assign po0607 = ~w6824;
assign po0608 = ~w6827;
assign po0609 = ~w6830;
assign po0610 = ~w6833;
assign po0611 = ~w6836;
assign po0612 = ~w6839;
assign po0613 = ~w6842;
assign po0614 = w6867;
assign po0615 = ~w6870;
assign po0616 = ~w6873;
assign po0617 = ~w6876;
assign po0618 = ~w6879;
assign po0619 = ~w6882;
assign po0620 = ~w6885;
assign po0621 = ~w6888;
assign po0622 = ~w6893;
assign po0623 = ~w6898;
assign po0624 = ~w6905;
assign po0625 = ~w6908;
assign po0626 = ~w6913;
assign po0627 = ~w6918;
assign po0628 = ~w6923;
assign po0629 = ~w6928;
assign po0630 = ~w6933;
assign po0631 = ~w6938;
assign po0632 = ~w6943;
assign po0633 = ~w6945;
assign po0634 = ~w6948;
assign po0635 = w6949;
assign po0636 = pi0583;
assign po0637 = w6259;
assign po0638 = ~w6952;
assign po0639 = ~w6955;
assign po0640 = ~w6958;
assign po0641 = ~w6961;
assign po0642 = ~w6964;
assign po0643 = ~w6967;
assign po0644 = ~w6970;
assign po0645 = ~w6973;
assign po0646 = ~w6976;
assign po0647 = ~w6979;
assign po0648 = ~w6982;
assign po0649 = ~w6985;
assign po0650 = ~w6988;
assign po0651 = ~w6991;
assign po0652 = ~w6994;
assign po0653 = ~w6997;
assign po0654 = ~w7000;
assign po0655 = ~w7003;
assign po0656 = ~w7006;
assign po0657 = ~w7009;
assign po0658 = ~w7012;
assign po0659 = ~w7015;
assign po0660 = ~w7018;
assign po0661 = ~w7021;
assign po0662 = ~w7024;
assign po0663 = ~w7027;
assign po0664 = ~w7030;
assign po0665 = ~w7033;
assign po0666 = ~w7036;
assign po0667 = ~w7039;
assign po0668 = ~w7042;
assign po0669 = ~w7045;
assign po0670 = ~w7048;
assign po0671 = ~w7051;
assign po0672 = ~w7054;
assign po0673 = ~w7057;
assign po0674 = ~w7060;
assign po0675 = ~w7063;
assign po0676 = ~w7066;
assign po0677 = ~w7069;
assign po0678 = ~w7072;
assign po0679 = ~w7075;
assign po0680 = ~w7078;
assign po0681 = ~w7081;
assign po0682 = ~w7084;
assign po0683 = ~w7087;
assign po0684 = ~w7090;
assign po0685 = ~w7093;
assign po0686 = ~w7096;
assign po0687 = ~w7099;
assign po0688 = ~w7102;
assign po0689 = ~w7105;
assign po0690 = ~w7108;
assign po0691 = ~w7111;
assign po0692 = ~w7114;
assign po0693 = ~w7117;
assign po0694 = ~w7120;
assign po0695 = ~w7123;
assign po0696 = ~w7126;
assign po0697 = ~w7129;
assign po0698 = ~w7132;
assign po0699 = ~w7135;
assign po0700 = ~w7138;
assign po0701 = ~w7141;
assign po0702 = ~w7144;
assign po0703 = ~w7147;
assign po0704 = ~w7150;
assign po0705 = ~w7153;
assign po0706 = ~w7156;
assign po0707 = ~w7159;
assign po0708 = ~w7162;
assign po0709 = ~w7165;
assign po0710 = ~w7168;
assign po0711 = ~w7171;
assign po0712 = ~w7174;
assign po0713 = ~w7177;
assign po0714 = ~w7180;
assign po0715 = ~w7183;
assign po0716 = ~w7186;
assign po0717 = ~w7189;
assign po0718 = ~w7192;
assign po0719 = ~w7195;
assign po0720 = ~w7198;
assign po0721 = ~w7201;
assign po0722 = ~w7204;
assign po0723 = ~w7207;
assign po0724 = w7216;
assign po0725 = ~w7219;
assign po0726 = ~w7222;
assign po0727 = ~w7225;
assign po0728 = ~w7228;
assign po0729 = ~w7231;
assign po0730 = ~w7234;
assign po0731 = ~w7237;
assign po0732 = ~w7240;
assign po0733 = ~w7243;
assign po0734 = ~w7246;
assign po0735 = ~w7249;
assign po0736 = ~w7252;
assign po0737 = ~w7255;
assign po0738 = ~w7258;
assign po0739 = ~w7261;
assign po0740 = w2568;
assign po0741 = ~w7264;
assign po0742 = ~w7267;
assign po0743 = ~w7270;
assign po0744 = ~w7273;
assign po0745 = w7280;
assign po0746 = ~w7301;
assign po0747 = ~w7306;
assign po0748 = w7311;
assign po0749 = w7316;
assign po0750 = ~w7745;
assign po0751 = w7753;
assign po0752 = w7761;
assign po0753 = w7770;
assign po0754 = w7777;
assign po0755 = ~w7783;
assign po0756 = w7789;
assign po0757 = w7794;
assign po0758 = w7798;
assign po0759 = ~w7801;
assign po0760 = w7813;
assign po0761 = w7821;
assign po0762 = w7825;
assign po0763 = ~w7831;
assign po0764 = w7835;
assign po0765 = w7839;
assign po0766 = w7843;
assign po0767 = w7847;
assign po0768 = w7851;
assign po0769 = w7855;
assign po0770 = w7859;
assign po0771 = ~w7865;
assign po0772 = ~w7870;
assign po0773 = ~w7876;
assign po0774 = ~w7882;
assign po0775 = w7886;
assign po0776 = w7890;
assign po0777 = w7894;
assign po0778 = w7898;
assign po0779 = w7902;
assign po0780 = w7906;
assign po0781 = w7915;
assign po0782 = w7924;
assign po0783 = w7928;
assign po0784 = w7932;
assign po0785 = w7936;
assign po0786 = w7940;
assign po0787 = w7944;
assign po0788 = w7948;
assign po0789 = w7952;
assign po0790 = w7956;
assign po0791 = w7960;
assign po0792 = w7964;
assign po0793 = w7968;
assign po0794 = w7972;
assign po0795 = w7976;
assign po0796 = w7980;
assign po0797 = w7984;
assign po0798 = w7988;
assign po0799 = w7992;
assign po0800 = w7996;
assign po0801 = w8000;
assign po0802 = w8004;
assign po0803 = w8008;
assign po0804 = w8012;
assign po0805 = w8016;
assign po0806 = w8020;
assign po0807 = w8024;
assign po0808 = w8028;
assign po0809 = w8032;
assign po0810 = w8036;
assign po0811 = w8040;
assign po0812 = w8044;
assign po0813 = w8048;
assign po0814 = w8052;
assign po0815 = w8056;
assign po0816 = ~w8072;
assign po0817 = w8076;
assign po0818 = w8080;
assign po0819 = w8084;
assign po0820 = ~w8128;
assign po0821 = ~w8166;
assign po0822 = w8170;
assign po0823 = ~w8208;
assign po0824 = ~w8246;
assign po0825 = ~w8284;
assign po0826 = w8288;
assign po0827 = ~w8322;
assign po0828 = ~w8354;
assign po0829 = ~w8392;
assign po0830 = ~w8430;
assign po0831 = ~w8468;
assign po0832 = ~w8506;
assign po0833 = ~w8544;
assign po0834 = ~w8576;
assign po0835 = ~w8608;
assign po0836 = ~w8646;
assign po0837 = w8650;
assign po0838 = w8654;
assign po0839 = ~w8686;
assign po0840 = w454;
assign po0841 = w8695;
assign po0842 = ~w8731;
assign po0843 = w8735;
assign po0844 = w8739;
assign po0845 = w8743;
assign po0846 = ~w8779;
assign po0847 = w8783;
assign po0848 = w8787;
assign po0849 = ~w8823;
assign po0850 = w8827;
assign po0851 = w8831;
assign po0852 = w8835;
assign po0853 = w8839;
assign po0854 = w8843;
assign po0855 = w8847;
assign po0856 = w8851;
assign po0857 = w8855;
assign po0858 = w8859;
assign po0859 = w8863;
assign po0860 = w8867;
assign po0861 = w8871;
assign po0862 = w8875;
assign po0863 = w8879;
assign po0864 = ~w8914;
assign po0865 = ~w8949;
assign po0866 = w8953;
assign po0867 = w8957;
assign po0868 = ~w8992;
assign po0869 = ~w9027;
assign po0870 = ~w9062;
assign po0871 = ~w9098;
assign po0872 = w9102;
assign po0873 = ~w9137;
assign po0874 = ~w9173;
assign po0875 = ~w9208;
assign po0876 = ~w9244;
assign po0877 = ~w9280;
assign po0878 = w9322;
assign po0879 = ~w9358;
assign po0880 = w9362;
assign po0881 = w9366;
assign po0882 = w9370;
assign po0883 = w9374;
assign po0884 = w9378;
assign po0885 = w9382;
assign po0886 = w9386;
assign po0887 = w9390;
assign po0888 = w9399;
assign po0889 = w9403;
assign po0890 = ~w9438;
assign po0891 = w9442;
assign po0892 = w9446;
assign po0893 = w9450;
assign po0894 = w9454;
assign po0895 = w9458;
assign po0896 = ~w9467;
assign po0897 = w7808;
assign po0898 = ~w9471;
assign po0899 = ~w9475;
assign po0900 = ~w9479;
assign po0901 = ~w9483;
assign po0902 = ~w9487;
assign po0903 = ~w9491;
assign po0904 = w9498;
assign po0905 = ~w9502;
assign po0906 = ~w9506;
assign po0907 = ~w9510;
assign po0908 = ~w9514;
assign po0909 = ~w9518;
assign po0910 = ~w9522;
assign po0911 = ~w9526;
assign po0912 = ~w9530;
assign po0913 = ~w9534;
assign po0914 = ~w9538;
assign po0915 = ~w9542;
assign po0916 = ~w9546;
assign po0917 = ~w9550;
assign po0918 = ~w9554;
assign po0919 = ~w9558;
assign po0920 = ~w9562;
assign po0921 = ~w9566;
assign po0922 = w9578;
assign po0923 = ~w9582;
assign po0924 = ~w9586;
assign po0925 = ~w9590;
assign po0926 = w9594;
assign po0927 = ~w9598;
assign po0928 = w9602;
assign po0929 = ~w9606;
assign po0930 = w9611;
assign po0931 = ~w9615;
assign po0932 = w9623;
assign po0933 = ~w9627;
assign po0934 = ~w9631;
assign po0935 = ~w9639;
assign po0936 = ~w9640;
assign po0937 = ~w9641;
assign po0938 = ~w9644;
assign po0939 = ~w9648;
assign po0940 = ~w9651;
assign po0941 = ~w9654;
assign po0942 = ~w9657;
assign po0943 = ~w9660;
assign po0944 = ~w9663;
assign po0945 = ~w9666;
assign po0946 = ~w9669;
assign po0947 = ~w9672;
assign po0948 = ~w9675;
assign po0949 = ~w9678;
assign po0950 = ~w1284;
assign po0951 = ~w9685;
assign po0952 = ~w9688;
assign po0953 = ~w9698;
assign po0954 = w7920;
assign po0955 = ~w9701;
assign po0956 = ~w9704;
assign po0957 = ~w9707;
assign po0958 = ~w9710;
assign po0959 = w9714;
assign po0960 = ~w9717;
assign po0961 = ~w9720;
assign po0962 = ~w9723;
assign po0963 = w9577;
assign po0964 = ~w9726;
assign po0965 = ~w9729;
assign po0966 = ~w9732;
assign po0967 = ~w9735;
assign po0968 = ~w9738;
assign po0969 = ~w9741;
assign po0970 = ~w9744;
assign po0971 = ~w9747;
assign po0972 = ~w9750;
assign po0973 = ~w9753;
assign po0974 = ~w9760;
assign po0975 = ~w9763;
assign po0976 = ~w9769;
assign po0977 = ~w9774;
assign po0978 = w9321;
assign po0979 = w9775;
assign po0980 = w8691;
assign po0981 = w9782;
assign po0982 = ~w9824;
assign po0983 = ~w9864;
assign po0984 = ~w9904;
assign po0985 = ~w9944;
assign po0986 = w9947;
assign po0987 = ~w9957;
assign po0988 = w9463;
assign po0989 = w9962;
assign po0990 = ~w9965;
assign po0991 = w9966;
assign po0992 = ~w9976;
assign po0993 = ~w9979;
assign po0994 = ~w9982;
assign po0995 = ~w9985;
assign po0996 = ~w9988;
assign po0997 = w9989;
assign po0998 = ~w9992;
assign po0999 = ~w9995;
assign po1000 = ~w9998;
assign po1001 = ~w10001;
assign po1002 = ~w10004;
assign po1003 = ~w10007;
assign po1004 = ~w10010;
assign po1005 = ~w10013;
assign po1006 = ~w10016;
assign po1007 = ~w10019;
assign po1008 = ~w10022;
assign po1009 = ~w10025;
assign po1010 = ~w10028;
assign po1011 = ~w10031;
assign po1012 = ~w10034;
assign po1013 = ~w10037;
assign po1014 = ~w10040;
assign po1015 = ~w10043;
assign po1016 = ~w10046;
assign po1017 = ~w10049;
assign po1018 = ~w10052;
assign po1019 = ~w10055;
assign po1020 = ~w10058;
assign po1021 = ~w10061;
assign po1022 = ~w10064;
assign po1023 = ~w10067;
assign po1024 = ~w10070;
assign po1025 = ~w10073;
assign po1026 = ~w10076;
assign po1027 = ~w10079;
assign po1028 = ~w10082;
assign po1029 = ~w10085;
assign po1030 = ~w10088;
assign po1031 = ~w10091;
assign po1032 = ~w10094;
assign po1033 = ~w10097;
assign po1034 = ~w10100;
assign po1035 = ~w10103;
assign po1036 = ~w10106;
assign po1037 = ~w10109;
assign po1038 = ~w529;
assign po1039 = ~w10115;
assign po1040 = ~w10119;
assign po1041 = ~w10123;
assign po1042 = ~w10127;
assign po1043 = ~w10131;
assign po1044 = ~w10135;
assign po1045 = ~w10139;
assign po1046 = ~w10143;
assign po1047 = ~w10147;
assign po1048 = ~w10151;
assign po1049 = ~w5355;
assign po1050 = ~w10155;
assign po1051 = ~w10159;
assign po1052 = ~w10163;
assign po1053 = pi0067;
assign po1054 = ~w10167;
assign po1055 = ~w10171;
assign po1056 = ~w10175;
assign po1057 = ~w2959;
assign po1058 = ~w10179;
assign po1059 = ~w10183;
assign po1060 = ~w10187;
assign po1061 = ~w10191;
assign po1062 = ~w10195;
assign po1063 = ~w10203;
assign po1064 = ~w10207;
assign po1065 = ~w10211;
assign po1066 = ~w10215;
assign po1067 = ~w10219;
assign po1068 = ~w10223;
assign po1069 = ~w10227;
assign po1070 = ~w10232;
assign po1071 = ~w10236;
assign po1072 = ~w10240;
assign po1073 = ~w10244;
assign po1074 = ~w10248;
assign po1075 = ~w10252;
assign po1076 = ~w10255;
assign po1077 = ~w10258;
assign po1078 = ~w10261;
assign po1079 = ~w10264;
assign po1080 = w10266;
assign po1081 = ~w10269;
assign po1082 = ~w10272;
assign po1083 = ~w10275;
assign po1084 = ~w10278;
assign po1085 = ~w10281;
assign po1086 = ~w10284;
assign po1087 = ~w10287;
assign po1088 = ~w10290;
assign po1089 = ~w10293;
assign po1090 = ~w10296;
assign po1091 = ~w10299;
assign po1092 = ~w10302;
assign po1093 = ~w10305;
assign po1094 = ~w10308;
assign po1095 = ~w10311;
assign po1096 = ~w10314;
assign po1097 = ~w10317;
assign po1098 = ~w10320;
assign po1099 = ~w10323;
assign po1100 = ~w10326;
assign po1101 = ~w10327;
assign po1102 = w10328;
assign po1103 = ~w10334;
assign po1104 = ~w10337;
assign po1105 = ~w10340;
assign po1106 = w10342;
assign po1107 = w10344;
assign po1108 = pi1134;
assign po1109 = pi0964;
assign po1110 = ~pi0954;
assign po1111 = pi0965;
assign po1112 = ~w10346;
assign po1113 = pi0991;
assign po1114 = pi0985;
assign po1115 = w10347;
assign po1116 = w10348;
assign po1117 = pi1014;
assign po1118 = w10349;
assign po1119 = pi1029;
assign po1120 = pi1004;
assign po1121 = pi1007;
assign po1122 = w10350;
assign po1123 = pi1135;
assign po1124 = w10351;
assign po1125 = w10352;
assign po1126 = w10353;
assign po1127 = w10354;
assign po1128 = w10355;
assign po1129 = w10356;
assign po1130 = ~pi0278;
assign po1131 = w10357;
assign po1132 = w10358;
assign po1133 = ~w10359;
assign po1134 = pi1064;
assign po1135 = w10360;
assign po1136 = pi0299;
assign po1137 = ~w10361;
assign po1138 = pi1075;
assign po1139 = pi1052;
assign po1140 = pi0771;
assign po1141 = pi0765;
assign po1142 = pi0605;
assign po1143 = pi0601;
assign po1144 = pi0278;
assign po1145 = pi0279;
assign po1146 = ~pi0915;
assign po1147 = ~pi0825;
assign po1148 = ~pi0826;
assign po1149 = ~pi0913;
assign po1150 = ~pi0894;
assign po1151 = ~pi0905;
assign po1152 = pi1095;
assign po1153 = ~pi0890;
assign po1154 = pi1094;
assign po1155 = ~pi0906;
assign po1156 = ~pi0896;
assign po1157 = ~pi0909;
assign po1158 = ~pi0911;
assign po1159 = ~pi0908;
assign po1160 = ~pi0891;
assign po1161 = ~pi0902;
assign po1162 = ~pi0903;
assign po1163 = ~pi0883;
assign po1164 = ~pi0888;
assign po1165 = ~pi0919;
assign po1166 = ~pi0886;
assign po1167 = ~pi0912;
assign po1168 = ~pi0895;
assign po1169 = ~pi0916;
assign po1170 = ~pi0889;
assign po1171 = ~pi0900;
assign po1172 = ~pi0885;
assign po1173 = ~pi0904;
assign po1174 = ~pi0899;
assign po1175 = ~pi0918;
assign po1176 = ~pi0898;
assign po1177 = ~pi0917;
assign po1178 = ~pi0827;
assign po1179 = ~pi0887;
assign po1180 = ~pi0884;
assign po1181 = ~pi0910;
assign po1182 = ~pi0828;
assign po1183 = ~pi0892;
assign po1184 = pi1187;
assign po1185 = pi1172;
assign po1186 = pi1170;
assign po1187 = pi1138;
assign po1188 = pi1177;
assign po1189 = pi1178;
assign po1190 = pi0863;
assign po1191 = pi1203;
assign po1192 = pi1185;
assign po1193 = pi1171;
assign po1194 = pi1192;
assign po1195 = pi1137;
assign po1196 = pi1186;
assign po1197 = pi1165;
assign po1198 = pi1164;
assign po1199 = pi1098;
assign po1200 = pi1183;
assign po1201 = pi0230;
assign po1202 = pi1169;
assign po1203 = pi1136;
assign po1204 = pi1181;
assign po1205 = pi0849;
assign po1206 = pi1193;
assign po1207 = pi1182;
assign po1208 = pi1168;
assign po1209 = pi1175;
assign po1210 = pi1191;
assign po1211 = pi1099;
assign po1212 = pi1174;
assign po1213 = pi1179;
assign po1214 = pi1202;
assign po1215 = pi1176;
assign po1216 = pi1173;
assign po1217 = pi1201;
assign po1218 = pi1167;
assign po1219 = pi0840;
assign po1220 = pi1189;
assign po1221 = pi1195;
assign po1222 = pi0864;
assign po1223 = pi1190;
assign po1224 = pi1188;
assign po1225 = pi1180;
assign po1226 = pi1194;
assign po1227 = pi1097;
assign po1228 = pi1166;
assign po1229 = pi1200;
assign po1230 = pi1184;
endmodule

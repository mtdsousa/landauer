module top (
            a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, b_8, b_9, b_10, b_11, b_12, b_13, b_14, b_15, b_16, b_17, b_18, b_19, b_20, b_21, b_22, b_23, b_24, b_25, b_26, b_27, b_28, b_29, b_30, b_31, b_32, b_33, b_34, b_35, b_36, b_37, b_38, b_39, b_40, b_41, b_42, b_43, b_44, b_45, b_46, b_47, b_48, b_49, b_50, b_51, b_52, b_53, b_54, b_55, b_56, b_57, b_58, b_59, b_60, b_61, b_62, b_63, 
            f_0, f_1, f_2, f_3, f_4, f_5, f_6, f_7, f_8, f_9, f_10, f_11, f_12, f_13, f_14, f_15, f_16, f_17, f_18, f_19, f_20, f_21, f_22, f_23, f_24, f_25, f_26, f_27, f_28, f_29, f_30, f_31, f_32, f_33, f_34, f_35, f_36, f_37, f_38, f_39, f_40, f_41, f_42, f_43, f_44, f_45, f_46, f_47, f_48, f_49, f_50, f_51, f_52, f_53, f_54, f_55, f_56, f_57, f_58, f_59, f_60, f_61, f_62, f_63, f_64, f_65, f_66, f_67, f_68, f_69, f_70, f_71, f_72, f_73, f_74, f_75, f_76, f_77, f_78, f_79, f_80, f_81, f_82, f_83, f_84, f_85, f_86, f_87, f_88, f_89, f_90, f_91, f_92, f_93, f_94, f_95, f_96, f_97, f_98, f_99, f_100, f_101, f_102, f_103, f_104, f_105, f_106, f_107, f_108, f_109, f_110, f_111, f_112, f_113, f_114, f_115, f_116, f_117, f_118, f_119, f_120, f_121, f_122, f_123, f_124, f_125, f_126, f_127);
input a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, b_8, b_9, b_10, b_11, b_12, b_13, b_14, b_15, b_16, b_17, b_18, b_19, b_20, b_21, b_22, b_23, b_24, b_25, b_26, b_27, b_28, b_29, b_30, b_31, b_32, b_33, b_34, b_35, b_36, b_37, b_38, b_39, b_40, b_41, b_42, b_43, b_44, b_45, b_46, b_47, b_48, b_49, b_50, b_51, b_52, b_53, b_54, b_55, b_56, b_57, b_58, b_59, b_60, b_61, b_62, b_63;
output f_0, f_1, f_2, f_3, f_4, f_5, f_6, f_7, f_8, f_9, f_10, f_11, f_12, f_13, f_14, f_15, f_16, f_17, f_18, f_19, f_20, f_21, f_22, f_23, f_24, f_25, f_26, f_27, f_28, f_29, f_30, f_31, f_32, f_33, f_34, f_35, f_36, f_37, f_38, f_39, f_40, f_41, f_42, f_43, f_44, f_45, f_46, f_47, f_48, f_49, f_50, f_51, f_52, f_53, f_54, f_55, f_56, f_57, f_58, f_59, f_60, f_61, f_62, f_63, f_64, f_65, f_66, f_67, f_68, f_69, f_70, f_71, f_72, f_73, f_74, f_75, f_76, f_77, f_78, f_79, f_80, f_81, f_82, f_83, f_84, f_85, f_86, f_87, f_88, f_89, f_90, f_91, f_92, f_93, f_94, f_95, f_96, f_97, f_98, f_99, f_100, f_101, f_102, f_103, f_104, f_105, f_106, f_107, f_108, f_109, f_110, f_111, f_112, f_113, f_114, f_115, f_116, f_117, f_118, f_119, f_120, f_121, f_122, f_123, f_124, f_125, f_126, f_127;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935;
assign w0 = a_0 & b_0;
assign w1 = a_2 & ~w0;
assign w2 = ~a_2 & ~w0;
assign w3 = ~w1 & ~w2;
assign w4 = ~a_0 & a_1;
assign w5 = b_0 & w4;
assign w6 = ~a_1 & a_2;
assign w7 = a_1 & ~a_2;
assign w8 = ~w6 & ~w7;
assign w9 = a_0 & w8;
assign w10 = w8 & w27388;
assign w11 = ~w5 & ~w10;
assign w12 = a_0 & ~w8;
assign w13 = b_0 & ~b_1;
assign w14 = ~b_0 & b_1;
assign w15 = ~w13 & ~w14;
assign w16 = w12 & ~w15;
assign w17 = w11 & ~w16;
assign w18 = a_2 & ~w17;
assign w19 = ~w17 & ~w18;
assign w20 = (w1 & w19) | (w1 & w27841) | (w19 & w27841);
assign w21 = ~w19 & w27842;
assign w22 = ~w20 & ~w21;
assign w23 = w8 & w27843;
assign w24 = ~w8 & w27389;
assign w25 = b_1 & w4;
assign w26 = ~w24 & ~w25;
assign w27 = ~w23 & w26;
assign w28 = b_0 & ~b_2;
assign w29 = b_1 & w28;
assign w30 = b_1 & ~b_2;
assign w31 = ~b_1 & b_2;
assign w32 = ~w30 & ~w31;
assign w33 = b_0 & b_1;
assign w34 = w32 & ~w33;
assign w35 = ~w29 & ~w34;
assign w36 = w12 & w35;
assign w37 = w27 & ~w36;
assign w38 = a_2 & ~w37;
assign w39 = w37 & a_2;
assign w40 = ~w37 & ~w38;
assign w41 = ~w39 & ~w40;
assign w42 = w20 & ~w41;
assign w43 = ~w20 & w41;
assign w44 = ~w42 & ~w43;
assign w45 = w8 & w27390;
assign w46 = ~w8 & w27325;
assign w47 = b_2 & w4;
assign w48 = ~w46 & ~w47;
assign w49 = ~w45 & w48;
assign w50 = b_1 & b_2;
assign w51 = ~w29 & ~w50;
assign w52 = ~b_2 & ~b_3;
assign w53 = b_2 & b_3;
assign w54 = ~w52 & ~w53;
assign w55 = ~w51 & w54;
assign w56 = w51 & ~w54;
assign w57 = ~w55 & ~w56;
assign w58 = w12 & w57;
assign w59 = w49 & ~w58;
assign w60 = (a_2 & w58) | (a_2 & w27326) | (w58 & w27326);
assign w61 = ~w58 & w38071;
assign w62 = ~w59 & ~w60;
assign w63 = a_2 & ~a_3;
assign w64 = ~a_2 & a_3;
assign w65 = ~w63 & ~w64;
assign w66 = b_0 & ~w65;
assign w67 = (w66 & w62) | (w66 & w38072) | (w62 & w38072);
assign w68 = ~w62 & w38073;
assign w69 = ~w67 & ~w68;
assign w70 = w42 & w69;
assign w71 = ~w42 & ~w69;
assign w72 = ~w70 & ~w71;
assign w73 = w8 & w27844;
assign w74 = ~w8 & w27845;
assign w75 = b_3 & w4;
assign w76 = ~w74 & ~w75;
assign w77 = ~w73 & w76;
assign w78 = (~w53 & w51) | (~w53 & w25349) | (w51 & w25349);
assign w79 = ~b_3 & ~b_4;
assign w80 = b_3 & b_4;
assign w81 = ~w79 & ~w80;
assign w82 = ~w78 & w81;
assign w83 = w78 & ~w81;
assign w84 = ~w82 & ~w83;
assign w85 = (w77 & ~w84) | (w77 & w27846) | (~w84 & w27846);
assign w86 = (w84 & w27847) | (w84 & w27848) | (w27847 & w27848);
assign w87 = (w27391 & ~w84) | (w27391 & w38074) | (~w84 & w38074);
assign w88 = ~w85 & ~w86;
assign w89 = ~w87 & ~w88;
assign w90 = (a_5 & w65) | (a_5 & w27849) | (w65 & w27849);
assign w91 = ~a_3 & a_4;
assign w92 = a_3 & ~a_4;
assign w93 = ~w91 & ~w92;
assign w94 = w65 & ~w93;
assign w95 = b_0 & w94;
assign w96 = ~a_4 & a_5;
assign w97 = a_4 & ~a_5;
assign w98 = ~w96 & ~w97;
assign w99 = ~w65 & w98;
assign w100 = b_1 & w99;
assign w101 = ~w95 & ~w100;
assign w102 = ~w65 & ~w98;
assign w103 = ~w15 & w102;
assign w104 = w101 & ~w103;
assign w105 = (a_5 & ~w101) | (a_5 & w25746) | (~w101 & w25746);
assign w106 = w101 & w26103;
assign w107 = ~w104 & ~w105;
assign w108 = (w90 & w107) | (w90 & w26104) | (w107 & w26104);
assign w109 = ~w107 & w27392;
assign w110 = ~w108 & ~w109;
assign w111 = ~w89 & w110;
assign w112 = w89 & w110;
assign w113 = ~w89 & ~w111;
assign w114 = ~w112 & ~w113;
assign w115 = (~w67 & ~w69) | (~w67 & w27393) | (~w69 & w27393);
assign w116 = ~w114 & ~w115;
assign w117 = w114 & w115;
assign w118 = ~w116 & ~w117;
assign w119 = w8 & w27850;
assign w120 = ~w8 & w27851;
assign w121 = b_4 & w4;
assign w122 = ~w120 & ~w121;
assign w123 = ~w119 & w122;
assign w124 = ~b_4 & ~b_5;
assign w125 = b_4 & b_5;
assign w126 = ~w124 & ~w125;
assign w127 = (~w78 & w25747) | (~w78 & w25748) | (w25747 & w25748);
assign w128 = (w78 & w25749) | (w78 & w25750) | (w25749 & w25750);
assign w129 = ~w127 & ~w128;
assign w130 = (w123 & ~w129) | (w123 & w27852) | (~w129 & w27852);
assign w131 = (w129 & w38075) | (w129 & w38076) | (w38075 & w38076);
assign w132 = (~w129 & w38077) | (~w129 & w38078) | (w38077 & w38078);
assign w133 = ~w130 & ~w131;
assign w134 = ~w132 & ~w133;
assign w135 = b_2 & w99;
assign w136 = w65 & ~w98;
assign w137 = w136 & w25350;
assign w138 = b_1 & w94;
assign w139 = ~w137 & ~w138;
assign w140 = w139 & w25751;
assign w141 = w139 & w25752;
assign w142 = ~w140 & ~w141;
assign w143 = a_5 & ~w142;
assign w144 = ~a_5 & w142;
assign w145 = ~w143 & ~w144;
assign w146 = w108 & ~w145;
assign w147 = ~w108 & w145;
assign w148 = ~w146 & ~w147;
assign w149 = ~w134 & w148;
assign w150 = w148 & ~w149;
assign w151 = ~w148 & ~w134;
assign w152 = ~w150 & ~w151;
assign w153 = (~w111 & w114) | (~w111 & w27394) | (w114 & w27394);
assign w154 = ~w152 & ~w153;
assign w155 = w152 & w153;
assign w156 = ~w154 & ~w155;
assign w157 = ~w149 & ~w154;
assign w158 = a_5 & ~a_6;
assign w159 = ~a_5 & a_6;
assign w160 = ~w158 & ~w159;
assign w161 = b_0 & ~w160;
assign w162 = ~w145 & w26105;
assign w163 = w146 & ~w162;
assign w164 = w161 & ~w162;
assign w165 = ~w163 & ~w164;
assign w166 = b_3 & w99;
assign w167 = w136 & w27011;
assign w168 = b_2 & w94;
assign w169 = ~w167 & ~w168;
assign w170 = ~w166 & w169;
assign w171 = w57 & w102;
assign w172 = w170 & ~w171;
assign w173 = a_5 & ~w172;
assign w174 = w172 & a_5;
assign w175 = ~w172 & ~w173;
assign w176 = ~w174 & ~w175;
assign w177 = ~w165 & w176;
assign w178 = w165 & ~w176;
assign w179 = ~w177 & ~w178;
assign w180 = w8 & w27853;
assign w181 = ~w8 & w27854;
assign w182 = b_5 & w4;
assign w183 = ~w181 & ~w182;
assign w184 = ~w180 & w183;
assign w185 = ~b_5 & ~b_6;
assign w186 = b_5 & b_6;
assign w187 = ~w185 & ~w186;
assign w188 = (w187 & w127) | (w187 & w26106) | (w127 & w26106);
assign w189 = ~w127 & w26107;
assign w190 = ~w188 & ~w189;
assign w191 = (w184 & ~w190) | (w184 & w27855) | (~w190 & w27855);
assign w192 = (w190 & w38079) | (w190 & w38080) | (w38079 & w38080);
assign w193 = (~w190 & w38081) | (~w190 & w38082) | (w38081 & w38082);
assign w194 = ~w191 & ~w192;
assign w195 = ~w193 & ~w194;
assign w196 = ~w179 & ~w195;
assign w197 = w179 & w195;
assign w198 = ~w196 & ~w197;
assign w199 = ~w157 & w198;
assign w200 = w157 & ~w198;
assign w201 = ~w199 & ~w200;
assign w202 = ~w196 & ~w199;
assign w203 = w8 & w27856;
assign w204 = ~w8 & w27857;
assign w205 = b_6 & w4;
assign w206 = ~w204 & ~w205;
assign w207 = ~w203 & w206;
assign w208 = ~b_6 & ~b_7;
assign w209 = b_6 & b_7;
assign w210 = ~w208 & ~w209;
assign w211 = (w127 & w26755) | (w127 & w26756) | (w26755 & w26756);
assign w212 = (~w127 & w27858) | (~w127 & w27859) | (w27858 & w27859);
assign w213 = ~w211 & ~w212;
assign w214 = (w207 & ~w213) | (w207 & w27860) | (~w213 & w27860);
assign w215 = (w213 & w38083) | (w213 & w38084) | (w38083 & w38084);
assign w216 = (~w213 & w38085) | (~w213 & w38086) | (w38085 & w38086);
assign w217 = ~w214 & ~w215;
assign w218 = ~w216 & ~w217;
assign w219 = b_4 & w99;
assign w220 = w136 & w26521;
assign w221 = b_3 & w94;
assign w222 = ~w220 & ~w221;
assign w223 = ~w219 & w222;
assign w224 = w84 & w102;
assign w225 = w223 & ~w224;
assign w226 = (a_5 & w224) | (a_5 & w26522) | (w224 & w26522);
assign w227 = ~w224 & w27012;
assign w228 = ~w225 & ~w226;
assign w229 = ~w227 & ~w228;
assign w230 = (a_8 & w160) | (a_8 & w27861) | (w160 & w27861);
assign w231 = ~a_6 & a_7;
assign w232 = a_6 & ~a_7;
assign w233 = ~w231 & ~w232;
assign w234 = w160 & ~w233;
assign w235 = b_0 & w234;
assign w236 = ~a_7 & a_8;
assign w237 = a_7 & ~a_8;
assign w238 = ~w236 & ~w237;
assign w239 = ~w160 & w238;
assign w240 = b_1 & w239;
assign w241 = ~w235 & ~w240;
assign w242 = ~w160 & ~w238;
assign w243 = ~w15 & w242;
assign w244 = w241 & ~w243;
assign w245 = (a_8 & ~w241) | (a_8 & w25753) | (~w241 & w25753);
assign w246 = w241 & w26108;
assign w247 = ~w244 & ~w245;
assign w248 = (w230 & w247) | (w230 & w26109) | (w247 & w26109);
assign w249 = ~w247 & w26757;
assign w250 = ~w248 & ~w249;
assign w251 = ~w229 & w250;
assign w252 = w229 & w250;
assign w253 = ~w229 & ~w251;
assign w254 = ~w252 & ~w253;
assign w255 = (~w162 & w165) | (~w162 & w26523) | (w165 & w26523);
assign w256 = ~w254 & ~w255;
assign w257 = w254 & w255;
assign w258 = ~w256 & ~w257;
assign w259 = ~w218 & w258;
assign w260 = w218 & ~w258;
assign w261 = ~w259 & ~w260;
assign w262 = (w261 & w199) | (w261 & w26758) | (w199 & w26758);
assign w263 = w202 & ~w261;
assign w264 = ~w262 & ~w263;
assign w265 = b_2 & w239;
assign w266 = w160 & ~w238;
assign w267 = w266 & w25351;
assign w268 = b_1 & w234;
assign w269 = ~w267 & ~w268;
assign w270 = ~w265 & w269;
assign w271 = w35 & w242;
assign w272 = w270 & ~w271;
assign w273 = (a_8 & ~w270) | (a_8 & w25754) | (~w270 & w25754);
assign w274 = w270 & w26110;
assign w275 = ~w272 & ~w273;
assign w276 = ~w274 & ~w275;
assign w277 = ~w248 & w276;
assign w278 = w248 & ~w276;
assign w279 = ~w277 & ~w278;
assign w280 = b_5 & w99;
assign w281 = w136 & w27013;
assign w282 = b_4 & w94;
assign w283 = ~w281 & ~w282;
assign w284 = ~w280 & w283;
assign w285 = w102 & w129;
assign w286 = w284 & ~w285;
assign w287 = (a_5 & w285) | (a_5 & w27014) | (w285 & w27014);
assign w288 = ~w285 & w38087;
assign w289 = ~w286 & ~w287;
assign w290 = ~w288 & ~w289;
assign w291 = w279 & ~w290;
assign w292 = w279 & ~w291;
assign w293 = ~w279 & ~w290;
assign w294 = ~w292 & ~w293;
assign w295 = ~w251 & ~w256;
assign w296 = w294 & w295;
assign w297 = ~w294 & ~w295;
assign w298 = ~w296 & ~w297;
assign w299 = w8 & w27862;
assign w300 = ~w8 & w27863;
assign w301 = b_7 & w4;
assign w302 = ~w300 & ~w301;
assign w303 = ~w299 & w302;
assign w304 = ~b_7 & ~b_8;
assign w305 = b_7 & b_8;
assign w306 = ~w304 & ~w305;
assign w307 = (w127 & w26879) | (w127 & w26880) | (w26879 & w26880);
assign w308 = (~w127 & w38088) | (~w127 & w38089) | (w38088 & w38089);
assign w309 = (w303 & ~w27866) | (w303 & w38090) | (~w27866 & w38090);
assign w310 = (w27866 & w38091) | (w27866 & w38092) | (w38091 & w38092);
assign w311 = (w27868 & ~w27866) | (w27868 & w38093) | (~w27866 & w38093);
assign w312 = ~w309 & ~w310;
assign w313 = ~w311 & ~w312;
assign w314 = w298 & ~w313;
assign w315 = w298 & ~w314;
assign w316 = ~w298 & ~w313;
assign w317 = ~w315 & ~w316;
assign w318 = (~w199 & w26881) | (~w199 & w26882) | (w26881 & w26882);
assign w319 = ~w317 & ~w318;
assign w320 = w317 & w318;
assign w321 = ~w319 & ~w320;
assign w322 = b_6 & w99;
assign w323 = w136 & w27869;
assign w324 = b_5 & w94;
assign w325 = ~w323 & ~w324;
assign w326 = ~w322 & w325;
assign w327 = (w326 & ~w190) | (w326 & w27870) | (~w190 & w27870);
assign w328 = (w190 & w38094) | (w190 & w38095) | (w38094 & w38095);
assign w329 = (~w190 & w38096) | (~w190 & w38097) | (w38096 & w38097);
assign w330 = ~w327 & ~w328;
assign w331 = ~w329 & ~w330;
assign w332 = a_8 & ~a_9;
assign w333 = ~a_8 & a_9;
assign w334 = ~w332 & ~w333;
assign w335 = b_0 & ~w334;
assign w336 = (w335 & w276) | (w335 & w26111) | (w276 & w26111);
assign w337 = ~w276 & w26112;
assign w338 = ~w336 & ~w337;
assign w339 = b_3 & w239;
assign w340 = w266 & w26524;
assign w341 = b_2 & w234;
assign w342 = ~w340 & ~w341;
assign w343 = ~w339 & w342;
assign w344 = w57 & w242;
assign w345 = w343 & ~w344;
assign w346 = a_8 & ~w345;
assign w347 = w345 & a_8;
assign w348 = ~w345 & ~w346;
assign w349 = ~w347 & ~w348;
assign w350 = ~w338 & ~w349;
assign w351 = w338 & w349;
assign w352 = ~w350 & ~w351;
assign w353 = ~w331 & w352;
assign w354 = w352 & ~w353;
assign w355 = ~w352 & ~w331;
assign w356 = ~w354 & ~w355;
assign w357 = (~w291 & w295) | (~w291 & w26760) | (w295 & w26760);
assign w358 = w356 & w357;
assign w359 = ~w356 & ~w357;
assign w360 = ~w358 & ~w359;
assign w361 = w8 & w27871;
assign w362 = ~w8 & w27872;
assign w363 = b_8 & w4;
assign w364 = ~w362 & ~w363;
assign w365 = ~w361 & w364;
assign w366 = ~b_8 & ~b_9;
assign w367 = b_8 & b_9;
assign w368 = ~w366 & ~w367;
assign w369 = (w368 & w307) | (w368 & w26883) | (w307 & w26883);
assign w370 = ~w307 & w27873;
assign w371 = ~w369 & ~w370;
assign w372 = (w365 & ~w371) | (w365 & w27874) | (~w371 & w27874);
assign w373 = (w371 & w38098) | (w371 & w38099) | (w38098 & w38099);
assign w374 = (~w371 & w38100) | (~w371 & w38101) | (w38100 & w38101);
assign w375 = ~w372 & ~w373;
assign w376 = ~w374 & ~w375;
assign w377 = w360 & ~w376;
assign w378 = w360 & ~w377;
assign w379 = ~w360 & ~w376;
assign w380 = ~w378 & ~w379;
assign w381 = (~w314 & w317) | (~w314 & w27327) | (w317 & w27327);
assign w382 = ~w380 & ~w381;
assign w383 = w380 & w381;
assign w384 = ~w382 & ~w383;
assign w385 = ~w377 & ~w382;
assign w386 = b_7 & w99;
assign w387 = w136 & w27875;
assign w388 = b_6 & w94;
assign w389 = ~w387 & ~w388;
assign w390 = ~w386 & w389;
assign w391 = (w390 & ~w213) | (w390 & w27876) | (~w213 & w27876);
assign w392 = (w213 & w38102) | (w213 & w38103) | (w38102 & w38103);
assign w393 = (~w213 & w38104) | (~w213 & w38105) | (w38104 & w38105);
assign w394 = ~w391 & ~w392;
assign w395 = ~w393 & ~w394;
assign w396 = ~w276 & w27877;
assign w397 = (~w396 & w338) | (~w396 & w27878) | (w338 & w27878);
assign w398 = b_4 & w239;
assign w399 = w266 & w26525;
assign w400 = b_3 & w234;
assign w401 = ~w399 & ~w400;
assign w402 = ~w398 & w401;
assign w403 = w84 & w242;
assign w404 = w402 & ~w403;
assign w405 = (a_8 & w403) | (a_8 & w26526) | (w403 & w26526);
assign w406 = ~w403 & w27015;
assign w407 = ~w404 & ~w405;
assign w408 = ~w406 & ~w407;
assign w409 = (a_11 & w334) | (a_11 & w27879) | (w334 & w27879);
assign w410 = ~a_9 & a_10;
assign w411 = a_9 & ~a_10;
assign w412 = ~w410 & ~w411;
assign w413 = w334 & ~w412;
assign w414 = b_0 & w413;
assign w415 = ~a_10 & a_11;
assign w416 = a_10 & ~a_11;
assign w417 = ~w415 & ~w416;
assign w418 = ~w334 & w417;
assign w419 = b_1 & w418;
assign w420 = ~w414 & ~w419;
assign w421 = ~w334 & ~w417;
assign w422 = ~w15 & w421;
assign w423 = w420 & ~w422;
assign w424 = (a_11 & ~w420) | (a_11 & w25352) | (~w420 & w25352);
assign w425 = w420 & w25755;
assign w426 = ~w423 & ~w424;
assign w427 = (w409 & w426) | (w409 & w25756) | (w426 & w25756);
assign w428 = ~w426 & w26761;
assign w429 = ~w427 & ~w428;
assign w430 = w408 & ~w429;
assign w431 = ~w408 & w429;
assign w432 = ~w430 & ~w431;
assign w433 = ~w397 & w432;
assign w434 = w397 & ~w432;
assign w435 = ~w433 & ~w434;
assign w436 = ~w395 & w435;
assign w437 = w435 & ~w436;
assign w438 = ~w435 & ~w395;
assign w439 = ~w437 & ~w438;
assign w440 = ~w353 & ~w359;
assign w441 = w439 & w440;
assign w442 = ~w439 & ~w440;
assign w443 = ~w441 & ~w442;
assign w444 = w8 & w27880;
assign w445 = ~w8 & w27881;
assign w446 = b_9 & w4;
assign w447 = ~w445 & ~w446;
assign w448 = ~w444 & w447;
assign w449 = ~b_9 & ~b_10;
assign w450 = b_9 & b_10;
assign w451 = ~w449 & ~w450;
assign w452 = (w307 & w27128) | (w307 & w27129) | (w27128 & w27129);
assign w453 = (~w307 & w27882) | (~w307 & w27883) | (w27882 & w27883);
assign w454 = ~w452 & ~w453;
assign w455 = (w448 & ~w454) | (w448 & w27884) | (~w454 & w27884);
assign w456 = (w454 & w38106) | (w454 & w38107) | (w38106 & w38107);
assign w457 = (~w454 & w38108) | (~w454 & w38109) | (w38108 & w38109);
assign w458 = ~w455 & ~w456;
assign w459 = ~w457 & ~w458;
assign w460 = ~w443 & w459;
assign w461 = w443 & ~w459;
assign w462 = ~w460 & ~w461;
assign w463 = ~w385 & w462;
assign w464 = w385 & ~w462;
assign w465 = ~w463 & ~w464;
assign w466 = (~w461 & w385) | (~w461 & w27395) | (w385 & w27395);
assign w467 = (~w436 & w440) | (~w436 & w27885) | (w440 & w27885);
assign w468 = b_8 & w99;
assign w469 = w136 & w27886;
assign w470 = b_7 & w94;
assign w471 = ~w469 & ~w470;
assign w472 = ~w468 & w471;
assign w473 = ~w308 & w27887;
assign w474 = (w472 & ~w27887) | (w472 & w38110) | (~w27887 & w38110);
assign w475 = (w27887 & w38111) | (w27887 & w38112) | (w38111 & w38112);
assign w476 = ~w473 & w27889;
assign w477 = ~w474 & ~w475;
assign w478 = ~w476 & ~w477;
assign w479 = (~w431 & w397) | (~w431 & w26527) | (w397 & w26527);
assign w480 = b_2 & w418;
assign w481 = w334 & ~w417;
assign w482 = w481 & w24984;
assign w483 = b_1 & w413;
assign w484 = ~w482 & ~w483;
assign w485 = ~w480 & w484;
assign w486 = w35 & w421;
assign w487 = w485 & ~w486;
assign w488 = (a_11 & ~w485) | (a_11 & w25353) | (~w485 & w25353);
assign w489 = w485 & w25757;
assign w490 = ~w487 & ~w488;
assign w491 = ~w489 & ~w490;
assign w492 = ~w427 & w491;
assign w493 = w427 & ~w491;
assign w494 = ~w492 & ~w493;
assign w495 = b_5 & w239;
assign w496 = w266 & w26762;
assign w497 = b_4 & w234;
assign w498 = ~w496 & ~w497;
assign w499 = ~w495 & w498;
assign w500 = w129 & w242;
assign w501 = w499 & ~w500;
assign w502 = (a_8 & w500) | (a_8 & w26763) | (w500 & w26763);
assign w503 = ~w500 & w38113;
assign w504 = ~w501 & ~w502;
assign w505 = ~w503 & ~w504;
assign w506 = w494 & ~w505;
assign w507 = w494 & ~w506;
assign w508 = ~w494 & ~w505;
assign w509 = ~w507 & ~w508;
assign w510 = ~w479 & ~w509;
assign w511 = w479 & w509;
assign w512 = ~w510 & ~w511;
assign w513 = ~w478 & w512;
assign w514 = ~w512 & ~w478;
assign w515 = w512 & ~w513;
assign w516 = ~w514 & ~w515;
assign w517 = ~w467 & ~w516;
assign w518 = ~w467 & ~w517;
assign w519 = w467 & ~w516;
assign w520 = w8 & w27890;
assign w521 = ~w8 & w27891;
assign w522 = b_10 & w4;
assign w523 = ~w521 & ~w522;
assign w524 = ~w520 & w523;
assign w525 = ~b_10 & ~b_11;
assign w526 = b_10 & b_11;
assign w527 = ~w525 & ~w526;
assign w528 = (w307 & w27892) | (w307 & w27893) | (w27892 & w27893);
assign w529 = (~w307 & w27894) | (~w307 & w27895) | (w27894 & w27895);
assign w530 = ~w528 & ~w529;
assign w531 = (w524 & ~w530) | (w524 & w27896) | (~w530 & w27896);
assign w532 = (w530 & w38114) | (w530 & w38115) | (w38114 & w38115);
assign w533 = (~w530 & w38116) | (~w530 & w38117) | (w38116 & w38117);
assign w534 = ~w531 & ~w532;
assign w535 = ~w533 & ~w534;
assign w536 = (w535 & w518) | (w535 & w27328) | (w518 & w27328);
assign w537 = ~w518 & w27329;
assign w538 = ~w536 & ~w537;
assign w539 = ~w466 & ~w538;
assign w540 = w466 & w538;
assign w541 = ~w539 & ~w540;
assign w542 = w8 & w27897;
assign w543 = ~w8 & w27898;
assign w544 = b_11 & w4;
assign w545 = ~w543 & ~w544;
assign w546 = ~w542 & w545;
assign w547 = ~b_11 & ~b_12;
assign w548 = b_11 & b_12;
assign w549 = ~w547 & ~w548;
assign w550 = (w307 & w27396) | (w307 & w27397) | (w27396 & w27397);
assign w551 = (~w307 & w27899) | (~w307 & w27900) | (w27899 & w27900);
assign w552 = ~w550 & ~w551;
assign w553 = (w546 & ~w552) | (w546 & w27901) | (~w552 & w27901);
assign w554 = (w552 & w38118) | (w552 & w38119) | (w38118 & w38119);
assign w555 = (~w552 & w38120) | (~w552 & w38121) | (w38120 & w38121);
assign w556 = ~w553 & ~w554;
assign w557 = ~w555 & ~w556;
assign w558 = b_6 & w239;
assign w559 = w266 & w27902;
assign w560 = b_5 & w234;
assign w561 = ~w559 & ~w560;
assign w562 = ~w558 & w561;
assign w563 = (w562 & ~w190) | (w562 & w27903) | (~w190 & w27903);
assign w564 = (w190 & w38122) | (w190 & w38123) | (w38122 & w38123);
assign w565 = (~w190 & w38124) | (~w190 & w38125) | (w38124 & w38125);
assign w566 = ~w563 & ~w564;
assign w567 = ~w565 & ~w566;
assign w568 = a_11 & ~a_12;
assign w569 = ~a_11 & a_12;
assign w570 = ~w568 & ~w569;
assign w571 = b_0 & ~w570;
assign w572 = (w571 & w491) | (w571 & w25758) | (w491 & w25758);
assign w573 = ~w491 & w25759;
assign w574 = ~w572 & ~w573;
assign w575 = b_3 & w418;
assign w576 = w481 & w26113;
assign w577 = b_2 & w413;
assign w578 = ~w576 & ~w577;
assign w579 = ~w575 & w578;
assign w580 = w57 & w421;
assign w581 = w579 & ~w580;
assign w582 = a_11 & ~w581;
assign w583 = w581 & a_11;
assign w584 = ~w581 & ~w582;
assign w585 = ~w583 & ~w584;
assign w586 = ~w574 & ~w585;
assign w587 = w574 & w585;
assign w588 = ~w586 & ~w587;
assign w589 = ~w567 & w588;
assign w590 = w588 & ~w589;
assign w591 = ~w588 & ~w567;
assign w592 = ~w590 & ~w591;
assign w593 = ~w506 & ~w510;
assign w594 = w592 & w593;
assign w595 = ~w592 & ~w593;
assign w596 = ~w594 & ~w595;
assign w597 = b_9 & w99;
assign w598 = w136 & w27904;
assign w599 = b_8 & w94;
assign w600 = ~w598 & ~w599;
assign w601 = ~w597 & w600;
assign w602 = (w601 & ~w371) | (w601 & w27905) | (~w371 & w27905);
assign w603 = (w371 & w38126) | (w371 & w38127) | (w38126 & w38127);
assign w604 = (~w371 & w38128) | (~w371 & w38129) | (w38128 & w38129);
assign w605 = ~w602 & ~w603;
assign w606 = ~w604 & ~w605;
assign w607 = ~w596 & w606;
assign w608 = w596 & ~w606;
assign w609 = ~w607 & ~w608;
assign w610 = (~w513 & w467) | (~w513 & w26884) | (w467 & w26884);
assign w611 = w609 & ~w610;
assign w612 = ~w609 & w610;
assign w613 = ~w611 & ~w612;
assign w614 = ~w557 & w613;
assign w615 = w613 & ~w614;
assign w616 = ~w613 & ~w557;
assign w617 = ~w615 & ~w616;
assign w618 = (~w535 & w518) | (~w535 & w27398) | (w518 & w27398);
assign w619 = (~w618 & w466) | (~w618 & w27201) | (w466 & w27201);
assign w620 = ~w617 & ~w619;
assign w621 = w617 & w619;
assign w622 = ~w620 & ~w621;
assign w623 = ~w614 & ~w620;
assign w624 = (~w608 & w610) | (~w608 & w27018) | (w610 & w27018);
assign w625 = b_7 & w239;
assign w626 = w266 & w27906;
assign w627 = b_6 & w234;
assign w628 = ~w626 & ~w627;
assign w629 = ~w625 & w628;
assign w630 = (w629 & ~w213) | (w629 & w27907) | (~w213 & w27907);
assign w631 = (w213 & w38130) | (w213 & w38131) | (w38130 & w38131);
assign w632 = (~w213 & w38132) | (~w213 & w38133) | (w38132 & w38133);
assign w633 = ~w630 & ~w631;
assign w634 = ~w632 & ~w633;
assign w635 = ~w491 & w27908;
assign w636 = (~w635 & w574) | (~w635 & w27909) | (w574 & w27909);
assign w637 = b_4 & w418;
assign w638 = w481 & w26114;
assign w639 = b_3 & w413;
assign w640 = ~w638 & ~w639;
assign w641 = ~w637 & w640;
assign w642 = w84 & w421;
assign w643 = w641 & ~w642;
assign w644 = (a_11 & w642) | (a_11 & w26115) | (w642 & w26115);
assign w645 = ~w642 & w26528;
assign w646 = ~w643 & ~w644;
assign w647 = ~w645 & ~w646;
assign w648 = (a_14 & w570) | (a_14 & w27910) | (w570 & w27910);
assign w649 = ~a_12 & a_13;
assign w650 = a_12 & ~a_13;
assign w651 = ~w649 & ~w650;
assign w652 = w570 & ~w651;
assign w653 = b_0 & w652;
assign w654 = ~a_13 & a_14;
assign w655 = a_13 & ~a_14;
assign w656 = ~w654 & ~w655;
assign w657 = ~w570 & w656;
assign w658 = b_1 & w657;
assign w659 = ~w653 & ~w658;
assign w660 = ~w570 & ~w656;
assign w661 = ~w15 & w660;
assign w662 = w659 & ~w661;
assign w663 = (a_14 & ~w659) | (a_14 & w25354) | (~w659 & w25354);
assign w664 = w659 & w25508;
assign w665 = ~w662 & ~w663;
assign w666 = (w648 & w665) | (w648 & w25509) | (w665 & w25509);
assign w667 = ~w665 & w26529;
assign w668 = ~w666 & ~w667;
assign w669 = w647 & ~w668;
assign w670 = ~w647 & w668;
assign w671 = ~w669 & ~w670;
assign w672 = ~w636 & w671;
assign w673 = w636 & ~w671;
assign w674 = ~w672 & ~w673;
assign w675 = ~w634 & w674;
assign w676 = w674 & ~w675;
assign w677 = ~w674 & ~w634;
assign w678 = ~w676 & ~w677;
assign w679 = ~w589 & ~w595;
assign w680 = w678 & w679;
assign w681 = ~w678 & ~w679;
assign w682 = ~w680 & ~w681;
assign w683 = b_10 & w99;
assign w684 = w136 & w27911;
assign w685 = b_9 & w94;
assign w686 = ~w684 & ~w685;
assign w687 = ~w683 & w686;
assign w688 = (w687 & ~w454) | (w687 & w27912) | (~w454 & w27912);
assign w689 = (w454 & w38134) | (w454 & w38135) | (w38134 & w38135);
assign w690 = (~w454 & w38136) | (~w454 & w38137) | (w38136 & w38137);
assign w691 = ~w688 & ~w689;
assign w692 = ~w690 & ~w691;
assign w693 = w682 & ~w692;
assign w694 = ~w682 & w692;
assign w695 = ~w624 & w27202;
assign w696 = ~w624 & ~w695;
assign w697 = ~w693 & ~w695;
assign w698 = ~w695 & w27202;
assign w699 = ~w696 & ~w698;
assign w700 = w8 & w27913;
assign w701 = ~w8 & w27914;
assign w702 = b_12 & w4;
assign w703 = ~w701 & ~w702;
assign w704 = ~w700 & w703;
assign w705 = (~w307 & w27453) | (~w307 & w27454) | (w27453 & w27454);
assign w706 = ~b_12 & ~b_13;
assign w707 = b_12 & b_13;
assign w708 = ~w706 & ~w707;
assign w709 = ~w705 & w708;
assign w710 = w705 & ~w708;
assign w711 = ~w709 & ~w710;
assign w712 = (w704 & ~w711) | (w704 & w27915) | (~w711 & w27915);
assign w713 = (w711 & w38138) | (w711 & w38139) | (w38138 & w38139);
assign w714 = (~w711 & w38140) | (~w711 & w38141) | (w38140 & w38141);
assign w715 = ~w712 & ~w713;
assign w716 = ~w714 & ~w715;
assign w717 = ~w699 & w716;
assign w718 = w699 & ~w716;
assign w719 = ~w717 & ~w718;
assign w720 = ~w623 & ~w719;
assign w721 = w623 & w719;
assign w722 = ~w720 & ~w721;
assign w723 = ~w699 & ~w716;
assign w724 = (~w723 & w623) | (~w723 & w27399) | (w623 & w27399);
assign w725 = w8 & w27916;
assign w726 = ~w8 & w27917;
assign w727 = b_13 & w4;
assign w728 = ~w726 & ~w727;
assign w729 = ~w725 & w728;
assign w730 = ~b_13 & ~b_14;
assign w731 = b_13 & b_14;
assign w732 = ~w730 & ~w731;
assign w733 = (~w705 & w27766) | (~w705 & w27767) | (w27766 & w27767);
assign w734 = (w705 & w27918) | (w705 & w27919) | (w27918 & w27919);
assign w735 = ~w733 & ~w734;
assign w736 = (w729 & ~w735) | (w729 & w27920) | (~w735 & w27920);
assign w737 = (w735 & w38142) | (w735 & w38143) | (w38142 & w38143);
assign w738 = (~w735 & w38144) | (~w735 & w38145) | (w38144 & w38145);
assign w739 = ~w736 & ~w737;
assign w740 = ~w738 & ~w739;
assign w741 = b_11 & w99;
assign w742 = w136 & w27921;
assign w743 = b_10 & w94;
assign w744 = ~w742 & ~w743;
assign w745 = ~w741 & w744;
assign w746 = (w745 & ~w530) | (w745 & w27922) | (~w530 & w27922);
assign w747 = (w530 & w38146) | (w530 & w38147) | (w38146 & w38147);
assign w748 = (~w530 & w38148) | (~w530 & w38149) | (w38148 & w38149);
assign w749 = ~w746 & ~w747;
assign w750 = ~w748 & ~w749;
assign w751 = (~w675 & w679) | (~w675 & w27923) | (w679 & w27923);
assign w752 = (~w670 & w636) | (~w670 & w26116) | (w636 & w26116);
assign w753 = b_2 & w657;
assign w754 = w570 & ~w656;
assign w755 = w754 & w24985;
assign w756 = b_1 & w652;
assign w757 = ~w755 & ~w756;
assign w758 = ~w753 & w757;
assign w759 = w35 & w660;
assign w760 = w758 & ~w759;
assign w761 = (a_14 & ~w758) | (a_14 & w25355) | (~w758 & w25355);
assign w762 = w758 & w25510;
assign w763 = ~w760 & ~w761;
assign w764 = ~w762 & ~w763;
assign w765 = ~w666 & w764;
assign w766 = w666 & ~w764;
assign w767 = ~w765 & ~w766;
assign w768 = b_5 & w418;
assign w769 = w481 & w26885;
assign w770 = b_4 & w413;
assign w771 = ~w769 & ~w770;
assign w772 = ~w768 & w771;
assign w773 = w129 & w421;
assign w774 = w772 & ~w773;
assign w775 = (a_11 & w773) | (a_11 & w26886) | (w773 & w26886);
assign w776 = ~w773 & w38150;
assign w777 = ~w774 & ~w775;
assign w778 = ~w776 & ~w777;
assign w779 = w767 & ~w778;
assign w780 = ~w767 & w778;
assign w781 = ~w752 & w26530;
assign w782 = ~w752 & ~w781;
assign w783 = (~w779 & w752) | (~w779 & w26764) | (w752 & w26764);
assign w784 = ~w780 & w783;
assign w785 = ~w782 & ~w784;
assign w786 = b_8 & w239;
assign w787 = w266 & w27924;
assign w788 = b_7 & w234;
assign w789 = ~w787 & ~w788;
assign w790 = ~w786 & w789;
assign w791 = ~w308 & w27925;
assign w792 = (w790 & ~w27925) | (w790 & w38151) | (~w27925 & w38151);
assign w793 = (w27925 & w38152) | (w27925 & w38153) | (w38152 & w38153);
assign w794 = ~w791 & w27927;
assign w795 = ~w792 & ~w793;
assign w796 = ~w794 & ~w795;
assign w797 = w785 & w796;
assign w798 = ~w785 & ~w796;
assign w799 = ~w797 & ~w798;
assign w800 = ~w751 & w799;
assign w801 = w751 & ~w799;
assign w802 = ~w800 & ~w801;
assign w803 = w750 & ~w802;
assign w804 = ~w750 & w802;
assign w805 = ~w803 & ~w804;
assign w806 = ~w697 & w805;
assign w807 = w697 & ~w805;
assign w808 = ~w806 & ~w807;
assign w809 = w740 & w808;
assign w810 = ~w740 & ~w808;
assign w811 = ~w809 & ~w810;
assign w812 = ~w724 & ~w811;
assign w813 = w724 & w811;
assign w814 = ~w812 & ~w813;
assign w815 = ~w740 & w808;
assign w816 = (~w815 & w724) | (~w815 & w27519) | (w724 & w27519);
assign w817 = w8 & w27928;
assign w818 = ~w8 & w27929;
assign w819 = b_14 & w4;
assign w820 = ~w818 & ~w819;
assign w821 = ~w817 & w820;
assign w822 = ~b_14 & ~b_15;
assign w823 = b_14 & b_15;
assign w824 = ~w822 & ~w823;
assign w825 = (~w705 & w27930) | (~w705 & w27931) | (w27930 & w27931);
assign w826 = (w705 & w27932) | (w705 & w27933) | (w27932 & w27933);
assign w827 = ~w825 & ~w826;
assign w828 = (w821 & ~w827) | (w821 & w27934) | (~w827 & w27934);
assign w829 = (w827 & w38154) | (w827 & w38155) | (w38154 & w38155);
assign w830 = (~w827 & w38156) | (~w827 & w38157) | (w38156 & w38157);
assign w831 = ~w828 & ~w829;
assign w832 = ~w830 & ~w831;
assign w833 = (~w804 & w697) | (~w804 & w27935) | (w697 & w27935);
assign w834 = b_12 & w99;
assign w835 = w136 & w27936;
assign w836 = b_11 & w94;
assign w837 = ~w835 & ~w836;
assign w838 = ~w834 & w837;
assign w839 = (w838 & ~w552) | (w838 & w27937) | (~w552 & w27937);
assign w840 = (w552 & w38158) | (w552 & w38159) | (w38158 & w38159);
assign w841 = (~w552 & w38160) | (~w552 & w38161) | (w38160 & w38161);
assign w842 = ~w839 & ~w840;
assign w843 = ~w841 & ~w842;
assign w844 = (~w798 & w751) | (~w798 & w26765) | (w751 & w26765);
assign w845 = b_9 & w239;
assign w846 = w266 & w27938;
assign w847 = b_8 & w234;
assign w848 = ~w846 & ~w847;
assign w849 = ~w845 & w848;
assign w850 = (w849 & ~w371) | (w849 & w27939) | (~w371 & w27939);
assign w851 = (w371 & w38162) | (w371 & w38163) | (w38162 & w38163);
assign w852 = (~w371 & w38164) | (~w371 & w38165) | (w38164 & w38165);
assign w853 = ~w850 & ~w851;
assign w854 = ~w852 & ~w853;
assign w855 = b_6 & w418;
assign w856 = w481 & w27940;
assign w857 = b_5 & w413;
assign w858 = ~w856 & ~w857;
assign w859 = ~w855 & w858;
assign w860 = (w859 & ~w190) | (w859 & w27941) | (~w190 & w27941);
assign w861 = (w190 & w38166) | (w190 & w38167) | (w38166 & w38167);
assign w862 = (~w190 & w38168) | (~w190 & w38169) | (w38168 & w38169);
assign w863 = ~w860 & ~w861;
assign w864 = ~w862 & ~w863;
assign w865 = a_14 & ~a_15;
assign w866 = ~a_14 & a_15;
assign w867 = ~w865 & ~w866;
assign w868 = b_0 & ~w867;
assign w869 = (w868 & w764) | (w868 & w25511) | (w764 & w25511);
assign w870 = ~w764 & w25512;
assign w871 = ~w869 & ~w870;
assign w872 = b_3 & w657;
assign w873 = w754 & w25760;
assign w874 = b_2 & w652;
assign w875 = ~w873 & ~w874;
assign w876 = ~w872 & w875;
assign w877 = w57 & w660;
assign w878 = w876 & ~w877;
assign w879 = a_14 & ~w878;
assign w880 = w878 & a_14;
assign w881 = ~w878 & ~w879;
assign w882 = ~w880 & ~w881;
assign w883 = ~w871 & ~w882;
assign w884 = w871 & w882;
assign w885 = ~w883 & ~w884;
assign w886 = ~w864 & w885;
assign w887 = w885 & ~w886;
assign w888 = ~w885 & ~w864;
assign w889 = ~w887 & ~w888;
assign w890 = ~w783 & ~w889;
assign w891 = w783 & w889;
assign w892 = ~w890 & ~w891;
assign w893 = ~w854 & w892;
assign w894 = ~w892 & ~w854;
assign w895 = w892 & ~w893;
assign w896 = ~w894 & ~w895;
assign w897 = ~w844 & ~w896;
assign w898 = w844 & w896;
assign w899 = ~w897 & ~w898;
assign w900 = ~w843 & w899;
assign w901 = ~w899 & ~w843;
assign w902 = w899 & ~w900;
assign w903 = ~w901 & ~w902;
assign w904 = ~w833 & ~w903;
assign w905 = w833 & w903;
assign w906 = ~w904 & ~w905;
assign w907 = ~w832 & w906;
assign w908 = ~w906 & ~w832;
assign w909 = w906 & ~w907;
assign w910 = ~w908 & ~w909;
assign w911 = ~w816 & ~w910;
assign w912 = w816 & ~w909;
assign w913 = ~w908 & w912;
assign w914 = ~w911 & ~w913;
assign w915 = (~w907 & w910) | (~w907 & w27520) | (w910 & w27520);
assign w916 = w8 & w27942;
assign w917 = ~w8 & w27943;
assign w918 = b_15 & w4;
assign w919 = ~w917 & ~w918;
assign w920 = ~w916 & w919;
assign w921 = ~b_15 & ~b_16;
assign w922 = b_15 & b_16;
assign w923 = ~w921 & ~w922;
assign w924 = (~w705 & w38170) | (~w705 & w38171) | (w38170 & w38171);
assign w925 = (w705 & w38172) | (w705 & w38173) | (w38172 & w38173);
assign w926 = ~w924 & ~w925;
assign w927 = (w920 & ~w926) | (w920 & w27946) | (~w926 & w27946);
assign w928 = (w926 & w38174) | (w926 & w38175) | (w38174 & w38175);
assign w929 = (~w926 & w38176) | (~w926 & w38177) | (w38176 & w38177);
assign w930 = ~w927 & ~w928;
assign w931 = ~w929 & ~w930;
assign w932 = (~w900 & w903) | (~w900 & w27947) | (w903 & w27947);
assign w933 = b_13 & w99;
assign w934 = w136 & w27948;
assign w935 = b_12 & w94;
assign w936 = ~w934 & ~w935;
assign w937 = ~w933 & w936;
assign w938 = (w937 & ~w711) | (w937 & w27949) | (~w711 & w27949);
assign w939 = (w711 & w38178) | (w711 & w38179) | (w38178 & w38179);
assign w940 = (~w711 & w38180) | (~w711 & w38181) | (w38180 & w38181);
assign w941 = ~w938 & ~w939;
assign w942 = ~w940 & ~w941;
assign w943 = b_10 & w239;
assign w944 = w266 & w27950;
assign w945 = b_9 & w234;
assign w946 = ~w944 & ~w945;
assign w947 = ~w943 & w946;
assign w948 = (w947 & ~w454) | (w947 & w27951) | (~w454 & w27951);
assign w949 = (w454 & w38182) | (w454 & w38183) | (w38182 & w38183);
assign w950 = (~w454 & w38184) | (~w454 & w38185) | (w38184 & w38185);
assign w951 = ~w948 & ~w949;
assign w952 = ~w950 & ~w951;
assign w953 = (~w886 & w889) | (~w886 & w26766) | (w889 & w26766);
assign w954 = b_7 & w418;
assign w955 = w481 & w27952;
assign w956 = b_6 & w413;
assign w957 = ~w955 & ~w956;
assign w958 = ~w954 & w957;
assign w959 = (w958 & ~w213) | (w958 & w27953) | (~w213 & w27953);
assign w960 = (w213 & w38186) | (w213 & w38187) | (w38186 & w38187);
assign w961 = (~w213 & w38188) | (~w213 & w38189) | (w38188 & w38189);
assign w962 = ~w959 & ~w960;
assign w963 = ~w961 & ~w962;
assign w964 = ~w764 & w27954;
assign w965 = (~w964 & w871) | (~w964 & w27955) | (w871 & w27955);
assign w966 = b_4 & w657;
assign w967 = w754 & w25761;
assign w968 = b_3 & w652;
assign w969 = ~w967 & ~w968;
assign w970 = ~w966 & w969;
assign w971 = w84 & w660;
assign w972 = w970 & ~w971;
assign w973 = (a_14 & w971) | (a_14 & w25762) | (w971 & w25762);
assign w974 = ~w971 & w26117;
assign w975 = ~w972 & ~w973;
assign w976 = ~w974 & ~w975;
assign w977 = (a_17 & w867) | (a_17 & w27956) | (w867 & w27956);
assign w978 = ~a_15 & a_16;
assign w979 = a_15 & ~a_16;
assign w980 = ~w978 & ~w979;
assign w981 = w867 & ~w980;
assign w982 = b_0 & w981;
assign w983 = ~a_16 & a_17;
assign w984 = a_16 & ~a_17;
assign w985 = ~w983 & ~w984;
assign w986 = ~w867 & w985;
assign w987 = b_1 & w986;
assign w988 = ~w982 & ~w987;
assign w989 = ~w867 & ~w985;
assign w990 = ~w15 & w989;
assign w991 = w988 & ~w990;
assign w992 = (a_17 & ~w988) | (a_17 & w25356) | (~w988 & w25356);
assign w993 = w988 & w25513;
assign w994 = ~w991 & ~w992;
assign w995 = (w977 & w994) | (w977 & w25514) | (w994 & w25514);
assign w996 = ~w994 & w26118;
assign w997 = ~w995 & ~w996;
assign w998 = w976 & ~w997;
assign w999 = ~w976 & w997;
assign w1000 = ~w998 & ~w999;
assign w1001 = ~w965 & w1000;
assign w1002 = w965 & ~w1000;
assign w1003 = ~w1001 & ~w1002;
assign w1004 = w963 & ~w1003;
assign w1005 = ~w963 & w1003;
assign w1006 = ~w1004 & ~w1005;
assign w1007 = ~w953 & w1006;
assign w1008 = w953 & ~w1006;
assign w1009 = ~w1007 & ~w1008;
assign w1010 = w952 & ~w1009;
assign w1011 = ~w952 & w1009;
assign w1012 = ~w1010 & ~w1011;
assign w1013 = (w1012 & w897) | (w1012 & w26887) | (w897 & w26887);
assign w1014 = ~w897 & w27400;
assign w1015 = ~w1013 & ~w1014;
assign w1016 = w942 & ~w1015;
assign w1017 = ~w942 & w1015;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = (w1018 & w904) | (w1018 & w27727) | (w904 & w27727);
assign w1020 = ~w904 & w27728;
assign w1021 = ~w1019 & ~w1020;
assign w1022 = w931 & w1021;
assign w1023 = ~w931 & ~w1021;
assign w1024 = ~w1022 & ~w1023;
assign w1025 = ~w915 & ~w1024;
assign w1026 = w915 & w1024;
assign w1027 = ~w1025 & ~w1026;
assign w1028 = w8 & w27957;
assign w1029 = ~w8 & w27958;
assign w1030 = b_16 & w4;
assign w1031 = ~w1029 & ~w1030;
assign w1032 = ~w1028 & w1031;
assign w1033 = ~b_16 & ~b_17;
assign w1034 = b_16 & b_17;
assign w1035 = ~w1033 & ~w1034;
assign w1036 = (~w705 & w38190) | (~w705 & w38191) | (w38190 & w38191);
assign w1037 = (w705 & w38192) | (w705 & w38193) | (w38192 & w38193);
assign w1038 = ~w1036 & ~w1037;
assign w1039 = (w1032 & ~w1038) | (w1032 & w27964) | (~w1038 & w27964);
assign w1040 = (w1038 & w38194) | (w1038 & w38195) | (w38194 & w38195);
assign w1041 = (~w1038 & w38196) | (~w1038 & w38197) | (w38196 & w38197);
assign w1042 = ~w1039 & ~w1040;
assign w1043 = ~w1041 & ~w1042;
assign w1044 = (~w1017 & w932) | (~w1017 & w27331) | (w932 & w27331);
assign w1045 = b_14 & w99;
assign w1046 = w136 & w27965;
assign w1047 = b_13 & w94;
assign w1048 = ~w1046 & ~w1047;
assign w1049 = ~w1045 & w1048;
assign w1050 = (w1049 & ~w735) | (w1049 & w27966) | (~w735 & w27966);
assign w1051 = (w735 & w38198) | (w735 & w38199) | (w38198 & w38199);
assign w1052 = (~w735 & w38200) | (~w735 & w38201) | (w38200 & w38201);
assign w1053 = ~w1050 & ~w1051;
assign w1054 = ~w1052 & ~w1053;
assign w1055 = ~w1011 & ~w1013;
assign w1056 = b_11 & w239;
assign w1057 = w266 & w27967;
assign w1058 = b_10 & w234;
assign w1059 = ~w1057 & ~w1058;
assign w1060 = ~w1056 & w1059;
assign w1061 = (w1060 & ~w530) | (w1060 & w27968) | (~w530 & w27968);
assign w1062 = (w530 & w38202) | (w530 & w38203) | (w38202 & w38203);
assign w1063 = (~w530 & w38204) | (~w530 & w38205) | (w38204 & w38205);
assign w1064 = ~w1061 & ~w1062;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = (~w1005 & w953) | (~w1005 & w27969) | (w953 & w27969);
assign w1067 = (~w999 & w965) | (~w999 & w25763) | (w965 & w25763);
assign w1068 = b_2 & w986;
assign w1069 = w867 & ~w985;
assign w1070 = w1069 & w24986;
assign w1071 = b_1 & w981;
assign w1072 = ~w1070 & ~w1071;
assign w1073 = ~w1068 & w1072;
assign w1074 = w35 & w989;
assign w1075 = w1073 & ~w1074;
assign w1076 = (a_17 & ~w1073) | (a_17 & w25357) | (~w1073 & w25357);
assign w1077 = w1073 & w25515;
assign w1078 = ~w1075 & ~w1076;
assign w1079 = ~w1077 & ~w1078;
assign w1080 = ~w995 & w1079;
assign w1081 = w995 & ~w1079;
assign w1082 = ~w1080 & ~w1081;
assign w1083 = b_5 & w657;
assign w1084 = w754 & w26767;
assign w1085 = b_4 & w652;
assign w1086 = ~w1084 & ~w1085;
assign w1087 = ~w1083 & w1086;
assign w1088 = w129 & w660;
assign w1089 = w1087 & ~w1088;
assign w1090 = (a_14 & w1088) | (a_14 & w26768) | (w1088 & w26768);
assign w1091 = ~w1088 & w38206;
assign w1092 = ~w1089 & ~w1090;
assign w1093 = ~w1091 & ~w1092;
assign w1094 = w1082 & ~w1093;
assign w1095 = ~w1082 & w1093;
assign w1096 = ~w1067 & w26119;
assign w1097 = ~w1067 & ~w1096;
assign w1098 = (~w1094 & w1067) | (~w1094 & w26531) | (w1067 & w26531);
assign w1099 = ~w1095 & w1098;
assign w1100 = ~w1097 & ~w1099;
assign w1101 = b_8 & w418;
assign w1102 = w481 & w27970;
assign w1103 = b_7 & w413;
assign w1104 = ~w1102 & ~w1103;
assign w1105 = ~w1101 & w1104;
assign w1106 = ~w308 & w27971;
assign w1107 = (w1105 & ~w27971) | (w1105 & w38207) | (~w27971 & w38207);
assign w1108 = (w27971 & w38208) | (w27971 & w38209) | (w38208 & w38209);
assign w1109 = ~w1106 & w27973;
assign w1110 = ~w1107 & ~w1108;
assign w1111 = ~w1109 & ~w1110;
assign w1112 = w1100 & w1111;
assign w1113 = ~w1100 & ~w1111;
assign w1114 = ~w1112 & ~w1113;
assign w1115 = ~w1066 & w1114;
assign w1116 = w1066 & ~w1114;
assign w1117 = ~w1115 & ~w1116;
assign w1118 = w1065 & ~w1117;
assign w1119 = ~w1065 & w1117;
assign w1120 = ~w1118 & ~w1119;
assign w1121 = ~w1055 & w1120;
assign w1122 = w1055 & ~w1120;
assign w1123 = ~w1121 & ~w1122;
assign w1124 = w1054 & ~w1123;
assign w1125 = ~w1054 & w1123;
assign w1126 = ~w1124 & ~w1125;
assign w1127 = ~w1044 & w1126;
assign w1128 = w1044 & ~w1126;
assign w1129 = ~w1127 & ~w1128;
assign w1130 = ~w1043 & w1129;
assign w1131 = w1129 & ~w1130;
assign w1132 = ~w1129 & ~w1043;
assign w1133 = ~w1131 & ~w1132;
assign w1134 = ~w931 & w1021;
assign w1135 = (~w1134 & w915) | (~w1134 & w27729) | (w915 & w27729);
assign w1136 = ~w1133 & ~w1135;
assign w1137 = w1133 & w1135;
assign w1138 = ~w1136 & ~w1137;
assign w1139 = (~w1125 & w1044) | (~w1125 & w27401) | (w1044 & w27401);
assign w1140 = b_15 & w99;
assign w1141 = w136 & w27974;
assign w1142 = b_14 & w94;
assign w1143 = ~w1141 & ~w1142;
assign w1144 = ~w1140 & w1143;
assign w1145 = (w1144 & ~w827) | (w1144 & w27975) | (~w827 & w27975);
assign w1146 = (w827 & w38210) | (w827 & w38211) | (w38210 & w38211);
assign w1147 = (~w827 & w38212) | (~w827 & w38213) | (w38212 & w38213);
assign w1148 = ~w1145 & ~w1146;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = (~w1119 & w1055) | (~w1119 & w27019) | (w1055 & w27019);
assign w1151 = b_12 & w239;
assign w1152 = w266 & w27976;
assign w1153 = b_11 & w234;
assign w1154 = ~w1152 & ~w1153;
assign w1155 = ~w1151 & w1154;
assign w1156 = (w1155 & ~w552) | (w1155 & w27977) | (~w552 & w27977);
assign w1157 = (w552 & w38214) | (w552 & w38215) | (w38214 & w38215);
assign w1158 = (~w552 & w38216) | (~w552 & w38217) | (w38216 & w38217);
assign w1159 = ~w1156 & ~w1157;
assign w1160 = ~w1158 & ~w1159;
assign w1161 = (~w1113 & ~w1114) | (~w1113 & w27978) | (~w1114 & w27978);
assign w1162 = b_6 & w657;
assign w1163 = w754 & w27979;
assign w1164 = b_5 & w652;
assign w1165 = ~w1163 & ~w1164;
assign w1166 = ~w1162 & w1165;
assign w1167 = (w1166 & ~w190) | (w1166 & w27980) | (~w190 & w27980);
assign w1168 = (w190 & w38218) | (w190 & w38219) | (w38218 & w38219);
assign w1169 = (~w190 & w38220) | (~w190 & w38221) | (w38220 & w38221);
assign w1170 = ~w1167 & ~w1168;
assign w1171 = ~w1169 & ~w1170;
assign w1172 = a_17 & ~a_18;
assign w1173 = ~a_17 & a_18;
assign w1174 = ~w1172 & ~w1173;
assign w1175 = b_0 & ~w1174;
assign w1176 = (w1175 & w1079) | (w1175 & w25516) | (w1079 & w25516);
assign w1177 = ~w1079 & w25517;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = b_3 & w986;
assign w1180 = w1069 & w25764;
assign w1181 = b_2 & w981;
assign w1182 = ~w1180 & ~w1181;
assign w1183 = ~w1179 & w1182;
assign w1184 = w57 & w989;
assign w1185 = w1183 & ~w1184;
assign w1186 = a_17 & ~w1185;
assign w1187 = w1185 & a_17;
assign w1188 = ~w1185 & ~w1186;
assign w1189 = ~w1187 & ~w1188;
assign w1190 = ~w1178 & ~w1189;
assign w1191 = w1178 & w1189;
assign w1192 = ~w1190 & ~w1191;
assign w1193 = ~w1171 & w1192;
assign w1194 = w1192 & ~w1193;
assign w1195 = ~w1192 & ~w1171;
assign w1196 = ~w1194 & ~w1195;
assign w1197 = ~w1098 & w1196;
assign w1198 = w1098 & ~w1196;
assign w1199 = ~w1197 & ~w1198;
assign w1200 = b_9 & w418;
assign w1201 = w481 & w27981;
assign w1202 = b_8 & w413;
assign w1203 = ~w1201 & ~w1202;
assign w1204 = ~w1200 & w1203;
assign w1205 = (w1204 & ~w371) | (w1204 & w27982) | (~w371 & w27982);
assign w1206 = (w371 & w38222) | (w371 & w38223) | (w38222 & w38223);
assign w1207 = (~w371 & w38224) | (~w371 & w38225) | (w38224 & w38225);
assign w1208 = ~w1205 & ~w1206;
assign w1209 = ~w1207 & ~w1208;
assign w1210 = ~w1199 & ~w1209;
assign w1211 = w1199 & w1209;
assign w1212 = ~w1210 & ~w1211;
assign w1213 = ~w1161 & w1212;
assign w1214 = w1161 & ~w1212;
assign w1215 = ~w1213 & ~w1214;
assign w1216 = w1160 & ~w1215;
assign w1217 = ~w1160 & w1215;
assign w1218 = ~w1216 & ~w1217;
assign w1219 = ~w1150 & w1218;
assign w1220 = w1150 & ~w1218;
assign w1221 = ~w1219 & ~w1220;
assign w1222 = ~w1149 & w1221;
assign w1223 = w1149 & ~w1221;
assign w1224 = ~w1222 & ~w1223;
assign w1225 = ~w1139 & w1224;
assign w1226 = w1139 & ~w1224;
assign w1227 = ~w1225 & ~w1226;
assign w1228 = w8 & w27983;
assign w1229 = ~w8 & w27984;
assign w1230 = b_17 & w4;
assign w1231 = ~w1229 & ~w1230;
assign w1232 = ~w1228 & w1231;
assign w1233 = ~b_17 & ~b_18;
assign w1234 = b_17 & b_18;
assign w1235 = ~w1233 & ~w1234;
assign w1236 = (~w705 & w38226) | (~w705 & w38227) | (w38226 & w38227);
assign w1237 = (w705 & w38228) | (w705 & w38229) | (w38228 & w38229);
assign w1238 = ~w1236 & ~w1237;
assign w1239 = (w1232 & ~w1238) | (w1232 & w27991) | (~w1238 & w27991);
assign w1240 = (w1238 & w38230) | (w1238 & w38231) | (w38230 & w38231);
assign w1241 = (~w1238 & w38232) | (~w1238 & w38233) | (w38232 & w38233);
assign w1242 = ~w1239 & ~w1240;
assign w1243 = ~w1241 & ~w1242;
assign w1244 = w1227 & ~w1243;
assign w1245 = w1227 & ~w1244;
assign w1246 = ~w1227 & ~w1243;
assign w1247 = ~w1245 & ~w1246;
assign w1248 = (~w1130 & w1133) | (~w1130 & w27730) | (w1133 & w27730);
assign w1249 = ~w1247 & ~w1248;
assign w1250 = w1247 & w1248;
assign w1251 = ~w1249 & ~w1250;
assign w1252 = b_16 & w99;
assign w1253 = w136 & w27992;
assign w1254 = b_15 & w94;
assign w1255 = ~w1253 & ~w1254;
assign w1256 = ~w1252 & w1255;
assign w1257 = (w1256 & ~w926) | (w1256 & w27993) | (~w926 & w27993);
assign w1258 = (w926 & w38234) | (w926 & w38235) | (w38234 & w38235);
assign w1259 = (~w926 & w38236) | (~w926 & w38237) | (w38236 & w38237);
assign w1260 = ~w1257 & ~w1258;
assign w1261 = ~w1259 & ~w1260;
assign w1262 = (~w1193 & w1196) | (~w1193 & w26532) | (w1196 & w26532);
assign w1263 = b_7 & w657;
assign w1264 = w754 & w27994;
assign w1265 = b_6 & w652;
assign w1266 = ~w1264 & ~w1265;
assign w1267 = ~w1263 & w1266;
assign w1268 = (w1267 & ~w213) | (w1267 & w27995) | (~w213 & w27995);
assign w1269 = (w213 & w38238) | (w213 & w38239) | (w38238 & w38239);
assign w1270 = (~w213 & w38240) | (~w213 & w38241) | (w38240 & w38241);
assign w1271 = ~w1268 & ~w1269;
assign w1272 = ~w1270 & ~w1271;
assign w1273 = ~w1079 & w27996;
assign w1274 = (~w1273 & w1178) | (~w1273 & w27997) | (w1178 & w27997);
assign w1275 = b_4 & w986;
assign w1276 = w1069 & w25765;
assign w1277 = b_3 & w981;
assign w1278 = ~w1276 & ~w1277;
assign w1279 = ~w1275 & w1278;
assign w1280 = w84 & w989;
assign w1281 = w1279 & ~w1280;
assign w1282 = (a_17 & w1280) | (a_17 & w25766) | (w1280 & w25766);
assign w1283 = ~w1280 & w26120;
assign w1284 = ~w1281 & ~w1282;
assign w1285 = ~w1283 & ~w1284;
assign w1286 = (a_20 & w1174) | (a_20 & w27998) | (w1174 & w27998);
assign w1287 = ~a_18 & a_19;
assign w1288 = a_18 & ~a_19;
assign w1289 = ~w1287 & ~w1288;
assign w1290 = w1174 & ~w1289;
assign w1291 = b_0 & w1290;
assign w1292 = ~a_19 & a_20;
assign w1293 = a_19 & ~a_20;
assign w1294 = ~w1292 & ~w1293;
assign w1295 = ~w1174 & w1294;
assign w1296 = b_1 & w1295;
assign w1297 = ~w1291 & ~w1296;
assign w1298 = ~w1174 & ~w1294;
assign w1299 = ~w15 & w1298;
assign w1300 = w1297 & ~w1299;
assign w1301 = (a_20 & ~w1297) | (a_20 & w25358) | (~w1297 & w25358);
assign w1302 = w1297 & w25518;
assign w1303 = ~w1300 & ~w1301;
assign w1304 = (w1286 & w1303) | (w1286 & w25519) | (w1303 & w25519);
assign w1305 = ~w1303 & w26121;
assign w1306 = ~w1304 & ~w1305;
assign w1307 = w1285 & w1306;
assign w1308 = ~w1285 & ~w1306;
assign w1309 = ~w1307 & ~w1308;
assign w1310 = ~w1274 & ~w1309;
assign w1311 = w1274 & w1309;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = ~w1272 & w1312;
assign w1314 = w1272 & ~w1312;
assign w1315 = ~w1313 & ~w1314;
assign w1316 = ~w1262 & w1315;
assign w1317 = w1262 & ~w1315;
assign w1318 = ~w1316 & ~w1317;
assign w1319 = b_10 & w418;
assign w1320 = w481 & w27999;
assign w1321 = b_9 & w413;
assign w1322 = ~w1320 & ~w1321;
assign w1323 = ~w1319 & w1322;
assign w1324 = (w1323 & ~w454) | (w1323 & w28000) | (~w454 & w28000);
assign w1325 = (w454 & w38242) | (w454 & w38243) | (w38242 & w38243);
assign w1326 = (~w454 & w38244) | (~w454 & w38245) | (w38244 & w38245);
assign w1327 = ~w1324 & ~w1325;
assign w1328 = ~w1326 & ~w1327;
assign w1329 = w1318 & ~w1328;
assign w1330 = w1318 & ~w1329;
assign w1331 = ~w1318 & ~w1328;
assign w1332 = ~w1330 & ~w1331;
assign w1333 = (~w1210 & w1161) | (~w1210 & w26888) | (w1161 & w26888);
assign w1334 = w1332 & w1333;
assign w1335 = ~w1332 & ~w1333;
assign w1336 = ~w1334 & ~w1335;
assign w1337 = b_13 & w239;
assign w1338 = w266 & w28001;
assign w1339 = b_12 & w234;
assign w1340 = ~w1338 & ~w1339;
assign w1341 = ~w1337 & w1340;
assign w1342 = (w1341 & ~w711) | (w1341 & w28002) | (~w711 & w28002);
assign w1343 = (w711 & w38246) | (w711 & w38247) | (w38246 & w38247);
assign w1344 = (~w711 & w38248) | (~w711 & w38249) | (w38248 & w38249);
assign w1345 = ~w1342 & ~w1343;
assign w1346 = ~w1344 & ~w1345;
assign w1347 = ~w1336 & w1346;
assign w1348 = w1336 & ~w1346;
assign w1349 = ~w1347 & ~w1348;
assign w1350 = (~w1217 & w1150) | (~w1217 & w28003) | (w1150 & w28003);
assign w1351 = w1349 & ~w1350;
assign w1352 = ~w1349 & w1350;
assign w1353 = ~w1351 & ~w1352;
assign w1354 = ~w1261 & w1353;
assign w1355 = w1353 & ~w1354;
assign w1356 = ~w1353 & ~w1261;
assign w1357 = ~w1355 & ~w1356;
assign w1358 = (~w1222 & w1139) | (~w1222 & w27521) | (w1139 & w27521);
assign w1359 = w1357 & w1358;
assign w1360 = ~w1357 & ~w1358;
assign w1361 = ~w1359 & ~w1360;
assign w1362 = w8 & w28004;
assign w1363 = ~w8 & w28005;
assign w1364 = b_18 & w4;
assign w1365 = ~w1363 & ~w1364;
assign w1366 = ~w1362 & w1365;
assign w1367 = ~b_18 & ~b_19;
assign w1368 = b_18 & b_19;
assign w1369 = ~w1367 & ~w1368;
assign w1370 = (~w705 & w38250) | (~w705 & w38251) | (w38250 & w38251);
assign w1371 = (w705 & w38252) | (w705 & w38253) | (w38252 & w38253);
assign w1372 = ~w1370 & ~w1371;
assign w1373 = (w1366 & ~w1372) | (w1366 & w28011) | (~w1372 & w28011);
assign w1374 = (w1372 & w38254) | (w1372 & w38255) | (w38254 & w38255);
assign w1375 = (~w1372 & w38256) | (~w1372 & w38257) | (w38256 & w38257);
assign w1376 = ~w1373 & ~w1374;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = w1361 & ~w1377;
assign w1379 = w1361 & ~w1378;
assign w1380 = ~w1361 & ~w1377;
assign w1381 = ~w1379 & ~w1380;
assign w1382 = ~w1244 & ~w1249;
assign w1383 = ~w1381 & ~w1382;
assign w1384 = w1381 & w1382;
assign w1385 = ~w1383 & ~w1384;
assign w1386 = (~w1354 & w1357) | (~w1354 & w27522) | (w1357 & w27522);
assign w1387 = b_17 & w99;
assign w1388 = w136 & w28012;
assign w1389 = b_16 & w94;
assign w1390 = ~w1388 & ~w1389;
assign w1391 = ~w1387 & w1390;
assign w1392 = (w1391 & ~w1038) | (w1391 & w28013) | (~w1038 & w28013);
assign w1393 = (w1038 & w38258) | (w1038 & w38259) | (w38258 & w38259);
assign w1394 = (~w1038 & w38260) | (~w1038 & w38261) | (w38260 & w38261);
assign w1395 = ~w1392 & ~w1393;
assign w1396 = ~w1394 & ~w1395;
assign w1397 = b_14 & w239;
assign w1398 = w266 & w28014;
assign w1399 = b_13 & w234;
assign w1400 = ~w1398 & ~w1399;
assign w1401 = ~w1397 & w1400;
assign w1402 = (w1401 & ~w735) | (w1401 & w28015) | (~w735 & w28015);
assign w1403 = (w735 & w38262) | (w735 & w38263) | (w38262 & w38263);
assign w1404 = (~w735 & w38264) | (~w735 & w38265) | (w38264 & w38265);
assign w1405 = ~w1402 & ~w1403;
assign w1406 = ~w1404 & ~w1405;
assign w1407 = ~w1329 & ~w1335;
assign w1408 = b_11 & w418;
assign w1409 = w481 & w28016;
assign w1410 = b_10 & w413;
assign w1411 = ~w1409 & ~w1410;
assign w1412 = ~w1408 & w1411;
assign w1413 = (w1412 & ~w530) | (w1412 & w28017) | (~w530 & w28017);
assign w1414 = (w530 & w38266) | (w530 & w38267) | (w38266 & w38267);
assign w1415 = (~w530 & w38268) | (~w530 & w38269) | (w38268 & w38269);
assign w1416 = ~w1413 & ~w1414;
assign w1417 = ~w1415 & ~w1416;
assign w1418 = (~w1313 & w1262) | (~w1313 & w28018) | (w1262 & w28018);
assign w1419 = ~w1285 & w1306;
assign w1420 = (~w1419 & w1274) | (~w1419 & w25767) | (w1274 & w25767);
assign w1421 = b_2 & w1295;
assign w1422 = w1174 & ~w1294;
assign w1423 = w1422 & w24987;
assign w1424 = b_1 & w1290;
assign w1425 = ~w1423 & ~w1424;
assign w1426 = ~w1421 & w1425;
assign w1427 = w35 & w1298;
assign w1428 = w1426 & ~w1427;
assign w1429 = (a_20 & ~w1426) | (a_20 & w25359) | (~w1426 & w25359);
assign w1430 = w1426 & w25520;
assign w1431 = ~w1428 & ~w1429;
assign w1432 = ~w1430 & ~w1431;
assign w1433 = ~w1304 & w1432;
assign w1434 = w1304 & ~w1432;
assign w1435 = ~w1433 & ~w1434;
assign w1436 = b_5 & w986;
assign w1437 = w1069 & w26769;
assign w1438 = b_4 & w981;
assign w1439 = ~w1437 & ~w1438;
assign w1440 = ~w1436 & w1439;
assign w1441 = w129 & w989;
assign w1442 = w1440 & ~w1441;
assign w1443 = (a_17 & w1441) | (a_17 & w26770) | (w1441 & w26770);
assign w1444 = ~w1441 & w38270;
assign w1445 = ~w1442 & ~w1443;
assign w1446 = ~w1444 & ~w1445;
assign w1447 = w1435 & ~w1446;
assign w1448 = ~w1435 & w1446;
assign w1449 = ~w1420 & w26122;
assign w1450 = ~w1420 & ~w1449;
assign w1451 = (~w1447 & w1420) | (~w1447 & w26533) | (w1420 & w26533);
assign w1452 = ~w1448 & w1451;
assign w1453 = ~w1450 & ~w1452;
assign w1454 = b_8 & w657;
assign w1455 = w754 & w28019;
assign w1456 = b_7 & w652;
assign w1457 = ~w1455 & ~w1456;
assign w1458 = ~w1454 & w1457;
assign w1459 = ~w308 & w28020;
assign w1460 = (w1458 & ~w28020) | (w1458 & w38271) | (~w28020 & w38271);
assign w1461 = (w28020 & w38272) | (w28020 & w38273) | (w38272 & w38273);
assign w1462 = ~w1459 & w28022;
assign w1463 = ~w1460 & ~w1461;
assign w1464 = ~w1462 & ~w1463;
assign w1465 = w1453 & w1464;
assign w1466 = ~w1453 & ~w1464;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = ~w1418 & w1467;
assign w1469 = w1418 & ~w1467;
assign w1470 = ~w1468 & ~w1469;
assign w1471 = w1417 & ~w1470;
assign w1472 = ~w1417 & w1470;
assign w1473 = ~w1471 & ~w1472;
assign w1474 = ~w1407 & w1473;
assign w1475 = w1407 & ~w1473;
assign w1476 = ~w1474 & ~w1475;
assign w1477 = ~w1406 & w1476;
assign w1478 = w1476 & ~w1477;
assign w1479 = ~w1476 & ~w1406;
assign w1480 = ~w1478 & ~w1479;
assign w1481 = (~w1348 & w1350) | (~w1348 & w27203) | (w1350 & w27203);
assign w1482 = ~w1480 & ~w1481;
assign w1483 = w1480 & w1481;
assign w1484 = ~w1482 & ~w1483;
assign w1485 = ~w1396 & w1484;
assign w1486 = ~w1484 & ~w1396;
assign w1487 = w1484 & ~w1485;
assign w1488 = ~w1486 & ~w1487;
assign w1489 = ~w1386 & ~w1488;
assign w1490 = w1488 & ~w1386;
assign w1491 = ~w1488 & ~w1489;
assign w1492 = ~w1490 & ~w1491;
assign w1493 = w8 & w28023;
assign w1494 = ~w8 & w28024;
assign w1495 = b_19 & w4;
assign w1496 = ~w1494 & ~w1495;
assign w1497 = ~w1493 & w1496;
assign w1498 = ~b_19 & ~b_20;
assign w1499 = b_19 & b_20;
assign w1500 = ~w1498 & ~w1499;
assign w1501 = (~w705 & w38274) | (~w705 & w38275) | (w38274 & w38275);
assign w1502 = (w705 & w38276) | (w705 & w38277) | (w38276 & w38277);
assign w1503 = ~w1501 & ~w1502;
assign w1504 = (w1497 & ~w1503) | (w1497 & w28027) | (~w1503 & w28027);
assign w1505 = (w1503 & w38278) | (w1503 & w38279) | (w38278 & w38279);
assign w1506 = (~w1503 & w38280) | (~w1503 & w38281) | (w38280 & w38281);
assign w1507 = ~w1504 & ~w1505;
assign w1508 = ~w1506 & ~w1507;
assign w1509 = (~w1508 & w1491) | (~w1508 & w27731) | (w1491 & w27731);
assign w1510 = ~w1492 & ~w1509;
assign w1511 = ~w1491 & w38282;
assign w1512 = ~w1510 & ~w1511;
assign w1513 = (~w1378 & w1382) | (~w1378 & w28028) | (w1382 & w28028);
assign w1514 = ~w1512 & ~w1513;
assign w1515 = w1512 & w1513;
assign w1516 = ~w1514 & ~w1515;
assign w1517 = (~w1477 & w1480) | (~w1477 & w27204) | (w1480 & w27204);
assign w1518 = b_15 & w239;
assign w1519 = w266 & w28029;
assign w1520 = b_14 & w234;
assign w1521 = ~w1519 & ~w1520;
assign w1522 = ~w1518 & w1521;
assign w1523 = (w1522 & ~w827) | (w1522 & w28030) | (~w827 & w28030);
assign w1524 = (w827 & w38283) | (w827 & w38284) | (w38283 & w38284);
assign w1525 = (~w827 & w38285) | (~w827 & w38286) | (w38285 & w38286);
assign w1526 = ~w1523 & ~w1524;
assign w1527 = ~w1525 & ~w1526;
assign w1528 = (~w1472 & w1407) | (~w1472 & w27020) | (w1407 & w27020);
assign w1529 = b_12 & w418;
assign w1530 = w481 & w28031;
assign w1531 = b_11 & w413;
assign w1532 = ~w1530 & ~w1531;
assign w1533 = ~w1529 & w1532;
assign w1534 = (w1533 & ~w552) | (w1533 & w28032) | (~w552 & w28032);
assign w1535 = (w552 & w38287) | (w552 & w38288) | (w38287 & w38288);
assign w1536 = (~w552 & w38289) | (~w552 & w38290) | (w38289 & w38290);
assign w1537 = ~w1534 & ~w1535;
assign w1538 = ~w1536 & ~w1537;
assign w1539 = (~w1466 & ~w1467) | (~w1466 & w28033) | (~w1467 & w28033);
assign w1540 = b_6 & w986;
assign w1541 = w1069 & w28034;
assign w1542 = b_5 & w981;
assign w1543 = ~w1541 & ~w1542;
assign w1544 = ~w1540 & w1543;
assign w1545 = (w1544 & ~w190) | (w1544 & w28035) | (~w190 & w28035);
assign w1546 = (w190 & w38291) | (w190 & w38292) | (w38291 & w38292);
assign w1547 = (~w190 & w38293) | (~w190 & w38294) | (w38293 & w38294);
assign w1548 = ~w1545 & ~w1546;
assign w1549 = ~w1547 & ~w1548;
assign w1550 = a_20 & ~a_21;
assign w1551 = ~a_20 & a_21;
assign w1552 = ~w1550 & ~w1551;
assign w1553 = b_0 & ~w1552;
assign w1554 = (w1553 & w1432) | (w1553 & w25521) | (w1432 & w25521);
assign w1555 = ~w1432 & w25522;
assign w1556 = ~w1554 & ~w1555;
assign w1557 = b_3 & w1295;
assign w1558 = w1422 & w25768;
assign w1559 = b_2 & w1290;
assign w1560 = ~w1558 & ~w1559;
assign w1561 = ~w1557 & w1560;
assign w1562 = w57 & w1298;
assign w1563 = w1561 & ~w1562;
assign w1564 = a_20 & ~w1563;
assign w1565 = w1563 & a_20;
assign w1566 = ~w1563 & ~w1564;
assign w1567 = ~w1565 & ~w1566;
assign w1568 = ~w1556 & ~w1567;
assign w1569 = w1556 & w1567;
assign w1570 = ~w1568 & ~w1569;
assign w1571 = ~w1549 & w1570;
assign w1572 = w1570 & ~w1571;
assign w1573 = ~w1570 & ~w1549;
assign w1574 = ~w1572 & ~w1573;
assign w1575 = ~w1451 & w1574;
assign w1576 = w1451 & ~w1574;
assign w1577 = ~w1575 & ~w1576;
assign w1578 = b_9 & w657;
assign w1579 = w754 & w28036;
assign w1580 = b_8 & w652;
assign w1581 = ~w1579 & ~w1580;
assign w1582 = ~w1578 & w1581;
assign w1583 = (w1582 & ~w371) | (w1582 & w28037) | (~w371 & w28037);
assign w1584 = (w371 & w38295) | (w371 & w38296) | (w38295 & w38296);
assign w1585 = (~w371 & w38297) | (~w371 & w38298) | (w38297 & w38298);
assign w1586 = ~w1583 & ~w1584;
assign w1587 = ~w1585 & ~w1586;
assign w1588 = ~w1577 & ~w1587;
assign w1589 = w1577 & w1587;
assign w1590 = ~w1588 & ~w1589;
assign w1591 = ~w1539 & w1590;
assign w1592 = w1539 & ~w1590;
assign w1593 = ~w1591 & ~w1592;
assign w1594 = w1538 & ~w1593;
assign w1595 = ~w1538 & w1593;
assign w1596 = ~w1594 & ~w1595;
assign w1597 = ~w1528 & w1596;
assign w1598 = w1528 & ~w1596;
assign w1599 = ~w1597 & ~w1598;
assign w1600 = ~w1527 & w1599;
assign w1601 = w1527 & ~w1599;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = ~w1517 & w1602;
assign w1604 = w1517 & ~w1602;
assign w1605 = ~w1603 & ~w1604;
assign w1606 = b_18 & w99;
assign w1607 = w136 & w28038;
assign w1608 = b_17 & w94;
assign w1609 = ~w1607 & ~w1608;
assign w1610 = ~w1606 & w1609;
assign w1611 = (w1610 & ~w1238) | (w1610 & w28039) | (~w1238 & w28039);
assign w1612 = (w1238 & w38299) | (w1238 & w38300) | (w38299 & w38300);
assign w1613 = (~w1238 & w38301) | (~w1238 & w38302) | (w38301 & w38302);
assign w1614 = ~w1611 & ~w1612;
assign w1615 = ~w1613 & ~w1614;
assign w1616 = w1605 & ~w1615;
assign w1617 = w1605 & ~w1616;
assign w1618 = ~w1605 & ~w1615;
assign w1619 = ~w1617 & ~w1618;
assign w1620 = (~w1485 & w1488) | (~w1485 & w27523) | (w1488 & w27523);
assign w1621 = w1619 & w1620;
assign w1622 = ~w1619 & ~w1620;
assign w1623 = ~w1621 & ~w1622;
assign w1624 = w8 & w28040;
assign w1625 = ~w8 & w28041;
assign w1626 = b_20 & w4;
assign w1627 = ~w1625 & ~w1626;
assign w1628 = ~w1624 & w1627;
assign w1629 = ~b_20 & ~b_21;
assign w1630 = b_20 & b_21;
assign w1631 = ~w1629 & ~w1630;
assign w1632 = (~w705 & w38303) | (~w705 & w38304) | (w38303 & w38304);
assign w1633 = (w705 & w38305) | (w705 & w38306) | (w38305 & w38306);
assign w1634 = ~w1632 & ~w1633;
assign w1635 = (w1628 & ~w1634) | (w1628 & w28048) | (~w1634 & w28048);
assign w1636 = (w1634 & w38307) | (w1634 & w38308) | (w38307 & w38308);
assign w1637 = (~w1634 & w38309) | (~w1634 & w38310) | (w38309 & w38310);
assign w1638 = ~w1635 & ~w1636;
assign w1639 = ~w1637 & ~w1638;
assign w1640 = w1623 & ~w1639;
assign w1641 = w1623 & ~w1640;
assign w1642 = ~w1623 & ~w1639;
assign w1643 = ~w1641 & ~w1642;
assign w1644 = (~w1509 & w1512) | (~w1509 & w28049) | (w1512 & w28049);
assign w1645 = ~w1643 & ~w1644;
assign w1646 = w1643 & w1644;
assign w1647 = ~w1645 & ~w1646;
assign w1648 = ~w1640 & ~w1645;
assign w1649 = (~w1600 & w1517) | (~w1600 & w27332) | (w1517 & w27332);
assign w1650 = b_16 & w239;
assign w1651 = w266 & w28050;
assign w1652 = b_15 & w234;
assign w1653 = ~w1651 & ~w1652;
assign w1654 = ~w1650 & w1653;
assign w1655 = (w1654 & ~w926) | (w1654 & w28051) | (~w926 & w28051);
assign w1656 = (w926 & w38311) | (w926 & w38312) | (w38311 & w38312);
assign w1657 = (~w926 & w38313) | (~w926 & w38314) | (w38313 & w38314);
assign w1658 = ~w1655 & ~w1656;
assign w1659 = ~w1657 & ~w1658;
assign w1660 = (~w1595 & w1528) | (~w1595 & w28052) | (w1528 & w28052);
assign w1661 = (~w1571 & w1574) | (~w1571 & w26534) | (w1574 & w26534);
assign w1662 = b_7 & w986;
assign w1663 = w1069 & w28053;
assign w1664 = b_6 & w981;
assign w1665 = ~w1663 & ~w1664;
assign w1666 = ~w1662 & w1665;
assign w1667 = (w1666 & ~w213) | (w1666 & w28054) | (~w213 & w28054);
assign w1668 = (w213 & w38315) | (w213 & w38316) | (w38315 & w38316);
assign w1669 = (~w213 & w38317) | (~w213 & w38318) | (w38317 & w38318);
assign w1670 = ~w1667 & ~w1668;
assign w1671 = ~w1669 & ~w1670;
assign w1672 = ~w1432 & w28055;
assign w1673 = (~w1672 & w1556) | (~w1672 & w28056) | (w1556 & w28056);
assign w1674 = b_4 & w1295;
assign w1675 = w1422 & w25769;
assign w1676 = b_3 & w1290;
assign w1677 = ~w1675 & ~w1676;
assign w1678 = ~w1674 & w1677;
assign w1679 = w84 & w1298;
assign w1680 = w1678 & ~w1679;
assign w1681 = (a_20 & w1679) | (a_20 & w25770) | (w1679 & w25770);
assign w1682 = ~w1679 & w26123;
assign w1683 = ~w1680 & ~w1681;
assign w1684 = ~w1682 & ~w1683;
assign w1685 = (a_23 & w1552) | (a_23 & w28057) | (w1552 & w28057);
assign w1686 = ~a_21 & a_22;
assign w1687 = a_21 & ~a_22;
assign w1688 = ~w1686 & ~w1687;
assign w1689 = w1552 & ~w1688;
assign w1690 = b_0 & w1689;
assign w1691 = ~a_22 & a_23;
assign w1692 = a_22 & ~a_23;
assign w1693 = ~w1691 & ~w1692;
assign w1694 = ~w1552 & w1693;
assign w1695 = b_1 & w1694;
assign w1696 = ~w1690 & ~w1695;
assign w1697 = ~w1552 & ~w1693;
assign w1698 = ~w15 & w1697;
assign w1699 = w1696 & ~w1698;
assign w1700 = (a_23 & ~w1696) | (a_23 & w25360) | (~w1696 & w25360);
assign w1701 = w1696 & w25523;
assign w1702 = ~w1699 & ~w1700;
assign w1703 = (w1685 & w1702) | (w1685 & w25524) | (w1702 & w25524);
assign w1704 = ~w1702 & w26124;
assign w1705 = ~w1703 & ~w1704;
assign w1706 = w1684 & w1705;
assign w1707 = ~w1684 & ~w1705;
assign w1708 = ~w1706 & ~w1707;
assign w1709 = ~w1673 & ~w1708;
assign w1710 = w1673 & w1708;
assign w1711 = ~w1709 & ~w1710;
assign w1712 = ~w1671 & w1711;
assign w1713 = w1671 & ~w1711;
assign w1714 = ~w1712 & ~w1713;
assign w1715 = ~w1661 & w1714;
assign w1716 = w1661 & ~w1714;
assign w1717 = ~w1715 & ~w1716;
assign w1718 = b_10 & w657;
assign w1719 = w754 & w28058;
assign w1720 = b_9 & w652;
assign w1721 = ~w1719 & ~w1720;
assign w1722 = ~w1718 & w1721;
assign w1723 = (w1722 & ~w454) | (w1722 & w28059) | (~w454 & w28059);
assign w1724 = (w454 & w38319) | (w454 & w38320) | (w38319 & w38320);
assign w1725 = (~w454 & w38321) | (~w454 & w38322) | (w38321 & w38322);
assign w1726 = ~w1723 & ~w1724;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = w1717 & ~w1727;
assign w1729 = w1717 & ~w1728;
assign w1730 = ~w1717 & ~w1727;
assign w1731 = ~w1729 & ~w1730;
assign w1732 = (~w1588 & w1539) | (~w1588 & w26771) | (w1539 & w26771);
assign w1733 = w1731 & w1732;
assign w1734 = ~w1731 & ~w1732;
assign w1735 = ~w1733 & ~w1734;
assign w1736 = b_13 & w418;
assign w1737 = w481 & w28060;
assign w1738 = b_12 & w413;
assign w1739 = ~w1737 & ~w1738;
assign w1740 = ~w1736 & w1739;
assign w1741 = (w1740 & ~w711) | (w1740 & w28061) | (~w711 & w28061);
assign w1742 = (w711 & w38323) | (w711 & w38324) | (w38323 & w38324);
assign w1743 = (~w711 & w38325) | (~w711 & w38326) | (w38325 & w38326);
assign w1744 = ~w1741 & ~w1742;
assign w1745 = ~w1743 & ~w1744;
assign w1746 = ~w1735 & w1745;
assign w1747 = w1735 & ~w1745;
assign w1748 = ~w1746 & ~w1747;
assign w1749 = ~w1660 & w1748;
assign w1750 = w1660 & ~w1748;
assign w1751 = ~w1749 & ~w1750;
assign w1752 = ~w1659 & w1751;
assign w1753 = w1659 & ~w1751;
assign w1754 = ~w1752 & ~w1753;
assign w1755 = ~w1649 & w1754;
assign w1756 = w1649 & ~w1754;
assign w1757 = ~w1755 & ~w1756;
assign w1758 = b_19 & w99;
assign w1759 = w136 & w28062;
assign w1760 = b_18 & w94;
assign w1761 = ~w1759 & ~w1760;
assign w1762 = ~w1758 & w1761;
assign w1763 = (w1762 & ~w1372) | (w1762 & w28063) | (~w1372 & w28063);
assign w1764 = (w1372 & w38327) | (w1372 & w38328) | (w38327 & w38328);
assign w1765 = (~w1372 & w38329) | (~w1372 & w38330) | (w38329 & w38330);
assign w1766 = ~w1763 & ~w1764;
assign w1767 = ~w1765 & ~w1766;
assign w1768 = w1757 & ~w1767;
assign w1769 = w1757 & ~w1768;
assign w1770 = ~w1757 & ~w1767;
assign w1771 = ~w1769 & ~w1770;
assign w1772 = ~w1616 & ~w1622;
assign w1773 = w1771 & w1772;
assign w1774 = ~w1771 & ~w1772;
assign w1775 = ~w1773 & ~w1774;
assign w1776 = w8 & w28064;
assign w1777 = ~w8 & w28065;
assign w1778 = b_21 & w4;
assign w1779 = ~w1777 & ~w1778;
assign w1780 = ~w1776 & w1779;
assign w1781 = ~b_21 & ~b_22;
assign w1782 = b_21 & b_22;
assign w1783 = ~w1781 & ~w1782;
assign w1784 = (~w705 & w38331) | (~w705 & w38332) | (w38331 & w38332);
assign w1785 = (w705 & w38333) | (w705 & w38334) | (w38333 & w38334);
assign w1786 = ~w1784 & ~w1785;
assign w1787 = (w1780 & ~w1786) | (w1780 & w28072) | (~w1786 & w28072);
assign w1788 = (w1786 & w38335) | (w1786 & w38336) | (w38335 & w38336);
assign w1789 = (~w1786 & w38337) | (~w1786 & w38338) | (w38337 & w38338);
assign w1790 = ~w1787 & ~w1788;
assign w1791 = ~w1789 & ~w1790;
assign w1792 = ~w1775 & w1791;
assign w1793 = w1775 & ~w1791;
assign w1794 = ~w1792 & ~w1793;
assign w1795 = ~w1648 & w1794;
assign w1796 = w1648 & ~w1794;
assign w1797 = ~w1795 & ~w1796;
assign w1798 = (~w1752 & w1649) | (~w1752 & w28073) | (w1649 & w28073);
assign w1799 = b_17 & w239;
assign w1800 = w266 & w28074;
assign w1801 = b_16 & w234;
assign w1802 = ~w1800 & ~w1801;
assign w1803 = ~w1799 & w1802;
assign w1804 = (w1803 & ~w1038) | (w1803 & w28075) | (~w1038 & w28075);
assign w1805 = (w1038 & w38339) | (w1038 & w38340) | (w38339 & w38340);
assign w1806 = (~w1038 & w38341) | (~w1038 & w38342) | (w38341 & w38342);
assign w1807 = ~w1804 & ~w1805;
assign w1808 = ~w1806 & ~w1807;
assign w1809 = b_14 & w418;
assign w1810 = w481 & w28076;
assign w1811 = b_13 & w413;
assign w1812 = ~w1810 & ~w1811;
assign w1813 = ~w1809 & w1812;
assign w1814 = (w1813 & ~w735) | (w1813 & w28077) | (~w735 & w28077);
assign w1815 = (w735 & w38343) | (w735 & w38344) | (w38343 & w38344);
assign w1816 = (~w735 & w38345) | (~w735 & w38346) | (w38345 & w38346);
assign w1817 = ~w1814 & ~w1815;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = ~w1728 & ~w1734;
assign w1820 = b_11 & w657;
assign w1821 = w754 & w28078;
assign w1822 = b_10 & w652;
assign w1823 = ~w1821 & ~w1822;
assign w1824 = ~w1820 & w1823;
assign w1825 = (w1824 & ~w530) | (w1824 & w28079) | (~w530 & w28079);
assign w1826 = (w530 & w38347) | (w530 & w38348) | (w38347 & w38348);
assign w1827 = (~w530 & w38349) | (~w530 & w38350) | (w38349 & w38350);
assign w1828 = ~w1825 & ~w1826;
assign w1829 = ~w1827 & ~w1828;
assign w1830 = (~w1712 & w1661) | (~w1712 & w28080) | (w1661 & w28080);
assign w1831 = ~w1684 & w1705;
assign w1832 = (~w1831 & w1673) | (~w1831 & w25771) | (w1673 & w25771);
assign w1833 = b_2 & w1694;
assign w1834 = w1552 & ~w1693;
assign w1835 = w1834 & w24988;
assign w1836 = b_1 & w1689;
assign w1837 = ~w1835 & ~w1836;
assign w1838 = ~w1833 & w1837;
assign w1839 = w35 & w1697;
assign w1840 = w1838 & ~w1839;
assign w1841 = (a_23 & ~w1838) | (a_23 & w25361) | (~w1838 & w25361);
assign w1842 = w1838 & w25525;
assign w1843 = ~w1840 & ~w1841;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = ~w1703 & w1844;
assign w1846 = w1703 & ~w1844;
assign w1847 = ~w1845 & ~w1846;
assign w1848 = b_5 & w1295;
assign w1849 = w1422 & w26772;
assign w1850 = b_4 & w1290;
assign w1851 = ~w1849 & ~w1850;
assign w1852 = ~w1848 & w1851;
assign w1853 = w129 & w1298;
assign w1854 = w1852 & ~w1853;
assign w1855 = (a_20 & w1853) | (a_20 & w26773) | (w1853 & w26773);
assign w1856 = ~w1853 & w38351;
assign w1857 = ~w1854 & ~w1855;
assign w1858 = ~w1856 & ~w1857;
assign w1859 = w1847 & ~w1858;
assign w1860 = ~w1847 & w1858;
assign w1861 = ~w1832 & w26125;
assign w1862 = ~w1832 & ~w1861;
assign w1863 = (~w1859 & w1832) | (~w1859 & w26535) | (w1832 & w26535);
assign w1864 = ~w1860 & w1863;
assign w1865 = ~w1862 & ~w1864;
assign w1866 = b_8 & w986;
assign w1867 = w1069 & w28081;
assign w1868 = b_7 & w981;
assign w1869 = ~w1867 & ~w1868;
assign w1870 = ~w1866 & w1869;
assign w1871 = ~w308 & w28082;
assign w1872 = (w1870 & ~w28082) | (w1870 & w38352) | (~w28082 & w38352);
assign w1873 = (w28082 & w38353) | (w28082 & w38354) | (w38353 & w38354);
assign w1874 = ~w1871 & w28084;
assign w1875 = ~w1872 & ~w1873;
assign w1876 = ~w1874 & ~w1875;
assign w1877 = w1865 & w1876;
assign w1878 = ~w1865 & ~w1876;
assign w1879 = ~w1877 & ~w1878;
assign w1880 = ~w1830 & w1879;
assign w1881 = w1830 & ~w1879;
assign w1882 = ~w1880 & ~w1881;
assign w1883 = w1829 & ~w1882;
assign w1884 = ~w1829 & w1882;
assign w1885 = ~w1883 & ~w1884;
assign w1886 = ~w1819 & w1885;
assign w1887 = w1819 & ~w1885;
assign w1888 = ~w1886 & ~w1887;
assign w1889 = ~w1818 & w1888;
assign w1890 = w1888 & ~w1889;
assign w1891 = ~w1888 & ~w1818;
assign w1892 = ~w1890 & ~w1891;
assign w1893 = (~w1747 & w1660) | (~w1747 & w27333) | (w1660 & w27333);
assign w1894 = ~w1892 & ~w1893;
assign w1895 = w1892 & w1893;
assign w1896 = ~w1894 & ~w1895;
assign w1897 = ~w1808 & w1896;
assign w1898 = ~w1896 & ~w1808;
assign w1899 = w1896 & ~w1897;
assign w1900 = ~w1898 & ~w1899;
assign w1901 = (~w1798 & w1899) | (~w1798 & w28085) | (w1899 & w28085);
assign w1902 = ~w1899 & w28086;
assign w1903 = ~w1900 & ~w1901;
assign w1904 = ~w1902 & ~w1903;
assign w1905 = b_20 & w99;
assign w1906 = w136 & w28087;
assign w1907 = b_19 & w94;
assign w1908 = ~w1906 & ~w1907;
assign w1909 = ~w1905 & w1908;
assign w1910 = (w1909 & ~w1503) | (w1909 & w28088) | (~w1503 & w28088);
assign w1911 = (w1503 & w38355) | (w1503 & w38356) | (w38355 & w38356);
assign w1912 = (~w1503 & w38357) | (~w1503 & w38358) | (w38357 & w38358);
assign w1913 = ~w1910 & ~w1911;
assign w1914 = ~w1912 & ~w1913;
assign w1915 = (~w1914 & w1903) | (~w1914 & w27524) | (w1903 & w27524);
assign w1916 = ~w1904 & ~w1915;
assign w1917 = ~w1914 & ~w1915;
assign w1918 = ~w1916 & ~w1917;
assign w1919 = (~w1768 & w1772) | (~w1768 & w27732) | (w1772 & w27732);
assign w1920 = w1918 & w1919;
assign w1921 = ~w1918 & ~w1919;
assign w1922 = ~w1920 & ~w1921;
assign w1923 = w8 & w28089;
assign w1924 = ~w8 & w28090;
assign w1925 = b_22 & w4;
assign w1926 = ~w1924 & ~w1925;
assign w1927 = ~w1923 & w1926;
assign w1928 = ~b_22 & ~b_23;
assign w1929 = b_22 & b_23;
assign w1930 = ~w1928 & ~w1929;
assign w1931 = (~w705 & w38359) | (~w705 & w38360) | (w38359 & w38360);
assign w1932 = (w705 & w38361) | (w705 & w38362) | (w38361 & w38362);
assign w1933 = ~w1931 & ~w1932;
assign w1934 = (w1927 & ~w1933) | (w1927 & w28096) | (~w1933 & w28096);
assign w1935 = (w1933 & w38363) | (w1933 & w38364) | (w38363 & w38364);
assign w1936 = (~w1933 & w38365) | (~w1933 & w38366) | (w38365 & w38366);
assign w1937 = ~w1934 & ~w1935;
assign w1938 = ~w1936 & ~w1937;
assign w1939 = w1922 & ~w1938;
assign w1940 = w1922 & ~w1939;
assign w1941 = ~w1922 & ~w1938;
assign w1942 = ~w1940 & ~w1941;
assign w1943 = (~w1793 & w1648) | (~w1793 & w28097) | (w1648 & w28097);
assign w1944 = ~w1942 & ~w1943;
assign w1945 = w1942 & w1943;
assign w1946 = ~w1944 & ~w1945;
assign w1947 = (~w1915 & w1918) | (~w1915 & w27733) | (w1918 & w27733);
assign w1948 = b_21 & w99;
assign w1949 = w136 & w28098;
assign w1950 = b_20 & w94;
assign w1951 = ~w1949 & ~w1950;
assign w1952 = ~w1948 & w1951;
assign w1953 = (w1952 & ~w1634) | (w1952 & w28099) | (~w1634 & w28099);
assign w1954 = (w1634 & w38367) | (w1634 & w38368) | (w38367 & w38368);
assign w1955 = (~w1634 & w38369) | (~w1634 & w38370) | (w38369 & w38370);
assign w1956 = ~w1953 & ~w1954;
assign w1957 = ~w1955 & ~w1956;
assign w1958 = (~w1897 & w1900) | (~w1897 & w27334) | (w1900 & w27334);
assign w1959 = b_15 & w418;
assign w1960 = w481 & w28100;
assign w1961 = b_14 & w413;
assign w1962 = ~w1960 & ~w1961;
assign w1963 = ~w1959 & w1962;
assign w1964 = (w1963 & ~w827) | (w1963 & w28101) | (~w827 & w28101);
assign w1965 = (w827 & w38371) | (w827 & w38372) | (w38371 & w38372);
assign w1966 = (~w827 & w38373) | (~w827 & w38374) | (w38373 & w38374);
assign w1967 = ~w1964 & ~w1965;
assign w1968 = ~w1966 & ~w1967;
assign w1969 = (~w1884 & w1819) | (~w1884 & w27021) | (w1819 & w27021);
assign w1970 = b_12 & w657;
assign w1971 = w754 & w28102;
assign w1972 = b_11 & w652;
assign w1973 = ~w1971 & ~w1972;
assign w1974 = ~w1970 & w1973;
assign w1975 = (w1974 & ~w552) | (w1974 & w28103) | (~w552 & w28103);
assign w1976 = (w552 & w38375) | (w552 & w38376) | (w38375 & w38376);
assign w1977 = (~w552 & w38377) | (~w552 & w38378) | (w38377 & w38378);
assign w1978 = ~w1975 & ~w1976;
assign w1979 = ~w1977 & ~w1978;
assign w1980 = (~w1878 & ~w1879) | (~w1878 & w28104) | (~w1879 & w28104);
assign w1981 = b_6 & w1295;
assign w1982 = w1422 & w28105;
assign w1983 = b_5 & w1290;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = ~w1981 & w1984;
assign w1986 = (w1985 & ~w190) | (w1985 & w28106) | (~w190 & w28106);
assign w1987 = (w190 & w38379) | (w190 & w38380) | (w38379 & w38380);
assign w1988 = (~w190 & w38381) | (~w190 & w38382) | (w38381 & w38382);
assign w1989 = ~w1986 & ~w1987;
assign w1990 = ~w1988 & ~w1989;
assign w1991 = a_23 & ~a_24;
assign w1992 = ~a_23 & a_24;
assign w1993 = ~w1991 & ~w1992;
assign w1994 = b_0 & ~w1993;
assign w1995 = (w1994 & w1844) | (w1994 & w25526) | (w1844 & w25526);
assign w1996 = ~w1844 & w25527;
assign w1997 = ~w1995 & ~w1996;
assign w1998 = b_3 & w1694;
assign w1999 = w1834 & w25772;
assign w2000 = b_2 & w1689;
assign w2001 = ~w1999 & ~w2000;
assign w2002 = ~w1998 & w2001;
assign w2003 = w57 & w1697;
assign w2004 = w2002 & ~w2003;
assign w2005 = a_23 & ~w2004;
assign w2006 = w2004 & a_23;
assign w2007 = ~w2004 & ~w2005;
assign w2008 = ~w2006 & ~w2007;
assign w2009 = ~w1997 & ~w2008;
assign w2010 = w1997 & w2008;
assign w2011 = ~w2009 & ~w2010;
assign w2012 = ~w1990 & w2011;
assign w2013 = w2011 & ~w2012;
assign w2014 = ~w2011 & ~w1990;
assign w2015 = ~w2013 & ~w2014;
assign w2016 = ~w1863 & w2015;
assign w2017 = w1863 & ~w2015;
assign w2018 = ~w2016 & ~w2017;
assign w2019 = b_9 & w986;
assign w2020 = w1069 & w28107;
assign w2021 = b_8 & w981;
assign w2022 = ~w2020 & ~w2021;
assign w2023 = ~w2019 & w2022;
assign w2024 = (w2023 & ~w371) | (w2023 & w28108) | (~w371 & w28108);
assign w2025 = (w371 & w38383) | (w371 & w38384) | (w38383 & w38384);
assign w2026 = (~w371 & w38385) | (~w371 & w38386) | (w38385 & w38386);
assign w2027 = ~w2024 & ~w2025;
assign w2028 = ~w2026 & ~w2027;
assign w2029 = ~w2018 & ~w2028;
assign w2030 = w2018 & w2028;
assign w2031 = ~w2029 & ~w2030;
assign w2032 = ~w1980 & w2031;
assign w2033 = w1980 & ~w2031;
assign w2034 = ~w2032 & ~w2033;
assign w2035 = w1979 & ~w2034;
assign w2036 = ~w1979 & w2034;
assign w2037 = ~w2035 & ~w2036;
assign w2038 = ~w1969 & w2037;
assign w2039 = w1969 & ~w2037;
assign w2040 = ~w2038 & ~w2039;
assign w2041 = ~w1968 & w2040;
assign w2042 = w2040 & ~w2041;
assign w2043 = ~w2040 & ~w1968;
assign w2044 = ~w2042 & ~w2043;
assign w2045 = (~w1889 & w1892) | (~w1889 & w27335) | (w1892 & w27335);
assign w2046 = w2044 & w2045;
assign w2047 = ~w2044 & ~w2045;
assign w2048 = ~w2046 & ~w2047;
assign w2049 = b_18 & w239;
assign w2050 = w266 & w28109;
assign w2051 = b_17 & w234;
assign w2052 = ~w2050 & ~w2051;
assign w2053 = ~w2049 & w2052;
assign w2054 = (w2053 & ~w1238) | (w2053 & w28110) | (~w1238 & w28110);
assign w2055 = (w1238 & w38387) | (w1238 & w38388) | (w38387 & w38388);
assign w2056 = (~w1238 & w38389) | (~w1238 & w38390) | (w38389 & w38390);
assign w2057 = ~w2054 & ~w2055;
assign w2058 = ~w2056 & ~w2057;
assign w2059 = ~w2048 & w2058;
assign w2060 = w2048 & ~w2058;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = ~w1958 & w2061;
assign w2063 = w1958 & ~w2061;
assign w2064 = ~w2062 & ~w2063;
assign w2065 = ~w1957 & w2064;
assign w2066 = ~w2064 & ~w1957;
assign w2067 = w2064 & ~w2065;
assign w2068 = ~w2066 & ~w2067;
assign w2069 = ~w1947 & ~w2068;
assign w2070 = w2068 & ~w1947;
assign w2071 = ~w2068 & ~w2069;
assign w2072 = ~w2070 & ~w2071;
assign w2073 = w8 & w28111;
assign w2074 = ~w8 & w28112;
assign w2075 = b_23 & w4;
assign w2076 = ~w2074 & ~w2075;
assign w2077 = ~w2073 & w2076;
assign w2078 = ~b_23 & ~b_24;
assign w2079 = b_23 & b_24;
assign w2080 = ~w2078 & ~w2079;
assign w2081 = (w2080 & w1931) | (w2080 & w28113) | (w1931 & w28113);
assign w2082 = ~w1931 & w28114;
assign w2083 = ~w2081 & ~w2082;
assign w2084 = (w2077 & ~w2083) | (w2077 & w28115) | (~w2083 & w28115);
assign w2085 = (w2083 & w38391) | (w2083 & w38392) | (w38391 & w38392);
assign w2086 = (~w2083 & w38393) | (~w2083 & w38394) | (w38393 & w38394);
assign w2087 = ~w2084 & ~w2085;
assign w2088 = ~w2086 & ~w2087;
assign w2089 = (~w2088 & w2071) | (~w2088 & w38395) | (w2071 & w38395);
assign w2090 = ~w2072 & ~w2089;
assign w2091 = ~w2071 & w38396;
assign w2092 = ~w2090 & ~w2091;
assign w2093 = ~w1939 & ~w1944;
assign w2094 = ~w2092 & ~w2093;
assign w2095 = w2092 & w2093;
assign w2096 = ~w2094 & ~w2095;
assign w2097 = (~w2089 & w2092) | (~w2089 & w28116) | (w2092 & w28116);
assign w2098 = w8 & w28117;
assign w2099 = ~w8 & w28118;
assign w2100 = b_24 & w4;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = ~w2098 & w2101;
assign w2103 = ~b_24 & ~b_25;
assign w2104 = b_24 & b_25;
assign w2105 = ~w2103 & ~w2104;
assign w2106 = (w1931 & w28121) | (w1931 & w28122) | (w28121 & w28122);
assign w2107 = (~w1931 & w28123) | (~w1931 & w28124) | (w28123 & w28124);
assign w2108 = ~w2106 & ~w2107;
assign w2109 = (w2102 & ~w2108) | (w2102 & w28125) | (~w2108 & w28125);
assign w2110 = (w2108 & w38397) | (w2108 & w38398) | (w38397 & w38398);
assign w2111 = (~w2108 & w38399) | (~w2108 & w38400) | (w38399 & w38400);
assign w2112 = ~w2109 & ~w2110;
assign w2113 = ~w2111 & ~w2112;
assign w2114 = (~w2065 & w2068) | (~w2065 & w38401) | (w2068 & w38401);
assign w2115 = b_16 & w418;
assign w2116 = w481 & w28126;
assign w2117 = b_15 & w413;
assign w2118 = ~w2116 & ~w2117;
assign w2119 = ~w2115 & w2118;
assign w2120 = (w2119 & ~w926) | (w2119 & w28127) | (~w926 & w28127);
assign w2121 = (w926 & w38402) | (w926 & w38403) | (w38402 & w38403);
assign w2122 = (~w926 & w38404) | (~w926 & w38405) | (w38404 & w38405);
assign w2123 = ~w2120 & ~w2121;
assign w2124 = ~w2122 & ~w2123;
assign w2125 = (~w2012 & w2015) | (~w2012 & w26536) | (w2015 & w26536);
assign w2126 = b_7 & w1295;
assign w2127 = w1422 & w28128;
assign w2128 = b_6 & w1290;
assign w2129 = ~w2127 & ~w2128;
assign w2130 = ~w2126 & w2129;
assign w2131 = (w2130 & ~w213) | (w2130 & w28129) | (~w213 & w28129);
assign w2132 = (w213 & w38406) | (w213 & w38407) | (w38406 & w38407);
assign w2133 = (~w213 & w38408) | (~w213 & w38409) | (w38408 & w38409);
assign w2134 = ~w2131 & ~w2132;
assign w2135 = ~w2133 & ~w2134;
assign w2136 = ~w1844 & w28130;
assign w2137 = (~w2136 & w1997) | (~w2136 & w28131) | (w1997 & w28131);
assign w2138 = b_4 & w1694;
assign w2139 = w1834 & w25773;
assign w2140 = b_3 & w1689;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = ~w2138 & w2141;
assign w2143 = w84 & w1697;
assign w2144 = w2142 & ~w2143;
assign w2145 = (a_23 & w2143) | (a_23 & w25774) | (w2143 & w25774);
assign w2146 = ~w2143 & w26126;
assign w2147 = ~w2144 & ~w2145;
assign w2148 = ~w2146 & ~w2147;
assign w2149 = (a_26 & w1993) | (a_26 & w28132) | (w1993 & w28132);
assign w2150 = ~a_24 & a_25;
assign w2151 = a_24 & ~a_25;
assign w2152 = ~w2150 & ~w2151;
assign w2153 = w1993 & ~w2152;
assign w2154 = b_0 & w2153;
assign w2155 = ~a_25 & a_26;
assign w2156 = a_25 & ~a_26;
assign w2157 = ~w2155 & ~w2156;
assign w2158 = ~w1993 & w2157;
assign w2159 = b_1 & w2158;
assign w2160 = ~w2154 & ~w2159;
assign w2161 = ~w1993 & ~w2157;
assign w2162 = ~w15 & w2161;
assign w2163 = w2160 & ~w2162;
assign w2164 = (a_26 & ~w2160) | (a_26 & w25362) | (~w2160 & w25362);
assign w2165 = w2160 & w25528;
assign w2166 = ~w2163 & ~w2164;
assign w2167 = (w2149 & w2166) | (w2149 & w25529) | (w2166 & w25529);
assign w2168 = ~w2166 & w26127;
assign w2169 = ~w2167 & ~w2168;
assign w2170 = w2148 & w2169;
assign w2171 = ~w2148 & ~w2169;
assign w2172 = ~w2170 & ~w2171;
assign w2173 = ~w2137 & ~w2172;
assign w2174 = w2137 & w2172;
assign w2175 = ~w2173 & ~w2174;
assign w2176 = ~w2135 & w2175;
assign w2177 = w2135 & ~w2175;
assign w2178 = ~w2176 & ~w2177;
assign w2179 = ~w2125 & w2178;
assign w2180 = w2125 & ~w2178;
assign w2181 = ~w2179 & ~w2180;
assign w2182 = b_10 & w986;
assign w2183 = w1069 & w28133;
assign w2184 = b_9 & w981;
assign w2185 = ~w2183 & ~w2184;
assign w2186 = ~w2182 & w2185;
assign w2187 = (w2186 & ~w454) | (w2186 & w28134) | (~w454 & w28134);
assign w2188 = (w454 & w38410) | (w454 & w38411) | (w38410 & w38411);
assign w2189 = (~w454 & w38412) | (~w454 & w38413) | (w38412 & w38413);
assign w2190 = ~w2187 & ~w2188;
assign w2191 = ~w2189 & ~w2190;
assign w2192 = w2181 & ~w2191;
assign w2193 = w2181 & ~w2192;
assign w2194 = ~w2181 & ~w2191;
assign w2195 = ~w2193 & ~w2194;
assign w2196 = (~w2029 & w1980) | (~w2029 & w26774) | (w1980 & w26774);
assign w2197 = w2195 & w2196;
assign w2198 = ~w2195 & ~w2196;
assign w2199 = ~w2197 & ~w2198;
assign w2200 = b_13 & w657;
assign w2201 = w754 & w28135;
assign w2202 = b_12 & w652;
assign w2203 = ~w2201 & ~w2202;
assign w2204 = ~w2200 & w2203;
assign w2205 = (w2204 & ~w711) | (w2204 & w28136) | (~w711 & w28136);
assign w2206 = (w711 & w38414) | (w711 & w38415) | (w38414 & w38415);
assign w2207 = (~w711 & w38416) | (~w711 & w38417) | (w38416 & w38417);
assign w2208 = ~w2205 & ~w2206;
assign w2209 = ~w2207 & ~w2208;
assign w2210 = ~w2199 & w2209;
assign w2211 = w2199 & ~w2209;
assign w2212 = ~w2210 & ~w2211;
assign w2213 = (~w2036 & w1969) | (~w2036 & w28137) | (w1969 & w28137);
assign w2214 = w2212 & ~w2213;
assign w2215 = ~w2212 & w2213;
assign w2216 = ~w2214 & ~w2215;
assign w2217 = ~w2124 & w2216;
assign w2218 = w2216 & ~w2217;
assign w2219 = ~w2216 & ~w2124;
assign w2220 = ~w2218 & ~w2219;
assign w2221 = ~w2041 & ~w2047;
assign w2222 = w2220 & w2221;
assign w2223 = ~w2220 & ~w2221;
assign w2224 = ~w2222 & ~w2223;
assign w2225 = b_19 & w239;
assign w2226 = w266 & w28138;
assign w2227 = b_18 & w234;
assign w2228 = ~w2226 & ~w2227;
assign w2229 = ~w2225 & w2228;
assign w2230 = (w2229 & ~w1372) | (w2229 & w28139) | (~w1372 & w28139);
assign w2231 = (w1372 & w38418) | (w1372 & w38419) | (w38418 & w38419);
assign w2232 = (~w1372 & w38420) | (~w1372 & w38421) | (w38420 & w38421);
assign w2233 = ~w2230 & ~w2231;
assign w2234 = ~w2232 & ~w2233;
assign w2235 = w2224 & ~w2234;
assign w2236 = w2224 & ~w2235;
assign w2237 = ~w2224 & ~w2234;
assign w2238 = ~w2236 & ~w2237;
assign w2239 = (~w2060 & w1958) | (~w2060 & w27402) | (w1958 & w27402);
assign w2240 = ~w2238 & ~w2239;
assign w2241 = ~w2238 & ~w2240;
assign w2242 = w2238 & ~w2239;
assign w2243 = b_22 & w99;
assign w2244 = w136 & w28140;
assign w2245 = b_21 & w94;
assign w2246 = ~w2244 & ~w2245;
assign w2247 = ~w2243 & w2246;
assign w2248 = (w2247 & ~w1786) | (w2247 & w28141) | (~w1786 & w28141);
assign w2249 = (w1786 & w38422) | (w1786 & w38423) | (w38422 & w38423);
assign w2250 = (~w1786 & w38424) | (~w1786 & w38425) | (w38424 & w38425);
assign w2251 = ~w2248 & ~w2249;
assign w2252 = ~w2250 & ~w2251;
assign w2253 = (w2252 & w2241) | (w2252 & w28142) | (w2241 & w28142);
assign w2254 = ~w2241 & w28143;
assign w2255 = ~w2253 & ~w2254;
assign w2256 = ~w2114 & ~w2255;
assign w2257 = w2114 & w2255;
assign w2258 = ~w2256 & ~w2257;
assign w2259 = ~w2113 & w2258;
assign w2260 = w2113 & ~w2258;
assign w2261 = ~w2259 & ~w2260;
assign w2262 = (~w28116 & w38426) | (~w28116 & w38427) | (w38426 & w38427);
assign w2263 = (w28116 & w38428) | (w28116 & w38429) | (w38428 & w38429);
assign w2264 = ~w2262 & ~w2263;
assign w2265 = (~w2259 & w2097) | (~w2259 & w28144) | (w2097 & w28144);
assign w2266 = (~w2252 & w2241) | (~w2252 & w28145) | (w2241 & w28145);
assign w2267 = ~w2256 & ~w2266;
assign w2268 = (~w2217 & w2221) | (~w2217 & w28146) | (w2221 & w28146);
assign w2269 = (~w2211 & w2213) | (~w2211 & w27403) | (w2213 & w27403);
assign w2270 = b_14 & w657;
assign w2271 = w754 & w28147;
assign w2272 = b_13 & w652;
assign w2273 = ~w2271 & ~w2272;
assign w2274 = ~w2270 & w2273;
assign w2275 = (w2274 & ~w735) | (w2274 & w28148) | (~w735 & w28148);
assign w2276 = (w735 & w38430) | (w735 & w38431) | (w38430 & w38431);
assign w2277 = (~w735 & w38432) | (~w735 & w38433) | (w38432 & w38433);
assign w2278 = ~w2275 & ~w2276;
assign w2279 = ~w2277 & ~w2278;
assign w2280 = b_11 & w986;
assign w2281 = w1069 & w28149;
assign w2282 = b_10 & w981;
assign w2283 = ~w2281 & ~w2282;
assign w2284 = ~w2280 & w2283;
assign w2285 = (w2284 & ~w530) | (w2284 & w28150) | (~w530 & w28150);
assign w2286 = (w530 & w38434) | (w530 & w38435) | (w38434 & w38435);
assign w2287 = (~w530 & w38436) | (~w530 & w38437) | (w38436 & w38437);
assign w2288 = ~w2285 & ~w2286;
assign w2289 = ~w2287 & ~w2288;
assign w2290 = (~w2176 & w2125) | (~w2176 & w28151) | (w2125 & w28151);
assign w2291 = ~w2148 & w2169;
assign w2292 = (~w2291 & w2137) | (~w2291 & w26775) | (w2137 & w26775);
assign w2293 = b_2 & w2158;
assign w2294 = w1993 & ~w2157;
assign w2295 = w2294 & w24989;
assign w2296 = b_1 & w2153;
assign w2297 = ~w2295 & ~w2296;
assign w2298 = ~w2293 & w2297;
assign w2299 = w35 & w2161;
assign w2300 = w2298 & ~w2299;
assign w2301 = (a_26 & ~w2298) | (a_26 & w24990) | (~w2298 & w24990);
assign w2302 = w2298 & w25363;
assign w2303 = ~w2300 & ~w2301;
assign w2304 = ~w2302 & ~w2303;
assign w2305 = ~w2167 & w2304;
assign w2306 = w2167 & ~w2304;
assign w2307 = ~w2305 & ~w2306;
assign w2308 = b_5 & w1694;
assign w2309 = w1834 & w28152;
assign w2310 = b_4 & w1689;
assign w2311 = ~w2309 & ~w2310;
assign w2312 = ~w2308 & w2311;
assign w2313 = w129 & w1697;
assign w2314 = w2312 & ~w2313;
assign w2315 = (a_23 & w2313) | (a_23 & w28153) | (w2313 & w28153);
assign w2316 = ~w2313 & w38438;
assign w2317 = ~w2314 & ~w2315;
assign w2318 = ~w2316 & ~w2317;
assign w2319 = w2307 & ~w2318;
assign w2320 = ~w2307 & w2318;
assign w2321 = (w2173 & w25775) | (w2173 & w25776) | (w25775 & w25776);
assign w2322 = ~w2292 & ~w2321;
assign w2323 = (~w25776 & w28154) | (~w25776 & w28155) | (w28154 & w28155);
assign w2324 = ~w25776 & w28156;
assign w2325 = b_8 & w1295;
assign w2326 = w1422 & w28157;
assign w2327 = b_7 & w1290;
assign w2328 = ~w2326 & ~w2327;
assign w2329 = ~w2325 & w2328;
assign w2330 = ~w308 & w28158;
assign w2331 = (w2329 & ~w28158) | (w2329 & w38439) | (~w28158 & w38439);
assign w2332 = (w28158 & w38440) | (w28158 & w38441) | (w38440 & w38441);
assign w2333 = ~w2330 & w28160;
assign w2334 = ~w2331 & ~w2332;
assign w2335 = ~w2333 & ~w2334;
assign w2336 = ~w2322 & w28161;
assign w2337 = (~w2335 & w2322) | (~w2335 & w28162) | (w2322 & w28162);
assign w2338 = ~w2336 & ~w2337;
assign w2339 = ~w2290 & w2338;
assign w2340 = w2290 & ~w2338;
assign w2341 = ~w2339 & ~w2340;
assign w2342 = w2289 & ~w2341;
assign w2343 = ~w2289 & w2341;
assign w2344 = ~w2342 & ~w2343;
assign w2345 = (w2344 & w2198) | (w2344 & w24992) | (w2198 & w24992);
assign w2346 = ~w2198 & w28163;
assign w2347 = ~w2345 & ~w2346;
assign w2348 = ~w2279 & w2347;
assign w2349 = w2347 & ~w2348;
assign w2350 = ~w2347 & ~w2279;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = ~w2269 & w2351;
assign w2353 = w2269 & ~w2351;
assign w2354 = ~w2352 & ~w2353;
assign w2355 = b_17 & w418;
assign w2356 = w481 & w28164;
assign w2357 = b_16 & w413;
assign w2358 = ~w2356 & ~w2357;
assign w2359 = ~w2355 & w2358;
assign w2360 = (w2359 & ~w1038) | (w2359 & w28165) | (~w1038 & w28165);
assign w2361 = (w1038 & w38442) | (w1038 & w38443) | (w38442 & w38443);
assign w2362 = (~w1038 & w38444) | (~w1038 & w38445) | (w38444 & w38445);
assign w2363 = ~w2360 & ~w2361;
assign w2364 = ~w2362 & ~w2363;
assign w2365 = ~w2354 & ~w2364;
assign w2366 = w2354 & w2364;
assign w2367 = ~w2365 & ~w2366;
assign w2368 = w2268 & ~w2367;
assign w2369 = (w2367 & w2223) | (w2367 & w24993) | (w2223 & w24993);
assign w2370 = ~w2368 & ~w2369;
assign w2371 = b_20 & w239;
assign w2372 = w266 & w28166;
assign w2373 = b_19 & w234;
assign w2374 = ~w2372 & ~w2373;
assign w2375 = ~w2371 & w2374;
assign w2376 = (w2375 & ~w1503) | (w2375 & w28167) | (~w1503 & w28167);
assign w2377 = (w1503 & w38446) | (w1503 & w38447) | (w38446 & w38447);
assign w2378 = (~w1503 & w38448) | (~w1503 & w38449) | (w38448 & w38449);
assign w2379 = ~w2376 & ~w2377;
assign w2380 = ~w2378 & ~w2379;
assign w2381 = w2370 & ~w2380;
assign w2382 = w2370 & ~w2381;
assign w2383 = ~w2370 & ~w2380;
assign w2384 = ~w2382 & ~w2383;
assign w2385 = (~w2235 & w2238) | (~w2235 & w27404) | (w2238 & w27404);
assign w2386 = w2384 & w2385;
assign w2387 = ~w2384 & ~w2385;
assign w2388 = ~w2386 & ~w2387;
assign w2389 = b_23 & w99;
assign w2390 = w136 & w28168;
assign w2391 = b_22 & w94;
assign w2392 = ~w2390 & ~w2391;
assign w2393 = ~w2389 & w2392;
assign w2394 = (w2393 & ~w1933) | (w2393 & w28169) | (~w1933 & w28169);
assign w2395 = (w1933 & w38450) | (w1933 & w38451) | (w38450 & w38451);
assign w2396 = (~w1933 & w38452) | (~w1933 & w38453) | (w38452 & w38453);
assign w2397 = ~w2394 & ~w2395;
assign w2398 = ~w2396 & ~w2397;
assign w2399 = w2388 & ~w2398;
assign w2400 = w2388 & ~w2399;
assign w2401 = ~w2388 & ~w2398;
assign w2402 = ~w2400 & ~w2401;
assign w2403 = ~w2267 & w2402;
assign w2404 = w2267 & ~w2402;
assign w2405 = ~w2403 & ~w2404;
assign w2406 = w8 & w28170;
assign w2407 = ~w8 & w28171;
assign w2408 = b_25 & w4;
assign w2409 = ~w2407 & ~w2408;
assign w2410 = ~w2406 & w2409;
assign w2411 = ~b_25 & ~b_26;
assign w2412 = b_25 & b_26;
assign w2413 = ~w2411 & ~w2412;
assign w2414 = (w1931 & w28174) | (w1931 & w28175) | (w28174 & w28175);
assign w2415 = (~w1931 & w28176) | (~w1931 & w28177) | (w28176 & w28177);
assign w2416 = ~w2414 & ~w2415;
assign w2417 = (w2410 & ~w2416) | (w2410 & w28178) | (~w2416 & w28178);
assign w2418 = (w2416 & w38454) | (w2416 & w38455) | (w38454 & w38455);
assign w2419 = (~w2416 & w38456) | (~w2416 & w38457) | (w38456 & w38457);
assign w2420 = ~w2417 & ~w2418;
assign w2421 = ~w2419 & ~w2420;
assign w2422 = ~w2405 & ~w2421;
assign w2423 = w2405 & w2421;
assign w2424 = ~w2422 & ~w2423;
assign w2425 = ~w2265 & w2424;
assign w2426 = w2265 & ~w2424;
assign w2427 = ~w2425 & ~w2426;
assign w2428 = (~w2422 & w2265) | (~w2422 & w38458) | (w2265 & w38458);
assign w2429 = b_24 & w99;
assign w2430 = w136 & w28179;
assign w2431 = b_23 & w94;
assign w2432 = ~w2430 & ~w2431;
assign w2433 = ~w2429 & w2432;
assign w2434 = (w2433 & ~w2083) | (w2433 & w28180) | (~w2083 & w28180);
assign w2435 = (w2083 & w38459) | (w2083 & w38460) | (w38459 & w38460);
assign w2436 = (~w2083 & w38461) | (~w2083 & w38462) | (w38461 & w38462);
assign w2437 = ~w2434 & ~w2435;
assign w2438 = ~w2436 & ~w2437;
assign w2439 = b_15 & w657;
assign w2440 = w754 & w28181;
assign w2441 = b_14 & w652;
assign w2442 = ~w2440 & ~w2441;
assign w2443 = ~w2439 & w2442;
assign w2444 = (w2443 & ~w827) | (w2443 & w28182) | (~w827 & w28182);
assign w2445 = (w827 & w38463) | (w827 & w38464) | (w38463 & w38464);
assign w2446 = (~w827 & w38465) | (~w827 & w38466) | (w38465 & w38466);
assign w2447 = ~w2444 & ~w2445;
assign w2448 = ~w2446 & ~w2447;
assign w2449 = (~w24992 & w26776) | (~w24992 & w26777) | (w26776 & w26777);
assign w2450 = b_12 & w986;
assign w2451 = w1069 & w28183;
assign w2452 = b_11 & w981;
assign w2453 = ~w2451 & ~w2452;
assign w2454 = ~w2450 & w2453;
assign w2455 = (w2454 & ~w552) | (w2454 & w28184) | (~w552 & w28184);
assign w2456 = (w552 & w38467) | (w552 & w38468) | (w38467 & w38468);
assign w2457 = (~w552 & w38469) | (~w552 & w38470) | (w38469 & w38470);
assign w2458 = ~w2455 & ~w2456;
assign w2459 = ~w2457 & ~w2458;
assign w2460 = ~w2337 & ~w2339;
assign w2461 = b_6 & w1694;
assign w2462 = w1834 & w28185;
assign w2463 = b_5 & w1689;
assign w2464 = ~w2462 & ~w2463;
assign w2465 = ~w2461 & w2464;
assign w2466 = (w2465 & ~w190) | (w2465 & w28186) | (~w190 & w28186);
assign w2467 = (w190 & w38471) | (w190 & w38472) | (w38471 & w38472);
assign w2468 = (~w190 & w38473) | (~w190 & w38474) | (w38473 & w38474);
assign w2469 = ~w2466 & ~w2467;
assign w2470 = ~w2468 & ~w2469;
assign w2471 = a_26 & ~a_27;
assign w2472 = ~a_26 & a_27;
assign w2473 = ~w2471 & ~w2472;
assign w2474 = b_0 & ~w2473;
assign w2475 = (w2474 & ~w2167) | (w2474 & w24994) | (~w2167 & w24994);
assign w2476 = w2167 & w24995;
assign w2477 = ~w2475 & ~w2476;
assign w2478 = b_3 & w2158;
assign w2479 = w2294 & w25530;
assign w2480 = b_2 & w2153;
assign w2481 = ~w2479 & ~w2480;
assign w2482 = ~w2478 & w2481;
assign w2483 = w57 & w2161;
assign w2484 = w2482 & ~w2483;
assign w2485 = a_26 & ~w2484;
assign w2486 = w2484 & a_26;
assign w2487 = ~w2484 & ~w2485;
assign w2488 = ~w2486 & ~w2487;
assign w2489 = ~w2477 & ~w2488;
assign w2490 = w2477 & w2488;
assign w2491 = ~w2489 & ~w2490;
assign w2492 = ~w2470 & w2491;
assign w2493 = w2491 & ~w2492;
assign w2494 = ~w2491 & ~w2470;
assign w2495 = ~w2493 & ~w2494;
assign w2496 = ~w2323 & w2495;
assign w2497 = w2323 & ~w2495;
assign w2498 = ~w2496 & ~w2497;
assign w2499 = b_9 & w1295;
assign w2500 = w1422 & w28187;
assign w2501 = b_8 & w1290;
assign w2502 = ~w2500 & ~w2501;
assign w2503 = ~w2499 & w2502;
assign w2504 = (w2503 & ~w371) | (w2503 & w28188) | (~w371 & w28188);
assign w2505 = (w371 & w38475) | (w371 & w38476) | (w38475 & w38476);
assign w2506 = (~w371 & w38477) | (~w371 & w38478) | (w38477 & w38478);
assign w2507 = ~w2504 & ~w2505;
assign w2508 = ~w2506 & ~w2507;
assign w2509 = ~w2498 & ~w2508;
assign w2510 = w2498 & w2508;
assign w2511 = ~w2509 & ~w2510;
assign w2512 = ~w2460 & w2511;
assign w2513 = w2460 & ~w2511;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = w2459 & ~w2514;
assign w2516 = ~w2459 & w2514;
assign w2517 = ~w2515 & ~w2516;
assign w2518 = ~w2449 & w2517;
assign w2519 = w2449 & ~w2517;
assign w2520 = ~w2518 & ~w2519;
assign w2521 = ~w2448 & w2520;
assign w2522 = w2520 & ~w2521;
assign w2523 = ~w2520 & ~w2448;
assign w2524 = ~w2522 & ~w2523;
assign w2525 = (~w2348 & w2269) | (~w2348 & w24996) | (w2269 & w24996);
assign w2526 = w2524 & w2525;
assign w2527 = ~w2524 & ~w2525;
assign w2528 = ~w2526 & ~w2527;
assign w2529 = b_18 & w418;
assign w2530 = w481 & w28189;
assign w2531 = b_17 & w413;
assign w2532 = ~w2530 & ~w2531;
assign w2533 = ~w2529 & w2532;
assign w2534 = (w2533 & ~w1238) | (w2533 & w24997) | (~w1238 & w24997);
assign w2535 = (w1238 & w28190) | (w1238 & w28191) | (w28190 & w28191);
assign w2536 = (~w1238 & w28192) | (~w1238 & w28193) | (w28192 & w28193);
assign w2537 = ~w2534 & ~w2535;
assign w2538 = ~w2536 & ~w2537;
assign w2539 = w2528 & ~w2538;
assign w2540 = w2528 & ~w2539;
assign w2541 = ~w2528 & ~w2538;
assign w2542 = ~w2540 & ~w2541;
assign w2543 = ~w2365 & ~w2369;
assign w2544 = w2542 & w2543;
assign w2545 = ~w2542 & ~w2543;
assign w2546 = ~w2544 & ~w2545;
assign w2547 = b_21 & w239;
assign w2548 = w266 & w28194;
assign w2549 = b_20 & w234;
assign w2550 = ~w2548 & ~w2549;
assign w2551 = ~w2547 & w2550;
assign w2552 = (w2551 & ~w1634) | (w2551 & w28195) | (~w1634 & w28195);
assign w2553 = (w1634 & w38479) | (w1634 & w38480) | (w38479 & w38480);
assign w2554 = (~w1634 & w38481) | (~w1634 & w38482) | (w38481 & w38482);
assign w2555 = ~w2552 & ~w2553;
assign w2556 = ~w2554 & ~w2555;
assign w2557 = ~w2546 & w2556;
assign w2558 = w2546 & ~w2556;
assign w2559 = ~w2557 & ~w2558;
assign w2560 = (~w2381 & w2384) | (~w2381 & w27405) | (w2384 & w27405);
assign w2561 = w2559 & ~w2560;
assign w2562 = ~w2559 & w2560;
assign w2563 = ~w2561 & ~w2562;
assign w2564 = ~w2438 & w2563;
assign w2565 = w2563 & ~w2564;
assign w2566 = ~w2563 & ~w2438;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = (~w2399 & w2267) | (~w2399 & w28196) | (w2267 & w28196);
assign w2569 = w2567 & w2568;
assign w2570 = ~w2567 & ~w2568;
assign w2571 = ~w2569 & ~w2570;
assign w2572 = w8 & w28197;
assign w2573 = ~w8 & w28198;
assign w2574 = b_26 & w4;
assign w2575 = ~w2573 & ~w2574;
assign w2576 = ~w2572 & w2575;
assign w2577 = ~b_26 & ~b_27;
assign w2578 = b_26 & b_27;
assign w2579 = ~w2577 & ~w2578;
assign w2580 = (w1931 & w28200) | (w1931 & w28201) | (w28200 & w28201);
assign w2581 = (~w1931 & w28202) | (~w1931 & w28203) | (w28202 & w28203);
assign w2582 = ~w2580 & ~w2581;
assign w2583 = (w2576 & ~w2582) | (w2576 & w28204) | (~w2582 & w28204);
assign w2584 = (w2582 & w38483) | (w2582 & w38484) | (w38483 & w38484);
assign w2585 = (~w2582 & w38485) | (~w2582 & w38486) | (w38485 & w38486);
assign w2586 = ~w2583 & ~w2584;
assign w2587 = ~w2585 & ~w2586;
assign w2588 = ~w2571 & w2587;
assign w2589 = w2571 & ~w2587;
assign w2590 = ~w2588 & ~w2589;
assign w2591 = ~w2428 & w2590;
assign w2592 = w2428 & ~w2590;
assign w2593 = ~w2591 & ~w2592;
assign w2594 = (~w2589 & w2428) | (~w2589 & w28205) | (w2428 & w28205);
assign w2595 = b_25 & w99;
assign w2596 = w136 & w28206;
assign w2597 = b_24 & w94;
assign w2598 = ~w2596 & ~w2597;
assign w2599 = ~w2595 & w2598;
assign w2600 = (w2599 & ~w2108) | (w2599 & w28207) | (~w2108 & w28207);
assign w2601 = (w2108 & w38487) | (w2108 & w38488) | (w38487 & w38488);
assign w2602 = (~w2108 & w38489) | (~w2108 & w38490) | (w38489 & w38490);
assign w2603 = ~w2600 & ~w2601;
assign w2604 = ~w2602 & ~w2603;
assign w2605 = ~w2323 & ~w2495;
assign w2606 = (~w2492 & w2495) | (~w2492 & w28208) | (w2495 & w28208);
assign w2607 = b_7 & w1694;
assign w2608 = w1834 & w28209;
assign w2609 = b_6 & w1689;
assign w2610 = ~w2608 & ~w2609;
assign w2611 = ~w2607 & w2610;
assign w2612 = (w2611 & ~w213) | (w2611 & w28210) | (~w213 & w28210);
assign w2613 = (w213 & w38491) | (w213 & w38492) | (w38491 & w38492);
assign w2614 = (~w213 & w38493) | (~w213 & w38494) | (w38493 & w38494);
assign w2615 = ~w2612 & ~w2613;
assign w2616 = ~w2614 & ~w2615;
assign w2617 = ~w2304 & w25531;
assign w2618 = (~w2617 & w2477) | (~w2617 & w25364) | (w2477 & w25364);
assign w2619 = b_4 & w2158;
assign w2620 = w2294 & w25532;
assign w2621 = b_3 & w2153;
assign w2622 = ~w2620 & ~w2621;
assign w2623 = ~w2619 & w2622;
assign w2624 = w84 & w2161;
assign w2625 = w2623 & ~w2624;
assign w2626 = (a_26 & w2624) | (a_26 & w24998) | (w2624 & w24998);
assign w2627 = ~w2624 & w25533;
assign w2628 = ~w2625 & ~w2626;
assign w2629 = ~w2627 & ~w2628;
assign w2630 = (a_29 & w2473) | (a_29 & w28211) | (w2473 & w28211);
assign w2631 = ~a_27 & a_28;
assign w2632 = a_27 & ~a_28;
assign w2633 = ~w2631 & ~w2632;
assign w2634 = w2473 & ~w2633;
assign w2635 = b_0 & w2634;
assign w2636 = ~a_28 & a_29;
assign w2637 = a_28 & ~a_29;
assign w2638 = ~w2636 & ~w2637;
assign w2639 = ~w2473 & w2638;
assign w2640 = b_1 & w2639;
assign w2641 = ~w2635 & ~w2640;
assign w2642 = ~w2473 & ~w2638;
assign w2643 = ~w15 & w2642;
assign w2644 = w2641 & ~w2643;
assign w2645 = (a_29 & ~w2641) | (a_29 & w25365) | (~w2641 & w25365);
assign w2646 = w2641 & w25534;
assign w2647 = ~w2644 & ~w2645;
assign w2648 = (w2630 & w2647) | (w2630 & w25535) | (w2647 & w25535);
assign w2649 = ~w2647 & w25536;
assign w2650 = ~w2648 & ~w2649;
assign w2651 = w2629 & w2650;
assign w2652 = ~w2629 & ~w2650;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = ~w2618 & ~w2653;
assign w2655 = w2618 & w2653;
assign w2656 = ~w2654 & ~w2655;
assign w2657 = ~w2616 & w2656;
assign w2658 = w2616 & ~w2656;
assign w2659 = ~w2657 & ~w2658;
assign w2660 = (w2659 & w2605) | (w2659 & w26537) | (w2605 & w26537);
assign w2661 = ~w2605 & w26538;
assign w2662 = ~w2660 & ~w2661;
assign w2663 = b_10 & w1295;
assign w2664 = w1422 & w28212;
assign w2665 = b_9 & w1290;
assign w2666 = ~w2664 & ~w2665;
assign w2667 = ~w2663 & w2666;
assign w2668 = (w2667 & ~w454) | (w2667 & w28213) | (~w454 & w28213);
assign w2669 = (w454 & w38495) | (w454 & w38496) | (w38495 & w38496);
assign w2670 = (~w454 & w38497) | (~w454 & w38498) | (w38497 & w38498);
assign w2671 = ~w2668 & ~w2669;
assign w2672 = ~w2670 & ~w2671;
assign w2673 = w2662 & ~w2672;
assign w2674 = w2662 & ~w2673;
assign w2675 = ~w2662 & ~w2672;
assign w2676 = ~w2674 & ~w2675;
assign w2677 = (~w2509 & w2460) | (~w2509 & w24999) | (w2460 & w24999);
assign w2678 = w2676 & w2677;
assign w2679 = ~w2676 & ~w2677;
assign w2680 = ~w2678 & ~w2679;
assign w2681 = b_13 & w986;
assign w2682 = w1069 & w28214;
assign w2683 = b_12 & w981;
assign w2684 = ~w2682 & ~w2683;
assign w2685 = ~w2681 & w2684;
assign w2686 = (w2685 & ~w711) | (w2685 & w25000) | (~w711 & w25000);
assign w2687 = (w711 & w28215) | (w711 & w28216) | (w28215 & w28216);
assign w2688 = (~w711 & w28217) | (~w711 & w28218) | (w28217 & w28218);
assign w2689 = ~w2686 & ~w2687;
assign w2690 = ~w2688 & ~w2689;
assign w2691 = w2680 & ~w2690;
assign w2692 = w2680 & ~w2691;
assign w2693 = ~w2680 & ~w2690;
assign w2694 = ~w2692 & ~w2693;
assign w2695 = (~w2516 & w2449) | (~w2516 & w25001) | (w2449 & w25001);
assign w2696 = ~w2694 & ~w2695;
assign w2697 = ~w2694 & ~w2696;
assign w2698 = w2694 & ~w2695;
assign w2699 = ~w2697 & ~w2698;
assign w2700 = b_16 & w657;
assign w2701 = w754 & w28219;
assign w2702 = b_15 & w652;
assign w2703 = ~w2701 & ~w2702;
assign w2704 = ~w2700 & w2703;
assign w2705 = (w2704 & ~w926) | (w2704 & w25002) | (~w926 & w25002);
assign w2706 = (w926 & w28220) | (w926 & w28221) | (w28220 & w28221);
assign w2707 = (~w926 & w28222) | (~w926 & w28223) | (w28222 & w28223);
assign w2708 = ~w2705 & ~w2706;
assign w2709 = ~w2707 & ~w2708;
assign w2710 = (~w2709 & w2697) | (~w2709 & w28224) | (w2697 & w28224);
assign w2711 = ~w2699 & ~w2710;
assign w2712 = ~w2697 & w28225;
assign w2713 = ~w2711 & ~w2712;
assign w2714 = (~w2521 & w2524) | (~w2521 & w28226) | (w2524 & w28226);
assign w2715 = w2713 & w2714;
assign w2716 = ~w2713 & ~w2714;
assign w2717 = ~w2715 & ~w2716;
assign w2718 = b_19 & w418;
assign w2719 = w481 & w28227;
assign w2720 = b_18 & w413;
assign w2721 = ~w2719 & ~w2720;
assign w2722 = ~w2718 & w2721;
assign w2723 = (w2722 & ~w1372) | (w2722 & w25003) | (~w1372 & w25003);
assign w2724 = (w1372 & w28228) | (w1372 & w28229) | (w28228 & w28229);
assign w2725 = (~w1372 & w28230) | (~w1372 & w28231) | (w28230 & w28231);
assign w2726 = ~w2723 & ~w2724;
assign w2727 = ~w2725 & ~w2726;
assign w2728 = w2717 & ~w2727;
assign w2729 = w2717 & ~w2728;
assign w2730 = ~w2717 & ~w2727;
assign w2731 = ~w2729 & ~w2730;
assign w2732 = (~w2539 & w2543) | (~w2539 & w25004) | (w2543 & w25004);
assign w2733 = w2731 & w2732;
assign w2734 = ~w2731 & ~w2732;
assign w2735 = ~w2733 & ~w2734;
assign w2736 = b_22 & w239;
assign w2737 = w266 & w28232;
assign w2738 = b_21 & w234;
assign w2739 = ~w2737 & ~w2738;
assign w2740 = ~w2736 & w2739;
assign w2741 = (w2740 & ~w1786) | (w2740 & w28233) | (~w1786 & w28233);
assign w2742 = (w1786 & w38499) | (w1786 & w38500) | (w38499 & w38500);
assign w2743 = (~w1786 & w38501) | (~w1786 & w38502) | (w38501 & w38502);
assign w2744 = ~w2741 & ~w2742;
assign w2745 = ~w2743 & ~w2744;
assign w2746 = ~w2735 & w2745;
assign w2747 = w2735 & ~w2745;
assign w2748 = ~w2746 & ~w2747;
assign w2749 = (~w2558 & w2560) | (~w2558 & w28234) | (w2560 & w28234);
assign w2750 = w2748 & ~w2749;
assign w2751 = ~w2748 & w2749;
assign w2752 = ~w2750 & ~w2751;
assign w2753 = ~w2604 & w2752;
assign w2754 = w2752 & ~w2753;
assign w2755 = ~w2752 & ~w2604;
assign w2756 = ~w2754 & ~w2755;
assign w2757 = (~w2564 & w2567) | (~w2564 & w38503) | (w2567 & w38503);
assign w2758 = w2756 & w2757;
assign w2759 = ~w2756 & ~w2757;
assign w2760 = ~w2758 & ~w2759;
assign w2761 = w8 & w28235;
assign w2762 = ~w8 & w28236;
assign w2763 = b_27 & w4;
assign w2764 = ~w2762 & ~w2763;
assign w2765 = ~w2761 & w2764;
assign w2766 = ~b_27 & ~b_28;
assign w2767 = b_27 & b_28;
assign w2768 = ~w2766 & ~w2767;
assign w2769 = (w1931 & w38504) | (w1931 & w38505) | (w38504 & w38505);
assign w2770 = (~w1931 & w38506) | (~w1931 & w38507) | (w38506 & w38507);
assign w2771 = ~w2769 & ~w2770;
assign w2772 = (w2765 & ~w2771) | (w2765 & w28239) | (~w2771 & w28239);
assign w2773 = (w2771 & w38508) | (w2771 & w38509) | (w38508 & w38509);
assign w2774 = (~w2771 & w38510) | (~w2771 & w38511) | (w38510 & w38511);
assign w2775 = ~w2772 & ~w2773;
assign w2776 = ~w2774 & ~w2775;
assign w2777 = ~w2760 & w2776;
assign w2778 = w2760 & ~w2776;
assign w2779 = ~w2777 & ~w2778;
assign w2780 = ~w2594 & w2779;
assign w2781 = w2594 & ~w2779;
assign w2782 = ~w2780 & ~w2781;
assign w2783 = (~w2753 & w2757) | (~w2753 & w28240) | (w2757 & w28240);
assign w2784 = b_26 & w99;
assign w2785 = w136 & w28241;
assign w2786 = b_25 & w94;
assign w2787 = ~w2785 & ~w2786;
assign w2788 = ~w2784 & w2787;
assign w2789 = (w2788 & ~w2416) | (w2788 & w28242) | (~w2416 & w28242);
assign w2790 = (w2416 & w38512) | (w2416 & w38513) | (w38512 & w38513);
assign w2791 = (~w2416 & w38514) | (~w2416 & w38515) | (w38514 & w38515);
assign w2792 = ~w2789 & ~w2790;
assign w2793 = ~w2791 & ~w2792;
assign w2794 = (~w2728 & w2731) | (~w2728 & w27406) | (w2731 & w27406);
assign w2795 = b_14 & w986;
assign w2796 = w1069 & w28243;
assign w2797 = b_13 & w981;
assign w2798 = ~w2796 & ~w2797;
assign w2799 = ~w2795 & w2798;
assign w2800 = (w2799 & ~w735) | (w2799 & w28244) | (~w735 & w28244);
assign w2801 = (w735 & w38516) | (w735 & w38517) | (w38516 & w38517);
assign w2802 = (~w735 & w38518) | (~w735 & w38519) | (w38518 & w38519);
assign w2803 = ~w2800 & ~w2801;
assign w2804 = ~w2802 & ~w2803;
assign w2805 = ~w2673 & ~w2679;
assign w2806 = b_11 & w1295;
assign w2807 = w1422 & w28245;
assign w2808 = b_10 & w1290;
assign w2809 = ~w2807 & ~w2808;
assign w2810 = ~w2806 & w2809;
assign w2811 = (w2810 & ~w530) | (w2810 & w28246) | (~w530 & w28246);
assign w2812 = (w530 & w38520) | (w530 & w38521) | (w38520 & w38521);
assign w2813 = (~w530 & w38522) | (~w530 & w38523) | (w38522 & w38523);
assign w2814 = ~w2811 & ~w2812;
assign w2815 = ~w2813 & ~w2814;
assign w2816 = (~w2657 & w2606) | (~w2657 & w25005) | (w2606 & w25005);
assign w2817 = ~w2629 & w2650;
assign w2818 = (~w2817 & w2618) | (~w2817 & w25006) | (w2618 & w25006);
assign w2819 = b_2 & w2639;
assign w2820 = w2473 & ~w2638;
assign w2821 = w2820 & w25007;
assign w2822 = b_1 & w2634;
assign w2823 = ~w2821 & ~w2822;
assign w2824 = ~w2819 & w2823;
assign w2825 = w35 & w2642;
assign w2826 = w2824 & ~w2825;
assign w2827 = (a_29 & ~w2824) | (a_29 & w25366) | (~w2824 & w25366);
assign w2828 = w2824 & w25537;
assign w2829 = ~w2826 & ~w2827;
assign w2830 = ~w2828 & ~w2829;
assign w2831 = ~w2648 & w2830;
assign w2832 = w2648 & ~w2830;
assign w2833 = ~w2831 & ~w2832;
assign w2834 = b_5 & w2158;
assign w2835 = w2294 & w26128;
assign w2836 = b_4 & w2153;
assign w2837 = ~w2835 & ~w2836;
assign w2838 = ~w2834 & w2837;
assign w2839 = w129 & w2161;
assign w2840 = w2838 & ~w2839;
assign w2841 = (a_26 & w2839) | (a_26 & w26129) | (w2839 & w26129);
assign w2842 = ~w2839 & w38524;
assign w2843 = ~w2840 & ~w2841;
assign w2844 = ~w2842 & ~w2843;
assign w2845 = w2833 & ~w2844;
assign w2846 = ~w2833 & w2844;
assign w2847 = ~w2818 & w25538;
assign w2848 = ~w2818 & ~w2847;
assign w2849 = (~w2845 & w2818) | (~w2845 & w25777) | (w2818 & w25777);
assign w2850 = ~w2846 & w2849;
assign w2851 = ~w2848 & ~w2850;
assign w2852 = b_8 & w1694;
assign w2853 = w1834 & w28247;
assign w2854 = b_7 & w1689;
assign w2855 = ~w2853 & ~w2854;
assign w2856 = ~w2852 & w2855;
assign w2857 = ~w308 & w28248;
assign w2858 = (w2856 & ~w28248) | (w2856 & w38525) | (~w28248 & w38525);
assign w2859 = (w28248 & w38526) | (w28248 & w38527) | (w38526 & w38527);
assign w2860 = ~w2857 & w28250;
assign w2861 = ~w2858 & ~w2859;
assign w2862 = ~w2860 & ~w2861;
assign w2863 = w2851 & w2862;
assign w2864 = ~w2851 & ~w2862;
assign w2865 = ~w2863 & ~w2864;
assign w2866 = ~w2816 & w2865;
assign w2867 = w2816 & ~w2865;
assign w2868 = ~w2866 & ~w2867;
assign w2869 = w2815 & ~w2868;
assign w2870 = ~w2815 & w2868;
assign w2871 = ~w2869 & ~w2870;
assign w2872 = ~w2805 & w2871;
assign w2873 = w2805 & ~w2871;
assign w2874 = ~w2872 & ~w2873;
assign w2875 = ~w2804 & w2874;
assign w2876 = w2874 & ~w2875;
assign w2877 = ~w2874 & ~w2804;
assign w2878 = ~w2876 & ~w2877;
assign w2879 = (~w2691 & w2694) | (~w2691 & w28251) | (w2694 & w28251);
assign w2880 = w2878 & w2879;
assign w2881 = ~w2878 & ~w2879;
assign w2882 = ~w2880 & ~w2881;
assign w2883 = b_17 & w657;
assign w2884 = w754 & w28252;
assign w2885 = b_16 & w652;
assign w2886 = ~w2884 & ~w2885;
assign w2887 = ~w2883 & w2886;
assign w2888 = (w2887 & ~w1038) | (w2887 & w25008) | (~w1038 & w25008);
assign w2889 = (w1038 & w28253) | (w1038 & w28254) | (w28253 & w28254);
assign w2890 = (~w1038 & w28255) | (~w1038 & w28256) | (w28255 & w28256);
assign w2891 = ~w2888 & ~w2889;
assign w2892 = ~w2890 & ~w2891;
assign w2893 = w2882 & ~w2892;
assign w2894 = w2882 & ~w2893;
assign w2895 = ~w2882 & ~w2892;
assign w2896 = ~w2894 & ~w2895;
assign w2897 = (~w2710 & w2714) | (~w2710 & w25009) | (w2714 & w25009);
assign w2898 = w2896 & w2897;
assign w2899 = ~w2896 & ~w2897;
assign w2900 = ~w2898 & ~w2899;
assign w2901 = b_20 & w418;
assign w2902 = w481 & w28257;
assign w2903 = b_19 & w413;
assign w2904 = ~w2902 & ~w2903;
assign w2905 = ~w2901 & w2904;
assign w2906 = (w2905 & ~w1503) | (w2905 & w28258) | (~w1503 & w28258);
assign w2907 = (w1503 & w38528) | (w1503 & w38529) | (w38528 & w38529);
assign w2908 = (~w1503 & w38530) | (~w1503 & w38531) | (w38530 & w38531);
assign w2909 = ~w2906 & ~w2907;
assign w2910 = ~w2908 & ~w2909;
assign w2911 = w2900 & ~w2910;
assign w2912 = ~w2900 & w2910;
assign w2913 = (w2734 & w27205) | (w2734 & w27206) | (w27205 & w27206);
assign w2914 = ~w2794 & ~w2913;
assign w2915 = (~w27206 & w28259) | (~w27206 & w28260) | (w28259 & w28260);
assign w2916 = ~w27206 & w28261;
assign w2917 = ~w2914 & ~w2916;
assign w2918 = b_23 & w239;
assign w2919 = w266 & w28262;
assign w2920 = b_22 & w234;
assign w2921 = ~w2919 & ~w2920;
assign w2922 = ~w2918 & w2921;
assign w2923 = (w2922 & ~w1933) | (w2922 & w28263) | (~w1933 & w28263);
assign w2924 = (w1933 & w38532) | (w1933 & w38533) | (w38532 & w38533);
assign w2925 = (~w1933 & w38534) | (~w1933 & w38535) | (w38534 & w38535);
assign w2926 = ~w2923 & ~w2924;
assign w2927 = ~w2925 & ~w2926;
assign w2928 = (~w2927 & w2914) | (~w2927 & w28264) | (w2914 & w28264);
assign w2929 = ~w2917 & ~w2928;
assign w2930 = ~w2914 & w28265;
assign w2931 = ~w2929 & ~w2930;
assign w2932 = ~w2747 & ~w2750;
assign w2933 = ~w2931 & ~w2932;
assign w2934 = w2931 & w2932;
assign w2935 = ~w2933 & ~w2934;
assign w2936 = ~w2793 & w2935;
assign w2937 = ~w2935 & ~w2793;
assign w2938 = w2935 & ~w2936;
assign w2939 = ~w2937 & ~w2938;
assign w2940 = ~w2783 & ~w2939;
assign w2941 = w2939 & ~w2783;
assign w2942 = ~w2939 & ~w2940;
assign w2943 = ~w2941 & ~w2942;
assign w2944 = w8 & w28266;
assign w2945 = ~w8 & w28267;
assign w2946 = b_28 & w4;
assign w2947 = ~w2945 & ~w2946;
assign w2948 = ~w2944 & w2947;
assign w2949 = ~b_28 & ~b_29;
assign w2950 = b_28 & b_29;
assign w2951 = ~w2949 & ~w2950;
assign w2952 = (w1931 & w38536) | (w1931 & w38537) | (w38536 & w38537);
assign w2953 = (~w1931 & w38538) | (~w1931 & w38539) | (w38538 & w38539);
assign w2954 = ~w2952 & ~w2953;
assign w2955 = (w2948 & ~w2954) | (w2948 & w28273) | (~w2954 & w28273);
assign w2956 = (w2954 & w38540) | (w2954 & w38541) | (w38540 & w38541);
assign w2957 = (~w2954 & w38542) | (~w2954 & w38543) | (w38542 & w38543);
assign w2958 = ~w2955 & ~w2956;
assign w2959 = ~w2957 & ~w2958;
assign w2960 = (~w2959 & w2942) | (~w2959 & w28274) | (w2942 & w28274);
assign w2961 = ~w2943 & ~w2960;
assign w2962 = ~w2942 & w38544;
assign w2963 = ~w2961 & ~w2962;
assign w2964 = (~w2778 & w2594) | (~w2778 & w38545) | (w2594 & w38545);
assign w2965 = ~w2963 & ~w2964;
assign w2966 = w2963 & w2964;
assign w2967 = ~w2965 & ~w2966;
assign w2968 = (~w2928 & w2931) | (~w2928 & w27407) | (w2931 & w27407);
assign w2969 = b_15 & w986;
assign w2970 = w1069 & w28275;
assign w2971 = b_14 & w981;
assign w2972 = ~w2970 & ~w2971;
assign w2973 = ~w2969 & w2972;
assign w2974 = (w2973 & ~w827) | (w2973 & w28276) | (~w827 & w28276);
assign w2975 = (w827 & w38546) | (w827 & w38547) | (w38546 & w38547);
assign w2976 = (~w827 & w38548) | (~w827 & w38549) | (w38548 & w38549);
assign w2977 = ~w2974 & ~w2975;
assign w2978 = ~w2976 & ~w2977;
assign w2979 = (~w2870 & w2805) | (~w2870 & w26778) | (w2805 & w26778);
assign w2980 = b_12 & w1295;
assign w2981 = w1422 & w28277;
assign w2982 = b_11 & w1290;
assign w2983 = ~w2981 & ~w2982;
assign w2984 = ~w2980 & w2983;
assign w2985 = (w2984 & ~w552) | (w2984 & w28278) | (~w552 & w28278);
assign w2986 = (w552 & w38550) | (w552 & w38551) | (w38550 & w38551);
assign w2987 = (~w552 & w38552) | (~w552 & w38553) | (w38552 & w38553);
assign w2988 = ~w2985 & ~w2986;
assign w2989 = ~w2987 & ~w2988;
assign w2990 = (~w2864 & ~w2865) | (~w2864 & w28279) | (~w2865 & w28279);
assign w2991 = b_6 & w2158;
assign w2992 = w2294 & w28280;
assign w2993 = b_5 & w2153;
assign w2994 = ~w2992 & ~w2993;
assign w2995 = ~w2991 & w2994;
assign w2996 = (w2995 & ~w190) | (w2995 & w28281) | (~w190 & w28281);
assign w2997 = (w190 & w38554) | (w190 & w38555) | (w38554 & w38555);
assign w2998 = (~w190 & w38556) | (~w190 & w38557) | (w38556 & w38557);
assign w2999 = ~w2996 & ~w2997;
assign w3000 = ~w2998 & ~w2999;
assign w3001 = a_29 & ~a_30;
assign w3002 = ~a_29 & a_30;
assign w3003 = ~w3001 & ~w3002;
assign w3004 = b_0 & ~w3003;
assign w3005 = (w3004 & w2830) | (w3004 & w25539) | (w2830 & w25539);
assign w3006 = ~w2830 & w25540;
assign w3007 = ~w3005 & ~w3006;
assign w3008 = b_3 & w2639;
assign w3009 = w2820 & w25778;
assign w3010 = b_2 & w2634;
assign w3011 = ~w3009 & ~w3010;
assign w3012 = ~w3008 & w3011;
assign w3013 = w57 & w2642;
assign w3014 = w3012 & ~w3013;
assign w3015 = a_29 & ~w3014;
assign w3016 = w3014 & a_29;
assign w3017 = ~w3014 & ~w3015;
assign w3018 = ~w3016 & ~w3017;
assign w3019 = ~w3007 & ~w3018;
assign w3020 = w3007 & w3018;
assign w3021 = ~w3019 & ~w3020;
assign w3022 = ~w3000 & w3021;
assign w3023 = w3021 & ~w3022;
assign w3024 = ~w3021 & ~w3000;
assign w3025 = ~w3023 & ~w3024;
assign w3026 = ~w2849 & w3025;
assign w3027 = w2849 & ~w3025;
assign w3028 = ~w3026 & ~w3027;
assign w3029 = b_9 & w1694;
assign w3030 = w1834 & w28282;
assign w3031 = b_8 & w1689;
assign w3032 = ~w3030 & ~w3031;
assign w3033 = ~w3029 & w3032;
assign w3034 = (w3033 & ~w371) | (w3033 & w28283) | (~w371 & w28283);
assign w3035 = (w371 & w38558) | (w371 & w38559) | (w38558 & w38559);
assign w3036 = (~w371 & w38560) | (~w371 & w38561) | (w38560 & w38561);
assign w3037 = ~w3034 & ~w3035;
assign w3038 = ~w3036 & ~w3037;
assign w3039 = ~w3028 & ~w3038;
assign w3040 = w3028 & w3038;
assign w3041 = ~w3039 & ~w3040;
assign w3042 = ~w2990 & w3041;
assign w3043 = w2990 & ~w3041;
assign w3044 = ~w3042 & ~w3043;
assign w3045 = w2989 & ~w3044;
assign w3046 = ~w2989 & w3044;
assign w3047 = ~w3045 & ~w3046;
assign w3048 = ~w2979 & w3047;
assign w3049 = w2979 & ~w3047;
assign w3050 = ~w3048 & ~w3049;
assign w3051 = ~w2978 & w3050;
assign w3052 = w3050 & ~w3051;
assign w3053 = ~w3050 & ~w2978;
assign w3054 = ~w3052 & ~w3053;
assign w3055 = (~w2875 & w2878) | (~w2875 & w28284) | (w2878 & w28284);
assign w3056 = w3054 & w3055;
assign w3057 = ~w3054 & ~w3055;
assign w3058 = ~w3056 & ~w3057;
assign w3059 = b_18 & w657;
assign w3060 = w754 & w28285;
assign w3061 = b_17 & w652;
assign w3062 = ~w3060 & ~w3061;
assign w3063 = ~w3059 & w3062;
assign w3064 = (w3063 & ~w1238) | (w3063 & w25010) | (~w1238 & w25010);
assign w3065 = (w1238 & w28286) | (w1238 & w28287) | (w28286 & w28287);
assign w3066 = (~w1238 & w28288) | (~w1238 & w28289) | (w28288 & w28289);
assign w3067 = ~w3064 & ~w3065;
assign w3068 = ~w3066 & ~w3067;
assign w3069 = w3058 & ~w3068;
assign w3070 = w3058 & ~w3069;
assign w3071 = ~w3058 & ~w3068;
assign w3072 = ~w3070 & ~w3071;
assign w3073 = (~w2893 & w2897) | (~w2893 & w26779) | (w2897 & w26779);
assign w3074 = w3072 & w3073;
assign w3075 = ~w3072 & ~w3073;
assign w3076 = ~w3074 & ~w3075;
assign w3077 = b_21 & w418;
assign w3078 = w481 & w28290;
assign w3079 = b_20 & w413;
assign w3080 = ~w3078 & ~w3079;
assign w3081 = ~w3077 & w3080;
assign w3082 = (w3081 & ~w1634) | (w3081 & w28291) | (~w1634 & w28291);
assign w3083 = (w1634 & w38562) | (w1634 & w38563) | (w38562 & w38563);
assign w3084 = (~w1634 & w38564) | (~w1634 & w38565) | (w38564 & w38565);
assign w3085 = ~w3082 & ~w3083;
assign w3086 = ~w3084 & ~w3085;
assign w3087 = w3076 & ~w3086;
assign w3088 = w3076 & ~w3087;
assign w3089 = ~w3076 & ~w3086;
assign w3090 = ~w3088 & ~w3089;
assign w3091 = ~w2915 & w3090;
assign w3092 = w2915 & ~w3090;
assign w3093 = ~w3091 & ~w3092;
assign w3094 = b_24 & w239;
assign w3095 = w266 & w28292;
assign w3096 = b_23 & w234;
assign w3097 = ~w3095 & ~w3096;
assign w3098 = ~w3094 & w3097;
assign w3099 = (w3098 & ~w2083) | (w3098 & w28293) | (~w2083 & w28293);
assign w3100 = (w2083 & w38566) | (w2083 & w38567) | (w38566 & w38567);
assign w3101 = (~w2083 & w38568) | (~w2083 & w38569) | (w38568 & w38569);
assign w3102 = ~w3099 & ~w3100;
assign w3103 = ~w3101 & ~w3102;
assign w3104 = ~w3093 & ~w3103;
assign w3105 = w3093 & w3103;
assign w3106 = ~w3104 & ~w3105;
assign w3107 = w2968 & ~w3106;
assign w3108 = ~w2968 & w3106;
assign w3109 = ~w3107 & ~w3108;
assign w3110 = b_27 & w99;
assign w3111 = w136 & w28294;
assign w3112 = b_26 & w94;
assign w3113 = ~w3111 & ~w3112;
assign w3114 = ~w3110 & w3113;
assign w3115 = (w3114 & ~w2582) | (w3114 & w28295) | (~w2582 & w28295);
assign w3116 = (w2582 & w38570) | (w2582 & w38571) | (w38570 & w38571);
assign w3117 = (~w2582 & w38572) | (~w2582 & w38573) | (w38572 & w38573);
assign w3118 = ~w3115 & ~w3116;
assign w3119 = ~w3117 & ~w3118;
assign w3120 = w3109 & ~w3119;
assign w3121 = w3109 & ~w3120;
assign w3122 = ~w3109 & ~w3119;
assign w3123 = ~w3121 & ~w3122;
assign w3124 = (~w2936 & w2939) | (~w2936 & w28296) | (w2939 & w28296);
assign w3125 = w3123 & w3124;
assign w3126 = ~w3123 & ~w3124;
assign w3127 = ~w3125 & ~w3126;
assign w3128 = w8 & w28297;
assign w3129 = ~w8 & w28298;
assign w3130 = b_29 & w4;
assign w3131 = ~w3129 & ~w3130;
assign w3132 = ~w3128 & w3131;
assign w3133 = ~b_29 & ~b_30;
assign w3134 = b_29 & b_30;
assign w3135 = ~w3133 & ~w3134;
assign w3136 = (w1931 & w38574) | (w1931 & w38575) | (w38574 & w38575);
assign w3137 = (~w1931 & w38576) | (~w1931 & w38577) | (w38576 & w38577);
assign w3138 = ~w3136 & ~w3137;
assign w3139 = (w3132 & ~w3138) | (w3132 & w28305) | (~w3138 & w28305);
assign w3140 = (w3138 & w38578) | (w3138 & w38579) | (w38578 & w38579);
assign w3141 = (~w3138 & w38580) | (~w3138 & w38581) | (w38580 & w38581);
assign w3142 = ~w3139 & ~w3140;
assign w3143 = ~w3141 & ~w3142;
assign w3144 = w3127 & ~w3143;
assign w3145 = w3127 & ~w3144;
assign w3146 = ~w3127 & ~w3143;
assign w3147 = ~w3145 & ~w3146;
assign w3148 = (~w2960 & w2963) | (~w2960 & w28306) | (w2963 & w28306);
assign w3149 = ~w3147 & ~w3148;
assign w3150 = w3147 & w3148;
assign w3151 = ~w3149 & ~w3150;
assign w3152 = b_16 & w986;
assign w3153 = w1069 & w28307;
assign w3154 = b_15 & w981;
assign w3155 = ~w3153 & ~w3154;
assign w3156 = ~w3152 & w3155;
assign w3157 = (w3156 & ~w926) | (w3156 & w28308) | (~w926 & w28308);
assign w3158 = (w926 & w38582) | (w926 & w38583) | (w38582 & w38583);
assign w3159 = (~w926 & w38584) | (~w926 & w38585) | (w38584 & w38585);
assign w3160 = ~w3157 & ~w3158;
assign w3161 = ~w3159 & ~w3160;
assign w3162 = (~w3022 & w3025) | (~w3022 & w26130) | (w3025 & w26130);
assign w3163 = b_7 & w2158;
assign w3164 = w2294 & w28309;
assign w3165 = b_6 & w2153;
assign w3166 = ~w3164 & ~w3165;
assign w3167 = ~w3163 & w3166;
assign w3168 = (w3167 & ~w213) | (w3167 & w28310) | (~w213 & w28310);
assign w3169 = (w213 & w38586) | (w213 & w38587) | (w38586 & w38587);
assign w3170 = (~w213 & w38588) | (~w213 & w38589) | (w38588 & w38589);
assign w3171 = ~w3168 & ~w3169;
assign w3172 = ~w3170 & ~w3171;
assign w3173 = ~w2830 & w28311;
assign w3174 = (~w3173 & w3007) | (~w3173 & w28312) | (w3007 & w28312);
assign w3175 = b_4 & w2639;
assign w3176 = w2820 & w25541;
assign w3177 = b_3 & w2634;
assign w3178 = ~w3176 & ~w3177;
assign w3179 = ~w3175 & w3178;
assign w3180 = w84 & w2642;
assign w3181 = w3179 & ~w3180;
assign w3182 = (a_29 & w3180) | (a_29 & w25542) | (w3180 & w25542);
assign w3183 = ~w3180 & w25779;
assign w3184 = ~w3181 & ~w3182;
assign w3185 = ~w3183 & ~w3184;
assign w3186 = (a_32 & w3003) | (a_32 & w28313) | (w3003 & w28313);
assign w3187 = ~a_30 & a_31;
assign w3188 = a_30 & ~a_31;
assign w3189 = ~w3187 & ~w3188;
assign w3190 = w3003 & ~w3189;
assign w3191 = b_0 & w3190;
assign w3192 = ~a_31 & a_32;
assign w3193 = a_31 & ~a_32;
assign w3194 = ~w3192 & ~w3193;
assign w3195 = ~w3003 & w3194;
assign w3196 = b_1 & w3195;
assign w3197 = ~w3191 & ~w3196;
assign w3198 = ~w3003 & ~w3194;
assign w3199 = ~w15 & w3198;
assign w3200 = w3197 & ~w3199;
assign w3201 = (a_32 & ~w3197) | (a_32 & w25543) | (~w3197 & w25543);
assign w3202 = w3197 & w25780;
assign w3203 = ~w3200 & ~w3201;
assign w3204 = (w3186 & w3203) | (w3186 & w25781) | (w3203 & w25781);
assign w3205 = ~w3203 & w25782;
assign w3206 = ~w3204 & ~w3205;
assign w3207 = w3185 & w3206;
assign w3208 = ~w3185 & ~w3206;
assign w3209 = ~w3207 & ~w3208;
assign w3210 = ~w3174 & ~w3209;
assign w3211 = w3174 & w3209;
assign w3212 = ~w3210 & ~w3211;
assign w3213 = ~w3172 & w3212;
assign w3214 = w3172 & ~w3212;
assign w3215 = ~w3213 & ~w3214;
assign w3216 = ~w3162 & w3215;
assign w3217 = w3162 & ~w3215;
assign w3218 = ~w3216 & ~w3217;
assign w3219 = b_10 & w1694;
assign w3220 = w1834 & w28314;
assign w3221 = b_9 & w1689;
assign w3222 = ~w3220 & ~w3221;
assign w3223 = ~w3219 & w3222;
assign w3224 = (w3223 & ~w454) | (w3223 & w25011) | (~w454 & w25011);
assign w3225 = (w454 & w28315) | (w454 & w28316) | (w28315 & w28316);
assign w3226 = (~w454 & w38590) | (~w454 & w38591) | (w38590 & w38591);
assign w3227 = ~w3224 & ~w3225;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = w3218 & ~w3228;
assign w3230 = w3218 & ~w3229;
assign w3231 = ~w3218 & ~w3228;
assign w3232 = ~w3230 & ~w3231;
assign w3233 = (~w3039 & w2990) | (~w3039 & w26131) | (w2990 & w26131);
assign w3234 = w3232 & w3233;
assign w3235 = ~w3232 & ~w3233;
assign w3236 = ~w3234 & ~w3235;
assign w3237 = b_13 & w1295;
assign w3238 = w1422 & w28317;
assign w3239 = b_12 & w1290;
assign w3240 = ~w3238 & ~w3239;
assign w3241 = ~w3237 & w3240;
assign w3242 = (w3241 & ~w711) | (w3241 & w28318) | (~w711 & w28318);
assign w3243 = (w711 & w38592) | (w711 & w38593) | (w38592 & w38593);
assign w3244 = (~w711 & w38594) | (~w711 & w38595) | (w38594 & w38595);
assign w3245 = ~w3242 & ~w3243;
assign w3246 = ~w3244 & ~w3245;
assign w3247 = ~w3236 & w3246;
assign w3248 = w3236 & ~w3246;
assign w3249 = ~w3247 & ~w3248;
assign w3250 = (~w3046 & w2979) | (~w3046 & w28319) | (w2979 & w28319);
assign w3251 = w3249 & ~w3250;
assign w3252 = ~w3249 & w3250;
assign w3253 = ~w3251 & ~w3252;
assign w3254 = ~w3161 & w3253;
assign w3255 = w3253 & ~w3254;
assign w3256 = ~w3253 & ~w3161;
assign w3257 = ~w3255 & ~w3256;
assign w3258 = (~w3051 & w3055) | (~w3051 & w26889) | (w3055 & w26889);
assign w3259 = w3257 & w3258;
assign w3260 = ~w3257 & ~w3258;
assign w3261 = ~w3259 & ~w3260;
assign w3262 = b_19 & w657;
assign w3263 = w754 & w28320;
assign w3264 = b_18 & w652;
assign w3265 = ~w3263 & ~w3264;
assign w3266 = ~w3262 & w3265;
assign w3267 = (w3266 & ~w1372) | (w3266 & w25012) | (~w1372 & w25012);
assign w3268 = (w1372 & w28321) | (w1372 & w28322) | (w28321 & w28322);
assign w3269 = (~w1372 & w28323) | (~w1372 & w28324) | (w28323 & w28324);
assign w3270 = ~w3267 & ~w3268;
assign w3271 = ~w3269 & ~w3270;
assign w3272 = w3261 & ~w3271;
assign w3273 = w3261 & ~w3272;
assign w3274 = ~w3261 & ~w3271;
assign w3275 = ~w3273 & ~w3274;
assign w3276 = (~w3069 & w3072) | (~w3069 & w27130) | (w3072 & w27130);
assign w3277 = w3275 & w3276;
assign w3278 = ~w3275 & ~w3276;
assign w3279 = ~w3277 & ~w3278;
assign w3280 = b_22 & w418;
assign w3281 = w481 & w28325;
assign w3282 = b_21 & w413;
assign w3283 = ~w3281 & ~w3282;
assign w3284 = ~w3280 & w3283;
assign w3285 = (w3284 & ~w1786) | (w3284 & w25013) | (~w1786 & w25013);
assign w3286 = (w1786 & w28326) | (w1786 & w28327) | (w28326 & w28327);
assign w3287 = (~w1786 & w28328) | (~w1786 & w28329) | (w28328 & w28329);
assign w3288 = ~w3285 & ~w3286;
assign w3289 = ~w3287 & ~w3288;
assign w3290 = w3279 & ~w3289;
assign w3291 = w3279 & ~w3290;
assign w3292 = ~w3279 & ~w3289;
assign w3293 = ~w3291 & ~w3292;
assign w3294 = ~w2915 & ~w3090;
assign w3295 = ~w3087 & ~w3294;
assign w3296 = w3293 & w3295;
assign w3297 = ~w3293 & ~w3295;
assign w3298 = ~w3296 & ~w3297;
assign w3299 = b_25 & w239;
assign w3300 = w266 & w28330;
assign w3301 = b_24 & w234;
assign w3302 = ~w3300 & ~w3301;
assign w3303 = ~w3299 & w3302;
assign w3304 = (w3303 & ~w2108) | (w3303 & w28331) | (~w2108 & w28331);
assign w3305 = (w2108 & w38596) | (w2108 & w38597) | (w38596 & w38597);
assign w3306 = (~w2108 & w38598) | (~w2108 & w38599) | (w38598 & w38599);
assign w3307 = ~w3304 & ~w3305;
assign w3308 = ~w3306 & ~w3307;
assign w3309 = w3298 & ~w3308;
assign w3310 = w3298 & ~w3309;
assign w3311 = ~w3298 & ~w3308;
assign w3312 = ~w3310 & ~w3311;
assign w3313 = (~w3104 & w2968) | (~w3104 & w28332) | (w2968 & w28332);
assign w3314 = w3312 & w3313;
assign w3315 = ~w3312 & ~w3313;
assign w3316 = ~w3314 & ~w3315;
assign w3317 = b_28 & w99;
assign w3318 = w136 & w28333;
assign w3319 = b_27 & w94;
assign w3320 = ~w3318 & ~w3319;
assign w3321 = ~w3317 & w3320;
assign w3322 = (w3321 & ~w2771) | (w3321 & w28334) | (~w2771 & w28334);
assign w3323 = (w2771 & w38600) | (w2771 & w38601) | (w38600 & w38601);
assign w3324 = (~w2771 & w38602) | (~w2771 & w38603) | (w38602 & w38603);
assign w3325 = ~w3322 & ~w3323;
assign w3326 = ~w3324 & ~w3325;
assign w3327 = w3316 & ~w3326;
assign w3328 = w3316 & ~w3327;
assign w3329 = ~w3316 & ~w3326;
assign w3330 = ~w3328 & ~w3329;
assign w3331 = (~w3120 & w3123) | (~w3120 & w38604) | (w3123 & w38604);
assign w3332 = w3330 & w3331;
assign w3333 = ~w3330 & ~w3331;
assign w3334 = ~w3332 & ~w3333;
assign w3335 = w8 & w28335;
assign w3336 = ~w8 & w28336;
assign w3337 = b_30 & w4;
assign w3338 = ~w3336 & ~w3337;
assign w3339 = ~w3335 & w3338;
assign w3340 = ~b_30 & ~b_31;
assign w3341 = b_30 & b_31;
assign w3342 = ~w3340 & ~w3341;
assign w3343 = (w1931 & w38605) | (w1931 & w38606) | (w38605 & w38606);
assign w3344 = (~w1931 & w38607) | (~w1931 & w38608) | (w38607 & w38608);
assign w3345 = ~w3343 & ~w3344;
assign w3346 = (w3339 & ~w3345) | (w3339 & w28342) | (~w3345 & w28342);
assign w3347 = (w3345 & w38609) | (w3345 & w38610) | (w38609 & w38610);
assign w3348 = (~w3345 & w38611) | (~w3345 & w38612) | (w38611 & w38612);
assign w3349 = ~w3346 & ~w3347;
assign w3350 = ~w3348 & ~w3349;
assign w3351 = w3334 & ~w3350;
assign w3352 = w3334 & ~w3351;
assign w3353 = ~w3334 & ~w3350;
assign w3354 = ~w3352 & ~w3353;
assign w3355 = (~w3144 & w3147) | (~w3144 & w38613) | (w3147 & w38613);
assign w3356 = ~w3354 & ~w3355;
assign w3357 = w3354 & w3355;
assign w3358 = ~w3356 & ~w3357;
assign w3359 = (~w3351 & w3354) | (~w3351 & w38614) | (w3354 & w38614);
assign w3360 = (~w3327 & w3330) | (~w3327 & w38615) | (w3330 & w38615);
assign w3361 = b_26 & w239;
assign w3362 = w266 & w28343;
assign w3363 = b_25 & w234;
assign w3364 = ~w3362 & ~w3363;
assign w3365 = ~w3361 & w3364;
assign w3366 = (w3365 & ~w2416) | (w3365 & w28344) | (~w2416 & w28344);
assign w3367 = (w2416 & w38616) | (w2416 & w38617) | (w38616 & w38617);
assign w3368 = (~w2416 & w38618) | (~w2416 & w38619) | (w38618 & w38619);
assign w3369 = ~w3366 & ~w3367;
assign w3370 = ~w3368 & ~w3369;
assign w3371 = (~w3290 & w3295) | (~w3290 & w25014) | (w3295 & w25014);
assign w3372 = (~w3272 & w3276) | (~w3272 & w27023) | (w3276 & w27023);
assign w3373 = b_17 & w986;
assign w3374 = w1069 & w28345;
assign w3375 = b_16 & w981;
assign w3376 = ~w3374 & ~w3375;
assign w3377 = ~w3373 & w3376;
assign w3378 = (w3377 & ~w1038) | (w3377 & w28346) | (~w1038 & w28346);
assign w3379 = (w1038 & w38620) | (w1038 & w38621) | (w38620 & w38621);
assign w3380 = (~w1038 & w38622) | (~w1038 & w38623) | (w38622 & w38623);
assign w3381 = ~w3378 & ~w3379;
assign w3382 = ~w3380 & ~w3381;
assign w3383 = (~w3248 & w3250) | (~w3248 & w26890) | (w3250 & w26890);
assign w3384 = ~w3229 & ~w3235;
assign w3385 = ~w3185 & w3206;
assign w3386 = (~w3385 & w3174) | (~w3385 & w25015) | (w3174 & w25015);
assign w3387 = b_2 & w3195;
assign w3388 = w3003 & ~w3194;
assign w3389 = w3388 & w25367;
assign w3390 = b_1 & w3190;
assign w3391 = ~w3389 & ~w3390;
assign w3392 = ~w3387 & w3391;
assign w3393 = w35 & w3198;
assign w3394 = w3392 & ~w3393;
assign w3395 = (a_32 & ~w3392) | (a_32 & w25544) | (~w3392 & w25544);
assign w3396 = w3392 & w25783;
assign w3397 = ~w3394 & ~w3395;
assign w3398 = ~w3396 & ~w3397;
assign w3399 = ~w3204 & w3398;
assign w3400 = w3204 & ~w3398;
assign w3401 = ~w3399 & ~w3400;
assign w3402 = b_5 & w2639;
assign w3403 = w2820 & w26539;
assign w3404 = b_4 & w2634;
assign w3405 = ~w3403 & ~w3404;
assign w3406 = ~w3402 & w3405;
assign w3407 = w129 & w2642;
assign w3408 = w3406 & ~w3407;
assign w3409 = (a_29 & w3407) | (a_29 & w26540) | (w3407 & w26540);
assign w3410 = ~w3407 & w38624;
assign w3411 = ~w3408 & ~w3409;
assign w3412 = ~w3410 & ~w3411;
assign w3413 = w3401 & ~w3412;
assign w3414 = ~w3401 & w3412;
assign w3415 = ~w3386 & w25784;
assign w3416 = ~w3386 & ~w3415;
assign w3417 = (~w3413 & w3386) | (~w3413 & w26132) | (w3386 & w26132);
assign w3418 = ~w3414 & w3417;
assign w3419 = ~w3416 & ~w3418;
assign w3420 = b_8 & w2158;
assign w3421 = w2294 & w28347;
assign w3422 = b_7 & w2153;
assign w3423 = ~w3421 & ~w3422;
assign w3424 = ~w3420 & w3423;
assign w3425 = ~w308 & w28348;
assign w3426 = (w3424 & ~w28348) | (w3424 & w38625) | (~w28348 & w38625);
assign w3427 = (w28348 & w38626) | (w28348 & w38627) | (w38626 & w38627);
assign w3428 = ~w3425 & w28350;
assign w3429 = ~w3426 & ~w3427;
assign w3430 = ~w3428 & ~w3429;
assign w3431 = ~w3419 & ~w3430;
assign w3432 = ~w3419 & ~w3431;
assign w3433 = w3419 & ~w3430;
assign w3434 = ~w3432 & ~w3433;
assign w3435 = (~w3213 & w3162) | (~w3213 & w28351) | (w3162 & w28351);
assign w3436 = ~w3432 & w28352;
assign w3437 = (~w3435 & w3432) | (~w3435 & w28353) | (w3432 & w28353);
assign w3438 = ~w3436 & ~w3437;
assign w3439 = b_11 & w1694;
assign w3440 = w1834 & w28354;
assign w3441 = b_10 & w1689;
assign w3442 = ~w3440 & ~w3441;
assign w3443 = ~w3439 & w3442;
assign w3444 = (w3443 & ~w530) | (w3443 & w28355) | (~w530 & w28355);
assign w3445 = (w530 & w38628) | (w530 & w38629) | (w38628 & w38629);
assign w3446 = (~w530 & w38630) | (~w530 & w38631) | (w38630 & w38631);
assign w3447 = ~w3444 & ~w3445;
assign w3448 = ~w3446 & ~w3447;
assign w3449 = w3438 & ~w3448;
assign w3450 = ~w3438 & w3448;
assign w3451 = ~w3384 & w25016;
assign w3452 = ~w3384 & ~w3451;
assign w3453 = (~w3449 & w3384) | (~w3449 & w28356) | (w3384 & w28356);
assign w3454 = w3384 & w25016;
assign w3455 = b_14 & w1295;
assign w3456 = w1422 & w28357;
assign w3457 = b_13 & w1290;
assign w3458 = ~w3456 & ~w3457;
assign w3459 = ~w3455 & w3458;
assign w3460 = (w3459 & ~w735) | (w3459 & w28358) | (~w735 & w28358);
assign w3461 = (w735 & w38632) | (w735 & w38633) | (w38632 & w38633);
assign w3462 = (~w735 & w38634) | (~w735 & w38635) | (w38634 & w38635);
assign w3463 = ~w3460 & ~w3461;
assign w3464 = ~w3462 & ~w3463;
assign w3465 = ~w3452 & w28359;
assign w3466 = (~w3464 & w3452) | (~w3464 & w28360) | (w3452 & w28360);
assign w3467 = ~w3465 & ~w3466;
assign w3468 = ~w3383 & w3467;
assign w3469 = w3383 & ~w3467;
assign w3470 = ~w3468 & ~w3469;
assign w3471 = ~w3382 & w3470;
assign w3472 = w3470 & ~w3471;
assign w3473 = ~w3470 & ~w3382;
assign w3474 = ~w3472 & ~w3473;
assign w3475 = ~w3254 & ~w3260;
assign w3476 = w3474 & w3475;
assign w3477 = ~w3474 & ~w3475;
assign w3478 = ~w3476 & ~w3477;
assign w3479 = b_20 & w657;
assign w3480 = w754 & w28361;
assign w3481 = b_19 & w652;
assign w3482 = ~w3480 & ~w3481;
assign w3483 = ~w3479 & w3482;
assign w3484 = (w3483 & ~w1503) | (w3483 & w28362) | (~w1503 & w28362);
assign w3485 = (w1503 & w38636) | (w1503 & w38637) | (w38636 & w38637);
assign w3486 = (~w1503 & w38638) | (~w1503 & w38639) | (w38638 & w38639);
assign w3487 = ~w3484 & ~w3485;
assign w3488 = ~w3486 & ~w3487;
assign w3489 = w3478 & ~w3488;
assign w3490 = ~w3478 & w3488;
assign w3491 = ~w3372 & w25017;
assign w3492 = ~w3372 & ~w3491;
assign w3493 = (~w3489 & w3372) | (~w3489 & w28363) | (w3372 & w28363);
assign w3494 = b_23 & w418;
assign w3495 = w481 & w28364;
assign w3496 = b_22 & w413;
assign w3497 = ~w3495 & ~w3496;
assign w3498 = ~w3494 & w3497;
assign w3499 = (w3498 & ~w1933) | (w3498 & w25018) | (~w1933 & w25018);
assign w3500 = (w1933 & w28365) | (w1933 & w28366) | (w28365 & w28366);
assign w3501 = (~w1933 & w28367) | (~w1933 & w28368) | (w28367 & w28368);
assign w3502 = ~w3499 & ~w3500;
assign w3503 = ~w3501 & ~w3502;
assign w3504 = ~w3492 & w27207;
assign w3505 = (~w3503 & w3492) | (~w3503 & w27208) | (w3492 & w27208);
assign w3506 = ~w3504 & ~w3505;
assign w3507 = (~w3295 & w38640) | (~w3295 & w38641) | (w38640 & w38641);
assign w3508 = (w3295 & w38642) | (w3295 & w38643) | (w38642 & w38643);
assign w3509 = ~w3507 & ~w3508;
assign w3510 = ~w3370 & w3509;
assign w3511 = w3509 & ~w3510;
assign w3512 = ~w3509 & ~w3370;
assign w3513 = ~w3511 & ~w3512;
assign w3514 = (~w3309 & w3312) | (~w3309 & w28369) | (w3312 & w28369);
assign w3515 = w3513 & w3514;
assign w3516 = ~w3513 & ~w3514;
assign w3517 = ~w3515 & ~w3516;
assign w3518 = b_29 & w99;
assign w3519 = w136 & w28370;
assign w3520 = b_28 & w94;
assign w3521 = ~w3519 & ~w3520;
assign w3522 = ~w3518 & w3521;
assign w3523 = (w3522 & ~w2954) | (w3522 & w28371) | (~w2954 & w28371);
assign w3524 = (w2954 & w38644) | (w2954 & w38645) | (w38644 & w38645);
assign w3525 = (~w2954 & w38646) | (~w2954 & w38647) | (w38646 & w38647);
assign w3526 = ~w3523 & ~w3524;
assign w3527 = ~w3525 & ~w3526;
assign w3528 = w3517 & ~w3527;
assign w3529 = ~w3517 & w3527;
assign w3530 = (w3333 & w28372) | (w3333 & w28373) | (w28372 & w28373);
assign w3531 = ~w3360 & ~w3530;
assign w3532 = ~w3528 & ~w3530;
assign w3533 = ~w3530 & w28372;
assign w3534 = ~w3531 & ~w3533;
assign w3535 = w8 & w28374;
assign w3536 = ~w8 & w28375;
assign w3537 = b_31 & w4;
assign w3538 = ~w3536 & ~w3537;
assign w3539 = ~w3535 & w3538;
assign w3540 = ~b_31 & ~b_32;
assign w3541 = b_31 & b_32;
assign w3542 = ~w3540 & ~w3541;
assign w3543 = (w1931 & w38648) | (w1931 & w38649) | (w38648 & w38649);
assign w3544 = (~w1931 & w38650) | (~w1931 & w38651) | (w38650 & w38651);
assign w3545 = ~w3543 & ~w3544;
assign w3546 = (w3539 & ~w3545) | (w3539 & w28381) | (~w3545 & w28381);
assign w3547 = (w3545 & w38652) | (w3545 & w38653) | (w38652 & w38653);
assign w3548 = (~w3545 & w38654) | (~w3545 & w38655) | (w38654 & w38655);
assign w3549 = ~w3546 & ~w3547;
assign w3550 = ~w3548 & ~w3549;
assign w3551 = ~w3534 & w3550;
assign w3552 = w3534 & ~w3550;
assign w3553 = ~w3551 & ~w3552;
assign w3554 = ~w3359 & ~w3553;
assign w3555 = w3359 & w3553;
assign w3556 = ~w3554 & ~w3555;
assign w3557 = ~w3534 & ~w3550;
assign w3558 = (~w3557 & w3359) | (~w3557 & w28382) | (w3359 & w28382);
assign w3559 = b_27 & w239;
assign w3560 = w266 & w28383;
assign w3561 = b_26 & w234;
assign w3562 = ~w3560 & ~w3561;
assign w3563 = ~w3559 & w3562;
assign w3564 = (w3563 & ~w2582) | (w3563 & w28384) | (~w2582 & w28384);
assign w3565 = (w2582 & w38656) | (w2582 & w38657) | (w38656 & w38657);
assign w3566 = (~w2582 & w38658) | (~w2582 & w38659) | (w38658 & w38659);
assign w3567 = ~w3564 & ~w3565;
assign w3568 = ~w3566 & ~w3567;
assign w3569 = (~w3505 & w3371) | (~w3505 & w25020) | (w3371 & w25020);
assign w3570 = ~w3471 & ~w3477;
assign w3571 = (~w3466 & ~w3467) | (~w3466 & w26891) | (~w3467 & w26891);
assign w3572 = b_15 & w1295;
assign w3573 = w1422 & w28385;
assign w3574 = b_14 & w1290;
assign w3575 = ~w3573 & ~w3574;
assign w3576 = ~w3572 & w3575;
assign w3577 = (w3576 & ~w827) | (w3576 & w28386) | (~w827 & w28386);
assign w3578 = (w827 & w38660) | (w827 & w38661) | (w38660 & w38661);
assign w3579 = (~w827 & w38662) | (~w827 & w38663) | (w38662 & w38663);
assign w3580 = ~w3577 & ~w3578;
assign w3581 = ~w3579 & ~w3580;
assign w3582 = (~w3431 & w3434) | (~w3431 & w25021) | (w3434 & w25021);
assign w3583 = b_6 & w2639;
assign w3584 = w2820 & w28387;
assign w3585 = b_5 & w2634;
assign w3586 = ~w3584 & ~w3585;
assign w3587 = ~w3583 & w3586;
assign w3588 = (w3587 & ~w190) | (w3587 & w28388) | (~w190 & w28388);
assign w3589 = (w190 & w38664) | (w190 & w38665) | (w38664 & w38665);
assign w3590 = (~w190 & w38666) | (~w190 & w38667) | (w38666 & w38667);
assign w3591 = ~w3588 & ~w3589;
assign w3592 = ~w3590 & ~w3591;
assign w3593 = a_32 & ~a_33;
assign w3594 = ~a_32 & a_33;
assign w3595 = ~w3593 & ~w3594;
assign w3596 = b_0 & ~w3595;
assign w3597 = (w3596 & w3398) | (w3596 & w25785) | (w3398 & w25785);
assign w3598 = ~w3398 & w25786;
assign w3599 = ~w3597 & ~w3598;
assign w3600 = b_3 & w3195;
assign w3601 = w3388 & w26133;
assign w3602 = b_2 & w3190;
assign w3603 = ~w3601 & ~w3602;
assign w3604 = ~w3600 & w3603;
assign w3605 = w57 & w3198;
assign w3606 = w3604 & ~w3605;
assign w3607 = a_32 & ~w3606;
assign w3608 = w3606 & a_32;
assign w3609 = ~w3606 & ~w3607;
assign w3610 = ~w3608 & ~w3609;
assign w3611 = ~w3599 & ~w3610;
assign w3612 = w3599 & w3610;
assign w3613 = ~w3611 & ~w3612;
assign w3614 = ~w3592 & w3613;
assign w3615 = w3613 & ~w3614;
assign w3616 = ~w3613 & ~w3592;
assign w3617 = ~w3615 & ~w3616;
assign w3618 = ~w3417 & w3617;
assign w3619 = w3417 & ~w3617;
assign w3620 = ~w3618 & ~w3619;
assign w3621 = b_9 & w2158;
assign w3622 = w2294 & w28389;
assign w3623 = b_8 & w2153;
assign w3624 = ~w3622 & ~w3623;
assign w3625 = ~w3621 & w3624;
assign w3626 = (w3625 & ~w371) | (w3625 & w28390) | (~w371 & w28390);
assign w3627 = (w371 & w38668) | (w371 & w38669) | (w38668 & w38669);
assign w3628 = (~w371 & w38670) | (~w371 & w38671) | (w38670 & w38671);
assign w3629 = ~w3626 & ~w3627;
assign w3630 = ~w3628 & ~w3629;
assign w3631 = ~w3620 & ~w3630;
assign w3632 = w3620 & w3630;
assign w3633 = ~w3631 & ~w3632;
assign w3634 = w3582 & ~w3633;
assign w3635 = ~w3582 & w3633;
assign w3636 = ~w3634 & ~w3635;
assign w3637 = b_12 & w1694;
assign w3638 = w1834 & w28391;
assign w3639 = b_11 & w1689;
assign w3640 = ~w3638 & ~w3639;
assign w3641 = ~w3637 & w3640;
assign w3642 = (w3641 & ~w552) | (w3641 & w25022) | (~w552 & w25022);
assign w3643 = (w552 & w28392) | (w552 & w28393) | (w28392 & w28393);
assign w3644 = (~w552 & w38672) | (~w552 & w38673) | (w38672 & w38673);
assign w3645 = ~w3642 & ~w3643;
assign w3646 = ~w3644 & ~w3645;
assign w3647 = ~w3636 & w3646;
assign w3648 = w3636 & ~w3646;
assign w3649 = ~w3647 & ~w3648;
assign w3650 = ~w3453 & w3649;
assign w3651 = w3453 & ~w3649;
assign w3652 = ~w3650 & ~w3651;
assign w3653 = ~w3581 & w3652;
assign w3654 = w3652 & ~w3653;
assign w3655 = ~w3652 & ~w3581;
assign w3656 = ~w3654 & ~w3655;
assign w3657 = ~w3571 & w3656;
assign w3658 = w3571 & ~w3656;
assign w3659 = ~w3657 & ~w3658;
assign w3660 = b_18 & w986;
assign w3661 = w1069 & w28394;
assign w3662 = b_17 & w981;
assign w3663 = ~w3661 & ~w3662;
assign w3664 = ~w3660 & w3663;
assign w3665 = (w3664 & ~w1238) | (w3664 & w28395) | (~w1238 & w28395);
assign w3666 = (w1238 & w38674) | (w1238 & w38675) | (w38674 & w38675);
assign w3667 = (~w1238 & w38676) | (~w1238 & w38677) | (w38676 & w38677);
assign w3668 = ~w3665 & ~w3666;
assign w3669 = ~w3667 & ~w3668;
assign w3670 = ~w3659 & ~w3669;
assign w3671 = w3659 & w3669;
assign w3672 = ~w3670 & ~w3671;
assign w3673 = w3570 & ~w3672;
assign w3674 = ~w3570 & w3672;
assign w3675 = ~w3673 & ~w3674;
assign w3676 = b_21 & w657;
assign w3677 = w754 & w28396;
assign w3678 = b_20 & w652;
assign w3679 = ~w3677 & ~w3678;
assign w3680 = ~w3676 & w3679;
assign w3681 = (w3680 & ~w1634) | (w3680 & w28397) | (~w1634 & w28397);
assign w3682 = (w1634 & w38678) | (w1634 & w38679) | (w38678 & w38679);
assign w3683 = (~w1634 & w38680) | (~w1634 & w38681) | (w38680 & w38681);
assign w3684 = ~w3681 & ~w3682;
assign w3685 = ~w3683 & ~w3684;
assign w3686 = w3675 & ~w3685;
assign w3687 = w3675 & ~w3686;
assign w3688 = ~w3675 & ~w3685;
assign w3689 = ~w3687 & ~w3688;
assign w3690 = ~w3493 & w3689;
assign w3691 = w3493 & ~w3689;
assign w3692 = ~w3690 & ~w3691;
assign w3693 = b_24 & w418;
assign w3694 = w481 & w28398;
assign w3695 = b_23 & w413;
assign w3696 = ~w3694 & ~w3695;
assign w3697 = ~w3693 & w3696;
assign w3698 = (w3697 & ~w2083) | (w3697 & w25023) | (~w2083 & w25023);
assign w3699 = (w2083 & w28399) | (w2083 & w28400) | (w28399 & w28400);
assign w3700 = (~w2083 & w28401) | (~w2083 & w28402) | (w28401 & w28402);
assign w3701 = ~w3698 & ~w3699;
assign w3702 = ~w3700 & ~w3701;
assign w3703 = w3692 & w3702;
assign w3704 = ~w3692 & ~w3702;
assign w3705 = ~w3703 & ~w3704;
assign w3706 = ~w3569 & w3705;
assign w3707 = w3569 & ~w3705;
assign w3708 = ~w3706 & ~w3707;
assign w3709 = ~w3568 & w3708;
assign w3710 = w3708 & ~w3709;
assign w3711 = ~w3708 & ~w3568;
assign w3712 = ~w3710 & ~w3711;
assign w3713 = (~w3510 & w3514) | (~w3510 & w27408) | (w3514 & w27408);
assign w3714 = w3712 & w3713;
assign w3715 = ~w3712 & ~w3713;
assign w3716 = ~w3714 & ~w3715;
assign w3717 = b_30 & w99;
assign w3718 = w136 & w28403;
assign w3719 = b_29 & w94;
assign w3720 = ~w3718 & ~w3719;
assign w3721 = ~w3717 & w3720;
assign w3722 = (w3721 & ~w3138) | (w3721 & w28404) | (~w3138 & w28404);
assign w3723 = (w3138 & w38682) | (w3138 & w38683) | (w38682 & w38683);
assign w3724 = (~w3138 & w38684) | (~w3138 & w38685) | (w38684 & w38685);
assign w3725 = ~w3722 & ~w3723;
assign w3726 = ~w3724 & ~w3725;
assign w3727 = w3716 & ~w3726;
assign w3728 = w3716 & ~w3727;
assign w3729 = ~w3716 & ~w3726;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = ~w3532 & w3730;
assign w3732 = w3532 & ~w3730;
assign w3733 = ~w3731 & ~w3732;
assign w3734 = w8 & w28405;
assign w3735 = ~w8 & w28406;
assign w3736 = b_32 & w4;
assign w3737 = ~w3735 & ~w3736;
assign w3738 = ~w3734 & w3737;
assign w3739 = ~b_32 & ~b_33;
assign w3740 = b_32 & b_33;
assign w3741 = ~w3739 & ~w3740;
assign w3742 = (w1931 & w38688) | (w1931 & w38689) | (w38688 & w38689);
assign w3743 = (~w1931 & w38690) | (~w1931 & w38691) | (w38690 & w38691);
assign w3744 = ~w3742 & ~w3743;
assign w3745 = (w3738 & ~w3744) | (w3738 & w28409) | (~w3744 & w28409);
assign w3746 = (w3744 & w38692) | (w3744 & w38693) | (w38692 & w38693);
assign w3747 = (~w3744 & w38694) | (~w3744 & w38695) | (w38694 & w38695);
assign w3748 = ~w3745 & ~w3746;
assign w3749 = ~w3747 & ~w3748;
assign w3750 = ~w3733 & ~w3749;
assign w3751 = w3733 & w3749;
assign w3752 = ~w3750 & ~w3751;
assign w3753 = ~w3558 & w3752;
assign w3754 = w3558 & ~w3752;
assign w3755 = ~w3753 & ~w3754;
assign w3756 = (~w3750 & w3558) | (~w3750 & w28410) | (w3558 & w28410);
assign w3757 = (~w3727 & w3532) | (~w3727 & w38696) | (w3532 & w38696);
assign w3758 = ~w3704 & ~w3706;
assign w3759 = (~w3648 & w3453) | (~w3648 & w25024) | (w3453 & w25024);
assign w3760 = b_10 & w2158;
assign w3761 = w2294 & w28411;
assign w3762 = b_9 & w2153;
assign w3763 = ~w3761 & ~w3762;
assign w3764 = ~w3760 & w3763;
assign w3765 = (w3764 & ~w454) | (w3764 & w28412) | (~w454 & w28412);
assign w3766 = (w454 & w38697) | (w454 & w38698) | (w38697 & w38698);
assign w3767 = (~w454 & w38699) | (~w454 & w38700) | (w38699 & w38700);
assign w3768 = ~w3765 & ~w3766;
assign w3769 = ~w3767 & ~w3768;
assign w3770 = (~w3614 & w3617) | (~w3614 & w26780) | (w3617 & w26780);
assign w3771 = b_7 & w2639;
assign w3772 = w2820 & w28413;
assign w3773 = b_6 & w2634;
assign w3774 = ~w3772 & ~w3773;
assign w3775 = ~w3771 & w3774;
assign w3776 = (w3775 & ~w213) | (w3775 & w28414) | (~w213 & w28414);
assign w3777 = (w213 & w38701) | (w213 & w38702) | (w38701 & w38702);
assign w3778 = (~w213 & w38703) | (~w213 & w38704) | (w38703 & w38704);
assign w3779 = ~w3776 & ~w3777;
assign w3780 = ~w3778 & ~w3779;
assign w3781 = ~w3398 & w28415;
assign w3782 = (~w3781 & w3599) | (~w3781 & w28416) | (w3599 & w28416);
assign w3783 = b_4 & w3195;
assign w3784 = w3388 & w26134;
assign w3785 = b_3 & w3190;
assign w3786 = ~w3784 & ~w3785;
assign w3787 = ~w3783 & w3786;
assign w3788 = w84 & w3198;
assign w3789 = w3787 & ~w3788;
assign w3790 = (a_32 & w3788) | (a_32 & w26135) | (w3788 & w26135);
assign w3791 = ~w3788 & w26541;
assign w3792 = ~w3789 & ~w3790;
assign w3793 = ~w3791 & ~w3792;
assign w3794 = (a_35 & w3595) | (a_35 & w28417) | (w3595 & w28417);
assign w3795 = ~a_33 & a_34;
assign w3796 = a_33 & ~a_34;
assign w3797 = ~w3795 & ~w3796;
assign w3798 = w3595 & ~w3797;
assign w3799 = b_0 & w3798;
assign w3800 = ~a_34 & a_35;
assign w3801 = a_34 & ~a_35;
assign w3802 = ~w3800 & ~w3801;
assign w3803 = ~w3595 & w3802;
assign w3804 = b_1 & w3803;
assign w3805 = ~w3799 & ~w3804;
assign w3806 = ~w3595 & ~w3802;
assign w3807 = ~w15 & w3806;
assign w3808 = w3805 & ~w3807;
assign w3809 = (a_35 & ~w3805) | (a_35 & w25545) | (~w3805 & w25545);
assign w3810 = w3805 & w25787;
assign w3811 = ~w3808 & ~w3809;
assign w3812 = (w3794 & w3811) | (w3794 & w25788) | (w3811 & w25788);
assign w3813 = ~w3811 & w26542;
assign w3814 = ~w3812 & ~w3813;
assign w3815 = w3793 & ~w3814;
assign w3816 = ~w3793 & w3814;
assign w3817 = ~w3815 & ~w3816;
assign w3818 = ~w3782 & w3817;
assign w3819 = w3782 & ~w3817;
assign w3820 = ~w3818 & ~w3819;
assign w3821 = w3780 & ~w3820;
assign w3822 = ~w3780 & w3820;
assign w3823 = ~w3821 & ~w3822;
assign w3824 = ~w3770 & w3823;
assign w3825 = w3770 & ~w3823;
assign w3826 = ~w3824 & ~w3825;
assign w3827 = ~w3769 & w3826;
assign w3828 = w3826 & ~w3827;
assign w3829 = ~w3826 & ~w3769;
assign w3830 = ~w3828 & ~w3829;
assign w3831 = (~w3631 & w3582) | (~w3631 & w26781) | (w3582 & w26781);
assign w3832 = w3830 & w3831;
assign w3833 = ~w3830 & ~w3831;
assign w3834 = ~w3832 & ~w3833;
assign w3835 = b_13 & w1694;
assign w3836 = w1834 & w28418;
assign w3837 = b_12 & w1689;
assign w3838 = ~w3836 & ~w3837;
assign w3839 = ~w3835 & w3838;
assign w3840 = (w3839 & ~w711) | (w3839 & w28419) | (~w711 & w28419);
assign w3841 = (w711 & w38705) | (w711 & w38706) | (w38705 & w38706);
assign w3842 = (~w711 & w38707) | (~w711 & w38708) | (w38707 & w38708);
assign w3843 = ~w3840 & ~w3841;
assign w3844 = ~w3842 & ~w3843;
assign w3845 = w3834 & ~w3844;
assign w3846 = ~w3834 & w3844;
assign w3847 = ~w3759 & w26543;
assign w3848 = ~w3759 & ~w3847;
assign w3849 = (~w3845 & w3759) | (~w3845 & w26782) | (w3759 & w26782);
assign w3850 = ~w3846 & w3849;
assign w3851 = ~w3848 & ~w3850;
assign w3852 = b_16 & w1295;
assign w3853 = w1422 & w28420;
assign w3854 = b_15 & w1290;
assign w3855 = ~w3853 & ~w3854;
assign w3856 = ~w3852 & w3855;
assign w3857 = (w3856 & ~w926) | (w3856 & w28421) | (~w926 & w28421);
assign w3858 = (w926 & w38709) | (w926 & w38710) | (w38709 & w38710);
assign w3859 = (~w926 & w38711) | (~w926 & w38712) | (w38711 & w38712);
assign w3860 = ~w3857 & ~w3858;
assign w3861 = ~w3859 & ~w3860;
assign w3862 = ~w3851 & ~w3861;
assign w3863 = ~w3851 & ~w3862;
assign w3864 = w3851 & ~w3861;
assign w3865 = ~w3863 & ~w3864;
assign w3866 = (~w3653 & w3656) | (~w3653 & w26892) | (w3656 & w26892);
assign w3867 = ~w3863 & w38713;
assign w3868 = (~w3866 & w3863) | (~w3866 & w38714) | (w3863 & w38714);
assign w3869 = ~w3867 & ~w3868;
assign w3870 = b_19 & w986;
assign w3871 = w1069 & w28422;
assign w3872 = b_18 & w981;
assign w3873 = ~w3871 & ~w3872;
assign w3874 = ~w3870 & w3873;
assign w3875 = (w3874 & ~w1372) | (w3874 & w25025) | (~w1372 & w25025);
assign w3876 = (w1372 & w28423) | (w1372 & w28424) | (w28423 & w28424);
assign w3877 = (~w1372 & w28425) | (~w1372 & w28426) | (w28425 & w28426);
assign w3878 = ~w3875 & ~w3876;
assign w3879 = ~w3877 & ~w3878;
assign w3880 = w3869 & ~w3879;
assign w3881 = w3869 & ~w3880;
assign w3882 = ~w3869 & ~w3879;
assign w3883 = ~w3881 & ~w3882;
assign w3884 = (~w3670 & w3570) | (~w3670 & w25026) | (w3570 & w25026);
assign w3885 = ~w3881 & w28427;
assign w3886 = (~w3884 & w3881) | (~w3884 & w28428) | (w3881 & w28428);
assign w3887 = ~w3885 & ~w3886;
assign w3888 = b_22 & w657;
assign w3889 = w754 & w28429;
assign w3890 = b_21 & w652;
assign w3891 = ~w3889 & ~w3890;
assign w3892 = ~w3888 & w3891;
assign w3893 = (w3892 & ~w1786) | (w3892 & w25027) | (~w1786 & w25027);
assign w3894 = (w1786 & w28430) | (w1786 & w28431) | (w28430 & w28431);
assign w3895 = (~w1786 & w28432) | (~w1786 & w28433) | (w28432 & w28433);
assign w3896 = ~w3893 & ~w3894;
assign w3897 = ~w3895 & ~w3896;
assign w3898 = w3887 & ~w3897;
assign w3899 = w3887 & ~w3898;
assign w3900 = ~w3887 & ~w3897;
assign w3901 = ~w3899 & ~w3900;
assign w3902 = (~w3686 & w3689) | (~w3686 & w25028) | (w3689 & w25028);
assign w3903 = w3901 & w3902;
assign w3904 = ~w3901 & ~w3902;
assign w3905 = ~w3903 & ~w3904;
assign w3906 = b_25 & w418;
assign w3907 = w481 & w28434;
assign w3908 = b_24 & w413;
assign w3909 = ~w3907 & ~w3908;
assign w3910 = ~w3906 & w3909;
assign w3911 = (w3910 & ~w2108) | (w3910 & w25029) | (~w2108 & w25029);
assign w3912 = (w2108 & w28435) | (w2108 & w28436) | (w28435 & w28436);
assign w3913 = (~w2108 & w28437) | (~w2108 & w28438) | (w28437 & w28438);
assign w3914 = ~w3911 & ~w3912;
assign w3915 = ~w3913 & ~w3914;
assign w3916 = w3905 & ~w3915;
assign w3917 = ~w3905 & w3915;
assign w3918 = ~w3758 & w25030;
assign w3919 = ~w3758 & ~w3918;
assign w3920 = ~w3916 & ~w3918;
assign w3921 = ~w3918 & w25030;
assign w3922 = ~w3919 & ~w3921;
assign w3923 = b_28 & w239;
assign w3924 = w266 & w28439;
assign w3925 = b_27 & w234;
assign w3926 = ~w3924 & ~w3925;
assign w3927 = ~w3923 & w3926;
assign w3928 = (w3927 & ~w2771) | (w3927 & w25031) | (~w2771 & w25031);
assign w3929 = (w2771 & w28440) | (w2771 & w28441) | (w28440 & w28441);
assign w3930 = (~w2771 & w28442) | (~w2771 & w28443) | (w28442 & w28443);
assign w3931 = ~w3928 & ~w3929;
assign w3932 = ~w3930 & ~w3931;
assign w3933 = ~w3922 & ~w3932;
assign w3934 = ~w3922 & ~w3933;
assign w3935 = w3922 & ~w3932;
assign w3936 = (~w3709 & w3713) | (~w3709 & w28444) | (w3713 & w28444);
assign w3937 = ~w3934 & w38715;
assign w3938 = (~w3936 & w3934) | (~w3936 & w38716) | (w3934 & w38716);
assign w3939 = ~w3937 & ~w3938;
assign w3940 = b_31 & w99;
assign w3941 = w136 & w28445;
assign w3942 = b_30 & w94;
assign w3943 = ~w3941 & ~w3942;
assign w3944 = ~w3940 & w3943;
assign w3945 = (w3944 & ~w3345) | (w3944 & w28446) | (~w3345 & w28446);
assign w3946 = (w3345 & w38717) | (w3345 & w38718) | (w38717 & w38718);
assign w3947 = (~w3345 & w38719) | (~w3345 & w38720) | (w38719 & w38720);
assign w3948 = ~w3945 & ~w3946;
assign w3949 = ~w3947 & ~w3948;
assign w3950 = w3939 & ~w3949;
assign w3951 = ~w3939 & w3949;
assign w3952 = (~w3532 & w38721) | (~w3532 & w38722) | (w38721 & w38722);
assign w3953 = ~w3950 & w3952;
assign w3954 = ~w3757 & ~w3953;
assign w3955 = ~w3952 & ~w3950;
assign w3956 = w28447 & ~w3952;
assign w3957 = w8 & w28448;
assign w3958 = ~w8 & w28449;
assign w3959 = b_33 & w4;
assign w3960 = ~w3958 & ~w3959;
assign w3961 = ~w3957 & w3960;
assign w3962 = ~b_33 & ~b_34;
assign w3963 = b_33 & b_34;
assign w3964 = ~w3962 & ~w3963;
assign w3965 = (w1931 & w38723) | (w1931 & w38724) | (w38723 & w38724);
assign w3966 = (~w1931 & w38725) | (~w1931 & w38726) | (w38725 & w38726);
assign w3967 = ~w3965 & ~w3966;
assign w3968 = (w3961 & ~w3967) | (w3961 & w28454) | (~w3967 & w28454);
assign w3969 = (w3967 & w38727) | (w3967 & w38728) | (w38727 & w38728);
assign w3970 = (~w3967 & w38729) | (~w3967 & w38730) | (w38729 & w38730);
assign w3971 = ~w3968 & ~w3969;
assign w3972 = ~w3970 & ~w3971;
assign w3973 = (w3972 & w3954) | (w3972 & w28455) | (w3954 & w28455);
assign w3974 = ~w3954 & w28456;
assign w3975 = ~w3973 & ~w3974;
assign w3976 = ~w3756 & ~w3975;
assign w3977 = w3756 & w3975;
assign w3978 = ~w3976 & ~w3977;
assign w3979 = (~w3972 & w3954) | (~w3972 & w28457) | (w3954 & w28457);
assign w3980 = (~w3979 & w3756) | (~w3979 & w38731) | (w3756 & w38731);
assign w3981 = b_29 & w239;
assign w3982 = w266 & w28458;
assign w3983 = b_28 & w234;
assign w3984 = ~w3982 & ~w3983;
assign w3985 = ~w3981 & w3984;
assign w3986 = (w3985 & ~w2954) | (w3985 & w25034) | (~w2954 & w25034);
assign w3987 = (w2954 & w28459) | (w2954 & w28460) | (w28459 & w28460);
assign w3988 = (~w2954 & w28461) | (~w2954 & w28462) | (w28461 & w28462);
assign w3989 = ~w3986 & ~w3987;
assign w3990 = ~w3988 & ~w3989;
assign w3991 = b_26 & w418;
assign w3992 = w481 & w28463;
assign w3993 = b_25 & w413;
assign w3994 = ~w3992 & ~w3993;
assign w3995 = ~w3991 & w3994;
assign w3996 = (w3995 & ~w2416) | (w3995 & w28464) | (~w2416 & w28464);
assign w3997 = (w2416 & w38732) | (w2416 & w38733) | (w38732 & w38733);
assign w3998 = (~w2416 & w38734) | (~w2416 & w38735) | (w38734 & w38735);
assign w3999 = ~w3996 & ~w3997;
assign w4000 = ~w3998 & ~w3999;
assign w4001 = (~w3898 & w3901) | (~w3898 & w27024) | (w3901 & w27024);
assign w4002 = (~w3880 & w3883) | (~w3880 & w26893) | (w3883 & w26893);
assign w4003 = b_17 & w1295;
assign w4004 = w1422 & w28465;
assign w4005 = b_16 & w1290;
assign w4006 = ~w4004 & ~w4005;
assign w4007 = ~w4003 & w4006;
assign w4008 = (w4007 & ~w1038) | (w4007 & w28466) | (~w1038 & w28466);
assign w4009 = (w1038 & w38736) | (w1038 & w38737) | (w38736 & w38737);
assign w4010 = (~w1038 & w38738) | (~w1038 & w38739) | (w38738 & w38739);
assign w4011 = ~w4008 & ~w4009;
assign w4012 = ~w4010 & ~w4011;
assign w4013 = ~w3827 & ~w3833;
assign w4014 = b_11 & w2158;
assign w4015 = w2294 & w28467;
assign w4016 = b_10 & w2153;
assign w4017 = ~w4015 & ~w4016;
assign w4018 = ~w4014 & w4017;
assign w4019 = (w4018 & ~w530) | (w4018 & w28468) | (~w530 & w28468);
assign w4020 = (w530 & w38740) | (w530 & w38741) | (w38740 & w38741);
assign w4021 = (~w530 & w38742) | (~w530 & w38743) | (w38742 & w38743);
assign w4022 = ~w4019 & ~w4020;
assign w4023 = ~w4021 & ~w4022;
assign w4024 = (~w3822 & w3770) | (~w3822 & w28469) | (w3770 & w28469);
assign w4025 = (~w3816 & w3782) | (~w3816 & w26136) | (w3782 & w26136);
assign w4026 = b_2 & w3803;
assign w4027 = w3595 & ~w3802;
assign w4028 = w4027 & w25368;
assign w4029 = b_1 & w3798;
assign w4030 = ~w4028 & ~w4029;
assign w4031 = ~w4026 & w4030;
assign w4032 = w35 & w3806;
assign w4033 = w4031 & ~w4032;
assign w4034 = (a_35 & ~w4031) | (a_35 & w25546) | (~w4031 & w25546);
assign w4035 = w4031 & w25789;
assign w4036 = ~w4033 & ~w4034;
assign w4037 = ~w4035 & ~w4036;
assign w4038 = ~w3812 & w4037;
assign w4039 = w3812 & ~w4037;
assign w4040 = ~w4038 & ~w4039;
assign w4041 = b_5 & w3195;
assign w4042 = w3388 & w26894;
assign w4043 = b_4 & w3190;
assign w4044 = ~w4042 & ~w4043;
assign w4045 = ~w4041 & w4044;
assign w4046 = w129 & w3198;
assign w4047 = w4045 & ~w4046;
assign w4048 = (a_32 & w4046) | (a_32 & w26895) | (w4046 & w26895);
assign w4049 = ~w4046 & w38744;
assign w4050 = ~w4047 & ~w4048;
assign w4051 = ~w4049 & ~w4050;
assign w4052 = w4040 & ~w4051;
assign w4053 = ~w4040 & w4051;
assign w4054 = ~w4025 & w26544;
assign w4055 = ~w4025 & ~w4054;
assign w4056 = (~w4052 & w4025) | (~w4052 & w26783) | (w4025 & w26783);
assign w4057 = ~w4053 & w4056;
assign w4058 = ~w4055 & ~w4057;
assign w4059 = b_8 & w2639;
assign w4060 = w2820 & w28470;
assign w4061 = b_7 & w2634;
assign w4062 = ~w4060 & ~w4061;
assign w4063 = ~w4059 & w4062;
assign w4064 = ~w308 & w28471;
assign w4065 = (w4063 & ~w28471) | (w4063 & w38745) | (~w28471 & w38745);
assign w4066 = (w28471 & w38746) | (w28471 & w38747) | (w38746 & w38747);
assign w4067 = ~w4064 & w28473;
assign w4068 = ~w4065 & ~w4066;
assign w4069 = ~w4067 & ~w4068;
assign w4070 = ~w4058 & ~w4069;
assign w4071 = ~w4058 & ~w4070;
assign w4072 = w4058 & ~w4069;
assign w4073 = ~w4071 & ~w4072;
assign w4074 = (~w4024 & w4071) | (~w4024 & w28474) | (w4071 & w28474);
assign w4075 = ~w4071 & w28475;
assign w4076 = ~w4074 & ~w4075;
assign w4077 = ~w4023 & w4076;
assign w4078 = ~w4076 & ~w4023;
assign w4079 = w4076 & ~w4077;
assign w4080 = ~w4078 & ~w4079;
assign w4081 = ~w4013 & ~w4080;
assign w4082 = ~w4080 & ~w4081;
assign w4083 = b_14 & w1694;
assign w4084 = w1834 & w28476;
assign w4085 = b_13 & w1689;
assign w4086 = ~w4084 & ~w4085;
assign w4087 = ~w4083 & w4086;
assign w4088 = (w4087 & ~w735) | (w4087 & w28477) | (~w735 & w28477);
assign w4089 = (w735 & w38748) | (w735 & w38749) | (w38748 & w38749);
assign w4090 = (~w735 & w38750) | (~w735 & w38751) | (w38750 & w38751);
assign w4091 = ~w4088 & ~w4089;
assign w4092 = ~w4090 & ~w4091;
assign w4093 = ~w4082 & w26896;
assign w4094 = (~w4092 & w4082) | (~w4092 & w26897) | (w4082 & w26897);
assign w4095 = ~w4093 & ~w4094;
assign w4096 = ~w3849 & w4095;
assign w4097 = w3849 & ~w4095;
assign w4098 = ~w4096 & ~w4097;
assign w4099 = ~w4012 & w4098;
assign w4100 = w4098 & ~w4099;
assign w4101 = ~w4098 & ~w4012;
assign w4102 = ~w4100 & ~w4101;
assign w4103 = (~w3862 & w3865) | (~w3862 & w26898) | (w3865 & w26898);
assign w4104 = w4102 & w4103;
assign w4105 = ~w4102 & ~w4103;
assign w4106 = ~w4104 & ~w4105;
assign w4107 = b_20 & w986;
assign w4108 = w1069 & w28478;
assign w4109 = b_19 & w981;
assign w4110 = ~w4108 & ~w4109;
assign w4111 = ~w4107 & w4110;
assign w4112 = (w4111 & ~w1503) | (w4111 & w28479) | (~w1503 & w28479);
assign w4113 = (w1503 & w38752) | (w1503 & w38753) | (w38752 & w38753);
assign w4114 = (~w1503 & w38754) | (~w1503 & w38755) | (w38754 & w38755);
assign w4115 = ~w4112 & ~w4113;
assign w4116 = ~w4114 & ~w4115;
assign w4117 = w4106 & ~w4116;
assign w4118 = ~w4106 & w4116;
assign w4119 = ~w4002 & w25035;
assign w4120 = ~w4002 & ~w4119;
assign w4121 = (~w4117 & w4002) | (~w4117 & w27025) | (w4002 & w27025);
assign w4122 = (w27025 & w25035) | (w27025 & w38756) | (w25035 & w38756);
assign w4123 = ~w4120 & ~w4122;
assign w4124 = b_23 & w657;
assign w4125 = w754 & w28480;
assign w4126 = b_22 & w652;
assign w4127 = ~w4125 & ~w4126;
assign w4128 = ~w4124 & w4127;
assign w4129 = (w4128 & ~w1933) | (w4128 & w28481) | (~w1933 & w28481);
assign w4130 = (w1933 & w38757) | (w1933 & w38758) | (w38757 & w38758);
assign w4131 = (~w1933 & w38759) | (~w1933 & w38760) | (w38759 & w38760);
assign w4132 = ~w4129 & ~w4130;
assign w4133 = ~w4131 & ~w4132;
assign w4134 = w4123 & w4133;
assign w4135 = ~w4123 & ~w4133;
assign w4136 = ~w4134 & ~w4135;
assign w4137 = ~w4001 & w4136;
assign w4138 = w4001 & ~w4136;
assign w4139 = ~w4137 & ~w4138;
assign w4140 = w4000 & ~w4139;
assign w4141 = ~w4000 & w4139;
assign w4142 = ~w4140 & ~w4141;
assign w4143 = ~w3920 & w4142;
assign w4144 = w3920 & ~w4142;
assign w4145 = ~w4143 & ~w4144;
assign w4146 = ~w3990 & w4145;
assign w4147 = w4145 & ~w4146;
assign w4148 = ~w4145 & ~w3990;
assign w4149 = ~w4147 & ~w4148;
assign w4150 = (~w3933 & w3936) | (~w3933 & w25036) | (w3936 & w25036);
assign w4151 = w4149 & w4150;
assign w4152 = ~w4149 & ~w4150;
assign w4153 = ~w4151 & ~w4152;
assign w4154 = b_32 & w99;
assign w4155 = w136 & w28482;
assign w4156 = b_31 & w94;
assign w4157 = ~w4155 & ~w4156;
assign w4158 = ~w4154 & w4157;
assign w4159 = (w4158 & ~w3545) | (w4158 & w28483) | (~w3545 & w28483);
assign w4160 = (w3545 & w38761) | (w3545 & w38762) | (w38761 & w38762);
assign w4161 = (~w3545 & w38763) | (~w3545 & w38764) | (w38763 & w38764);
assign w4162 = ~w4159 & ~w4160;
assign w4163 = ~w4161 & ~w4162;
assign w4164 = w4153 & ~w4163;
assign w4165 = ~w4153 & w4163;
assign w4166 = (w3952 & w28484) | (w3952 & ~w4165) | (w28484 & ~w4165);
assign w4167 = (w28484 & w28485) | (w28484 & w38765) | (w28485 & w38765);
assign w4168 = ~w3955 & ~w4167;
assign w4169 = (~w28484 & w38766) | (~w28484 & w38767) | (w38766 & w38767);
assign w4170 = w28485 & ~w4166;
assign w4171 = w8 & w28486;
assign w4172 = ~w8 & w28487;
assign w4173 = b_34 & w4;
assign w4174 = ~w4172 & ~w4173;
assign w4175 = ~w4171 & w4174;
assign w4176 = ~b_34 & ~b_35;
assign w4177 = b_34 & b_35;
assign w4178 = ~w4176 & ~w4177;
assign w4179 = (w1931 & w38768) | (w1931 & w38769) | (w38768 & w38769);
assign w4180 = (~w1931 & w38770) | (~w1931 & w38771) | (w38770 & w38771);
assign w4181 = ~w4179 & ~w4180;
assign w4182 = (w4175 & ~w4181) | (w4175 & w28494) | (~w4181 & w28494);
assign w4183 = (w4181 & w38772) | (w4181 & w38773) | (w38772 & w38773);
assign w4184 = (~w4181 & w38774) | (~w4181 & w38775) | (w38774 & w38775);
assign w4185 = ~w4182 & ~w4183;
assign w4186 = ~w4184 & ~w4185;
assign w4187 = (w4186 & w4168) | (w4186 & w28495) | (w4168 & w28495);
assign w4188 = ~w4168 & w28496;
assign w4189 = ~w4187 & ~w4188;
assign w4190 = ~w3980 & ~w4189;
assign w4191 = w3980 & w4189;
assign w4192 = ~w4190 & ~w4191;
assign w4193 = b_33 & w99;
assign w4194 = w136 & w28497;
assign w4195 = b_32 & w94;
assign w4196 = ~w4194 & ~w4195;
assign w4197 = ~w4193 & w4196;
assign w4198 = (w4197 & ~w3744) | (w4197 & w28498) | (~w3744 & w28498);
assign w4199 = (w3744 & w38776) | (w3744 & w38777) | (w38776 & w38777);
assign w4200 = (~w3744 & w38778) | (~w3744 & w38779) | (w38778 & w38779);
assign w4201 = ~w4198 & ~w4199;
assign w4202 = ~w4200 & ~w4201;
assign w4203 = (~w4146 & w4150) | (~w4146 & w27409) | (w4150 & w27409);
assign w4204 = (~w4141 & w3920) | (~w4141 & w27336) | (w3920 & w27336);
assign w4205 = b_27 & w418;
assign w4206 = w481 & w28499;
assign w4207 = b_26 & w413;
assign w4208 = ~w4206 & ~w4207;
assign w4209 = ~w4205 & w4208;
assign w4210 = (w4209 & ~w2582) | (w4209 & w28500) | (~w2582 & w28500);
assign w4211 = (w2582 & w38780) | (w2582 & w38781) | (w38780 & w38781);
assign w4212 = (~w2582 & w38782) | (~w2582 & w38783) | (w38782 & w38783);
assign w4213 = ~w4210 & ~w4211;
assign w4214 = ~w4212 & ~w4213;
assign w4215 = (~w4135 & ~w4136) | (~w4135 & w28501) | (~w4136 & w28501);
assign w4216 = (~w4099 & w4103) | (~w4099 & w28502) | (w4103 & w28502);
assign w4217 = (~w4094 & ~w4095) | (~w4094 & w27026) | (~w4095 & w27026);
assign w4218 = b_15 & w1694;
assign w4219 = w1834 & w28503;
assign w4220 = b_14 & w1689;
assign w4221 = ~w4219 & ~w4220;
assign w4222 = ~w4218 & w4221;
assign w4223 = (w4222 & ~w827) | (w4222 & w28504) | (~w827 & w28504);
assign w4224 = (w827 & w38784) | (w827 & w38785) | (w38784 & w38785);
assign w4225 = (~w827 & w38786) | (~w827 & w38787) | (w38786 & w38787);
assign w4226 = ~w4223 & ~w4224;
assign w4227 = ~w4225 & ~w4226;
assign w4228 = (~w4070 & w4073) | (~w4070 & w26899) | (w4073 & w26899);
assign w4229 = b_6 & w3195;
assign w4230 = w3388 & w28505;
assign w4231 = b_5 & w3190;
assign w4232 = ~w4230 & ~w4231;
assign w4233 = ~w4229 & w4232;
assign w4234 = (w4233 & ~w190) | (w4233 & w28506) | (~w190 & w28506);
assign w4235 = (w190 & w38788) | (w190 & w38789) | (w38788 & w38789);
assign w4236 = (~w190 & w38790) | (~w190 & w38791) | (w38790 & w38791);
assign w4237 = ~w4234 & ~w4235;
assign w4238 = ~w4236 & ~w4237;
assign w4239 = a_35 & ~a_36;
assign w4240 = ~a_35 & a_36;
assign w4241 = ~w4239 & ~w4240;
assign w4242 = b_0 & ~w4241;
assign w4243 = (w4242 & w4037) | (w4242 & w25790) | (w4037 & w25790);
assign w4244 = ~w4037 & w25791;
assign w4245 = ~w4243 & ~w4244;
assign w4246 = b_3 & w3803;
assign w4247 = w4027 & w26137;
assign w4248 = b_2 & w3798;
assign w4249 = ~w4247 & ~w4248;
assign w4250 = ~w4246 & w4249;
assign w4251 = w57 & w3806;
assign w4252 = w4250 & ~w4251;
assign w4253 = a_35 & ~w4252;
assign w4254 = w4252 & a_35;
assign w4255 = ~w4252 & ~w4253;
assign w4256 = ~w4254 & ~w4255;
assign w4257 = ~w4245 & ~w4256;
assign w4258 = w4245 & w4256;
assign w4259 = ~w4257 & ~w4258;
assign w4260 = ~w4238 & w4259;
assign w4261 = w4259 & ~w4260;
assign w4262 = ~w4259 & ~w4238;
assign w4263 = ~w4261 & ~w4262;
assign w4264 = ~w4056 & w4263;
assign w4265 = w4056 & ~w4263;
assign w4266 = ~w4264 & ~w4265;
assign w4267 = b_9 & w2639;
assign w4268 = w2820 & w28507;
assign w4269 = b_8 & w2634;
assign w4270 = ~w4268 & ~w4269;
assign w4271 = ~w4267 & w4270;
assign w4272 = (w4271 & ~w371) | (w4271 & w28508) | (~w371 & w28508);
assign w4273 = (w371 & w38792) | (w371 & w38793) | (w38792 & w38793);
assign w4274 = (~w371 & w38794) | (~w371 & w38795) | (w38794 & w38795);
assign w4275 = ~w4272 & ~w4273;
assign w4276 = ~w4274 & ~w4275;
assign w4277 = ~w4266 & ~w4276;
assign w4278 = w4266 & w4276;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = w4228 & ~w4279;
assign w4281 = ~w4228 & w4279;
assign w4282 = ~w4280 & ~w4281;
assign w4283 = b_12 & w2158;
assign w4284 = w2294 & w28509;
assign w4285 = b_11 & w2153;
assign w4286 = ~w4284 & ~w4285;
assign w4287 = ~w4283 & w4286;
assign w4288 = (w4287 & ~w552) | (w4287 & w28510) | (~w552 & w28510);
assign w4289 = (w552 & w38796) | (w552 & w38797) | (w38796 & w38797);
assign w4290 = (~w552 & w38798) | (~w552 & w38799) | (w38798 & w38799);
assign w4291 = ~w4288 & ~w4289;
assign w4292 = ~w4290 & ~w4291;
assign w4293 = ~w4282 & w4292;
assign w4294 = w4282 & ~w4292;
assign w4295 = ~w4293 & ~w4294;
assign w4296 = (~w4077 & w4080) | (~w4077 & w26900) | (w4080 & w26900);
assign w4297 = w4295 & ~w4296;
assign w4298 = ~w4295 & w4296;
assign w4299 = ~w4297 & ~w4298;
assign w4300 = ~w4227 & w4299;
assign w4301 = w4299 & ~w4300;
assign w4302 = ~w4299 & ~w4227;
assign w4303 = ~w4301 & ~w4302;
assign w4304 = ~w4217 & w4303;
assign w4305 = w4217 & ~w4303;
assign w4306 = ~w4304 & ~w4305;
assign w4307 = b_18 & w1295;
assign w4308 = w1422 & w28511;
assign w4309 = b_17 & w1290;
assign w4310 = ~w4308 & ~w4309;
assign w4311 = ~w4307 & w4310;
assign w4312 = (w4311 & ~w1238) | (w4311 & w28512) | (~w1238 & w28512);
assign w4313 = (w1238 & w38800) | (w1238 & w38801) | (w38800 & w38801);
assign w4314 = (~w1238 & w38802) | (~w1238 & w38803) | (w38802 & w38803);
assign w4315 = ~w4312 & ~w4313;
assign w4316 = ~w4314 & ~w4315;
assign w4317 = ~w4306 & ~w4316;
assign w4318 = w4306 & w4316;
assign w4319 = ~w4317 & ~w4318;
assign w4320 = w4216 & ~w4319;
assign w4321 = ~w4216 & w4319;
assign w4322 = ~w4320 & ~w4321;
assign w4323 = b_21 & w986;
assign w4324 = w1069 & w28513;
assign w4325 = b_20 & w981;
assign w4326 = ~w4324 & ~w4325;
assign w4327 = ~w4323 & w4326;
assign w4328 = (w4327 & ~w1634) | (w4327 & w28514) | (~w1634 & w28514);
assign w4329 = (w1634 & w38804) | (w1634 & w38805) | (w38804 & w38805);
assign w4330 = (~w1634 & w38806) | (~w1634 & w38807) | (w38806 & w38807);
assign w4331 = ~w4328 & ~w4329;
assign w4332 = ~w4330 & ~w4331;
assign w4333 = w4322 & ~w4332;
assign w4334 = w4322 & ~w4333;
assign w4335 = ~w4322 & ~w4332;
assign w4336 = ~w4334 & ~w4335;
assign w4337 = ~w4121 & w4336;
assign w4338 = w4121 & ~w4336;
assign w4339 = ~w4337 & ~w4338;
assign w4340 = b_24 & w657;
assign w4341 = w754 & w28515;
assign w4342 = b_23 & w652;
assign w4343 = ~w4341 & ~w4342;
assign w4344 = ~w4340 & w4343;
assign w4345 = (w4344 & ~w2083) | (w4344 & w28516) | (~w2083 & w28516);
assign w4346 = (w2083 & w38808) | (w2083 & w38809) | (w38808 & w38809);
assign w4347 = (~w2083 & w38810) | (~w2083 & w38811) | (w38810 & w38811);
assign w4348 = ~w4345 & ~w4346;
assign w4349 = ~w4347 & ~w4348;
assign w4350 = w4339 & w4349;
assign w4351 = ~w4339 & ~w4349;
assign w4352 = ~w4350 & ~w4351;
assign w4353 = ~w4215 & w4352;
assign w4354 = w4215 & ~w4352;
assign w4355 = ~w4353 & ~w4354;
assign w4356 = ~w4214 & w4355;
assign w4357 = w4355 & ~w4356;
assign w4358 = ~w4355 & ~w4214;
assign w4359 = ~w4357 & ~w4358;
assign w4360 = ~w4204 & w4359;
assign w4361 = w4204 & ~w4359;
assign w4362 = ~w4360 & ~w4361;
assign w4363 = b_30 & w239;
assign w4364 = w266 & w28517;
assign w4365 = b_29 & w234;
assign w4366 = ~w4364 & ~w4365;
assign w4367 = ~w4363 & w4366;
assign w4368 = (w4367 & ~w3138) | (w4367 & w28518) | (~w3138 & w28518);
assign w4369 = (w3138 & w38812) | (w3138 & w38813) | (w38812 & w38813);
assign w4370 = (~w3138 & w38814) | (~w3138 & w38815) | (w38814 & w38815);
assign w4371 = ~w4368 & ~w4369;
assign w4372 = ~w4370 & ~w4371;
assign w4373 = w4362 & w4372;
assign w4374 = ~w4362 & ~w4372;
assign w4375 = ~w4373 & ~w4374;
assign w4376 = ~w4203 & w4375;
assign w4377 = w4203 & ~w4375;
assign w4378 = ~w4376 & ~w4377;
assign w4379 = ~w4202 & w4378;
assign w4380 = w4202 & ~w4378;
assign w4381 = ~w4379 & ~w4380;
assign w4382 = ~w4169 & w4381;
assign w4383 = w4169 & ~w4381;
assign w4384 = ~w4382 & ~w4383;
assign w4385 = w8 & w28519;
assign w4386 = ~w8 & w28520;
assign w4387 = b_35 & w4;
assign w4388 = ~w4386 & ~w4387;
assign w4389 = ~w4385 & w4388;
assign w4390 = ~b_35 & ~b_36;
assign w4391 = b_35 & b_36;
assign w4392 = ~w4390 & ~w4391;
assign w4393 = (w1931 & w38816) | (w1931 & w38817) | (w38816 & w38817);
assign w4394 = (~w1931 & w38818) | (~w1931 & w38819) | (w38818 & w38819);
assign w4395 = ~w4393 & ~w4394;
assign w4396 = (w4389 & ~w4395) | (w4389 & w28526) | (~w4395 & w28526);
assign w4397 = (w4395 & w38820) | (w4395 & w38821) | (w38820 & w38821);
assign w4398 = (~w4395 & w38822) | (~w4395 & w38823) | (w38822 & w38823);
assign w4399 = ~w4396 & ~w4397;
assign w4400 = ~w4398 & ~w4399;
assign w4401 = w4384 & ~w4400;
assign w4402 = w4384 & ~w4401;
assign w4403 = ~w4384 & ~w4400;
assign w4404 = ~w4402 & ~w4403;
assign w4405 = (~w4186 & w4168) | (~w4186 & w28527) | (w4168 & w28527);
assign w4406 = ~w4190 & ~w4405;
assign w4407 = ~w4404 & ~w4406;
assign w4408 = w4404 & w4406;
assign w4409 = ~w4407 & ~w4408;
assign w4410 = (~w4401 & w4406) | (~w4401 & w28528) | (w4406 & w28528);
assign w4411 = b_34 & w99;
assign w4412 = w136 & w28529;
assign w4413 = b_33 & w94;
assign w4414 = ~w4412 & ~w4413;
assign w4415 = ~w4411 & w4414;
assign w4416 = (w4415 & ~w3967) | (w4415 & w28530) | (~w3967 & w28530);
assign w4417 = (w3967 & w38824) | (w3967 & w38825) | (w38824 & w38825);
assign w4418 = (~w3967 & w38826) | (~w3967 & w38827) | (w38826 & w38827);
assign w4419 = ~w4416 & ~w4417;
assign w4420 = ~w4418 & ~w4419;
assign w4421 = (~w4374 & w4203) | (~w4374 & w27525) | (w4203 & w27525);
assign w4422 = b_31 & w239;
assign w4423 = w266 & w28531;
assign w4424 = b_30 & w234;
assign w4425 = ~w4423 & ~w4424;
assign w4426 = ~w4422 & w4425;
assign w4427 = (w4426 & ~w3345) | (w4426 & w28532) | (~w3345 & w28532);
assign w4428 = (w3345 & w38828) | (w3345 & w38829) | (w38828 & w38829);
assign w4429 = (~w3345 & w38830) | (~w3345 & w38831) | (w38830 & w38831);
assign w4430 = ~w4427 & ~w4428;
assign w4431 = ~w4429 & ~w4430;
assign w4432 = (~w4356 & w4359) | (~w4356 & w27337) | (w4359 & w27337);
assign w4433 = (~w4351 & w4215) | (~w4351 & w27131) | (w4215 & w27131);
assign w4434 = b_16 & w1694;
assign w4435 = w1834 & w28533;
assign w4436 = b_15 & w1689;
assign w4437 = ~w4435 & ~w4436;
assign w4438 = ~w4434 & w4437;
assign w4439 = (w4438 & ~w926) | (w4438 & w28534) | (~w926 & w28534);
assign w4440 = (w926 & w38832) | (w926 & w38833) | (w38832 & w38833);
assign w4441 = (~w926 & w38834) | (~w926 & w38835) | (w38834 & w38835);
assign w4442 = ~w4439 & ~w4440;
assign w4443 = ~w4441 & ~w4442;
assign w4444 = (~w4294 & w4296) | (~w4294 & w27027) | (w4296 & w27027);
assign w4445 = b_13 & w2158;
assign w4446 = w2294 & w28535;
assign w4447 = b_12 & w2153;
assign w4448 = ~w4446 & ~w4447;
assign w4449 = ~w4445 & w4448;
assign w4450 = (w4449 & ~w711) | (w4449 & w28536) | (~w711 & w28536);
assign w4451 = (w711 & w38836) | (w711 & w38837) | (w38836 & w38837);
assign w4452 = (~w711 & w38838) | (~w711 & w38839) | (w38838 & w38839);
assign w4453 = ~w4450 & ~w4451;
assign w4454 = ~w4452 & ~w4453;
assign w4455 = (~w4277 & w4228) | (~w4277 & w27028) | (w4228 & w27028);
assign w4456 = b_10 & w2639;
assign w4457 = w2820 & w28537;
assign w4458 = b_9 & w2634;
assign w4459 = ~w4457 & ~w4458;
assign w4460 = ~w4456 & w4459;
assign w4461 = (w4460 & ~w454) | (w4460 & w28538) | (~w454 & w28538);
assign w4462 = (w454 & w38840) | (w454 & w38841) | (w38840 & w38841);
assign w4463 = (~w454 & w38842) | (~w454 & w38843) | (w38842 & w38843);
assign w4464 = ~w4461 & ~w4462;
assign w4465 = ~w4463 & ~w4464;
assign w4466 = (~w4260 & w4263) | (~w4260 & w26784) | (w4263 & w26784);
assign w4467 = b_7 & w3195;
assign w4468 = w3388 & w28539;
assign w4469 = b_6 & w3190;
assign w4470 = ~w4468 & ~w4469;
assign w4471 = ~w4467 & w4470;
assign w4472 = (w4471 & ~w213) | (w4471 & w28540) | (~w213 & w28540);
assign w4473 = (w213 & w38844) | (w213 & w38845) | (w38844 & w38845);
assign w4474 = (~w213 & w38846) | (~w213 & w38847) | (w38846 & w38847);
assign w4475 = ~w4472 & ~w4473;
assign w4476 = ~w4474 & ~w4475;
assign w4477 = ~w4037 & w28541;
assign w4478 = (~w4477 & w4245) | (~w4477 & w28542) | (w4245 & w28542);
assign w4479 = b_4 & w3803;
assign w4480 = w4027 & w26138;
assign w4481 = b_3 & w3798;
assign w4482 = ~w4480 & ~w4481;
assign w4483 = ~w4479 & w4482;
assign w4484 = w84 & w3806;
assign w4485 = w4483 & ~w4484;
assign w4486 = (a_35 & w4484) | (a_35 & w26139) | (w4484 & w26139);
assign w4487 = ~w4484 & w26545;
assign w4488 = ~w4485 & ~w4486;
assign w4489 = ~w4487 & ~w4488;
assign w4490 = (a_38 & w4241) | (a_38 & w28543) | (w4241 & w28543);
assign w4491 = ~a_36 & a_37;
assign w4492 = a_36 & ~a_37;
assign w4493 = ~w4491 & ~w4492;
assign w4494 = w4241 & ~w4493;
assign w4495 = b_0 & w4494;
assign w4496 = ~a_37 & a_38;
assign w4497 = a_37 & ~a_38;
assign w4498 = ~w4496 & ~w4497;
assign w4499 = ~w4241 & w4498;
assign w4500 = b_1 & w4499;
assign w4501 = ~w4495 & ~w4500;
assign w4502 = ~w4241 & ~w4498;
assign w4503 = ~w15 & w4502;
assign w4504 = w4501 & ~w4503;
assign w4505 = (a_38 & ~w4501) | (a_38 & w25547) | (~w4501 & w25547);
assign w4506 = w4501 & w25792;
assign w4507 = ~w4504 & ~w4505;
assign w4508 = (w4490 & w4507) | (w4490 & w25793) | (w4507 & w25793);
assign w4509 = ~w4507 & w26546;
assign w4510 = ~w4508 & ~w4509;
assign w4511 = w4489 & ~w4510;
assign w4512 = ~w4489 & w4510;
assign w4513 = ~w4511 & ~w4512;
assign w4514 = ~w4478 & w4513;
assign w4515 = w4478 & ~w4513;
assign w4516 = ~w4514 & ~w4515;
assign w4517 = w4476 & ~w4516;
assign w4518 = ~w4476 & w4516;
assign w4519 = ~w4517 & ~w4518;
assign w4520 = ~w4466 & w4519;
assign w4521 = w4466 & ~w4519;
assign w4522 = ~w4520 & ~w4521;
assign w4523 = w4465 & ~w4522;
assign w4524 = ~w4465 & w4522;
assign w4525 = ~w4523 & ~w4524;
assign w4526 = ~w4455 & w4525;
assign w4527 = w4455 & ~w4525;
assign w4528 = ~w4526 & ~w4527;
assign w4529 = w4454 & ~w4528;
assign w4530 = ~w4454 & w4528;
assign w4531 = ~w4529 & ~w4530;
assign w4532 = ~w4444 & w4531;
assign w4533 = w4444 & ~w4531;
assign w4534 = ~w4532 & ~w4533;
assign w4535 = ~w4443 & w4534;
assign w4536 = w4534 & ~w4535;
assign w4537 = ~w4534 & ~w4443;
assign w4538 = ~w4536 & ~w4537;
assign w4539 = (~w4300 & w4303) | (~w4300 & w27029) | (w4303 & w27029);
assign w4540 = w4538 & w4539;
assign w4541 = ~w4538 & ~w4539;
assign w4542 = ~w4540 & ~w4541;
assign w4543 = b_19 & w1295;
assign w4544 = w1422 & w28544;
assign w4545 = b_18 & w1290;
assign w4546 = ~w4544 & ~w4545;
assign w4547 = ~w4543 & w4546;
assign w4548 = (w4547 & ~w1372) | (w4547 & w28545) | (~w1372 & w28545);
assign w4549 = (w1372 & w38848) | (w1372 & w38849) | (w38848 & w38849);
assign w4550 = (~w1372 & w38850) | (~w1372 & w38851) | (w38850 & w38851);
assign w4551 = ~w4548 & ~w4549;
assign w4552 = ~w4550 & ~w4551;
assign w4553 = w4542 & ~w4552;
assign w4554 = w4542 & ~w4553;
assign w4555 = ~w4542 & ~w4552;
assign w4556 = ~w4554 & ~w4555;
assign w4557 = (~w4317 & w4216) | (~w4317 & w27030) | (w4216 & w27030);
assign w4558 = w4556 & w4557;
assign w4559 = ~w4556 & ~w4557;
assign w4560 = ~w4558 & ~w4559;
assign w4561 = b_22 & w986;
assign w4562 = w1069 & w28546;
assign w4563 = b_21 & w981;
assign w4564 = ~w4562 & ~w4563;
assign w4565 = ~w4561 & w4564;
assign w4566 = (w4565 & ~w1786) | (w4565 & w28547) | (~w1786 & w28547);
assign w4567 = (w1786 & w38852) | (w1786 & w38853) | (w38852 & w38853);
assign w4568 = (~w1786 & w38854) | (~w1786 & w38855) | (w38854 & w38855);
assign w4569 = ~w4566 & ~w4567;
assign w4570 = ~w4568 & ~w4569;
assign w4571 = w4560 & ~w4570;
assign w4572 = w4560 & ~w4571;
assign w4573 = ~w4560 & ~w4570;
assign w4574 = ~w4572 & ~w4573;
assign w4575 = (~w4333 & w4336) | (~w4333 & w27132) | (w4336 & w27132);
assign w4576 = w4574 & w4575;
assign w4577 = ~w4574 & ~w4575;
assign w4578 = ~w4576 & ~w4577;
assign w4579 = b_25 & w657;
assign w4580 = w754 & w28548;
assign w4581 = b_24 & w652;
assign w4582 = ~w4580 & ~w4581;
assign w4583 = ~w4579 & w4582;
assign w4584 = (w4583 & ~w2108) | (w4583 & w28549) | (~w2108 & w28549);
assign w4585 = (w2108 & w38856) | (w2108 & w38857) | (w38856 & w38857);
assign w4586 = (~w2108 & w38858) | (~w2108 & w38859) | (w38858 & w38859);
assign w4587 = ~w4584 & ~w4585;
assign w4588 = ~w4586 & ~w4587;
assign w4589 = w4578 & ~w4588;
assign w4590 = ~w4578 & w4588;
assign w4591 = ~w4433 & w27209;
assign w4592 = ~w4433 & ~w4591;
assign w4593 = (~w4589 & w4433) | (~w4589 & w27338) | (w4433 & w27338);
assign w4594 = (w27338 & w27209) | (w27338 & w28550) | (w27209 & w28550);
assign w4595 = ~w4592 & ~w4594;
assign w4596 = b_28 & w418;
assign w4597 = w481 & w28551;
assign w4598 = b_27 & w413;
assign w4599 = ~w4597 & ~w4598;
assign w4600 = ~w4596 & w4599;
assign w4601 = (w4600 & ~w2771) | (w4600 & w28552) | (~w2771 & w28552);
assign w4602 = (w2771 & w38860) | (w2771 & w38861) | (w38860 & w38861);
assign w4603 = (~w2771 & w38862) | (~w2771 & w38863) | (w38862 & w38863);
assign w4604 = ~w4601 & ~w4602;
assign w4605 = ~w4603 & ~w4604;
assign w4606 = w4595 & w4605;
assign w4607 = ~w4595 & ~w4605;
assign w4608 = ~w4606 & ~w4607;
assign w4609 = ~w4432 & w4608;
assign w4610 = w4432 & ~w4608;
assign w4611 = ~w4609 & ~w4610;
assign w4612 = w4431 & ~w4611;
assign w4613 = ~w4431 & w4611;
assign w4614 = ~w4612 & ~w4613;
assign w4615 = ~w4421 & w4614;
assign w4616 = w4421 & ~w4614;
assign w4617 = ~w4615 & ~w4616;
assign w4618 = ~w4420 & w4617;
assign w4619 = w4617 & ~w4618;
assign w4620 = ~w4617 & ~w4420;
assign w4621 = ~w4619 & ~w4620;
assign w4622 = (~w4379 & w4169) | (~w4379 & w28553) | (w4169 & w28553);
assign w4623 = w4621 & w4622;
assign w4624 = ~w4621 & ~w4622;
assign w4625 = ~w4623 & ~w4624;
assign w4626 = w8 & w28554;
assign w4627 = ~w8 & w28555;
assign w4628 = b_36 & w4;
assign w4629 = ~w4627 & ~w4628;
assign w4630 = ~w4626 & w4629;
assign w4631 = ~b_36 & ~b_37;
assign w4632 = b_36 & b_37;
assign w4633 = ~w4631 & ~w4632;
assign w4634 = (w1931 & w38864) | (w1931 & w38865) | (w38864 & w38865);
assign w4635 = (~w1931 & w38866) | (~w1931 & w38867) | (w38866 & w38867);
assign w4636 = ~w4634 & ~w4635;
assign w4637 = (w4630 & ~w4636) | (w4630 & w28561) | (~w4636 & w28561);
assign w4638 = (w4636 & w38868) | (w4636 & w38869) | (w38868 & w38869);
assign w4639 = (~w4636 & w38870) | (~w4636 & w38871) | (w38870 & w38871);
assign w4640 = ~w4637 & ~w4638;
assign w4641 = ~w4639 & ~w4640;
assign w4642 = ~w4625 & w4641;
assign w4643 = w4625 & ~w4641;
assign w4644 = ~w4642 & ~w4643;
assign w4645 = ~w4410 & w4644;
assign w4646 = w4410 & ~w4644;
assign w4647 = ~w4645 & ~w4646;
assign w4648 = w8 & w28562;
assign w4649 = ~w8 & w28563;
assign w4650 = b_37 & w4;
assign w4651 = ~w4649 & ~w4650;
assign w4652 = ~w4648 & w4651;
assign w4653 = ~b_37 & ~b_38;
assign w4654 = b_37 & b_38;
assign w4655 = ~w4653 & ~w4654;
assign w4656 = (w1931 & w38872) | (w1931 & w38873) | (w38872 & w38873);
assign w4657 = (~w1931 & w38874) | (~w1931 & w38875) | (w38874 & w38875);
assign w4658 = ~w4656 & ~w4657;
assign w4659 = (w4652 & ~w4658) | (w4652 & w28569) | (~w4658 & w28569);
assign w4660 = (w4658 & w38876) | (w4658 & w38877) | (w38876 & w38877);
assign w4661 = (~w4658 & w38878) | (~w4658 & w38879) | (w38878 & w38879);
assign w4662 = ~w4659 & ~w4660;
assign w4663 = ~w4661 & ~w4662;
assign w4664 = (~w4618 & w4621) | (~w4618 & w28570) | (w4621 & w28570);
assign w4665 = b_35 & w99;
assign w4666 = w136 & w28571;
assign w4667 = b_34 & w94;
assign w4668 = ~w4666 & ~w4667;
assign w4669 = ~w4665 & w4668;
assign w4670 = (w4669 & ~w4181) | (w4669 & w28572) | (~w4181 & w28572);
assign w4671 = (w4181 & w38880) | (w4181 & w38881) | (w38880 & w38881);
assign w4672 = (~w4181 & w38882) | (~w4181 & w38883) | (w38882 & w38883);
assign w4673 = ~w4670 & ~w4671;
assign w4674 = ~w4672 & ~w4673;
assign w4675 = (~w4613 & w4421) | (~w4613 & w27734) | (w4421 & w27734);
assign w4676 = b_32 & w239;
assign w4677 = w266 & w28573;
assign w4678 = b_31 & w234;
assign w4679 = ~w4677 & ~w4678;
assign w4680 = ~w4676 & w4679;
assign w4681 = (w4680 & ~w3545) | (w4680 & w28574) | (~w3545 & w28574);
assign w4682 = (w3545 & w38884) | (w3545 & w38885) | (w38884 & w38885);
assign w4683 = (~w3545 & w38886) | (~w3545 & w38887) | (w38886 & w38887);
assign w4684 = ~w4681 & ~w4682;
assign w4685 = ~w4683 & ~w4684;
assign w4686 = (~w4607 & w4432) | (~w4607 & w28575) | (w4432 & w28575);
assign w4687 = b_29 & w418;
assign w4688 = w481 & w28576;
assign w4689 = b_28 & w413;
assign w4690 = ~w4688 & ~w4689;
assign w4691 = ~w4687 & w4690;
assign w4692 = (w4691 & ~w2954) | (w4691 & w28577) | (~w2954 & w28577);
assign w4693 = (w2954 & w38888) | (w2954 & w38889) | (w38888 & w38889);
assign w4694 = (~w2954 & w38890) | (~w2954 & w38891) | (w38890 & w38891);
assign w4695 = ~w4692 & ~w4693;
assign w4696 = ~w4694 & ~w4695;
assign w4697 = ~w4571 & ~w4577;
assign w4698 = b_17 & w1694;
assign w4699 = w1834 & w28578;
assign w4700 = b_16 & w1689;
assign w4701 = ~w4699 & ~w4700;
assign w4702 = ~w4698 & w4701;
assign w4703 = (w4702 & ~w1038) | (w4702 & w28579) | (~w1038 & w28579);
assign w4704 = (w1038 & w38892) | (w1038 & w38893) | (w38892 & w38893);
assign w4705 = (~w1038 & w38894) | (~w1038 & w38895) | (w38894 & w38895);
assign w4706 = ~w4703 & ~w4704;
assign w4707 = ~w4705 & ~w4706;
assign w4708 = (~w4530 & w4444) | (~w4530 & w27133) | (w4444 & w27133);
assign w4709 = (~w4524 & w4455) | (~w4524 & w27134) | (w4455 & w27134);
assign w4710 = b_11 & w2639;
assign w4711 = w2820 & w28580;
assign w4712 = b_10 & w2634;
assign w4713 = ~w4711 & ~w4712;
assign w4714 = ~w4710 & w4713;
assign w4715 = (w4714 & ~w530) | (w4714 & w28581) | (~w530 & w28581);
assign w4716 = (w530 & w38896) | (w530 & w38897) | (w38896 & w38897);
assign w4717 = (~w530 & w38898) | (~w530 & w38899) | (w38898 & w38899);
assign w4718 = ~w4715 & ~w4716;
assign w4719 = ~w4717 & ~w4718;
assign w4720 = (~w4518 & w4466) | (~w4518 & w28582) | (w4466 & w28582);
assign w4721 = (~w4512 & w4478) | (~w4512 & w26140) | (w4478 & w26140);
assign w4722 = b_2 & w4499;
assign w4723 = w4241 & ~w4498;
assign w4724 = w4723 & w25369;
assign w4725 = b_1 & w4494;
assign w4726 = ~w4724 & ~w4725;
assign w4727 = ~w4722 & w4726;
assign w4728 = w35 & w4502;
assign w4729 = w4727 & ~w4728;
assign w4730 = (a_38 & ~w4727) | (a_38 & w25548) | (~w4727 & w25548);
assign w4731 = w4727 & w25794;
assign w4732 = ~w4729 & ~w4730;
assign w4733 = ~w4731 & ~w4732;
assign w4734 = ~w4508 & w4733;
assign w4735 = w4508 & ~w4733;
assign w4736 = ~w4734 & ~w4735;
assign w4737 = b_5 & w3803;
assign w4738 = w4027 & w26547;
assign w4739 = b_4 & w3798;
assign w4740 = ~w4738 & ~w4739;
assign w4741 = ~w4737 & w4740;
assign w4742 = w129 & w3806;
assign w4743 = w4741 & ~w4742;
assign w4744 = (a_35 & w4742) | (a_35 & w26548) | (w4742 & w26548);
assign w4745 = ~w4742 & w38900;
assign w4746 = ~w4743 & ~w4744;
assign w4747 = ~w4745 & ~w4746;
assign w4748 = w4736 & ~w4747;
assign w4749 = w4736 & ~w4748;
assign w4750 = ~w4736 & ~w4747;
assign w4751 = ~w4749 & ~w4750;
assign w4752 = ~w4721 & w4751;
assign w4753 = w4721 & ~w4751;
assign w4754 = ~w4752 & ~w4753;
assign w4755 = b_8 & w3195;
assign w4756 = w3388 & w28583;
assign w4757 = b_7 & w3190;
assign w4758 = ~w4756 & ~w4757;
assign w4759 = ~w4755 & w4758;
assign w4760 = ~w308 & w28584;
assign w4761 = (w4759 & ~w28584) | (w4759 & w38901) | (~w28584 & w38901);
assign w4762 = (w28584 & w38902) | (w28584 & w38903) | (w38902 & w38903);
assign w4763 = ~w4760 & w28586;
assign w4764 = ~w4761 & ~w4762;
assign w4765 = ~w4763 & ~w4764;
assign w4766 = ~w4754 & ~w4765;
assign w4767 = w4754 & w4765;
assign w4768 = ~w4766 & ~w4767;
assign w4769 = ~w4720 & w4768;
assign w4770 = w4720 & ~w4768;
assign w4771 = ~w4769 & ~w4770;
assign w4772 = ~w4719 & w4771;
assign w4773 = ~w4771 & ~w4719;
assign w4774 = w4771 & ~w4772;
assign w4775 = ~w4773 & ~w4774;
assign w4776 = ~w4709 & ~w4775;
assign w4777 = ~w4775 & ~w4776;
assign w4778 = b_14 & w2158;
assign w4779 = w2294 & w28587;
assign w4780 = b_13 & w2153;
assign w4781 = ~w4779 & ~w4780;
assign w4782 = ~w4778 & w4781;
assign w4783 = (w4782 & ~w735) | (w4782 & w28588) | (~w735 & w28588);
assign w4784 = (w735 & w38904) | (w735 & w38905) | (w38904 & w38905);
assign w4785 = (~w735 & w38906) | (~w735 & w38907) | (w38906 & w38907);
assign w4786 = ~w4783 & ~w4784;
assign w4787 = ~w4785 & ~w4786;
assign w4788 = ~w4777 & w27135;
assign w4789 = (~w4787 & w4777) | (~w4787 & w27136) | (w4777 & w27136);
assign w4790 = ~w4788 & ~w4789;
assign w4791 = ~w4708 & w4790;
assign w4792 = w4708 & ~w4790;
assign w4793 = ~w4791 & ~w4792;
assign w4794 = ~w4707 & w4793;
assign w4795 = w4793 & ~w4794;
assign w4796 = ~w4793 & ~w4707;
assign w4797 = ~w4795 & ~w4796;
assign w4798 = (~w4535 & w4538) | (~w4535 & w38908) | (w4538 & w38908);
assign w4799 = w4797 & w4798;
assign w4800 = ~w4797 & ~w4798;
assign w4801 = ~w4799 & ~w4800;
assign w4802 = b_20 & w1295;
assign w4803 = w1422 & w28589;
assign w4804 = b_19 & w1290;
assign w4805 = ~w4803 & ~w4804;
assign w4806 = ~w4802 & w4805;
assign w4807 = (w4806 & ~w1503) | (w4806 & w28590) | (~w1503 & w28590);
assign w4808 = (w1503 & w38909) | (w1503 & w38910) | (w38909 & w38910);
assign w4809 = (~w1503 & w38911) | (~w1503 & w38912) | (w38911 & w38912);
assign w4810 = ~w4807 & ~w4808;
assign w4811 = ~w4809 & ~w4810;
assign w4812 = w4801 & ~w4811;
assign w4813 = w4801 & ~w4812;
assign w4814 = ~w4801 & ~w4811;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = (~w4553 & w4556) | (~w4553 & w38913) | (w4556 & w38913);
assign w4817 = w4815 & w4816;
assign w4818 = ~w4815 & ~w4816;
assign w4819 = ~w4817 & ~w4818;
assign w4820 = b_23 & w986;
assign w4821 = w1069 & w28591;
assign w4822 = b_22 & w981;
assign w4823 = ~w4821 & ~w4822;
assign w4824 = ~w4820 & w4823;
assign w4825 = (w4824 & ~w1933) | (w4824 & w28592) | (~w1933 & w28592);
assign w4826 = (w1933 & w38914) | (w1933 & w38915) | (w38914 & w38915);
assign w4827 = (~w1933 & w38916) | (~w1933 & w38917) | (w38916 & w38917);
assign w4828 = ~w4825 & ~w4826;
assign w4829 = ~w4827 & ~w4828;
assign w4830 = w4819 & ~w4829;
assign w4831 = ~w4819 & w4829;
assign w4832 = (w4577 & w27339) | (w4577 & w27340) | (w27339 & w27340);
assign w4833 = ~w4697 & ~w4832;
assign w4834 = (~w4577 & w38918) | (~w4577 & w38919) | (w38918 & w38919);
assign w4835 = ~w4577 & w38920;
assign w4836 = b_26 & w657;
assign w4837 = w754 & w28593;
assign w4838 = b_25 & w652;
assign w4839 = ~w4837 & ~w4838;
assign w4840 = ~w4836 & w4839;
assign w4841 = (w4840 & ~w2416) | (w4840 & w28594) | (~w2416 & w28594);
assign w4842 = (w2416 & w38921) | (w2416 & w38922) | (w38921 & w38922);
assign w4843 = (~w2416 & w38923) | (~w2416 & w38924) | (w38923 & w38924);
assign w4844 = ~w4841 & ~w4842;
assign w4845 = ~w4843 & ~w4844;
assign w4846 = ~w4833 & w38925;
assign w4847 = (~w4845 & w4833) | (~w4845 & w38926) | (w4833 & w38926);
assign w4848 = ~w4846 & ~w4847;
assign w4849 = ~w4593 & w4848;
assign w4850 = w4593 & ~w4848;
assign w4851 = ~w4849 & ~w4850;
assign w4852 = w4696 & ~w4851;
assign w4853 = ~w4696 & w4851;
assign w4854 = ~w4852 & ~w4853;
assign w4855 = ~w4686 & w4854;
assign w4856 = w4686 & ~w4854;
assign w4857 = ~w4855 & ~w4856;
assign w4858 = w4685 & ~w4857;
assign w4859 = ~w4685 & w4857;
assign w4860 = ~w4858 & ~w4859;
assign w4861 = ~w4675 & w4860;
assign w4862 = w4675 & ~w4860;
assign w4863 = ~w4861 & ~w4862;
assign w4864 = w4674 & ~w4863;
assign w4865 = ~w4674 & w4863;
assign w4866 = ~w4864 & ~w4865;
assign w4867 = ~w4664 & w4866;
assign w4868 = w4664 & ~w4866;
assign w4869 = ~w4867 & ~w4868;
assign w4870 = ~w4663 & w4869;
assign w4871 = w4869 & ~w4870;
assign w4872 = ~w4869 & ~w4663;
assign w4873 = ~w4871 & ~w4872;
assign w4874 = (~w4643 & w4410) | (~w4643 & w28595) | (w4410 & w28595);
assign w4875 = ~w4873 & ~w4874;
assign w4876 = w4873 & w4874;
assign w4877 = ~w4875 & ~w4876;
assign w4878 = w8 & w28596;
assign w4879 = ~w8 & w28597;
assign w4880 = b_38 & w4;
assign w4881 = ~w4879 & ~w4880;
assign w4882 = ~w4878 & w4881;
assign w4883 = ~b_38 & ~b_39;
assign w4884 = b_38 & b_39;
assign w4885 = ~w4883 & ~w4884;
assign w4886 = (w4885 & w4656) | (w4885 & w28598) | (w4656 & w28598);
assign w4887 = ~w4656 & w28599;
assign w4888 = ~w4886 & ~w4887;
assign w4889 = (w4882 & ~w4888) | (w4882 & w28600) | (~w4888 & w28600);
assign w4890 = (w4888 & w38927) | (w4888 & w38928) | (w38927 & w38928);
assign w4891 = (~w4888 & w38929) | (~w4888 & w38930) | (w38929 & w38930);
assign w4892 = ~w4889 & ~w4890;
assign w4893 = ~w4891 & ~w4892;
assign w4894 = (~w4865 & w4664) | (~w4865 & w38931) | (w4664 & w38931);
assign w4895 = (~w4859 & w4675) | (~w4859 & w28601) | (w4675 & w28601);
assign w4896 = b_33 & w239;
assign w4897 = w266 & w28602;
assign w4898 = b_32 & w234;
assign w4899 = ~w4897 & ~w4898;
assign w4900 = ~w4896 & w4899;
assign w4901 = (w4900 & ~w3744) | (w4900 & w25037) | (~w3744 & w25037);
assign w4902 = (w3744 & w28603) | (w3744 & w28604) | (w28603 & w28604);
assign w4903 = (~w3744 & w28605) | (~w3744 & w28606) | (w28605 & w28606);
assign w4904 = ~w4901 & ~w4902;
assign w4905 = ~w4903 & ~w4904;
assign w4906 = (~w4853 & w4686) | (~w4853 & w25038) | (w4686 & w25038);
assign w4907 = (~w4847 & w4593) | (~w4847 & w38932) | (w4593 & w38932);
assign w4908 = b_27 & w657;
assign w4909 = w754 & w28607;
assign w4910 = b_26 & w652;
assign w4911 = ~w4909 & ~w4910;
assign w4912 = ~w4908 & w4911;
assign w4913 = (w4912 & ~w2582) | (w4912 & w28608) | (~w2582 & w28608);
assign w4914 = (w2582 & w38933) | (w2582 & w38934) | (w38933 & w38934);
assign w4915 = (~w2582 & w38935) | (~w2582 & w38936) | (w38935 & w38936);
assign w4916 = ~w4913 & ~w4914;
assign w4917 = ~w4915 & ~w4916;
assign w4918 = (~w4794 & w4798) | (~w4794 & w27137) | (w4798 & w27137);
assign w4919 = (~w4789 & w4708) | (~w4789 & w28609) | (w4708 & w28609);
assign w4920 = b_15 & w2158;
assign w4921 = w2294 & w28610;
assign w4922 = b_14 & w2153;
assign w4923 = ~w4921 & ~w4922;
assign w4924 = ~w4920 & w4923;
assign w4925 = (w4924 & ~w827) | (w4924 & w28611) | (~w827 & w28611);
assign w4926 = (w827 & w38937) | (w827 & w38938) | (w38937 & w38938);
assign w4927 = (~w827 & w38939) | (~w827 & w38940) | (w38939 & w38940);
assign w4928 = ~w4925 & ~w4926;
assign w4929 = ~w4927 & ~w4928;
assign w4930 = b_6 & w3803;
assign w4931 = w4027 & w28612;
assign w4932 = b_5 & w3798;
assign w4933 = ~w4931 & ~w4932;
assign w4934 = ~w4930 & w4933;
assign w4935 = (w4934 & ~w190) | (w4934 & w28613) | (~w190 & w28613);
assign w4936 = (w190 & w38941) | (w190 & w38942) | (w38941 & w38942);
assign w4937 = (~w190 & w38943) | (~w190 & w38944) | (w38943 & w38944);
assign w4938 = ~w4935 & ~w4936;
assign w4939 = ~w4937 & ~w4938;
assign w4940 = a_38 & ~a_39;
assign w4941 = ~a_38 & a_39;
assign w4942 = ~w4940 & ~w4941;
assign w4943 = b_0 & ~w4942;
assign w4944 = (w4943 & w4733) | (w4943 & w25795) | (w4733 & w25795);
assign w4945 = ~w4733 & w25796;
assign w4946 = ~w4944 & ~w4945;
assign w4947 = b_3 & w4499;
assign w4948 = w4723 & w26141;
assign w4949 = b_2 & w4494;
assign w4950 = ~w4948 & ~w4949;
assign w4951 = ~w4947 & w4950;
assign w4952 = w57 & w4502;
assign w4953 = w4951 & ~w4952;
assign w4954 = a_38 & ~w4953;
assign w4955 = w4953 & a_38;
assign w4956 = ~w4953 & ~w4954;
assign w4957 = ~w4955 & ~w4956;
assign w4958 = ~w4946 & ~w4957;
assign w4959 = w4946 & w4957;
assign w4960 = ~w4958 & ~w4959;
assign w4961 = ~w4939 & w4960;
assign w4962 = w4960 & ~w4961;
assign w4963 = ~w4960 & ~w4939;
assign w4964 = ~w4962 & ~w4963;
assign w4965 = ~w4721 & ~w4751;
assign w4966 = ~w4748 & ~w4965;
assign w4967 = w4964 & w4966;
assign w4968 = ~w4964 & ~w4966;
assign w4969 = ~w4967 & ~w4968;
assign w4970 = b_9 & w3195;
assign w4971 = w3388 & w28614;
assign w4972 = b_8 & w3190;
assign w4973 = ~w4971 & ~w4972;
assign w4974 = ~w4970 & w4973;
assign w4975 = (w4974 & ~w371) | (w4974 & w28615) | (~w371 & w28615);
assign w4976 = (w371 & w38945) | (w371 & w38946) | (w38945 & w38946);
assign w4977 = (~w371 & w38947) | (~w371 & w38948) | (w38947 & w38948);
assign w4978 = ~w4975 & ~w4976;
assign w4979 = ~w4977 & ~w4978;
assign w4980 = w4969 & ~w4979;
assign w4981 = w4969 & ~w4980;
assign w4982 = ~w4969 & ~w4979;
assign w4983 = ~w4981 & ~w4982;
assign w4984 = (~w4766 & w4720) | (~w4766 & w26901) | (w4720 & w26901);
assign w4985 = w4983 & w4984;
assign w4986 = ~w4983 & ~w4984;
assign w4987 = ~w4985 & ~w4986;
assign w4988 = b_12 & w2639;
assign w4989 = w2820 & w28616;
assign w4990 = b_11 & w2634;
assign w4991 = ~w4989 & ~w4990;
assign w4992 = ~w4988 & w4991;
assign w4993 = (w4992 & ~w552) | (w4992 & w28617) | (~w552 & w28617);
assign w4994 = (w552 & w38949) | (w552 & w38950) | (w38949 & w38950);
assign w4995 = (~w552 & w38951) | (~w552 & w38952) | (w38951 & w38952);
assign w4996 = ~w4993 & ~w4994;
assign w4997 = ~w4995 & ~w4996;
assign w4998 = ~w4987 & w4997;
assign w4999 = w4987 & ~w4997;
assign w5000 = ~w4998 & ~w4999;
assign w5001 = (~w4772 & w4775) | (~w4772 & w27138) | (w4775 & w27138);
assign w5002 = w5000 & ~w5001;
assign w5003 = ~w5000 & w5001;
assign w5004 = ~w5002 & ~w5003;
assign w5005 = ~w4929 & w5004;
assign w5006 = w5004 & ~w5005;
assign w5007 = ~w5004 & ~w4929;
assign w5008 = ~w5006 & ~w5007;
assign w5009 = ~w4919 & w5008;
assign w5010 = w4919 & ~w5008;
assign w5011 = ~w5009 & ~w5010;
assign w5012 = b_18 & w1694;
assign w5013 = w1834 & w28618;
assign w5014 = b_17 & w1689;
assign w5015 = ~w5013 & ~w5014;
assign w5016 = ~w5012 & w5015;
assign w5017 = (w5016 & ~w1238) | (w5016 & w28619) | (~w1238 & w28619);
assign w5018 = (w1238 & w38953) | (w1238 & w38954) | (w38953 & w38954);
assign w5019 = (~w1238 & w38955) | (~w1238 & w38956) | (w38955 & w38956);
assign w5020 = ~w5017 & ~w5018;
assign w5021 = ~w5019 & ~w5020;
assign w5022 = ~w5011 & ~w5021;
assign w5023 = w5011 & w5021;
assign w5024 = ~w5022 & ~w5023;
assign w5025 = w4918 & ~w5024;
assign w5026 = ~w4918 & w5024;
assign w5027 = ~w5025 & ~w5026;
assign w5028 = b_21 & w1295;
assign w5029 = w1422 & w28620;
assign w5030 = b_20 & w1290;
assign w5031 = ~w5029 & ~w5030;
assign w5032 = ~w5028 & w5031;
assign w5033 = (w5032 & ~w1634) | (w5032 & w28621) | (~w1634 & w28621);
assign w5034 = (w1634 & w38957) | (w1634 & w38958) | (w38957 & w38958);
assign w5035 = (~w1634 & w38959) | (~w1634 & w38960) | (w38959 & w38960);
assign w5036 = ~w5033 & ~w5034;
assign w5037 = ~w5035 & ~w5036;
assign w5038 = w5027 & ~w5037;
assign w5039 = w5027 & ~w5038;
assign w5040 = ~w5027 & ~w5037;
assign w5041 = ~w5039 & ~w5040;
assign w5042 = ~w4812 & ~w4818;
assign w5043 = w5041 & w5042;
assign w5044 = ~w5041 & ~w5042;
assign w5045 = ~w5043 & ~w5044;
assign w5046 = b_24 & w986;
assign w5047 = w1069 & w28622;
assign w5048 = b_23 & w981;
assign w5049 = ~w5047 & ~w5048;
assign w5050 = ~w5046 & w5049;
assign w5051 = (w5050 & ~w2083) | (w5050 & w28623) | (~w2083 & w28623);
assign w5052 = (w2083 & w38961) | (w2083 & w38962) | (w38961 & w38962);
assign w5053 = (~w2083 & w38963) | (~w2083 & w38964) | (w38963 & w38964);
assign w5054 = ~w5051 & ~w5052;
assign w5055 = ~w5053 & ~w5054;
assign w5056 = ~w5045 & w5055;
assign w5057 = w5045 & ~w5055;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = ~w4834 & w5058;
assign w5060 = w4834 & ~w5058;
assign w5061 = ~w5059 & ~w5060;
assign w5062 = ~w4917 & w5061;
assign w5063 = w5061 & ~w5062;
assign w5064 = ~w5061 & ~w4917;
assign w5065 = ~w5063 & ~w5064;
assign w5066 = ~w4907 & w5065;
assign w5067 = w4907 & ~w5065;
assign w5068 = ~w5066 & ~w5067;
assign w5069 = b_30 & w418;
assign w5070 = w481 & w28624;
assign w5071 = b_29 & w413;
assign w5072 = ~w5070 & ~w5071;
assign w5073 = ~w5069 & w5072;
assign w5074 = (w5073 & ~w3138) | (w5073 & w28625) | (~w3138 & w28625);
assign w5075 = (w3138 & w38965) | (w3138 & w38966) | (w38965 & w38966);
assign w5076 = (~w3138 & w38967) | (~w3138 & w38968) | (w38967 & w38968);
assign w5077 = ~w5074 & ~w5075;
assign w5078 = ~w5076 & ~w5077;
assign w5079 = ~w5068 & ~w5078;
assign w5080 = w5068 & w5078;
assign w5081 = ~w5079 & ~w5080;
assign w5082 = ~w4906 & w5081;
assign w5083 = w4906 & ~w5081;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = ~w4905 & w5084;
assign w5086 = w4905 & w5084;
assign w5087 = ~w5084 & ~w4905;
assign w5088 = ~w5086 & ~w5087;
assign w5089 = ~w4895 & w5088;
assign w5090 = w4895 & ~w5088;
assign w5091 = ~w5089 & ~w5090;
assign w5092 = b_36 & w99;
assign w5093 = w136 & w28626;
assign w5094 = b_35 & w94;
assign w5095 = ~w5093 & ~w5094;
assign w5096 = ~w5092 & w5095;
assign w5097 = (w5096 & ~w4395) | (w5096 & w28627) | (~w4395 & w28627);
assign w5098 = (w4395 & w38969) | (w4395 & w38970) | (w38969 & w38970);
assign w5099 = (~w4395 & w38971) | (~w4395 & w38972) | (w38971 & w38972);
assign w5100 = ~w5097 & ~w5098;
assign w5101 = ~w5099 & ~w5100;
assign w5102 = w5091 & w5101;
assign w5103 = ~w5091 & ~w5101;
assign w5104 = ~w5102 & ~w5103;
assign w5105 = (w5104 & w4867) | (w5104 & w25039) | (w4867 & w25039);
assign w5106 = w4894 & ~w5104;
assign w5107 = ~w5105 & ~w5106;
assign w5108 = ~w5105 & w38973;
assign w5109 = w5107 & ~w5108;
assign w5110 = (~w4893 & w5105) | (~w4893 & w38974) | (w5105 & w38974);
assign w5111 = ~w5109 & ~w5110;
assign w5112 = ~w4870 & ~w4875;
assign w5113 = ~w5111 & ~w5112;
assign w5114 = w5111 & w5112;
assign w5115 = ~w5113 & ~w5114;
assign w5116 = (~w5108 & w5112) | (~w5108 & w38975) | (w5112 & w38975);
assign w5117 = (~w25039 & w28628) | (~w25039 & w28629) | (w28628 & w28629);
assign w5118 = b_37 & w99;
assign w5119 = w136 & w28630;
assign w5120 = b_36 & w94;
assign w5121 = ~w5119 & ~w5120;
assign w5122 = ~w5118 & w5121;
assign w5123 = (w5122 & ~w4636) | (w5122 & w28631) | (~w4636 & w28631);
assign w5124 = (w4636 & w38976) | (w4636 & w38977) | (w38976 & w38977);
assign w5125 = (~w4636 & w38978) | (~w4636 & w38979) | (w38978 & w38979);
assign w5126 = ~w5123 & ~w5124;
assign w5127 = ~w5125 & ~w5126;
assign w5128 = (~w5085 & w4895) | (~w5085 & w28632) | (w4895 & w28632);
assign w5129 = b_34 & w239;
assign w5130 = w266 & w28633;
assign w5131 = b_33 & w234;
assign w5132 = ~w5130 & ~w5131;
assign w5133 = ~w5129 & w5132;
assign w5134 = (w5133 & ~w3967) | (w5133 & w28634) | (~w3967 & w28634);
assign w5135 = (w3967 & w38980) | (w3967 & w38981) | (w38980 & w38981);
assign w5136 = (~w3967 & w38982) | (~w3967 & w38983) | (w38982 & w38983);
assign w5137 = ~w5134 & ~w5135;
assign w5138 = ~w5136 & ~w5137;
assign w5139 = (~w5079 & w4906) | (~w5079 & w27410) | (w4906 & w27410);
assign w5140 = ~w4907 & ~w5065;
assign w5141 = ~w5062 & ~w5140;
assign w5142 = b_28 & w657;
assign w5143 = w754 & w28635;
assign w5144 = b_27 & w652;
assign w5145 = ~w5143 & ~w5144;
assign w5146 = ~w5142 & w5145;
assign w5147 = (w5146 & ~w2771) | (w5146 & w28636) | (~w2771 & w28636);
assign w5148 = (w2771 & w38984) | (w2771 & w38985) | (w38984 & w38985);
assign w5149 = (~w2771 & w38986) | (~w2771 & w38987) | (w38986 & w38987);
assign w5150 = ~w5147 & ~w5148;
assign w5151 = ~w5149 & ~w5150;
assign w5152 = b_16 & w2158;
assign w5153 = w2294 & w28637;
assign w5154 = b_15 & w2153;
assign w5155 = ~w5153 & ~w5154;
assign w5156 = ~w5152 & w5155;
assign w5157 = (w5156 & ~w926) | (w5156 & w28638) | (~w926 & w28638);
assign w5158 = (w926 & w38988) | (w926 & w38989) | (w38988 & w38989);
assign w5159 = (~w926 & w38990) | (~w926 & w38991) | (w38990 & w38991);
assign w5160 = ~w5157 & ~w5158;
assign w5161 = ~w5159 & ~w5160;
assign w5162 = ~w4999 & ~w5002;
assign w5163 = (~w4980 & w4983) | (~w4980 & w26902) | (w4983 & w26902);
assign w5164 = b_7 & w3803;
assign w5165 = w4027 & w28639;
assign w5166 = b_6 & w3798;
assign w5167 = ~w5165 & ~w5166;
assign w5168 = ~w5164 & w5167;
assign w5169 = (w5168 & ~w213) | (w5168 & w28640) | (~w213 & w28640);
assign w5170 = (w213 & w38992) | (w213 & w38993) | (w38992 & w38993);
assign w5171 = (~w213 & w38994) | (~w213 & w38995) | (w38994 & w38995);
assign w5172 = ~w5169 & ~w5170;
assign w5173 = ~w5171 & ~w5172;
assign w5174 = ~w4733 & w28641;
assign w5175 = (~w5174 & w4946) | (~w5174 & w28642) | (w4946 & w28642);
assign w5176 = b_4 & w4499;
assign w5177 = w4723 & w26142;
assign w5178 = b_3 & w4494;
assign w5179 = ~w5177 & ~w5178;
assign w5180 = ~w5176 & w5179;
assign w5181 = w84 & w4502;
assign w5182 = w5180 & ~w5181;
assign w5183 = (a_38 & w5181) | (a_38 & w26143) | (w5181 & w26143);
assign w5184 = ~w5181 & w26549;
assign w5185 = ~w5182 & ~w5183;
assign w5186 = ~w5184 & ~w5185;
assign w5187 = (a_41 & w4942) | (a_41 & w28643) | (w4942 & w28643);
assign w5188 = ~a_39 & a_40;
assign w5189 = a_39 & ~a_40;
assign w5190 = ~w5188 & ~w5189;
assign w5191 = w4942 & ~w5190;
assign w5192 = b_0 & w5191;
assign w5193 = ~a_40 & a_41;
assign w5194 = a_40 & ~a_41;
assign w5195 = ~w5193 & ~w5194;
assign w5196 = ~w4942 & w5195;
assign w5197 = b_1 & w5196;
assign w5198 = ~w5192 & ~w5197;
assign w5199 = ~w4942 & ~w5195;
assign w5200 = ~w15 & w5199;
assign w5201 = w5198 & ~w5200;
assign w5202 = (a_41 & ~w5198) | (a_41 & w25549) | (~w5198 & w25549);
assign w5203 = w5198 & w25797;
assign w5204 = ~w5201 & ~w5202;
assign w5205 = (w5187 & w5204) | (w5187 & w25798) | (w5204 & w25798);
assign w5206 = ~w5204 & w26550;
assign w5207 = ~w5205 & ~w5206;
assign w5208 = w5186 & ~w5207;
assign w5209 = ~w5186 & w5207;
assign w5210 = ~w5208 & ~w5209;
assign w5211 = ~w5175 & w5210;
assign w5212 = w5175 & ~w5210;
assign w5213 = ~w5211 & ~w5212;
assign w5214 = ~w5173 & w5213;
assign w5215 = w5213 & ~w5214;
assign w5216 = ~w5213 & ~w5173;
assign w5217 = ~w5215 & ~w5216;
assign w5218 = ~w4961 & ~w4968;
assign w5219 = w5217 & w5218;
assign w5220 = ~w5217 & ~w5218;
assign w5221 = ~w5219 & ~w5220;
assign w5222 = b_10 & w3195;
assign w5223 = w3388 & w28644;
assign w5224 = b_9 & w3190;
assign w5225 = ~w5223 & ~w5224;
assign w5226 = ~w5222 & w5225;
assign w5227 = (w5226 & ~w454) | (w5226 & w28645) | (~w454 & w28645);
assign w5228 = (w454 & w38996) | (w454 & w38997) | (w38996 & w38997);
assign w5229 = (~w454 & w38998) | (~w454 & w38999) | (w38998 & w38999);
assign w5230 = ~w5227 & ~w5228;
assign w5231 = ~w5229 & ~w5230;
assign w5232 = w5221 & ~w5231;
assign w5233 = ~w5221 & w5231;
assign w5234 = ~w5163 & w27031;
assign w5235 = ~w5163 & ~w5234;
assign w5236 = ~w5232 & ~w5234;
assign w5237 = ~w5234 & w27031;
assign w5238 = ~w5235 & ~w5237;
assign w5239 = b_13 & w2639;
assign w5240 = w2820 & w28646;
assign w5241 = b_12 & w2634;
assign w5242 = ~w5240 & ~w5241;
assign w5243 = ~w5239 & w5242;
assign w5244 = (w5243 & ~w711) | (w5243 & w28647) | (~w711 & w28647);
assign w5245 = (w711 & w39000) | (w711 & w39001) | (w39000 & w39001);
assign w5246 = (~w711 & w39002) | (~w711 & w39003) | (w39002 & w39003);
assign w5247 = ~w5244 & ~w5245;
assign w5248 = ~w5246 & ~w5247;
assign w5249 = w5238 & w5248;
assign w5250 = ~w5238 & ~w5248;
assign w5251 = ~w5249 & ~w5250;
assign w5252 = ~w5162 & w5251;
assign w5253 = w5162 & ~w5251;
assign w5254 = ~w5252 & ~w5253;
assign w5255 = ~w5161 & w5254;
assign w5256 = w5254 & ~w5255;
assign w5257 = ~w5254 & ~w5161;
assign w5258 = ~w5256 & ~w5257;
assign w5259 = (~w5005 & w5008) | (~w5005 & w28648) | (w5008 & w28648);
assign w5260 = w5258 & w5259;
assign w5261 = ~w5258 & ~w5259;
assign w5262 = ~w5260 & ~w5261;
assign w5263 = b_19 & w1694;
assign w5264 = w1834 & w28649;
assign w5265 = b_18 & w1689;
assign w5266 = ~w5264 & ~w5265;
assign w5267 = ~w5263 & w5266;
assign w5268 = (w5267 & ~w1372) | (w5267 & w28650) | (~w1372 & w28650);
assign w5269 = (w1372 & w39004) | (w1372 & w39005) | (w39004 & w39005);
assign w5270 = (~w1372 & w39006) | (~w1372 & w39007) | (w39006 & w39007);
assign w5271 = ~w5268 & ~w5269;
assign w5272 = ~w5270 & ~w5271;
assign w5273 = w5262 & ~w5272;
assign w5274 = w5262 & ~w5273;
assign w5275 = ~w5262 & ~w5272;
assign w5276 = ~w5274 & ~w5275;
assign w5277 = (~w5022 & w4918) | (~w5022 & w27211) | (w4918 & w27211);
assign w5278 = w5276 & w5277;
assign w5279 = ~w5276 & ~w5277;
assign w5280 = ~w5278 & ~w5279;
assign w5281 = b_22 & w1295;
assign w5282 = w1422 & w28651;
assign w5283 = b_21 & w1290;
assign w5284 = ~w5282 & ~w5283;
assign w5285 = ~w5281 & w5284;
assign w5286 = (w5285 & ~w1786) | (w5285 & w28652) | (~w1786 & w28652);
assign w5287 = (w1786 & w39008) | (w1786 & w39009) | (w39008 & w39009);
assign w5288 = (~w1786 & w39010) | (~w1786 & w39011) | (w39010 & w39011);
assign w5289 = ~w5286 & ~w5287;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = w5280 & ~w5290;
assign w5292 = w5280 & ~w5291;
assign w5293 = ~w5280 & ~w5290;
assign w5294 = ~w5292 & ~w5293;
assign w5295 = (~w5038 & w5042) | (~w5038 & w27139) | (w5042 & w27139);
assign w5296 = w5294 & w5295;
assign w5297 = ~w5294 & ~w5295;
assign w5298 = ~w5296 & ~w5297;
assign w5299 = b_25 & w986;
assign w5300 = w1069 & w28653;
assign w5301 = b_24 & w981;
assign w5302 = ~w5300 & ~w5301;
assign w5303 = ~w5299 & w5302;
assign w5304 = (w5303 & ~w2108) | (w5303 & w28654) | (~w2108 & w28654);
assign w5305 = (w2108 & w39012) | (w2108 & w39013) | (w39012 & w39013);
assign w5306 = (~w2108 & w39014) | (~w2108 & w39015) | (w39014 & w39015);
assign w5307 = ~w5304 & ~w5305;
assign w5308 = ~w5306 & ~w5307;
assign w5309 = w5298 & ~w5308;
assign w5310 = w5298 & ~w5309;
assign w5311 = ~w5298 & ~w5308;
assign w5312 = ~w5310 & ~w5311;
assign w5313 = ~w5057 & ~w5059;
assign w5314 = ~w5312 & ~w5313;
assign w5315 = w5312 & w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = ~w5151 & w5316;
assign w5318 = ~w5316 & ~w5151;
assign w5319 = w5316 & ~w5317;
assign w5320 = ~w5318 & ~w5319;
assign w5321 = ~w5141 & ~w5320;
assign w5322 = w5320 & ~w5141;
assign w5323 = ~w5320 & ~w5321;
assign w5324 = b_31 & w418;
assign w5325 = w481 & w28655;
assign w5326 = b_30 & w413;
assign w5327 = ~w5325 & ~w5326;
assign w5328 = ~w5324 & w5327;
assign w5329 = (w5328 & ~w3345) | (w5328 & w28656) | (~w3345 & w28656);
assign w5330 = (w3345 & w39016) | (w3345 & w39017) | (w39016 & w39017);
assign w5331 = (~w3345 & w39018) | (~w3345 & w39019) | (w39018 & w39019);
assign w5332 = ~w5329 & ~w5330;
assign w5333 = ~w5331 & ~w5332;
assign w5334 = ~w5323 & w39020;
assign w5335 = (~w5333 & w5323) | (~w5333 & w39021) | (w5323 & w39021);
assign w5336 = ~w5334 & ~w5335;
assign w5337 = ~w5139 & w5336;
assign w5338 = w5139 & ~w5336;
assign w5339 = ~w5337 & ~w5338;
assign w5340 = w5138 & ~w5339;
assign w5341 = ~w5138 & w5339;
assign w5342 = ~w5340 & ~w5341;
assign w5343 = ~w5128 & w5342;
assign w5344 = w5128 & ~w5342;
assign w5345 = ~w5343 & ~w5344;
assign w5346 = ~w5127 & w5345;
assign w5347 = w5345 & ~w5346;
assign w5348 = ~w5345 & ~w5127;
assign w5349 = ~w5347 & ~w5348;
assign w5350 = ~w5117 & w5349;
assign w5351 = w5117 & ~w5349;
assign w5352 = ~w5350 & ~w5351;
assign w5353 = w8 & w28657;
assign w5354 = ~w8 & w28658;
assign w5355 = b_39 & w4;
assign w5356 = ~w5354 & ~w5355;
assign w5357 = ~w5353 & w5356;
assign w5358 = ~b_39 & ~b_40;
assign w5359 = b_39 & b_40;
assign w5360 = ~w5358 & ~w5359;
assign w5361 = (w4656 & w28661) | (w4656 & w28662) | (w28661 & w28662);
assign w5362 = (~w4656 & w28663) | (~w4656 & w28664) | (w28663 & w28664);
assign w5363 = ~w5361 & ~w5362;
assign w5364 = (w5357 & ~w5363) | (w5357 & w28665) | (~w5363 & w28665);
assign w5365 = (w5363 & w39022) | (w5363 & w39023) | (w39022 & w39023);
assign w5366 = (~w5363 & w39024) | (~w5363 & w39025) | (w39024 & w39025);
assign w5367 = ~w5364 & ~w5365;
assign w5368 = ~w5366 & ~w5367;
assign w5369 = ~w5352 & ~w5368;
assign w5370 = w5352 & w5368;
assign w5371 = ~w5369 & ~w5370;
assign w5372 = ~w5116 & w5371;
assign w5373 = w5116 & ~w5371;
assign w5374 = ~w5372 & ~w5373;
assign w5375 = (~w5369 & w5116) | (~w5369 & w28666) | (w5116 & w28666);
assign w5376 = ~w5117 & ~w5349;
assign w5377 = (~w5346 & w5349) | (~w5346 & w28667) | (w5349 & w28667);
assign w5378 = (~w5341 & ~w5342) | (~w5341 & w28668) | (~w5342 & w28668);
assign w5379 = b_35 & w239;
assign w5380 = w266 & w28669;
assign w5381 = b_34 & w234;
assign w5382 = ~w5380 & ~w5381;
assign w5383 = ~w5379 & w5382;
assign w5384 = (w5383 & ~w4181) | (w5383 & w25040) | (~w4181 & w25040);
assign w5385 = (w4181 & w28670) | (w4181 & w28671) | (w28670 & w28671);
assign w5386 = (~w4181 & w28672) | (~w4181 & w28673) | (w28672 & w28673);
assign w5387 = ~w5384 & ~w5385;
assign w5388 = ~w5386 & ~w5387;
assign w5389 = (~w5335 & ~w5336) | (~w5335 & w27411) | (~w5336 & w27411);
assign w5390 = b_32 & w418;
assign w5391 = w481 & w28674;
assign w5392 = b_31 & w413;
assign w5393 = ~w5391 & ~w5392;
assign w5394 = ~w5390 & w5393;
assign w5395 = (w5394 & ~w3545) | (w5394 & w25041) | (~w3545 & w25041);
assign w5396 = (w3545 & w28675) | (w3545 & w28676) | (w28675 & w28676);
assign w5397 = (~w3545 & w28677) | (~w3545 & w28678) | (w28677 & w28678);
assign w5398 = ~w5395 & ~w5396;
assign w5399 = ~w5397 & ~w5398;
assign w5400 = (~w5317 & w5320) | (~w5317 & w39026) | (w5320 & w39026);
assign w5401 = b_29 & w657;
assign w5402 = w754 & w28679;
assign w5403 = b_28 & w652;
assign w5404 = ~w5402 & ~w5403;
assign w5405 = ~w5401 & w5404;
assign w5406 = (w5405 & ~w2954) | (w5405 & w28680) | (~w2954 & w28680);
assign w5407 = (w2954 & w39027) | (w2954 & w39028) | (w39027 & w39028);
assign w5408 = (~w2954 & w39029) | (~w2954 & w39030) | (w39029 & w39030);
assign w5409 = ~w5406 & ~w5407;
assign w5410 = ~w5408 & ~w5409;
assign w5411 = (~w5309 & w5312) | (~w5309 & w39031) | (w5312 & w39031);
assign w5412 = (~w5291 & w5294) | (~w5291 & w39032) | (w5294 & w39032);
assign w5413 = b_20 & w1694;
assign w5414 = w1834 & w28681;
assign w5415 = b_19 & w1689;
assign w5416 = ~w5414 & ~w5415;
assign w5417 = ~w5413 & w5416;
assign w5418 = (w5417 & ~w1503) | (w5417 & w28682) | (~w1503 & w28682);
assign w5419 = (w1503 & w39033) | (w1503 & w39034) | (w39033 & w39034);
assign w5420 = (~w1503 & w39035) | (~w1503 & w39036) | (w39035 & w39036);
assign w5421 = ~w5418 & ~w5419;
assign w5422 = ~w5420 & ~w5421;
assign w5423 = (~w5255 & w5258) | (~w5255 & w28683) | (w5258 & w28683);
assign w5424 = b_17 & w2158;
assign w5425 = w2294 & w28684;
assign w5426 = b_16 & w2153;
assign w5427 = ~w5425 & ~w5426;
assign w5428 = ~w5424 & w5427;
assign w5429 = (w5428 & ~w1038) | (w5428 & w28685) | (~w1038 & w28685);
assign w5430 = (w1038 & w39037) | (w1038 & w39038) | (w39037 & w39038);
assign w5431 = (~w1038 & w39039) | (~w1038 & w39040) | (w39039 & w39040);
assign w5432 = ~w5429 & ~w5430;
assign w5433 = ~w5431 & ~w5432;
assign w5434 = ~w5250 & ~w5252;
assign w5435 = b_14 & w2639;
assign w5436 = w2820 & w28686;
assign w5437 = b_13 & w2634;
assign w5438 = ~w5436 & ~w5437;
assign w5439 = ~w5435 & w5438;
assign w5440 = (w5439 & ~w735) | (w5439 & w28687) | (~w735 & w28687);
assign w5441 = (w735 & w39041) | (w735 & w39042) | (w39041 & w39042);
assign w5442 = (~w735 & w39043) | (~w735 & w39044) | (w39043 & w39044);
assign w5443 = ~w5440 & ~w5441;
assign w5444 = ~w5442 & ~w5443;
assign w5445 = (~w5214 & w5218) | (~w5214 & w28688) | (w5218 & w28688);
assign w5446 = b_8 & w3803;
assign w5447 = w4027 & w28689;
assign w5448 = b_7 & w3798;
assign w5449 = ~w5447 & ~w5448;
assign w5450 = ~w5446 & w5449;
assign w5451 = ~w308 & w28690;
assign w5452 = (w5450 & ~w28690) | (w5450 & w39045) | (~w28690 & w39045);
assign w5453 = (w28690 & w39046) | (w28690 & w39047) | (w39046 & w39047);
assign w5454 = ~w5451 & w28692;
assign w5455 = ~w5452 & ~w5453;
assign w5456 = ~w5454 & ~w5455;
assign w5457 = (~w5209 & w5175) | (~w5209 & w26144) | (w5175 & w26144);
assign w5458 = b_2 & w5196;
assign w5459 = w4942 & ~w5195;
assign w5460 = w5459 & w25370;
assign w5461 = b_1 & w5191;
assign w5462 = ~w5460 & ~w5461;
assign w5463 = ~w5458 & w5462;
assign w5464 = w35 & w5199;
assign w5465 = w5463 & ~w5464;
assign w5466 = (a_41 & ~w5463) | (a_41 & w25550) | (~w5463 & w25550);
assign w5467 = w5463 & w25799;
assign w5468 = ~w5465 & ~w5466;
assign w5469 = ~w5467 & ~w5468;
assign w5470 = ~w5205 & w5469;
assign w5471 = w5205 & ~w5469;
assign w5472 = ~w5470 & ~w5471;
assign w5473 = b_5 & w4499;
assign w5474 = w4723 & w26551;
assign w5475 = b_4 & w4494;
assign w5476 = ~w5474 & ~w5475;
assign w5477 = ~w5473 & w5476;
assign w5478 = w129 & w4502;
assign w5479 = w5477 & ~w5478;
assign w5480 = (a_38 & w5478) | (a_38 & w26552) | (w5478 & w26552);
assign w5481 = ~w5478 & w39048;
assign w5482 = ~w5479 & ~w5480;
assign w5483 = ~w5481 & ~w5482;
assign w5484 = w5472 & ~w5483;
assign w5485 = w5472 & ~w5484;
assign w5486 = ~w5472 & ~w5483;
assign w5487 = ~w5485 & ~w5486;
assign w5488 = ~w5457 & ~w5487;
assign w5489 = w5457 & w5487;
assign w5490 = ~w5488 & ~w5489;
assign w5491 = ~w5456 & w5490;
assign w5492 = ~w5490 & ~w5456;
assign w5493 = w5490 & ~w5491;
assign w5494 = ~w5492 & ~w5493;
assign w5495 = ~w5445 & ~w5494;
assign w5496 = ~w5445 & ~w5495;
assign w5497 = b_11 & w3195;
assign w5498 = w3388 & w28693;
assign w5499 = b_10 & w3190;
assign w5500 = ~w5498 & ~w5499;
assign w5501 = ~w5497 & w5500;
assign w5502 = (w5501 & ~w530) | (w5501 & w28694) | (~w530 & w28694);
assign w5503 = (w530 & w39049) | (w530 & w39050) | (w39049 & w39050);
assign w5504 = (~w530 & w39051) | (~w530 & w39052) | (w39051 & w39052);
assign w5505 = ~w5502 & ~w5503;
assign w5506 = ~w5504 & ~w5505;
assign w5507 = ~w5496 & w27032;
assign w5508 = (~w5506 & w5496) | (~w5506 & w27033) | (w5496 & w27033);
assign w5509 = ~w5507 & ~w5508;
assign w5510 = ~w5236 & w5509;
assign w5511 = w5236 & ~w5509;
assign w5512 = ~w5510 & ~w5511;
assign w5513 = w5444 & ~w5512;
assign w5514 = ~w5444 & w5512;
assign w5515 = ~w5513 & ~w5514;
assign w5516 = ~w5434 & w5515;
assign w5517 = w5434 & ~w5515;
assign w5518 = ~w5516 & ~w5517;
assign w5519 = w5433 & ~w5518;
assign w5520 = ~w5433 & w5518;
assign w5521 = ~w5519 & ~w5520;
assign w5522 = ~w5423 & w5521;
assign w5523 = w5423 & ~w5521;
assign w5524 = ~w5522 & ~w5523;
assign w5525 = ~w5422 & w5524;
assign w5526 = w5524 & ~w5525;
assign w5527 = ~w5524 & ~w5422;
assign w5528 = ~w5526 & ~w5527;
assign w5529 = (~w5273 & w5276) | (~w5273 & w27212) | (w5276 & w27212);
assign w5530 = w5528 & w5529;
assign w5531 = ~w5528 & ~w5529;
assign w5532 = ~w5530 & ~w5531;
assign w5533 = b_23 & w1295;
assign w5534 = w1422 & w28695;
assign w5535 = b_22 & w1290;
assign w5536 = ~w5534 & ~w5535;
assign w5537 = ~w5533 & w5536;
assign w5538 = (w5537 & ~w1933) | (w5537 & w28696) | (~w1933 & w28696);
assign w5539 = (w1933 & w39053) | (w1933 & w39054) | (w39053 & w39054);
assign w5540 = (~w1933 & w39055) | (~w1933 & w39056) | (w39055 & w39056);
assign w5541 = ~w5538 & ~w5539;
assign w5542 = ~w5540 & ~w5541;
assign w5543 = w5532 & ~w5542;
assign w5544 = ~w5532 & w5542;
assign w5545 = (w5297 & w27341) | (w5297 & w27342) | (w27341 & w27342);
assign w5546 = ~w5412 & ~w5545;
assign w5547 = (~w5297 & w28697) | (~w5297 & w28698) | (w28697 & w28698);
assign w5548 = ~w5297 & w28699;
assign w5549 = b_26 & w986;
assign w5550 = w1069 & w28700;
assign w5551 = b_25 & w981;
assign w5552 = ~w5550 & ~w5551;
assign w5553 = ~w5549 & w5552;
assign w5554 = (w5553 & ~w2416) | (w5553 & w28701) | (~w2416 & w28701);
assign w5555 = (w2416 & w39057) | (w2416 & w39058) | (w39057 & w39058);
assign w5556 = (~w2416 & w39059) | (~w2416 & w39060) | (w39059 & w39060);
assign w5557 = ~w5554 & ~w5555;
assign w5558 = ~w5556 & ~w5557;
assign w5559 = ~w5546 & w28702;
assign w5560 = (~w5558 & w5546) | (~w5558 & w28703) | (w5546 & w28703);
assign w5561 = ~w5559 & ~w5560;
assign w5562 = (w5561 & w5314) | (w5561 & w28704) | (w5314 & w28704);
assign w5563 = ~w5314 & w28705;
assign w5564 = ~w5562 & ~w5563;
assign w5565 = w5410 & ~w5564;
assign w5566 = ~w5410 & w5564;
assign w5567 = ~w5565 & ~w5566;
assign w5568 = (w5567 & w5321) | (w5567 & w28706) | (w5321 & w28706);
assign w5569 = ~w5321 & w28707;
assign w5570 = ~w5568 & ~w5569;
assign w5571 = w5399 & ~w5570;
assign w5572 = ~w5399 & w5570;
assign w5573 = ~w5571 & ~w5572;
assign w5574 = ~w5389 & w5573;
assign w5575 = w5389 & ~w5573;
assign w5576 = ~w5574 & ~w5575;
assign w5577 = ~w5388 & w5576;
assign w5578 = w5576 & ~w5577;
assign w5579 = ~w5576 & ~w5388;
assign w5580 = ~w5578 & ~w5579;
assign w5581 = ~w5378 & w5580;
assign w5582 = w5378 & ~w5580;
assign w5583 = ~w5581 & ~w5582;
assign w5584 = b_38 & w99;
assign w5585 = w136 & w28708;
assign w5586 = b_37 & w94;
assign w5587 = ~w5585 & ~w5586;
assign w5588 = ~w5584 & w5587;
assign w5589 = (w5588 & ~w4658) | (w5588 & w28709) | (~w4658 & w28709);
assign w5590 = (w4658 & w39061) | (w4658 & w39062) | (w39061 & w39062);
assign w5591 = (~w4658 & w39063) | (~w4658 & w39064) | (w39063 & w39064);
assign w5592 = ~w5589 & ~w5590;
assign w5593 = ~w5591 & ~w5592;
assign w5594 = ~w5583 & ~w5593;
assign w5595 = w5583 & w5593;
assign w5596 = ~w5594 & ~w5595;
assign w5597 = w5377 & ~w5596;
assign w5598 = (w5596 & w5376) | (w5596 & w25042) | (w5376 & w25042);
assign w5599 = w8 & w28710;
assign w5600 = ~w8 & w28711;
assign w5601 = b_40 & w4;
assign w5602 = ~w5600 & ~w5601;
assign w5603 = ~w5599 & w5602;
assign w5604 = ~b_40 & ~b_41;
assign w5605 = b_40 & b_41;
assign w5606 = ~w5604 & ~w5605;
assign w5607 = (w4656 & w28714) | (w4656 & w28715) | (w28714 & w28715);
assign w5608 = (~w4656 & w28716) | (~w4656 & w28717) | (w28716 & w28717);
assign w5609 = ~w5607 & ~w5608;
assign w5610 = (w5603 & ~w5609) | (w5603 & w28718) | (~w5609 & w28718);
assign w5611 = (w5609 & w39065) | (w5609 & w39066) | (w39065 & w39066);
assign w5612 = (~w5609 & w39067) | (~w5609 & w39068) | (w39067 & w39068);
assign w5613 = ~w5610 & ~w5611;
assign w5614 = ~w5612 & ~w5613;
assign w5615 = (w5614 & w5598) | (w5614 & w28719) | (w5598 & w28719);
assign w5616 = ~w5598 & w28720;
assign w5617 = ~w5615 & ~w5616;
assign w5618 = (w5617 & w5372) | (w5617 & w25043) | (w5372 & w25043);
assign w5619 = w5375 & ~w5617;
assign w5620 = ~w5618 & ~w5619;
assign w5621 = (~w25042 & w28721) | (~w25042 & w28722) | (w28721 & w28722);
assign w5622 = b_39 & w99;
assign w5623 = w136 & w28723;
assign w5624 = b_38 & w94;
assign w5625 = ~w5623 & ~w5624;
assign w5626 = ~w5622 & w5625;
assign w5627 = (w5626 & ~w4888) | (w5626 & w28724) | (~w4888 & w28724);
assign w5628 = (w4888 & w39069) | (w4888 & w39070) | (w39069 & w39070);
assign w5629 = (~w4888 & w39071) | (~w4888 & w39072) | (w39071 & w39072);
assign w5630 = ~w5627 & ~w5628;
assign w5631 = ~w5629 & ~w5630;
assign w5632 = (~w5577 & w5580) | (~w5577 & w28725) | (w5580 & w28725);
assign w5633 = ~w5572 & ~w5574;
assign w5634 = b_33 & w418;
assign w5635 = w481 & w28726;
assign w5636 = b_32 & w413;
assign w5637 = ~w5635 & ~w5636;
assign w5638 = ~w5634 & w5637;
assign w5639 = (w5638 & ~w3744) | (w5638 & w25044) | (~w3744 & w25044);
assign w5640 = (w3744 & w28727) | (w3744 & w28728) | (w28727 & w28728);
assign w5641 = (~w3744 & w28729) | (~w3744 & w28730) | (w28729 & w28730);
assign w5642 = ~w5639 & ~w5640;
assign w5643 = ~w5641 & ~w5642;
assign w5644 = (~w5566 & w5400) | (~w5566 & w27412) | (w5400 & w27412);
assign w5645 = (~w5560 & w5411) | (~w5560 & w27413) | (w5411 & w27413);
assign w5646 = b_27 & w986;
assign w5647 = w1069 & w28731;
assign w5648 = b_26 & w981;
assign w5649 = ~w5647 & ~w5648;
assign w5650 = ~w5646 & w5649;
assign w5651 = (w5650 & ~w2582) | (w5650 & w28732) | (~w2582 & w28732);
assign w5652 = (w2582 & w39073) | (w2582 & w39074) | (w39073 & w39074);
assign w5653 = (~w2582 & w39075) | (~w2582 & w39076) | (w39075 & w39076);
assign w5654 = ~w5651 & ~w5652;
assign w5655 = ~w5653 & ~w5654;
assign w5656 = b_21 & w1694;
assign w5657 = w1834 & w28733;
assign w5658 = b_20 & w1689;
assign w5659 = ~w5657 & ~w5658;
assign w5660 = ~w5656 & w5659;
assign w5661 = (w5660 & ~w1634) | (w5660 & w28734) | (~w1634 & w28734);
assign w5662 = (w1634 & w39077) | (w1634 & w39078) | (w39077 & w39078);
assign w5663 = (~w1634 & w39079) | (~w1634 & w39080) | (w39079 & w39080);
assign w5664 = ~w5661 & ~w5662;
assign w5665 = ~w5663 & ~w5664;
assign w5666 = (~w5520 & w5423) | (~w5520 & w27214) | (w5423 & w27214);
assign w5667 = (~w5514 & w5434) | (~w5514 & w27215) | (w5434 & w27215);
assign w5668 = (~w5508 & w5236) | (~w5508 & w28735) | (w5236 & w28735);
assign w5669 = b_12 & w3195;
assign w5670 = w3388 & w28736;
assign w5671 = b_11 & w3190;
assign w5672 = ~w5670 & ~w5671;
assign w5673 = ~w5669 & w5672;
assign w5674 = (w5673 & ~w552) | (w5673 & w28737) | (~w552 & w28737);
assign w5675 = (w552 & w39081) | (w552 & w39082) | (w39081 & w39082);
assign w5676 = (~w552 & w39083) | (~w552 & w39084) | (w39083 & w39084);
assign w5677 = ~w5674 & ~w5675;
assign w5678 = ~w5676 & ~w5677;
assign w5679 = (~w5491 & w5445) | (~w5491 & w26553) | (w5445 & w26553);
assign w5680 = b_6 & w4499;
assign w5681 = w4723 & w28738;
assign w5682 = b_5 & w4494;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = ~w5680 & w5683;
assign w5685 = (w5684 & ~w190) | (w5684 & w28739) | (~w190 & w28739);
assign w5686 = (w190 & w39085) | (w190 & w39086) | (w39085 & w39086);
assign w5687 = (~w190 & w39087) | (~w190 & w39088) | (w39087 & w39088);
assign w5688 = ~w5685 & ~w5686;
assign w5689 = ~w5687 & ~w5688;
assign w5690 = a_41 & ~a_42;
assign w5691 = ~a_41 & a_42;
assign w5692 = ~w5690 & ~w5691;
assign w5693 = b_0 & ~w5692;
assign w5694 = (w5693 & w5469) | (w5693 & w25800) | (w5469 & w25800);
assign w5695 = ~w5469 & w25801;
assign w5696 = ~w5694 & ~w5695;
assign w5697 = b_3 & w5196;
assign w5698 = w5459 & w26145;
assign w5699 = b_2 & w5191;
assign w5700 = ~w5698 & ~w5699;
assign w5701 = ~w5697 & w5700;
assign w5702 = w57 & w5199;
assign w5703 = w5701 & ~w5702;
assign w5704 = a_41 & ~w5703;
assign w5705 = w5703 & a_41;
assign w5706 = ~w5703 & ~w5704;
assign w5707 = ~w5705 & ~w5706;
assign w5708 = ~w5696 & ~w5707;
assign w5709 = w5696 & w5707;
assign w5710 = ~w5708 & ~w5709;
assign w5711 = ~w5689 & w5710;
assign w5712 = w5710 & ~w5711;
assign w5713 = ~w5710 & ~w5689;
assign w5714 = ~w5712 & ~w5713;
assign w5715 = ~w5484 & ~w5488;
assign w5716 = w5714 & w5715;
assign w5717 = ~w5714 & ~w5715;
assign w5718 = ~w5716 & ~w5717;
assign w5719 = b_9 & w3803;
assign w5720 = w4027 & w28740;
assign w5721 = b_8 & w3798;
assign w5722 = ~w5720 & ~w5721;
assign w5723 = ~w5719 & w5722;
assign w5724 = (w5723 & ~w371) | (w5723 & w28741) | (~w371 & w28741);
assign w5725 = (w371 & w39089) | (w371 & w39090) | (w39089 & w39090);
assign w5726 = (~w371 & w39091) | (~w371 & w39092) | (w39091 & w39092);
assign w5727 = ~w5724 & ~w5725;
assign w5728 = ~w5726 & ~w5727;
assign w5729 = ~w5718 & w5728;
assign w5730 = w5718 & ~w5728;
assign w5731 = ~w5729 & ~w5730;
assign w5732 = ~w5679 & w5731;
assign w5733 = w5679 & ~w5731;
assign w5734 = ~w5732 & ~w5733;
assign w5735 = ~w5678 & w5734;
assign w5736 = ~w5734 & ~w5678;
assign w5737 = w5734 & ~w5735;
assign w5738 = ~w5736 & ~w5737;
assign w5739 = ~w5668 & ~w5738;
assign w5740 = ~w5668 & ~w5739;
assign w5741 = ~w5738 & ~w5739;
assign w5742 = ~w5740 & ~w5741;
assign w5743 = b_15 & w2639;
assign w5744 = w2820 & w28742;
assign w5745 = b_14 & w2634;
assign w5746 = ~w5744 & ~w5745;
assign w5747 = ~w5743 & w5746;
assign w5748 = (w5747 & ~w827) | (w5747 & w28743) | (~w827 & w28743);
assign w5749 = (w827 & w39093) | (w827 & w39094) | (w39093 & w39094);
assign w5750 = (~w827 & w39095) | (~w827 & w39096) | (w39095 & w39096);
assign w5751 = ~w5748 & ~w5749;
assign w5752 = ~w5750 & ~w5751;
assign w5753 = ~w5742 & ~w5752;
assign w5754 = ~w5742 & ~w5753;
assign w5755 = w5742 & ~w5752;
assign w5756 = ~w5754 & ~w5755;
assign w5757 = ~w5754 & w27216;
assign w5758 = (w5667 & w5754) | (w5667 & w27217) | (w5754 & w27217);
assign w5759 = ~w5757 & ~w5758;
assign w5760 = b_18 & w2158;
assign w5761 = w2294 & w28744;
assign w5762 = b_17 & w2153;
assign w5763 = ~w5761 & ~w5762;
assign w5764 = ~w5760 & w5763;
assign w5765 = (w5764 & ~w1238) | (w5764 & w28745) | (~w1238 & w28745);
assign w5766 = (w1238 & w39097) | (w1238 & w39098) | (w39097 & w39098);
assign w5767 = (~w1238 & w39099) | (~w1238 & w39100) | (w39099 & w39100);
assign w5768 = ~w5765 & ~w5766;
assign w5769 = ~w5767 & ~w5768;
assign w5770 = ~w5759 & ~w5769;
assign w5771 = w5759 & w5769;
assign w5772 = ~w5770 & ~w5771;
assign w5773 = ~w5666 & w5772;
assign w5774 = w5666 & ~w5772;
assign w5775 = ~w5773 & ~w5774;
assign w5776 = ~w5665 & w5775;
assign w5777 = w5775 & ~w5776;
assign w5778 = ~w5775 & ~w5665;
assign w5779 = ~w5777 & ~w5778;
assign w5780 = (~w5525 & w5528) | (~w5525 & w27218) | (w5528 & w27218);
assign w5781 = w5779 & w5780;
assign w5782 = ~w5779 & ~w5780;
assign w5783 = ~w5781 & ~w5782;
assign w5784 = b_24 & w1295;
assign w5785 = w1422 & w28746;
assign w5786 = b_23 & w1290;
assign w5787 = ~w5785 & ~w5786;
assign w5788 = ~w5784 & w5787;
assign w5789 = (w5788 & ~w2083) | (w5788 & w28747) | (~w2083 & w28747);
assign w5790 = (w2083 & w39101) | (w2083 & w39102) | (w39101 & w39102);
assign w5791 = (~w2083 & w39103) | (~w2083 & w39104) | (w39103 & w39104);
assign w5792 = ~w5789 & ~w5790;
assign w5793 = ~w5791 & ~w5792;
assign w5794 = ~w5783 & w5793;
assign w5795 = w5783 & ~w5793;
assign w5796 = ~w5794 & ~w5795;
assign w5797 = ~w5547 & w5796;
assign w5798 = w5547 & ~w5796;
assign w5799 = ~w5797 & ~w5798;
assign w5800 = ~w5655 & w5799;
assign w5801 = w5799 & ~w5800;
assign w5802 = ~w5799 & ~w5655;
assign w5803 = ~w5801 & ~w5802;
assign w5804 = ~w5645 & w5803;
assign w5805 = w5645 & ~w5803;
assign w5806 = ~w5804 & ~w5805;
assign w5807 = b_30 & w657;
assign w5808 = w754 & w28748;
assign w5809 = b_29 & w652;
assign w5810 = ~w5808 & ~w5809;
assign w5811 = ~w5807 & w5810;
assign w5812 = (w5811 & ~w3138) | (w5811 & w28749) | (~w3138 & w28749);
assign w5813 = (w3138 & w39105) | (w3138 & w39106) | (w39105 & w39106);
assign w5814 = (~w3138 & w39107) | (~w3138 & w39108) | (w39107 & w39108);
assign w5815 = ~w5812 & ~w5813;
assign w5816 = ~w5814 & ~w5815;
assign w5817 = ~w5806 & ~w5816;
assign w5818 = w5806 & w5816;
assign w5819 = ~w5817 & ~w5818;
assign w5820 = ~w5644 & w5819;
assign w5821 = w5644 & ~w5819;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = ~w5643 & w5822;
assign w5824 = w5822 & ~w5823;
assign w5825 = ~w5822 & ~w5643;
assign w5826 = ~w5824 & ~w5825;
assign w5827 = ~w5633 & w5826;
assign w5828 = w5633 & ~w5826;
assign w5829 = ~w5827 & ~w5828;
assign w5830 = b_36 & w239;
assign w5831 = w266 & w28750;
assign w5832 = b_35 & w234;
assign w5833 = ~w5831 & ~w5832;
assign w5834 = ~w5830 & w5833;
assign w5835 = (w5834 & ~w4395) | (w5834 & w25045) | (~w4395 & w25045);
assign w5836 = (w4395 & w28751) | (w4395 & w28752) | (w28751 & w28752);
assign w5837 = (~w4395 & w28753) | (~w4395 & w28754) | (w28753 & w28754);
assign w5838 = ~w5835 & ~w5836;
assign w5839 = ~w5837 & ~w5838;
assign w5840 = w5829 & w5839;
assign w5841 = ~w5829 & ~w5839;
assign w5842 = ~w5840 & ~w5841;
assign w5843 = ~w5632 & w5842;
assign w5844 = w5632 & ~w5842;
assign w5845 = ~w5843 & ~w5844;
assign w5846 = ~w5631 & w5845;
assign w5847 = ~w5845 & ~w5631;
assign w5848 = w5845 & ~w5846;
assign w5849 = ~w5847 & ~w5848;
assign w5850 = ~w5621 & ~w5849;
assign w5851 = w5849 & ~w5621;
assign w5852 = ~w5849 & ~w5850;
assign w5853 = ~w5851 & ~w5852;
assign w5854 = w8 & w28755;
assign w5855 = ~w8 & w28756;
assign w5856 = b_41 & w4;
assign w5857 = ~w5855 & ~w5856;
assign w5858 = ~w5854 & w5857;
assign w5859 = ~b_41 & ~b_42;
assign w5860 = b_41 & b_42;
assign w5861 = ~w5859 & ~w5860;
assign w5862 = (w4656 & w28758) | (w4656 & w28759) | (w28758 & w28759);
assign w5863 = (~w4656 & w28760) | (~w4656 & w28761) | (w28760 & w28761);
assign w5864 = ~w5862 & ~w5863;
assign w5865 = (w5858 & ~w5864) | (w5858 & w28762) | (~w5864 & w28762);
assign w5866 = (w5864 & w39109) | (w5864 & w39110) | (w39109 & w39110);
assign w5867 = (~w5864 & w39111) | (~w5864 & w39112) | (w39111 & w39112);
assign w5868 = ~w5865 & ~w5866;
assign w5869 = ~w5867 & ~w5868;
assign w5870 = (~w5869 & w5852) | (~w5869 & w39113) | (w5852 & w39113);
assign w5871 = ~w5853 & ~w5870;
assign w5872 = ~w5852 & w39114;
assign w5873 = ~w5871 & ~w5872;
assign w5874 = (~w25043 & w39115) | (~w25043 & w39116) | (w39115 & w39116);
assign w5875 = ~w5873 & ~w5874;
assign w5876 = w5873 & w5874;
assign w5877 = ~w5875 & ~w5876;
assign w5878 = w8 & w28763;
assign w5879 = ~w8 & w28764;
assign w5880 = b_42 & w4;
assign w5881 = ~w5879 & ~w5880;
assign w5882 = ~w5878 & w5881;
assign w5883 = ~b_42 & ~b_43;
assign w5884 = b_42 & b_43;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = (w4656 & w28766) | (w4656 & w28767) | (w28766 & w28767);
assign w5887 = (~w4656 & w28768) | (~w4656 & w28769) | (w28768 & w28769);
assign w5888 = ~w5886 & ~w5887;
assign w5889 = (w5882 & ~w5888) | (w5882 & w28770) | (~w5888 & w28770);
assign w5890 = (w5888 & w39117) | (w5888 & w39118) | (w39117 & w39118);
assign w5891 = (~w5888 & w39119) | (~w5888 & w39120) | (w39119 & w39120);
assign w5892 = ~w5889 & ~w5890;
assign w5893 = ~w5891 & ~w5892;
assign w5894 = (~w5846 & w5849) | (~w5846 & w39121) | (w5849 & w39121);
assign w5895 = (~w5841 & w5632) | (~w5841 & w25046) | (w5632 & w25046);
assign w5896 = b_34 & w418;
assign w5897 = w481 & w28771;
assign w5898 = b_33 & w413;
assign w5899 = ~w5897 & ~w5898;
assign w5900 = ~w5896 & w5899;
assign w5901 = (w5900 & ~w3967) | (w5900 & w28772) | (~w3967 & w28772);
assign w5902 = (w3967 & w39122) | (w3967 & w39123) | (w39122 & w39123);
assign w5903 = (~w3967 & w39124) | (~w3967 & w39125) | (w39124 & w39125);
assign w5904 = ~w5901 & ~w5902;
assign w5905 = ~w5903 & ~w5904;
assign w5906 = (~w5817 & w5644) | (~w5817 & w27526) | (w5644 & w27526);
assign w5907 = (~w5800 & w5645) | (~w5800 & w28773) | (w5645 & w28773);
assign w5908 = b_28 & w986;
assign w5909 = w1069 & w28774;
assign w5910 = b_27 & w981;
assign w5911 = ~w5909 & ~w5910;
assign w5912 = ~w5908 & w5911;
assign w5913 = (w5912 & ~w2771) | (w5912 & w28775) | (~w2771 & w28775);
assign w5914 = (w2771 & w39126) | (w2771 & w39127) | (w39126 & w39127);
assign w5915 = (~w2771 & w39128) | (~w2771 & w39129) | (w39128 & w39129);
assign w5916 = ~w5913 & ~w5914;
assign w5917 = ~w5915 & ~w5916;
assign w5918 = b_16 & w2639;
assign w5919 = w2820 & w28776;
assign w5920 = b_15 & w2634;
assign w5921 = ~w5919 & ~w5920;
assign w5922 = ~w5918 & w5921;
assign w5923 = (w5922 & ~w926) | (w5922 & w28777) | (~w926 & w28777);
assign w5924 = (w926 & w39130) | (w926 & w39131) | (w39130 & w39131);
assign w5925 = (~w926 & w39132) | (~w926 & w39133) | (w39132 & w39133);
assign w5926 = ~w5923 & ~w5924;
assign w5927 = ~w5925 & ~w5926;
assign w5928 = ~w5735 & ~w5739;
assign w5929 = (~w5730 & w5679) | (~w5730 & w26785) | (w5679 & w26785);
assign w5930 = b_7 & w4499;
assign w5931 = w4723 & w28778;
assign w5932 = b_6 & w4494;
assign w5933 = ~w5931 & ~w5932;
assign w5934 = ~w5930 & w5933;
assign w5935 = (w5934 & ~w213) | (w5934 & w28779) | (~w213 & w28779);
assign w5936 = (w213 & w39134) | (w213 & w39135) | (w39134 & w39135);
assign w5937 = (~w213 & w39136) | (~w213 & w39137) | (w39136 & w39137);
assign w5938 = ~w5935 & ~w5936;
assign w5939 = ~w5937 & ~w5938;
assign w5940 = ~w5469 & w28780;
assign w5941 = (~w5940 & w5696) | (~w5940 & w28781) | (w5696 & w28781);
assign w5942 = b_4 & w5196;
assign w5943 = w5459 & w26146;
assign w5944 = b_3 & w5191;
assign w5945 = ~w5943 & ~w5944;
assign w5946 = ~w5942 & w5945;
assign w5947 = w84 & w5199;
assign w5948 = w5946 & ~w5947;
assign w5949 = (a_41 & w5947) | (a_41 & w26147) | (w5947 & w26147);
assign w5950 = ~w5947 & w26554;
assign w5951 = ~w5948 & ~w5949;
assign w5952 = ~w5950 & ~w5951;
assign w5953 = (a_44 & w5692) | (a_44 & w28782) | (w5692 & w28782);
assign w5954 = ~a_42 & a_43;
assign w5955 = a_42 & ~a_43;
assign w5956 = ~w5954 & ~w5955;
assign w5957 = w5692 & ~w5956;
assign w5958 = b_0 & w5957;
assign w5959 = ~a_43 & a_44;
assign w5960 = a_43 & ~a_44;
assign w5961 = ~w5959 & ~w5960;
assign w5962 = ~w5692 & w5961;
assign w5963 = b_1 & w5962;
assign w5964 = ~w5958 & ~w5963;
assign w5965 = ~w5692 & ~w5961;
assign w5966 = ~w15 & w5965;
assign w5967 = w5964 & ~w5966;
assign w5968 = (a_44 & ~w5964) | (a_44 & w25551) | (~w5964 & w25551);
assign w5969 = w5964 & w25802;
assign w5970 = ~w5967 & ~w5968;
assign w5971 = (w5953 & w5970) | (w5953 & w25803) | (w5970 & w25803);
assign w5972 = ~w5970 & w26555;
assign w5973 = ~w5971 & ~w5972;
assign w5974 = w5952 & ~w5973;
assign w5975 = ~w5952 & w5973;
assign w5976 = ~w5974 & ~w5975;
assign w5977 = ~w5941 & w5976;
assign w5978 = w5941 & ~w5976;
assign w5979 = ~w5977 & ~w5978;
assign w5980 = ~w5939 & w5979;
assign w5981 = w5979 & ~w5980;
assign w5982 = ~w5979 & ~w5939;
assign w5983 = ~w5981 & ~w5982;
assign w5984 = ~w5711 & ~w5717;
assign w5985 = w5983 & w5984;
assign w5986 = ~w5983 & ~w5984;
assign w5987 = ~w5985 & ~w5986;
assign w5988 = b_10 & w3803;
assign w5989 = w4027 & w28783;
assign w5990 = b_9 & w3798;
assign w5991 = ~w5989 & ~w5990;
assign w5992 = ~w5988 & w5991;
assign w5993 = (w5992 & ~w454) | (w5992 & w28784) | (~w454 & w28784);
assign w5994 = (w454 & w39138) | (w454 & w39139) | (w39138 & w39139);
assign w5995 = (~w454 & w39140) | (~w454 & w39141) | (w39140 & w39141);
assign w5996 = ~w5993 & ~w5994;
assign w5997 = ~w5995 & ~w5996;
assign w5998 = w5987 & ~w5997;
assign w5999 = ~w5987 & w5997;
assign w6000 = ~w5929 & w26903;
assign w6001 = ~w5929 & ~w6000;
assign w6002 = ~w5998 & ~w6000;
assign w6003 = ~w6000 & w26903;
assign w6004 = ~w6001 & ~w6003;
assign w6005 = b_13 & w3195;
assign w6006 = w3388 & w28785;
assign w6007 = b_12 & w3190;
assign w6008 = ~w6006 & ~w6007;
assign w6009 = ~w6005 & w6008;
assign w6010 = (w6009 & ~w711) | (w6009 & w28786) | (~w711 & w28786);
assign w6011 = (w711 & w39142) | (w711 & w39143) | (w39142 & w39143);
assign w6012 = (~w711 & w39144) | (~w711 & w39145) | (w39144 & w39145);
assign w6013 = ~w6010 & ~w6011;
assign w6014 = ~w6012 & ~w6013;
assign w6015 = w6004 & w6014;
assign w6016 = ~w6004 & ~w6014;
assign w6017 = ~w6015 & ~w6016;
assign w6018 = ~w5928 & w6017;
assign w6019 = w5928 & ~w6017;
assign w6020 = ~w6018 & ~w6019;
assign w6021 = ~w5927 & w6020;
assign w6022 = w6020 & ~w6021;
assign w6023 = ~w6020 & ~w5927;
assign w6024 = ~w6022 & ~w6023;
assign w6025 = (~w5753 & w5756) | (~w5753 & w27140) | (w5756 & w27140);
assign w6026 = w6024 & w6025;
assign w6027 = ~w6024 & ~w6025;
assign w6028 = ~w6026 & ~w6027;
assign w6029 = b_19 & w2158;
assign w6030 = w2294 & w28787;
assign w6031 = b_18 & w2153;
assign w6032 = ~w6030 & ~w6031;
assign w6033 = ~w6029 & w6032;
assign w6034 = (w6033 & ~w1372) | (w6033 & w28788) | (~w1372 & w28788);
assign w6035 = (w1372 & w39146) | (w1372 & w39147) | (w39146 & w39147);
assign w6036 = (~w1372 & w39148) | (~w1372 & w39149) | (w39148 & w39149);
assign w6037 = ~w6034 & ~w6035;
assign w6038 = ~w6036 & ~w6037;
assign w6039 = w6028 & ~w6038;
assign w6040 = w6028 & ~w6039;
assign w6041 = ~w6028 & ~w6038;
assign w6042 = ~w6040 & ~w6041;
assign w6043 = ~w5770 & ~w5773;
assign w6044 = w6042 & w6043;
assign w6045 = ~w6042 & ~w6043;
assign w6046 = ~w6044 & ~w6045;
assign w6047 = b_22 & w1694;
assign w6048 = w1834 & w28789;
assign w6049 = b_21 & w1689;
assign w6050 = ~w6048 & ~w6049;
assign w6051 = ~w6047 & w6050;
assign w6052 = (w6051 & ~w1786) | (w6051 & w28790) | (~w1786 & w28790);
assign w6053 = (w1786 & w39150) | (w1786 & w39151) | (w39150 & w39151);
assign w6054 = (~w1786 & w39152) | (~w1786 & w39153) | (w39152 & w39153);
assign w6055 = ~w6052 & ~w6053;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = w6046 & ~w6056;
assign w6058 = w6046 & ~w6057;
assign w6059 = ~w6046 & ~w6056;
assign w6060 = ~w6058 & ~w6059;
assign w6061 = ~w5776 & ~w5782;
assign w6062 = w6060 & w6061;
assign w6063 = ~w6060 & ~w6061;
assign w6064 = ~w6062 & ~w6063;
assign w6065 = b_25 & w1295;
assign w6066 = w1422 & w28791;
assign w6067 = b_24 & w1290;
assign w6068 = ~w6066 & ~w6067;
assign w6069 = ~w6065 & w6068;
assign w6070 = (w6069 & ~w2108) | (w6069 & w28792) | (~w2108 & w28792);
assign w6071 = (w2108 & w39154) | (w2108 & w39155) | (w39154 & w39155);
assign w6072 = (~w2108 & w39156) | (~w2108 & w39157) | (w39156 & w39157);
assign w6073 = ~w6070 & ~w6071;
assign w6074 = ~w6072 & ~w6073;
assign w6075 = w6064 & ~w6074;
assign w6076 = w6064 & ~w6075;
assign w6077 = ~w6064 & ~w6074;
assign w6078 = ~w6076 & ~w6077;
assign w6079 = (~w5795 & w5547) | (~w5795 & w27527) | (w5547 & w27527);
assign w6080 = (~w6079 & w6076) | (~w6079 & w27528) | (w6076 & w27528);
assign w6081 = ~w6076 & w27529;
assign w6082 = ~w6080 & ~w6081;
assign w6083 = ~w5917 & w6082;
assign w6084 = ~w6082 & ~w5917;
assign w6085 = w6082 & ~w6083;
assign w6086 = ~w6084 & ~w6085;
assign w6087 = (~w5907 & w6085) | (~w5907 & w39158) | (w6085 & w39158);
assign w6088 = ~w6086 & ~w6087;
assign w6089 = b_31 & w657;
assign w6090 = w754 & w28793;
assign w6091 = b_30 & w652;
assign w6092 = ~w6090 & ~w6091;
assign w6093 = ~w6089 & w6092;
assign w6094 = (w6093 & ~w3345) | (w6093 & w28794) | (~w3345 & w28794);
assign w6095 = (w3345 & w39159) | (w3345 & w39160) | (w39159 & w39160);
assign w6096 = (~w3345 & w39161) | (~w3345 & w39162) | (w39161 & w39162);
assign w6097 = ~w6094 & ~w6095;
assign w6098 = ~w6096 & ~w6097;
assign w6099 = ~w6088 & w27414;
assign w6100 = (~w6098 & w6088) | (~w6098 & w27415) | (w6088 & w27415);
assign w6101 = ~w6099 & ~w6100;
assign w6102 = ~w5906 & w6101;
assign w6103 = w5906 & ~w6101;
assign w6104 = ~w6102 & ~w6103;
assign w6105 = ~w5905 & w6104;
assign w6106 = w6104 & ~w6105;
assign w6107 = ~w6104 & ~w5905;
assign w6108 = ~w6106 & ~w6107;
assign w6109 = ~w5633 & ~w5826;
assign w6110 = ~w5823 & ~w6109;
assign w6111 = w6108 & w6110;
assign w6112 = ~w6108 & ~w6110;
assign w6113 = ~w6111 & ~w6112;
assign w6114 = b_37 & w239;
assign w6115 = w266 & w28795;
assign w6116 = b_36 & w234;
assign w6117 = ~w6115 & ~w6116;
assign w6118 = ~w6114 & w6117;
assign w6119 = (w6118 & ~w4636) | (w6118 & w28796) | (~w4636 & w28796);
assign w6120 = (w4636 & w39163) | (w4636 & w39164) | (w39163 & w39164);
assign w6121 = (~w4636 & w39165) | (~w4636 & w39166) | (w39165 & w39166);
assign w6122 = ~w6119 & ~w6120;
assign w6123 = ~w6121 & ~w6122;
assign w6124 = w6113 & ~w6123;
assign w6125 = ~w6113 & w6123;
assign w6126 = ~w5895 & w28797;
assign w6127 = ~w5895 & ~w6126;
assign w6128 = ~w6124 & ~w6126;
assign w6129 = ~w6126 & w28797;
assign w6130 = ~w6127 & ~w6129;
assign w6131 = b_40 & w99;
assign w6132 = w136 & w28798;
assign w6133 = b_39 & w94;
assign w6134 = ~w6132 & ~w6133;
assign w6135 = ~w6131 & w6134;
assign w6136 = (w6135 & ~w5363) | (w6135 & w28799) | (~w5363 & w28799);
assign w6137 = (w5363 & w39167) | (w5363 & w39168) | (w39167 & w39168);
assign w6138 = (~w5363 & w39169) | (~w5363 & w39170) | (w39169 & w39170);
assign w6139 = ~w6136 & ~w6137;
assign w6140 = ~w6138 & ~w6139;
assign w6141 = w6130 & w6140;
assign w6142 = ~w6130 & ~w6140;
assign w6143 = ~w6141 & ~w6142;
assign w6144 = ~w5894 & w6143;
assign w6145 = w5894 & ~w6143;
assign w6146 = ~w6144 & ~w6145;
assign w6147 = ~w5893 & w6146;
assign w6148 = w6146 & ~w6147;
assign w6149 = ~w6146 & ~w5893;
assign w6150 = ~w6148 & ~w6149;
assign w6151 = (~w5870 & w5873) | (~w5870 & w28800) | (w5873 & w28800);
assign w6152 = ~w6150 & ~w6151;
assign w6153 = w6150 & w6151;
assign w6154 = ~w6152 & ~w6153;
assign w6155 = ~w6147 & ~w6152;
assign w6156 = ~w6142 & ~w6144;
assign w6157 = b_41 & w99;
assign w6158 = w136 & w28801;
assign w6159 = b_40 & w94;
assign w6160 = ~w6158 & ~w6159;
assign w6161 = ~w6157 & w6160;
assign w6162 = (w6161 & ~w5609) | (w6161 & w28802) | (~w5609 & w28802);
assign w6163 = (w5609 & w39171) | (w5609 & w39172) | (w39171 & w39172);
assign w6164 = (~w5609 & w39173) | (~w5609 & w39174) | (w39173 & w39174);
assign w6165 = ~w6162 & ~w6163;
assign w6166 = ~w6164 & ~w6165;
assign w6167 = b_35 & w418;
assign w6168 = w481 & w28803;
assign w6169 = b_34 & w413;
assign w6170 = ~w6168 & ~w6169;
assign w6171 = ~w6167 & w6170;
assign w6172 = (w6171 & ~w4181) | (w6171 & w28804) | (~w4181 & w28804);
assign w6173 = (w4181 & w39175) | (w4181 & w39176) | (w39175 & w39176);
assign w6174 = (~w4181 & w39177) | (~w4181 & w39178) | (w39177 & w39178);
assign w6175 = ~w6172 & ~w6173;
assign w6176 = ~w6174 & ~w6175;
assign w6177 = (~w6100 & ~w6101) | (~w6100 & w27530) | (~w6101 & w27530);
assign w6178 = b_32 & w657;
assign w6179 = w754 & w28805;
assign w6180 = b_31 & w652;
assign w6181 = ~w6179 & ~w6180;
assign w6182 = ~w6178 & w6181;
assign w6183 = (w6182 & ~w3545) | (w6182 & w28806) | (~w3545 & w28806);
assign w6184 = (w3545 & w39179) | (w3545 & w39180) | (w39179 & w39180);
assign w6185 = (~w3545 & w39181) | (~w3545 & w39182) | (w39181 & w39182);
assign w6186 = ~w6183 & ~w6184;
assign w6187 = ~w6185 & ~w6186;
assign w6188 = (~w6083 & w6086) | (~w6083 & w27416) | (w6086 & w27416);
assign w6189 = b_29 & w986;
assign w6190 = w1069 & w28807;
assign w6191 = b_28 & w981;
assign w6192 = ~w6190 & ~w6191;
assign w6193 = ~w6189 & w6192;
assign w6194 = (w6193 & ~w2954) | (w6193 & w28808) | (~w2954 & w28808);
assign w6195 = (w2954 & w39183) | (w2954 & w39184) | (w39183 & w39184);
assign w6196 = (~w2954 & w39185) | (~w2954 & w39186) | (w39185 & w39186);
assign w6197 = ~w6194 & ~w6195;
assign w6198 = ~w6196 & ~w6197;
assign w6199 = (~w6075 & w6078) | (~w6075 & w27417) | (w6078 & w27417);
assign w6200 = (~w6057 & w6060) | (~w6057 & w27219) | (w6060 & w27219);
assign w6201 = b_20 & w2158;
assign w6202 = w2294 & w28809;
assign w6203 = b_19 & w2153;
assign w6204 = ~w6202 & ~w6203;
assign w6205 = ~w6201 & w6204;
assign w6206 = (w6205 & ~w1503) | (w6205 & w28810) | (~w1503 & w28810);
assign w6207 = (w1503 & w39187) | (w1503 & w39188) | (w39187 & w39188);
assign w6208 = (~w1503 & w39189) | (~w1503 & w39190) | (w39189 & w39190);
assign w6209 = ~w6206 & ~w6207;
assign w6210 = ~w6208 & ~w6209;
assign w6211 = b_17 & w2639;
assign w6212 = w2820 & w28811;
assign w6213 = b_16 & w2634;
assign w6214 = ~w6212 & ~w6213;
assign w6215 = ~w6211 & w6214;
assign w6216 = (w6215 & ~w1038) | (w6215 & w28812) | (~w1038 & w28812);
assign w6217 = (w1038 & w39191) | (w1038 & w39192) | (w39191 & w39192);
assign w6218 = (~w1038 & w39193) | (~w1038 & w39194) | (w39193 & w39194);
assign w6219 = ~w6216 & ~w6217;
assign w6220 = ~w6218 & ~w6219;
assign w6221 = (~w6016 & w5928) | (~w6016 & w27141) | (w5928 & w27141);
assign w6222 = b_14 & w3195;
assign w6223 = w3388 & w28813;
assign w6224 = b_13 & w3190;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = ~w6222 & w6225;
assign w6227 = (w6226 & ~w735) | (w6226 & w28814) | (~w735 & w28814);
assign w6228 = (w735 & w39195) | (w735 & w39196) | (w39195 & w39196);
assign w6229 = (~w735 & w39197) | (~w735 & w39198) | (w39197 & w39198);
assign w6230 = ~w6227 & ~w6228;
assign w6231 = ~w6229 & ~w6230;
assign w6232 = (~w5980 & w5984) | (~w5980 & w28815) | (w5984 & w28815);
assign w6233 = b_8 & w4499;
assign w6234 = w4723 & w28816;
assign w6235 = b_7 & w4494;
assign w6236 = ~w6234 & ~w6235;
assign w6237 = ~w6233 & w6236;
assign w6238 = ~w308 & w28817;
assign w6239 = (w6237 & ~w28817) | (w6237 & w39199) | (~w28817 & w39199);
assign w6240 = (w28817 & w39200) | (w28817 & w39201) | (w39200 & w39201);
assign w6241 = ~w6238 & w28819;
assign w6242 = ~w6239 & ~w6240;
assign w6243 = ~w6241 & ~w6242;
assign w6244 = (~w5975 & w5941) | (~w5975 & w26148) | (w5941 & w26148);
assign w6245 = b_2 & w5962;
assign w6246 = w5692 & ~w5961;
assign w6247 = w6246 & w25371;
assign w6248 = b_1 & w5957;
assign w6249 = ~w6247 & ~w6248;
assign w6250 = ~w6245 & w6249;
assign w6251 = w35 & w5965;
assign w6252 = w6250 & ~w6251;
assign w6253 = (a_44 & ~w6250) | (a_44 & w25552) | (~w6250 & w25552);
assign w6254 = w6250 & w25804;
assign w6255 = ~w6252 & ~w6253;
assign w6256 = ~w6254 & ~w6255;
assign w6257 = ~w5971 & w6256;
assign w6258 = w5971 & ~w6256;
assign w6259 = ~w6257 & ~w6258;
assign w6260 = b_5 & w5196;
assign w6261 = w5459 & w26556;
assign w6262 = b_4 & w5191;
assign w6263 = ~w6261 & ~w6262;
assign w6264 = ~w6260 & w6263;
assign w6265 = w129 & w5199;
assign w6266 = w6264 & ~w6265;
assign w6267 = (a_41 & w6265) | (a_41 & w26557) | (w6265 & w26557);
assign w6268 = ~w6265 & w39202;
assign w6269 = ~w6266 & ~w6267;
assign w6270 = ~w6268 & ~w6269;
assign w6271 = w6259 & ~w6270;
assign w6272 = w6259 & ~w6271;
assign w6273 = ~w6259 & ~w6270;
assign w6274 = ~w6272 & ~w6273;
assign w6275 = ~w6244 & ~w6274;
assign w6276 = w6244 & w6274;
assign w6277 = ~w6275 & ~w6276;
assign w6278 = ~w6243 & w6277;
assign w6279 = ~w6277 & ~w6243;
assign w6280 = w6277 & ~w6278;
assign w6281 = ~w6279 & ~w6280;
assign w6282 = ~w6232 & ~w6281;
assign w6283 = ~w6232 & ~w6282;
assign w6284 = b_11 & w3803;
assign w6285 = w4027 & w28820;
assign w6286 = b_10 & w3798;
assign w6287 = ~w6285 & ~w6286;
assign w6288 = ~w6284 & w6287;
assign w6289 = (w6288 & ~w530) | (w6288 & w28821) | (~w530 & w28821);
assign w6290 = (w530 & w39203) | (w530 & w39204) | (w39203 & w39204);
assign w6291 = (~w530 & w39205) | (~w530 & w39206) | (w39205 & w39206);
assign w6292 = ~w6289 & ~w6290;
assign w6293 = ~w6291 & ~w6292;
assign w6294 = ~w6283 & w26904;
assign w6295 = (~w6293 & w6283) | (~w6293 & w26905) | (w6283 & w26905);
assign w6296 = ~w6294 & ~w6295;
assign w6297 = ~w6002 & w6296;
assign w6298 = w6002 & ~w6296;
assign w6299 = ~w6297 & ~w6298;
assign w6300 = w6231 & ~w6299;
assign w6301 = ~w6231 & w6299;
assign w6302 = ~w6300 & ~w6301;
assign w6303 = ~w6221 & w6302;
assign w6304 = w6221 & ~w6302;
assign w6305 = ~w6303 & ~w6304;
assign w6306 = w6220 & ~w6305;
assign w6307 = ~w6220 & w6305;
assign w6308 = ~w6306 & ~w6307;
assign w6309 = (w6308 & w6027) | (w6308 & w27220) | (w6027 & w27220);
assign w6310 = ~w6027 & w27221;
assign w6311 = ~w6309 & ~w6310;
assign w6312 = ~w6210 & w6311;
assign w6313 = w6311 & ~w6312;
assign w6314 = ~w6311 & ~w6210;
assign w6315 = ~w6313 & ~w6314;
assign w6316 = (~w6039 & w6042) | (~w6039 & w27222) | (w6042 & w27222);
assign w6317 = w6315 & w6316;
assign w6318 = ~w6315 & ~w6316;
assign w6319 = ~w6317 & ~w6318;
assign w6320 = b_23 & w1694;
assign w6321 = w1834 & w28822;
assign w6322 = b_22 & w1689;
assign w6323 = ~w6321 & ~w6322;
assign w6324 = ~w6320 & w6323;
assign w6325 = (w6324 & ~w1933) | (w6324 & w28823) | (~w1933 & w28823);
assign w6326 = (w1933 & w39207) | (w1933 & w39208) | (w39207 & w39208);
assign w6327 = (~w1933 & w39209) | (~w1933 & w39210) | (w39209 & w39210);
assign w6328 = ~w6325 & ~w6326;
assign w6329 = ~w6327 & ~w6328;
assign w6330 = w6319 & ~w6329;
assign w6331 = ~w6319 & w6329;
assign w6332 = ~w6200 & w27343;
assign w6333 = ~w6200 & ~w6332;
assign w6334 = (~w6330 & w6200) | (~w6330 & w27418) | (w6200 & w27418);
assign w6335 = (w27418 & w27343) | (w27418 & w39211) | (w27343 & w39211);
assign w6336 = ~w6333 & ~w6335;
assign w6337 = b_26 & w1295;
assign w6338 = w1422 & w28824;
assign w6339 = b_25 & w1290;
assign w6340 = ~w6338 & ~w6339;
assign w6341 = ~w6337 & w6340;
assign w6342 = (w6341 & ~w2416) | (w6341 & w28825) | (~w2416 & w28825);
assign w6343 = (w2416 & w39212) | (w2416 & w39213) | (w39212 & w39213);
assign w6344 = (~w2416 & w39214) | (~w2416 & w39215) | (w39214 & w39215);
assign w6345 = ~w6342 & ~w6343;
assign w6346 = ~w6344 & ~w6345;
assign w6347 = w6336 & w6346;
assign w6348 = ~w6336 & ~w6346;
assign w6349 = ~w6347 & ~w6348;
assign w6350 = ~w6199 & w6349;
assign w6351 = w6199 & ~w6349;
assign w6352 = ~w6350 & ~w6351;
assign w6353 = w6198 & ~w6352;
assign w6354 = ~w6198 & w6352;
assign w6355 = ~w6353 & ~w6354;
assign w6356 = ~w6188 & w6355;
assign w6357 = w6188 & ~w6355;
assign w6358 = ~w6356 & ~w6357;
assign w6359 = w6187 & ~w6358;
assign w6360 = ~w6187 & w6358;
assign w6361 = ~w6359 & ~w6360;
assign w6362 = ~w6177 & w6361;
assign w6363 = w6177 & ~w6361;
assign w6364 = ~w6362 & ~w6363;
assign w6365 = ~w6176 & w6364;
assign w6366 = w6364 & ~w6365;
assign w6367 = ~w6364 & ~w6176;
assign w6368 = ~w6366 & ~w6367;
assign w6369 = (~w6105 & w6110) | (~w6105 & w27735) | (w6110 & w27735);
assign w6370 = w6368 & w6369;
assign w6371 = ~w6368 & ~w6369;
assign w6372 = ~w6370 & ~w6371;
assign w6373 = b_38 & w239;
assign w6374 = w266 & w28826;
assign w6375 = b_37 & w234;
assign w6376 = ~w6374 & ~w6375;
assign w6377 = ~w6373 & w6376;
assign w6378 = (w6377 & ~w4658) | (w6377 & w25047) | (~w4658 & w25047);
assign w6379 = (w4658 & w28827) | (w4658 & w28828) | (w28827 & w28828);
assign w6380 = (~w4658 & w28829) | (~w4658 & w28830) | (w28829 & w28830);
assign w6381 = ~w6378 & ~w6379;
assign w6382 = ~w6380 & ~w6381;
assign w6383 = w6372 & ~w6382;
assign w6384 = w6372 & ~w6383;
assign w6385 = ~w6372 & ~w6382;
assign w6386 = ~w6384 & ~w6385;
assign w6387 = ~w6128 & ~w6386;
assign w6388 = w6128 & w6386;
assign w6389 = ~w6387 & ~w6388;
assign w6390 = ~w6166 & w6389;
assign w6391 = ~w6389 & ~w6166;
assign w6392 = w6389 & ~w6390;
assign w6393 = ~w6391 & ~w6392;
assign w6394 = ~w6156 & ~w6393;
assign w6395 = ~w6156 & ~w6394;
assign w6396 = ~w6393 & ~w6394;
assign w6397 = ~w6395 & ~w6396;
assign w6398 = w8 & w28831;
assign w6399 = ~w8 & w28832;
assign w6400 = b_43 & w4;
assign w6401 = ~w6399 & ~w6400;
assign w6402 = ~w6398 & w6401;
assign w6403 = ~b_43 & ~b_44;
assign w6404 = b_43 & b_44;
assign w6405 = ~w6403 & ~w6404;
assign w6406 = (w4656 & w28834) | (w4656 & w28835) | (w28834 & w28835);
assign w6407 = (~w4656 & w28836) | (~w4656 & w28837) | (w28836 & w28837);
assign w6408 = ~w6406 & ~w6407;
assign w6409 = (w6402 & ~w6408) | (w6402 & w28838) | (~w6408 & w28838);
assign w6410 = (w6408 & w39216) | (w6408 & w39217) | (w39216 & w39217);
assign w6411 = (~w6408 & w39218) | (~w6408 & w39219) | (w39218 & w39219);
assign w6412 = ~w6409 & ~w6410;
assign w6413 = ~w6411 & ~w6412;
assign w6414 = ~w6397 & w6413;
assign w6415 = w6397 & ~w6413;
assign w6416 = ~w6414 & ~w6415;
assign w6417 = ~w6155 & ~w6416;
assign w6418 = w6155 & w6416;
assign w6419 = ~w6417 & ~w6418;
assign w6420 = ~w6397 & ~w6413;
assign w6421 = ~w6417 & ~w6420;
assign w6422 = (~w6365 & w6369) | (~w6365 & w27531) | (w6369 & w27531);
assign w6423 = (~w6360 & w6177) | (~w6360 & w28839) | (w6177 & w28839);
assign w6424 = b_33 & w657;
assign w6425 = w754 & w28840;
assign w6426 = b_32 & w652;
assign w6427 = ~w6425 & ~w6426;
assign w6428 = ~w6424 & w6427;
assign w6429 = (w6428 & ~w3744) | (w6428 & w28841) | (~w3744 & w28841);
assign w6430 = (w3744 & w39220) | (w3744 & w39221) | (w39220 & w39221);
assign w6431 = (~w3744 & w39222) | (~w3744 & w39223) | (w39222 & w39223);
assign w6432 = ~w6429 & ~w6430;
assign w6433 = ~w6431 & ~w6432;
assign w6434 = (~w6354 & w6188) | (~w6354 & w27532) | (w6188 & w27532);
assign w6435 = (~w6348 & ~w6349) | (~w6348 & w28842) | (~w6349 & w28842);
assign w6436 = b_27 & w1295;
assign w6437 = w1422 & w28843;
assign w6438 = b_26 & w1290;
assign w6439 = ~w6437 & ~w6438;
assign w6440 = ~w6436 & w6439;
assign w6441 = (w6440 & ~w2582) | (w6440 & w28844) | (~w2582 & w28844);
assign w6442 = (w2582 & w39224) | (w2582 & w39225) | (w39224 & w39225);
assign w6443 = (~w2582 & w39226) | (~w2582 & w39227) | (w39226 & w39227);
assign w6444 = ~w6441 & ~w6442;
assign w6445 = ~w6443 & ~w6444;
assign w6446 = b_21 & w2158;
assign w6447 = w2294 & w28845;
assign w6448 = b_20 & w2153;
assign w6449 = ~w6447 & ~w6448;
assign w6450 = ~w6446 & w6449;
assign w6451 = (w6450 & ~w1634) | (w6450 & w28846) | (~w1634 & w28846);
assign w6452 = (w1634 & w39228) | (w1634 & w39229) | (w39228 & w39229);
assign w6453 = (~w1634 & w39230) | (~w1634 & w39231) | (w39230 & w39231);
assign w6454 = ~w6451 & ~w6452;
assign w6455 = ~w6453 & ~w6454;
assign w6456 = (~w27220 & w28847) | (~w27220 & w28848) | (w28847 & w28848);
assign w6457 = (~w6301 & w6221) | (~w6301 & w27223) | (w6221 & w27223);
assign w6458 = (~w6295 & w6002) | (~w6295 & w28849) | (w6002 & w28849);
assign w6459 = b_12 & w3803;
assign w6460 = w4027 & w28850;
assign w6461 = b_11 & w3798;
assign w6462 = ~w6460 & ~w6461;
assign w6463 = ~w6459 & w6462;
assign w6464 = (w6463 & ~w552) | (w6463 & w28851) | (~w552 & w28851);
assign w6465 = (w552 & w39232) | (w552 & w39233) | (w39232 & w39233);
assign w6466 = (~w552 & w39234) | (~w552 & w39235) | (w39234 & w39235);
assign w6467 = ~w6464 & ~w6465;
assign w6468 = ~w6466 & ~w6467;
assign w6469 = (~w6278 & w6232) | (~w6278 & w26558) | (w6232 & w26558);
assign w6470 = b_6 & w5196;
assign w6471 = w5459 & w28852;
assign w6472 = b_5 & w5191;
assign w6473 = ~w6471 & ~w6472;
assign w6474 = ~w6470 & w6473;
assign w6475 = (w6474 & ~w190) | (w6474 & w28853) | (~w190 & w28853);
assign w6476 = (w190 & w39236) | (w190 & w39237) | (w39236 & w39237);
assign w6477 = (~w190 & w39238) | (~w190 & w39239) | (w39238 & w39239);
assign w6478 = ~w6475 & ~w6476;
assign w6479 = ~w6477 & ~w6478;
assign w6480 = a_44 & ~a_45;
assign w6481 = ~a_44 & a_45;
assign w6482 = ~w6480 & ~w6481;
assign w6483 = b_0 & ~w6482;
assign w6484 = (w6483 & w6256) | (w6483 & w25805) | (w6256 & w25805);
assign w6485 = ~w6256 & w25806;
assign w6486 = ~w6484 & ~w6485;
assign w6487 = b_3 & w5962;
assign w6488 = w6246 & w26149;
assign w6489 = b_2 & w5957;
assign w6490 = ~w6488 & ~w6489;
assign w6491 = ~w6487 & w6490;
assign w6492 = w57 & w5965;
assign w6493 = w6491 & ~w6492;
assign w6494 = a_44 & ~w6493;
assign w6495 = w6493 & a_44;
assign w6496 = ~w6493 & ~w6494;
assign w6497 = ~w6495 & ~w6496;
assign w6498 = ~w6486 & ~w6497;
assign w6499 = w6486 & w6497;
assign w6500 = ~w6498 & ~w6499;
assign w6501 = ~w6479 & w6500;
assign w6502 = w6500 & ~w6501;
assign w6503 = ~w6500 & ~w6479;
assign w6504 = ~w6502 & ~w6503;
assign w6505 = ~w6271 & ~w6275;
assign w6506 = w6504 & w6505;
assign w6507 = ~w6504 & ~w6505;
assign w6508 = ~w6506 & ~w6507;
assign w6509 = b_9 & w4499;
assign w6510 = w4723 & w28854;
assign w6511 = b_8 & w4494;
assign w6512 = ~w6510 & ~w6511;
assign w6513 = ~w6509 & w6512;
assign w6514 = (w6513 & ~w371) | (w6513 & w28855) | (~w371 & w28855);
assign w6515 = (w371 & w39240) | (w371 & w39241) | (w39240 & w39241);
assign w6516 = (~w371 & w39242) | (~w371 & w39243) | (w39242 & w39243);
assign w6517 = ~w6514 & ~w6515;
assign w6518 = ~w6516 & ~w6517;
assign w6519 = ~w6508 & w6518;
assign w6520 = w6508 & ~w6518;
assign w6521 = ~w6519 & ~w6520;
assign w6522 = ~w6469 & w6521;
assign w6523 = w6469 & ~w6521;
assign w6524 = ~w6522 & ~w6523;
assign w6525 = ~w6468 & w6524;
assign w6526 = ~w6524 & ~w6468;
assign w6527 = w6524 & ~w6525;
assign w6528 = ~w6526 & ~w6527;
assign w6529 = ~w6458 & ~w6528;
assign w6530 = ~w6458 & ~w6529;
assign w6531 = ~w6528 & ~w6529;
assign w6532 = ~w6530 & ~w6531;
assign w6533 = b_15 & w3195;
assign w6534 = w3388 & w28856;
assign w6535 = b_14 & w3190;
assign w6536 = ~w6534 & ~w6535;
assign w6537 = ~w6533 & w6536;
assign w6538 = (w6537 & ~w827) | (w6537 & w28857) | (~w827 & w28857);
assign w6539 = (w827 & w39244) | (w827 & w39245) | (w39244 & w39245);
assign w6540 = (~w827 & w39246) | (~w827 & w39247) | (w39246 & w39247);
assign w6541 = ~w6538 & ~w6539;
assign w6542 = ~w6540 & ~w6541;
assign w6543 = ~w6532 & ~w6542;
assign w6544 = ~w6532 & ~w6543;
assign w6545 = w6532 & ~w6542;
assign w6546 = ~w6544 & ~w6545;
assign w6547 = ~w6544 & w27224;
assign w6548 = (w6457 & w6544) | (w6457 & w27225) | (w6544 & w27225);
assign w6549 = ~w6547 & ~w6548;
assign w6550 = b_18 & w2639;
assign w6551 = w2820 & w28858;
assign w6552 = b_17 & w2634;
assign w6553 = ~w6551 & ~w6552;
assign w6554 = ~w6550 & w6553;
assign w6555 = (w6554 & ~w1238) | (w6554 & w28859) | (~w1238 & w28859);
assign w6556 = (w1238 & w39248) | (w1238 & w39249) | (w39248 & w39249);
assign w6557 = (~w1238 & w39250) | (~w1238 & w39251) | (w39250 & w39251);
assign w6558 = ~w6555 & ~w6556;
assign w6559 = ~w6557 & ~w6558;
assign w6560 = ~w6549 & ~w6559;
assign w6561 = w6549 & w6559;
assign w6562 = ~w6560 & ~w6561;
assign w6563 = ~w6456 & w6562;
assign w6564 = w6456 & ~w6562;
assign w6565 = ~w6563 & ~w6564;
assign w6566 = ~w6455 & w6565;
assign w6567 = w6565 & ~w6566;
assign w6568 = ~w6565 & ~w6455;
assign w6569 = ~w6567 & ~w6568;
assign w6570 = (~w6312 & w6315) | (~w6312 & w39252) | (w6315 & w39252);
assign w6571 = w6569 & w6570;
assign w6572 = ~w6569 & ~w6570;
assign w6573 = ~w6571 & ~w6572;
assign w6574 = b_24 & w1694;
assign w6575 = w1834 & w28860;
assign w6576 = b_23 & w1689;
assign w6577 = ~w6575 & ~w6576;
assign w6578 = ~w6574 & w6577;
assign w6579 = (w6578 & ~w2083) | (w6578 & w28861) | (~w2083 & w28861);
assign w6580 = (w2083 & w39253) | (w2083 & w39254) | (w39253 & w39254);
assign w6581 = (~w2083 & w39255) | (~w2083 & w39256) | (w39255 & w39256);
assign w6582 = ~w6579 & ~w6580;
assign w6583 = ~w6581 & ~w6582;
assign w6584 = ~w6573 & w6583;
assign w6585 = w6573 & ~w6583;
assign w6586 = ~w6584 & ~w6585;
assign w6587 = ~w6334 & w6586;
assign w6588 = w6334 & ~w6586;
assign w6589 = ~w6587 & ~w6588;
assign w6590 = ~w6445 & w6589;
assign w6591 = w6589 & ~w6590;
assign w6592 = ~w6589 & ~w6445;
assign w6593 = ~w6591 & ~w6592;
assign w6594 = ~w6435 & w6593;
assign w6595 = w6435 & ~w6593;
assign w6596 = ~w6594 & ~w6595;
assign w6597 = b_30 & w986;
assign w6598 = w1069 & w28862;
assign w6599 = b_29 & w981;
assign w6600 = ~w6598 & ~w6599;
assign w6601 = ~w6597 & w6600;
assign w6602 = (w6601 & ~w3138) | (w6601 & w28863) | (~w3138 & w28863);
assign w6603 = (w3138 & w39257) | (w3138 & w39258) | (w39257 & w39258);
assign w6604 = (~w3138 & w39259) | (~w3138 & w39260) | (w39259 & w39260);
assign w6605 = ~w6602 & ~w6603;
assign w6606 = ~w6604 & ~w6605;
assign w6607 = ~w6596 & ~w6606;
assign w6608 = w6596 & w6606;
assign w6609 = ~w6607 & ~w6608;
assign w6610 = ~w6434 & w6609;
assign w6611 = w6434 & ~w6609;
assign w6612 = ~w6610 & ~w6611;
assign w6613 = ~w6433 & w6612;
assign w6614 = w6612 & ~w6613;
assign w6615 = ~w6612 & ~w6433;
assign w6616 = ~w6614 & ~w6615;
assign w6617 = ~w6423 & w6616;
assign w6618 = w6423 & ~w6616;
assign w6619 = ~w6617 & ~w6618;
assign w6620 = b_36 & w418;
assign w6621 = w481 & w28864;
assign w6622 = b_35 & w413;
assign w6623 = ~w6621 & ~w6622;
assign w6624 = ~w6620 & w6623;
assign w6625 = (w6624 & ~w4395) | (w6624 & w28865) | (~w4395 & w28865);
assign w6626 = (w4395 & w39261) | (w4395 & w39262) | (w39261 & w39262);
assign w6627 = (~w4395 & w39263) | (~w4395 & w39264) | (w39263 & w39264);
assign w6628 = ~w6625 & ~w6626;
assign w6629 = ~w6627 & ~w6628;
assign w6630 = ~w6619 & ~w6629;
assign w6631 = w6619 & w6629;
assign w6632 = ~w6630 & ~w6631;
assign w6633 = w6422 & ~w6632;
assign w6634 = ~w6422 & w6632;
assign w6635 = ~w6633 & ~w6634;
assign w6636 = b_39 & w239;
assign w6637 = w266 & w28866;
assign w6638 = b_38 & w234;
assign w6639 = ~w6637 & ~w6638;
assign w6640 = ~w6636 & w6639;
assign w6641 = (w6640 & ~w4888) | (w6640 & w25048) | (~w4888 & w25048);
assign w6642 = (w4888 & w28867) | (w4888 & w28868) | (w28867 & w28868);
assign w6643 = (~w4888 & w28869) | (~w4888 & w28870) | (w28869 & w28870);
assign w6644 = ~w6641 & ~w6642;
assign w6645 = ~w6643 & ~w6644;
assign w6646 = w6635 & ~w6645;
assign w6647 = w6635 & ~w6646;
assign w6648 = ~w6635 & ~w6645;
assign w6649 = ~w6647 & ~w6648;
assign w6650 = ~w6383 & ~w6387;
assign w6651 = w6649 & w6650;
assign w6652 = ~w6649 & ~w6650;
assign w6653 = ~w6651 & ~w6652;
assign w6654 = b_42 & w99;
assign w6655 = w136 & w28871;
assign w6656 = b_41 & w94;
assign w6657 = ~w6655 & ~w6656;
assign w6658 = ~w6654 & w6657;
assign w6659 = (w6658 & ~w5864) | (w6658 & w28872) | (~w5864 & w28872);
assign w6660 = (w5864 & w39265) | (w5864 & w39266) | (w39265 & w39266);
assign w6661 = (~w5864 & w39267) | (~w5864 & w39268) | (w39267 & w39268);
assign w6662 = ~w6659 & ~w6660;
assign w6663 = ~w6661 & ~w6662;
assign w6664 = w6653 & ~w6663;
assign w6665 = w6653 & ~w6664;
assign w6666 = ~w6653 & ~w6663;
assign w6667 = ~w6665 & ~w6666;
assign w6668 = (~w6390 & w6156) | (~w6390 & w25049) | (w6156 & w25049);
assign w6669 = w6667 & w6668;
assign w6670 = ~w6667 & ~w6668;
assign w6671 = ~w6669 & ~w6670;
assign w6672 = w8 & w28873;
assign w6673 = ~w8 & w28874;
assign w6674 = b_44 & w4;
assign w6675 = ~w6673 & ~w6674;
assign w6676 = ~w6672 & w6675;
assign w6677 = ~b_44 & ~b_45;
assign w6678 = b_44 & b_45;
assign w6679 = ~w6677 & ~w6678;
assign w6680 = (w4656 & w39269) | (w4656 & w39270) | (w39269 & w39270);
assign w6681 = (~w4656 & w39271) | (~w4656 & w39272) | (w39271 & w39272);
assign w6682 = ~w6680 & ~w6681;
assign w6683 = (w6676 & ~w6682) | (w6676 & w28877) | (~w6682 & w28877);
assign w6684 = (w6682 & w39273) | (w6682 & w39274) | (w39273 & w39274);
assign w6685 = (~w6682 & w39275) | (~w6682 & w39276) | (w39275 & w39276);
assign w6686 = ~w6683 & ~w6684;
assign w6687 = ~w6685 & ~w6686;
assign w6688 = ~w6671 & w6687;
assign w6689 = w6671 & ~w6687;
assign w6690 = ~w6688 & ~w6689;
assign w6691 = (w6690 & w6417) | (w6690 & w25050) | (w6417 & w25050);
assign w6692 = w6421 & ~w6690;
assign w6693 = ~w6691 & ~w6692;
assign w6694 = (~w6646 & w6650) | (~w6646 & w39277) | (w6650 & w39277);
assign w6695 = b_34 & w657;
assign w6696 = w754 & w28878;
assign w6697 = b_33 & w652;
assign w6698 = ~w6696 & ~w6697;
assign w6699 = ~w6695 & w6698;
assign w6700 = (w6699 & ~w3967) | (w6699 & w28879) | (~w3967 & w28879);
assign w6701 = (w3967 & w39278) | (w3967 & w39279) | (w39278 & w39279);
assign w6702 = (~w3967 & w39280) | (~w3967 & w39281) | (w39280 & w39281);
assign w6703 = ~w6700 & ~w6701;
assign w6704 = ~w6702 & ~w6703;
assign w6705 = (~w6607 & w6434) | (~w6607 & w28880) | (w6434 & w28880);
assign w6706 = (~w6590 & w6435) | (~w6590 & w27533) | (w6435 & w27533);
assign w6707 = b_28 & w1295;
assign w6708 = w1422 & w28881;
assign w6709 = b_27 & w1290;
assign w6710 = ~w6708 & ~w6709;
assign w6711 = ~w6707 & w6710;
assign w6712 = (w6711 & ~w2771) | (w6711 & w28882) | (~w2771 & w28882);
assign w6713 = (w2771 & w39282) | (w2771 & w39283) | (w39282 & w39283);
assign w6714 = (~w2771 & w39284) | (~w2771 & w39285) | (w39284 & w39285);
assign w6715 = ~w6712 & ~w6713;
assign w6716 = ~w6714 & ~w6715;
assign w6717 = b_16 & w3195;
assign w6718 = w3388 & w28883;
assign w6719 = b_15 & w3190;
assign w6720 = ~w6718 & ~w6719;
assign w6721 = ~w6717 & w6720;
assign w6722 = (w6721 & ~w926) | (w6721 & w28884) | (~w926 & w28884);
assign w6723 = (w926 & w39286) | (w926 & w39287) | (w39286 & w39287);
assign w6724 = (~w926 & w39288) | (~w926 & w39289) | (w39288 & w39289);
assign w6725 = ~w6722 & ~w6723;
assign w6726 = ~w6724 & ~w6725;
assign w6727 = ~w6525 & ~w6529;
assign w6728 = (~w6520 & w6469) | (~w6520 & w26786) | (w6469 & w26786);
assign w6729 = b_7 & w5196;
assign w6730 = w5459 & w28885;
assign w6731 = b_6 & w5191;
assign w6732 = ~w6730 & ~w6731;
assign w6733 = ~w6729 & w6732;
assign w6734 = (w6733 & ~w213) | (w6733 & w28886) | (~w213 & w28886);
assign w6735 = (w213 & w39290) | (w213 & w39291) | (w39290 & w39291);
assign w6736 = (~w213 & w39292) | (~w213 & w39293) | (w39292 & w39293);
assign w6737 = ~w6734 & ~w6735;
assign w6738 = ~w6736 & ~w6737;
assign w6739 = ~w6256 & w28887;
assign w6740 = (~w6739 & w6486) | (~w6739 & w28888) | (w6486 & w28888);
assign w6741 = b_4 & w5962;
assign w6742 = w6246 & w26150;
assign w6743 = b_3 & w5957;
assign w6744 = ~w6742 & ~w6743;
assign w6745 = ~w6741 & w6744;
assign w6746 = w84 & w5965;
assign w6747 = w6745 & ~w6746;
assign w6748 = (a_44 & w6746) | (a_44 & w26151) | (w6746 & w26151);
assign w6749 = ~w6746 & w27034;
assign w6750 = ~w6747 & ~w6748;
assign w6751 = ~w6749 & ~w6750;
assign w6752 = (a_47 & w6482) | (a_47 & w28889) | (w6482 & w28889);
assign w6753 = ~a_45 & a_46;
assign w6754 = a_45 & ~a_46;
assign w6755 = ~w6753 & ~w6754;
assign w6756 = w6482 & ~w6755;
assign w6757 = b_0 & w6756;
assign w6758 = ~a_46 & a_47;
assign w6759 = a_46 & ~a_47;
assign w6760 = ~w6758 & ~w6759;
assign w6761 = ~w6482 & w6760;
assign w6762 = b_1 & w6761;
assign w6763 = ~w6757 & ~w6762;
assign w6764 = ~w6482 & ~w6760;
assign w6765 = ~w15 & w6764;
assign w6766 = w6763 & ~w6765;
assign w6767 = (a_47 & ~w6763) | (a_47 & w25807) | (~w6763 & w25807);
assign w6768 = w6763 & w26152;
assign w6769 = ~w6766 & ~w6767;
assign w6770 = (w6752 & w6769) | (w6752 & w26153) | (w6769 & w26153);
assign w6771 = ~w6769 & w26787;
assign w6772 = ~w6770 & ~w6771;
assign w6773 = w6751 & ~w6772;
assign w6774 = ~w6751 & w6772;
assign w6775 = ~w6773 & ~w6774;
assign w6776 = ~w6740 & w6775;
assign w6777 = w6740 & ~w6775;
assign w6778 = ~w6776 & ~w6777;
assign w6779 = ~w6738 & w6778;
assign w6780 = w6778 & ~w6779;
assign w6781 = ~w6778 & ~w6738;
assign w6782 = ~w6780 & ~w6781;
assign w6783 = ~w6501 & ~w6507;
assign w6784 = w6782 & w6783;
assign w6785 = ~w6782 & ~w6783;
assign w6786 = ~w6784 & ~w6785;
assign w6787 = b_10 & w4499;
assign w6788 = w4723 & w28890;
assign w6789 = b_9 & w4494;
assign w6790 = ~w6788 & ~w6789;
assign w6791 = ~w6787 & w6790;
assign w6792 = (w6791 & ~w454) | (w6791 & w28891) | (~w454 & w28891);
assign w6793 = (w454 & w39294) | (w454 & w39295) | (w39294 & w39295);
assign w6794 = (~w454 & w39296) | (~w454 & w39297) | (w39296 & w39297);
assign w6795 = ~w6792 & ~w6793;
assign w6796 = ~w6794 & ~w6795;
assign w6797 = w6786 & ~w6796;
assign w6798 = ~w6786 & w6796;
assign w6799 = ~w6728 & w26906;
assign w6800 = ~w6728 & ~w6799;
assign w6801 = ~w6797 & ~w6799;
assign w6802 = ~w6799 & w26906;
assign w6803 = ~w6800 & ~w6802;
assign w6804 = b_13 & w3803;
assign w6805 = w4027 & w28892;
assign w6806 = b_12 & w3798;
assign w6807 = ~w6805 & ~w6806;
assign w6808 = ~w6804 & w6807;
assign w6809 = (w6808 & ~w711) | (w6808 & w28893) | (~w711 & w28893);
assign w6810 = (w711 & w39298) | (w711 & w39299) | (w39298 & w39299);
assign w6811 = (~w711 & w39300) | (~w711 & w39301) | (w39300 & w39301);
assign w6812 = ~w6809 & ~w6810;
assign w6813 = ~w6811 & ~w6812;
assign w6814 = w6803 & w6813;
assign w6815 = ~w6803 & ~w6813;
assign w6816 = ~w6814 & ~w6815;
assign w6817 = ~w6727 & w6816;
assign w6818 = w6727 & ~w6816;
assign w6819 = ~w6817 & ~w6818;
assign w6820 = ~w6726 & w6819;
assign w6821 = w6819 & ~w6820;
assign w6822 = ~w6819 & ~w6726;
assign w6823 = ~w6821 & ~w6822;
assign w6824 = (~w6543 & w6546) | (~w6543 & w27142) | (w6546 & w27142);
assign w6825 = w6823 & w6824;
assign w6826 = ~w6823 & ~w6824;
assign w6827 = ~w6825 & ~w6826;
assign w6828 = b_19 & w2639;
assign w6829 = w2820 & w28894;
assign w6830 = b_18 & w2634;
assign w6831 = ~w6829 & ~w6830;
assign w6832 = ~w6828 & w6831;
assign w6833 = (w6832 & ~w1372) | (w6832 & w28895) | (~w1372 & w28895);
assign w6834 = (w1372 & w39302) | (w1372 & w39303) | (w39302 & w39303);
assign w6835 = (~w1372 & w39304) | (~w1372 & w39305) | (w39304 & w39305);
assign w6836 = ~w6833 & ~w6834;
assign w6837 = ~w6835 & ~w6836;
assign w6838 = w6827 & ~w6837;
assign w6839 = w6827 & ~w6838;
assign w6840 = ~w6827 & ~w6837;
assign w6841 = ~w6839 & ~w6840;
assign w6842 = (~w6560 & w6456) | (~w6560 & w25051) | (w6456 & w25051);
assign w6843 = w6841 & w6842;
assign w6844 = ~w6841 & ~w6842;
assign w6845 = ~w6843 & ~w6844;
assign w6846 = b_22 & w2158;
assign w6847 = w2294 & w28896;
assign w6848 = b_21 & w2153;
assign w6849 = ~w6847 & ~w6848;
assign w6850 = ~w6846 & w6849;
assign w6851 = (w6850 & ~w1786) | (w6850 & w28897) | (~w1786 & w28897);
assign w6852 = (w1786 & w39306) | (w1786 & w39307) | (w39306 & w39307);
assign w6853 = (~w1786 & w39308) | (~w1786 & w39309) | (w39308 & w39309);
assign w6854 = ~w6851 & ~w6852;
assign w6855 = ~w6853 & ~w6854;
assign w6856 = w6845 & ~w6855;
assign w6857 = w6845 & ~w6856;
assign w6858 = ~w6845 & ~w6855;
assign w6859 = ~w6857 & ~w6858;
assign w6860 = (~w6566 & w6570) | (~w6566 & w28898) | (w6570 & w28898);
assign w6861 = w6859 & w6860;
assign w6862 = ~w6859 & ~w6860;
assign w6863 = ~w6861 & ~w6862;
assign w6864 = b_25 & w1694;
assign w6865 = w1834 & w28899;
assign w6866 = b_24 & w1689;
assign w6867 = ~w6865 & ~w6866;
assign w6868 = ~w6864 & w6867;
assign w6869 = (w6868 & ~w2108) | (w6868 & w28900) | (~w2108 & w28900);
assign w6870 = (w2108 & w39310) | (w2108 & w39311) | (w39310 & w39311);
assign w6871 = (~w2108 & w39312) | (~w2108 & w39313) | (w39312 & w39313);
assign w6872 = ~w6869 & ~w6870;
assign w6873 = ~w6871 & ~w6872;
assign w6874 = w6863 & ~w6873;
assign w6875 = w6863 & ~w6874;
assign w6876 = ~w6863 & ~w6873;
assign w6877 = ~w6875 & ~w6876;
assign w6878 = (~w6585 & w6334) | (~w6585 & w39314) | (w6334 & w39314);
assign w6879 = ~w6877 & ~w6878;
assign w6880 = w6877 & w6878;
assign w6881 = ~w6879 & ~w6880;
assign w6882 = ~w6716 & w6881;
assign w6883 = ~w6881 & ~w6716;
assign w6884 = w6881 & ~w6882;
assign w6885 = ~w6883 & ~w6884;
assign w6886 = ~w6706 & ~w6885;
assign w6887 = ~w6885 & ~w6886;
assign w6888 = b_31 & w986;
assign w6889 = w1069 & w28901;
assign w6890 = b_30 & w981;
assign w6891 = ~w6889 & ~w6890;
assign w6892 = ~w6888 & w6891;
assign w6893 = (w6892 & ~w3345) | (w6892 & w28902) | (~w3345 & w28902);
assign w6894 = (w3345 & w39315) | (w3345 & w39316) | (w39315 & w39316);
assign w6895 = (~w3345 & w39317) | (~w3345 & w39318) | (w39317 & w39318);
assign w6896 = ~w6893 & ~w6894;
assign w6897 = ~w6895 & ~w6896;
assign w6898 = ~w6887 & w27534;
assign w6899 = (~w6897 & w6887) | (~w6897 & w27535) | (w6887 & w27535);
assign w6900 = ~w6898 & ~w6899;
assign w6901 = ~w6705 & w6900;
assign w6902 = w6705 & ~w6900;
assign w6903 = ~w6901 & ~w6902;
assign w6904 = ~w6704 & w6903;
assign w6905 = w6903 & ~w6904;
assign w6906 = ~w6903 & ~w6704;
assign w6907 = ~w6905 & ~w6906;
assign w6908 = (~w6613 & w6616) | (~w6613 & w28903) | (w6616 & w28903);
assign w6909 = w6907 & w6908;
assign w6910 = ~w6907 & ~w6908;
assign w6911 = ~w6909 & ~w6910;
assign w6912 = b_37 & w418;
assign w6913 = w481 & w28904;
assign w6914 = b_36 & w413;
assign w6915 = ~w6913 & ~w6914;
assign w6916 = ~w6912 & w6915;
assign w6917 = (w6916 & ~w4636) | (w6916 & w28905) | (~w4636 & w28905);
assign w6918 = (w4636 & w39319) | (w4636 & w39320) | (w39319 & w39320);
assign w6919 = (~w4636 & w39321) | (~w4636 & w39322) | (w39321 & w39322);
assign w6920 = ~w6917 & ~w6918;
assign w6921 = ~w6919 & ~w6920;
assign w6922 = w6911 & ~w6921;
assign w6923 = w6911 & ~w6922;
assign w6924 = ~w6911 & ~w6921;
assign w6925 = ~w6923 & ~w6924;
assign w6926 = (~w6630 & w6422) | (~w6630 & w27736) | (w6422 & w27736);
assign w6927 = w6925 & w6926;
assign w6928 = ~w6925 & ~w6926;
assign w6929 = ~w6927 & ~w6928;
assign w6930 = b_40 & w239;
assign w6931 = w266 & w28906;
assign w6932 = b_39 & w234;
assign w6933 = ~w6931 & ~w6932;
assign w6934 = ~w6930 & w6933;
assign w6935 = (w6934 & ~w5363) | (w6934 & w28907) | (~w5363 & w28907);
assign w6936 = (w5363 & w39323) | (w5363 & w39324) | (w39323 & w39324);
assign w6937 = (~w5363 & w39325) | (~w5363 & w39326) | (w39325 & w39326);
assign w6938 = ~w6935 & ~w6936;
assign w6939 = ~w6937 & ~w6938;
assign w6940 = w6929 & ~w6939;
assign w6941 = ~w6929 & w6939;
assign w6942 = (~w28908 & w39327) | (~w28908 & w39328) | (w39327 & w39328);
assign w6943 = (~w28908 & w39329) | (~w28908 & w39330) | (w39329 & w39330);
assign w6944 = ~w28908 & w39331;
assign w6945 = ~w6942 & ~w6944;
assign w6946 = b_43 & w99;
assign w6947 = w136 & w28909;
assign w6948 = b_42 & w94;
assign w6949 = ~w6947 & ~w6948;
assign w6950 = ~w6946 & w6949;
assign w6951 = (w6950 & ~w5888) | (w6950 & w28910) | (~w5888 & w28910);
assign w6952 = (w5888 & w39332) | (w5888 & w39333) | (w39332 & w39333);
assign w6953 = (~w5888 & w39334) | (~w5888 & w39335) | (w39334 & w39335);
assign w6954 = ~w6951 & ~w6952;
assign w6955 = ~w6953 & ~w6954;
assign w6956 = ~w6945 & ~w6955;
assign w6957 = ~w6945 & ~w6956;
assign w6958 = w6945 & ~w6955;
assign w6959 = ~w6957 & ~w6958;
assign w6960 = (~w6664 & w6667) | (~w6664 & w39336) | (w6667 & w39336);
assign w6961 = w6959 & w6960;
assign w6962 = ~w6959 & ~w6960;
assign w6963 = ~w6961 & ~w6962;
assign w6964 = w8 & w28911;
assign w6965 = ~w8 & w28912;
assign w6966 = b_45 & w4;
assign w6967 = ~w6965 & ~w6966;
assign w6968 = ~w6964 & w6967;
assign w6969 = ~b_45 & ~b_46;
assign w6970 = b_45 & b_46;
assign w6971 = ~w6969 & ~w6970;
assign w6972 = (w4656 & w39337) | (w4656 & w39338) | (w39337 & w39338);
assign w6973 = (~w4656 & w39339) | (~w4656 & w39340) | (w39339 & w39340);
assign w6974 = ~w6972 & ~w6973;
assign w6975 = (w6968 & ~w6974) | (w6968 & w28919) | (~w6974 & w28919);
assign w6976 = (w6974 & w39341) | (w6974 & w39342) | (w39341 & w39342);
assign w6977 = (~w6974 & w39343) | (~w6974 & w39344) | (w39343 & w39344);
assign w6978 = ~w6975 & ~w6976;
assign w6979 = ~w6977 & ~w6978;
assign w6980 = w6963 & ~w6979;
assign w6981 = w6963 & ~w6980;
assign w6982 = ~w6963 & ~w6979;
assign w6983 = ~w6981 & ~w6982;
assign w6984 = (~w25050 & w28920) | (~w25050 & w28921) | (w28920 & w28921);
assign w6985 = ~w6983 & ~w6984;
assign w6986 = w6983 & w6984;
assign w6987 = ~w6985 & ~w6986;
assign w6988 = w8 & w28922;
assign w6989 = ~w8 & w28923;
assign w6990 = b_46 & w4;
assign w6991 = ~w6989 & ~w6990;
assign w6992 = ~w6988 & w6991;
assign w6993 = ~b_46 & ~b_47;
assign w6994 = b_46 & b_47;
assign w6995 = ~w6993 & ~w6994;
assign w6996 = (w4656 & w39345) | (w4656 & w39346) | (w39345 & w39346);
assign w6997 = (~w4656 & w39347) | (~w4656 & w39348) | (w39347 & w39348);
assign w6998 = ~w6996 & ~w6997;
assign w6999 = (w6992 & ~w6998) | (w6992 & w28930) | (~w6998 & w28930);
assign w7000 = (w6998 & w39349) | (w6998 & w39350) | (w39349 & w39350);
assign w7001 = (~w6998 & w39351) | (~w6998 & w39352) | (w39351 & w39352);
assign w7002 = ~w6999 & ~w7000;
assign w7003 = ~w7001 & ~w7002;
assign w7004 = (~w6956 & w6959) | (~w6956 & w39353) | (w6959 & w39353);
assign w7005 = b_35 & w657;
assign w7006 = w754 & w28931;
assign w7007 = b_34 & w652;
assign w7008 = ~w7006 & ~w7007;
assign w7009 = ~w7005 & w7008;
assign w7010 = (w7009 & ~w4181) | (w7009 & w28932) | (~w4181 & w28932);
assign w7011 = (w4181 & w39354) | (w4181 & w39355) | (w39354 & w39355);
assign w7012 = (~w4181 & w39356) | (~w4181 & w39357) | (w39356 & w39357);
assign w7013 = ~w7010 & ~w7011;
assign w7014 = ~w7012 & ~w7013;
assign w7015 = ~w6899 & ~w6901;
assign w7016 = b_32 & w986;
assign w7017 = w1069 & w28933;
assign w7018 = b_31 & w981;
assign w7019 = ~w7017 & ~w7018;
assign w7020 = ~w7016 & w7019;
assign w7021 = (w7020 & ~w3545) | (w7020 & w28934) | (~w3545 & w28934);
assign w7022 = (w3545 & w39358) | (w3545 & w39359) | (w39358 & w39359);
assign w7023 = (~w3545 & w39360) | (~w3545 & w39361) | (w39360 & w39361);
assign w7024 = ~w7021 & ~w7022;
assign w7025 = ~w7023 & ~w7024;
assign w7026 = (~w6882 & w6885) | (~w6882 & w27536) | (w6885 & w27536);
assign w7027 = b_29 & w1295;
assign w7028 = w1422 & w28935;
assign w7029 = b_28 & w1290;
assign w7030 = ~w7028 & ~w7029;
assign w7031 = ~w7027 & w7030;
assign w7032 = (w7031 & ~w2954) | (w7031 & w28936) | (~w2954 & w28936);
assign w7033 = (w2954 & w39362) | (w2954 & w39363) | (w39362 & w39363);
assign w7034 = (~w2954 & w39364) | (~w2954 & w39365) | (w39364 & w39365);
assign w7035 = ~w7032 & ~w7033;
assign w7036 = ~w7034 & ~w7035;
assign w7037 = (~w6874 & w6877) | (~w6874 & w27537) | (w6877 & w27537);
assign w7038 = (~w6856 & w6860) | (~w6856 & w25053) | (w6860 & w25053);
assign w7039 = (~w6820 & w6824) | (~w6820 & w25054) | (w6824 & w25054);
assign w7040 = b_17 & w3195;
assign w7041 = w3388 & w28937;
assign w7042 = b_16 & w3190;
assign w7043 = ~w7041 & ~w7042;
assign w7044 = ~w7040 & w7043;
assign w7045 = (w7044 & ~w1038) | (w7044 & w28938) | (~w1038 & w28938);
assign w7046 = (w1038 & w39366) | (w1038 & w39367) | (w39366 & w39367);
assign w7047 = (~w1038 & w39368) | (~w1038 & w39369) | (w39368 & w39369);
assign w7048 = ~w7045 & ~w7046;
assign w7049 = ~w7047 & ~w7048;
assign w7050 = (~w6815 & w6727) | (~w6815 & w27035) | (w6727 & w27035);
assign w7051 = b_14 & w3803;
assign w7052 = w4027 & w28939;
assign w7053 = b_13 & w3798;
assign w7054 = ~w7052 & ~w7053;
assign w7055 = ~w7051 & w7054;
assign w7056 = (w7055 & ~w735) | (w7055 & w28940) | (~w735 & w28940);
assign w7057 = (w735 & w39370) | (w735 & w39371) | (w39370 & w39371);
assign w7058 = (~w735 & w39372) | (~w735 & w39373) | (w39372 & w39373);
assign w7059 = ~w7056 & ~w7057;
assign w7060 = ~w7058 & ~w7059;
assign w7061 = (~w6779 & w6783) | (~w6779 & w28941) | (w6783 & w28941);
assign w7062 = b_8 & w5196;
assign w7063 = w5459 & w28942;
assign w7064 = b_7 & w5191;
assign w7065 = ~w7063 & ~w7064;
assign w7066 = ~w7062 & w7065;
assign w7067 = ~w308 & w28943;
assign w7068 = (w7066 & ~w28943) | (w7066 & w39374) | (~w28943 & w39374);
assign w7069 = (w28943 & w39375) | (w28943 & w39376) | (w39375 & w39376);
assign w7070 = ~w7067 & w28945;
assign w7071 = ~w7068 & ~w7069;
assign w7072 = ~w7070 & ~w7071;
assign w7073 = (~w6774 & w6740) | (~w6774 & w26154) | (w6740 & w26154);
assign w7074 = b_2 & w6761;
assign w7075 = w6482 & ~w6760;
assign w7076 = w7075 & w25553;
assign w7077 = b_1 & w6756;
assign w7078 = ~w7076 & ~w7077;
assign w7079 = ~w7074 & w7078;
assign w7080 = w35 & w6764;
assign w7081 = w7079 & ~w7080;
assign w7082 = (a_47 & ~w7079) | (a_47 & w25808) | (~w7079 & w25808);
assign w7083 = w7079 & w26155;
assign w7084 = ~w7081 & ~w7082;
assign w7085 = ~w7083 & ~w7084;
assign w7086 = ~w6770 & w7085;
assign w7087 = w6770 & ~w7085;
assign w7088 = ~w7086 & ~w7087;
assign w7089 = b_5 & w5962;
assign w7090 = w6246 & w26788;
assign w7091 = b_4 & w5957;
assign w7092 = ~w7090 & ~w7091;
assign w7093 = ~w7089 & w7092;
assign w7094 = w129 & w5965;
assign w7095 = w7093 & ~w7094;
assign w7096 = (a_44 & w7094) | (a_44 & w26789) | (w7094 & w26789);
assign w7097 = ~w7094 & w39377;
assign w7098 = ~w7095 & ~w7096;
assign w7099 = ~w7097 & ~w7098;
assign w7100 = w7088 & ~w7099;
assign w7101 = w7088 & ~w7100;
assign w7102 = ~w7088 & ~w7099;
assign w7103 = ~w7101 & ~w7102;
assign w7104 = ~w7073 & ~w7103;
assign w7105 = w7073 & w7103;
assign w7106 = ~w7104 & ~w7105;
assign w7107 = ~w7072 & w7106;
assign w7108 = ~w7106 & ~w7072;
assign w7109 = w7106 & ~w7107;
assign w7110 = ~w7108 & ~w7109;
assign w7111 = ~w7061 & ~w7110;
assign w7112 = ~w7061 & ~w7111;
assign w7113 = b_11 & w4499;
assign w7114 = w4723 & w28946;
assign w7115 = b_10 & w4494;
assign w7116 = ~w7114 & ~w7115;
assign w7117 = ~w7113 & w7116;
assign w7118 = (w7117 & ~w530) | (w7117 & w28947) | (~w530 & w28947);
assign w7119 = (w530 & w39378) | (w530 & w39379) | (w39378 & w39379);
assign w7120 = (~w530 & w39380) | (~w530 & w39381) | (w39380 & w39381);
assign w7121 = ~w7118 & ~w7119;
assign w7122 = ~w7120 & ~w7121;
assign w7123 = ~w7112 & w26907;
assign w7124 = (~w7122 & w7112) | (~w7122 & w26908) | (w7112 & w26908);
assign w7125 = ~w7123 & ~w7124;
assign w7126 = ~w6801 & w7125;
assign w7127 = w6801 & ~w7125;
assign w7128 = ~w7126 & ~w7127;
assign w7129 = ~w7060 & w7128;
assign w7130 = w7128 & ~w7129;
assign w7131 = ~w7128 & ~w7060;
assign w7132 = ~w7130 & ~w7131;
assign w7133 = ~w7050 & ~w7132;
assign w7134 = w7050 & w7132;
assign w7135 = ~w7133 & ~w7134;
assign w7136 = ~w7049 & w7135;
assign w7137 = ~w7135 & ~w7049;
assign w7138 = w7135 & ~w7136;
assign w7139 = ~w7137 & ~w7138;
assign w7140 = w7139 & ~w7039;
assign w7141 = w7039 & ~w7139;
assign w7142 = ~w7140 & ~w7141;
assign w7143 = b_20 & w2639;
assign w7144 = w2820 & w28948;
assign w7145 = b_19 & w2634;
assign w7146 = ~w7144 & ~w7145;
assign w7147 = ~w7143 & w7146;
assign w7148 = (w7147 & ~w1503) | (w7147 & w28949) | (~w1503 & w28949);
assign w7149 = (w1503 & w39382) | (w1503 & w39383) | (w39382 & w39383);
assign w7150 = (~w1503 & w39384) | (~w1503 & w39385) | (w39384 & w39385);
assign w7151 = ~w7148 & ~w7149;
assign w7152 = ~w7150 & ~w7151;
assign w7153 = (~w7152 & w7140) | (~w7152 & w27143) | (w7140 & w27143);
assign w7154 = ~w7142 & ~w7153;
assign w7155 = ~w27143 & w28950;
assign w7156 = ~w7154 & ~w7155;
assign w7157 = (~w6838 & w6841) | (~w6838 & w27226) | (w6841 & w27226);
assign w7158 = w7156 & w7157;
assign w7159 = ~w7156 & ~w7157;
assign w7160 = ~w7158 & ~w7159;
assign w7161 = b_23 & w2158;
assign w7162 = w2294 & w28951;
assign w7163 = b_22 & w2153;
assign w7164 = ~w7162 & ~w7163;
assign w7165 = ~w7161 & w7164;
assign w7166 = (w7165 & ~w1933) | (w7165 & w28952) | (~w1933 & w28952);
assign w7167 = (w1933 & w39386) | (w1933 & w39387) | (w39386 & w39387);
assign w7168 = (~w1933 & w39388) | (~w1933 & w39389) | (w39388 & w39389);
assign w7169 = ~w7166 & ~w7167;
assign w7170 = ~w7168 & ~w7169;
assign w7171 = w7160 & ~w7170;
assign w7172 = ~w7160 & w7170;
assign w7173 = ~w7038 & w25055;
assign w7174 = ~w7038 & ~w7173;
assign w7175 = (~w7171 & w7038) | (~w7171 & w27227) | (w7038 & w27227);
assign w7176 = (w27227 & w25055) | (w27227 & w28953) | (w25055 & w28953);
assign w7177 = ~w7174 & ~w7176;
assign w7178 = b_26 & w1694;
assign w7179 = w1834 & w28954;
assign w7180 = b_25 & w1689;
assign w7181 = ~w7179 & ~w7180;
assign w7182 = ~w7178 & w7181;
assign w7183 = (w7182 & ~w2416) | (w7182 & w28955) | (~w2416 & w28955);
assign w7184 = (w2416 & w39390) | (w2416 & w39391) | (w39390 & w39391);
assign w7185 = (~w2416 & w39392) | (~w2416 & w39393) | (w39392 & w39393);
assign w7186 = ~w7183 & ~w7184;
assign w7187 = ~w7185 & ~w7186;
assign w7188 = w7177 & w7187;
assign w7189 = ~w7177 & ~w7187;
assign w7190 = ~w7188 & ~w7189;
assign w7191 = ~w7037 & w7190;
assign w7192 = w7037 & ~w7190;
assign w7193 = ~w7191 & ~w7192;
assign w7194 = w7036 & ~w7193;
assign w7195 = ~w7036 & w7193;
assign w7196 = ~w7194 & ~w7195;
assign w7197 = (w7196 & w6886) | (w7196 & w25056) | (w6886 & w25056);
assign w7198 = w7026 & ~w7196;
assign w7199 = ~w7197 & ~w7198;
assign w7200 = w7025 & ~w7199;
assign w7201 = ~w7025 & w7199;
assign w7202 = ~w7200 & ~w7201;
assign w7203 = ~w7015 & w7202;
assign w7204 = w7015 & ~w7202;
assign w7205 = ~w7203 & ~w7204;
assign w7206 = ~w7014 & w7205;
assign w7207 = w7205 & ~w7206;
assign w7208 = ~w7205 & ~w7014;
assign w7209 = ~w7207 & ~w7208;
assign w7210 = ~w6904 & ~w6910;
assign w7211 = w7209 & w7210;
assign w7212 = ~w7209 & ~w7210;
assign w7213 = ~w7211 & ~w7212;
assign w7214 = b_38 & w418;
assign w7215 = w481 & w28956;
assign w7216 = b_37 & w413;
assign w7217 = ~w7215 & ~w7216;
assign w7218 = ~w7214 & w7217;
assign w7219 = (w7218 & ~w4658) | (w7218 & w25057) | (~w4658 & w25057);
assign w7220 = (w4658 & w28957) | (w4658 & w28958) | (w28957 & w28958);
assign w7221 = (~w4658 & w28959) | (~w4658 & w28960) | (w28959 & w28960);
assign w7222 = ~w7219 & ~w7220;
assign w7223 = ~w7221 & ~w7222;
assign w7224 = w7213 & ~w7223;
assign w7225 = w7213 & ~w7224;
assign w7226 = ~w7213 & ~w7223;
assign w7227 = ~w7225 & ~w7226;
assign w7228 = (~w6922 & w6925) | (~w6922 & w27737) | (w6925 & w27737);
assign w7229 = w7227 & w7228;
assign w7230 = ~w7227 & ~w7228;
assign w7231 = ~w7229 & ~w7230;
assign w7232 = b_41 & w239;
assign w7233 = w266 & w28961;
assign w7234 = b_40 & w234;
assign w7235 = ~w7233 & ~w7234;
assign w7236 = ~w7232 & w7235;
assign w7237 = (w7236 & ~w5609) | (w7236 & w28962) | (~w5609 & w28962);
assign w7238 = (w5609 & w39394) | (w5609 & w39395) | (w39394 & w39395);
assign w7239 = (~w5609 & w39396) | (~w5609 & w39397) | (w39396 & w39397);
assign w7240 = ~w7237 & ~w7238;
assign w7241 = ~w7239 & ~w7240;
assign w7242 = w7231 & ~w7241;
assign w7243 = ~w7231 & w7241;
assign w7244 = ~w6943 & w25058;
assign w7245 = ~w6943 & ~w7244;
assign w7246 = (~w7242 & w6943) | (~w7242 & w28963) | (w6943 & w28963);
assign w7247 = (w28963 & w25058) | (w28963 & w39398) | (w25058 & w39398);
assign w7248 = ~w7245 & ~w7247;
assign w7249 = b_44 & w99;
assign w7250 = w136 & w28964;
assign w7251 = b_43 & w94;
assign w7252 = ~w7250 & ~w7251;
assign w7253 = ~w7249 & w7252;
assign w7254 = (w7253 & ~w6408) | (w7253 & w28965) | (~w6408 & w28965);
assign w7255 = (w6408 & w39399) | (w6408 & w39400) | (w39399 & w39400);
assign w7256 = (~w6408 & w39401) | (~w6408 & w39402) | (w39401 & w39402);
assign w7257 = ~w7254 & ~w7255;
assign w7258 = ~w7256 & ~w7257;
assign w7259 = w7248 & w7258;
assign w7260 = ~w7248 & ~w7258;
assign w7261 = ~w7259 & ~w7260;
assign w7262 = (w7261 & w6962) | (w7261 & w25059) | (w6962 & w25059);
assign w7263 = w7004 & ~w7261;
assign w7264 = ~w7262 & ~w7263;
assign w7265 = ~w7262 & w39403;
assign w7266 = w7264 & ~w7265;
assign w7267 = (~w7003 & w7262) | (~w7003 & w39404) | (w7262 & w39404);
assign w7268 = ~w7266 & ~w7267;
assign w7269 = (~w6980 & w6983) | (~w6980 & w28966) | (w6983 & w28966);
assign w7270 = ~w7268 & ~w7269;
assign w7271 = w7268 & w7269;
assign w7272 = ~w7270 & ~w7271;
assign w7273 = (~w7265 & w7268) | (~w7265 & w28967) | (w7268 & w28967);
assign w7274 = w8 & w28968;
assign w7275 = ~w8 & w28969;
assign w7276 = b_47 & w4;
assign w7277 = ~w7275 & ~w7276;
assign w7278 = ~w7274 & w7277;
assign w7279 = ~b_47 & ~b_48;
assign w7280 = b_47 & b_48;
assign w7281 = ~w7279 & ~w7280;
assign w7282 = (w4656 & w39405) | (w4656 & w39406) | (w39405 & w39406);
assign w7283 = (~w4656 & w39407) | (~w4656 & w39408) | (w39407 & w39408);
assign w7284 = ~w7282 & ~w7283;
assign w7285 = (w7278 & ~w7284) | (w7278 & w28976) | (~w7284 & w28976);
assign w7286 = (w7284 & w39409) | (w7284 & w39410) | (w39409 & w39410);
assign w7287 = (~w7284 & w39411) | (~w7284 & w39412) | (w39411 & w39412);
assign w7288 = ~w7285 & ~w7286;
assign w7289 = ~w7287 & ~w7288;
assign w7290 = (~w25059 & w28977) | (~w25059 & w28978) | (w28977 & w28978);
assign w7291 = (~w7201 & w7015) | (~w7201 & w25061) | (w7015 & w25061);
assign w7292 = b_33 & w986;
assign w7293 = w1069 & w28979;
assign w7294 = b_32 & w981;
assign w7295 = ~w7293 & ~w7294;
assign w7296 = ~w7292 & w7295;
assign w7297 = (w7296 & ~w3744) | (w7296 & w28980) | (~w3744 & w28980);
assign w7298 = (w3744 & w39413) | (w3744 & w39414) | (w39413 & w39414);
assign w7299 = (~w3744 & w39415) | (~w3744 & w39416) | (w39415 & w39416);
assign w7300 = ~w7297 & ~w7298;
assign w7301 = ~w7299 & ~w7300;
assign w7302 = (~w7189 & w7037) | (~w7189 & w25062) | (w7037 & w25062);
assign w7303 = b_27 & w1694;
assign w7304 = w1834 & w28981;
assign w7305 = b_26 & w1689;
assign w7306 = ~w7304 & ~w7305;
assign w7307 = ~w7303 & w7306;
assign w7308 = (w7307 & ~w2582) | (w7307 & w28982) | (~w2582 & w28982);
assign w7309 = (w2582 & w39417) | (w2582 & w39418) | (w39417 & w39418);
assign w7310 = (~w2582 & w39419) | (~w2582 & w39420) | (w39419 & w39420);
assign w7311 = ~w7308 & ~w7309;
assign w7312 = ~w7310 & ~w7311;
assign w7313 = ~w7129 & ~w7133;
assign w7314 = b_15 & w3803;
assign w7315 = w4027 & w28983;
assign w7316 = b_14 & w3798;
assign w7317 = ~w7315 & ~w7316;
assign w7318 = ~w7314 & w7317;
assign w7319 = (w7318 & ~w827) | (w7318 & w28984) | (~w827 & w28984);
assign w7320 = (w827 & w39421) | (w827 & w39422) | (w39421 & w39422);
assign w7321 = (~w827 & w39423) | (~w827 & w39424) | (w39423 & w39424);
assign w7322 = ~w7319 & ~w7320;
assign w7323 = ~w7321 & ~w7322;
assign w7324 = (~w7124 & w6801) | (~w7124 & w28985) | (w6801 & w28985);
assign w7325 = b_12 & w4499;
assign w7326 = w4723 & w28986;
assign w7327 = b_11 & w4494;
assign w7328 = ~w7326 & ~w7327;
assign w7329 = ~w7325 & w7328;
assign w7330 = (w7329 & ~w552) | (w7329 & w28987) | (~w552 & w28987);
assign w7331 = (w552 & w39425) | (w552 & w39426) | (w39425 & w39426);
assign w7332 = (~w552 & w39427) | (~w552 & w39428) | (w39427 & w39428);
assign w7333 = ~w7330 & ~w7331;
assign w7334 = ~w7332 & ~w7333;
assign w7335 = (~w7107 & w7061) | (~w7107 & w26559) | (w7061 & w26559);
assign w7336 = b_6 & w5962;
assign w7337 = w6246 & w28988;
assign w7338 = b_5 & w5957;
assign w7339 = ~w7337 & ~w7338;
assign w7340 = ~w7336 & w7339;
assign w7341 = (w7340 & ~w190) | (w7340 & w28989) | (~w190 & w28989);
assign w7342 = (w190 & w39429) | (w190 & w39430) | (w39429 & w39430);
assign w7343 = (~w190 & w39431) | (~w190 & w39432) | (w39431 & w39432);
assign w7344 = ~w7341 & ~w7342;
assign w7345 = ~w7343 & ~w7344;
assign w7346 = a_47 & ~a_48;
assign w7347 = ~a_47 & a_48;
assign w7348 = ~w7346 & ~w7347;
assign w7349 = b_0 & ~w7348;
assign w7350 = (w7349 & w7085) | (w7349 & w26156) | (w7085 & w26156);
assign w7351 = ~w7085 & w26157;
assign w7352 = ~w7350 & ~w7351;
assign w7353 = b_3 & w6761;
assign w7354 = w7075 & w26560;
assign w7355 = b_2 & w6756;
assign w7356 = ~w7354 & ~w7355;
assign w7357 = ~w7353 & w7356;
assign w7358 = w57 & w6764;
assign w7359 = w7357 & ~w7358;
assign w7360 = a_47 & ~w7359;
assign w7361 = w7359 & a_47;
assign w7362 = ~w7359 & ~w7360;
assign w7363 = ~w7361 & ~w7362;
assign w7364 = ~w7352 & ~w7363;
assign w7365 = w7352 & w7363;
assign w7366 = ~w7364 & ~w7365;
assign w7367 = ~w7345 & w7366;
assign w7368 = w7366 & ~w7367;
assign w7369 = ~w7366 & ~w7345;
assign w7370 = ~w7368 & ~w7369;
assign w7371 = ~w7100 & ~w7104;
assign w7372 = w7370 & w7371;
assign w7373 = ~w7370 & ~w7371;
assign w7374 = ~w7372 & ~w7373;
assign w7375 = b_9 & w5196;
assign w7376 = w5459 & w28990;
assign w7377 = b_8 & w5191;
assign w7378 = ~w7376 & ~w7377;
assign w7379 = ~w7375 & w7378;
assign w7380 = (w7379 & ~w371) | (w7379 & w28991) | (~w371 & w28991);
assign w7381 = (w371 & w39433) | (w371 & w39434) | (w39433 & w39434);
assign w7382 = (~w371 & w39435) | (~w371 & w39436) | (w39435 & w39436);
assign w7383 = ~w7380 & ~w7381;
assign w7384 = ~w7382 & ~w7383;
assign w7385 = ~w7374 & w7384;
assign w7386 = w7374 & ~w7384;
assign w7387 = ~w7385 & ~w7386;
assign w7388 = ~w7335 & w7387;
assign w7389 = w7335 & ~w7387;
assign w7390 = ~w7388 & ~w7389;
assign w7391 = ~w7334 & w7390;
assign w7392 = ~w7390 & ~w7334;
assign w7393 = w7390 & ~w7391;
assign w7394 = ~w7392 & ~w7393;
assign w7395 = (~w7394 & w7126) | (~w7394 & w26561) | (w7126 & w26561);
assign w7396 = w7324 & w7394;
assign w7397 = ~w7395 & ~w7396;
assign w7398 = ~w7323 & w7397;
assign w7399 = w7323 & ~w7397;
assign w7400 = ~w7398 & ~w7399;
assign w7401 = (w7400 & w7133) | (w7400 & w28992) | (w7133 & w28992);
assign w7402 = ~w7133 & w28993;
assign w7403 = ~w7401 & ~w7402;
assign w7404 = b_18 & w3195;
assign w7405 = w3388 & w28994;
assign w7406 = b_17 & w3190;
assign w7407 = ~w7405 & ~w7406;
assign w7408 = ~w7404 & w7407;
assign w7409 = (w7408 & ~w1238) | (w7408 & w28995) | (~w1238 & w28995);
assign w7410 = (w1238 & w39437) | (w1238 & w39438) | (w39437 & w39438);
assign w7411 = (~w1238 & w39439) | (~w1238 & w39440) | (w39439 & w39440);
assign w7412 = ~w7409 & ~w7410;
assign w7413 = ~w7411 & ~w7412;
assign w7414 = w7403 & ~w7413;
assign w7415 = w7403 & ~w7414;
assign w7416 = ~w7403 & ~w7413;
assign w7417 = ~w7415 & ~w7416;
assign w7418 = (~w7136 & w7039) | (~w7136 & w27144) | (w7039 & w27144);
assign w7419 = w7417 & w7418;
assign w7420 = ~w7417 & ~w7418;
assign w7421 = ~w7419 & ~w7420;
assign w7422 = b_21 & w2639;
assign w7423 = w2820 & w28996;
assign w7424 = b_20 & w2634;
assign w7425 = ~w7423 & ~w7424;
assign w7426 = ~w7422 & w7425;
assign w7427 = (w7426 & ~w1634) | (w7426 & w28997) | (~w1634 & w28997);
assign w7428 = (w1634 & w39441) | (w1634 & w39442) | (w39441 & w39442);
assign w7429 = (~w1634 & w39443) | (~w1634 & w39444) | (w39443 & w39444);
assign w7430 = ~w7427 & ~w7428;
assign w7431 = ~w7429 & ~w7430;
assign w7432 = w7421 & ~w7431;
assign w7433 = w7421 & ~w7432;
assign w7434 = ~w7421 & ~w7431;
assign w7435 = ~w7433 & ~w7434;
assign w7436 = (~w7153 & w7156) | (~w7153 & w27228) | (w7156 & w27228);
assign w7437 = w7435 & w7436;
assign w7438 = ~w7435 & ~w7436;
assign w7439 = ~w7437 & ~w7438;
assign w7440 = b_24 & w2158;
assign w7441 = w2294 & w28998;
assign w7442 = b_23 & w2153;
assign w7443 = ~w7441 & ~w7442;
assign w7444 = ~w7440 & w7443;
assign w7445 = (w7444 & ~w2083) | (w7444 & w28999) | (~w2083 & w28999);
assign w7446 = (w2083 & w39445) | (w2083 & w39446) | (w39445 & w39446);
assign w7447 = (~w2083 & w39447) | (~w2083 & w39448) | (w39447 & w39448);
assign w7448 = ~w7445 & ~w7446;
assign w7449 = ~w7447 & ~w7448;
assign w7450 = ~w7439 & w7449;
assign w7451 = w7439 & ~w7449;
assign w7452 = ~w7450 & ~w7451;
assign w7453 = ~w7175 & w7452;
assign w7454 = w7175 & ~w7452;
assign w7455 = ~w7453 & ~w7454;
assign w7456 = ~w7312 & w7455;
assign w7457 = w7455 & ~w7456;
assign w7458 = ~w7455 & ~w7312;
assign w7459 = ~w7457 & ~w7458;
assign w7460 = ~w7302 & w7459;
assign w7461 = w7302 & ~w7459;
assign w7462 = ~w7460 & ~w7461;
assign w7463 = b_30 & w1295;
assign w7464 = w1422 & w29000;
assign w7465 = b_29 & w1290;
assign w7466 = ~w7464 & ~w7465;
assign w7467 = ~w7463 & w7466;
assign w7468 = (w7467 & ~w3138) | (w7467 & w29001) | (~w3138 & w29001);
assign w7469 = (w3138 & w39449) | (w3138 & w39450) | (w39449 & w39450);
assign w7470 = (~w3138 & w39451) | (~w3138 & w39452) | (w39451 & w39452);
assign w7471 = ~w7468 & ~w7469;
assign w7472 = ~w7470 & ~w7471;
assign w7473 = ~w7462 & ~w7472;
assign w7474 = w7462 & w7472;
assign w7475 = ~w7473 & ~w7474;
assign w7476 = (w7475 & w7197) | (w7475 & w26562) | (w7197 & w26562);
assign w7477 = ~w7197 & w26563;
assign w7478 = ~w7476 & ~w7477;
assign w7479 = ~w7301 & w7478;
assign w7480 = w7301 & w7478;
assign w7481 = ~w7478 & ~w7301;
assign w7482 = ~w7480 & ~w7481;
assign w7483 = ~w7291 & w7482;
assign w7484 = w7291 & ~w7482;
assign w7485 = ~w7483 & ~w7484;
assign w7486 = b_36 & w657;
assign w7487 = w754 & w29002;
assign w7488 = b_35 & w652;
assign w7489 = ~w7487 & ~w7488;
assign w7490 = ~w7486 & w7489;
assign w7491 = (w7490 & ~w4395) | (w7490 & w26564) | (~w4395 & w26564);
assign w7492 = (w4395 & w29003) | (w4395 & w29004) | (w29003 & w29004);
assign w7493 = (~w4395 & w29005) | (~w4395 & w29006) | (w29005 & w29006);
assign w7494 = ~w7491 & ~w7492;
assign w7495 = ~w7493 & ~w7494;
assign w7496 = ~w7485 & ~w7495;
assign w7497 = w7485 & w7495;
assign w7498 = ~w7496 & ~w7497;
assign w7499 = ~w7212 & w25063;
assign w7500 = (w7498 & w7212) | (w7498 & w25064) | (w7212 & w25064);
assign w7501 = ~w7499 & ~w7500;
assign w7502 = b_39 & w418;
assign w7503 = w481 & w29007;
assign w7504 = b_38 & w413;
assign w7505 = ~w7503 & ~w7504;
assign w7506 = ~w7502 & w7505;
assign w7507 = (w7506 & ~w4888) | (w7506 & w25065) | (~w4888 & w25065);
assign w7508 = (w4888 & w26565) | (w4888 & w26566) | (w26565 & w26566);
assign w7509 = (~w4888 & w29008) | (~w4888 & w29009) | (w29008 & w29009);
assign w7510 = ~w7507 & ~w7508;
assign w7511 = ~w7509 & ~w7510;
assign w7512 = w7501 & ~w7511;
assign w7513 = w7501 & ~w7512;
assign w7514 = ~w7501 & ~w7511;
assign w7515 = ~w7513 & ~w7514;
assign w7516 = (~w7224 & w7227) | (~w7224 & w27738) | (w7227 & w27738);
assign w7517 = w7515 & w7516;
assign w7518 = ~w7515 & ~w7516;
assign w7519 = ~w7517 & ~w7518;
assign w7520 = b_42 & w239;
assign w7521 = w266 & w29010;
assign w7522 = b_41 & w234;
assign w7523 = ~w7521 & ~w7522;
assign w7524 = ~w7520 & w7523;
assign w7525 = (w7524 & ~w5864) | (w7524 & w25066) | (~w5864 & w25066);
assign w7526 = (w5864 & w29011) | (w5864 & w29012) | (w29011 & w29012);
assign w7527 = (~w5864 & w29013) | (~w5864 & w29014) | (w29013 & w29014);
assign w7528 = ~w7525 & ~w7526;
assign w7529 = ~w7527 & ~w7528;
assign w7530 = w7519 & ~w7529;
assign w7531 = w7519 & ~w7530;
assign w7532 = ~w7519 & ~w7529;
assign w7533 = ~w7531 & ~w7532;
assign w7534 = ~w7246 & w7533;
assign w7535 = w7246 & ~w7533;
assign w7536 = ~w7534 & ~w7535;
assign w7537 = b_45 & w99;
assign w7538 = w136 & w29015;
assign w7539 = b_44 & w94;
assign w7540 = ~w7538 & ~w7539;
assign w7541 = ~w7537 & w7540;
assign w7542 = (w7541 & ~w6682) | (w7541 & w29016) | (~w6682 & w29016);
assign w7543 = (w6682 & w39453) | (w6682 & w39454) | (w39453 & w39454);
assign w7544 = (~w6682 & w39455) | (~w6682 & w39456) | (w39455 & w39456);
assign w7545 = ~w7542 & ~w7543;
assign w7546 = ~w7544 & ~w7545;
assign w7547 = ~w7536 & ~w7546;
assign w7548 = w7536 & w7546;
assign w7549 = ~w7547 & ~w7548;
assign w7550 = (w6962 & w27145) | (w6962 & w27146) | (w27145 & w27146);
assign w7551 = (w7289 & w7550) | (w7289 & w29017) | (w7550 & w29017);
assign w7552 = ~w7550 & w29018;
assign w7553 = ~w7551 & ~w7552;
assign w7554 = (w7553 & w7270) | (w7553 & w26568) | (w7270 & w26568);
assign w7555 = w7273 & ~w7553;
assign w7556 = ~w7554 & ~w7555;
assign w7557 = (~w26568 & w39457) | (~w26568 & w39458) | (w39457 & w39458);
assign w7558 = (~w7456 & w7302) | (~w7456 & w26569) | (w7302 & w26569);
assign w7559 = b_28 & w1694;
assign w7560 = w1834 & w29019;
assign w7561 = b_27 & w1689;
assign w7562 = ~w7560 & ~w7561;
assign w7563 = ~w7559 & w7562;
assign w7564 = (w7563 & ~w2771) | (w7563 & w29020) | (~w2771 & w29020);
assign w7565 = (w2771 & w39459) | (w2771 & w39460) | (w39459 & w39460);
assign w7566 = (~w2771 & w39461) | (~w2771 & w39462) | (w39461 & w39462);
assign w7567 = ~w7564 & ~w7565;
assign w7568 = ~w7566 & ~w7567;
assign w7569 = b_16 & w3803;
assign w7570 = w4027 & w29021;
assign w7571 = b_15 & w3798;
assign w7572 = ~w7570 & ~w7571;
assign w7573 = ~w7569 & w7572;
assign w7574 = (w7573 & ~w926) | (w7573 & w29022) | (~w926 & w29022);
assign w7575 = (w926 & w39463) | (w926 & w39464) | (w39463 & w39464);
assign w7576 = (~w926 & w39465) | (~w926 & w39466) | (w39465 & w39466);
assign w7577 = ~w7574 & ~w7575;
assign w7578 = ~w7576 & ~w7577;
assign w7579 = (~w26561 & w26790) | (~w26561 & w26791) | (w26790 & w26791);
assign w7580 = (~w7386 & w7335) | (~w7386 & w26570) | (w7335 & w26570);
assign w7581 = b_7 & w5962;
assign w7582 = w6246 & w29023;
assign w7583 = b_6 & w5957;
assign w7584 = ~w7582 & ~w7583;
assign w7585 = ~w7581 & w7584;
assign w7586 = (w7585 & ~w213) | (w7585 & w29024) | (~w213 & w29024);
assign w7587 = (w213 & w39467) | (w213 & w39468) | (w39467 & w39468);
assign w7588 = (~w213 & w39469) | (~w213 & w39470) | (w39469 & w39470);
assign w7589 = ~w7586 & ~w7587;
assign w7590 = ~w7588 & ~w7589;
assign w7591 = ~w7085 & w29025;
assign w7592 = (~w7591 & w7352) | (~w7591 & w29026) | (w7352 & w29026);
assign w7593 = b_4 & w6761;
assign w7594 = w7075 & w26571;
assign w7595 = b_3 & w6756;
assign w7596 = ~w7594 & ~w7595;
assign w7597 = ~w7593 & w7596;
assign w7598 = w84 & w6764;
assign w7599 = w7597 & ~w7598;
assign w7600 = (a_47 & w7598) | (a_47 & w26572) | (w7598 & w26572);
assign w7601 = ~w7598 & w27419;
assign w7602 = ~w7599 & ~w7600;
assign w7603 = ~w7601 & ~w7602;
assign w7604 = (a_50 & w7348) | (a_50 & w29027) | (w7348 & w29027);
assign w7605 = ~a_48 & a_49;
assign w7606 = a_48 & ~a_49;
assign w7607 = ~w7605 & ~w7606;
assign w7608 = w7348 & ~w7607;
assign w7609 = b_0 & w7608;
assign w7610 = ~a_49 & a_50;
assign w7611 = a_49 & ~a_50;
assign w7612 = ~w7610 & ~w7611;
assign w7613 = ~w7348 & w7612;
assign w7614 = b_1 & w7613;
assign w7615 = ~w7609 & ~w7614;
assign w7616 = ~w7348 & ~w7612;
assign w7617 = ~w15 & w7616;
assign w7618 = w7615 & ~w7617;
assign w7619 = (a_50 & ~w7615) | (a_50 & w25554) | (~w7615 & w25554);
assign w7620 = w7615 & w25809;
assign w7621 = ~w7618 & ~w7619;
assign w7622 = (w7604 & w7621) | (w7604 & w25810) | (w7621 & w25810);
assign w7623 = ~w7621 & w27147;
assign w7624 = ~w7622 & ~w7623;
assign w7625 = w7603 & ~w7624;
assign w7626 = ~w7603 & w7624;
assign w7627 = ~w7625 & ~w7626;
assign w7628 = ~w7592 & w7627;
assign w7629 = w7592 & ~w7627;
assign w7630 = ~w7628 & ~w7629;
assign w7631 = ~w7590 & w7630;
assign w7632 = w7630 & ~w7631;
assign w7633 = ~w7630 & ~w7590;
assign w7634 = ~w7632 & ~w7633;
assign w7635 = ~w7367 & ~w7373;
assign w7636 = w7634 & w7635;
assign w7637 = ~w7634 & ~w7635;
assign w7638 = ~w7636 & ~w7637;
assign w7639 = b_10 & w5196;
assign w7640 = w5459 & w29028;
assign w7641 = b_9 & w5191;
assign w7642 = ~w7640 & ~w7641;
assign w7643 = ~w7639 & w7642;
assign w7644 = (w7643 & ~w454) | (w7643 & w29029) | (~w454 & w29029);
assign w7645 = (w454 & w39471) | (w454 & w39472) | (w39471 & w39472);
assign w7646 = (~w454 & w39473) | (~w454 & w39474) | (w39473 & w39474);
assign w7647 = ~w7644 & ~w7645;
assign w7648 = ~w7646 & ~w7647;
assign w7649 = w7638 & ~w7648;
assign w7650 = ~w7638 & w7648;
assign w7651 = ~w7580 & w26792;
assign w7652 = ~w7580 & ~w7651;
assign w7653 = ~w7649 & ~w7651;
assign w7654 = ~w7651 & w26792;
assign w7655 = ~w7652 & ~w7654;
assign w7656 = b_13 & w4499;
assign w7657 = w4723 & w29030;
assign w7658 = b_12 & w4494;
assign w7659 = ~w7657 & ~w7658;
assign w7660 = ~w7656 & w7659;
assign w7661 = (w7660 & ~w711) | (w7660 & w29031) | (~w711 & w29031);
assign w7662 = (w711 & w39475) | (w711 & w39476) | (w39475 & w39476);
assign w7663 = (~w711 & w39477) | (~w711 & w39478) | (w39477 & w39478);
assign w7664 = ~w7661 & ~w7662;
assign w7665 = ~w7663 & ~w7664;
assign w7666 = w7655 & w7665;
assign w7667 = ~w7655 & ~w7665;
assign w7668 = ~w7666 & ~w7667;
assign w7669 = ~w7579 & w7668;
assign w7670 = w7579 & ~w7668;
assign w7671 = ~w7669 & ~w7670;
assign w7672 = ~w7578 & w7671;
assign w7673 = w7671 & ~w7672;
assign w7674 = ~w7671 & ~w7578;
assign w7675 = ~w7673 & ~w7674;
assign w7676 = (~w7398 & w7313) | (~w7398 & w26573) | (w7313 & w26573);
assign w7677 = w7675 & w7676;
assign w7678 = ~w7675 & ~w7676;
assign w7679 = ~w7677 & ~w7678;
assign w7680 = b_19 & w3195;
assign w7681 = w3388 & w29032;
assign w7682 = b_18 & w3190;
assign w7683 = ~w7681 & ~w7682;
assign w7684 = ~w7680 & w7683;
assign w7685 = (w7684 & ~w1372) | (w7684 & w29033) | (~w1372 & w29033);
assign w7686 = (w1372 & w39479) | (w1372 & w39480) | (w39479 & w39480);
assign w7687 = (~w1372 & w39481) | (~w1372 & w39482) | (w39481 & w39482);
assign w7688 = ~w7685 & ~w7686;
assign w7689 = ~w7687 & ~w7688;
assign w7690 = w7679 & ~w7689;
assign w7691 = w7679 & ~w7690;
assign w7692 = ~w7679 & ~w7689;
assign w7693 = ~w7691 & ~w7692;
assign w7694 = (~w7414 & w7417) | (~w7414 & w27344) | (w7417 & w27344);
assign w7695 = w7693 & w7694;
assign w7696 = ~w7693 & ~w7694;
assign w7697 = ~w7695 & ~w7696;
assign w7698 = b_22 & w2639;
assign w7699 = w2820 & w29034;
assign w7700 = b_21 & w2634;
assign w7701 = ~w7699 & ~w7700;
assign w7702 = ~w7698 & w7701;
assign w7703 = (w7702 & ~w1786) | (w7702 & w29035) | (~w1786 & w29035);
assign w7704 = (w1786 & w39483) | (w1786 & w39484) | (w39483 & w39484);
assign w7705 = (~w1786 & w39485) | (~w1786 & w39486) | (w39485 & w39486);
assign w7706 = ~w7703 & ~w7704;
assign w7707 = ~w7705 & ~w7706;
assign w7708 = w7697 & ~w7707;
assign w7709 = w7697 & ~w7708;
assign w7710 = ~w7697 & ~w7707;
assign w7711 = ~w7709 & ~w7710;
assign w7712 = (~w7432 & w7436) | (~w7432 & w26574) | (w7436 & w26574);
assign w7713 = w7711 & w7712;
assign w7714 = ~w7711 & ~w7712;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = b_25 & w2158;
assign w7717 = w2294 & w29036;
assign w7718 = b_24 & w2153;
assign w7719 = ~w7717 & ~w7718;
assign w7720 = ~w7716 & w7719;
assign w7721 = (w7720 & ~w2108) | (w7720 & w29037) | (~w2108 & w29037);
assign w7722 = (w2108 & w39487) | (w2108 & w39488) | (w39487 & w39488);
assign w7723 = (~w2108 & w39489) | (~w2108 & w39490) | (w39489 & w39490);
assign w7724 = ~w7721 & ~w7722;
assign w7725 = ~w7723 & ~w7724;
assign w7726 = w7715 & ~w7725;
assign w7727 = w7715 & ~w7726;
assign w7728 = ~w7715 & ~w7725;
assign w7729 = ~w7727 & ~w7728;
assign w7730 = (~w7451 & w7175) | (~w7451 & w26575) | (w7175 & w26575);
assign w7731 = ~w7729 & ~w7730;
assign w7732 = w7729 & w7730;
assign w7733 = ~w7731 & ~w7732;
assign w7734 = ~w7568 & w7733;
assign w7735 = ~w7733 & ~w7568;
assign w7736 = w7733 & ~w7734;
assign w7737 = ~w7735 & ~w7736;
assign w7738 = w7737 & ~w7558;
assign w7739 = w7558 & ~w7737;
assign w7740 = ~w7738 & ~w7739;
assign w7741 = b_31 & w1295;
assign w7742 = w1422 & w29038;
assign w7743 = b_30 & w1290;
assign w7744 = ~w7742 & ~w7743;
assign w7745 = ~w7741 & w7744;
assign w7746 = (w7745 & ~w3345) | (w7745 & w29039) | (~w3345 & w29039);
assign w7747 = (w3345 & w39491) | (w3345 & w39492) | (w39491 & w39492);
assign w7748 = (~w3345 & w39493) | (~w3345 & w39494) | (w39493 & w39494);
assign w7749 = ~w7746 & ~w7747;
assign w7750 = ~w7748 & ~w7749;
assign w7751 = (~w7750 & w7738) | (~w7750 & w27148) | (w7738 & w27148);
assign w7752 = ~w7740 & ~w7751;
assign w7753 = ~w27148 & w29040;
assign w7754 = ~w7752 & ~w7753;
assign w7755 = (~w26562 & w27538) | (~w26562 & w27539) | (w27538 & w27539);
assign w7756 = w7754 & w7755;
assign w7757 = ~w7754 & ~w7755;
assign w7758 = ~w7756 & ~w7757;
assign w7759 = b_34 & w986;
assign w7760 = w1069 & w29041;
assign w7761 = b_33 & w981;
assign w7762 = ~w7760 & ~w7761;
assign w7763 = ~w7759 & w7762;
assign w7764 = (w7763 & ~w3967) | (w7763 & w29042) | (~w3967 & w29042);
assign w7765 = (w3967 & w39495) | (w3967 & w39496) | (w39495 & w39496);
assign w7766 = (~w3967 & w39497) | (~w3967 & w39498) | (w39497 & w39498);
assign w7767 = ~w7764 & ~w7765;
assign w7768 = ~w7766 & ~w7767;
assign w7769 = w7758 & ~w7768;
assign w7770 = w7758 & ~w7769;
assign w7771 = ~w7758 & ~w7768;
assign w7772 = ~w7770 & ~w7771;
assign w7773 = (~w7479 & w7291) | (~w7479 & w27149) | (w7291 & w27149);
assign w7774 = w7772 & w7773;
assign w7775 = ~w7772 & ~w7773;
assign w7776 = ~w7774 & ~w7775;
assign w7777 = b_37 & w657;
assign w7778 = w754 & w29043;
assign w7779 = b_36 & w652;
assign w7780 = ~w7778 & ~w7779;
assign w7781 = ~w7777 & w7780;
assign w7782 = (w7781 & ~w4636) | (w7781 & w26576) | (~w4636 & w26576);
assign w7783 = (w4636 & w29044) | (w4636 & w29045) | (w29044 & w29045);
assign w7784 = (~w4636 & w29046) | (~w4636 & w29047) | (w29046 & w29047);
assign w7785 = ~w7782 & ~w7783;
assign w7786 = ~w7784 & ~w7785;
assign w7787 = w7776 & ~w7786;
assign w7788 = w7776 & ~w7787;
assign w7789 = ~w7776 & ~w7786;
assign w7790 = ~w7788 & ~w7789;
assign w7791 = (~w25064 & w29048) | (~w25064 & w29049) | (w29048 & w29049);
assign w7792 = w7790 & w7791;
assign w7793 = ~w7790 & ~w7791;
assign w7794 = ~w7792 & ~w7793;
assign w7795 = b_40 & w418;
assign w7796 = w481 & w29050;
assign w7797 = b_39 & w413;
assign w7798 = ~w7796 & ~w7797;
assign w7799 = ~w7795 & w7798;
assign w7800 = (w7799 & ~w5363) | (w7799 & w25067) | (~w5363 & w25067);
assign w7801 = (w5363 & w26577) | (w5363 & w26578) | (w26577 & w26578);
assign w7802 = (~w5363 & w29051) | (~w5363 & w29052) | (w29051 & w29052);
assign w7803 = ~w7800 & ~w7801;
assign w7804 = ~w7802 & ~w7803;
assign w7805 = w7794 & ~w7804;
assign w7806 = w7794 & ~w7805;
assign w7807 = ~w7794 & ~w7804;
assign w7808 = ~w7806 & ~w7807;
assign w7809 = (~w7512 & w7516) | (~w7512 & w25068) | (w7516 & w25068);
assign w7810 = w7808 & w7809;
assign w7811 = ~w7808 & ~w7809;
assign w7812 = ~w7810 & ~w7811;
assign w7813 = b_43 & w239;
assign w7814 = w266 & w29053;
assign w7815 = b_42 & w234;
assign w7816 = ~w7814 & ~w7815;
assign w7817 = ~w7813 & w7816;
assign w7818 = (w7817 & ~w5888) | (w7817 & w25069) | (~w5888 & w25069);
assign w7819 = (w5888 & w29054) | (w5888 & w29055) | (w29054 & w29055);
assign w7820 = (~w5888 & w29056) | (~w5888 & w29057) | (w29056 & w29057);
assign w7821 = ~w7818 & ~w7819;
assign w7822 = ~w7820 & ~w7821;
assign w7823 = w7812 & ~w7822;
assign w7824 = w7812 & ~w7823;
assign w7825 = ~w7812 & ~w7822;
assign w7826 = ~w7824 & ~w7825;
assign w7827 = (~w7530 & w7533) | (~w7530 & w29058) | (w7533 & w29058);
assign w7828 = w7826 & w7827;
assign w7829 = (~w7246 & w27150) | (~w7246 & w27151) | (w27150 & w27151);
assign w7830 = ~w7828 & ~w7829;
assign w7831 = b_46 & w99;
assign w7832 = w136 & w29059;
assign w7833 = b_45 & w94;
assign w7834 = ~w7832 & ~w7833;
assign w7835 = ~w7831 & w7834;
assign w7836 = (w7835 & ~w6974) | (w7835 & w29060) | (~w6974 & w29060);
assign w7837 = (w6974 & w39499) | (w6974 & w39500) | (w39499 & w39500);
assign w7838 = (~w6974 & w39501) | (~w6974 & w39502) | (w39501 & w39502);
assign w7839 = ~w7836 & ~w7837;
assign w7840 = ~w7838 & ~w7839;
assign w7841 = ~w7829 & w29061;
assign w7842 = w7830 & ~w7841;
assign w7843 = (~w7840 & ~w29061) | (~w7840 & w39503) | (~w29061 & w39503);
assign w7844 = ~w7842 & ~w7843;
assign w7845 = ~w7547 & ~w7550;
assign w7846 = w7844 & w7845;
assign w7847 = ~w7844 & ~w7845;
assign w7848 = ~w7846 & ~w7847;
assign w7849 = w8 & w29062;
assign w7850 = ~w8 & w29063;
assign w7851 = b_48 & w4;
assign w7852 = ~w7850 & ~w7851;
assign w7853 = ~w7849 & w7852;
assign w7854 = ~b_48 & ~b_49;
assign w7855 = b_48 & b_49;
assign w7856 = ~w7854 & ~w7855;
assign w7857 = (w4656 & w39504) | (w4656 & w39505) | (w39504 & w39505);
assign w7858 = (~w4656 & w39506) | (~w4656 & w39507) | (w39506 & w39507);
assign w7859 = ~w7857 & ~w7858;
assign w7860 = (w7853 & ~w7859) | (w7853 & w29070) | (~w7859 & w29070);
assign w7861 = (w7859 & w39508) | (w7859 & w39509) | (w39508 & w39509);
assign w7862 = (~w7859 & w39510) | (~w7859 & w39511) | (w39510 & w39511);
assign w7863 = ~w7860 & ~w7861;
assign w7864 = ~w7862 & ~w7863;
assign w7865 = ~w7848 & w7864;
assign w7866 = w7848 & ~w7864;
assign w7867 = ~w7865 & ~w7866;
assign w7868 = ~w7557 & w7867;
assign w7869 = w7557 & ~w7867;
assign w7870 = ~w7868 & ~w7869;
assign w7871 = ~w7823 & ~w7829;
assign w7872 = b_35 & w986;
assign w7873 = w1069 & w29071;
assign w7874 = b_34 & w981;
assign w7875 = ~w7873 & ~w7874;
assign w7876 = ~w7872 & w7875;
assign w7877 = (w7876 & ~w4181) | (w7876 & w29072) | (~w4181 & w29072);
assign w7878 = (w4181 & w39512) | (w4181 & w39513) | (w39512 & w39513);
assign w7879 = (~w4181 & w39514) | (~w4181 & w39515) | (w39514 & w39515);
assign w7880 = ~w7877 & ~w7878;
assign w7881 = ~w7879 & ~w7880;
assign w7882 = (~w7751 & w7755) | (~w7751 & w27152) | (w7755 & w27152);
assign w7883 = b_32 & w1295;
assign w7884 = w1422 & w29073;
assign w7885 = b_31 & w1290;
assign w7886 = ~w7884 & ~w7885;
assign w7887 = ~w7883 & w7886;
assign w7888 = (w7887 & ~w3545) | (w7887 & w29074) | (~w3545 & w29074);
assign w7889 = (w3545 & w39516) | (w3545 & w39517) | (w39516 & w39517);
assign w7890 = (~w3545 & w39518) | (~w3545 & w39519) | (w39518 & w39519);
assign w7891 = ~w7888 & ~w7889;
assign w7892 = ~w7890 & ~w7891;
assign w7893 = (~w7734 & w7558) | (~w7734 & w27153) | (w7558 & w27153);
assign w7894 = b_29 & w1694;
assign w7895 = w1834 & w29075;
assign w7896 = b_28 & w1689;
assign w7897 = ~w7895 & ~w7896;
assign w7898 = ~w7894 & w7897;
assign w7899 = (w7898 & ~w2954) | (w7898 & w29076) | (~w2954 & w29076);
assign w7900 = (w2954 & w39520) | (w2954 & w39521) | (w39520 & w39521);
assign w7901 = (~w2954 & w39522) | (~w2954 & w39523) | (w39522 & w39523);
assign w7902 = ~w7899 & ~w7900;
assign w7903 = ~w7901 & ~w7902;
assign w7904 = (~w7726 & w7729) | (~w7726 & w27229) | (w7729 & w27229);
assign w7905 = (~w7708 & w7711) | (~w7708 & w39524) | (w7711 & w39524);
assign w7906 = ~w7672 & ~w7678;
assign w7907 = b_17 & w3803;
assign w7908 = w4027 & w29077;
assign w7909 = b_16 & w3798;
assign w7910 = ~w7908 & ~w7909;
assign w7911 = ~w7907 & w7910;
assign w7912 = (w7911 & ~w1038) | (w7911 & w29078) | (~w1038 & w29078);
assign w7913 = (w1038 & w39525) | (w1038 & w39526) | (w39525 & w39526);
assign w7914 = (~w1038 & w39527) | (~w1038 & w39528) | (w39527 & w39528);
assign w7915 = ~w7912 & ~w7913;
assign w7916 = ~w7914 & ~w7915;
assign w7917 = (~w7667 & ~w7668) | (~w7667 & w37616) | (~w7668 & w37616);
assign w7918 = b_14 & w4499;
assign w7919 = w4723 & w29079;
assign w7920 = b_13 & w4494;
assign w7921 = ~w7919 & ~w7920;
assign w7922 = ~w7918 & w7921;
assign w7923 = (w7922 & ~w735) | (w7922 & w29080) | (~w735 & w29080);
assign w7924 = (w735 & w39529) | (w735 & w39530) | (w39529 & w39530);
assign w7925 = (~w735 & w39531) | (~w735 & w39532) | (w39531 & w39532);
assign w7926 = ~w7923 & ~w7924;
assign w7927 = ~w7925 & ~w7926;
assign w7928 = (~w7631 & w7635) | (~w7631 & w29081) | (w7635 & w29081);
assign w7929 = b_8 & w5962;
assign w7930 = w6246 & w29082;
assign w7931 = b_7 & w5957;
assign w7932 = ~w7930 & ~w7931;
assign w7933 = ~w7929 & w7932;
assign w7934 = ~w308 & w29083;
assign w7935 = (w7933 & ~w29083) | (w7933 & w39533) | (~w29083 & w39533);
assign w7936 = (w29083 & w39534) | (w29083 & w39535) | (w39534 & w39535);
assign w7937 = ~w7934 & w29085;
assign w7938 = ~w7935 & ~w7936;
assign w7939 = ~w7937 & ~w7938;
assign w7940 = b_2 & w7613;
assign w7941 = w7348 & ~w7612;
assign w7942 = w7941 & w25372;
assign w7943 = b_1 & w7608;
assign w7944 = ~w7942 & ~w7943;
assign w7945 = ~w7940 & w7944;
assign w7946 = w35 & w7616;
assign w7947 = w7945 & ~w7946;
assign w7948 = (a_50 & ~w7945) | (a_50 & w25373) | (~w7945 & w25373);
assign w7949 = w7945 & w25555;
assign w7950 = ~w7947 & ~w7948;
assign w7951 = ~w7949 & ~w7950;
assign w7952 = ~w7622 & w7951;
assign w7953 = w7622 & ~w7951;
assign w7954 = ~w7952 & ~w7953;
assign w7955 = b_5 & w6761;
assign w7956 = w7075 & w26158;
assign w7957 = b_4 & w6756;
assign w7958 = ~w7956 & ~w7957;
assign w7959 = ~w7955 & w7958;
assign w7960 = w129 & w6764;
assign w7961 = w7959 & ~w7960;
assign w7962 = (a_47 & w7960) | (a_47 & w26159) | (w7960 & w26159);
assign w7963 = ~w7960 & w39536;
assign w7964 = ~w7961 & ~w7962;
assign w7965 = ~w7963 & ~w7964;
assign w7966 = w7954 & ~w7965;
assign w7967 = w7954 & ~w7966;
assign w7968 = ~w7954 & ~w7965;
assign w7969 = ~w7967 & ~w7968;
assign w7970 = (~w7969 & w7628) | (~w7969 & w25374) | (w7628 & w25374);
assign w7971 = ~w7628 & w25375;
assign w7972 = ~w7970 & ~w7971;
assign w7973 = ~w7939 & w7972;
assign w7974 = ~w7972 & ~w7939;
assign w7975 = w7972 & ~w7973;
assign w7976 = ~w7974 & ~w7975;
assign w7977 = ~w7928 & ~w7976;
assign w7978 = ~w7928 & ~w7977;
assign w7979 = b_11 & w5196;
assign w7980 = w5459 & w29086;
assign w7981 = b_10 & w5191;
assign w7982 = ~w7980 & ~w7981;
assign w7983 = ~w7979 & w7982;
assign w7984 = (w7983 & ~w530) | (w7983 & w29087) | (~w530 & w29087);
assign w7985 = (w530 & w39537) | (w530 & w39538) | (w39537 & w39538);
assign w7986 = (~w530 & w39539) | (~w530 & w39540) | (w39539 & w39540);
assign w7987 = ~w7984 & ~w7985;
assign w7988 = ~w7986 & ~w7987;
assign w7989 = ~w7978 & w27036;
assign w7990 = (~w7988 & w7978) | (~w7988 & w27037) | (w7978 & w27037);
assign w7991 = ~w7989 & ~w7990;
assign w7992 = (w7991 & w7651) | (w7991 & w25376) | (w7651 & w25376);
assign w7993 = w7653 & ~w7991;
assign w7994 = ~w7992 & ~w7993;
assign w7995 = ~w7992 & w26793;
assign w7996 = w7994 & ~w7995;
assign w7997 = (~w7927 & w7992) | (~w7927 & w27345) | (w7992 & w27345);
assign w7998 = ~w7996 & ~w7997;
assign w7999 = ~w7917 & ~w7998;
assign w8000 = w7917 & w7998;
assign w8001 = ~w7999 & ~w8000;
assign w8002 = ~w7916 & w8001;
assign w8003 = ~w8001 & ~w7916;
assign w8004 = w8001 & ~w8002;
assign w8005 = ~w8003 & ~w8004;
assign w8006 = ~w7906 & ~w8005;
assign w8007 = ~w7906 & ~w8006;
assign w8008 = w7906 & ~w8005;
assign w8009 = ~w8007 & ~w8008;
assign w8010 = b_20 & w3195;
assign w8011 = w3388 & w29088;
assign w8012 = b_19 & w3190;
assign w8013 = ~w8011 & ~w8012;
assign w8014 = ~w8010 & w8013;
assign w8015 = (w8014 & ~w1503) | (w8014 & w29089) | (~w1503 & w29089);
assign w8016 = (w1503 & w39541) | (w1503 & w39542) | (w39541 & w39542);
assign w8017 = (~w1503 & w39543) | (~w1503 & w39544) | (w39543 & w39544);
assign w8018 = ~w8015 & ~w8016;
assign w8019 = ~w8017 & ~w8018;
assign w8020 = (~w8019 & w8007) | (~w8019 & w37617) | (w8007 & w37617);
assign w8021 = ~w8009 & ~w8020;
assign w8022 = ~w8007 & w39545;
assign w8023 = ~w8021 & ~w8022;
assign w8024 = (~w7690 & w7694) | (~w7690 & w27154) | (w7694 & w27154);
assign w8025 = ~w8021 & w27739;
assign w8026 = (~w8024 & w8021) | (~w8024 & w27740) | (w8021 & w27740);
assign w8027 = ~w8025 & ~w8026;
assign w8028 = b_23 & w2639;
assign w8029 = w2820 & w29090;
assign w8030 = b_22 & w2634;
assign w8031 = ~w8029 & ~w8030;
assign w8032 = ~w8028 & w8031;
assign w8033 = (w8032 & ~w1933) | (w8032 & w29091) | (~w1933 & w29091);
assign w8034 = (w1933 & w39546) | (w1933 & w39547) | (w39546 & w39547);
assign w8035 = (~w1933 & w39548) | (~w1933 & w39549) | (w39548 & w39549);
assign w8036 = ~w8033 & ~w8034;
assign w8037 = ~w8035 & ~w8036;
assign w8038 = w8027 & ~w8037;
assign w8039 = ~w8027 & w8037;
assign w8040 = (w7714 & w27155) | (w7714 & w27156) | (w27155 & w27156);
assign w8041 = ~w7905 & ~w8040;
assign w8042 = ~w8038 & ~w8040;
assign w8043 = ~w8040 & w27156;
assign w8044 = ~w8041 & ~w8043;
assign w8045 = b_26 & w2158;
assign w8046 = w2294 & w29092;
assign w8047 = b_25 & w2153;
assign w8048 = ~w8046 & ~w8047;
assign w8049 = ~w8045 & w8048;
assign w8050 = (w8049 & ~w2416) | (w8049 & w29093) | (~w2416 & w29093);
assign w8051 = (w2416 & w39550) | (w2416 & w39551) | (w39550 & w39551);
assign w8052 = (~w2416 & w39552) | (~w2416 & w39553) | (w39552 & w39553);
assign w8053 = ~w8050 & ~w8051;
assign w8054 = ~w8052 & ~w8053;
assign w8055 = w8044 & w8054;
assign w8056 = ~w8044 & ~w8054;
assign w8057 = ~w8055 & ~w8056;
assign w8058 = ~w7904 & w8057;
assign w8059 = w7904 & ~w8057;
assign w8060 = ~w8058 & ~w8059;
assign w8061 = w7903 & ~w8060;
assign w8062 = ~w7903 & w8060;
assign w8063 = ~w8061 & ~w8062;
assign w8064 = ~w7893 & w8063;
assign w8065 = w7893 & ~w8063;
assign w8066 = ~w8064 & ~w8065;
assign w8067 = w7892 & ~w8066;
assign w8068 = ~w7892 & w8066;
assign w8069 = ~w8067 & ~w8068;
assign w8070 = (w8069 & w7757) | (w8069 & w25378) | (w7757 & w25378);
assign w8071 = ~w7757 & w25379;
assign w8072 = ~w8070 & ~w8071;
assign w8073 = ~w7881 & w8072;
assign w8074 = w8072 & ~w8073;
assign w8075 = ~w8072 & ~w7881;
assign w8076 = ~w8074 & ~w8075;
assign w8077 = (~w7769 & w7773) | (~w7769 & w26581) | (w7773 & w26581);
assign w8078 = w8076 & w8077;
assign w8079 = ~w8076 & ~w8077;
assign w8080 = ~w8078 & ~w8079;
assign w8081 = b_38 & w657;
assign w8082 = w754 & w29094;
assign w8083 = b_37 & w652;
assign w8084 = ~w8082 & ~w8083;
assign w8085 = ~w8081 & w8084;
assign w8086 = (w8085 & ~w4658) | (w8085 & w25380) | (~w4658 & w25380);
assign w8087 = (w4658 & w29095) | (w4658 & w29096) | (w29095 & w29096);
assign w8088 = (~w4658 & w29097) | (~w4658 & w29098) | (w29097 & w29098);
assign w8089 = ~w8086 & ~w8087;
assign w8090 = ~w8088 & ~w8089;
assign w8091 = w8080 & ~w8090;
assign w8092 = w8080 & ~w8091;
assign w8093 = ~w8080 & ~w8090;
assign w8094 = ~w8092 & ~w8093;
assign w8095 = (~w7787 & w7791) | (~w7787 & w27157) | (w7791 & w27157);
assign w8096 = w8094 & w8095;
assign w8097 = ~w8094 & ~w8095;
assign w8098 = ~w8096 & ~w8097;
assign w8099 = b_41 & w418;
assign w8100 = w481 & w29099;
assign w8101 = b_40 & w413;
assign w8102 = ~w8100 & ~w8101;
assign w8103 = ~w8099 & w8102;
assign w8104 = (w8103 & ~w5609) | (w8103 & w25070) | (~w5609 & w25070);
assign w8105 = (w5609 & w25381) | (w5609 & w25382) | (w25381 & w25382);
assign w8106 = (~w5609 & w29100) | (~w5609 & w29101) | (w29100 & w29101);
assign w8107 = ~w8104 & ~w8105;
assign w8108 = ~w8106 & ~w8107;
assign w8109 = w8098 & ~w8108;
assign w8110 = w8098 & ~w8109;
assign w8111 = ~w8098 & ~w8108;
assign w8112 = ~w8110 & ~w8111;
assign w8113 = (~w7805 & w7808) | (~w7805 & w27741) | (w7808 & w27741);
assign w8114 = w8112 & w8113;
assign w8115 = ~w8112 & ~w8113;
assign w8116 = ~w8114 & ~w8115;
assign w8117 = b_44 & w239;
assign w8118 = w266 & w29102;
assign w8119 = b_43 & w234;
assign w8120 = ~w8118 & ~w8119;
assign w8121 = ~w8117 & w8120;
assign w8122 = (w8121 & ~w6408) | (w8121 & w25383) | (~w6408 & w25383);
assign w8123 = (w6408 & w29103) | (w6408 & w29104) | (w29103 & w29104);
assign w8124 = (~w6408 & w29105) | (~w6408 & w29106) | (w29105 & w29106);
assign w8125 = ~w8122 & ~w8123;
assign w8126 = ~w8124 & ~w8125;
assign w8127 = w8116 & ~w8126;
assign w8128 = ~w8116 & w8126;
assign w8129 = (w25071 & w7829) | (w25071 & w27742) | (w7829 & w27742);
assign w8130 = ~w7871 & ~w8129;
assign w8131 = (~w7829 & w27743) | (~w7829 & w27744) | (w27743 & w27744);
assign w8132 = ~w8128 & w8131;
assign w8133 = ~w8130 & ~w8132;
assign w8134 = b_47 & w99;
assign w8135 = w136 & w29107;
assign w8136 = b_46 & w94;
assign w8137 = ~w8135 & ~w8136;
assign w8138 = ~w8134 & w8137;
assign w8139 = (w8138 & ~w6998) | (w8138 & w25384) | (~w6998 & w25384);
assign w8140 = (w6998 & w29108) | (w6998 & w29109) | (w29108 & w29109);
assign w8141 = (~w6998 & w29110) | (~w6998 & w29111) | (w29110 & w29111);
assign w8142 = ~w8139 & ~w8140;
assign w8143 = ~w8141 & ~w8142;
assign w8144 = ~w8133 & ~w8143;
assign w8145 = ~w8133 & ~w8144;
assign w8146 = w8133 & ~w8143;
assign w8147 = ~w8145 & ~w8146;
assign w8148 = (~w7841 & w7845) | (~w7841 & w25072) | (w7845 & w25072);
assign w8149 = w8147 & w8148;
assign w8150 = ~w8147 & ~w8148;
assign w8151 = ~w8149 & ~w8150;
assign w8152 = w8 & w29112;
assign w8153 = ~w8 & w29113;
assign w8154 = b_49 & w4;
assign w8155 = ~w8153 & ~w8154;
assign w8156 = ~w8152 & w8155;
assign w8157 = ~b_49 & ~b_50;
assign w8158 = b_49 & b_50;
assign w8159 = ~w8157 & ~w8158;
assign w8160 = (w4656 & w39554) | (w4656 & w39555) | (w39554 & w39555);
assign w8161 = (~w4656 & w39556) | (~w4656 & w39557) | (w39556 & w39557);
assign w8162 = ~w8160 & ~w8161;
assign w8163 = (w8156 & ~w8162) | (w8156 & w29119) | (~w8162 & w29119);
assign w8164 = (w8162 & w39558) | (w8162 & w39559) | (w39558 & w39559);
assign w8165 = (~w8162 & w39560) | (~w8162 & w39561) | (w39560 & w39561);
assign w8166 = ~w8163 & ~w8164;
assign w8167 = ~w8165 & ~w8166;
assign w8168 = w8151 & ~w8167;
assign w8169 = w8151 & ~w8168;
assign w8170 = ~w8151 & ~w8167;
assign w8171 = ~w8169 & ~w8170;
assign w8172 = (~w7270 & w27158) | (~w7270 & w27159) | (w27158 & w27159);
assign w8173 = ~w8171 & ~w8172;
assign w8174 = w8171 & w8172;
assign w8175 = ~w8173 & ~w8174;
assign w8176 = w8 & w29120;
assign w8177 = ~w8 & w29121;
assign w8178 = b_50 & w4;
assign w8179 = ~w8177 & ~w8178;
assign w8180 = ~w8176 & w8179;
assign w8181 = ~b_50 & ~b_51;
assign w8182 = b_50 & b_51;
assign w8183 = ~w8181 & ~w8182;
assign w8184 = (w4656 & w39562) | (w4656 & w39563) | (w39562 & w39563);
assign w8185 = (~w4656 & w39564) | (~w4656 & w39565) | (w39564 & w39565);
assign w8186 = ~w8184 & ~w8185;
assign w8187 = (w8180 & ~w8186) | (w8180 & w29127) | (~w8186 & w29127);
assign w8188 = (w8186 & w39566) | (w8186 & w39567) | (w39566 & w39567);
assign w8189 = (~w8186 & w39568) | (~w8186 & w39569) | (w39568 & w39569);
assign w8190 = ~w8187 & ~w8188;
assign w8191 = ~w8189 & ~w8190;
assign w8192 = (~w8144 & w8147) | (~w8144 & w29128) | (w8147 & w29128);
assign w8193 = b_45 & w239;
assign w8194 = w266 & w29129;
assign w8195 = b_44 & w234;
assign w8196 = ~w8194 & ~w8195;
assign w8197 = ~w8193 & w8196;
assign w8198 = (w8197 & ~w6682) | (w8197 & w25389) | (~w6682 & w25389);
assign w8199 = (w6682 & w26584) | (w6682 & w26585) | (w26584 & w26585);
assign w8200 = (~w6682 & w29130) | (~w6682 & w29131) | (w29130 & w29131);
assign w8201 = ~w8198 & ~w8199;
assign w8202 = ~w8200 & ~w8201;
assign w8203 = (~w8068 & w7882) | (~w8068 & w25073) | (w7882 & w25073);
assign w8204 = b_33 & w1295;
assign w8205 = w1422 & w29132;
assign w8206 = b_32 & w1290;
assign w8207 = ~w8205 & ~w8206;
assign w8208 = ~w8204 & w8207;
assign w8209 = (w8208 & ~w3744) | (w8208 & w25390) | (~w3744 & w25390);
assign w8210 = (w3744 & w26586) | (w3744 & w26587) | (w26586 & w26587);
assign w8211 = (~w3744 & w29133) | (~w3744 & w29134) | (w29133 & w29134);
assign w8212 = ~w8209 & ~w8210;
assign w8213 = ~w8211 & ~w8212;
assign w8214 = (~w8062 & w7893) | (~w8062 & w25391) | (w7893 & w25391);
assign w8215 = (~w8056 & ~w8057) | (~w8056 & w25074) | (~w8057 & w25074);
assign w8216 = b_27 & w2158;
assign w8217 = w2294 & w29135;
assign w8218 = b_26 & w2153;
assign w8219 = ~w8217 & ~w8218;
assign w8220 = ~w8216 & w8219;
assign w8221 = (w8220 & ~w2582) | (w8220 & w29136) | (~w2582 & w29136);
assign w8222 = (w2582 & w39570) | (w2582 & w39571) | (w39570 & w39571);
assign w8223 = (~w2582 & w39572) | (~w2582 & w39573) | (w39572 & w39573);
assign w8224 = ~w8221 & ~w8222;
assign w8225 = ~w8223 & ~w8224;
assign w8226 = (~w8002 & w7906) | (~w8002 & w25392) | (w7906 & w25392);
assign w8227 = b_18 & w3803;
assign w8228 = w4027 & w29137;
assign w8229 = b_17 & w3798;
assign w8230 = ~w8228 & ~w8229;
assign w8231 = ~w8227 & w8230;
assign w8232 = (w8231 & ~w1238) | (w8231 & w29138) | (~w1238 & w29138);
assign w8233 = (w1238 & w39574) | (w1238 & w39575) | (w39574 & w39575);
assign w8234 = (~w1238 & w39576) | (~w1238 & w39577) | (w39576 & w39577);
assign w8235 = ~w8232 & ~w8233;
assign w8236 = ~w8234 & ~w8235;
assign w8237 = (~w7995 & w7998) | (~w7995 & w26910) | (w7998 & w26910);
assign w8238 = b_15 & w4499;
assign w8239 = w4723 & w29139;
assign w8240 = b_14 & w4494;
assign w8241 = ~w8239 & ~w8240;
assign w8242 = ~w8238 & w8241;
assign w8243 = (w8242 & ~w827) | (w8242 & w29140) | (~w827 & w29140);
assign w8244 = (w827 & w39578) | (w827 & w39579) | (w39578 & w39579);
assign w8245 = (~w827 & w39580) | (~w827 & w39581) | (w39580 & w39581);
assign w8246 = ~w8243 & ~w8244;
assign w8247 = ~w8245 & ~w8246;
assign w8248 = (~w25376 & w26588) | (~w25376 & w26589) | (w26588 & w26589);
assign w8249 = b_12 & w5196;
assign w8250 = w5459 & w29141;
assign w8251 = b_11 & w5191;
assign w8252 = ~w8250 & ~w8251;
assign w8253 = ~w8249 & w8252;
assign w8254 = (w8253 & ~w552) | (w8253 & w29142) | (~w552 & w29142);
assign w8255 = (w552 & w39582) | (w552 & w39583) | (w39582 & w39583);
assign w8256 = (~w552 & w39584) | (~w552 & w39585) | (w39584 & w39585);
assign w8257 = ~w8254 & ~w8255;
assign w8258 = ~w8256 & ~w8257;
assign w8259 = b_6 & w6761;
assign w8260 = w7075 & w29143;
assign w8261 = b_5 & w6756;
assign w8262 = ~w8260 & ~w8261;
assign w8263 = ~w8259 & w8262;
assign w8264 = (w8263 & ~w190) | (w8263 & w29144) | (~w190 & w29144);
assign w8265 = (w190 & w39586) | (w190 & w39587) | (w39586 & w39587);
assign w8266 = (~w190 & w39588) | (~w190 & w39589) | (w39588 & w39589);
assign w8267 = ~w8264 & ~w8265;
assign w8268 = ~w8266 & ~w8267;
assign w8269 = a_50 & ~a_51;
assign w8270 = ~a_50 & a_51;
assign w8271 = ~w8269 & ~w8270;
assign w8272 = b_0 & ~w8271;
assign w8273 = (w8272 & ~w7622) | (w8272 & w25394) | (~w7622 & w25394);
assign w8274 = w7622 & w25395;
assign w8275 = ~w8273 & ~w8274;
assign w8276 = b_3 & w7613;
assign w8277 = w7941 & w25811;
assign w8278 = b_2 & w7608;
assign w8279 = ~w8277 & ~w8278;
assign w8280 = ~w8276 & w8279;
assign w8281 = w57 & w7616;
assign w8282 = w8280 & ~w8281;
assign w8283 = a_50 & ~w8282;
assign w8284 = w8282 & a_50;
assign w8285 = ~w8282 & ~w8283;
assign w8286 = ~w8284 & ~w8285;
assign w8287 = ~w8275 & ~w8286;
assign w8288 = w8275 & w8286;
assign w8289 = ~w8287 & ~w8288;
assign w8290 = ~w8268 & w8289;
assign w8291 = w8289 & ~w8290;
assign w8292 = ~w8289 & ~w8268;
assign w8293 = ~w8291 & ~w8292;
assign w8294 = (~w25374 & w26160) | (~w25374 & w26161) | (w26160 & w26161);
assign w8295 = w8293 & w8294;
assign w8296 = ~w8293 & ~w8294;
assign w8297 = ~w8295 & ~w8296;
assign w8298 = b_9 & w5962;
assign w8299 = w6246 & w29145;
assign w8300 = b_8 & w5957;
assign w8301 = ~w8299 & ~w8300;
assign w8302 = ~w8298 & w8301;
assign w8303 = (w8302 & ~w371) | (w8302 & w29146) | (~w371 & w29146);
assign w8304 = (w371 & w39590) | (w371 & w39591) | (w39590 & w39591);
assign w8305 = (~w371 & w39592) | (~w371 & w39593) | (w39592 & w39593);
assign w8306 = ~w8303 & ~w8304;
assign w8307 = ~w8305 & ~w8306;
assign w8308 = ~w8297 & w8307;
assign w8309 = w8297 & ~w8307;
assign w8310 = ~w8308 & ~w8309;
assign w8311 = (~w25393 & w26162) | (~w25393 & w26163) | (w26162 & w26163);
assign w8312 = (w25393 & w26794) | (w25393 & w26795) | (w26794 & w26795);
assign w8313 = ~w8311 & ~w8312;
assign w8314 = ~w8258 & w8313;
assign w8315 = ~w8313 & ~w8258;
assign w8316 = w8313 & ~w8314;
assign w8317 = ~w8315 & ~w8316;
assign w8318 = ~w8248 & ~w8317;
assign w8319 = w8248 & w8317;
assign w8320 = ~w8318 & ~w8319;
assign w8321 = ~w8247 & w8320;
assign w8322 = w8247 & ~w8320;
assign w8323 = ~w8321 & ~w8322;
assign w8324 = ~w8237 & w8323;
assign w8325 = w8237 & ~w8323;
assign w8326 = ~w8324 & ~w8325;
assign w8327 = ~w8236 & w8326;
assign w8328 = w8236 & ~w8326;
assign w8329 = ~w8327 & ~w8328;
assign w8330 = (~w25392 & w26911) | (~w25392 & w26912) | (w26911 & w26912);
assign w8331 = w8226 & ~w8329;
assign w8332 = ~w8330 & ~w8331;
assign w8333 = b_21 & w3195;
assign w8334 = w3388 & w29147;
assign w8335 = b_20 & w3190;
assign w8336 = ~w8334 & ~w8335;
assign w8337 = ~w8333 & w8336;
assign w8338 = (w8337 & ~w1634) | (w8337 & w29148) | (~w1634 & w29148);
assign w8339 = (w1634 & w39594) | (w1634 & w39595) | (w39594 & w39595);
assign w8340 = (~w1634 & w39596) | (~w1634 & w39597) | (w39596 & w39597);
assign w8341 = ~w8338 & ~w8339;
assign w8342 = ~w8340 & ~w8341;
assign w8343 = w8332 & ~w8342;
assign w8344 = w8332 & ~w8343;
assign w8345 = ~w8332 & ~w8342;
assign w8346 = ~w8344 & ~w8345;
assign w8347 = (~w8020 & w8023) | (~w8020 & w27160) | (w8023 & w27160);
assign w8348 = w8346 & w8347;
assign w8349 = ~w8346 & ~w8347;
assign w8350 = ~w8348 & ~w8349;
assign w8351 = b_24 & w2639;
assign w8352 = w2820 & w29149;
assign w8353 = b_23 & w2634;
assign w8354 = ~w8352 & ~w8353;
assign w8355 = ~w8351 & w8354;
assign w8356 = (w8355 & ~w2083) | (w8355 & w29150) | (~w2083 & w29150);
assign w8357 = (w2083 & w39598) | (w2083 & w39599) | (w39598 & w39599);
assign w8358 = (~w2083 & w39600) | (~w2083 & w39601) | (w39600 & w39601);
assign w8359 = ~w8356 & ~w8357;
assign w8360 = ~w8358 & ~w8359;
assign w8361 = ~w8350 & w8360;
assign w8362 = w8350 & ~w8360;
assign w8363 = ~w8361 & ~w8362;
assign w8364 = ~w8042 & w8363;
assign w8365 = w8042 & ~w8363;
assign w8366 = ~w8364 & ~w8365;
assign w8367 = ~w8225 & w8366;
assign w8368 = w8366 & ~w8367;
assign w8369 = ~w8366 & ~w8225;
assign w8370 = ~w8368 & ~w8369;
assign w8371 = ~w8215 & w8370;
assign w8372 = w8215 & ~w8370;
assign w8373 = ~w8371 & ~w8372;
assign w8374 = b_30 & w1694;
assign w8375 = w1834 & w29151;
assign w8376 = b_29 & w1689;
assign w8377 = ~w8375 & ~w8376;
assign w8378 = ~w8374 & w8377;
assign w8379 = (w8378 & ~w3138) | (w8378 & w29152) | (~w3138 & w29152);
assign w8380 = (w3138 & w39602) | (w3138 & w39603) | (w39602 & w39603);
assign w8381 = (~w3138 & w39604) | (~w3138 & w39605) | (w39604 & w39605);
assign w8382 = ~w8379 & ~w8380;
assign w8383 = ~w8381 & ~w8382;
assign w8384 = ~w8373 & ~w8383;
assign w8385 = w8373 & w8383;
assign w8386 = ~w8384 & ~w8385;
assign w8387 = ~w8214 & w8386;
assign w8388 = w8214 & ~w8386;
assign w8389 = ~w8387 & ~w8388;
assign w8390 = ~w8213 & w8389;
assign w8391 = w8389 & ~w8390;
assign w8392 = ~w8389 & ~w8213;
assign w8393 = ~w8391 & ~w8392;
assign w8394 = ~w8203 & w8393;
assign w8395 = w8203 & ~w8393;
assign w8396 = ~w8394 & ~w8395;
assign w8397 = b_36 & w986;
assign w8398 = w1069 & w29153;
assign w8399 = b_35 & w981;
assign w8400 = ~w8398 & ~w8399;
assign w8401 = ~w8397 & w8400;
assign w8402 = (w8401 & ~w4395) | (w8401 & w25396) | (~w4395 & w25396);
assign w8403 = (w4395 & w29154) | (w4395 & w29155) | (w29154 & w29155);
assign w8404 = (~w4395 & w29156) | (~w4395 & w29157) | (w29156 & w29157);
assign w8405 = ~w8402 & ~w8403;
assign w8406 = ~w8404 & ~w8405;
assign w8407 = ~w8396 & ~w8406;
assign w8408 = w8396 & w8406;
assign w8409 = ~w8407 & ~w8408;
assign w8410 = ~w8079 & w25075;
assign w8411 = (w8409 & w8079) | (w8409 & w25076) | (w8079 & w25076);
assign w8412 = ~w8410 & ~w8411;
assign w8413 = b_39 & w657;
assign w8414 = w754 & w29158;
assign w8415 = b_38 & w652;
assign w8416 = ~w8414 & ~w8415;
assign w8417 = ~w8413 & w8416;
assign w8418 = (w8417 & ~w4888) | (w8417 & w25077) | (~w4888 & w25077);
assign w8419 = (w4888 & w25397) | (w4888 & w25398) | (w25397 & w25398);
assign w8420 = (~w4888 & w29159) | (~w4888 & w29160) | (w29159 & w29160);
assign w8421 = ~w8418 & ~w8419;
assign w8422 = ~w8420 & ~w8421;
assign w8423 = w8412 & ~w8422;
assign w8424 = w8412 & ~w8423;
assign w8425 = ~w8412 & ~w8422;
assign w8426 = ~w8424 & ~w8425;
assign w8427 = (~w8091 & w8095) | (~w8091 & w26590) | (w8095 & w26590);
assign w8428 = w8426 & w8427;
assign w8429 = ~w8426 & ~w8427;
assign w8430 = ~w8428 & ~w8429;
assign w8431 = b_42 & w418;
assign w8432 = w481 & w29161;
assign w8433 = b_41 & w413;
assign w8434 = ~w8432 & ~w8433;
assign w8435 = ~w8431 & w8434;
assign w8436 = (w8435 & ~w5864) | (w8435 & w25078) | (~w5864 & w25078);
assign w8437 = (w5864 & w25399) | (w5864 & w25400) | (w25399 & w25400);
assign w8438 = (~w5864 & w29162) | (~w5864 & w29163) | (w29162 & w29163);
assign w8439 = ~w8436 & ~w8437;
assign w8440 = ~w8438 & ~w8439;
assign w8441 = ~w8430 & w8440;
assign w8442 = w8430 & ~w8440;
assign w8443 = ~w8441 & ~w8442;
assign w8444 = (~w8109 & w8113) | (~w8109 & w27161) | (w8113 & w27161);
assign w8445 = w8443 & ~w8444;
assign w8446 = ~w8443 & w8444;
assign w8447 = ~w8445 & ~w8446;
assign w8448 = ~w8202 & w8447;
assign w8449 = w8447 & ~w8448;
assign w8450 = ~w8447 & ~w8202;
assign w8451 = ~w8449 & ~w8450;
assign w8452 = ~w8131 & w8451;
assign w8453 = w8131 & ~w8451;
assign w8454 = ~w8452 & ~w8453;
assign w8455 = b_48 & w99;
assign w8456 = w136 & w29164;
assign w8457 = b_47 & w94;
assign w8458 = ~w8456 & ~w8457;
assign w8459 = ~w8455 & w8458;
assign w8460 = (w8459 & ~w7284) | (w8459 & w29165) | (~w7284 & w29165);
assign w8461 = (w7284 & w39606) | (w7284 & w39607) | (w39606 & w39607);
assign w8462 = (~w7284 & w39608) | (~w7284 & w39609) | (w39608 & w39609);
assign w8463 = ~w8460 & ~w8461;
assign w8464 = ~w8462 & ~w8463;
assign w8465 = w8454 & w8464;
assign w8466 = ~w8454 & ~w8464;
assign w8467 = ~w8465 & ~w8466;
assign w8468 = ~w8192 & w8467;
assign w8469 = w8192 & ~w8467;
assign w8470 = ~w8468 & ~w8469;
assign w8471 = ~w8191 & w8470;
assign w8472 = w8191 & ~w8470;
assign w8473 = ~w8471 & ~w8472;
assign w8474 = (w8473 & w8173) | (w8473 & w29166) | (w8173 & w29166);
assign w8475 = ~w8173 & w29167;
assign w8476 = ~w8474 & ~w8475;
assign w8477 = (~w8466 & w8192) | (~w8466 & w29168) | (w8192 & w29168);
assign w8478 = (~w8442 & w8444) | (~w8442 & w25079) | (w8444 & w25079);
assign w8479 = (~w8367 & w8215) | (~w8367 & w27162) | (w8215 & w27162);
assign w8480 = (~w8362 & w8042) | (~w8362 & w27346) | (w8042 & w27346);
assign w8481 = ~w8327 & ~w8330;
assign w8482 = b_16 & w4499;
assign w8483 = w4723 & w29169;
assign w8484 = b_15 & w4494;
assign w8485 = ~w8483 & ~w8484;
assign w8486 = ~w8482 & w8485;
assign w8487 = (w8486 & ~w926) | (w8486 & w29170) | (~w926 & w29170);
assign w8488 = (w926 & w39610) | (w926 & w39611) | (w39610 & w39611);
assign w8489 = (~w926 & w39612) | (~w926 & w39613) | (w39612 & w39613);
assign w8490 = ~w8487 & ~w8488;
assign w8491 = ~w8489 & ~w8490;
assign w8492 = (~w8314 & w8248) | (~w8314 & w26796) | (w8248 & w26796);
assign w8493 = ~w8309 & ~w8311;
assign w8494 = b_7 & w6761;
assign w8495 = w7075 & w29171;
assign w8496 = b_6 & w6756;
assign w8497 = ~w8495 & ~w8496;
assign w8498 = ~w8494 & w8497;
assign w8499 = (w8498 & ~w213) | (w8498 & w29172) | (~w213 & w29172);
assign w8500 = (w213 & w39614) | (w213 & w39615) | (w39614 & w39615);
assign w8501 = (~w213 & w39616) | (~w213 & w39617) | (w39616 & w39617);
assign w8502 = ~w8499 & ~w8500;
assign w8503 = ~w8501 & ~w8502;
assign w8504 = ~w7951 & w25812;
assign w8505 = (~w8504 & w8275) | (~w8504 & w25556) | (w8275 & w25556);
assign w8506 = b_4 & w7613;
assign w8507 = w7941 & w25813;
assign w8508 = b_3 & w7608;
assign w8509 = ~w8507 & ~w8508;
assign w8510 = ~w8506 & w8509;
assign w8511 = w84 & w7616;
assign w8512 = w8510 & ~w8511;
assign w8513 = (a_50 & w8511) | (a_50 & w25814) | (w8511 & w25814);
assign w8514 = ~w8511 & w26164;
assign w8515 = ~w8512 & ~w8513;
assign w8516 = ~w8514 & ~w8515;
assign w8517 = (a_53 & w8271) | (a_53 & w29173) | (w8271 & w29173);
assign w8518 = ~a_51 & a_52;
assign w8519 = a_51 & ~a_52;
assign w8520 = ~w8518 & ~w8519;
assign w8521 = w8271 & ~w8520;
assign w8522 = b_0 & w8521;
assign w8523 = ~a_52 & a_53;
assign w8524 = a_52 & ~a_53;
assign w8525 = ~w8523 & ~w8524;
assign w8526 = ~w8271 & w8525;
assign w8527 = b_1 & w8526;
assign w8528 = ~w8522 & ~w8527;
assign w8529 = ~w8271 & ~w8525;
assign w8530 = ~w15 & w8529;
assign w8531 = w8528 & ~w8530;
assign w8532 = (a_53 & ~w8528) | (a_53 & w25557) | (~w8528 & w25557);
assign w8533 = w8528 & w25815;
assign w8534 = ~w8531 & ~w8532;
assign w8535 = (w8517 & w8534) | (w8517 & w25816) | (w8534 & w25816);
assign w8536 = ~w8534 & w26165;
assign w8537 = ~w8535 & ~w8536;
assign w8538 = w8516 & ~w8537;
assign w8539 = ~w8516 & w8537;
assign w8540 = ~w8538 & ~w8539;
assign w8541 = ~w8505 & w8540;
assign w8542 = w8505 & ~w8540;
assign w8543 = ~w8541 & ~w8542;
assign w8544 = ~w8503 & w8543;
assign w8545 = w8543 & ~w8544;
assign w8546 = ~w8543 & ~w8503;
assign w8547 = ~w8545 & ~w8546;
assign w8548 = (~w8290 & w8293) | (~w8290 & w27038) | (w8293 & w27038);
assign w8549 = w8547 & w8548;
assign w8550 = ~w8547 & ~w8548;
assign w8551 = ~w8549 & ~w8550;
assign w8552 = b_10 & w5962;
assign w8553 = w6246 & w29174;
assign w8554 = b_9 & w5957;
assign w8555 = ~w8553 & ~w8554;
assign w8556 = ~w8552 & w8555;
assign w8557 = (w8556 & ~w454) | (w8556 & w29175) | (~w454 & w29175);
assign w8558 = (w454 & w39618) | (w454 & w39619) | (w39618 & w39619);
assign w8559 = (~w454 & w39620) | (~w454 & w39621) | (w39620 & w39621);
assign w8560 = ~w8557 & ~w8558;
assign w8561 = ~w8559 & ~w8560;
assign w8562 = w8551 & ~w8561;
assign w8563 = ~w8551 & w8561;
assign w8564 = (w8311 & w26797) | (w8311 & w27039) | (w26797 & w27039);
assign w8565 = ~w8493 & ~w8564;
assign w8566 = (~w8311 & w27040) | (~w8311 & w27041) | (w27040 & w27041);
assign w8567 = (~w8311 & w27230) | (~w8311 & w27231) | (w27230 & w27231);
assign w8568 = b_13 & w5196;
assign w8569 = w5459 & w29176;
assign w8570 = b_12 & w5191;
assign w8571 = ~w8569 & ~w8570;
assign w8572 = ~w8568 & w8571;
assign w8573 = (w8572 & ~w711) | (w8572 & w29177) | (~w711 & w29177);
assign w8574 = (w711 & w39622) | (w711 & w39623) | (w39622 & w39623);
assign w8575 = (~w711 & w39624) | (~w711 & w39625) | (w39624 & w39625);
assign w8576 = ~w8573 & ~w8574;
assign w8577 = ~w8575 & ~w8576;
assign w8578 = ~w8565 & w26798;
assign w8579 = (~w8577 & w8565) | (~w8577 & w26799) | (w8565 & w26799);
assign w8580 = ~w8578 & ~w8579;
assign w8581 = ~w8492 & w8580;
assign w8582 = w8492 & ~w8580;
assign w8583 = ~w8581 & ~w8582;
assign w8584 = ~w8491 & w8583;
assign w8585 = w8583 & ~w8584;
assign w8586 = ~w8583 & ~w8491;
assign w8587 = ~w8585 & ~w8586;
assign w8588 = ~w8321 & ~w8324;
assign w8589 = w8587 & w8588;
assign w8590 = ~w8587 & ~w8588;
assign w8591 = ~w8589 & ~w8590;
assign w8592 = b_19 & w3803;
assign w8593 = w4027 & w29178;
assign w8594 = b_18 & w3798;
assign w8595 = ~w8593 & ~w8594;
assign w8596 = ~w8592 & w8595;
assign w8597 = (w8596 & ~w1372) | (w8596 & w29179) | (~w1372 & w29179);
assign w8598 = (w1372 & w39626) | (w1372 & w39627) | (w39626 & w39627);
assign w8599 = (~w1372 & w39628) | (~w1372 & w39629) | (w39628 & w39629);
assign w8600 = ~w8597 & ~w8598;
assign w8601 = ~w8599 & ~w8600;
assign w8602 = w8591 & ~w8601;
assign w8603 = ~w8591 & w8601;
assign w8604 = (w8330 & w27042) | (w8330 & w27043) | (w27042 & w27043);
assign w8605 = ~w8481 & ~w8604;
assign w8606 = ~w8602 & ~w8604;
assign w8607 = ~w8604 & w27043;
assign w8608 = ~w8605 & ~w8607;
assign w8609 = b_22 & w3195;
assign w8610 = w3388 & w29180;
assign w8611 = b_21 & w3190;
assign w8612 = ~w8610 & ~w8611;
assign w8613 = ~w8609 & w8612;
assign w8614 = (w8613 & ~w1786) | (w8613 & w29181) | (~w1786 & w29181);
assign w8615 = (w1786 & w39630) | (w1786 & w39631) | (w39630 & w39631);
assign w8616 = (~w1786 & w39632) | (~w1786 & w39633) | (w39632 & w39633);
assign w8617 = ~w8614 & ~w8615;
assign w8618 = ~w8616 & ~w8617;
assign w8619 = ~w8608 & ~w8618;
assign w8620 = ~w8608 & ~w8619;
assign w8621 = w8608 & ~w8618;
assign w8622 = ~w8620 & ~w8621;
assign w8623 = (~w8343 & w8347) | (~w8343 & w26801) | (w8347 & w26801);
assign w8624 = w8622 & w8623;
assign w8625 = ~w8622 & ~w8623;
assign w8626 = ~w8624 & ~w8625;
assign w8627 = b_25 & w2639;
assign w8628 = w2820 & w29182;
assign w8629 = b_24 & w2634;
assign w8630 = ~w8628 & ~w8629;
assign w8631 = ~w8627 & w8630;
assign w8632 = (w8631 & ~w2108) | (w8631 & w29183) | (~w2108 & w29183);
assign w8633 = (w2108 & w39634) | (w2108 & w39635) | (w39634 & w39635);
assign w8634 = (~w2108 & w39636) | (~w2108 & w39637) | (w39636 & w39637);
assign w8635 = ~w8632 & ~w8633;
assign w8636 = ~w8634 & ~w8635;
assign w8637 = w8626 & ~w8636;
assign w8638 = w8626 & ~w8637;
assign w8639 = ~w8626 & ~w8636;
assign w8640 = ~w8638 & ~w8639;
assign w8641 = ~w8480 & w8640;
assign w8642 = w8480 & ~w8640;
assign w8643 = ~w8641 & ~w8642;
assign w8644 = b_28 & w2158;
assign w8645 = w2294 & w29184;
assign w8646 = b_27 & w2153;
assign w8647 = ~w8645 & ~w8646;
assign w8648 = ~w8644 & w8647;
assign w8649 = (w8648 & ~w2771) | (w8648 & w29185) | (~w2771 & w29185);
assign w8650 = (w2771 & w39638) | (w2771 & w39639) | (w39638 & w39639);
assign w8651 = (~w2771 & w39640) | (~w2771 & w39641) | (w39640 & w39641);
assign w8652 = ~w8649 & ~w8650;
assign w8653 = ~w8651 & ~w8652;
assign w8654 = ~w8643 & ~w8653;
assign w8655 = w8643 & w8653;
assign w8656 = ~w8654 & ~w8655;
assign w8657 = w8479 & ~w8656;
assign w8658 = ~w8479 & w8656;
assign w8659 = ~w8657 & ~w8658;
assign w8660 = b_31 & w1694;
assign w8661 = w1834 & w29186;
assign w8662 = b_30 & w1689;
assign w8663 = ~w8661 & ~w8662;
assign w8664 = ~w8660 & w8663;
assign w8665 = (w8664 & ~w3345) | (w8664 & w26592) | (~w3345 & w26592);
assign w8666 = (w3345 & w29187) | (w3345 & w29188) | (w29187 & w29188);
assign w8667 = (~w3345 & w29189) | (~w3345 & w29190) | (w29189 & w29190);
assign w8668 = ~w8665 & ~w8666;
assign w8669 = ~w8667 & ~w8668;
assign w8670 = w8659 & ~w8669;
assign w8671 = w8659 & ~w8670;
assign w8672 = ~w8659 & ~w8669;
assign w8673 = ~w8671 & ~w8672;
assign w8674 = (~w8384 & w8214) | (~w8384 & w26802) | (w8214 & w26802);
assign w8675 = w8673 & w8674;
assign w8676 = ~w8673 & ~w8674;
assign w8677 = ~w8675 & ~w8676;
assign w8678 = b_34 & w1295;
assign w8679 = w1422 & w29191;
assign w8680 = b_33 & w1290;
assign w8681 = ~w8679 & ~w8680;
assign w8682 = ~w8678 & w8681;
assign w8683 = (w8682 & ~w3967) | (w8682 & w26593) | (~w3967 & w26593);
assign w8684 = (w3967 & w29192) | (w3967 & w29193) | (w29192 & w29193);
assign w8685 = (~w3967 & w29194) | (~w3967 & w29195) | (w29194 & w29195);
assign w8686 = ~w8683 & ~w8684;
assign w8687 = ~w8685 & ~w8686;
assign w8688 = w8677 & ~w8687;
assign w8689 = w8677 & ~w8688;
assign w8690 = ~w8677 & ~w8687;
assign w8691 = ~w8689 & ~w8690;
assign w8692 = (~w8390 & w8203) | (~w8390 & w25401) | (w8203 & w25401);
assign w8693 = w8691 & w8692;
assign w8694 = ~w8691 & ~w8692;
assign w8695 = ~w8693 & ~w8694;
assign w8696 = b_37 & w986;
assign w8697 = w1069 & w29196;
assign w8698 = b_36 & w981;
assign w8699 = ~w8697 & ~w8698;
assign w8700 = ~w8696 & w8699;
assign w8701 = (w8700 & ~w4636) | (w8700 & w25402) | (~w4636 & w25402);
assign w8702 = (w4636 & w26594) | (w4636 & w26595) | (w26594 & w26595);
assign w8703 = (~w4636 & w29197) | (~w4636 & w29198) | (w29197 & w29198);
assign w8704 = ~w8701 & ~w8702;
assign w8705 = ~w8703 & ~w8704;
assign w8706 = w8695 & ~w8705;
assign w8707 = w8695 & ~w8706;
assign w8708 = ~w8695 & ~w8705;
assign w8709 = ~w8707 & ~w8708;
assign w8710 = (~w8079 & w27163) | (~w8079 & w27164) | (w27163 & w27164);
assign w8711 = w8709 & w8710;
assign w8712 = ~w8709 & ~w8710;
assign w8713 = ~w8711 & ~w8712;
assign w8714 = b_40 & w657;
assign w8715 = w754 & w29199;
assign w8716 = b_39 & w652;
assign w8717 = ~w8715 & ~w8716;
assign w8718 = ~w8714 & w8717;
assign w8719 = (w8718 & ~w5363) | (w8718 & w25080) | (~w5363 & w25080);
assign w8720 = (w5363 & w25403) | (w5363 & w25404) | (w25403 & w25404);
assign w8721 = (~w5363 & w29200) | (~w5363 & w29201) | (w29200 & w29201);
assign w8722 = ~w8719 & ~w8720;
assign w8723 = ~w8721 & ~w8722;
assign w8724 = w8713 & ~w8723;
assign w8725 = w8713 & ~w8724;
assign w8726 = ~w8713 & ~w8723;
assign w8727 = ~w8725 & ~w8726;
assign w8728 = (~w8423 & w8427) | (~w8423 & w25081) | (w8427 & w25081);
assign w8729 = w8727 & w8728;
assign w8730 = ~w8727 & ~w8728;
assign w8731 = ~w8729 & ~w8730;
assign w8732 = b_43 & w418;
assign w8733 = w481 & w29202;
assign w8734 = b_42 & w413;
assign w8735 = ~w8733 & ~w8734;
assign w8736 = ~w8732 & w8735;
assign w8737 = (w8736 & ~w5888) | (w8736 & w25405) | (~w5888 & w25405);
assign w8738 = (w5888 & w26596) | (w5888 & w26597) | (w26596 & w26597);
assign w8739 = (~w5888 & w29203) | (~w5888 & w29204) | (w29203 & w29204);
assign w8740 = ~w8737 & ~w8738;
assign w8741 = ~w8739 & ~w8740;
assign w8742 = w8731 & ~w8741;
assign w8743 = ~w8731 & w8741;
assign w8744 = (~w8444 & w26803) | (~w8444 & w26804) | (w26803 & w26804);
assign w8745 = (~w8742 & w8478) | (~w8742 & w26598) | (w8478 & w26598);
assign w8746 = w25406 & w8478;
assign w8747 = (~w8746 & w8744) | (~w8746 & w27540) | (w8744 & w27540);
assign w8748 = b_46 & w239;
assign w8749 = w266 & w29205;
assign w8750 = b_45 & w234;
assign w8751 = ~w8749 & ~w8750;
assign w8752 = ~w8748 & w8751;
assign w8753 = (w8752 & ~w6974) | (w8752 & w25407) | (~w6974 & w25407);
assign w8754 = (w6974 & w26599) | (w6974 & w26600) | (w26599 & w26600);
assign w8755 = (~w6974 & w29206) | (~w6974 & w29207) | (w29206 & w29207);
assign w8756 = ~w8753 & ~w8754;
assign w8757 = ~w8755 & ~w8756;
assign w8758 = (~w27540 & w27745) | (~w27540 & w27746) | (w27745 & w27746);
assign w8759 = ~w8747 & ~w8758;
assign w8760 = (~w27746 & w39642) | (~w27746 & w39643) | (w39642 & w39643);
assign w8761 = ~w8759 & ~w8760;
assign w8762 = (~w8448 & w8131) | (~w8448 & w29208) | (w8131 & w29208);
assign w8763 = w8761 & w8762;
assign w8764 = ~w8761 & ~w8762;
assign w8765 = ~w8763 & ~w8764;
assign w8766 = b_49 & w99;
assign w8767 = w136 & w29209;
assign w8768 = b_48 & w94;
assign w8769 = ~w8767 & ~w8768;
assign w8770 = ~w8766 & w8769;
assign w8771 = (w8770 & ~w7859) | (w8770 & w29210) | (~w7859 & w29210);
assign w8772 = (w7859 & w39644) | (w7859 & w39645) | (w39644 & w39645);
assign w8773 = (~w7859 & w39646) | (~w7859 & w39647) | (w39646 & w39647);
assign w8774 = ~w8771 & ~w8772;
assign w8775 = ~w8773 & ~w8774;
assign w8776 = w8765 & ~w8775;
assign w8777 = w8765 & ~w8776;
assign w8778 = ~w8765 & ~w8775;
assign w8779 = ~w8777 & ~w8778;
assign w8780 = ~w8477 & w8779;
assign w8781 = w8477 & ~w8779;
assign w8782 = ~w8780 & ~w8781;
assign w8783 = w8 & w29211;
assign w8784 = ~w8 & w29212;
assign w8785 = b_51 & w4;
assign w8786 = ~w8784 & ~w8785;
assign w8787 = ~w8783 & w8786;
assign w8788 = ~b_51 & ~b_52;
assign w8789 = b_51 & b_52;
assign w8790 = ~w8788 & ~w8789;
assign w8791 = (w4656 & w39648) | (w4656 & w39649) | (w39648 & w39649);
assign w8792 = (~w4656 & w39650) | (~w4656 & w39651) | (w39650 & w39651);
assign w8793 = ~w8791 & ~w8792;
assign w8794 = (w8787 & ~w8793) | (w8787 & w29218) | (~w8793 & w29218);
assign w8795 = (w8793 & w39652) | (w8793 & w39653) | (w39652 & w39653);
assign w8796 = (~w8793 & w39654) | (~w8793 & w39655) | (w39654 & w39655);
assign w8797 = ~w8794 & ~w8795;
assign w8798 = ~w8796 & ~w8797;
assign w8799 = ~w8782 & ~w8798;
assign w8800 = w8782 & w8798;
assign w8801 = ~w8799 & ~w8800;
assign w8802 = (w8801 & w8474) | (w8801 & w26805) | (w8474 & w26805);
assign w8803 = ~w8474 & w29219;
assign w8804 = ~w8802 & ~w8803;
assign w8805 = ~w8799 & ~w8802;
assign w8806 = (~w8776 & w8477) | (~w8776 & w29220) | (w8477 & w29220);
assign w8807 = b_35 & w1295;
assign w8808 = w1422 & w29221;
assign w8809 = b_34 & w1290;
assign w8810 = ~w8808 & ~w8809;
assign w8811 = ~w8807 & w8810;
assign w8812 = (w8811 & ~w4181) | (w8811 & w26601) | (~w4181 & w26601);
assign w8813 = (w4181 & w29222) | (w4181 & w29223) | (w29222 & w29223);
assign w8814 = (~w4181 & w29224) | (~w4181 & w29225) | (w29224 & w29225);
assign w8815 = ~w8812 & ~w8813;
assign w8816 = ~w8814 & ~w8815;
assign w8817 = (~w8670 & w8673) | (~w8670 & w26806) | (w8673 & w26806);
assign w8818 = b_32 & w1694;
assign w8819 = w1834 & w29226;
assign w8820 = b_31 & w1689;
assign w8821 = ~w8819 & ~w8820;
assign w8822 = ~w8818 & w8821;
assign w8823 = (w8822 & ~w3545) | (w8822 & w26602) | (~w3545 & w26602);
assign w8824 = (w3545 & w29227) | (w3545 & w29228) | (w29227 & w29228);
assign w8825 = (~w3545 & w29229) | (~w3545 & w29230) | (w29229 & w29230);
assign w8826 = ~w8823 & ~w8824;
assign w8827 = ~w8825 & ~w8826;
assign w8828 = (~w8654 & w8479) | (~w8654 & w26807) | (w8479 & w26807);
assign w8829 = b_29 & w2158;
assign w8830 = w2294 & w29231;
assign w8831 = b_28 & w2153;
assign w8832 = ~w8830 & ~w8831;
assign w8833 = ~w8829 & w8832;
assign w8834 = (w8833 & ~w2954) | (w8833 & w29232) | (~w2954 & w29232);
assign w8835 = (w2954 & w39656) | (w2954 & w39657) | (w39656 & w39657);
assign w8836 = (~w2954 & w39658) | (~w2954 & w39659) | (w39658 & w39659);
assign w8837 = ~w8834 & ~w8835;
assign w8838 = ~w8836 & ~w8837;
assign w8839 = (~w8637 & w8480) | (~w8637 & w26808) | (w8480 & w26808);
assign w8840 = (~w8619 & w8622) | (~w8619 & w39660) | (w8622 & w39660);
assign w8841 = b_23 & w3195;
assign w8842 = w3388 & w29233;
assign w8843 = b_22 & w3190;
assign w8844 = ~w8842 & ~w8843;
assign w8845 = ~w8841 & w8844;
assign w8846 = (w8845 & ~w1933) | (w8845 & w29234) | (~w1933 & w29234);
assign w8847 = (w1933 & w39661) | (w1933 & w39662) | (w39661 & w39662);
assign w8848 = (~w1933 & w39663) | (~w1933 & w39664) | (w39663 & w39664);
assign w8849 = ~w8846 & ~w8847;
assign w8850 = ~w8848 & ~w8849;
assign w8851 = (~w8584 & w8588) | (~w8584 & w26809) | (w8588 & w26809);
assign w8852 = b_17 & w4499;
assign w8853 = w4723 & w29235;
assign w8854 = b_16 & w4494;
assign w8855 = ~w8853 & ~w8854;
assign w8856 = ~w8852 & w8855;
assign w8857 = (w8856 & ~w1038) | (w8856 & w29236) | (~w1038 & w29236);
assign w8858 = (w1038 & w39665) | (w1038 & w39666) | (w39665 & w39666);
assign w8859 = (~w1038 & w39667) | (~w1038 & w39668) | (w39667 & w39668);
assign w8860 = ~w8857 & ~w8858;
assign w8861 = ~w8859 & ~w8860;
assign w8862 = (~w8579 & w8492) | (~w8579 & w26810) | (w8492 & w26810);
assign w8863 = b_14 & w5196;
assign w8864 = w5459 & w29237;
assign w8865 = b_13 & w5191;
assign w8866 = ~w8864 & ~w8865;
assign w8867 = ~w8863 & w8866;
assign w8868 = (w8867 & ~w735) | (w8867 & w29238) | (~w735 & w29238);
assign w8869 = (w735 & w39669) | (w735 & w39670) | (w39669 & w39670);
assign w8870 = (~w735 & w39671) | (~w735 & w39672) | (w39671 & w39672);
assign w8871 = ~w8868 & ~w8869;
assign w8872 = ~w8870 & ~w8871;
assign w8873 = b_11 & w5962;
assign w8874 = w6246 & w29239;
assign w8875 = b_10 & w5957;
assign w8876 = ~w8874 & ~w8875;
assign w8877 = ~w8873 & w8876;
assign w8878 = (w8877 & ~w530) | (w8877 & w29240) | (~w530 & w29240);
assign w8879 = (w530 & w39673) | (w530 & w39674) | (w39673 & w39674);
assign w8880 = (~w530 & w39675) | (~w530 & w39676) | (w39675 & w39676);
assign w8881 = ~w8878 & ~w8879;
assign w8882 = ~w8880 & ~w8881;
assign w8883 = (~w8544 & w8548) | (~w8544 & w26603) | (w8548 & w26603);
assign w8884 = ~w8539 & ~w8541;
assign w8885 = b_2 & w8526;
assign w8886 = w8271 & ~w8525;
assign w8887 = w8886 & w25408;
assign w8888 = b_1 & w8521;
assign w8889 = ~w8887 & ~w8888;
assign w8890 = ~w8885 & w8889;
assign w8891 = w35 & w8529;
assign w8892 = w8890 & ~w8891;
assign w8893 = (a_53 & ~w8890) | (a_53 & w25558) | (~w8890 & w25558);
assign w8894 = w8890 & w25817;
assign w8895 = ~w8892 & ~w8893;
assign w8896 = ~w8894 & ~w8895;
assign w8897 = ~w8535 & w8896;
assign w8898 = w8535 & ~w8896;
assign w8899 = ~w8897 & ~w8898;
assign w8900 = b_5 & w7613;
assign w8901 = w7941 & w26166;
assign w8902 = b_4 & w7608;
assign w8903 = ~w8901 & ~w8902;
assign w8904 = ~w8900 & w8903;
assign w8905 = w129 & w7616;
assign w8906 = w8904 & ~w8905;
assign w8907 = (a_50 & w8905) | (a_50 & w26167) | (w8905 & w26167);
assign w8908 = ~w8905 & w39677;
assign w8909 = ~w8906 & ~w8907;
assign w8910 = ~w8908 & ~w8909;
assign w8911 = w8899 & ~w8910;
assign w8912 = ~w8899 & w8910;
assign w8913 = (~w8912 & w8541) | (~w8912 & w25559) | (w8541 & w25559);
assign w8914 = ~w8911 & w8913;
assign w8915 = ~w8884 & ~w8914;
assign w8916 = ~w8913 & ~w8911;
assign w8917 = b_8 & w6761;
assign w8918 = w7075 & w29241;
assign w8919 = b_7 & w6756;
assign w8920 = ~w8918 & ~w8919;
assign w8921 = ~w8917 & w8920;
assign w8922 = ~w308 & w29242;
assign w8923 = (w8921 & ~w29242) | (w8921 & w39678) | (~w29242 & w39678);
assign w8924 = (w29242 & w39679) | (w29242 & w39680) | (w39679 & w39680);
assign w8925 = ~w8922 & w29244;
assign w8926 = ~w8923 & ~w8924;
assign w8927 = ~w8925 & ~w8926;
assign w8928 = ~w8915 & w26605;
assign w8929 = (~w8927 & w8915) | (~w8927 & w26606) | (w8915 & w26606);
assign w8930 = ~w8928 & ~w8929;
assign w8931 = ~w8883 & w8930;
assign w8932 = w8883 & ~w8930;
assign w8933 = ~w8931 & ~w8932;
assign w8934 = w8882 & ~w8933;
assign w8935 = ~w8882 & w8933;
assign w8936 = ~w8934 & ~w8935;
assign w8937 = ~w8566 & w8936;
assign w8938 = w8566 & ~w8936;
assign w8939 = ~w8937 & ~w8938;
assign w8940 = ~w8872 & w8939;
assign w8941 = w8939 & ~w8940;
assign w8942 = ~w8939 & ~w8872;
assign w8943 = ~w8941 & ~w8942;
assign w8944 = ~w8862 & ~w8943;
assign w8945 = w8862 & w8943;
assign w8946 = ~w8944 & ~w8945;
assign w8947 = ~w8861 & w8946;
assign w8948 = ~w8946 & ~w8861;
assign w8949 = w8946 & ~w8947;
assign w8950 = ~w8948 & ~w8949;
assign w8951 = ~w8851 & ~w8950;
assign w8952 = ~w8851 & ~w8951;
assign w8953 = w8851 & ~w8950;
assign w8954 = ~w8952 & ~w8953;
assign w8955 = b_20 & w3803;
assign w8956 = w4027 & w29245;
assign w8957 = b_19 & w3798;
assign w8958 = ~w8956 & ~w8957;
assign w8959 = ~w8955 & w8958;
assign w8960 = (w8959 & ~w1503) | (w8959 & w29246) | (~w1503 & w29246);
assign w8961 = (w1503 & w39681) | (w1503 & w39682) | (w39681 & w39682);
assign w8962 = (~w1503 & w39683) | (~w1503 & w39684) | (w39683 & w39684);
assign w8963 = ~w8960 & ~w8961;
assign w8964 = ~w8962 & ~w8963;
assign w8965 = (~w8964 & w8952) | (~w8964 & w26913) | (w8952 & w26913);
assign w8966 = ~w8954 & ~w8965;
assign w8967 = ~w26913 & w27044;
assign w8968 = ~w8966 & ~w8967;
assign w8969 = (~w8606 & w8966) | (~w8606 & w27165) | (w8966 & w27165);
assign w8970 = w8606 & w8968;
assign w8971 = ~w8969 & ~w8970;
assign w8972 = ~w8969 & w27232;
assign w8973 = ~w8971 & ~w8850;
assign w8974 = w8971 & ~w8972;
assign w8975 = ~w8973 & ~w8974;
assign w8976 = (~w8975 & w8625) | (~w8975 & w25560) | (w8625 & w25560);
assign w8977 = ~w8840 & ~w8976;
assign w8978 = b_26 & w2639;
assign w8979 = w2820 & w29247;
assign w8980 = b_25 & w2634;
assign w8981 = ~w8979 & ~w8980;
assign w8982 = ~w8978 & w8981;
assign w8983 = (w8982 & ~w2416) | (w8982 & w29248) | (~w2416 & w29248);
assign w8984 = (w2416 & w39685) | (w2416 & w39686) | (w39685 & w39686);
assign w8985 = (~w2416 & w39687) | (~w2416 & w39688) | (w39687 & w39688);
assign w8986 = ~w8983 & ~w8984;
assign w8987 = ~w8985 & ~w8986;
assign w8988 = ~w8977 & w27046;
assign w8989 = (~w8987 & w8977) | (~w8987 & w27047) | (w8977 & w27047);
assign w8990 = ~w8988 & ~w8989;
assign w8991 = ~w8839 & w8990;
assign w8992 = w8839 & ~w8990;
assign w8993 = ~w8991 & ~w8992;
assign w8994 = w8838 & ~w8993;
assign w8995 = ~w8838 & w8993;
assign w8996 = ~w8994 & ~w8995;
assign w8997 = ~w8828 & w8996;
assign w8998 = w8828 & ~w8996;
assign w8999 = ~w8997 & ~w8998;
assign w9000 = w8827 & ~w8999;
assign w9001 = ~w8827 & w8999;
assign w9002 = ~w9000 & ~w9001;
assign w9003 = (~w26806 & w27166) | (~w26806 & w27167) | (w27166 & w27167);
assign w9004 = (w26806 & w27168) | (w26806 & w27169) | (w27168 & w27169);
assign w9005 = ~w9003 & ~w9004;
assign w9006 = ~w8816 & w9005;
assign w9007 = w9005 & ~w9006;
assign w9008 = ~w9005 & ~w8816;
assign w9009 = ~w9007 & ~w9008;
assign w9010 = (~w8688 & w8691) | (~w8688 & w27420) | (w8691 & w27420);
assign w9011 = w9009 & w9010;
assign w9012 = ~w9009 & ~w9010;
assign w9013 = ~w9011 & ~w9012;
assign w9014 = b_38 & w986;
assign w9015 = w1069 & w29249;
assign w9016 = b_37 & w981;
assign w9017 = ~w9015 & ~w9016;
assign w9018 = ~w9014 & w9017;
assign w9019 = (w9018 & ~w4658) | (w9018 & w25409) | (~w4658 & w25409);
assign w9020 = (w4658 & w25561) | (w4658 & w25562) | (w25561 & w25562);
assign w9021 = (~w4658 & w29250) | (~w4658 & w29251) | (w29250 & w29251);
assign w9022 = ~w9019 & ~w9020;
assign w9023 = ~w9021 & ~w9022;
assign w9024 = w9013 & ~w9023;
assign w9025 = w9013 & ~w9024;
assign w9026 = ~w9013 & ~w9023;
assign w9027 = ~w9025 & ~w9026;
assign w9028 = (~w8706 & w8710) | (~w8706 & w25410) | (w8710 & w25410);
assign w9029 = w9027 & w9028;
assign w9030 = ~w9027 & ~w9028;
assign w9031 = ~w9029 & ~w9030;
assign w9032 = b_41 & w657;
assign w9033 = w754 & w29252;
assign w9034 = b_40 & w652;
assign w9035 = ~w9033 & ~w9034;
assign w9036 = ~w9032 & w9035;
assign w9037 = (w9036 & ~w5609) | (w9036 & w25082) | (~w5609 & w25082);
assign w9038 = (w5609 & w25411) | (w5609 & w25412) | (w25411 & w25412);
assign w9039 = (~w5609 & w25563) | (~w5609 & w25564) | (w25563 & w25564);
assign w9040 = ~w9037 & ~w9038;
assign w9041 = ~w9039 & ~w9040;
assign w9042 = w9031 & ~w9041;
assign w9043 = w9041 & w9031;
assign w9044 = ~w9031 & ~w9041;
assign w9045 = ~w9043 & ~w9044;
assign w9046 = (~w8724 & w8727) | (~w8724 & w27421) | (w8727 & w27421);
assign w9047 = w9045 & w9046;
assign w9048 = ~w9045 & ~w9046;
assign w9049 = ~w9047 & ~w9048;
assign w9050 = b_44 & w418;
assign w9051 = w481 & w29253;
assign w9052 = b_43 & w413;
assign w9053 = ~w9051 & ~w9052;
assign w9054 = ~w9050 & w9053;
assign w9055 = (w9054 & ~w6408) | (w9054 & w25413) | (~w6408 & w25413);
assign w9056 = (w6408 & w26607) | (w6408 & w26608) | (w26607 & w26608);
assign w9057 = (~w6408 & w29254) | (~w6408 & w29255) | (w29254 & w29255);
assign w9058 = ~w9055 & ~w9056;
assign w9059 = ~w9057 & ~w9058;
assign w9060 = w9049 & ~w9059;
assign w9061 = ~w9049 & w9059;
assign w9062 = ~w8745 & w25083;
assign w9063 = ~w8745 & ~w9062;
assign w9064 = (~w9060 & w8745) | (~w9060 & w26811) | (w8745 & w26811);
assign w9065 = (w26811 & w25083) | (w26811 & w27747) | (w25083 & w27747);
assign w9066 = ~w9063 & ~w9065;
assign w9067 = b_47 & w239;
assign w9068 = w266 & w29256;
assign w9069 = b_46 & w234;
assign w9070 = ~w9068 & ~w9069;
assign w9071 = ~w9067 & w9070;
assign w9072 = (w9071 & ~w6998) | (w9071 & w25414) | (~w6998 & w25414);
assign w9073 = (w6998 & w26609) | (w6998 & w26610) | (w26609 & w26610);
assign w9074 = (~w6998 & w29257) | (~w6998 & w29258) | (w29257 & w29258);
assign w9075 = ~w9072 & ~w9073;
assign w9076 = ~w9074 & ~w9075;
assign w9077 = (~w9076 & w9063) | (~w9076 & w39689) | (w9063 & w39689);
assign w9078 = ~w9066 & ~w9077;
assign w9079 = ~w9063 & w39690;
assign w9080 = ~w9078 & ~w9079;
assign w9081 = (~w8758 & w8761) | (~w8758 & w39691) | (w8761 & w39691);
assign w9082 = w9080 & w9081;
assign w9083 = ~w9080 & ~w9081;
assign w9084 = ~w9082 & ~w9083;
assign w9085 = b_50 & w99;
assign w9086 = w136 & w29259;
assign w9087 = b_49 & w94;
assign w9088 = ~w9086 & ~w9087;
assign w9089 = ~w9085 & w9088;
assign w9090 = (w9089 & ~w8162) | (w9089 & w29260) | (~w8162 & w29260);
assign w9091 = (w8162 & w39692) | (w8162 & w39693) | (w39692 & w39693);
assign w9092 = (~w8162 & w39694) | (~w8162 & w39695) | (w39694 & w39695);
assign w9093 = ~w9090 & ~w9091;
assign w9094 = ~w9092 & ~w9093;
assign w9095 = w9084 & ~w9094;
assign w9096 = ~w9084 & w9094;
assign w9097 = (~w8477 & w26812) | (~w8477 & w26813) | (w26812 & w26813);
assign w9098 = (~w26812 & w29262) | (~w26812 & w29263) | (w29262 & w29263);
assign w9099 = (~w26812 & w39696) | (~w26812 & w39697) | (w39696 & w39697);
assign w9100 = w8 & w29264;
assign w9101 = ~w8 & w29265;
assign w9102 = b_52 & w4;
assign w9103 = ~w9101 & ~w9102;
assign w9104 = ~w9100 & w9103;
assign w9105 = ~b_52 & ~b_53;
assign w9106 = b_52 & b_53;
assign w9107 = ~w9105 & ~w9106;
assign w9108 = (w4656 & w39698) | (w4656 & w39699) | (w39698 & w39699);
assign w9109 = (~w6406 & w29269) | (~w6406 & w29270) | (w29269 & w29270);
assign w9110 = ~w9108 & ~w9109;
assign w9111 = (w9109 & w39700) | (w9109 & w39701) | (w39700 & w39701);
assign w9112 = a_2 & ~w9111;
assign w9113 = w9111 & a_2;
assign w9114 = ~w9111 & ~w9112;
assign w9115 = ~w9113 & ~w9114;
assign w9116 = (w9115 & w9099) | (w9115 & w29272) | (w9099 & w29272);
assign w9117 = ~w9099 & w29273;
assign w9118 = ~w9116 & ~w9117;
assign w9119 = (~w9118 & w8802) | (~w9118 & w39702) | (w8802 & w39702);
assign w9120 = ~w8802 & w39703;
assign w9121 = ~w9119 & ~w9120;
assign w9122 = (~w9115 & w9099) | (~w9115 & w29274) | (w9099 & w29274);
assign w9123 = (~w9122 & w8805) | (~w9122 & w25085) | (w8805 & w25085);
assign w9124 = w8 & w29275;
assign w9125 = ~w8 & w29276;
assign w9126 = b_53 & w4;
assign w9127 = ~w9125 & ~w9126;
assign w9128 = ~w9124 & w9127;
assign w9129 = ~b_53 & ~b_54;
assign w9130 = b_53 & b_54;
assign w9131 = ~w9129 & ~w9130;
assign w9132 = (w4656 & w39704) | (w4656 & w39705) | (w39704 & w39705);
assign w9133 = (~w4656 & w39706) | (~w4656 & w39707) | (w39706 & w39707);
assign w9134 = ~w9132 & ~w9133;
assign w9135 = (w9128 & ~w9134) | (w9128 & w29282) | (~w9134 & w29282);
assign w9136 = (w9134 & w39708) | (w9134 & w39709) | (w39708 & w39709);
assign w9137 = (~w9134 & w39710) | (~w9134 & w39711) | (w39710 & w39711);
assign w9138 = ~w9135 & ~w9136;
assign w9139 = ~w9137 & ~w9138;
assign w9140 = b_45 & w418;
assign w9141 = w481 & w29283;
assign w9142 = b_44 & w413;
assign w9143 = ~w9141 & ~w9142;
assign w9144 = ~w9140 & w9143;
assign w9145 = (w9144 & ~w6682) | (w9144 & w25415) | (~w6682 & w25415);
assign w9146 = (w6682 & w25568) | (w6682 & w25569) | (w25568 & w25569);
assign w9147 = (~w6682 & w26611) | (~w6682 & w26612) | (w26611 & w26612);
assign w9148 = ~w9145 & ~w9146;
assign w9149 = ~w9147 & ~w9148;
assign w9150 = (~w9042 & w9046) | (~w9042 & w25416) | (w9046 & w25416);
assign w9151 = (~w9006 & w9010) | (~w9006 & w26816) | (w9010 & w26816);
assign w9152 = (~w9001 & w8817) | (~w9001 & w25570) | (w8817 & w25570);
assign w9153 = (~w8995 & w8828) | (~w8995 & w25571) | (w8828 & w25571);
assign w9154 = b_30 & w2158;
assign w9155 = w2294 & w29284;
assign w9156 = b_29 & w2153;
assign w9157 = ~w9155 & ~w9156;
assign w9158 = ~w9154 & w9157;
assign w9159 = (w9158 & ~w3138) | (w9158 & w29285) | (~w3138 & w29285);
assign w9160 = (w3138 & w39712) | (w3138 & w39713) | (w39712 & w39713);
assign w9161 = (~w3138 & w39714) | (~w3138 & w39715) | (w39714 & w39715);
assign w9162 = ~w9159 & ~w9160;
assign w9163 = ~w9161 & ~w9162;
assign w9164 = (~w8989 & w8839) | (~w8989 & w25572) | (w8839 & w25572);
assign w9165 = b_27 & w2639;
assign w9166 = w2820 & w29286;
assign w9167 = b_26 & w2634;
assign w9168 = ~w9166 & ~w9167;
assign w9169 = ~w9165 & w9168;
assign w9170 = (w9169 & ~w2582) | (w9169 & w29287) | (~w2582 & w29287);
assign w9171 = (w2582 & w39716) | (w2582 & w39717) | (w39716 & w39717);
assign w9172 = (~w2582 & w39718) | (~w2582 & w39719) | (w39718 & w39719);
assign w9173 = ~w9170 & ~w9171;
assign w9174 = ~w9172 & ~w9173;
assign w9175 = b_24 & w3195;
assign w9176 = w3388 & w29288;
assign w9177 = b_23 & w3190;
assign w9178 = ~w9176 & ~w9177;
assign w9179 = ~w9175 & w9178;
assign w9180 = (w9179 & ~w2083) | (w9179 & w29289) | (~w2083 & w29289);
assign w9181 = (w2083 & w39720) | (w2083 & w39721) | (w39720 & w39721);
assign w9182 = (~w2083 & w39722) | (~w2083 & w39723) | (w39722 & w39723);
assign w9183 = ~w9180 & ~w9181;
assign w9184 = ~w9182 & ~w9183;
assign w9185 = (~w8965 & w8968) | (~w8965 & w27048) | (w8968 & w27048);
assign w9186 = b_21 & w3803;
assign w9187 = w4027 & w29290;
assign w9188 = b_20 & w3798;
assign w9189 = ~w9187 & ~w9188;
assign w9190 = ~w9186 & w9189;
assign w9191 = (w9190 & ~w1634) | (w9190 & w29291) | (~w1634 & w29291);
assign w9192 = (w1634 & w39724) | (w1634 & w39725) | (w39724 & w39725);
assign w9193 = (~w1634 & w39726) | (~w1634 & w39727) | (w39726 & w39727);
assign w9194 = ~w9191 & ~w9192;
assign w9195 = ~w9193 & ~w9194;
assign w9196 = (~w8947 & w8851) | (~w8947 & w25573) | (w8851 & w25573);
assign w9197 = b_18 & w4499;
assign w9198 = w4723 & w29292;
assign w9199 = b_17 & w4494;
assign w9200 = ~w9198 & ~w9199;
assign w9201 = ~w9197 & w9200;
assign w9202 = (w9201 & ~w1238) | (w9201 & w25574) | (~w1238 & w25574);
assign w9203 = (w1238 & w29293) | (w1238 & w29294) | (w29293 & w29294);
assign w9204 = (~w1238 & w29295) | (~w1238 & w29296) | (w29295 & w29296);
assign w9205 = ~w9202 & ~w9203;
assign w9206 = ~w9204 & ~w9205;
assign w9207 = (~w8940 & w8862) | (~w8940 & w25575) | (w8862 & w25575);
assign w9208 = b_15 & w5196;
assign w9209 = w5459 & w29297;
assign w9210 = b_14 & w5191;
assign w9211 = ~w9209 & ~w9210;
assign w9212 = ~w9208 & w9211;
assign w9213 = (w9212 & ~w827) | (w9212 & w29298) | (~w827 & w29298);
assign w9214 = (w827 & w39728) | (w827 & w39729) | (w39728 & w39729);
assign w9215 = (~w827 & w39730) | (~w827 & w39731) | (w39730 & w39731);
assign w9216 = ~w9213 & ~w9214;
assign w9217 = ~w9215 & ~w9216;
assign w9218 = (~w8935 & w8566) | (~w8935 & w26817) | (w8566 & w26817);
assign w9219 = b_12 & w5962;
assign w9220 = w6246 & w29299;
assign w9221 = b_11 & w5957;
assign w9222 = ~w9220 & ~w9221;
assign w9223 = ~w9219 & w9222;
assign w9224 = (w9223 & ~w552) | (w9223 & w29300) | (~w552 & w29300);
assign w9225 = (w552 & w39732) | (w552 & w39733) | (w39732 & w39733);
assign w9226 = (~w552 & w39734) | (~w552 & w39735) | (w39734 & w39735);
assign w9227 = ~w9224 & ~w9225;
assign w9228 = ~w9226 & ~w9227;
assign w9229 = (~w8929 & w8883) | (~w8929 & w25576) | (w8883 & w25576);
assign w9230 = b_9 & w6761;
assign w9231 = w7075 & w29301;
assign w9232 = b_8 & w6756;
assign w9233 = ~w9231 & ~w9232;
assign w9234 = ~w9230 & w9233;
assign w9235 = (w9234 & ~w371) | (w9234 & w29302) | (~w371 & w29302);
assign w9236 = (w371 & w39736) | (w371 & w39737) | (w39736 & w39737);
assign w9237 = (~w371 & w39738) | (~w371 & w39739) | (w39738 & w39739);
assign w9238 = ~w9235 & ~w9236;
assign w9239 = ~w9237 & ~w9238;
assign w9240 = b_6 & w7613;
assign w9241 = w7941 & w29303;
assign w9242 = b_5 & w7608;
assign w9243 = ~w9241 & ~w9242;
assign w9244 = ~w9240 & w9243;
assign w9245 = (w9244 & ~w190) | (w9244 & w29304) | (~w190 & w29304);
assign w9246 = (w190 & w39740) | (w190 & w39741) | (w39740 & w39741);
assign w9247 = (~w190 & w39742) | (~w190 & w39743) | (w39742 & w39743);
assign w9248 = ~w9245 & ~w9246;
assign w9249 = ~w9247 & ~w9248;
assign w9250 = a_53 & ~a_54;
assign w9251 = ~a_53 & a_54;
assign w9252 = ~w9250 & ~w9251;
assign w9253 = b_0 & ~w9252;
assign w9254 = (w9253 & w8896) | (w9253 & w25818) | (w8896 & w25818);
assign w9255 = ~w8896 & w25819;
assign w9256 = ~w9254 & ~w9255;
assign w9257 = b_3 & w8526;
assign w9258 = w8886 & w25820;
assign w9259 = b_2 & w8521;
assign w9260 = ~w9258 & ~w9259;
assign w9261 = ~w9257 & w9260;
assign w9262 = w57 & w8529;
assign w9263 = w9261 & ~w9262;
assign w9264 = a_53 & ~w9263;
assign w9265 = w9263 & a_53;
assign w9266 = ~w9263 & ~w9264;
assign w9267 = ~w9265 & ~w9266;
assign w9268 = ~w9256 & ~w9267;
assign w9269 = w9256 & w9267;
assign w9270 = ~w9268 & ~w9269;
assign w9271 = ~w9249 & w9270;
assign w9272 = w9270 & ~w9271;
assign w9273 = ~w9270 & ~w9249;
assign w9274 = ~w9272 & ~w9273;
assign w9275 = ~w8916 & ~w9274;
assign w9276 = w8916 & w9274;
assign w9277 = ~w9275 & ~w9276;
assign w9278 = ~w9239 & w9277;
assign w9279 = ~w9277 & ~w9239;
assign w9280 = w9277 & ~w9278;
assign w9281 = ~w9279 & ~w9280;
assign w9282 = ~w9229 & ~w9281;
assign w9283 = w9229 & ~w9280;
assign w9284 = ~w9279 & w9283;
assign w9285 = ~w9282 & ~w9284;
assign w9286 = ~w9228 & w9285;
assign w9287 = ~w9285 & ~w9228;
assign w9288 = w9285 & ~w9286;
assign w9289 = ~w9287 & ~w9288;
assign w9290 = (~w9218 & w9288) | (~w9218 & w27347) | (w9288 & w27347);
assign w9291 = ~w9288 & w27348;
assign w9292 = ~w9290 & ~w9291;
assign w9293 = ~w9217 & w9292;
assign w9294 = w9217 & ~w9292;
assign w9295 = ~w9293 & ~w9294;
assign w9296 = ~w9207 & w9295;
assign w9297 = w9207 & ~w9295;
assign w9298 = ~w9296 & ~w9297;
assign w9299 = ~w9206 & w9298;
assign w9300 = ~w9298 & ~w9206;
assign w9301 = w9298 & ~w9299;
assign w9302 = ~w9300 & ~w9301;
assign w9303 = ~w9196 & ~w9302;
assign w9304 = w9196 & w9302;
assign w9305 = ~w9303 & ~w9304;
assign w9306 = ~w9195 & w9305;
assign w9307 = w9195 & ~w9305;
assign w9308 = ~w9306 & ~w9307;
assign w9309 = (~w8968 & w27170) | (~w8968 & w27171) | (w27170 & w27171);
assign w9310 = (w8968 & w27172) | (w8968 & w27173) | (w27172 & w27173);
assign w9311 = ~w9309 & ~w9310;
assign w9312 = ~w9184 & w9311;
assign w9313 = w9184 & ~w9311;
assign w9314 = ~w9312 & ~w9313;
assign w9315 = (~w8840 & w27422) | (~w8840 & w27423) | (w27422 & w27423);
assign w9316 = (w8840 & w27424) | (w8840 & w27425) | (w27424 & w27425);
assign w9317 = ~w9315 & ~w9316;
assign w9318 = ~w9174 & w9317;
assign w9319 = w9174 & ~w9317;
assign w9320 = ~w9318 & ~w9319;
assign w9321 = ~w9164 & w9320;
assign w9322 = w9164 & ~w9320;
assign w9323 = ~w9321 & ~w9322;
assign w9324 = ~w9163 & w9323;
assign w9325 = w9163 & ~w9323;
assign w9326 = ~w9324 & ~w9325;
assign w9327 = ~w9153 & w9326;
assign w9328 = w9153 & ~w9326;
assign w9329 = ~w9327 & ~w9328;
assign w9330 = b_33 & w1694;
assign w9331 = w1834 & w29305;
assign w9332 = b_32 & w1689;
assign w9333 = ~w9331 & ~w9332;
assign w9334 = ~w9330 & w9333;
assign w9335 = (w9334 & ~w3744) | (w9334 & w25577) | (~w3744 & w25577);
assign w9336 = (w3744 & w26613) | (w3744 & w26614) | (w26613 & w26614);
assign w9337 = (~w3744 & w29306) | (~w3744 & w29307) | (w29306 & w29307);
assign w9338 = ~w9335 & ~w9336;
assign w9339 = ~w9337 & ~w9338;
assign w9340 = w9329 & ~w9339;
assign w9341 = w9329 & ~w9340;
assign w9342 = ~w9329 & ~w9339;
assign w9343 = ~w9341 & ~w9342;
assign w9344 = ~w9152 & w9343;
assign w9345 = w9152 & ~w9343;
assign w9346 = ~w9344 & ~w9345;
assign w9347 = b_36 & w1295;
assign w9348 = w1422 & w29308;
assign w9349 = b_35 & w1290;
assign w9350 = ~w9348 & ~w9349;
assign w9351 = ~w9347 & w9350;
assign w9352 = (w9351 & ~w4395) | (w9351 & w26615) | (~w4395 & w26615);
assign w9353 = (w4395 & w29309) | (w4395 & w29310) | (w29309 & w29310);
assign w9354 = (~w4395 & w29311) | (~w4395 & w29312) | (w29311 & w29312);
assign w9355 = ~w9352 & ~w9353;
assign w9356 = ~w9354 & ~w9355;
assign w9357 = ~w9346 & ~w9356;
assign w9358 = w9346 & w9356;
assign w9359 = ~w9357 & ~w9358;
assign w9360 = w9151 & ~w9359;
assign w9361 = ~w9151 & w9359;
assign w9362 = ~w9360 & ~w9361;
assign w9363 = b_39 & w986;
assign w9364 = w1069 & w29313;
assign w9365 = b_38 & w981;
assign w9366 = ~w9364 & ~w9365;
assign w9367 = ~w9363 & w9366;
assign w9368 = (w9367 & ~w4888) | (w9367 & w25417) | (~w4888 & w25417);
assign w9369 = (w4888 & w25578) | (w4888 & w25579) | (w25578 & w25579);
assign w9370 = (~w4888 & w29314) | (~w4888 & w29315) | (w29314 & w29315);
assign w9371 = ~w9368 & ~w9369;
assign w9372 = ~w9370 & ~w9371;
assign w9373 = w9362 & ~w9372;
assign w9374 = w9362 & ~w9373;
assign w9375 = ~w9362 & ~w9372;
assign w9376 = ~w9374 & ~w9375;
assign w9377 = (~w9024 & w9027) | (~w9024 & w27233) | (w9027 & w27233);
assign w9378 = w9376 & w9377;
assign w9379 = ~w9376 & ~w9377;
assign w9380 = ~w9378 & ~w9379;
assign w9381 = b_42 & w657;
assign w9382 = w754 & w29316;
assign w9383 = b_41 & w652;
assign w9384 = ~w9382 & ~w9383;
assign w9385 = ~w9381 & w9384;
assign w9386 = (w9385 & ~w5864) | (w9385 & w25087) | (~w5864 & w25087);
assign w9387 = (w5864 & w25418) | (w5864 & w25419) | (w25418 & w25419);
assign w9388 = (~w5864 & w25580) | (~w5864 & w25581) | (w25580 & w25581);
assign w9389 = ~w9386 & ~w9387;
assign w9390 = ~w9388 & ~w9389;
assign w9391 = ~w9380 & w9390;
assign w9392 = w9380 & ~w9390;
assign w9393 = ~w9391 & ~w9392;
assign w9394 = ~w9150 & w9393;
assign w9395 = w9150 & ~w9393;
assign w9396 = ~w9394 & ~w9395;
assign w9397 = ~w9149 & w9396;
assign w9398 = ~w9396 & ~w9149;
assign w9399 = w9149 & w9396;
assign w9400 = ~w9398 & ~w9399;
assign w9401 = ~w9064 & ~w9400;
assign w9402 = ~w9064 & ~w9401;
assign w9403 = w9064 & ~w9400;
assign w9404 = ~w9402 & ~w9403;
assign w9405 = b_48 & w239;
assign w9406 = w266 & w29317;
assign w9407 = b_47 & w234;
assign w9408 = ~w9406 & ~w9407;
assign w9409 = ~w9405 & w9408;
assign w9410 = (w9409 & ~w7284) | (w9409 & w26616) | (~w7284 & w26616);
assign w9411 = (w7284 & w29318) | (w7284 & w29319) | (w29318 & w29319);
assign w9412 = (~w7284 & w29320) | (~w7284 & w29321) | (w29320 & w29321);
assign w9413 = ~w9410 & ~w9411;
assign w9414 = ~w9412 & ~w9413;
assign w9415 = (~w9414 & w9402) | (~w9414 & w27748) | (w9402 & w27748);
assign w9416 = ~w9404 & ~w9415;
assign w9417 = ~w9414 & ~w9415;
assign w9418 = ~w9416 & ~w9417;
assign w9419 = ~w9077 & ~w9083;
assign w9420 = ~w9083 & w29322;
assign w9421 = (~w9418 & w9083) | (~w9418 & w29323) | (w9083 & w29323);
assign w9422 = ~w9420 & ~w9421;
assign w9423 = b_51 & w99;
assign w9424 = w136 & w29324;
assign w9425 = b_50 & w94;
assign w9426 = ~w9424 & ~w9425;
assign w9427 = ~w9423 & w9426;
assign w9428 = (w9427 & ~w8186) | (w9427 & w29325) | (~w8186 & w29325);
assign w9429 = (w8186 & w39744) | (w8186 & w39745) | (w39744 & w39745);
assign w9430 = (~w8186 & w39746) | (~w8186 & w39747) | (w39746 & w39747);
assign w9431 = ~w9428 & ~w9429;
assign w9432 = ~w9430 & ~w9431;
assign w9433 = ~w9422 & w9432;
assign w9434 = w9422 & ~w9432;
assign w9435 = ~w9433 & ~w9434;
assign w9436 = (w9435 & w9097) | (w9435 & w27049) | (w9097 & w27049);
assign w9437 = w9098 & ~w9435;
assign w9438 = ~w9436 & ~w9437;
assign w9439 = ~w9139 & w9438;
assign w9440 = w9139 & ~w9438;
assign w9441 = ~w9439 & ~w9440;
assign w9442 = (~w8805 & w25582) | (~w8805 & w25583) | (w25582 & w25583);
assign w9443 = w9123 & ~w9441;
assign w9444 = ~w9442 & ~w9443;
assign w9445 = (~w9097 & w29326) | (~w9097 & w29327) | (w29326 & w29327);
assign w9446 = b_52 & w99;
assign w9447 = w136 & w29328;
assign w9448 = b_51 & w94;
assign w9449 = ~w9447 & ~w9448;
assign w9450 = ~w9446 & w9449;
assign w9451 = (w9450 & ~w8793) | (w9450 & w29329) | (~w8793 & w29329);
assign w9452 = (w8793 & w39748) | (w8793 & w39749) | (w39748 & w39749);
assign w9453 = (~w8793 & w39750) | (~w8793 & w39751) | (w39750 & w39751);
assign w9454 = ~w9451 & ~w9452;
assign w9455 = ~w9453 & ~w9454;
assign w9456 = b_49 & w239;
assign w9457 = w266 & w29330;
assign w9458 = b_48 & w234;
assign w9459 = ~w9457 & ~w9458;
assign w9460 = ~w9456 & w9459;
assign w9461 = (w9460 & ~w7859) | (w9460 & w25420) | (~w7859 & w25420);
assign w9462 = (w7859 & w29331) | (w7859 & w29332) | (w29331 & w29332);
assign w9463 = (~w7859 & w29333) | (~w7859 & w29334) | (w29333 & w29334);
assign w9464 = ~w9461 & ~w9462;
assign w9465 = ~w9463 & ~w9464;
assign w9466 = (~w9397 & w9064) | (~w9397 & w27749) | (w9064 & w27749);
assign w9467 = (~w9392 & w9150) | (~w9392 & w25088) | (w9150 & w25088);
assign w9468 = (~w9299 & w9196) | (~w9299 & w25089) | (w9196 & w25089);
assign w9469 = b_16 & w5196;
assign w9470 = w5459 & w29335;
assign w9471 = b_15 & w5191;
assign w9472 = ~w9470 & ~w9471;
assign w9473 = ~w9469 & w9472;
assign w9474 = (w9473 & ~w926) | (w9473 & w29336) | (~w926 & w29336);
assign w9475 = (w926 & w39752) | (w926 & w39753) | (w39752 & w39753);
assign w9476 = (~w926 & w39754) | (~w926 & w39755) | (w39754 & w39755);
assign w9477 = ~w9474 & ~w9475;
assign w9478 = ~w9476 & ~w9477;
assign w9479 = (~w9286 & w9289) | (~w9286 & w26914) | (w9289 & w26914);
assign w9480 = b_13 & w5962;
assign w9481 = w6246 & w29337;
assign w9482 = b_12 & w5957;
assign w9483 = ~w9481 & ~w9482;
assign w9484 = ~w9480 & w9483;
assign w9485 = (w9484 & ~w711) | (w9484 & w29338) | (~w711 & w29338);
assign w9486 = (w711 & w39756) | (w711 & w39757) | (w39756 & w39757);
assign w9487 = (~w711 & w39758) | (~w711 & w39759) | (w39758 & w39759);
assign w9488 = ~w9485 & ~w9486;
assign w9489 = ~w9487 & ~w9488;
assign w9490 = (~w9278 & w9281) | (~w9278 & w26617) | (w9281 & w26617);
assign w9491 = b_10 & w6761;
assign w9492 = w7075 & w29339;
assign w9493 = b_9 & w6756;
assign w9494 = ~w9492 & ~w9493;
assign w9495 = ~w9491 & w9494;
assign w9496 = (w9495 & ~w454) | (w9495 & w29340) | (~w454 & w29340);
assign w9497 = (w454 & w39760) | (w454 & w39761) | (w39760 & w39761);
assign w9498 = (~w454 & w39762) | (~w454 & w39763) | (w39762 & w39763);
assign w9499 = ~w9496 & ~w9497;
assign w9500 = ~w9498 & ~w9499;
assign w9501 = (~w9271 & w9274) | (~w9271 & w26168) | (w9274 & w26168);
assign w9502 = b_7 & w7613;
assign w9503 = w7941 & w29341;
assign w9504 = b_6 & w7608;
assign w9505 = ~w9503 & ~w9504;
assign w9506 = ~w9502 & w9505;
assign w9507 = (w9506 & ~w213) | (w9506 & w29342) | (~w213 & w29342);
assign w9508 = (w213 & w39764) | (w213 & w39765) | (w39764 & w39765);
assign w9509 = (~w213 & w39766) | (~w213 & w39767) | (w39766 & w39767);
assign w9510 = ~w9507 & ~w9508;
assign w9511 = ~w9509 & ~w9510;
assign w9512 = ~w8896 & w25821;
assign w9513 = (~w9512 & w9256) | (~w9512 & w25584) | (w9256 & w25584);
assign w9514 = b_4 & w8526;
assign w9515 = w8886 & w25822;
assign w9516 = b_3 & w8521;
assign w9517 = ~w9515 & ~w9516;
assign w9518 = ~w9514 & w9517;
assign w9519 = w84 & w8529;
assign w9520 = w9518 & ~w9519;
assign w9521 = (a_53 & w9519) | (a_53 & w25823) | (w9519 & w25823);
assign w9522 = ~w9519 & w26169;
assign w9523 = ~w9520 & ~w9521;
assign w9524 = ~w9522 & ~w9523;
assign w9525 = (a_56 & w9252) | (a_56 & w29343) | (w9252 & w29343);
assign w9526 = ~a_54 & a_55;
assign w9527 = a_54 & ~a_55;
assign w9528 = ~w9526 & ~w9527;
assign w9529 = w9252 & ~w9528;
assign w9530 = b_0 & w9529;
assign w9531 = ~a_55 & a_56;
assign w9532 = a_55 & ~a_56;
assign w9533 = ~w9531 & ~w9532;
assign w9534 = ~w9252 & w9533;
assign w9535 = b_1 & w9534;
assign w9536 = ~w9530 & ~w9535;
assign w9537 = ~w9252 & ~w9533;
assign w9538 = ~w15 & w9537;
assign w9539 = w9536 & ~w9538;
assign w9540 = (a_56 & ~w9536) | (a_56 & w25824) | (~w9536 & w25824);
assign w9541 = w9536 & w26170;
assign w9542 = ~w9539 & ~w9540;
assign w9543 = (w9525 & w9542) | (w9525 & w26171) | (w9542 & w26171);
assign w9544 = ~w9542 & w26172;
assign w9545 = ~w9543 & ~w9544;
assign w9546 = w9524 & ~w9545;
assign w9547 = ~w9524 & w9545;
assign w9548 = ~w9546 & ~w9547;
assign w9549 = ~w9513 & w9548;
assign w9550 = w9513 & ~w9548;
assign w9551 = ~w9549 & ~w9550;
assign w9552 = w9511 & ~w9551;
assign w9553 = ~w9511 & w9551;
assign w9554 = ~w9552 & ~w9553;
assign w9555 = ~w9501 & w9554;
assign w9556 = w9501 & ~w9554;
assign w9557 = ~w9555 & ~w9556;
assign w9558 = w9500 & ~w9557;
assign w9559 = ~w9500 & w9557;
assign w9560 = ~w9558 & ~w9559;
assign w9561 = ~w9490 & w9560;
assign w9562 = w9490 & ~w9560;
assign w9563 = ~w9561 & ~w9562;
assign w9564 = w9489 & ~w9563;
assign w9565 = ~w9489 & w9563;
assign w9566 = ~w9564 & ~w9565;
assign w9567 = ~w9479 & w9566;
assign w9568 = w9479 & ~w9566;
assign w9569 = ~w9567 & ~w9568;
assign w9570 = ~w9478 & w9569;
assign w9571 = w9569 & ~w9570;
assign w9572 = ~w9569 & ~w9478;
assign w9573 = ~w9571 & ~w9572;
assign w9574 = (~w9293 & w9207) | (~w9293 & w26915) | (w9207 & w26915);
assign w9575 = w9573 & w9574;
assign w9576 = ~w9573 & ~w9574;
assign w9577 = ~w9575 & ~w9576;
assign w9578 = b_19 & w4499;
assign w9579 = w4723 & w29344;
assign w9580 = b_18 & w4494;
assign w9581 = ~w9579 & ~w9580;
assign w9582 = ~w9578 & w9581;
assign w9583 = (w9582 & ~w1372) | (w9582 & w29345) | (~w1372 & w29345);
assign w9584 = (w1372 & w39768) | (w1372 & w39769) | (w39768 & w39769);
assign w9585 = (~w1372 & w39770) | (~w1372 & w39771) | (w39770 & w39771);
assign w9586 = ~w9583 & ~w9584;
assign w9587 = ~w9585 & ~w9586;
assign w9588 = w9577 & ~w9587;
assign w9589 = ~w9577 & w9587;
assign w9590 = (~w25089 & w26818) | (~w25089 & w26819) | (w26818 & w26819);
assign w9591 = (~w9468 & ~w9590) | (~w9468 & w27051) | (~w9590 & w27051);
assign w9592 = (~w26819 & w27349) | (~w26819 & w27350) | (w27349 & w27350);
assign w9593 = w27052 & ~w9590;
assign w9594 = ~w9591 & ~w9593;
assign w9595 = b_22 & w3803;
assign w9596 = w4027 & w29346;
assign w9597 = b_21 & w3798;
assign w9598 = ~w9596 & ~w9597;
assign w9599 = ~w9595 & w9598;
assign w9600 = (w9599 & ~w1786) | (w9599 & w29347) | (~w1786 & w29347);
assign w9601 = (w1786 & w39772) | (w1786 & w39773) | (w39772 & w39773);
assign w9602 = (~w1786 & w39774) | (~w1786 & w39775) | (w39774 & w39775);
assign w9603 = ~w9600 & ~w9601;
assign w9604 = ~w9602 & ~w9603;
assign w9605 = ~w9594 & ~w9604;
assign w9606 = ~w9594 & ~w9605;
assign w9607 = w9594 & ~w9604;
assign w9608 = ~w9606 & ~w9607;
assign w9609 = (~w9306 & w9185) | (~w9306 & w27053) | (w9185 & w27053);
assign w9610 = ~w9606 & w27351;
assign w9611 = (~w9609 & w9606) | (~w9609 & w27352) | (w9606 & w27352);
assign w9612 = ~w9610 & ~w9611;
assign w9613 = b_25 & w3195;
assign w9614 = w3388 & w29348;
assign w9615 = b_24 & w3190;
assign w9616 = ~w9614 & ~w9615;
assign w9617 = ~w9613 & w9616;
assign w9618 = (w9617 & ~w2108) | (w9617 & w29349) | (~w2108 & w29349);
assign w9619 = (w2108 & w39776) | (w2108 & w39777) | (w39776 & w39777);
assign w9620 = (~w2108 & w39778) | (~w2108 & w39779) | (w39778 & w39779);
assign w9621 = ~w9618 & ~w9619;
assign w9622 = ~w9620 & ~w9621;
assign w9623 = w9612 & ~w9622;
assign w9624 = w9612 & ~w9623;
assign w9625 = ~w9612 & ~w9622;
assign w9626 = ~w9624 & ~w9625;
assign w9627 = (w8840 & w25585) | (w8840 & w25586) | (w25585 & w25586);
assign w9628 = w9626 & w9627;
assign w9629 = ~w9626 & ~w9627;
assign w9630 = ~w9628 & ~w9629;
assign w9631 = b_28 & w2639;
assign w9632 = w2820 & w29350;
assign w9633 = b_27 & w2634;
assign w9634 = ~w9632 & ~w9633;
assign w9635 = ~w9631 & w9634;
assign w9636 = (w9635 & ~w2771) | (w9635 & w26618) | (~w2771 & w26618);
assign w9637 = (w2771 & w29351) | (w2771 & w29352) | (w29351 & w29352);
assign w9638 = (~w2771 & w29353) | (~w2771 & w29354) | (w29353 & w29354);
assign w9639 = ~w9636 & ~w9637;
assign w9640 = ~w9638 & ~w9639;
assign w9641 = w9630 & ~w9640;
assign w9642 = w9630 & ~w9641;
assign w9643 = ~w9630 & ~w9640;
assign w9644 = ~w9642 & ~w9643;
assign w9645 = (~w9318 & w9164) | (~w9318 & w27054) | (w9164 & w27054);
assign w9646 = w9644 & w9645;
assign w9647 = ~w9644 & ~w9645;
assign w9648 = ~w9646 & ~w9647;
assign w9649 = b_31 & w2158;
assign w9650 = w2294 & w29355;
assign w9651 = b_30 & w2153;
assign w9652 = ~w9650 & ~w9651;
assign w9653 = ~w9649 & w9652;
assign w9654 = (w9653 & ~w3345) | (w9653 & w26619) | (~w3345 & w26619);
assign w9655 = (w3345 & w29356) | (w3345 & w29357) | (w29356 & w29357);
assign w9656 = (~w3345 & w29358) | (~w3345 & w29359) | (w29358 & w29359);
assign w9657 = ~w9654 & ~w9655;
assign w9658 = ~w9656 & ~w9657;
assign w9659 = w9648 & ~w9658;
assign w9660 = w9648 & ~w9659;
assign w9661 = ~w9648 & ~w9658;
assign w9662 = ~w9660 & ~w9661;
assign w9663 = (~w9324 & w9153) | (~w9324 & w27055) | (w9153 & w27055);
assign w9664 = w9662 & w9663;
assign w9665 = ~w9662 & ~w9663;
assign w9666 = ~w9664 & ~w9665;
assign w9667 = b_34 & w1694;
assign w9668 = w1834 & w29360;
assign w9669 = b_33 & w1689;
assign w9670 = ~w9668 & ~w9669;
assign w9671 = ~w9667 & w9670;
assign w9672 = (w9671 & ~w3967) | (w9671 & w26620) | (~w3967 & w26620);
assign w9673 = (w3967 & w29361) | (w3967 & w29362) | (w29361 & w29362);
assign w9674 = (~w3967 & w29363) | (~w3967 & w29364) | (w29363 & w29364);
assign w9675 = ~w9672 & ~w9673;
assign w9676 = ~w9674 & ~w9675;
assign w9677 = w9666 & ~w9676;
assign w9678 = w9666 & ~w9677;
assign w9679 = ~w9666 & ~w9676;
assign w9680 = ~w9678 & ~w9679;
assign w9681 = (~w9340 & w9152) | (~w9340 & w27174) | (w9152 & w27174);
assign w9682 = w9680 & w9681;
assign w9683 = ~w9680 & ~w9681;
assign w9684 = ~w9682 & ~w9683;
assign w9685 = b_37 & w1295;
assign w9686 = w1422 & w29365;
assign w9687 = b_36 & w1290;
assign w9688 = ~w9686 & ~w9687;
assign w9689 = ~w9685 & w9688;
assign w9690 = (w9689 & ~w4636) | (w9689 & w25587) | (~w4636 & w25587);
assign w9691 = (w4636 & w26621) | (w4636 & w26622) | (w26621 & w26622);
assign w9692 = (~w4636 & w29366) | (~w4636 & w29367) | (w29366 & w29367);
assign w9693 = ~w9690 & ~w9691;
assign w9694 = ~w9692 & ~w9693;
assign w9695 = w9684 & ~w9694;
assign w9696 = w9684 & ~w9695;
assign w9697 = ~w9684 & ~w9694;
assign w9698 = ~w9696 & ~w9697;
assign w9699 = (~w9357 & w9151) | (~w9357 & w25588) | (w9151 & w25588);
assign w9700 = w9698 & w9699;
assign w9701 = ~w9698 & ~w9699;
assign w9702 = ~w9700 & ~w9701;
assign w9703 = b_40 & w986;
assign w9704 = w1069 & w29368;
assign w9705 = b_39 & w981;
assign w9706 = ~w9704 & ~w9705;
assign w9707 = ~w9703 & w9706;
assign w9708 = (w9707 & ~w5363) | (w9707 & w25421) | (~w5363 & w25421);
assign w9709 = (w5363 & w25589) | (w5363 & w25590) | (w25589 & w25590);
assign w9710 = (~w5363 & w26623) | (~w5363 & w26624) | (w26623 & w26624);
assign w9711 = ~w9708 & ~w9709;
assign w9712 = ~w9710 & ~w9711;
assign w9713 = w9702 & ~w9712;
assign w9714 = w9712 & w9702;
assign w9715 = ~w9702 & ~w9712;
assign w9716 = ~w9714 & ~w9715;
assign w9717 = (~w9373 & w9377) | (~w9373 & w26820) | (w9377 & w26820);
assign w9718 = w9716 & w9717;
assign w9719 = ~w9716 & ~w9717;
assign w9720 = ~w9718 & ~w9719;
assign w9721 = b_43 & w657;
assign w9722 = w754 & w29369;
assign w9723 = b_42 & w652;
assign w9724 = ~w9722 & ~w9723;
assign w9725 = ~w9721 & w9724;
assign w9726 = (w9725 & ~w5888) | (w9725 & w25091) | (~w5888 & w25091);
assign w9727 = (w5888 & w25422) | (w5888 & w25423) | (w25422 & w25423);
assign w9728 = (~w5888 & w25591) | (~w5888 & w25592) | (w25591 & w25592);
assign w9729 = ~w9726 & ~w9727;
assign w9730 = ~w9728 & ~w9729;
assign w9731 = w9720 & ~w9730;
assign w9732 = ~w9720 & w9730;
assign w9733 = ~w9467 & w25092;
assign w9734 = ~w9467 & ~w9733;
assign w9735 = (~w9731 & w9467) | (~w9731 & w27056) | (w9467 & w27056);
assign w9736 = b_46 & w418;
assign w9737 = w481 & w29370;
assign w9738 = b_45 & w413;
assign w9739 = ~w9737 & ~w9738;
assign w9740 = ~w9736 & w9739;
assign w9741 = (w9740 & ~w6974) | (w9740 & w25424) | (~w6974 & w25424);
assign w9742 = (w6974 & w25593) | (w6974 & w25594) | (w25593 & w25594);
assign w9743 = (~w6974 & w26625) | (~w6974 & w26626) | (w26625 & w26626);
assign w9744 = ~w9741 & ~w9742;
assign w9745 = ~w9743 & ~w9744;
assign w9746 = ~w9734 & w27828;
assign w9747 = (~w9745 & w9734) | (~w9745 & w27829) | (w9734 & w27829);
assign w9748 = ~w9746 & ~w9747;
assign w9749 = ~w9466 & w9748;
assign w9750 = w9466 & ~w9748;
assign w9751 = ~w9749 & ~w9750;
assign w9752 = w9465 & ~w9751;
assign w9753 = ~w9465 & w9751;
assign w9754 = ~w9752 & ~w9753;
assign w9755 = (w9754 & w9421) | (w9754 & w25093) | (w9421 & w25093);
assign w9756 = (w9419 & w29371) | (w9419 & w29372) | (w29371 & w29372);
assign w9757 = ~w9755 & ~w9756;
assign w9758 = ~w9455 & w9757;
assign w9759 = w9757 & ~w9758;
assign w9760 = ~w9757 & ~w9455;
assign w9761 = ~w9759 & ~w9760;
assign w9762 = ~w9445 & w9761;
assign w9763 = w9445 & ~w9761;
assign w9764 = ~w9762 & ~w9763;
assign w9765 = w8 & w29373;
assign w9766 = ~w8 & w29374;
assign w9767 = b_54 & w4;
assign w9768 = ~w9766 & ~w9767;
assign w9769 = ~w9765 & w9768;
assign w9770 = (~w6406 & w29375) | (~w6406 & w29376) | (w29375 & w29376);
assign w9771 = ~b_54 & ~b_55;
assign w9772 = b_54 & b_55;
assign w9773 = ~w9771 & ~w9772;
assign w9774 = (w6406 & w39780) | (w6406 & w39781) | (w39780 & w39781);
assign w9775 = (~w6406 & w39782) | (~w6406 & w39783) | (w39782 & w39783);
assign w9776 = ~w9774 & ~w9775;
assign w9777 = (w9769 & ~w9776) | (w9769 & w29377) | (~w9776 & w29377);
assign w9778 = (w9776 & w39784) | (w9776 & w39785) | (w39784 & w39785);
assign w9779 = (~w9776 & w39786) | (~w9776 & w39787) | (w39786 & w39787);
assign w9780 = ~w9777 & ~w9778;
assign w9781 = ~w9779 & ~w9780;
assign w9782 = ~w9764 & ~w9781;
assign w9783 = w9764 & w9781;
assign w9784 = ~w9782 & ~w9783;
assign w9785 = (w9784 & w9442) | (w9784 & w25095) | (w9442 & w25095);
assign w9786 = ~w9442 & w29378;
assign w9787 = ~w9785 & ~w9786;
assign w9788 = w8 & w29379;
assign w9789 = ~w8 & w29380;
assign w9790 = b_55 & w4;
assign w9791 = ~w9789 & ~w9790;
assign w9792 = ~w9788 & w9791;
assign w9793 = ~b_55 & ~b_56;
assign w9794 = b_55 & b_56;
assign w9795 = ~w9793 & ~w9794;
assign w9796 = (w6406 & w39788) | (w6406 & w39789) | (w39788 & w39789);
assign w9797 = (~w6406 & w39790) | (~w6406 & w39791) | (w39790 & w39791);
assign w9798 = ~w9796 & ~w9797;
assign w9799 = (w9792 & ~w9798) | (w9792 & w29386) | (~w9798 & w29386);
assign w9800 = (w9798 & w39792) | (w9798 & w39793) | (w39792 & w39793);
assign w9801 = (~w9798 & w39794) | (~w9798 & w39795) | (w39794 & w39795);
assign w9802 = ~w9799 & ~w9800;
assign w9803 = ~w9801 & ~w9802;
assign w9804 = (~w9758 & w9445) | (~w9758 & w25096) | (w9445 & w25096);
assign w9805 = ~w9753 & ~w9755;
assign w9806 = b_50 & w239;
assign w9807 = w266 & w29387;
assign w9808 = b_49 & w234;
assign w9809 = ~w9807 & ~w9808;
assign w9810 = ~w9806 & w9809;
assign w9811 = (w9810 & ~w8162) | (w9810 & w29388) | (~w8162 & w29388);
assign w9812 = (w8162 & w39796) | (w8162 & w39797) | (w39796 & w39797);
assign w9813 = (~w8162 & w39798) | (~w8162 & w39799) | (w39798 & w39799);
assign w9814 = ~w9811 & ~w9812;
assign w9815 = ~w9813 & ~w9814;
assign w9816 = (~w9747 & w9466) | (~w9747 & w25097) | (w9466 & w25097);
assign w9817 = b_35 & w1694;
assign w9818 = w1834 & w29389;
assign w9819 = b_34 & w1689;
assign w9820 = ~w9818 & ~w9819;
assign w9821 = ~w9817 & w9820;
assign w9822 = (w9821 & ~w4181) | (w9821 & w25595) | (~w4181 & w25595);
assign w9823 = (w4181 & w26627) | (w4181 & w26628) | (w26627 & w26628);
assign w9824 = (~w4181 & w29390) | (~w4181 & w29391) | (w29390 & w29391);
assign w9825 = ~w9822 & ~w9823;
assign w9826 = ~w9824 & ~w9825;
assign w9827 = b_32 & w2158;
assign w9828 = w2294 & w29392;
assign w9829 = b_31 & w2153;
assign w9830 = ~w9828 & ~w9829;
assign w9831 = ~w9827 & w9830;
assign w9832 = (w9831 & ~w3545) | (w9831 & w25596) | (~w3545 & w25596);
assign w9833 = (w3545 & w26629) | (w3545 & w26630) | (w26629 & w26630);
assign w9834 = (~w3545 & w29393) | (~w3545 & w29394) | (w29393 & w29394);
assign w9835 = ~w9832 & ~w9833;
assign w9836 = ~w9834 & ~w9835;
assign w9837 = (~w9641 & w9645) | (~w9641 & w25098) | (w9645 & w25098);
assign w9838 = ~w9623 & ~w9629;
assign w9839 = (~w9605 & w9608) | (~w9605 & w27234) | (w9608 & w27234);
assign w9840 = (~w9570 & w9573) | (~w9570 & w27353) | (w9573 & w27353);
assign w9841 = b_17 & w5196;
assign w9842 = w5459 & w29395;
assign w9843 = b_16 & w5191;
assign w9844 = ~w9842 & ~w9843;
assign w9845 = ~w9841 & w9844;
assign w9846 = (w9845 & ~w1038) | (w9845 & w29396) | (~w1038 & w29396);
assign w9847 = (w1038 & w39800) | (w1038 & w39801) | (w39800 & w39801);
assign w9848 = (~w1038 & w39802) | (~w1038 & w39803) | (w39802 & w39803);
assign w9849 = ~w9846 & ~w9847;
assign w9850 = ~w9848 & ~w9849;
assign w9851 = (~w9565 & w9479) | (~w9565 & w27057) | (w9479 & w27057);
assign w9852 = b_14 & w5962;
assign w9853 = w6246 & w29397;
assign w9854 = b_13 & w5957;
assign w9855 = ~w9853 & ~w9854;
assign w9856 = ~w9852 & w9855;
assign w9857 = (w9856 & ~w735) | (w9856 & w29398) | (~w735 & w29398);
assign w9858 = (w735 & w39804) | (w735 & w39805) | (w39804 & w39805);
assign w9859 = (~w735 & w39806) | (~w735 & w39807) | (w39806 & w39807);
assign w9860 = ~w9857 & ~w9858;
assign w9861 = ~w9859 & ~w9860;
assign w9862 = (~w9559 & w9490) | (~w9559 & w26821) | (w9490 & w26821);
assign w9863 = b_11 & w6761;
assign w9864 = w7075 & w29399;
assign w9865 = b_10 & w6756;
assign w9866 = ~w9864 & ~w9865;
assign w9867 = ~w9863 & w9866;
assign w9868 = (w9867 & ~w530) | (w9867 & w29400) | (~w530 & w29400);
assign w9869 = (w530 & w39808) | (w530 & w39809) | (w39808 & w39809);
assign w9870 = (~w530 & w39810) | (~w530 & w39811) | (w39810 & w39811);
assign w9871 = ~w9868 & ~w9869;
assign w9872 = ~w9870 & ~w9871;
assign w9873 = (~w9553 & w9501) | (~w9553 & w26631) | (w9501 & w26631);
assign w9874 = ~w9547 & ~w9549;
assign w9875 = b_2 & w9534;
assign w9876 = w9252 & ~w9533;
assign w9877 = w9876 & w25597;
assign w9878 = b_1 & w9529;
assign w9879 = ~w9877 & ~w9878;
assign w9880 = ~w9875 & w9879;
assign w9881 = w35 & w9537;
assign w9882 = w9880 & ~w9881;
assign w9883 = (a_56 & ~w9880) | (a_56 & w25825) | (~w9880 & w25825);
assign w9884 = w9880 & w26173;
assign w9885 = ~w9882 & ~w9883;
assign w9886 = ~w9884 & ~w9885;
assign w9887 = ~w9543 & w9886;
assign w9888 = w9543 & ~w9886;
assign w9889 = ~w9887 & ~w9888;
assign w9890 = b_5 & w8526;
assign w9891 = w8886 & w26174;
assign w9892 = b_4 & w8521;
assign w9893 = ~w9891 & ~w9892;
assign w9894 = ~w9890 & w9893;
assign w9895 = w129 & w8529;
assign w9896 = w9894 & ~w9895;
assign w9897 = (a_53 & w9895) | (a_53 & w26175) | (w9895 & w26175);
assign w9898 = ~w9895 & w39812;
assign w9899 = ~w9896 & ~w9897;
assign w9900 = ~w9898 & ~w9899;
assign w9901 = w9889 & ~w9900;
assign w9902 = ~w9889 & w9900;
assign w9903 = (~w9902 & w9549) | (~w9902 & w25826) | (w9549 & w25826);
assign w9904 = ~w9901 & w9903;
assign w9905 = ~w9874 & ~w9904;
assign w9906 = ~w9903 & ~w9901;
assign w9907 = b_8 & w7613;
assign w9908 = w7941 & w29401;
assign w9909 = b_7 & w7608;
assign w9910 = ~w9908 & ~w9909;
assign w9911 = ~w9907 & w9910;
assign w9912 = ~w308 & w29402;
assign w9913 = (w9911 & ~w29402) | (w9911 & w39813) | (~w29402 & w39813);
assign w9914 = (w29402 & w39814) | (w29402 & w39815) | (w39814 & w39815);
assign w9915 = ~w9912 & w29404;
assign w9916 = ~w9913 & ~w9914;
assign w9917 = ~w9915 & ~w9916;
assign w9918 = ~w9905 & w26633;
assign w9919 = (~w9917 & w9905) | (~w9917 & w26634) | (w9905 & w26634);
assign w9920 = ~w9918 & ~w9919;
assign w9921 = ~w9873 & w9920;
assign w9922 = w9873 & ~w9920;
assign w9923 = ~w9921 & ~w9922;
assign w9924 = w9872 & ~w9923;
assign w9925 = ~w9872 & w9923;
assign w9926 = ~w9924 & ~w9925;
assign w9927 = ~w9862 & w9926;
assign w9928 = w9862 & ~w9926;
assign w9929 = ~w9927 & ~w9928;
assign w9930 = ~w9861 & w9929;
assign w9931 = w9929 & ~w9930;
assign w9932 = ~w9929 & ~w9861;
assign w9933 = ~w9931 & ~w9932;
assign w9934 = ~w9851 & ~w9933;
assign w9935 = w9851 & w9933;
assign w9936 = ~w9934 & ~w9935;
assign w9937 = ~w9850 & w9936;
assign w9938 = ~w9936 & ~w9850;
assign w9939 = w9936 & ~w9937;
assign w9940 = ~w9938 & ~w9939;
assign w9941 = ~w9840 & ~w9940;
assign w9942 = ~w9840 & ~w9941;
assign w9943 = w9840 & ~w9940;
assign w9944 = ~w9942 & ~w9943;
assign w9945 = b_20 & w4499;
assign w9946 = w4723 & w29405;
assign w9947 = b_19 & w4494;
assign w9948 = ~w9946 & ~w9947;
assign w9949 = ~w9945 & w9948;
assign w9950 = (w9949 & ~w1503) | (w9949 & w29406) | (~w1503 & w29406);
assign w9951 = (w1503 & w39816) | (w1503 & w39817) | (w39816 & w39817);
assign w9952 = (~w1503 & w39818) | (~w1503 & w39819) | (w39818 & w39819);
assign w9953 = ~w9950 & ~w9951;
assign w9954 = ~w9952 & ~w9953;
assign w9955 = (~w9954 & w9942) | (~w9954 & w27058) | (w9942 & w27058);
assign w9956 = ~w9944 & ~w9955;
assign w9957 = ~w9942 & w27426;
assign w9958 = ~w9956 & ~w9957;
assign w9959 = ~w9592 & w9958;
assign w9960 = w9592 & ~w9958;
assign w9961 = ~w9959 & ~w9960;
assign w9962 = b_23 & w3803;
assign w9963 = w4027 & w29407;
assign w9964 = b_22 & w3798;
assign w9965 = ~w9963 & ~w9964;
assign w9966 = ~w9962 & w9965;
assign w9967 = (w9966 & ~w1933) | (w9966 & w29408) | (~w1933 & w29408);
assign w9968 = (w1933 & w39820) | (w1933 & w39821) | (w39820 & w39821);
assign w9969 = (~w1933 & w39822) | (~w1933 & w39823) | (w39822 & w39823);
assign w9970 = ~w9967 & ~w9968;
assign w9971 = ~w9969 & ~w9970;
assign w9972 = ~w9961 & ~w9971;
assign w9973 = w9961 & w9971;
assign w9974 = ~w9972 & ~w9973;
assign w9975 = w9839 & ~w9974;
assign w9976 = (w9974 & w9611) | (w9974 & w25827) | (w9611 & w25827);
assign w9977 = ~w9975 & ~w9976;
assign w9978 = b_26 & w3195;
assign w9979 = w3388 & w29409;
assign w9980 = b_25 & w3190;
assign w9981 = ~w9979 & ~w9980;
assign w9982 = ~w9978 & w9981;
assign w9983 = (w9982 & ~w2416) | (w9982 & w25828) | (~w2416 & w25828);
assign w9984 = (w2416 & w29410) | (w2416 & w29411) | (w29410 & w29411);
assign w9985 = (~w2416 & w29412) | (~w2416 & w29413) | (w29412 & w29413);
assign w9986 = ~w9983 & ~w9984;
assign w9987 = ~w9985 & ~w9986;
assign w9988 = ~w9976 & w27235;
assign w9989 = (w9987 & w9976) | (w9987 & w27236) | (w9976 & w27236);
assign w9990 = (w9629 & w25829) | (w9629 & w25830) | (w25829 & w25830);
assign w9991 = ~w9838 & ~w9990;
assign w9992 = (~w9629 & w27059) | (~w9629 & w27060) | (w27059 & w27060);
assign w9993 = w27237 & w27060;
assign w9994 = ~w9991 & ~w9993;
assign w9995 = b_29 & w2639;
assign w9996 = w2820 & w29414;
assign w9997 = b_28 & w2634;
assign w9998 = ~w9996 & ~w9997;
assign w9999 = ~w9995 & w9998;
assign w10000 = (w9999 & ~w2954) | (w9999 & w29415) | (~w2954 & w29415);
assign w10001 = (w2954 & w39824) | (w2954 & w39825) | (w39824 & w39825);
assign w10002 = (~w2954 & w39826) | (~w2954 & w39827) | (w39826 & w39827);
assign w10003 = ~w10000 & ~w10001;
assign w10004 = ~w10002 & ~w10003;
assign w10005 = w9994 & w10004;
assign w10006 = ~w9994 & ~w10004;
assign w10007 = ~w10005 & ~w10006;
assign w10008 = ~w9837 & w10007;
assign w10009 = w9837 & ~w10007;
assign w10010 = ~w10008 & ~w10009;
assign w10011 = w9836 & ~w10010;
assign w10012 = ~w9836 & w10010;
assign w10013 = ~w10011 & ~w10012;
assign w10014 = (w10013 & w9665) | (w10013 & w25100) | (w9665 & w25100);
assign w10015 = ~w9665 & w25101;
assign w10016 = ~w10014 & ~w10015;
assign w10017 = ~w9826 & w10016;
assign w10018 = w10016 & ~w10017;
assign w10019 = ~w10016 & ~w9826;
assign w10020 = ~w10018 & ~w10019;
assign w10021 = (~w9677 & w9681) | (~w9677 & w27061) | (w9681 & w27061);
assign w10022 = w10020 & w10021;
assign w10023 = ~w10020 & ~w10021;
assign w10024 = ~w10022 & ~w10023;
assign w10025 = b_38 & w1295;
assign w10026 = w1422 & w29416;
assign w10027 = b_37 & w1290;
assign w10028 = ~w10026 & ~w10027;
assign w10029 = ~w10025 & w10028;
assign w10030 = (w10029 & ~w4658) | (w10029 & w25598) | (~w4658 & w25598);
assign w10031 = (w4658 & w25831) | (w4658 & w25832) | (w25831 & w25832);
assign w10032 = (~w4658 & w29417) | (~w4658 & w29418) | (w29417 & w29418);
assign w10033 = ~w10030 & ~w10031;
assign w10034 = ~w10032 & ~w10033;
assign w10035 = w10024 & ~w10034;
assign w10036 = w10024 & ~w10035;
assign w10037 = ~w10024 & ~w10034;
assign w10038 = ~w10036 & ~w10037;
assign w10039 = (~w9695 & w9698) | (~w9695 & w27750) | (w9698 & w27750);
assign w10040 = w10038 & w10039;
assign w10041 = ~w10038 & ~w10039;
assign w10042 = ~w10040 & ~w10041;
assign w10043 = b_41 & w986;
assign w10044 = w1069 & w29419;
assign w10045 = b_40 & w981;
assign w10046 = ~w10044 & ~w10045;
assign w10047 = ~w10043 & w10046;
assign w10048 = (w10047 & ~w5609) | (w10047 & w25425) | (~w5609 & w25425);
assign w10049 = (w5609 & w25599) | (w5609 & w25600) | (w25599 & w25600);
assign w10050 = (~w5609 & w25833) | (~w5609 & w25834) | (w25833 & w25834);
assign w10051 = ~w10048 & ~w10049;
assign w10052 = ~w10050 & ~w10051;
assign w10053 = w10042 & ~w10052;
assign w10054 = w10052 & w10042;
assign w10055 = ~w10042 & ~w10052;
assign w10056 = ~w10054 & ~w10055;
assign w10057 = (~w9713 & w9717) | (~w9713 & w25601) | (w9717 & w25601);
assign w10058 = w10056 & w10057;
assign w10059 = ~w10056 & ~w10057;
assign w10060 = ~w10058 & ~w10059;
assign w10061 = b_44 & w657;
assign w10062 = w754 & w29420;
assign w10063 = b_43 & w652;
assign w10064 = ~w10062 & ~w10063;
assign w10065 = ~w10061 & w10064;
assign w10066 = (w10065 & ~w6408) | (w10065 & w25102) | (~w6408 & w25102);
assign w10067 = (w6408 & w25426) | (w6408 & w25427) | (w25426 & w25427);
assign w10068 = (~w6408 & w25602) | (~w6408 & w25603) | (w25602 & w25603);
assign w10069 = ~w10066 & ~w10067;
assign w10070 = ~w10068 & ~w10069;
assign w10071 = w10060 & ~w10070;
assign w10072 = ~w10060 & w10070;
assign w10073 = ~w9735 & w25103;
assign w10074 = ~w9735 & ~w10073;
assign w10075 = ~w10071 & ~w10073;
assign w10076 = ~w10073 & w25103;
assign w10077 = ~w10074 & ~w10076;
assign w10078 = b_47 & w418;
assign w10079 = w481 & w29421;
assign w10080 = b_46 & w413;
assign w10081 = ~w10079 & ~w10080;
assign w10082 = ~w10078 & w10081;
assign w10083 = (w10082 & ~w6998) | (w10082 & w25104) | (~w6998 & w25104);
assign w10084 = (w6998 & w25428) | (w6998 & w25429) | (w25428 & w25429);
assign w10085 = (~w6998 & w25604) | (~w6998 & w25605) | (w25604 & w25605);
assign w10086 = ~w10083 & ~w10084;
assign w10087 = ~w10085 & ~w10086;
assign w10088 = ~w10077 & ~w10087;
assign w10089 = w10087 & ~w10077;
assign w10090 = w10077 & ~w10087;
assign w10091 = ~w10089 & ~w10090;
assign w10092 = ~w9816 & ~w10091;
assign w10093 = w9816 & w10091;
assign w10094 = ~w10092 & ~w10093;
assign w10095 = ~w9815 & w10094;
assign w10096 = ~w10094 & ~w9815;
assign w10097 = w10094 & ~w10095;
assign w10098 = ~w10096 & ~w10097;
assign w10099 = ~w9805 & ~w10098;
assign w10100 = ~w9805 & ~w10099;
assign w10101 = b_53 & w99;
assign w10102 = w136 & w29422;
assign w10103 = b_52 & w94;
assign w10104 = ~w10102 & ~w10103;
assign w10105 = ~w10101 & w10104;
assign w10106 = (w9109 & w39828) | (w9109 & w39829) | (w39828 & w39829);
assign w10107 = a_5 & ~w10106;
assign w10108 = w10106 & a_5;
assign w10109 = ~w10106 & ~w10107;
assign w10110 = ~w10108 & ~w10109;
assign w10111 = ~w10100 & w25835;
assign w10112 = (~w10110 & w10100) | (~w10110 & w25836) | (w10100 & w25836);
assign w10113 = ~w10111 & ~w10112;
assign w10114 = ~w9804 & w10113;
assign w10115 = w9804 & ~w10113;
assign w10116 = ~w10114 & ~w10115;
assign w10117 = ~w9803 & w10116;
assign w10118 = w10116 & ~w10117;
assign w10119 = ~w10116 & ~w9803;
assign w10120 = ~w10118 & ~w10119;
assign w10121 = (~w9442 & w27062) | (~w9442 & w27063) | (w27062 & w27063);
assign w10122 = ~w10120 & ~w10121;
assign w10123 = w10120 & w10121;
assign w10124 = ~w10122 & ~w10123;
assign w10125 = (~w10112 & w9804) | (~w10112 & w25105) | (w9804 & w25105);
assign w10126 = b_54 & w99;
assign w10127 = w136 & w29424;
assign w10128 = b_53 & w94;
assign w10129 = ~w10127 & ~w10128;
assign w10130 = ~w10126 & w10129;
assign w10131 = (w10130 & ~w9134) | (w10130 & w29425) | (~w9134 & w29425);
assign w10132 = (w9134 & w39830) | (w9134 & w39831) | (w39830 & w39831);
assign w10133 = (~w9134 & w39832) | (~w9134 & w39833) | (w39832 & w39833);
assign w10134 = ~w10131 & ~w10132;
assign w10135 = ~w10133 & ~w10134;
assign w10136 = (~w10095 & w9805) | (~w10095 & w25106) | (w9805 & w25106);
assign w10137 = b_51 & w239;
assign w10138 = w266 & w29426;
assign w10139 = b_50 & w234;
assign w10140 = ~w10138 & ~w10139;
assign w10141 = ~w10137 & w10140;
assign w10142 = (w10141 & ~w8186) | (w10141 & w29427) | (~w8186 & w29427);
assign w10143 = (w8186 & w39834) | (w8186 & w39835) | (w39834 & w39835);
assign w10144 = (~w8186 & w39836) | (~w8186 & w39837) | (w39836 & w39837);
assign w10145 = ~w10142 & ~w10143;
assign w10146 = ~w10144 & ~w10145;
assign w10147 = (~w10088 & w10091) | (~w10088 & w25606) | (w10091 & w25606);
assign w10148 = b_48 & w418;
assign w10149 = w481 & w29428;
assign w10150 = b_47 & w413;
assign w10151 = ~w10149 & ~w10150;
assign w10152 = ~w10148 & w10151;
assign w10153 = (w10152 & ~w7284) | (w10152 & w25430) | (~w7284 & w25430);
assign w10154 = (w7284 & w25607) | (w7284 & w25608) | (w25607 & w25608);
assign w10155 = (~w7284 & w25837) | (~w7284 & w25838) | (w25837 & w25838);
assign w10156 = ~w10153 & ~w10154;
assign w10157 = ~w10155 & ~w10156;
assign w10158 = b_45 & w657;
assign w10159 = w754 & w29429;
assign w10160 = b_44 & w652;
assign w10161 = ~w10159 & ~w10160;
assign w10162 = ~w10158 & w10161;
assign w10163 = (w10162 & ~w6682) | (w10162 & w25431) | (~w6682 & w25431);
assign w10164 = (w6682 & w25609) | (w6682 & w25610) | (w25609 & w25610);
assign w10165 = (~w6682 & w25839) | (~w6682 & w25840) | (w25839 & w25840);
assign w10166 = ~w10163 & ~w10164;
assign w10167 = ~w10165 & ~w10166;
assign w10168 = (~w10053 & w10057) | (~w10053 & w27751) | (w10057 & w27751);
assign w10169 = (~w10017 & w10021) | (~w10017 & w25107) | (w10021 & w25107);
assign w10170 = ~w10012 & ~w10014;
assign w10171 = (~w10006 & ~w10007) | (~w10006 & w27175) | (~w10007 & w27175);
assign w10172 = b_30 & w2639;
assign w10173 = w2820 & w29430;
assign w10174 = b_29 & w2634;
assign w10175 = ~w10173 & ~w10174;
assign w10176 = ~w10172 & w10175;
assign w10177 = (w10176 & ~w3138) | (w10176 & w29431) | (~w3138 & w29431);
assign w10178 = (w3138 & w39838) | (w3138 & w39839) | (w39838 & w39839);
assign w10179 = (~w3138 & w39840) | (~w3138 & w39841) | (w39840 & w39841);
assign w10180 = ~w10177 & ~w10178;
assign w10181 = ~w10179 & ~w10180;
assign w10182 = (~w9955 & w9958) | (~w9955 & w27176) | (w9958 & w27176);
assign w10183 = b_21 & w4499;
assign w10184 = w4723 & w29432;
assign w10185 = b_20 & w4494;
assign w10186 = ~w10184 & ~w10185;
assign w10187 = ~w10183 & w10186;
assign w10188 = (w10187 & ~w1634) | (w10187 & w29433) | (~w1634 & w29433);
assign w10189 = (w1634 & w39842) | (w1634 & w39843) | (w39842 & w39843);
assign w10190 = (~w1634 & w39844) | (~w1634 & w39845) | (w39844 & w39845);
assign w10191 = ~w10188 & ~w10189;
assign w10192 = ~w10190 & ~w10191;
assign w10193 = (~w9937 & w9840) | (~w9937 & w27064) | (w9840 & w27064);
assign w10194 = b_18 & w5196;
assign w10195 = w5459 & w29434;
assign w10196 = b_17 & w5191;
assign w10197 = ~w10195 & ~w10196;
assign w10198 = ~w10194 & w10197;
assign w10199 = (w10198 & ~w1238) | (w10198 & w25841) | (~w1238 & w25841);
assign w10200 = (w1238 & w29435) | (w1238 & w29436) | (w29435 & w29436);
assign w10201 = (~w1238 & w29437) | (~w1238 & w29438) | (w29437 & w29438);
assign w10202 = ~w10199 & ~w10200;
assign w10203 = ~w10201 & ~w10202;
assign w10204 = (~w9930 & w9851) | (~w9930 & w25842) | (w9851 & w25842);
assign w10205 = b_15 & w5962;
assign w10206 = w6246 & w29439;
assign w10207 = b_14 & w5957;
assign w10208 = ~w10206 & ~w10207;
assign w10209 = ~w10205 & w10208;
assign w10210 = (w10209 & ~w827) | (w10209 & w29440) | (~w827 & w29440);
assign w10211 = (w827 & w39846) | (w827 & w39847) | (w39846 & w39847);
assign w10212 = (~w827 & w39848) | (~w827 & w39849) | (w39848 & w39849);
assign w10213 = ~w10210 & ~w10211;
assign w10214 = ~w10212 & ~w10213;
assign w10215 = (~w9925 & w9862) | (~w9925 & w25843) | (w9862 & w25843);
assign w10216 = b_12 & w6761;
assign w10217 = w7075 & w29441;
assign w10218 = b_11 & w6756;
assign w10219 = ~w10217 & ~w10218;
assign w10220 = ~w10216 & w10219;
assign w10221 = (w10220 & ~w552) | (w10220 & w29442) | (~w552 & w29442);
assign w10222 = (w552 & w39850) | (w552 & w39851) | (w39850 & w39851);
assign w10223 = (~w552 & w39852) | (~w552 & w39853) | (w39852 & w39853);
assign w10224 = ~w10221 & ~w10222;
assign w10225 = ~w10223 & ~w10224;
assign w10226 = ~w9919 & ~w9921;
assign w10227 = b_6 & w8526;
assign w10228 = w8886 & w29443;
assign w10229 = b_5 & w8521;
assign w10230 = ~w10228 & ~w10229;
assign w10231 = ~w10227 & w10230;
assign w10232 = (w10231 & ~w190) | (w10231 & w29444) | (~w190 & w29444);
assign w10233 = (w190 & w39854) | (w190 & w39855) | (w39854 & w39855);
assign w10234 = (~w190 & w39856) | (~w190 & w39857) | (w39856 & w39857);
assign w10235 = ~w10232 & ~w10233;
assign w10236 = ~w10234 & ~w10235;
assign w10237 = a_56 & ~a_57;
assign w10238 = ~a_56 & a_57;
assign w10239 = ~w10237 & ~w10238;
assign w10240 = b_0 & ~w10239;
assign w10241 = (w10240 & w9886) | (w10240 & w26176) | (w9886 & w26176);
assign w10242 = ~w9886 & w26177;
assign w10243 = ~w10241 & ~w10242;
assign w10244 = b_3 & w9534;
assign w10245 = w9876 & w26178;
assign w10246 = b_2 & w9529;
assign w10247 = ~w10245 & ~w10246;
assign w10248 = ~w10244 & w10247;
assign w10249 = w57 & w9537;
assign w10250 = w10248 & ~w10249;
assign w10251 = a_56 & ~w10250;
assign w10252 = w10250 & a_56;
assign w10253 = ~w10250 & ~w10251;
assign w10254 = ~w10252 & ~w10253;
assign w10255 = ~w10243 & ~w10254;
assign w10256 = w10243 & w10254;
assign w10257 = ~w10255 & ~w10256;
assign w10258 = ~w10236 & w10257;
assign w10259 = w10257 & ~w10258;
assign w10260 = ~w10257 & ~w10236;
assign w10261 = ~w10259 & ~w10260;
assign w10262 = ~w9906 & w10261;
assign w10263 = w9906 & ~w10261;
assign w10264 = ~w10262 & ~w10263;
assign w10265 = b_9 & w7613;
assign w10266 = w7941 & w29445;
assign w10267 = b_8 & w7608;
assign w10268 = ~w10266 & ~w10267;
assign w10269 = ~w10265 & w10268;
assign w10270 = (w10269 & ~w371) | (w10269 & w29446) | (~w371 & w29446);
assign w10271 = (w371 & w39858) | (w371 & w39859) | (w39858 & w39859);
assign w10272 = (~w371 & w39860) | (~w371 & w39861) | (w39860 & w39861);
assign w10273 = ~w10270 & ~w10271;
assign w10274 = ~w10272 & ~w10273;
assign w10275 = ~w10264 & ~w10274;
assign w10276 = w10264 & w10274;
assign w10277 = ~w10275 & ~w10276;
assign w10278 = ~w10226 & w10277;
assign w10279 = w10226 & ~w10277;
assign w10280 = ~w10278 & ~w10279;
assign w10281 = w10225 & ~w10280;
assign w10282 = ~w10225 & w10280;
assign w10283 = ~w10281 & ~w10282;
assign w10284 = ~w10215 & w10283;
assign w10285 = w10215 & ~w10283;
assign w10286 = ~w10284 & ~w10285;
assign w10287 = ~w10214 & w10286;
assign w10288 = w10214 & ~w10286;
assign w10289 = ~w10287 & ~w10288;
assign w10290 = (~w25842 & w27065) | (~w25842 & w27066) | (w27065 & w27066);
assign w10291 = (w25842 & w27067) | (w25842 & w27068) | (w27067 & w27068);
assign w10292 = ~w10290 & ~w10291;
assign w10293 = ~w10203 & w10292;
assign w10294 = ~w10292 & ~w10203;
assign w10295 = w10292 & ~w10293;
assign w10296 = ~w10294 & ~w10295;
assign w10297 = ~w10193 & ~w10296;
assign w10298 = w10193 & w10296;
assign w10299 = ~w10297 & ~w10298;
assign w10300 = ~w10192 & w10299;
assign w10301 = w10192 & ~w10299;
assign w10302 = ~w10300 & ~w10301;
assign w10303 = ~w10182 & w10302;
assign w10304 = w10182 & ~w10302;
assign w10305 = ~w10303 & ~w10304;
assign w10306 = b_24 & w3803;
assign w10307 = w4027 & w29447;
assign w10308 = b_23 & w3798;
assign w10309 = ~w10307 & ~w10308;
assign w10310 = ~w10306 & w10309;
assign w10311 = (w10310 & ~w2083) | (w10310 & w29448) | (~w2083 & w29448);
assign w10312 = (w2083 & w39862) | (w2083 & w39863) | (w39862 & w39863);
assign w10313 = (~w2083 & w39864) | (~w2083 & w39865) | (w39864 & w39865);
assign w10314 = ~w10311 & ~w10312;
assign w10315 = ~w10313 & ~w10314;
assign w10316 = w10305 & ~w10315;
assign w10317 = w10305 & ~w10316;
assign w10318 = ~w10305 & ~w10315;
assign w10319 = ~w10317 & ~w10318;
assign w10320 = (~w25827 & w27177) | (~w25827 & w27178) | (w27177 & w27178);
assign w10321 = w10319 & w10320;
assign w10322 = ~w10319 & ~w10320;
assign w10323 = ~w10321 & ~w10322;
assign w10324 = b_27 & w3195;
assign w10325 = w3388 & w29449;
assign w10326 = b_26 & w3190;
assign w10327 = ~w10325 & ~w10326;
assign w10328 = ~w10324 & w10327;
assign w10329 = (w10328 & ~w2582) | (w10328 & w29450) | (~w2582 & w29450);
assign w10330 = (w2582 & w39866) | (w2582 & w39867) | (w39866 & w39867);
assign w10331 = (~w2582 & w39868) | (~w2582 & w39869) | (w39868 & w39869);
assign w10332 = ~w10329 & ~w10330;
assign w10333 = ~w10331 & ~w10332;
assign w10334 = ~w10323 & w10333;
assign w10335 = w10323 & ~w10333;
assign w10336 = ~w10334 & ~w10335;
assign w10337 = ~w9992 & w10336;
assign w10338 = w9992 & ~w10336;
assign w10339 = ~w10337 & ~w10338;
assign w10340 = ~w10181 & w10339;
assign w10341 = w10181 & ~w10339;
assign w10342 = ~w10340 & ~w10341;
assign w10343 = (~w27175 & w27541) | (~w27175 & w27542) | (w27541 & w27542);
assign w10344 = (w27175 & w27543) | (w27175 & w27544) | (w27543 & w27544);
assign w10345 = ~w10343 & ~w10344;
assign w10346 = b_33 & w2158;
assign w10347 = w2294 & w29451;
assign w10348 = b_32 & w2153;
assign w10349 = ~w10347 & ~w10348;
assign w10350 = ~w10346 & w10349;
assign w10351 = (w10350 & ~w3744) | (w10350 & w25611) | (~w3744 & w25611);
assign w10352 = (w3744 & w25844) | (w3744 & w25845) | (w25844 & w25845);
assign w10353 = (~w3744 & w29452) | (~w3744 & w29453) | (w29452 & w29453);
assign w10354 = ~w10351 & ~w10352;
assign w10355 = ~w10353 & ~w10354;
assign w10356 = w10345 & ~w10355;
assign w10357 = w10345 & ~w10356;
assign w10358 = ~w10345 & ~w10355;
assign w10359 = ~w10357 & ~w10358;
assign w10360 = ~w10170 & w10359;
assign w10361 = w10170 & ~w10359;
assign w10362 = ~w10360 & ~w10361;
assign w10363 = b_36 & w1694;
assign w10364 = w1834 & w29454;
assign w10365 = b_35 & w1689;
assign w10366 = ~w10364 & ~w10365;
assign w10367 = ~w10363 & w10366;
assign w10368 = (w10367 & ~w4395) | (w10367 & w25846) | (~w4395 & w25846);
assign w10369 = (w4395 & w29455) | (w4395 & w29456) | (w29455 & w29456);
assign w10370 = (~w4395 & w29457) | (~w4395 & w29458) | (w29457 & w29458);
assign w10371 = ~w10368 & ~w10369;
assign w10372 = ~w10370 & ~w10371;
assign w10373 = ~w10362 & ~w10372;
assign w10374 = w10362 & w10372;
assign w10375 = ~w10373 & ~w10374;
assign w10376 = w10169 & ~w10375;
assign w10377 = ~w10169 & w10375;
assign w10378 = ~w10376 & ~w10377;
assign w10379 = b_39 & w1295;
assign w10380 = w1422 & w29459;
assign w10381 = b_38 & w1290;
assign w10382 = ~w10380 & ~w10381;
assign w10383 = ~w10379 & w10382;
assign w10384 = (w10383 & ~w4888) | (w10383 & w25432) | (~w4888 & w25432);
assign w10385 = (w4888 & w25612) | (w4888 & w25613) | (w25612 & w25613);
assign w10386 = (~w4888 & w25847) | (~w4888 & w25848) | (w25847 & w25848);
assign w10387 = ~w10384 & ~w10385;
assign w10388 = ~w10386 & ~w10387;
assign w10389 = w10378 & ~w10388;
assign w10390 = w10388 & w10378;
assign w10391 = ~w10378 & ~w10388;
assign w10392 = ~w10390 & ~w10391;
assign w10393 = (~w10035 & w10039) | (~w10035 & w27069) | (w10039 & w27069);
assign w10394 = w10392 & w10393;
assign w10395 = ~w10392 & ~w10393;
assign w10396 = ~w10394 & ~w10395;
assign w10397 = b_42 & w986;
assign w10398 = w1069 & w29460;
assign w10399 = b_41 & w981;
assign w10400 = ~w10398 & ~w10399;
assign w10401 = ~w10397 & w10400;
assign w10402 = (w10401 & ~w5864) | (w10401 & w25614) | (~w5864 & w25614);
assign w10403 = (w5864 & w25849) | (w5864 & w25850) | (w25849 & w25850);
assign w10404 = (~w5864 & w26635) | (~w5864 & w26636) | (w26635 & w26636);
assign w10405 = ~w10402 & ~w10403;
assign w10406 = ~w10404 & ~w10405;
assign w10407 = ~w10396 & w10406;
assign w10408 = w10396 & ~w10406;
assign w10409 = ~w10407 & ~w10408;
assign w10410 = ~w10168 & w10409;
assign w10411 = w10168 & ~w10409;
assign w10412 = ~w10410 & ~w10411;
assign w10413 = (w10412 & w10166) | (w10412 & w26822) | (w10166 & w26822);
assign w10414 = (~w26822 & w27427) | (~w26822 & w27428) | (w27427 & w27428);
assign w10415 = w10167 & w10412;
assign w10416 = ~w10414 & ~w10415;
assign w10417 = ~w10075 & ~w10416;
assign w10418 = w10075 & w10416;
assign w10419 = ~w10417 & ~w10418;
assign w10420 = ~w10157 & w10419;
assign w10421 = ~w10419 & ~w10157;
assign w10422 = w10157 & w10419;
assign w10423 = ~w10421 & ~w10422;
assign w10424 = ~w10147 & ~w10423;
assign w10425 = w10147 & w10423;
assign w10426 = ~w10424 & ~w10425;
assign w10427 = ~w10146 & w10426;
assign w10428 = ~w10426 & ~w10146;
assign w10429 = w10426 & ~w10427;
assign w10430 = ~w10428 & ~w10429;
assign w10431 = ~w10136 & ~w10430;
assign w10432 = w10136 & w10430;
assign w10433 = ~w10431 & ~w10432;
assign w10434 = ~w10135 & w10433;
assign w10435 = ~w10433 & ~w10135;
assign w10436 = w10433 & ~w10434;
assign w10437 = ~w10435 & ~w10436;
assign w10438 = ~w10125 & ~w10437;
assign w10439 = ~w10125 & ~w10438;
assign w10440 = w10125 & ~w10437;
assign w10441 = ~w10439 & ~w10440;
assign w10442 = w8 & w29461;
assign w10443 = ~w8 & w29462;
assign w10444 = b_56 & w4;
assign w10445 = ~w10443 & ~w10444;
assign w10446 = ~w10442 & w10445;
assign w10447 = ~b_56 & ~b_57;
assign w10448 = b_56 & b_57;
assign w10449 = ~w10447 & ~w10448;
assign w10450 = (w6406 & w39870) | (w6406 & w39871) | (w39870 & w39871);
assign w10451 = (~w6406 & w39872) | (~w6406 & w39873) | (w39872 & w39873);
assign w10452 = ~w10450 & ~w10451;
assign w10453 = (w10446 & ~w10452) | (w10446 & w29469) | (~w10452 & w29469);
assign w10454 = (w10452 & w39874) | (w10452 & w39875) | (w39874 & w39875);
assign w10455 = (~w10452 & w39876) | (~w10452 & w39877) | (w39876 & w39877);
assign w10456 = ~w10453 & ~w10454;
assign w10457 = ~w10455 & ~w10456;
assign w10458 = (~w10457 & w10439) | (~w10457 & w25853) | (w10439 & w25853);
assign w10459 = ~w10441 & ~w10458;
assign w10460 = ~w10439 & w39878;
assign w10461 = ~w10459 & ~w10460;
assign w10462 = (~w10117 & w10121) | (~w10117 & w25108) | (w10121 & w25108);
assign w10463 = ~w10461 & ~w10462;
assign w10464 = w10461 & w10462;
assign w10465 = ~w10463 & ~w10464;
assign w10466 = w8 & w29470;
assign w10467 = ~w8 & w29471;
assign w10468 = b_57 & w4;
assign w10469 = ~w10467 & ~w10468;
assign w10470 = ~w10466 & w10469;
assign w10471 = ~b_57 & ~b_58;
assign w10472 = b_57 & b_58;
assign w10473 = ~w10471 & ~w10472;
assign w10474 = (w6406 & w39879) | (w6406 & w39880) | (w39879 & w39880);
assign w10475 = (~w6406 & w39881) | (~w6406 & w39882) | (w39881 & w39882);
assign w10476 = ~w10474 & ~w10475;
assign w10477 = (w10470 & ~w10476) | (w10470 & w29478) | (~w10476 & w29478);
assign w10478 = (w10476 & w39883) | (w10476 & w39884) | (w39883 & w39884);
assign w10479 = (~w10476 & w39885) | (~w10476 & w39886) | (w39885 & w39886);
assign w10480 = ~w10477 & ~w10478;
assign w10481 = ~w10479 & ~w10480;
assign w10482 = b_55 & w99;
assign w10483 = w136 & w29479;
assign w10484 = b_54 & w94;
assign w10485 = ~w10483 & ~w10484;
assign w10486 = ~w10482 & w10485;
assign w10487 = (w10486 & ~w9776) | (w10486 & w29480) | (~w9776 & w29480);
assign w10488 = (w9776 & w39887) | (w9776 & w39888) | (w39887 & w39888);
assign w10489 = (~w9776 & w39889) | (~w9776 & w39890) | (w39889 & w39890);
assign w10490 = ~w10487 & ~w10488;
assign w10491 = ~w10489 & ~w10490;
assign w10492 = b_52 & w239;
assign w10493 = w266 & w29481;
assign w10494 = b_51 & w234;
assign w10495 = ~w10493 & ~w10494;
assign w10496 = ~w10492 & w10495;
assign w10497 = (w10496 & ~w8793) | (w10496 & w25855) | (~w8793 & w25855);
assign w10498 = (w8793 & w29482) | (w8793 & w29483) | (w29482 & w29483);
assign w10499 = (~w8793 & w29484) | (~w8793 & w29485) | (w29484 & w29485);
assign w10500 = ~w10497 & ~w10498;
assign w10501 = ~w10499 & ~w10500;
assign w10502 = (~w10420 & w10147) | (~w10420 & w27429) | (w10147 & w27429);
assign w10503 = b_49 & w418;
assign w10504 = w481 & w29486;
assign w10505 = b_48 & w413;
assign w10506 = ~w10504 & ~w10505;
assign w10507 = ~w10503 & w10506;
assign w10508 = (w10507 & ~w7859) | (w10507 & w25615) | (~w7859 & w25615);
assign w10509 = (w7859 & w25856) | (w7859 & w25857) | (w25856 & w25857);
assign w10510 = (~w7859 & w29487) | (~w7859 & w29488) | (w29487 & w29488);
assign w10511 = ~w10508 & ~w10509;
assign w10512 = ~w10510 & ~w10511;
assign w10513 = (~w10413 & w10416) | (~w10413 & w25858) | (w10416 & w25858);
assign w10514 = (~w10408 & w10168) | (~w10408 & w27830) | (w10168 & w27830);
assign w10515 = (~w10340 & w10171) | (~w10340 & w27238) | (w10171 & w27238);
assign w10516 = (~w10335 & w9992) | (~w10335 & w27239) | (w9992 & w27239);
assign w10517 = (~w10293 & w10193) | (~w10293 & w25859) | (w10193 & w25859);
assign w10518 = ~w10282 & ~w10284;
assign w10519 = b_10 & w7613;
assign w10520 = w7941 & w29489;
assign w10521 = b_9 & w7608;
assign w10522 = ~w10520 & ~w10521;
assign w10523 = ~w10519 & w10522;
assign w10524 = (w10523 & ~w454) | (w10523 & w29490) | (~w454 & w29490);
assign w10525 = (w454 & w39891) | (w454 & w39892) | (w39891 & w39892);
assign w10526 = (~w454 & w39893) | (~w454 & w39894) | (w39893 & w39894);
assign w10527 = ~w10524 & ~w10525;
assign w10528 = ~w10526 & ~w10527;
assign w10529 = ~w9906 & ~w10261;
assign w10530 = b_7 & w8526;
assign w10531 = w8886 & w29491;
assign w10532 = b_6 & w8521;
assign w10533 = ~w10531 & ~w10532;
assign w10534 = ~w10530 & w10533;
assign w10535 = (w10534 & ~w213) | (w10534 & w29492) | (~w213 & w29492);
assign w10536 = (w213 & w39895) | (w213 & w39896) | (w39895 & w39896);
assign w10537 = (~w213 & w39897) | (~w213 & w39898) | (w39897 & w39898);
assign w10538 = ~w10535 & ~w10536;
assign w10539 = ~w10537 & ~w10538;
assign w10540 = ~w9886 & w26179;
assign w10541 = (~w10540 & w10243) | (~w10540 & w25860) | (w10243 & w25860);
assign w10542 = b_4 & w9534;
assign w10543 = w9876 & w26180;
assign w10544 = b_3 & w9529;
assign w10545 = ~w10543 & ~w10544;
assign w10546 = ~w10542 & w10545;
assign w10547 = w84 & w9537;
assign w10548 = w10546 & ~w10547;
assign w10549 = (a_56 & w10547) | (a_56 & w26181) | (w10547 & w26181);
assign w10550 = ~w10547 & w27354;
assign w10551 = ~w10548 & ~w10549;
assign w10552 = ~w10550 & ~w10551;
assign w10553 = (a_59 & w10239) | (a_59 & w29493) | (w10239 & w29493);
assign w10554 = ~a_57 & a_58;
assign w10555 = a_57 & ~a_58;
assign w10556 = ~w10554 & ~w10555;
assign w10557 = w10239 & ~w10556;
assign w10558 = b_0 & w10557;
assign w10559 = ~a_58 & a_59;
assign w10560 = a_58 & ~a_59;
assign w10561 = ~w10559 & ~w10560;
assign w10562 = ~w10239 & w10561;
assign w10563 = b_1 & w10562;
assign w10564 = ~w10558 & ~w10563;
assign w10565 = ~w10239 & ~w10561;
assign w10566 = ~w15 & w10565;
assign w10567 = w10564 & ~w10566;
assign w10568 = (a_59 & ~w10564) | (a_59 & w26182) | (~w10564 & w26182);
assign w10569 = w10564 & w27355;
assign w10570 = ~w10567 & ~w10568;
assign w10571 = (w10553 & w10570) | (w10553 & w27356) | (w10570 & w27356);
assign w10572 = ~w10570 & w27357;
assign w10573 = ~w10571 & ~w10572;
assign w10574 = w10552 & ~w10573;
assign w10575 = ~w10552 & w10573;
assign w10576 = ~w10574 & ~w10575;
assign w10577 = ~w10541 & w10576;
assign w10578 = w10541 & ~w10576;
assign w10579 = ~w10577 & ~w10578;
assign w10580 = w10539 & ~w10579;
assign w10581 = ~w10539 & w10579;
assign w10582 = ~w10580 & ~w10581;
assign w10583 = (w10582 & w10529) | (w10582 & w26183) | (w10529 & w26183);
assign w10584 = ~w10529 & w26184;
assign w10585 = ~w10583 & ~w10584;
assign w10586 = ~w10528 & w10585;
assign w10587 = w10528 & w10585;
assign w10588 = ~w10585 & ~w10528;
assign w10589 = ~w10587 & ~w10588;
assign w10590 = (~w10275 & w10226) | (~w10275 & w26185) | (w10226 & w26185);
assign w10591 = w10589 & w10590;
assign w10592 = ~w10589 & ~w10590;
assign w10593 = ~w10591 & ~w10592;
assign w10594 = b_13 & w6761;
assign w10595 = w7075 & w29494;
assign w10596 = b_12 & w6756;
assign w10597 = ~w10595 & ~w10596;
assign w10598 = ~w10594 & w10597;
assign w10599 = (w10598 & ~w711) | (w10598 & w29495) | (~w711 & w29495);
assign w10600 = (w711 & w39899) | (w711 & w39900) | (w39899 & w39900);
assign w10601 = (~w711 & w39901) | (~w711 & w39902) | (w39901 & w39902);
assign w10602 = ~w10599 & ~w10600;
assign w10603 = ~w10601 & ~w10602;
assign w10604 = w10593 & ~w10603;
assign w10605 = ~w10593 & w10603;
assign w10606 = ~w10518 & w26186;
assign w10607 = ~w10518 & ~w10606;
assign w10608 = ~w10604 & ~w10606;
assign w10609 = ~w10606 & w26186;
assign w10610 = ~w10607 & ~w10609;
assign w10611 = b_16 & w5962;
assign w10612 = w6246 & w29496;
assign w10613 = b_15 & w5957;
assign w10614 = ~w10612 & ~w10613;
assign w10615 = ~w10611 & w10614;
assign w10616 = (w10615 & ~w926) | (w10615 & w29497) | (~w926 & w29497);
assign w10617 = (w926 & w39903) | (w926 & w39904) | (w39903 & w39904);
assign w10618 = (~w926 & w39905) | (~w926 & w39906) | (w39905 & w39906);
assign w10619 = ~w10616 & ~w10617;
assign w10620 = ~w10618 & ~w10619;
assign w10621 = ~w10610 & ~w10620;
assign w10622 = ~w10610 & ~w10621;
assign w10623 = w10610 & ~w10620;
assign w10624 = ~w10622 & ~w10623;
assign w10625 = (~w10287 & w10204) | (~w10287 & w26187) | (w10204 & w26187);
assign w10626 = ~w10622 & w27358;
assign w10627 = (~w10625 & w10622) | (~w10625 & w27359) | (w10622 & w27359);
assign w10628 = ~w10626 & ~w10627;
assign w10629 = b_19 & w5196;
assign w10630 = w5459 & w29498;
assign w10631 = b_18 & w5191;
assign w10632 = ~w10630 & ~w10631;
assign w10633 = ~w10629 & w10632;
assign w10634 = (w10633 & ~w1372) | (w10633 & w29499) | (~w1372 & w29499);
assign w10635 = (w1372 & w39907) | (w1372 & w39908) | (w39907 & w39908);
assign w10636 = (~w1372 & w39909) | (~w1372 & w39910) | (w39909 & w39910);
assign w10637 = ~w10634 & ~w10635;
assign w10638 = ~w10636 & ~w10637;
assign w10639 = w10628 & ~w10638;
assign w10640 = ~w10628 & w10638;
assign w10641 = ~w10517 & w26188;
assign w10642 = ~w10517 & ~w10641;
assign w10643 = ~w10639 & ~w10641;
assign w10644 = ~w10641 & w26188;
assign w10645 = ~w10642 & ~w10644;
assign w10646 = b_22 & w4499;
assign w10647 = w4723 & w29500;
assign w10648 = b_21 & w4494;
assign w10649 = ~w10647 & ~w10648;
assign w10650 = ~w10646 & w10649;
assign w10651 = (w10650 & ~w1786) | (w10650 & w29501) | (~w1786 & w29501);
assign w10652 = (w1786 & w39911) | (w1786 & w39912) | (w39911 & w39912);
assign w10653 = (~w1786 & w39913) | (~w1786 & w39914) | (w39913 & w39914);
assign w10654 = ~w10651 & ~w10652;
assign w10655 = ~w10653 & ~w10654;
assign w10656 = ~w10645 & ~w10655;
assign w10657 = ~w10645 & ~w10656;
assign w10658 = w10645 & ~w10655;
assign w10659 = ~w10657 & ~w10658;
assign w10660 = (~w10300 & w10182) | (~w10300 & w27240) | (w10182 & w27240);
assign w10661 = w10659 & w10660;
assign w10662 = ~w10659 & ~w10660;
assign w10663 = ~w10661 & ~w10662;
assign w10664 = b_25 & w3803;
assign w10665 = w4027 & w29502;
assign w10666 = b_24 & w3798;
assign w10667 = ~w10665 & ~w10666;
assign w10668 = ~w10664 & w10667;
assign w10669 = (w10668 & ~w2108) | (w10668 & w26189) | (~w2108 & w26189);
assign w10670 = (w2108 & w29503) | (w2108 & w29504) | (w29503 & w29504);
assign w10671 = (~w2108 & w29505) | (~w2108 & w29506) | (w29505 & w29506);
assign w10672 = ~w10669 & ~w10670;
assign w10673 = ~w10671 & ~w10672;
assign w10674 = w10663 & ~w10673;
assign w10675 = w10663 & ~w10674;
assign w10676 = ~w10663 & ~w10673;
assign w10677 = ~w10675 & ~w10676;
assign w10678 = ~w10316 & ~w10322;
assign w10679 = w10677 & w10678;
assign w10680 = ~w10677 & ~w10678;
assign w10681 = ~w10679 & ~w10680;
assign w10682 = b_28 & w3195;
assign w10683 = w3388 & w29507;
assign w10684 = b_27 & w3190;
assign w10685 = ~w10683 & ~w10684;
assign w10686 = ~w10682 & w10685;
assign w10687 = (w10686 & ~w2771) | (w10686 & w25861) | (~w2771 & w25861);
assign w10688 = (w2771 & w26190) | (w2771 & w26191) | (w26190 & w26191);
assign w10689 = (~w2771 & w29508) | (~w2771 & w29509) | (w29508 & w29509);
assign w10690 = ~w10687 & ~w10688;
assign w10691 = ~w10689 & ~w10690;
assign w10692 = w10681 & ~w10691;
assign w10693 = w10681 & ~w10692;
assign w10694 = ~w10681 & ~w10691;
assign w10695 = ~w10693 & ~w10694;
assign w10696 = ~w10516 & w10695;
assign w10697 = w10516 & ~w10695;
assign w10698 = ~w10696 & ~w10697;
assign w10699 = b_31 & w2639;
assign w10700 = w2820 & w29510;
assign w10701 = b_30 & w2634;
assign w10702 = ~w10700 & ~w10701;
assign w10703 = ~w10699 & w10702;
assign w10704 = (w10703 & ~w3345) | (w10703 & w26192) | (~w3345 & w26192);
assign w10705 = (w3345 & w29511) | (w3345 & w29512) | (w29511 & w29512);
assign w10706 = (~w3345 & w29513) | (~w3345 & w29514) | (w29513 & w29514);
assign w10707 = ~w10704 & ~w10705;
assign w10708 = ~w10706 & ~w10707;
assign w10709 = ~w10698 & ~w10708;
assign w10710 = w10698 & w10708;
assign w10711 = ~w10709 & ~w10710;
assign w10712 = w10515 & ~w10711;
assign w10713 = ~w10515 & w10711;
assign w10714 = ~w10712 & ~w10713;
assign w10715 = b_34 & w2158;
assign w10716 = w2294 & w29515;
assign w10717 = b_33 & w2153;
assign w10718 = ~w10716 & ~w10717;
assign w10719 = ~w10715 & w10718;
assign w10720 = (w10719 & ~w3967) | (w10719 & w25862) | (~w3967 & w25862);
assign w10721 = (w3967 & w26193) | (w3967 & w26194) | (w26193 & w26194);
assign w10722 = (~w3967 & w29516) | (~w3967 & w29517) | (w29516 & w29517);
assign w10723 = ~w10720 & ~w10721;
assign w10724 = ~w10722 & ~w10723;
assign w10725 = w10714 & ~w10724;
assign w10726 = w10714 & ~w10725;
assign w10727 = ~w10714 & ~w10724;
assign w10728 = ~w10726 & ~w10727;
assign w10729 = (~w10356 & w10170) | (~w10356 & w25863) | (w10170 & w25863);
assign w10730 = w10728 & w10729;
assign w10731 = ~w10728 & ~w10729;
assign w10732 = ~w10730 & ~w10731;
assign w10733 = b_37 & w1694;
assign w10734 = w1834 & w29518;
assign w10735 = b_36 & w1689;
assign w10736 = ~w10734 & ~w10735;
assign w10737 = ~w10733 & w10736;
assign w10738 = (w10737 & ~w4636) | (w10737 & w25616) | (~w4636 & w25616);
assign w10739 = (w4636 & w25864) | (w4636 & w25865) | (w25864 & w25865);
assign w10740 = (~w4636 & w29519) | (~w4636 & w29520) | (w29519 & w29520);
assign w10741 = ~w10738 & ~w10739;
assign w10742 = ~w10740 & ~w10741;
assign w10743 = w10732 & ~w10742;
assign w10744 = w10732 & ~w10743;
assign w10745 = ~w10732 & ~w10742;
assign w10746 = ~w10744 & ~w10745;
assign w10747 = (~w10373 & w10169) | (~w10373 & w25866) | (w10169 & w25866);
assign w10748 = w10746 & w10747;
assign w10749 = ~w10746 & ~w10747;
assign w10750 = ~w10748 & ~w10749;
assign w10751 = b_40 & w1295;
assign w10752 = w1422 & w29521;
assign w10753 = b_39 & w1290;
assign w10754 = ~w10752 & ~w10753;
assign w10755 = ~w10751 & w10754;
assign w10756 = (w10755 & ~w5363) | (w10755 & w25433) | (~w5363 & w25433);
assign w10757 = (w5363 & w25617) | (w5363 & w25618) | (w25617 & w25618);
assign w10758 = (~w5363 & w25867) | (~w5363 & w25868) | (w25867 & w25868);
assign w10759 = ~w10756 & ~w10757;
assign w10760 = ~w10758 & ~w10759;
assign w10761 = w10750 & ~w10760;
assign w10762 = w10760 & w10750;
assign w10763 = ~w10750 & ~w10760;
assign w10764 = ~w10762 & ~w10763;
assign w10765 = (~w10389 & w10393) | (~w10389 & w25109) | (w10393 & w25109);
assign w10766 = w10764 & w10765;
assign w10767 = ~w10764 & ~w10765;
assign w10768 = ~w10766 & ~w10767;
assign w10769 = b_43 & w986;
assign w10770 = w1069 & w29522;
assign w10771 = b_42 & w981;
assign w10772 = ~w10770 & ~w10771;
assign w10773 = ~w10769 & w10772;
assign w10774 = (w10773 & ~w5888) | (w10773 & w25619) | (~w5888 & w25619);
assign w10775 = (w5888 & w25869) | (w5888 & w25870) | (w25869 & w25870);
assign w10776 = (~w5888 & w26195) | (~w5888 & w26196) | (w26195 & w26196);
assign w10777 = ~w10774 & ~w10775;
assign w10778 = ~w10776 & ~w10777;
assign w10779 = w10768 & ~w10778;
assign w10780 = ~w10768 & w10778;
assign w10781 = (w10410 & w25871) | (w10410 & w25872) | (w25871 & w25872);
assign w10782 = ~w10514 & ~w10781;
assign w10783 = (~w25871 & w27241) | (~w25871 & w27242) | (w27241 & w27242);
assign w10784 = ~w10781 & w25872;
assign w10785 = ~w10782 & ~w10784;
assign w10786 = b_46 & w657;
assign w10787 = w754 & w29523;
assign w10788 = b_45 & w652;
assign w10789 = ~w10787 & ~w10788;
assign w10790 = ~w10786 & w10789;
assign w10791 = (w10790 & ~w6974) | (w10790 & w25620) | (~w6974 & w25620);
assign w10792 = (w6974 & w25873) | (w6974 & w25874) | (w25873 & w25874);
assign w10793 = (~w6974 & w26197) | (~w6974 & w26198) | (w26197 & w26198);
assign w10794 = ~w10791 & ~w10792;
assign w10795 = ~w10793 & ~w10794;
assign w10796 = w10785 & w10795;
assign w10797 = ~w10785 & ~w10795;
assign w10798 = ~w10796 & ~w10797;
assign w10799 = ~w10513 & w10798;
assign w10800 = w10513 & ~w10798;
assign w10801 = ~w10799 & ~w10800;
assign w10802 = w10512 & ~w10801;
assign w10803 = ~w10512 & w10801;
assign w10804 = ~w10802 & ~w10803;
assign w10805 = (w10804 & w10424) | (w10804 & w26637) | (w10424 & w26637);
assign w10806 = ~w10424 & w26638;
assign w10807 = ~w10805 & ~w10806;
assign w10808 = w10501 & ~w10807;
assign w10809 = ~w10501 & w10807;
assign w10810 = ~w10808 & ~w10809;
assign w10811 = (w10810 & w10431) | (w10810 & w25111) | (w10431 & w25111);
assign w10812 = ~w10431 & w29524;
assign w10813 = ~w10811 & ~w10812;
assign w10814 = w10491 & ~w10813;
assign w10815 = ~w10491 & w10813;
assign w10816 = ~w10814 & ~w10815;
assign w10817 = (~w25854 & w29525) | (~w25854 & w29526) | (w29525 & w29526);
assign w10818 = (w25854 & w29527) | (w25854 & w29528) | (w29527 & w29528);
assign w10819 = ~w10817 & ~w10818;
assign w10820 = ~w10481 & w10819;
assign w10821 = w10819 & ~w10820;
assign w10822 = ~w10819 & ~w10481;
assign w10823 = ~w10821 & ~w10822;
assign w10824 = (~w10458 & w10461) | (~w10458 & w39915) | (w10461 & w39915);
assign w10825 = ~w10823 & ~w10824;
assign w10826 = w10823 & w10824;
assign w10827 = ~w10825 & ~w10826;
assign w10828 = (~w10820 & w10824) | (~w10820 & w25112) | (w10824 & w25112);
assign w10829 = ~w10815 & ~w10817;
assign w10830 = (~w10431 & w26639) | (~w10431 & w26640) | (w26639 & w26640);
assign w10831 = b_53 & w239;
assign w10832 = w266 & w29529;
assign w10833 = b_52 & w234;
assign w10834 = ~w10832 & ~w10833;
assign w10835 = ~w10831 & w10834;
assign w10836 = (w9109 & w39916) | (w9109 & w39917) | (w39916 & w39917);
assign w10837 = a_8 & ~w10836;
assign w10838 = w10836 & a_8;
assign w10839 = ~w10836 & ~w10837;
assign w10840 = ~w10838 & ~w10839;
assign w10841 = (~w10803 & w10502) | (~w10803 & w25875) | (w10502 & w25875);
assign w10842 = b_50 & w418;
assign w10843 = w481 & w29531;
assign w10844 = b_49 & w413;
assign w10845 = ~w10843 & ~w10844;
assign w10846 = ~w10842 & w10845;
assign w10847 = (w10846 & ~w8162) | (w10846 & w25876) | (~w8162 & w25876);
assign w10848 = (w8162 & w26199) | (w8162 & w26200) | (w26199 & w26200);
assign w10849 = (~w8162 & w29532) | (~w8162 & w29533) | (w29532 & w29533);
assign w10850 = ~w10847 & ~w10848;
assign w10851 = ~w10849 & ~w10850;
assign w10852 = ~w10761 & ~w10767;
assign w10853 = b_35 & w2158;
assign w10854 = w2294 & w29534;
assign w10855 = b_34 & w2153;
assign w10856 = ~w10854 & ~w10855;
assign w10857 = ~w10853 & w10856;
assign w10858 = (w10857 & ~w4181) | (w10857 & w25877) | (~w4181 & w25877);
assign w10859 = (w4181 & w26201) | (w4181 & w26202) | (w26201 & w26202);
assign w10860 = (~w4181 & w29535) | (~w4181 & w29536) | (w29535 & w29536);
assign w10861 = ~w10858 & ~w10859;
assign w10862 = ~w10860 & ~w10861;
assign w10863 = (~w10709 & w10515) | (~w10709 & w26203) | (w10515 & w26203);
assign w10864 = ~w10516 & ~w10695;
assign w10865 = (~w10692 & w10695) | (~w10692 & w27430) | (w10695 & w27430);
assign w10866 = (~w10656 & w10659) | (~w10656 & w27243) | (w10659 & w27243);
assign w10867 = (~w10621 & w10624) | (~w10621 & w25113) | (w10624 & w25113);
assign w10868 = b_17 & w5962;
assign w10869 = w6246 & w29537;
assign w10870 = b_16 & w5957;
assign w10871 = ~w10869 & ~w10870;
assign w10872 = ~w10868 & w10871;
assign w10873 = (w10872 & ~w1038) | (w10872 & w25878) | (~w1038 & w25878);
assign w10874 = (w1038 & w26204) | (w1038 & w26205) | (w26204 & w26205);
assign w10875 = (~w1038 & w29538) | (~w1038 & w29539) | (w29538 & w29539);
assign w10876 = ~w10873 & ~w10874;
assign w10877 = ~w10875 & ~w10876;
assign w10878 = b_14 & w6761;
assign w10879 = w7075 & w29540;
assign w10880 = b_13 & w6756;
assign w10881 = ~w10879 & ~w10880;
assign w10882 = ~w10878 & w10881;
assign w10883 = (w10882 & ~w735) | (w10882 & w26206) | (~w735 & w26206);
assign w10884 = (w735 & w29541) | (w735 & w29542) | (w29541 & w29542);
assign w10885 = (~w735 & w29543) | (~w735 & w29544) | (w29543 & w29544);
assign w10886 = ~w10883 & ~w10884;
assign w10887 = ~w10885 & ~w10886;
assign w10888 = (~w10586 & w10590) | (~w10586 & w26916) | (w10590 & w26916);
assign w10889 = b_11 & w7613;
assign w10890 = w7941 & w29545;
assign w10891 = b_10 & w7608;
assign w10892 = ~w10890 & ~w10891;
assign w10893 = ~w10889 & w10892;
assign w10894 = (w10893 & ~w530) | (w10893 & w29546) | (~w530 & w29546);
assign w10895 = (w530 & w39918) | (w530 & w39919) | (w39918 & w39919);
assign w10896 = (~w530 & w39920) | (~w530 & w39921) | (w39920 & w39921);
assign w10897 = ~w10894 & ~w10895;
assign w10898 = ~w10896 & ~w10897;
assign w10899 = ~w10581 & ~w10583;
assign w10900 = ~w10575 & ~w10577;
assign w10901 = b_2 & w10562;
assign w10902 = w10239 & ~w10561;
assign w10903 = w10902 & w26207;
assign w10904 = b_1 & w10557;
assign w10905 = ~w10903 & ~w10904;
assign w10906 = ~w10901 & w10905;
assign w10907 = w35 & w10565;
assign w10908 = w10906 & ~w10907;
assign w10909 = (a_59 & ~w10906) | (a_59 & w26641) | (~w10906 & w26641);
assign w10910 = w10906 & w27360;
assign w10911 = ~w10908 & ~w10909;
assign w10912 = ~w10910 & ~w10911;
assign w10913 = ~w10571 & w10912;
assign w10914 = w10571 & ~w10912;
assign w10915 = ~w10913 & ~w10914;
assign w10916 = b_5 & w9534;
assign w10917 = w9876 & w26823;
assign w10918 = b_4 & w9529;
assign w10919 = ~w10917 & ~w10918;
assign w10920 = ~w10916 & w10919;
assign w10921 = w129 & w9537;
assign w10922 = w10920 & ~w10921;
assign w10923 = (a_56 & w10921) | (a_56 & w26824) | (w10921 & w26824);
assign w10924 = ~w10921 & w39922;
assign w10925 = ~w10922 & ~w10923;
assign w10926 = ~w10924 & ~w10925;
assign w10927 = w10915 & ~w10926;
assign w10928 = ~w10915 & w10926;
assign w10929 = ~w10900 & w26208;
assign w10930 = ~w10900 & ~w10929;
assign w10931 = (~w10927 & w10900) | (~w10927 & w26642) | (w10900 & w26642);
assign w10932 = ~w10928 & w10931;
assign w10933 = ~w10930 & ~w10932;
assign w10934 = b_8 & w8526;
assign w10935 = w8886 & w29547;
assign w10936 = b_7 & w8521;
assign w10937 = ~w10935 & ~w10936;
assign w10938 = ~w10934 & w10937;
assign w10939 = ~w308 & w29548;
assign w10940 = (w10938 & ~w29548) | (w10938 & w39923) | (~w29548 & w39923);
assign w10941 = (w29548 & w39924) | (w29548 & w39925) | (w39924 & w39925);
assign w10942 = ~w10939 & w29550;
assign w10943 = ~w10940 & ~w10941;
assign w10944 = ~w10942 & ~w10943;
assign w10945 = w10933 & w10944;
assign w10946 = ~w10933 & ~w10944;
assign w10947 = ~w10945 & ~w10946;
assign w10948 = ~w10899 & w10947;
assign w10949 = w10899 & ~w10947;
assign w10950 = ~w10948 & ~w10949;
assign w10951 = w10898 & ~w10950;
assign w10952 = ~w10898 & w10950;
assign w10953 = ~w10951 & ~w10952;
assign w10954 = ~w10888 & w10953;
assign w10955 = w10888 & ~w10953;
assign w10956 = ~w10954 & ~w10955;
assign w10957 = ~w10887 & w10956;
assign w10958 = w10956 & ~w10957;
assign w10959 = ~w10956 & ~w10887;
assign w10960 = ~w10958 & ~w10959;
assign w10961 = ~w10608 & ~w10960;
assign w10962 = w10608 & w10960;
assign w10963 = ~w10961 & ~w10962;
assign w10964 = ~w10877 & w10963;
assign w10965 = ~w10963 & ~w10877;
assign w10966 = w10963 & ~w10964;
assign w10967 = ~w10965 & ~w10966;
assign w10968 = ~w10867 & ~w10967;
assign w10969 = ~w10867 & ~w10968;
assign w10970 = ~w10967 & ~w10968;
assign w10971 = ~w10969 & ~w10970;
assign w10972 = b_20 & w5196;
assign w10973 = w5459 & w29551;
assign w10974 = b_19 & w5191;
assign w10975 = ~w10973 & ~w10974;
assign w10976 = ~w10972 & w10975;
assign w10977 = (w10976 & ~w1503) | (w10976 & w29552) | (~w1503 & w29552);
assign w10978 = (w1503 & w39926) | (w1503 & w39927) | (w39926 & w39927);
assign w10979 = (~w1503 & w39928) | (~w1503 & w39929) | (w39928 & w39929);
assign w10980 = ~w10977 & ~w10978;
assign w10981 = ~w10979 & ~w10980;
assign w10982 = ~w10971 & ~w10981;
assign w10983 = ~w10971 & ~w10982;
assign w10984 = w10971 & ~w10981;
assign w10985 = ~w10983 & ~w10984;
assign w10986 = ~w10983 & w27361;
assign w10987 = (w10643 & w10983) | (w10643 & w27362) | (w10983 & w27362);
assign w10988 = ~w10986 & ~w10987;
assign w10989 = b_23 & w4499;
assign w10990 = w4723 & w29553;
assign w10991 = b_22 & w4494;
assign w10992 = ~w10990 & ~w10991;
assign w10993 = ~w10989 & w10992;
assign w10994 = (w10993 & ~w1933) | (w10993 & w29554) | (~w1933 & w29554);
assign w10995 = (w1933 & w39930) | (w1933 & w39931) | (w39930 & w39931);
assign w10996 = (~w1933 & w39932) | (~w1933 & w39933) | (w39932 & w39933);
assign w10997 = ~w10994 & ~w10995;
assign w10998 = ~w10996 & ~w10997;
assign w10999 = ~w10988 & ~w10998;
assign w11000 = w10988 & w10998;
assign w11001 = ~w10999 & ~w11000;
assign w11002 = w10866 & ~w11001;
assign w11003 = ~w10866 & w11001;
assign w11004 = ~w11002 & ~w11003;
assign w11005 = b_26 & w3803;
assign w11006 = w4027 & w29555;
assign w11007 = b_25 & w3798;
assign w11008 = ~w11006 & ~w11007;
assign w11009 = ~w11005 & w11008;
assign w11010 = (w11009 & ~w2416) | (w11009 & w26209) | (~w2416 & w26209);
assign w11011 = (w2416 & w29556) | (w2416 & w29557) | (w29556 & w29557);
assign w11012 = (~w2416 & w29558) | (~w2416 & w29559) | (w29558 & w29559);
assign w11013 = ~w11010 & ~w11011;
assign w11014 = ~w11012 & ~w11013;
assign w11015 = w11004 & ~w11014;
assign w11016 = w11004 & ~w11015;
assign w11017 = ~w11004 & ~w11014;
assign w11018 = ~w11016 & ~w11017;
assign w11019 = (~w10674 & w10678) | (~w10674 & w26210) | (w10678 & w26210);
assign w11020 = w11018 & w11019;
assign w11021 = ~w11018 & ~w11019;
assign w11022 = ~w11020 & ~w11021;
assign w11023 = b_29 & w3195;
assign w11024 = w3388 & w29560;
assign w11025 = b_28 & w3190;
assign w11026 = ~w11024 & ~w11025;
assign w11027 = ~w11023 & w11026;
assign w11028 = (w11027 & ~w2954) | (w11027 & w25879) | (~w2954 & w25879);
assign w11029 = (w2954 & w26211) | (w2954 & w26212) | (w26211 & w26212);
assign w11030 = (~w2954 & w29561) | (~w2954 & w29562) | (w29561 & w29562);
assign w11031 = ~w11028 & ~w11029;
assign w11032 = ~w11030 & ~w11031;
assign w11033 = w11022 & ~w11032;
assign w11034 = ~w11022 & w11032;
assign w11035 = (w10864 & w26213) | (w10864 & w26214) | (w26213 & w26214);
assign w11036 = ~w10865 & ~w11035;
assign w11037 = (~w10864 & w27545) | (~w10864 & w27546) | (w27545 & w27546);
assign w11038 = ~w10864 & w27431;
assign w11039 = b_32 & w2639;
assign w11040 = w2820 & w29563;
assign w11041 = b_31 & w2634;
assign w11042 = ~w11040 & ~w11041;
assign w11043 = ~w11039 & w11042;
assign w11044 = (w11043 & ~w3545) | (w11043 & w26215) | (~w3545 & w26215);
assign w11045 = (w3545 & w29564) | (w3545 & w29565) | (w29564 & w29565);
assign w11046 = (~w3545 & w29566) | (~w3545 & w29567) | (w29566 & w29567);
assign w11047 = ~w11044 & ~w11045;
assign w11048 = ~w11046 & ~w11047;
assign w11049 = ~w11036 & w27432;
assign w11050 = (~w11048 & w11036) | (~w11048 & w27433) | (w11036 & w27433);
assign w11051 = ~w11049 & ~w11050;
assign w11052 = ~w10863 & w11051;
assign w11053 = w10863 & ~w11051;
assign w11054 = ~w11052 & ~w11053;
assign w11055 = ~w10862 & w11054;
assign w11056 = w11054 & ~w11055;
assign w11057 = ~w11054 & ~w10862;
assign w11058 = ~w11056 & ~w11057;
assign w11059 = (~w10725 & w10729) | (~w10725 & w27244) | (w10729 & w27244);
assign w11060 = w11058 & w11059;
assign w11061 = ~w11058 & ~w11059;
assign w11062 = ~w11060 & ~w11061;
assign w11063 = b_38 & w1694;
assign w11064 = w1834 & w29568;
assign w11065 = b_37 & w1689;
assign w11066 = ~w11064 & ~w11065;
assign w11067 = ~w11063 & w11066;
assign w11068 = (w11067 & ~w4658) | (w11067 & w25621) | (~w4658 & w25621);
assign w11069 = (w4658 & w25880) | (w4658 & w25881) | (w25880 & w25881);
assign w11070 = (~w4658 & w29569) | (~w4658 & w29570) | (w29569 & w29570);
assign w11071 = ~w11068 & ~w11069;
assign w11072 = ~w11070 & ~w11071;
assign w11073 = w11062 & ~w11072;
assign w11074 = w11062 & ~w11073;
assign w11075 = ~w11062 & ~w11072;
assign w11076 = ~w11074 & ~w11075;
assign w11077 = (~w10743 & w10746) | (~w10743 & w27245) | (w10746 & w27245);
assign w11078 = w11076 & w11077;
assign w11079 = ~w11076 & ~w11077;
assign w11080 = ~w11078 & ~w11079;
assign w11081 = b_41 & w1295;
assign w11082 = w1422 & w29571;
assign w11083 = b_40 & w1290;
assign w11084 = ~w11082 & ~w11083;
assign w11085 = ~w11081 & w11084;
assign w11086 = (w11085 & ~w5609) | (w11085 & w25434) | (~w5609 & w25434);
assign w11087 = (w5609 & w25622) | (w5609 & w25623) | (w25622 & w25623);
assign w11088 = (~w5609 & w25882) | (~w5609 & w25883) | (w25882 & w25883);
assign w11089 = ~w11086 & ~w11087;
assign w11090 = ~w11088 & ~w11089;
assign w11091 = w11080 & ~w11090;
assign w11092 = ~w11080 & w11090;
assign w11093 = (~w11092 & w10767) | (~w11092 & w25115) | (w10767 & w25115);
assign w11094 = (w10767 & w26216) | (w10767 & w26217) | (w26216 & w26217);
assign w11095 = ~w10852 & ~w11094;
assign w11096 = (~w10767 & w26643) | (~w10767 & w26644) | (w26643 & w26644);
assign w11097 = w26217 & ~w11093;
assign w11098 = b_44 & w986;
assign w11099 = w1069 & w29572;
assign w11100 = b_43 & w981;
assign w11101 = ~w11099 & ~w11100;
assign w11102 = ~w11098 & w11101;
assign w11103 = (w11102 & ~w6408) | (w11102 & w25624) | (~w6408 & w25624);
assign w11104 = (w6408 & w25884) | (w6408 & w25885) | (w25884 & w25885);
assign w11105 = (~w6408 & w26218) | (~w6408 & w26219) | (w26218 & w26219);
assign w11106 = ~w11103 & ~w11104;
assign w11107 = ~w11105 & ~w11106;
assign w11108 = (~w11107 & w11095) | (~w11107 & w27752) | (w11095 & w27752);
assign w11109 = (w11107 & w11095) | (w11107 & w27831) | (w11095 & w27831);
assign w11110 = ~w11095 & w27832;
assign w11111 = ~w11109 & ~w11110;
assign w11112 = ~w10783 & w11111;
assign w11113 = w10783 & ~w11111;
assign w11114 = ~w11112 & ~w11113;
assign w11115 = b_47 & w657;
assign w11116 = w754 & w29573;
assign w11117 = b_46 & w652;
assign w11118 = ~w11116 & ~w11117;
assign w11119 = ~w11115 & w11118;
assign w11120 = (w11119 & ~w6998) | (w11119 & w25435) | (~w6998 & w25435);
assign w11121 = (w6998 & w25625) | (w6998 & w25626) | (w25625 & w25626);
assign w11122 = (~w6998 & w25886) | (~w6998 & w25887) | (w25886 & w25887);
assign w11123 = ~w11120 & ~w11121;
assign w11124 = ~w11122 & ~w11123;
assign w11125 = ~w11114 & ~w11124;
assign w11126 = w11114 & w11124;
assign w11127 = ~w11125 & ~w11126;
assign w11128 = (~w27179 & w27833) | (~w27179 & w27834) | (w27833 & w27834);
assign w11129 = (w27179 & w27835) | (w27179 & w27836) | (w27835 & w27836);
assign w11130 = ~w11128 & ~w11129;
assign w11131 = ~w10851 & w11130;
assign w11132 = w11130 & ~w11131;
assign w11133 = ~w11130 & ~w10851;
assign w11134 = ~w11132 & ~w11133;
assign w11135 = ~w10841 & ~w11134;
assign w11136 = w10841 & w11134;
assign w11137 = ~w11135 & ~w11136;
assign w11138 = ~w10840 & w11137;
assign w11139 = ~w11137 & ~w10840;
assign w11140 = w11137 & ~w11138;
assign w11141 = ~w11139 & ~w11140;
assign w11142 = ~w10830 & ~w11141;
assign w11143 = ~w10830 & ~w11142;
assign w11144 = w10830 & ~w11141;
assign w11145 = ~w11143 & ~w11144;
assign w11146 = b_56 & w99;
assign w11147 = w136 & w29574;
assign w11148 = b_55 & w94;
assign w11149 = ~w11147 & ~w11148;
assign w11150 = ~w11146 & w11149;
assign w11151 = (w11150 & ~w9798) | (w11150 & w29575) | (~w9798 & w29575);
assign w11152 = (w9798 & w39934) | (w9798 & w39935) | (w39934 & w39935);
assign w11153 = (~w9798 & w39936) | (~w9798 & w39937) | (w39936 & w39937);
assign w11154 = ~w11151 & ~w11152;
assign w11155 = ~w11153 & ~w11154;
assign w11156 = (~w11155 & w11143) | (~w11155 & w26220) | (w11143 & w26220);
assign w11157 = ~w11145 & ~w11156;
assign w11158 = ~w11143 & w39938;
assign w11159 = w8 & w29576;
assign w11160 = ~w8 & w29577;
assign w11161 = b_58 & w4;
assign w11162 = ~w11160 & ~w11161;
assign w11163 = ~w11159 & w11162;
assign w11164 = ~b_58 & ~b_59;
assign w11165 = b_58 & b_59;
assign w11166 = ~w11164 & ~w11165;
assign w11167 = (w6406 & w39939) | (w6406 & w39940) | (w39939 & w39940);
assign w11168 = (~w6406 & w39941) | (~w6406 & w39942) | (w39941 & w39942);
assign w11169 = ~w11167 & ~w11168;
assign w11170 = (w11163 & ~w11169) | (w11163 & w29584) | (~w11169 & w29584);
assign w11171 = (w11169 & w39943) | (w11169 & w39944) | (w39943 & w39944);
assign w11172 = (~w11169 & w39945) | (~w11169 & w39946) | (w39945 & w39946);
assign w11173 = ~w11170 & ~w11171;
assign w11174 = ~w11172 & ~w11173;
assign w11175 = (w11174 & w11157) | (w11174 & w39947) | (w11157 & w39947);
assign w11176 = ~w11157 & w39948;
assign w11177 = ~w11175 & ~w11176;
assign w11178 = ~w10829 & ~w11177;
assign w11179 = w11177 & ~w10829;
assign w11180 = ~w11177 & ~w11178;
assign w11181 = ~w11179 & ~w11180;
assign w11182 = ~w10828 & ~w11181;
assign w11183 = (w29586 & w39949) | (w29586 & w39950) | (w39949 & w39950);
assign w11184 = ~w11182 & ~w11183;
assign w11185 = (~w11157 & w39951) | (~w11157 & w39952) | (w39951 & w39952);
assign w11186 = b_60 & w9;
assign w11187 = ~w8 & w29589;
assign w11188 = b_59 & w4;
assign w11189 = ~w11187 & ~w11188;
assign w11190 = ~w11186 & w11189;
assign w11191 = ~b_59 & ~b_60;
assign w11192 = b_59 & b_60;
assign w11193 = ~w11191 & ~w11192;
assign w11194 = (w6406 & w39953) | (w6406 & w39954) | (w39953 & w39954);
assign w11195 = (~w6406 & w39955) | (~w6406 & w39956) | (w39955 & w39956);
assign w11196 = ~w11194 & ~w11195;
assign w11197 = (w11190 & ~w11196) | (w11190 & w29595) | (~w11196 & w29595);
assign w11198 = (w11196 & w39957) | (w11196 & w39958) | (w39957 & w39958);
assign w11199 = (~w11196 & w39959) | (~w11196 & w39960) | (w39959 & w39960);
assign w11200 = ~w11197 & ~w11198;
assign w11201 = ~w11199 & ~w11200;
assign w11202 = b_57 & w99;
assign w11203 = w136 & w29596;
assign w11204 = b_56 & w94;
assign w11205 = ~w11203 & ~w11204;
assign w11206 = ~w11202 & w11205;
assign w11207 = (w11206 & ~w10452) | (w11206 & w29597) | (~w10452 & w29597);
assign w11208 = (w10452 & w39961) | (w10452 & w39962) | (w39961 & w39962);
assign w11209 = (~w10452 & w39963) | (~w10452 & w39964) | (w39963 & w39964);
assign w11210 = ~w11207 & ~w11208;
assign w11211 = ~w11209 & ~w11210;
assign w11212 = (~w11138 & w10830) | (~w11138 & w26225) | (w10830 & w26225);
assign w11213 = b_54 & w239;
assign w11214 = w266 & w29598;
assign w11215 = b_53 & w234;
assign w11216 = ~w11214 & ~w11215;
assign w11217 = ~w11213 & w11216;
assign w11218 = (w11217 & ~w9134) | (w11217 & w29599) | (~w9134 & w29599);
assign w11219 = (w9134 & w39965) | (w9134 & w39966) | (w39965 & w39966);
assign w11220 = (~w9134 & w39967) | (~w9134 & w39968) | (w39967 & w39968);
assign w11221 = ~w11218 & ~w11219;
assign w11222 = ~w11220 & ~w11221;
assign w11223 = (~w11131 & w11134) | (~w11131 & w27547) | (w11134 & w27547);
assign w11224 = b_51 & w418;
assign w11225 = w481 & w29600;
assign w11226 = b_50 & w413;
assign w11227 = ~w11225 & ~w11226;
assign w11228 = ~w11224 & w11227;
assign w11229 = (w11228 & ~w8186) | (w11228 & w25888) | (~w8186 & w25888);
assign w11230 = (w8186 & w26226) | (w8186 & w26227) | (w26226 & w26227);
assign w11231 = (~w8186 & w29601) | (~w8186 & w29602) | (w29601 & w29602);
assign w11232 = ~w11229 & ~w11230;
assign w11233 = ~w11231 & ~w11232;
assign w11234 = (~w11125 & ~w11127) | (~w11125 & w27180) | (~w11127 & w27180);
assign w11235 = b_48 & w657;
assign w11236 = w754 & w29603;
assign w11237 = b_47 & w652;
assign w11238 = ~w11236 & ~w11237;
assign w11239 = ~w11235 & w11238;
assign w11240 = (w11239 & ~w7284) | (w11239 & w25627) | (~w7284 & w25627);
assign w11241 = (w7284 & w25889) | (w7284 & w25890) | (w25889 & w25890);
assign w11242 = (~w7284 & w26228) | (~w7284 & w26229) | (w26228 & w26229);
assign w11243 = ~w11240 & ~w11241;
assign w11244 = ~w11242 & ~w11243;
assign w11245 = (~w11108 & w11111) | (~w11108 & w25119) | (w11111 & w25119);
assign w11246 = b_45 & w986;
assign w11247 = w1069 & w29604;
assign w11248 = b_44 & w981;
assign w11249 = ~w11247 & ~w11248;
assign w11250 = ~w11246 & w11249;
assign w11251 = (w11250 & ~w6682) | (w11250 & w25628) | (~w6682 & w25628);
assign w11252 = (w6682 & w25891) | (w6682 & w25892) | (w25891 & w25892);
assign w11253 = (~w6682 & w26230) | (~w6682 & w26231) | (w26230 & w26231);
assign w11254 = ~w11251 & ~w11252;
assign w11255 = ~w11253 & ~w11254;
assign w11256 = (~w11055 & w11058) | (~w11055 & w27434) | (w11058 & w27434);
assign w11257 = (~w11050 & w10863) | (~w11050 & w27548) | (w10863 & w27548);
assign w11258 = b_33 & w2639;
assign w11259 = w2820 & w29605;
assign w11260 = b_32 & w2634;
assign w11261 = ~w11259 & ~w11260;
assign w11262 = ~w11258 & w11261;
assign w11263 = (w11262 & ~w3744) | (w11262 & w25629) | (~w3744 & w25629);
assign w11264 = (w3744 & w25893) | (w3744 & w25894) | (w25893 & w25894);
assign w11265 = (~w3744 & w26232) | (~w3744 & w26233) | (w26232 & w26233);
assign w11266 = ~w11263 & ~w11264;
assign w11267 = ~w11265 & ~w11266;
assign w11268 = (~w10982 & w10985) | (~w10982 & w27181) | (w10985 & w27181);
assign w11269 = b_21 & w5196;
assign w11270 = w5459 & w29606;
assign w11271 = b_20 & w5191;
assign w11272 = ~w11270 & ~w11271;
assign w11273 = ~w11269 & w11272;
assign w11274 = (w11273 & ~w1634) | (w11273 & w29607) | (~w1634 & w29607);
assign w11275 = (w1634 & w39969) | (w1634 & w39970) | (w39969 & w39970);
assign w11276 = (~w1634 & w39971) | (~w1634 & w39972) | (w39971 & w39972);
assign w11277 = ~w11274 & ~w11275;
assign w11278 = ~w11276 & ~w11277;
assign w11279 = (~w10964 & w10867) | (~w10964 & w25120) | (w10867 & w25120);
assign w11280 = b_18 & w5962;
assign w11281 = w6246 & w29608;
assign w11282 = b_17 & w5957;
assign w11283 = ~w11281 & ~w11282;
assign w11284 = ~w11280 & w11283;
assign w11285 = (w11284 & ~w1238) | (w11284 & w25895) | (~w1238 & w25895);
assign w11286 = (w1238 & w26234) | (w1238 & w26235) | (w26234 & w26235);
assign w11287 = (~w1238 & w29609) | (~w1238 & w29610) | (w29609 & w29610);
assign w11288 = ~w11285 & ~w11286;
assign w11289 = ~w11287 & ~w11288;
assign w11290 = (~w10957 & w10960) | (~w10957 & w26825) | (w10960 & w26825);
assign w11291 = b_15 & w6761;
assign w11292 = w7075 & w29611;
assign w11293 = b_14 & w6756;
assign w11294 = ~w11292 & ~w11293;
assign w11295 = ~w11291 & w11294;
assign w11296 = (w11295 & ~w827) | (w11295 & w29612) | (~w827 & w29612);
assign w11297 = (w827 & w39973) | (w827 & w39974) | (w39973 & w39974);
assign w11298 = (~w827 & w39975) | (~w827 & w39976) | (w39975 & w39976);
assign w11299 = ~w11296 & ~w11297;
assign w11300 = ~w11298 & ~w11299;
assign w11301 = (~w10952 & w10888) | (~w10952 & w26645) | (w10888 & w26645);
assign w11302 = b_12 & w7613;
assign w11303 = w7941 & w29613;
assign w11304 = b_11 & w7608;
assign w11305 = ~w11303 & ~w11304;
assign w11306 = ~w11302 & w11305;
assign w11307 = (w11306 & ~w552) | (w11306 & w29614) | (~w552 & w29614);
assign w11308 = (w552 & w39977) | (w552 & w39978) | (w39977 & w39978);
assign w11309 = (~w552 & w39979) | (~w552 & w39980) | (w39979 & w39980);
assign w11310 = ~w11307 & ~w11308;
assign w11311 = ~w11309 & ~w11310;
assign w11312 = ~w10946 & ~w10948;
assign w11313 = b_6 & w9534;
assign w11314 = w9876 & w29615;
assign w11315 = b_5 & w9529;
assign w11316 = ~w11314 & ~w11315;
assign w11317 = ~w11313 & w11316;
assign w11318 = (w11317 & ~w190) | (w11317 & w29616) | (~w190 & w29616);
assign w11319 = (w190 & w39981) | (w190 & w39982) | (w39981 & w39982);
assign w11320 = (~w190 & w39983) | (~w190 & w39984) | (w39983 & w39984);
assign w11321 = ~w11318 & ~w11319;
assign w11322 = ~w11320 & ~w11321;
assign w11323 = a_59 & ~a_60;
assign w11324 = ~a_59 & a_60;
assign w11325 = ~w11323 & ~w11324;
assign w11326 = b_0 & ~w11325;
assign w11327 = (w11326 & w10912) | (w11326 & w27455) | (w10912 & w27455);
assign w11328 = ~w10912 & w27456;
assign w11329 = ~w11327 & ~w11328;
assign w11330 = b_3 & w10562;
assign w11331 = w10902 & w26917;
assign w11332 = b_2 & w10557;
assign w11333 = ~w11331 & ~w11332;
assign w11334 = ~w11330 & w11333;
assign w11335 = w57 & w10565;
assign w11336 = w11334 & ~w11335;
assign w11337 = a_59 & ~w11336;
assign w11338 = w11336 & a_59;
assign w11339 = ~w11336 & ~w11337;
assign w11340 = ~w11338 & ~w11339;
assign w11341 = ~w11329 & ~w11340;
assign w11342 = w11329 & w11340;
assign w11343 = ~w11341 & ~w11342;
assign w11344 = ~w11322 & w11343;
assign w11345 = w11343 & ~w11344;
assign w11346 = ~w11343 & ~w11322;
assign w11347 = ~w11345 & w26826;
assign w11348 = (w10931 & w11345) | (w10931 & w26827) | (w11345 & w26827);
assign w11349 = ~w11347 & ~w11348;
assign w11350 = b_9 & w8526;
assign w11351 = w8886 & w29617;
assign w11352 = b_8 & w8521;
assign w11353 = ~w11351 & ~w11352;
assign w11354 = ~w11350 & w11353;
assign w11355 = (w11354 & ~w371) | (w11354 & w29618) | (~w371 & w29618);
assign w11356 = (w371 & w39985) | (w371 & w39986) | (w39985 & w39986);
assign w11357 = (~w371 & w39987) | (~w371 & w39988) | (w39987 & w39988);
assign w11358 = ~w11355 & ~w11356;
assign w11359 = ~w11357 & ~w11358;
assign w11360 = ~w11349 & ~w11359;
assign w11361 = w11349 & w11359;
assign w11362 = ~w11360 & ~w11361;
assign w11363 = ~w11312 & w11362;
assign w11364 = w11312 & ~w11362;
assign w11365 = ~w11363 & ~w11364;
assign w11366 = w11311 & ~w11365;
assign w11367 = ~w11311 & w11365;
assign w11368 = ~w11366 & ~w11367;
assign w11369 = ~w11301 & w11368;
assign w11370 = w11301 & ~w11368;
assign w11371 = ~w11369 & ~w11370;
assign w11372 = ~w11300 & w11371;
assign w11373 = w11300 & ~w11371;
assign w11374 = ~w11372 & ~w11373;
assign w11375 = ~w11290 & w11374;
assign w11376 = w11290 & ~w11374;
assign w11377 = ~w11375 & ~w11376;
assign w11378 = ~w11289 & w11377;
assign w11379 = ~w11377 & ~w11289;
assign w11380 = w11377 & ~w11378;
assign w11381 = ~w11379 & ~w11380;
assign w11382 = ~w11279 & ~w11381;
assign w11383 = w11279 & w11381;
assign w11384 = ~w11382 & ~w11383;
assign w11385 = ~w11278 & w11384;
assign w11386 = w11278 & ~w11384;
assign w11387 = ~w11385 & ~w11386;
assign w11388 = (~w10985 & w27457) | (~w10985 & w27458) | (w27457 & w27458);
assign w11389 = (w10985 & w27459) | (w10985 & w27460) | (w27459 & w27460);
assign w11390 = ~w11388 & ~w11389;
assign w11391 = b_24 & w4499;
assign w11392 = w4723 & w29619;
assign w11393 = b_23 & w4494;
assign w11394 = ~w11392 & ~w11393;
assign w11395 = ~w11391 & w11394;
assign w11396 = (w11395 & ~w2083) | (w11395 & w26236) | (~w2083 & w26236);
assign w11397 = (w2083 & w29620) | (w2083 & w29621) | (w29620 & w29621);
assign w11398 = (~w2083 & w29622) | (~w2083 & w29623) | (w29622 & w29623);
assign w11399 = ~w11396 & ~w11397;
assign w11400 = ~w11398 & ~w11399;
assign w11401 = w11390 & ~w11400;
assign w11402 = w11390 & ~w11401;
assign w11403 = ~w11390 & ~w11400;
assign w11404 = ~w11402 & ~w11403;
assign w11405 = (~w10999 & w10866) | (~w10999 & w25121) | (w10866 & w25121);
assign w11406 = w11404 & w11405;
assign w11407 = ~w11404 & ~w11405;
assign w11408 = ~w11406 & ~w11407;
assign w11409 = b_27 & w3803;
assign w11410 = w4027 & w29624;
assign w11411 = b_26 & w3798;
assign w11412 = ~w11410 & ~w11411;
assign w11413 = ~w11409 & w11412;
assign w11414 = (w11413 & ~w2582) | (w11413 & w25896) | (~w2582 & w25896);
assign w11415 = (w2582 & w26237) | (w2582 & w26238) | (w26237 & w26238);
assign w11416 = (~w2582 & w29625) | (~w2582 & w29626) | (w29625 & w29626);
assign w11417 = ~w11414 & ~w11415;
assign w11418 = ~w11416 & ~w11417;
assign w11419 = w11408 & ~w11418;
assign w11420 = w11408 & ~w11419;
assign w11421 = ~w11408 & ~w11418;
assign w11422 = ~w11420 & ~w11421;
assign w11423 = (~w11015 & w11019) | (~w11015 & w27246) | (w11019 & w27246);
assign w11424 = w11422 & w11423;
assign w11425 = ~w11422 & ~w11423;
assign w11426 = ~w11424 & ~w11425;
assign w11427 = b_30 & w3195;
assign w11428 = w3388 & w29627;
assign w11429 = b_29 & w3190;
assign w11430 = ~w11428 & ~w11429;
assign w11431 = ~w11427 & w11430;
assign w11432 = (w11431 & ~w3138) | (w11431 & w26239) | (~w3138 & w26239);
assign w11433 = (w3138 & w29628) | (w3138 & w29629) | (w29628 & w29629);
assign w11434 = (~w3138 & w29630) | (~w3138 & w29631) | (w29630 & w29631);
assign w11435 = ~w11432 & ~w11433;
assign w11436 = ~w11434 & ~w11435;
assign w11437 = ~w11426 & w11436;
assign w11438 = w11426 & ~w11436;
assign w11439 = ~w11437 & ~w11438;
assign w11440 = ~w11037 & w11439;
assign w11441 = w11037 & ~w11439;
assign w11442 = ~w11440 & ~w11441;
assign w11443 = ~w11267 & w11442;
assign w11444 = w11267 & w11442;
assign w11445 = ~w11442 & ~w11267;
assign w11446 = ~w11444 & ~w11445;
assign w11447 = ~w11257 & w11446;
assign w11448 = w11257 & ~w11446;
assign w11449 = ~w11447 & ~w11448;
assign w11450 = b_36 & w2158;
assign w11451 = w2294 & w29632;
assign w11452 = b_35 & w2153;
assign w11453 = ~w11451 & ~w11452;
assign w11454 = ~w11450 & w11453;
assign w11455 = (w11454 & ~w4395) | (w11454 & w25897) | (~w4395 & w25897);
assign w11456 = (w4395 & w26240) | (w4395 & w26241) | (w26240 & w26241);
assign w11457 = (~w4395 & w29633) | (~w4395 & w29634) | (w29633 & w29634);
assign w11458 = ~w11455 & ~w11456;
assign w11459 = ~w11457 & ~w11458;
assign w11460 = ~w11449 & ~w11459;
assign w11461 = w11449 & w11459;
assign w11462 = ~w11460 & ~w11461;
assign w11463 = w11256 & ~w11462;
assign w11464 = ~w11256 & w11462;
assign w11465 = ~w11463 & ~w11464;
assign w11466 = b_39 & w1694;
assign w11467 = w1834 & w29635;
assign w11468 = b_38 & w1689;
assign w11469 = ~w11467 & ~w11468;
assign w11470 = ~w11466 & w11469;
assign w11471 = (w11470 & ~w4888) | (w11470 & w25630) | (~w4888 & w25630);
assign w11472 = (w4888 & w25898) | (w4888 & w25899) | (w25898 & w25899);
assign w11473 = (~w4888 & w29636) | (~w4888 & w29637) | (w29636 & w29637);
assign w11474 = ~w11471 & ~w11472;
assign w11475 = ~w11473 & ~w11474;
assign w11476 = w11465 & ~w11475;
assign w11477 = w11465 & ~w11476;
assign w11478 = ~w11465 & ~w11475;
assign w11479 = ~w11477 & ~w11478;
assign w11480 = (~w11073 & w11076) | (~w11073 & w27435) | (w11076 & w27435);
assign w11481 = w11479 & w11480;
assign w11482 = ~w11479 & ~w11480;
assign w11483 = ~w11481 & ~w11482;
assign w11484 = b_42 & w1295;
assign w11485 = w1422 & w29638;
assign w11486 = b_41 & w1290;
assign w11487 = ~w11485 & ~w11486;
assign w11488 = ~w11484 & w11487;
assign w11489 = (w11488 & ~w5864) | (w11488 & w25631) | (~w5864 & w25631);
assign w11490 = (w5864 & w25900) | (w5864 & w25901) | (w25900 & w25901);
assign w11491 = (~w5864 & w26242) | (~w5864 & w26243) | (w26242 & w26243);
assign w11492 = ~w11489 & ~w11490;
assign w11493 = ~w11491 & ~w11492;
assign w11494 = ~w11483 & w11493;
assign w11495 = w11483 & ~w11493;
assign w11496 = ~w11494 & ~w11495;
assign w11497 = ~w11096 & w11496;
assign w11498 = w11096 & ~w11496;
assign w11499 = ~w11497 & ~w11498;
assign w11500 = (w11499 & w11254) | (w11499 & w26244) | (w11254 & w26244);
assign w11501 = (~w26244 & w27753) | (~w26244 & w27754) | (w27753 & w27754);
assign w11502 = ~w26244 & w27436;
assign w11503 = ~w11501 & ~w11502;
assign w11504 = ~w11245 & ~w11503;
assign w11505 = w11245 & w11503;
assign w11506 = ~w11504 & ~w11505;
assign w11507 = ~w11244 & w11506;
assign w11508 = ~w11506 & ~w11244;
assign w11509 = w11244 & w11506;
assign w11510 = ~w11508 & ~w11509;
assign w11511 = ~w11234 & ~w11510;
assign w11512 = w11234 & w11510;
assign w11513 = ~w11511 & ~w11512;
assign w11514 = ~w11233 & w11513;
assign w11515 = ~w11513 & ~w11233;
assign w11516 = w11513 & ~w11514;
assign w11517 = ~w11515 & ~w11516;
assign w11518 = ~w11223 & ~w11517;
assign w11519 = w11223 & w11517;
assign w11520 = ~w11518 & ~w11519;
assign w11521 = ~w11222 & w11520;
assign w11522 = w11222 & ~w11520;
assign w11523 = ~w11521 & ~w11522;
assign w11524 = ~w11212 & w11523;
assign w11525 = w11212 & ~w11523;
assign w11526 = ~w11524 & ~w11525;
assign w11527 = ~w11211 & w11526;
assign w11528 = w11211 & ~w11526;
assign w11529 = ~w11527 & ~w11528;
assign w11530 = ~w11201 & w11529;
assign w11531 = w11201 & ~w11529;
assign w11532 = ~w11530 & ~w11531;
assign w11533 = ~w11185 & w11532;
assign w11534 = w11185 & ~w11532;
assign w11535 = ~w11533 & ~w11534;
assign w11536 = (~w10828 & w26245) | (~w10828 & w26246) | (w26245 & w26246);
assign w11537 = (w10828 & w39989) | (w10828 & w39990) | (w39989 & w39990);
assign w11538 = ~w11536 & ~w11537;
assign w11539 = b_55 & w239;
assign w11540 = w266 & w29639;
assign w11541 = b_54 & w234;
assign w11542 = ~w11540 & ~w11541;
assign w11543 = ~w11539 & w11542;
assign w11544 = (w11543 & ~w9776) | (w11543 & w29640) | (~w9776 & w29640);
assign w11545 = (w9776 & w39991) | (w9776 & w39992) | (w39991 & w39992);
assign w11546 = (~w9776 & w39993) | (~w9776 & w39994) | (w39993 & w39994);
assign w11547 = ~w11544 & ~w11545;
assign w11548 = ~w11546 & ~w11547;
assign w11549 = ~w11514 & ~w11518;
assign w11550 = b_52 & w418;
assign w11551 = w481 & w29641;
assign w11552 = b_51 & w413;
assign w11553 = ~w11551 & ~w11552;
assign w11554 = ~w11550 & w11553;
assign w11555 = (w11554 & ~w8793) | (w11554 & w26247) | (~w8793 & w26247);
assign w11556 = (w8793 & w29642) | (w8793 & w29643) | (w29642 & w29643);
assign w11557 = (~w8793 & w29644) | (~w8793 & w29645) | (w29644 & w29645);
assign w11558 = ~w11555 & ~w11556;
assign w11559 = ~w11557 & ~w11558;
assign w11560 = (~w11507 & w11510) | (~w11507 & w27182) | (w11510 & w27182);
assign w11561 = b_49 & w657;
assign w11562 = w754 & w29646;
assign w11563 = b_48 & w652;
assign w11564 = ~w11562 & ~w11563;
assign w11565 = ~w11561 & w11564;
assign w11566 = (w11565 & ~w7859) | (w11565 & w25902) | (~w7859 & w25902);
assign w11567 = (w7859 & w26248) | (w7859 & w26249) | (w26248 & w26249);
assign w11568 = (~w7859 & w26828) | (~w7859 & w26829) | (w26828 & w26829);
assign w11569 = ~w11566 & ~w11567;
assign w11570 = ~w11568 & ~w11569;
assign w11571 = ~w11500 & ~w11504;
assign w11572 = (~w11495 & w11096) | (~w11495 & w27437) | (w11096 & w27437);
assign w11573 = (~w11443 & w11257) | (~w11443 & w25123) | (w11257 & w25123);
assign w11574 = ~w11438 & ~w11440;
assign w11575 = (~w11378 & w11279) | (~w11378 & w26830) | (w11279 & w26830);
assign w11576 = ~w11367 & ~w11369;
assign w11577 = b_10 & w8526;
assign w11578 = w8886 & w29647;
assign w11579 = b_9 & w8521;
assign w11580 = ~w11578 & ~w11579;
assign w11581 = ~w11577 & w11580;
assign w11582 = (w11581 & ~w454) | (w11581 & w29648) | (~w454 & w29648);
assign w11583 = (w454 & w39995) | (w454 & w39996) | (w39995 & w39996);
assign w11584 = (~w454 & w39997) | (~w454 & w39998) | (w39997 & w39998);
assign w11585 = ~w11582 & ~w11583;
assign w11586 = ~w11584 & ~w11585;
assign w11587 = (~w26831 & w27461) | (~w26831 & w27462) | (w27461 & w27462);
assign w11588 = b_7 & w9534;
assign w11589 = w9876 & w29649;
assign w11590 = b_6 & w9529;
assign w11591 = ~w11589 & ~w11590;
assign w11592 = ~w11588 & w11591;
assign w11593 = (w11592 & ~w213) | (w11592 & w29650) | (~w213 & w29650);
assign w11594 = (w213 & w39999) | (w213 & w40000) | (w39999 & w40000);
assign w11595 = (~w213 & w40001) | (~w213 & w40002) | (w40001 & w40002);
assign w11596 = ~w11593 & ~w11594;
assign w11597 = ~w11595 & ~w11596;
assign w11598 = ~w10912 & w29651;
assign w11599 = (~w11598 & w11329) | (~w11598 & w26832) | (w11329 & w26832);
assign w11600 = b_4 & w10562;
assign w11601 = w10902 & w26918;
assign w11602 = b_3 & w10557;
assign w11603 = ~w11601 & ~w11602;
assign w11604 = ~w11600 & w11603;
assign w11605 = w84 & w10565;
assign w11606 = w11604 & ~w11605;
assign w11607 = (a_59 & w11605) | (a_59 & w26919) | (w11605 & w26919);
assign w11608 = ~w11605 & w40003;
assign w11609 = ~w11606 & ~w11607;
assign w11610 = ~w11608 & ~w11609;
assign w11611 = (a_62 & w11325) | (a_62 & w29652) | (w11325 & w29652);
assign w11612 = ~a_60 & a_61;
assign w11613 = a_60 & ~a_61;
assign w11614 = ~w11612 & ~w11613;
assign w11615 = w11325 & ~w11614;
assign w11616 = b_0 & w11615;
assign w11617 = ~a_61 & a_62;
assign w11618 = a_61 & ~a_62;
assign w11619 = ~w11617 & ~w11618;
assign w11620 = ~w11325 & w11619;
assign w11621 = b_1 & w11620;
assign w11622 = ~w11616 & ~w11621;
assign w11623 = ~w11325 & ~w11619;
assign w11624 = ~w15 & w11623;
assign w11625 = w11622 & ~w11624;
assign w11626 = (a_62 & ~w11622) | (a_62 & w26920) | (~w11622 & w26920);
assign w11627 = w11622 & w27463;
assign w11628 = ~w11625 & ~w11626;
assign w11629 = (w11611 & w11628) | (w11611 & w27464) | (w11628 & w27464);
assign w11630 = ~w11628 & w29653;
assign w11631 = ~w11629 & ~w11630;
assign w11632 = w11610 & ~w11631;
assign w11633 = ~w11610 & w11631;
assign w11634 = ~w11632 & ~w11633;
assign w11635 = ~w11599 & w11634;
assign w11636 = w11599 & ~w11634;
assign w11637 = ~w11635 & ~w11636;
assign w11638 = w11597 & ~w11637;
assign w11639 = ~w11597 & w11637;
assign w11640 = ~w11638 & ~w11639;
assign w11641 = ~w11587 & w11640;
assign w11642 = w11587 & ~w11640;
assign w11643 = ~w11641 & ~w11642;
assign w11644 = ~w11586 & w11643;
assign w11645 = w11643 & ~w11644;
assign w11646 = ~w11643 & ~w11586;
assign w11647 = ~w11645 & ~w11646;
assign w11648 = (~w11360 & w11312) | (~w11360 & w26921) | (w11312 & w26921);
assign w11649 = w11647 & w11648;
assign w11650 = ~w11647 & ~w11648;
assign w11651 = ~w11649 & ~w11650;
assign w11652 = b_13 & w7613;
assign w11653 = w7941 & w29654;
assign w11654 = b_12 & w7608;
assign w11655 = ~w11653 & ~w11654;
assign w11656 = ~w11652 & w11655;
assign w11657 = (w11656 & ~w711) | (w11656 & w29655) | (~w711 & w29655);
assign w11658 = (w711 & w40004) | (w711 & w40005) | (w40004 & w40005);
assign w11659 = (~w711 & w40006) | (~w711 & w40007) | (w40006 & w40007);
assign w11660 = ~w11657 & ~w11658;
assign w11661 = ~w11659 & ~w11660;
assign w11662 = w11651 & ~w11661;
assign w11663 = ~w11651 & w11661;
assign w11664 = ~w11576 & w26833;
assign w11665 = ~w11576 & ~w11664;
assign w11666 = (~w11662 & w11576) | (~w11662 & w27465) | (w11576 & w27465);
assign w11667 = w11576 & w26833;
assign w11668 = ~w11665 & ~w11667;
assign w11669 = b_16 & w6761;
assign w11670 = w7075 & w29656;
assign w11671 = b_15 & w6756;
assign w11672 = ~w11670 & ~w11671;
assign w11673 = ~w11669 & w11672;
assign w11674 = (w11673 & ~w926) | (w11673 & w29657) | (~w926 & w29657);
assign w11675 = (w926 & w40008) | (w926 & w40009) | (w40008 & w40009);
assign w11676 = (~w926 & w40010) | (~w926 & w40011) | (w40010 & w40011);
assign w11677 = ~w11674 & ~w11675;
assign w11678 = ~w11676 & ~w11677;
assign w11679 = (~w11678 & w11665) | (~w11678 & w27466) | (w11665 & w27466);
assign w11680 = ~w11668 & ~w11679;
assign w11681 = ~w11665 & w27467;
assign w11682 = ~w11680 & ~w11681;
assign w11683 = (~w11372 & w11290) | (~w11372 & w27183) | (w11290 & w27183);
assign w11684 = ~w11680 & w27184;
assign w11685 = (~w11683 & w11680) | (~w11683 & w27185) | (w11680 & w27185);
assign w11686 = ~w11684 & ~w11685;
assign w11687 = b_19 & w5962;
assign w11688 = w6246 & w29658;
assign w11689 = b_18 & w5957;
assign w11690 = ~w11688 & ~w11689;
assign w11691 = ~w11687 & w11690;
assign w11692 = (w11691 & ~w1372) | (w11691 & w29659) | (~w1372 & w29659);
assign w11693 = (w1372 & w40012) | (w1372 & w40013) | (w40012 & w40013);
assign w11694 = (~w1372 & w40014) | (~w1372 & w40015) | (w40014 & w40015);
assign w11695 = ~w11692 & ~w11693;
assign w11696 = ~w11694 & ~w11695;
assign w11697 = w11686 & ~w11696;
assign w11698 = ~w11686 & w11696;
assign w11699 = ~w26922 & ~w11575;
assign w11700 = (~w11697 & ~w26922) | (~w11697 & w27549) | (~w26922 & w27549);
assign w11701 = w11575 & w26922;
assign w11702 = ~w11699 & ~w11701;
assign w11703 = b_22 & w5196;
assign w11704 = w5459 & w29660;
assign w11705 = b_21 & w5191;
assign w11706 = ~w11704 & ~w11705;
assign w11707 = ~w11703 & w11706;
assign w11708 = (w11707 & ~w1786) | (w11707 & w29661) | (~w1786 & w29661);
assign w11709 = (w1786 & w40016) | (w1786 & w40017) | (w40016 & w40017);
assign w11710 = (~w1786 & w40018) | (~w1786 & w40019) | (w40018 & w40019);
assign w11711 = ~w11708 & ~w11709;
assign w11712 = ~w11710 & ~w11711;
assign w11713 = (~w11712 & w11699) | (~w11712 & w27186) | (w11699 & w27186);
assign w11714 = ~w11702 & ~w11713;
assign w11715 = ~w11712 & ~w11713;
assign w11716 = ~w11714 & ~w11715;
assign w11717 = (~w11385 & w11268) | (~w11385 & w27247) | (w11268 & w27247);
assign w11718 = w11716 & w11717;
assign w11719 = ~w11716 & ~w11717;
assign w11720 = ~w11718 & ~w11719;
assign w11721 = b_25 & w4499;
assign w11722 = w4723 & w29662;
assign w11723 = b_24 & w4494;
assign w11724 = ~w11722 & ~w11723;
assign w11725 = ~w11721 & w11724;
assign w11726 = (w11725 & ~w2108) | (w11725 & w26250) | (~w2108 & w26250);
assign w11727 = (w2108 & w29663) | (w2108 & w29664) | (w29663 & w29664);
assign w11728 = (~w2108 & w29665) | (~w2108 & w29666) | (w29665 & w29666);
assign w11729 = ~w11726 & ~w11727;
assign w11730 = ~w11728 & ~w11729;
assign w11731 = w11720 & ~w11730;
assign w11732 = w11720 & ~w11731;
assign w11733 = ~w11720 & ~w11730;
assign w11734 = ~w11732 & ~w11733;
assign w11735 = (~w11401 & w11404) | (~w11401 & w27363) | (w11404 & w27363);
assign w11736 = w11734 & w11735;
assign w11737 = ~w11734 & ~w11735;
assign w11738 = ~w11736 & ~w11737;
assign w11739 = b_28 & w3803;
assign w11740 = w4027 & w29667;
assign w11741 = b_27 & w3798;
assign w11742 = ~w11740 & ~w11741;
assign w11743 = ~w11739 & w11742;
assign w11744 = (w11743 & ~w2771) | (w11743 & w25903) | (~w2771 & w25903);
assign w11745 = (w2771 & w26251) | (w2771 & w26252) | (w26251 & w26252);
assign w11746 = (~w2771 & w29668) | (~w2771 & w29669) | (w29668 & w29669);
assign w11747 = ~w11744 & ~w11745;
assign w11748 = ~w11746 & ~w11747;
assign w11749 = w11738 & ~w11748;
assign w11750 = w11738 & ~w11749;
assign w11751 = ~w11738 & ~w11748;
assign w11752 = ~w11750 & ~w11751;
assign w11753 = (~w11419 & w11423) | (~w11419 & w25124) | (w11423 & w25124);
assign w11754 = w11752 & w11753;
assign w11755 = ~w11752 & ~w11753;
assign w11756 = ~w11754 & ~w11755;
assign w11757 = b_31 & w3195;
assign w11758 = w3388 & w29670;
assign w11759 = b_30 & w3190;
assign w11760 = ~w11758 & ~w11759;
assign w11761 = ~w11757 & w11760;
assign w11762 = (w11761 & ~w3345) | (w11761 & w25632) | (~w3345 & w25632);
assign w11763 = (w3345 & w25904) | (w3345 & w25905) | (w25904 & w25905);
assign w11764 = (~w3345 & w26253) | (~w3345 & w26254) | (w26253 & w26254);
assign w11765 = ~w11762 & ~w11763;
assign w11766 = ~w11764 & ~w11765;
assign w11767 = w11756 & ~w11766;
assign w11768 = w11766 & w11756;
assign w11769 = ~w11756 & ~w11766;
assign w11770 = ~w11768 & ~w11769;
assign w11771 = ~w11574 & w11770;
assign w11772 = w11574 & ~w11770;
assign w11773 = ~w11771 & ~w11772;
assign w11774 = b_34 & w2639;
assign w11775 = w2820 & w29671;
assign w11776 = b_33 & w2634;
assign w11777 = ~w11775 & ~w11776;
assign w11778 = ~w11774 & w11777;
assign w11779 = (w11778 & ~w3967) | (w11778 & w26255) | (~w3967 & w26255);
assign w11780 = (w3967 & w29672) | (w3967 & w29673) | (w29672 & w29673);
assign w11781 = (~w3967 & w29674) | (~w3967 & w29675) | (w29674 & w29675);
assign w11782 = ~w11779 & ~w11780;
assign w11783 = ~w11781 & ~w11782;
assign w11784 = ~w11773 & ~w11783;
assign w11785 = w11773 & w11783;
assign w11786 = ~w11784 & ~w11785;
assign w11787 = w11573 & ~w11786;
assign w11788 = ~w11573 & w11786;
assign w11789 = ~w11787 & ~w11788;
assign w11790 = b_37 & w2158;
assign w11791 = w2294 & w29676;
assign w11792 = b_36 & w2153;
assign w11793 = ~w11791 & ~w11792;
assign w11794 = ~w11790 & w11793;
assign w11795 = (w11794 & ~w4636) | (w11794 & w25633) | (~w4636 & w25633);
assign w11796 = (w4636 & w25906) | (w4636 & w25907) | (w25906 & w25907);
assign w11797 = (~w4636 & w26256) | (~w4636 & w26257) | (w26256 & w26257);
assign w11798 = ~w11795 & ~w11796;
assign w11799 = ~w11797 & ~w11798;
assign w11800 = w11789 & ~w11799;
assign w11801 = w11789 & ~w11800;
assign w11802 = ~w11789 & ~w11799;
assign w11803 = ~w11801 & ~w11802;
assign w11804 = (~w11460 & w11256) | (~w11460 & w25125) | (w11256 & w25125);
assign w11805 = w11803 & w11804;
assign w11806 = ~w11803 & ~w11804;
assign w11807 = ~w11805 & ~w11806;
assign w11808 = b_40 & w1694;
assign w11809 = w1834 & w29677;
assign w11810 = b_39 & w1689;
assign w11811 = ~w11809 & ~w11810;
assign w11812 = ~w11808 & w11811;
assign w11813 = (w11812 & ~w5363) | (w11812 & w25436) | (~w5363 & w25436);
assign w11814 = (w5363 & w25634) | (w5363 & w25635) | (w25634 & w25635);
assign w11815 = (~w5363 & w25908) | (~w5363 & w25909) | (w25908 & w25909);
assign w11816 = ~w11813 & ~w11814;
assign w11817 = ~w11815 & ~w11816;
assign w11818 = w11807 & ~w11817;
assign w11819 = w11817 & w11807;
assign w11820 = ~w11807 & ~w11817;
assign w11821 = ~w11819 & ~w11820;
assign w11822 = ~w11476 & ~w11482;
assign w11823 = ~w11482 & w29678;
assign w11824 = (~w11821 & w11482) | (~w11821 & w29679) | (w11482 & w29679);
assign w11825 = ~w11823 & ~w11824;
assign w11826 = b_43 & w1295;
assign w11827 = w1422 & w29680;
assign w11828 = b_42 & w1290;
assign w11829 = ~w11827 & ~w11828;
assign w11830 = ~w11826 & w11829;
assign w11831 = (w11830 & ~w5888) | (w11830 & w25910) | (~w5888 & w25910);
assign w11832 = (w5888 & w26258) | (w5888 & w26259) | (w26258 & w26259);
assign w11833 = (~w5888 & w26646) | (~w5888 & w26647) | (w26646 & w26647);
assign w11834 = ~w11831 & ~w11832;
assign w11835 = ~w11833 & ~w11834;
assign w11836 = w11825 & ~w11835;
assign w11837 = ~w11825 & w11835;
assign w11838 = ~w11572 & w26260;
assign w11839 = ~w11572 & ~w11838;
assign w11840 = (~w11836 & w11572) | (~w11836 & w29681) | (w11572 & w29681);
assign w11841 = (w26648 & w26260) | (w26648 & w27364) | (w26260 & w27364);
assign w11842 = b_46 & w986;
assign w11843 = w1069 & w29682;
assign w11844 = b_45 & w981;
assign w11845 = ~w11843 & ~w11844;
assign w11846 = ~w11842 & w11845;
assign w11847 = (w11846 & ~w6974) | (w11846 & w25911) | (~w6974 & w25911);
assign w11848 = (w6974 & w26261) | (w6974 & w26262) | (w26261 & w26262);
assign w11849 = (~w6974 & w26649) | (~w6974 & w26650) | (w26649 & w26650);
assign w11850 = ~w11847 & ~w11848;
assign w11851 = ~w11849 & ~w11850;
assign w11852 = ~w11839 & w37618;
assign w11853 = (~w11851 & w11839) | (~w11851 & w37619) | (w11839 & w37619);
assign w11854 = ~w11852 & ~w11853;
assign w11855 = ~w11571 & w11854;
assign w11856 = w11571 & ~w11854;
assign w11857 = ~w11855 & ~w11856;
assign w11858 = w11570 & ~w11857;
assign w11859 = ~w11570 & w11857;
assign w11860 = ~w11858 & ~w11859;
assign w11861 = (w11860 & w11511) | (w11860 & w26651) | (w11511 & w26651);
assign w11862 = ~w11511 & w26652;
assign w11863 = ~w11861 & ~w11862;
assign w11864 = w11559 & ~w11863;
assign w11865 = ~w11559 & w11863;
assign w11866 = ~w11864 & ~w11865;
assign w11867 = (w11866 & w11518) | (w11866 & w26653) | (w11518 & w26653);
assign w11868 = ~w11518 & w26654;
assign w11869 = ~w11867 & ~w11868;
assign w11870 = ~w11548 & w11869;
assign w11871 = w11869 & ~w11870;
assign w11872 = ~w11869 & ~w11548;
assign w11873 = ~w11871 & ~w11872;
assign w11874 = (~w11521 & w11212) | (~w11521 & w26655) | (w11212 & w26655);
assign w11875 = w11873 & w11874;
assign w11876 = ~w11873 & ~w11874;
assign w11877 = ~w11875 & ~w11876;
assign w11878 = b_58 & w99;
assign w11879 = w136 & w29683;
assign w11880 = b_57 & w94;
assign w11881 = ~w11879 & ~w11880;
assign w11882 = ~w11878 & w11881;
assign w11883 = (w11882 & ~w10476) | (w11882 & w29684) | (~w10476 & w29684);
assign w11884 = (w10476 & w40020) | (w10476 & w40021) | (w40020 & w40021);
assign w11885 = (~w10476 & w40022) | (~w10476 & w40023) | (w40022 & w40023);
assign w11886 = ~w11883 & ~w11884;
assign w11887 = ~w11885 & ~w11886;
assign w11888 = ~w11877 & w11887;
assign w11889 = w11877 & ~w11887;
assign w11890 = ~w11888 & ~w11889;
assign w11891 = w8 & w29685;
assign w11892 = ~w8 & w29686;
assign w11893 = b_60 & w4;
assign w11894 = ~w11892 & ~w11893;
assign w11895 = ~w11891 & w11894;
assign w11896 = ~b_60 & ~b_61;
assign w11897 = b_60 & b_61;
assign w11898 = ~w11896 & ~w11897;
assign w11899 = (w6406 & w40024) | (w6406 & w40025) | (w40024 & w40025);
assign w11900 = (~w6406 & w40026) | (~w6406 & w40027) | (w40026 & w40027);
assign w11901 = ~w11899 & ~w11900;
assign w11902 = (w11895 & ~w11901) | (w11895 & w29692) | (~w11901 & w29692);
assign w11903 = (w11901 & w40028) | (w11901 & w40029) | (w40028 & w40029);
assign w11904 = (~w11901 & w40030) | (~w11901 & w40031) | (w40030 & w40031);
assign w11905 = ~w11902 & ~w11903;
assign w11906 = ~w11904 & ~w11905;
assign w11907 = w11890 & ~w11906;
assign w11908 = w11890 & ~w11907;
assign w11909 = (~w11527 & ~w11529) | (~w11527 & w29693) | (~w11529 & w29693);
assign w11910 = ~w11908 & w26834;
assign w11911 = (~w11909 & w11908) | (~w11909 & w26835) | (w11908 & w26835);
assign w11912 = ~w11910 & ~w11911;
assign w11913 = ~w11533 & ~w11536;
assign w11914 = (w11912 & w11536) | (w11912 & w26656) | (w11536 & w26656);
assign w11915 = ~w11912 & w11913;
assign w11916 = ~w11914 & ~w11915;
assign w11917 = (~w26656 & w29694) | (~w26656 & w29695) | (w29694 & w29695);
assign w11918 = (~w11889 & ~w11890) | (~w11889 & w29696) | (~w11890 & w29696);
assign w11919 = (~w11865 & w11549) | (~w11865 & w26263) | (w11549 & w26263);
assign w11920 = (~w11859 & w11560) | (~w11859 & w26264) | (w11560 & w26264);
assign w11921 = b_50 & w657;
assign w11922 = w754 & w29697;
assign w11923 = b_49 & w652;
assign w11924 = ~w11922 & ~w11923;
assign w11925 = ~w11921 & w11924;
assign w11926 = (w11925 & ~w8162) | (w11925 & w25912) | (~w8162 & w25912);
assign w11927 = (w8162 & w26265) | (w8162 & w26266) | (w26265 & w26266);
assign w11928 = (~w8162 & w29698) | (~w8162 & w29699) | (w29698 & w29699);
assign w11929 = ~w11926 & ~w11927;
assign w11930 = ~w11928 & ~w11929;
assign w11931 = (~w11818 & w11822) | (~w11818 & w25126) | (w11822 & w25126);
assign w11932 = (~w11767 & w11574) | (~w11767 & w25127) | (w11574 & w25127);
assign w11933 = (~w11713 & w11716) | (~w11713 & w27248) | (w11716 & w27248);
assign w11934 = (~w11679 & w11682) | (~w11679 & w27070) | (w11682 & w27070);
assign w11935 = b_17 & w6761;
assign w11936 = w7075 & w29700;
assign w11937 = b_16 & w6756;
assign w11938 = ~w11936 & ~w11937;
assign w11939 = ~w11935 & w11938;
assign w11940 = (w11939 & ~w1038) | (w11939 & w29701) | (~w1038 & w29701);
assign w11941 = (w1038 & w40032) | (w1038 & w40033) | (w40032 & w40033);
assign w11942 = (~w1038 & w40034) | (~w1038 & w40035) | (w40034 & w40035);
assign w11943 = ~w11940 & ~w11941;
assign w11944 = ~w11942 & ~w11943;
assign w11945 = b_14 & w7613;
assign w11946 = w7941 & w29702;
assign w11947 = b_13 & w7608;
assign w11948 = ~w11946 & ~w11947;
assign w11949 = ~w11945 & w11948;
assign w11950 = (w11949 & ~w735) | (w11949 & w29703) | (~w735 & w29703);
assign w11951 = (w735 & w40036) | (w735 & w40037) | (w40036 & w40037);
assign w11952 = (~w735 & w40038) | (~w735 & w40039) | (w40038 & w40039);
assign w11953 = ~w11950 & ~w11951;
assign w11954 = ~w11952 & ~w11953;
assign w11955 = (~w11644 & w11647) | (~w11644 & w27071) | (w11647 & w27071);
assign w11956 = b_11 & w8526;
assign w11957 = w8886 & w29704;
assign w11958 = b_10 & w8521;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = ~w11956 & w11959;
assign w11961 = (w11960 & ~w530) | (w11960 & w29705) | (~w530 & w29705);
assign w11962 = (w530 & w40040) | (w530 & w40041) | (w40040 & w40041);
assign w11963 = (~w530 & w40042) | (~w530 & w40043) | (w40042 & w40043);
assign w11964 = ~w11961 & ~w11962;
assign w11965 = ~w11963 & ~w11964;
assign w11966 = (~w11639 & w11587) | (~w11639 & w27187) | (w11587 & w27187);
assign w11967 = (~w11633 & w11599) | (~w11633 & w26923) | (w11599 & w26923);
assign w11968 = b_2 & w11620;
assign w11969 = w11325 & ~w11619;
assign w11970 = w11969 & w26924;
assign w11971 = b_1 & w11615;
assign w11972 = ~w11970 & ~w11971;
assign w11973 = ~w11968 & w11972;
assign w11974 = w35 & w11623;
assign w11975 = w11973 & ~w11974;
assign w11976 = (a_62 & ~w11973) | (a_62 & w26925) | (~w11973 & w26925);
assign w11977 = w11973 & w27468;
assign w11978 = ~w11975 & ~w11976;
assign w11979 = ~w11977 & ~w11978;
assign w11980 = ~w11629 & w11979;
assign w11981 = w11629 & ~w11979;
assign w11982 = ~w11980 & ~w11981;
assign w11983 = b_5 & w10562;
assign w11984 = w10902 & w29706;
assign w11985 = b_4 & w10557;
assign w11986 = ~w11984 & ~w11985;
assign w11987 = ~w11983 & w11986;
assign w11988 = w129 & w10565;
assign w11989 = w11987 & ~w11988;
assign w11990 = (a_59 & w11988) | (a_59 & w29707) | (w11988 & w29707);
assign w11991 = ~w11988 & w40044;
assign w11992 = ~w11989 & ~w11990;
assign w11993 = ~w11991 & ~w11992;
assign w11994 = w11982 & ~w11993;
assign w11995 = ~w11982 & w11993;
assign w11996 = ~w11967 & w26926;
assign w11997 = ~w11967 & ~w11996;
assign w11998 = (~w11994 & w11967) | (~w11994 & w27188) | (w11967 & w27188);
assign w11999 = ~w11995 & w11998;
assign w12000 = ~w11997 & ~w11999;
assign w12001 = b_8 & w9534;
assign w12002 = w9876 & w29708;
assign w12003 = b_7 & w9529;
assign w12004 = ~w12002 & ~w12003;
assign w12005 = ~w12001 & w12004;
assign w12006 = ~w308 & w29709;
assign w12007 = (w12005 & ~w29709) | (w12005 & w40045) | (~w29709 & w40045);
assign w12008 = (w29709 & w40046) | (w29709 & w40047) | (w40046 & w40047);
assign w12009 = ~w12006 & w29711;
assign w12010 = ~w12007 & ~w12008;
assign w12011 = ~w12009 & ~w12010;
assign w12012 = w12000 & w12011;
assign w12013 = ~w12000 & ~w12011;
assign w12014 = ~w12012 & ~w12013;
assign w12015 = ~w11966 & w12014;
assign w12016 = w11966 & ~w12014;
assign w12017 = ~w12015 & ~w12016;
assign w12018 = w11965 & ~w12017;
assign w12019 = ~w11965 & w12017;
assign w12020 = ~w12018 & ~w12019;
assign w12021 = ~w11955 & w12020;
assign w12022 = w11955 & ~w12020;
assign w12023 = ~w12021 & ~w12022;
assign w12024 = ~w11954 & w12023;
assign w12025 = w12023 & ~w12024;
assign w12026 = ~w12023 & ~w11954;
assign w12027 = ~w12025 & ~w12026;
assign w12028 = ~w11666 & ~w12027;
assign w12029 = w11666 & w12027;
assign w12030 = ~w12028 & ~w12029;
assign w12031 = ~w11944 & w12030;
assign w12032 = ~w12030 & ~w11944;
assign w12033 = w12030 & ~w12031;
assign w12034 = ~w12032 & ~w12033;
assign w12035 = ~w11934 & ~w12034;
assign w12036 = w12034 & ~w11934;
assign w12037 = ~w12034 & ~w12035;
assign w12038 = ~w12036 & ~w12037;
assign w12039 = b_20 & w5962;
assign w12040 = w6246 & w29712;
assign w12041 = b_19 & w5957;
assign w12042 = ~w12040 & ~w12041;
assign w12043 = ~w12039 & w12042;
assign w12044 = (w12043 & ~w1503) | (w12043 & w29713) | (~w1503 & w29713);
assign w12045 = (w1503 & w40048) | (w1503 & w40049) | (w40048 & w40049);
assign w12046 = (~w1503 & w40050) | (~w1503 & w40051) | (w40050 & w40051);
assign w12047 = ~w12044 & ~w12045;
assign w12048 = ~w12046 & ~w12047;
assign w12049 = (~w12048 & w12037) | (~w12048 & w27469) | (w12037 & w27469);
assign w12050 = ~w12038 & ~w12049;
assign w12051 = ~w12037 & w27470;
assign w12052 = ~w12050 & w27189;
assign w12053 = (w11700 & w12050) | (w11700 & w27190) | (w12050 & w27190);
assign w12054 = ~w12052 & ~w12053;
assign w12055 = b_23 & w5196;
assign w12056 = w5459 & w29714;
assign w12057 = b_22 & w5191;
assign w12058 = ~w12056 & ~w12057;
assign w12059 = ~w12055 & w12058;
assign w12060 = (w12059 & ~w1933) | (w12059 & w29715) | (~w1933 & w29715);
assign w12061 = (w1933 & w40052) | (w1933 & w40053) | (w40052 & w40053);
assign w12062 = (~w1933 & w40054) | (~w1933 & w40055) | (w40054 & w40055);
assign w12063 = ~w12060 & ~w12061;
assign w12064 = ~w12062 & ~w12063;
assign w12065 = ~w12054 & ~w12064;
assign w12066 = w12054 & w12064;
assign w12067 = ~w12065 & ~w12066;
assign w12068 = w11933 & ~w12067;
assign w12069 = ~w11933 & w12067;
assign w12070 = ~w12068 & ~w12069;
assign w12071 = b_26 & w4499;
assign w12072 = w4723 & w29716;
assign w12073 = b_25 & w4494;
assign w12074 = ~w12072 & ~w12073;
assign w12075 = ~w12071 & w12074;
assign w12076 = (w12075 & ~w2416) | (w12075 & w26267) | (~w2416 & w26267);
assign w12077 = (w2416 & w29717) | (w2416 & w29718) | (w29717 & w29718);
assign w12078 = (~w2416 & w29719) | (~w2416 & w29720) | (w29719 & w29720);
assign w12079 = ~w12076 & ~w12077;
assign w12080 = ~w12078 & ~w12079;
assign w12081 = w12070 & ~w12080;
assign w12082 = w12070 & ~w12081;
assign w12083 = ~w12070 & ~w12080;
assign w12084 = ~w12082 & ~w12083;
assign w12085 = (~w11731 & w11734) | (~w11731 & w27550) | (w11734 & w27550);
assign w12086 = w12084 & w12085;
assign w12087 = ~w12084 & ~w12085;
assign w12088 = ~w12086 & ~w12087;
assign w12089 = b_29 & w3803;
assign w12090 = w4027 & w29721;
assign w12091 = b_28 & w3798;
assign w12092 = ~w12090 & ~w12091;
assign w12093 = ~w12089 & w12092;
assign w12094 = (w12093 & ~w2954) | (w12093 & w25913) | (~w2954 & w25913);
assign w12095 = (w2954 & w26268) | (w2954 & w26269) | (w26268 & w26269);
assign w12096 = (~w2954 & w29722) | (~w2954 & w29723) | (w29722 & w29723);
assign w12097 = ~w12094 & ~w12095;
assign w12098 = ~w12096 & ~w12097;
assign w12099 = w12088 & ~w12098;
assign w12100 = w12088 & ~w12099;
assign w12101 = ~w12088 & ~w12098;
assign w12102 = ~w12100 & ~w12101;
assign w12103 = (~w11749 & w11752) | (~w11749 & w27471) | (w11752 & w27471);
assign w12104 = w12102 & w12103;
assign w12105 = ~w12102 & ~w12103;
assign w12106 = ~w12104 & ~w12105;
assign w12107 = b_32 & w3195;
assign w12108 = w3388 & w29724;
assign w12109 = b_31 & w3190;
assign w12110 = ~w12108 & ~w12109;
assign w12111 = ~w12107 & w12110;
assign w12112 = (w12111 & ~w3545) | (w12111 & w25914) | (~w3545 & w25914);
assign w12113 = (w3545 & w26270) | (w3545 & w26271) | (w26270 & w26271);
assign w12114 = (~w3545 & w29725) | (~w3545 & w29726) | (w29725 & w29726);
assign w12115 = ~w12112 & ~w12113;
assign w12116 = ~w12114 & ~w12115;
assign w12117 = w12106 & ~w12116;
assign w12118 = ~w12106 & w12116;
assign w12119 = ~w11932 & w25128;
assign w12120 = ~w11932 & ~w12119;
assign w12121 = (~w12117 & w11932) | (~w12117 & w26272) | (w11932 & w26272);
assign w12122 = (w26272 & w25128) | (w26272 & w27249) | (w25128 & w27249);
assign w12123 = ~w12120 & ~w12122;
assign w12124 = b_35 & w2639;
assign w12125 = w2820 & w29727;
assign w12126 = b_34 & w2634;
assign w12127 = ~w12125 & ~w12126;
assign w12128 = ~w12124 & w12127;
assign w12129 = (w12128 & ~w4181) | (w12128 & w26273) | (~w4181 & w26273);
assign w12130 = (w4181 & w29728) | (w4181 & w29729) | (w29728 & w29729);
assign w12131 = (~w4181 & w29730) | (~w4181 & w29731) | (w29730 & w29731);
assign w12132 = ~w12129 & ~w12130;
assign w12133 = ~w12131 & ~w12132;
assign w12134 = (~w12133 & w12120) | (~w12133 & w27755) | (w12120 & w27755);
assign w12135 = ~w12123 & ~w12134;
assign w12136 = ~w12120 & w27756;
assign w12137 = ~w12135 & ~w12136;
assign w12138 = (~w11784 & w11573) | (~w11784 & w26274) | (w11573 & w26274);
assign w12139 = ~w12135 & w27551;
assign w12140 = (~w12138 & w12135) | (~w12138 & w27552) | (w12135 & w27552);
assign w12141 = ~w12139 & ~w12140;
assign w12142 = b_38 & w2158;
assign w12143 = w2294 & w29732;
assign w12144 = b_37 & w2153;
assign w12145 = ~w12143 & ~w12144;
assign w12146 = ~w12142 & w12145;
assign w12147 = (w12146 & ~w4658) | (w12146 & w25915) | (~w4658 & w25915);
assign w12148 = (w4658 & w26275) | (w4658 & w26276) | (w26275 & w26276);
assign w12149 = (~w4658 & w29733) | (~w4658 & w29734) | (w29733 & w29734);
assign w12150 = ~w12147 & ~w12148;
assign w12151 = ~w12149 & ~w12150;
assign w12152 = w12141 & ~w12151;
assign w12153 = w12141 & ~w12152;
assign w12154 = ~w12141 & ~w12151;
assign w12155 = ~w12153 & ~w12154;
assign w12156 = (~w11800 & w11803) | (~w11800 & w26277) | (w11803 & w26277);
assign w12157 = w12155 & w12156;
assign w12158 = ~w12155 & ~w12156;
assign w12159 = ~w12157 & ~w12158;
assign w12160 = b_41 & w1694;
assign w12161 = w1834 & w29735;
assign w12162 = b_40 & w1689;
assign w12163 = ~w12161 & ~w12162;
assign w12164 = ~w12160 & w12163;
assign w12165 = (w12164 & ~w5609) | (w12164 & w25636) | (~w5609 & w25636);
assign w12166 = (w5609 & w25916) | (w5609 & w25917) | (w25916 & w25917);
assign w12167 = (~w5609 & w26278) | (~w5609 & w26279) | (w26278 & w26279);
assign w12168 = ~w12165 & ~w12166;
assign w12169 = ~w12167 & ~w12168;
assign w12170 = w12159 & ~w12169;
assign w12171 = ~w12159 & w12169;
assign w12172 = ~w11931 & w25129;
assign w12173 = ~w11931 & ~w12172;
assign w12174 = (~w12170 & w11931) | (~w12170 & w25918) | (w11931 & w25918);
assign w12175 = (w25918 & w25129) | (w25918 & w26280) | (w25129 & w26280);
assign w12176 = ~w12173 & ~w12175;
assign w12177 = b_44 & w1295;
assign w12178 = w1422 & w29736;
assign w12179 = b_43 & w1290;
assign w12180 = ~w12178 & ~w12179;
assign w12181 = ~w12177 & w12180;
assign w12182 = (w12181 & ~w6408) | (w12181 & w25637) | (~w6408 & w25637);
assign w12183 = (w6408 & w25919) | (w6408 & w25920) | (w25919 & w25920);
assign w12184 = (~w6408 & w26281) | (~w6408 & w26282) | (w26281 & w26282);
assign w12185 = ~w12182 & ~w12183;
assign w12186 = ~w12184 & ~w12185;
assign w12187 = ~w12176 & ~w12186;
assign w12188 = w12186 & ~w12176;
assign w12189 = w12176 & ~w12186;
assign w12190 = ~w12188 & ~w12189;
assign w12191 = ~w11840 & w12190;
assign w12192 = w11840 & ~w12190;
assign w12193 = ~w12191 & ~w12192;
assign w12194 = b_47 & w986;
assign w12195 = w1069 & w29737;
assign w12196 = b_46 & w981;
assign w12197 = ~w12195 & ~w12196;
assign w12198 = ~w12194 & w12197;
assign w12199 = (w12198 & ~w6998) | (w12198 & w25437) | (~w6998 & w25437);
assign w12200 = (w6998 & w25638) | (w6998 & w25639) | (w25638 & w25639);
assign w12201 = (~w6998 & w25921) | (~w6998 & w25922) | (w25921 & w25922);
assign w12202 = ~w12199 & ~w12200;
assign w12203 = ~w12201 & ~w12202;
assign w12204 = ~w12193 & ~w12203;
assign w12205 = w12193 & w12203;
assign w12206 = ~w12204 & ~w12205;
assign w12207 = (w12206 & w11855) | (w12206 & w25130) | (w11855 & w25130);
assign w12208 = ~w12206 & w26283;
assign w12209 = ~w12207 & ~w12208;
assign w12210 = ~w12207 & w26284;
assign w12211 = w12209 & ~w12210;
assign w12212 = (~w11930 & w12207) | (~w11930 & w26657) | (w12207 & w26657);
assign w12213 = ~w12211 & ~w12212;
assign w12214 = ~w11920 & w12213;
assign w12215 = w11920 & ~w12213;
assign w12216 = ~w12214 & ~w12215;
assign w12217 = b_53 & w418;
assign w12218 = w481 & w29738;
assign w12219 = b_52 & w413;
assign w12220 = ~w12218 & ~w12219;
assign w12221 = ~w12217 & w12220;
assign w12222 = (w9109 & w40056) | (w9109 & w40057) | (w40056 & w40057);
assign w12223 = a_11 & ~w12222;
assign w12224 = w12222 & a_11;
assign w12225 = ~w12222 & ~w12223;
assign w12226 = ~w12224 & ~w12225;
assign w12227 = ~w12216 & ~w12226;
assign w12228 = w12216 & w12226;
assign w12229 = ~w12227 & ~w12228;
assign w12230 = ~w11919 & w12229;
assign w12231 = w11919 & ~w12229;
assign w12232 = ~w12230 & ~w12231;
assign w12233 = b_56 & w239;
assign w12234 = w266 & w29740;
assign w12235 = b_55 & w234;
assign w12236 = ~w12234 & ~w12235;
assign w12237 = ~w12233 & w12236;
assign w12238 = (w12237 & ~w9798) | (w12237 & w29741) | (~w9798 & w29741);
assign w12239 = (w9798 & w40058) | (w9798 & w40059) | (w40058 & w40059);
assign w12240 = (~w9798 & w40060) | (~w9798 & w40061) | (w40060 & w40061);
assign w12241 = ~w12238 & ~w12239;
assign w12242 = ~w12240 & ~w12241;
assign w12243 = ~w12232 & w12242;
assign w12244 = w12232 & ~w12242;
assign w12245 = ~w12243 & ~w12244;
assign w12246 = b_59 & w99;
assign w12247 = w136 & w29742;
assign w12248 = b_58 & w94;
assign w12249 = ~w12247 & ~w12248;
assign w12250 = ~w12246 & w12249;
assign w12251 = (w12250 & ~w25438) | (w12250 & w29743) | (~w25438 & w29743);
assign w12252 = a_5 & ~w12251;
assign w12253 = w12251 & a_5;
assign w12254 = ~w12251 & ~w12252;
assign w12255 = ~w12253 & ~w12254;
assign w12256 = w12245 & ~w12255;
assign w12257 = w12245 & ~w12256;
assign w12258 = ~w12245 & ~w12255;
assign w12259 = (~w11870 & w11873) | (~w11870 & w29744) | (w11873 & w29744);
assign w12260 = ~w12257 & w25439;
assign w12261 = (~w12259 & w12257) | (~w12259 & w25440) | (w12257 & w25440);
assign w12262 = ~w12260 & ~w12261;
assign w12263 = w8 & w29745;
assign w12264 = ~w8 & w29746;
assign w12265 = b_61 & w4;
assign w12266 = ~w12264 & ~w12265;
assign w12267 = ~w12263 & w12266;
assign w12268 = ~b_61 & ~b_62;
assign w12269 = b_61 & b_62;
assign w12270 = ~w12268 & ~w12269;
assign w12271 = (w6406 & w40062) | (w6406 & w40063) | (w40062 & w40063);
assign w12272 = (~w6406 & w40064) | (~w6406 & w40065) | (w40064 & w40065);
assign w12273 = ~w12271 & ~w12272;
assign w12274 = (w12267 & ~w12273) | (w12267 & w29752) | (~w12273 & w29752);
assign w12275 = (w12273 & w40066) | (w12273 & w40067) | (w40066 & w40067);
assign w12276 = (~w12273 & w40068) | (~w12273 & w40069) | (w40068 & w40069);
assign w12277 = ~w12274 & ~w12275;
assign w12278 = ~w12276 & ~w12277;
assign w12279 = ~w12262 & w12278;
assign w12280 = w12262 & ~w12278;
assign w12281 = ~w12279 & ~w12280;
assign w12282 = ~w11918 & w12281;
assign w12283 = w11918 & ~w12281;
assign w12284 = ~w12282 & ~w12283;
assign w12285 = (w12284 & w11914) | (w12284 & w25131) | (w11914 & w25131);
assign w12286 = w11917 & ~w12284;
assign w12287 = ~w12285 & ~w12286;
assign w12288 = (~w12210 & w11920) | (~w12210 & w25132) | (w11920 & w25132);
assign w12289 = b_51 & w657;
assign w12290 = w754 & w29753;
assign w12291 = b_50 & w652;
assign w12292 = ~w12290 & ~w12291;
assign w12293 = ~w12289 & w12292;
assign w12294 = (w12293 & ~w8186) | (w12293 & w26285) | (~w8186 & w26285);
assign w12295 = (w8186 & w29754) | (w8186 & w29755) | (w29754 & w29755);
assign w12296 = (~w8186 & w29756) | (~w8186 & w29757) | (w29756 & w29757);
assign w12297 = ~w12294 & ~w12295;
assign w12298 = ~w12296 & ~w12297;
assign w12299 = (~w25130 & w25923) | (~w25130 & w25924) | (w25923 & w25924);
assign w12300 = b_48 & w986;
assign w12301 = w1069 & w29758;
assign w12302 = b_47 & w981;
assign w12303 = ~w12301 & ~w12302;
assign w12304 = ~w12300 & w12303;
assign w12305 = (w12304 & ~w7284) | (w12304 & w25640) | (~w7284 & w25640);
assign w12306 = (w7284 & w25925) | (w7284 & w25926) | (w25925 & w25926);
assign w12307 = (~w7284 & w26286) | (~w7284 & w26287) | (w26286 & w26287);
assign w12308 = ~w12305 & ~w12306;
assign w12309 = ~w12307 & ~w12308;
assign w12310 = (~w11840 & w12189) | (~w11840 & w26658) | (w12189 & w26658);
assign w12311 = (~w12187 & w12190) | (~w12187 & w26288) | (w12190 & w26288);
assign w12312 = b_45 & w1295;
assign w12313 = w1422 & w29759;
assign w12314 = b_44 & w1290;
assign w12315 = ~w12313 & ~w12314;
assign w12316 = ~w12312 & w12315;
assign w12317 = (w12316 & ~w6682) | (w12316 & w25443) | (~w6682 & w25443);
assign w12318 = (w6682 & w25641) | (w6682 & w25642) | (w25641 & w25642);
assign w12319 = (~w6682 & w25927) | (~w6682 & w25928) | (w25927 & w25928);
assign w12320 = ~w12317 & ~w12318;
assign w12321 = ~w12319 & ~w12320;
assign w12322 = b_42 & w1694;
assign w12323 = w1834 & w29760;
assign w12324 = b_41 & w1689;
assign w12325 = ~w12323 & ~w12324;
assign w12326 = ~w12322 & w12325;
assign w12327 = (w12326 & ~w5864) | (w12326 & w25643) | (~w5864 & w25643);
assign w12328 = (w5864 & w25929) | (w5864 & w25930) | (w25929 & w25930);
assign w12329 = (~w5864 & w29761) | (~w5864 & w29762) | (w29761 & w29762);
assign w12330 = ~w12327 & ~w12328;
assign w12331 = ~w12329 & ~w12330;
assign w12332 = (~w12152 & w12155) | (~w12152 & w25444) | (w12155 & w25444);
assign w12333 = (~w12134 & w12137) | (~w12134 & w25445) | (w12137 & w25445);
assign w12334 = b_33 & w3195;
assign w12335 = w3388 & w29763;
assign w12336 = b_32 & w3190;
assign w12337 = ~w12335 & ~w12336;
assign w12338 = ~w12334 & w12337;
assign w12339 = (w12338 & ~w3744) | (w12338 & w25644) | (~w3744 & w25644);
assign w12340 = (w3744 & w25931) | (w3744 & w25932) | (w25931 & w25932);
assign w12341 = (~w3744 & w29764) | (~w3744 & w29765) | (w29764 & w29765);
assign w12342 = ~w12339 & ~w12340;
assign w12343 = ~w12341 & ~w12342;
assign w12344 = (~w26927 & w27072) | (~w26927 & w27073) | (w27072 & w27073);
assign w12345 = b_21 & w5962;
assign w12346 = w6246 & w29766;
assign w12347 = b_20 & w5957;
assign w12348 = ~w12346 & ~w12347;
assign w12349 = ~w12345 & w12348;
assign w12350 = (w12349 & ~w1634) | (w12349 & w29767) | (~w1634 & w29767);
assign w12351 = (w1634 & w40070) | (w1634 & w40071) | (w40070 & w40071);
assign w12352 = (~w1634 & w40072) | (~w1634 & w40073) | (w40072 & w40073);
assign w12353 = ~w12350 & ~w12351;
assign w12354 = ~w12352 & ~w12353;
assign w12355 = (~w12031 & w12034) | (~w12031 & w27472) | (w12034 & w27472);
assign w12356 = b_15 & w7613;
assign w12357 = w7941 & w29768;
assign w12358 = b_14 & w7608;
assign w12359 = ~w12357 & ~w12358;
assign w12360 = ~w12356 & w12359;
assign w12361 = (w12360 & ~w827) | (w12360 & w29769) | (~w827 & w29769);
assign w12362 = (w827 & w40074) | (w827 & w40075) | (w40074 & w40075);
assign w12363 = (~w827 & w40076) | (~w827 & w40077) | (w40076 & w40077);
assign w12364 = ~w12361 & ~w12362;
assign w12365 = ~w12363 & ~w12364;
assign w12366 = (~w12019 & w11955) | (~w12019 & w27365) | (w11955 & w27365);
assign w12367 = (~w12013 & ~w12014) | (~w12013 & w29770) | (~w12014 & w29770);
assign w12368 = b_9 & w9534;
assign w12369 = w9876 & w29771;
assign w12370 = b_8 & w9529;
assign w12371 = ~w12369 & ~w12370;
assign w12372 = ~w12368 & w12371;
assign w12373 = (w12372 & ~w371) | (w12372 & w29772) | (~w371 & w29772);
assign w12374 = (w371 & w40078) | (w371 & w40079) | (w40078 & w40079);
assign w12375 = (~w371 & w40080) | (~w371 & w40081) | (w40080 & w40081);
assign w12376 = ~w12373 & ~w12374;
assign w12377 = ~w12375 & ~w12376;
assign w12378 = a_62 & ~a_63;
assign w12379 = ~a_62 & a_63;
assign w12380 = ~w12378 & ~w12379;
assign w12381 = b_0 & ~w12380;
assign w12382 = ~w11979 & w27473;
assign w12383 = w11981 & ~w12382;
assign w12384 = (w12381 & w11979) | (w12381 & w27474) | (w11979 & w27474);
assign w12385 = ~w12383 & ~w12384;
assign w12386 = b_3 & w11620;
assign w12387 = w11969 & w27191;
assign w12388 = b_2 & w11615;
assign w12389 = ~w12387 & ~w12388;
assign w12390 = ~w12386 & w12389;
assign w12391 = w57 & w11623;
assign w12392 = w12390 & ~w12391;
assign w12393 = a_62 & ~w12392;
assign w12394 = w12392 & a_62;
assign w12395 = ~w12392 & ~w12393;
assign w12396 = ~w12394 & ~w12395;
assign w12397 = (~w12396 & w12383) | (~w12396 & w27074) | (w12383 & w27074);
assign w12398 = ~w12385 & ~w12397;
assign w12399 = ~w12396 & ~w12397;
assign w12400 = ~w12398 & ~w12399;
assign w12401 = b_6 & w10562;
assign w12402 = w10902 & w29773;
assign w12403 = b_5 & w10557;
assign w12404 = ~w12402 & ~w12403;
assign w12405 = ~w12401 & w12404;
assign w12406 = (w12405 & ~w190) | (w12405 & w29774) | (~w190 & w29774);
assign w12407 = (w190 & w40082) | (w190 & w40083) | (w40082 & w40083);
assign w12408 = (~w190 & w40084) | (~w190 & w40085) | (w40084 & w40085);
assign w12409 = ~w12406 & ~w12407;
assign w12410 = ~w12408 & ~w12409;
assign w12411 = w12400 & w12410;
assign w12412 = ~w12400 & ~w12410;
assign w12413 = ~w12411 & ~w12412;
assign w12414 = ~w11998 & w12413;
assign w12415 = w11998 & ~w12413;
assign w12416 = ~w12414 & ~w12415;
assign w12417 = ~w12377 & w12416;
assign w12418 = w12416 & ~w12417;
assign w12419 = ~w12416 & ~w12377;
assign w12420 = ~w12418 & ~w12419;
assign w12421 = ~w12367 & w12420;
assign w12422 = w12367 & ~w12420;
assign w12423 = ~w12421 & ~w12422;
assign w12424 = b_12 & w8526;
assign w12425 = w8886 & w29775;
assign w12426 = b_11 & w8521;
assign w12427 = ~w12425 & ~w12426;
assign w12428 = ~w12424 & w12427;
assign w12429 = (w12428 & ~w552) | (w12428 & w29776) | (~w552 & w29776);
assign w12430 = (w552 & w40086) | (w552 & w40087) | (w40086 & w40087);
assign w12431 = (~w552 & w40088) | (~w552 & w40089) | (w40088 & w40089);
assign w12432 = ~w12429 & ~w12430;
assign w12433 = ~w12431 & ~w12432;
assign w12434 = w12423 & w12433;
assign w12435 = ~w12423 & ~w12433;
assign w12436 = ~w12434 & ~w12435;
assign w12437 = ~w12366 & w12436;
assign w12438 = w12366 & ~w12436;
assign w12439 = ~w12437 & ~w12438;
assign w12440 = ~w12365 & w12439;
assign w12441 = w12439 & ~w12440;
assign w12442 = ~w12439 & ~w12365;
assign w12443 = ~w12441 & ~w12442;
assign w12444 = (~w12024 & w12027) | (~w12024 & w27475) | (w12027 & w27475);
assign w12445 = w12443 & w12444;
assign w12446 = ~w12443 & ~w12444;
assign w12447 = ~w12445 & ~w12446;
assign w12448 = b_18 & w6761;
assign w12449 = w7075 & w29777;
assign w12450 = b_17 & w6756;
assign w12451 = ~w12449 & ~w12450;
assign w12452 = ~w12448 & w12451;
assign w12453 = (w12452 & ~w1238) | (w12452 & w29778) | (~w1238 & w29778);
assign w12454 = (w1238 & w40090) | (w1238 & w40091) | (w40090 & w40091);
assign w12455 = (~w1238 & w40092) | (~w1238 & w40093) | (w40092 & w40093);
assign w12456 = ~w12453 & ~w12454;
assign w12457 = ~w12455 & ~w12456;
assign w12458 = ~w12447 & w12457;
assign w12459 = w12447 & ~w12457;
assign w12460 = ~w12458 & ~w12459;
assign w12461 = ~w12355 & w12460;
assign w12462 = w12355 & ~w12460;
assign w12463 = ~w12461 & ~w12462;
assign w12464 = ~w12354 & w12463;
assign w12465 = w12354 & ~w12463;
assign w12466 = ~w12464 & ~w12465;
assign w12467 = ~w12344 & w12466;
assign w12468 = w12344 & ~w12466;
assign w12469 = ~w12467 & ~w12468;
assign w12470 = b_24 & w5196;
assign w12471 = w5459 & w29779;
assign w12472 = b_23 & w5191;
assign w12473 = ~w12471 & ~w12472;
assign w12474 = ~w12470 & w12473;
assign w12475 = (w12474 & ~w2083) | (w12474 & w29780) | (~w2083 & w29780);
assign w12476 = (w2083 & w40094) | (w2083 & w40095) | (w40094 & w40095);
assign w12477 = (~w2083 & w40096) | (~w2083 & w40097) | (w40096 & w40097);
assign w12478 = ~w12475 & ~w12476;
assign w12479 = ~w12477 & ~w12478;
assign w12480 = w12469 & ~w12479;
assign w12481 = w12469 & ~w12480;
assign w12482 = ~w12469 & ~w12479;
assign w12483 = ~w12481 & ~w12482;
assign w12484 = (~w12065 & ~w12067) | (~w12065 & w27476) | (~w12067 & w27476);
assign w12485 = w12483 & w12484;
assign w12486 = ~w12483 & ~w12484;
assign w12487 = ~w12485 & ~w12486;
assign w12488 = b_27 & w4499;
assign w12489 = w4723 & w29781;
assign w12490 = b_26 & w4494;
assign w12491 = ~w12489 & ~w12490;
assign w12492 = ~w12488 & w12491;
assign w12493 = (w12492 & ~w2582) | (w12492 & w26289) | (~w2582 & w26289);
assign w12494 = (w2582 & w29782) | (w2582 & w29783) | (w29782 & w29783);
assign w12495 = (~w2582 & w29784) | (~w2582 & w29785) | (w29784 & w29785);
assign w12496 = ~w12493 & ~w12494;
assign w12497 = ~w12495 & ~w12496;
assign w12498 = w12487 & ~w12497;
assign w12499 = w12487 & ~w12498;
assign w12500 = ~w12487 & ~w12497;
assign w12501 = ~w12499 & ~w12500;
assign w12502 = ~w12081 & ~w12087;
assign w12503 = w12501 & w12502;
assign w12504 = ~w12501 & ~w12502;
assign w12505 = ~w12503 & ~w12504;
assign w12506 = b_30 & w3803;
assign w12507 = w4027 & w29786;
assign w12508 = b_29 & w3798;
assign w12509 = ~w12507 & ~w12508;
assign w12510 = ~w12506 & w12509;
assign w12511 = (w12510 & ~w3138) | (w12510 & w25933) | (~w3138 & w25933);
assign w12512 = (w3138 & w26290) | (w3138 & w26291) | (w26290 & w26291);
assign w12513 = (~w3138 & w29787) | (~w3138 & w29788) | (w29787 & w29788);
assign w12514 = ~w12511 & ~w12512;
assign w12515 = ~w12513 & ~w12514;
assign w12516 = ~w12505 & w12515;
assign w12517 = w12505 & ~w12515;
assign w12518 = ~w12516 & ~w12517;
assign w12519 = (~w12099 & w12102) | (~w12099 & w27477) | (w12102 & w27477);
assign w12520 = w12518 & ~w12519;
assign w12521 = ~w12518 & w12519;
assign w12522 = ~w12520 & ~w12521;
assign w12523 = ~w12343 & w12522;
assign w12524 = w12522 & ~w12523;
assign w12525 = ~w12522 & ~w12343;
assign w12526 = ~w12524 & ~w12525;
assign w12527 = ~w12121 & w12526;
assign w12528 = w12121 & ~w12526;
assign w12529 = ~w12527 & ~w12528;
assign w12530 = b_36 & w2639;
assign w12531 = w2820 & w29789;
assign w12532 = b_35 & w2634;
assign w12533 = ~w12531 & ~w12532;
assign w12534 = ~w12530 & w12533;
assign w12535 = (w12534 & ~w4395) | (w12534 & w25934) | (~w4395 & w25934);
assign w12536 = (w4395 & w29790) | (w4395 & w29791) | (w29790 & w29791);
assign w12537 = (~w4395 & w29792) | (~w4395 & w29793) | (w29792 & w29793);
assign w12538 = ~w12535 & ~w12536;
assign w12539 = ~w12537 & ~w12538;
assign w12540 = ~w12529 & ~w12539;
assign w12541 = w12529 & w12539;
assign w12542 = ~w12540 & ~w12541;
assign w12543 = w12333 & ~w12542;
assign w12544 = ~w12333 & w12542;
assign w12545 = ~w12543 & ~w12544;
assign w12546 = b_39 & w2158;
assign w12547 = w2294 & w29794;
assign w12548 = b_38 & w2153;
assign w12549 = ~w12547 & ~w12548;
assign w12550 = ~w12546 & w12549;
assign w12551 = (w12550 & ~w4888) | (w12550 & w25645) | (~w4888 & w25645);
assign w12552 = (w4888 & w25935) | (w4888 & w25936) | (w25935 & w25936);
assign w12553 = (~w4888 & w26292) | (~w4888 & w26293) | (w26292 & w26293);
assign w12554 = ~w12551 & ~w12552;
assign w12555 = ~w12553 & ~w12554;
assign w12556 = ~w12545 & w12555;
assign w12557 = w12545 & ~w12555;
assign w12558 = ~w12556 & ~w12557;
assign w12559 = ~w12332 & w12558;
assign w12560 = w12332 & ~w12558;
assign w12561 = ~w12559 & ~w12560;
assign w12562 = ~w12331 & w12561;
assign w12563 = ~w12561 & ~w12331;
assign w12564 = w12561 & ~w12562;
assign w12565 = ~w12563 & ~w12564;
assign w12566 = ~w12174 & ~w12565;
assign w12567 = w12174 & w12565;
assign w12568 = ~w12566 & ~w12567;
assign w12569 = ~w12321 & w12568;
assign w12570 = ~w12568 & ~w12321;
assign w12571 = w12321 & w12568;
assign w12572 = ~w12570 & ~w12571;
assign w12573 = ~w12311 & ~w12572;
assign w12574 = ~w12310 & w27553;
assign w12575 = ~w12573 & ~w12574;
assign w12576 = ~w12574 & w29795;
assign w12577 = (~w12309 & w12574) | (~w12309 & w29796) | (w12574 & w29796);
assign w12578 = w12575 & ~w12576;
assign w12579 = ~w12577 & ~w12578;
assign w12580 = ~w12299 & ~w12579;
assign w12581 = w12299 & w12579;
assign w12582 = ~w12580 & ~w12581;
assign w12583 = ~w12298 & w12582;
assign w12584 = w12298 & ~w12582;
assign w12585 = ~w12583 & ~w12584;
assign w12586 = ~w12288 & w12585;
assign w12587 = w12288 & ~w12585;
assign w12588 = ~w12586 & ~w12587;
assign w12589 = b_54 & w418;
assign w12590 = w481 & w29797;
assign w12591 = b_53 & w413;
assign w12592 = ~w12590 & ~w12591;
assign w12593 = ~w12589 & w12592;
assign w12594 = (w12593 & ~w9134) | (w12593 & w26294) | (~w9134 & w26294);
assign w12595 = (w9134 & w29798) | (w9134 & w29799) | (w29798 & w29799);
assign w12596 = (~w9134 & w29800) | (~w9134 & w29801) | (w29800 & w29801);
assign w12597 = ~w12594 & ~w12595;
assign w12598 = ~w12596 & ~w12597;
assign w12599 = w12588 & ~w12598;
assign w12600 = w12588 & ~w12599;
assign w12601 = ~w12588 & ~w12598;
assign w12602 = ~w12600 & ~w12601;
assign w12603 = (~w12227 & w11919) | (~w12227 & w25133) | (w11919 & w25133);
assign w12604 = w12602 & w12603;
assign w12605 = ~w12602 & ~w12603;
assign w12606 = ~w12604 & ~w12605;
assign w12607 = b_57 & w239;
assign w12608 = w266 & w29802;
assign w12609 = b_56 & w234;
assign w12610 = ~w12608 & ~w12609;
assign w12611 = ~w12607 & w12610;
assign w12612 = (w12611 & ~w10452) | (w12611 & w29803) | (~w10452 & w29803);
assign w12613 = (w10452 & w40098) | (w10452 & w40099) | (w40098 & w40099);
assign w12614 = (~w10452 & w40100) | (~w10452 & w40101) | (w40100 & w40101);
assign w12615 = ~w12612 & ~w12613;
assign w12616 = ~w12614 & ~w12615;
assign w12617 = w12606 & ~w12616;
assign w12618 = w12606 & ~w12617;
assign w12619 = b_60 & w99;
assign w12620 = w136 & w29804;
assign w12621 = b_59 & w94;
assign w12622 = ~w12620 & ~w12621;
assign w12623 = ~w12619 & w12622;
assign w12624 = (w12623 & ~w11196) | (w12623 & w27554) | (~w11196 & w27554);
assign w12625 = (w11196 & w29805) | (w11196 & w29806) | (w29805 & w29806);
assign w12626 = (~w11196 & w29807) | (~w11196 & w29808) | (w29807 & w29808);
assign w12627 = ~w12624 & ~w12625;
assign w12628 = ~w12626 & ~w12627;
assign w12629 = (w12628 & w12618) | (w12628 & w26295) | (w12618 & w26295);
assign w12630 = ~w12618 & w26296;
assign w12631 = ~w12629 & ~w12630;
assign w12632 = (~w12244 & ~w12245) | (~w12244 & w29809) | (~w12245 & w29809);
assign w12633 = w12631 & w12632;
assign w12634 = ~w12631 & ~w12632;
assign w12635 = ~w12633 & ~w12634;
assign w12636 = w8 & w29810;
assign w12637 = ~w8 & w29811;
assign w12638 = b_62 & w4;
assign w12639 = ~w12637 & ~w12638;
assign w12640 = ~w12636 & w12639;
assign w12641 = b_62 & ~b_63;
assign w12642 = ~b_62 & b_63;
assign w12643 = ~w12641 & ~w12642;
assign w12644 = (w6406 & w40102) | (w6406 & w40103) | (w40102 & w40103);
assign w12645 = (~w6406 & w40104) | (~w6406 & w40105) | (w40104 & w40105);
assign w12646 = ~w12644 & ~w12645;
assign w12647 = (w12640 & ~w12646) | (w12640 & w29817) | (~w12646 & w29817);
assign w12648 = (w12646 & w40106) | (w12646 & w40107) | (w40106 & w40107);
assign w12649 = (~w12646 & w40108) | (~w12646 & w40109) | (w40108 & w40109);
assign w12650 = ~w12647 & ~w12648;
assign w12651 = ~w12649 & ~w12650;
assign w12652 = w12635 & ~w12651;
assign w12653 = w12635 & ~w12652;
assign w12654 = ~w12635 & ~w12651;
assign w12655 = ~w12653 & ~w12654;
assign w12656 = (~w12261 & ~w12262) | (~w12261 & w26836) | (~w12262 & w26836);
assign w12657 = (~w12656 & w12653) | (~w12656 & w25135) | (w12653 & w25135);
assign w12658 = ~w12655 & ~w12657;
assign w12659 = ~w12656 & ~w12657;
assign w12660 = ~w12658 & ~w12659;
assign w12661 = (~w11914 & w25447) | (~w11914 & w25448) | (w25447 & w25448);
assign w12662 = ~w12660 & ~w12661;
assign w12663 = w12660 & w12661;
assign w12664 = ~w12662 & ~w12663;
assign w12665 = (~w12657 & w12661) | (~w12657 & w25136) | (w12661 & w25136);
assign w12666 = (~w12634 & ~w12635) | (~w12634 & w29818) | (~w12635 & w29818);
assign w12667 = ~w8 & w29819;
assign w12668 = b_63 & w4;
assign w12669 = ~w12667 & ~w12668;
assign w12670 = (w6406 & w40110) | (w6406 & w40111) | (w40110 & w40111);
assign w12671 = b_63 & ~w12670;
assign w12672 = (w12 & w12671) | (w12 & w29824) | (w12671 & w29824);
assign w12673 = w12669 & ~w12672;
assign w12674 = (a_2 & w12672) | (a_2 & w29825) | (w12672 & w29825);
assign w12675 = ~w12672 & w29826;
assign w12676 = ~w12673 & ~w12674;
assign w12677 = ~w12675 & ~w12676;
assign w12678 = (~w12628 & w12618) | (~w12628 & w27837) | (w12618 & w27837);
assign w12679 = (~w12618 & w40112) | (~w12618 & w40113) | (w40112 & w40113);
assign w12680 = (~w12599 & w12602) | (~w12599 & w26297) | (w12602 & w26297);
assign w12681 = b_55 & w418;
assign w12682 = w481 & w29827;
assign w12683 = b_54 & w413;
assign w12684 = ~w12682 & ~w12683;
assign w12685 = ~w12681 & w12684;
assign w12686 = (w12685 & ~w9776) | (w12685 & w29828) | (~w9776 & w29828);
assign w12687 = (w9776 & w40114) | (w9776 & w40115) | (w40114 & w40115);
assign w12688 = (~w9776 & w40116) | (~w9776 & w40117) | (w40116 & w40117);
assign w12689 = ~w12686 & ~w12687;
assign w12690 = ~w12688 & ~w12689;
assign w12691 = (~w12583 & ~w12585) | (~w12583 & w27838) | (~w12585 & w27838);
assign w12692 = b_52 & w657;
assign w12693 = w754 & w29829;
assign w12694 = b_51 & w652;
assign w12695 = ~w12693 & ~w12694;
assign w12696 = ~w12692 & w12695;
assign w12697 = (w12696 & ~w8793) | (w12696 & w26298) | (~w8793 & w26298);
assign w12698 = (w8793 & w29830) | (w8793 & w29831) | (w29830 & w29831);
assign w12699 = (~w8793 & w29832) | (~w8793 & w29833) | (w29832 & w29833);
assign w12700 = ~w12697 & ~w12698;
assign w12701 = ~w12699 & ~w12700;
assign w12702 = (~w12576 & w12579) | (~w12576 & w27781) | (w12579 & w27781);
assign w12703 = b_49 & w986;
assign w12704 = w1069 & w29834;
assign w12705 = b_48 & w981;
assign w12706 = ~w12704 & ~w12705;
assign w12707 = ~w12703 & w12706;
assign w12708 = (w12707 & ~w7859) | (w12707 & w25646) | (~w7859 & w25646);
assign w12709 = (w7859 & w25937) | (w7859 & w25938) | (w25937 & w25938);
assign w12710 = (~w7859 & w26299) | (~w7859 & w26300) | (w26299 & w26300);
assign w12711 = ~w12708 & ~w12709;
assign w12712 = ~w12710 & ~w12711;
assign w12713 = (~w12569 & w12311) | (~w12569 & w25449) | (w12311 & w25449);
assign w12714 = b_46 & w1295;
assign w12715 = w1422 & w29835;
assign w12716 = b_45 & w1290;
assign w12717 = ~w12715 & ~w12716;
assign w12718 = ~w12714 & w12717;
assign w12719 = (w12718 & ~w6974) | (w12718 & w25647) | (~w6974 & w25647);
assign w12720 = (w6974 & w25939) | (w6974 & w25940) | (w25939 & w25940);
assign w12721 = (~w6974 & w26301) | (~w6974 & w26302) | (w26301 & w26302);
assign w12722 = ~w12719 & ~w12720;
assign w12723 = ~w12721 & ~w12722;
assign w12724 = ~w12562 & ~w12566;
assign w12725 = b_34 & w3195;
assign w12726 = w3388 & w29836;
assign w12727 = b_33 & w3190;
assign w12728 = ~w12726 & ~w12727;
assign w12729 = ~w12725 & w12728;
assign w12730 = (w12729 & ~w3967) | (w12729 & w25941) | (~w3967 & w25941);
assign w12731 = (w3967 & w29837) | (w3967 & w29838) | (w29837 & w29838);
assign w12732 = (~w3967 & w29839) | (~w3967 & w29840) | (w29839 & w29840);
assign w12733 = ~w12730 & ~w12731;
assign w12734 = ~w12732 & ~w12733;
assign w12735 = b_22 & w5962;
assign w12736 = w6246 & w29841;
assign w12737 = b_21 & w5957;
assign w12738 = ~w12736 & ~w12737;
assign w12739 = ~w12735 & w12738;
assign w12740 = (w12739 & ~w1786) | (w12739 & w29842) | (~w1786 & w29842);
assign w12741 = (w1786 & w40118) | (w1786 & w40119) | (w40118 & w40119);
assign w12742 = (~w1786 & w40120) | (~w1786 & w40121) | (w40120 & w40121);
assign w12743 = ~w12740 & ~w12741;
assign w12744 = ~w12742 & ~w12743;
assign w12745 = b_16 & w7613;
assign w12746 = w7941 & w29843;
assign w12747 = b_15 & w7608;
assign w12748 = ~w12746 & ~w12747;
assign w12749 = ~w12745 & w12748;
assign w12750 = (w12749 & ~w926) | (w12749 & w29844) | (~w926 & w29844);
assign w12751 = (w926 & w40122) | (w926 & w40123) | (w40122 & w40123);
assign w12752 = (~w926 & w40124) | (~w926 & w40125) | (w40124 & w40125);
assign w12753 = ~w12750 & ~w12751;
assign w12754 = ~w12752 & ~w12753;
assign w12755 = b_10 & w9534;
assign w12756 = w9876 & w29845;
assign w12757 = b_9 & w9529;
assign w12758 = ~w12756 & ~w12757;
assign w12759 = ~w12755 & w12758;
assign w12760 = (w12759 & ~w454) | (w12759 & w29846) | (~w454 & w29846);
assign w12761 = (w454 & w40126) | (w454 & w40127) | (w40126 & w40127);
assign w12762 = (~w454 & w40128) | (~w454 & w40129) | (w40128 & w40129);
assign w12763 = ~w12760 & ~w12761;
assign w12764 = ~w12762 & ~w12763;
assign w12765 = (~w12412 & ~w12413) | (~w12412 & w27192) | (~w12413 & w27192);
assign w12766 = w12380 & w29847;
assign w12767 = b_1 & ~w12380;
assign w12768 = ~w12766 & ~w12767;
assign w12769 = b_4 & w11620;
assign w12770 = w11969 & w27250;
assign w12771 = b_3 & w11615;
assign w12772 = ~w12770 & ~w12771;
assign w12773 = ~w12769 & w12772;
assign w12774 = w84 & w11623;
assign w12775 = w12773 & ~w12774;
assign w12776 = (a_62 & w12774) | (a_62 & w27251) | (w12774 & w27251);
assign w12777 = ~w12774 & w40130;
assign w12778 = ~w12775 & ~w12776;
assign w12779 = ~w12777 & ~w12778;
assign w12780 = (~w12768 & w12778) | (~w12768 & w40131) | (w12778 & w40131);
assign w12781 = ~w12778 & w40132;
assign w12782 = ~w12779 & ~w12780;
assign w12783 = ~w12781 & ~w12782;
assign w12784 = ~w12382 & ~w12397;
assign w12785 = w12783 & w12784;
assign w12786 = ~w12783 & ~w12784;
assign w12787 = ~w12785 & ~w12786;
assign w12788 = b_7 & w10562;
assign w12789 = w10902 & w29848;
assign w12790 = b_6 & w10557;
assign w12791 = ~w12789 & ~w12790;
assign w12792 = ~w12788 & w12791;
assign w12793 = (w12792 & ~w213) | (w12792 & w29849) | (~w213 & w29849);
assign w12794 = (w213 & w40133) | (w213 & w40134) | (w40133 & w40134);
assign w12795 = (~w213 & w40135) | (~w213 & w40136) | (w40135 & w40136);
assign w12796 = ~w12793 & ~w12794;
assign w12797 = ~w12795 & ~w12796;
assign w12798 = ~w12787 & w12797;
assign w12799 = w12787 & ~w12797;
assign w12800 = ~w12798 & ~w12799;
assign w12801 = ~w12765 & w12800;
assign w12802 = w12765 & ~w12800;
assign w12803 = ~w12801 & ~w12802;
assign w12804 = ~w12764 & w12803;
assign w12805 = w12803 & ~w12804;
assign w12806 = ~w12803 & ~w12764;
assign w12807 = ~w12805 & ~w12806;
assign w12808 = (~w12417 & w12420) | (~w12417 & w27366) | (w12420 & w27366);
assign w12809 = w12807 & w12808;
assign w12810 = ~w12807 & ~w12808;
assign w12811 = ~w12809 & ~w12810;
assign w12812 = b_13 & w8526;
assign w12813 = w8886 & w29850;
assign w12814 = b_12 & w8521;
assign w12815 = ~w12813 & ~w12814;
assign w12816 = ~w12812 & w12815;
assign w12817 = (w12816 & ~w711) | (w12816 & w29851) | (~w711 & w29851);
assign w12818 = (w711 & w40137) | (w711 & w40138) | (w40137 & w40138);
assign w12819 = (~w711 & w40139) | (~w711 & w40140) | (w40139 & w40140);
assign w12820 = ~w12817 & ~w12818;
assign w12821 = ~w12819 & ~w12820;
assign w12822 = ~w12811 & w12821;
assign w12823 = w12811 & ~w12821;
assign w12824 = ~w12822 & ~w12823;
assign w12825 = (~w12435 & ~w12436) | (~w12435 & w27367) | (~w12436 & w27367);
assign w12826 = w12824 & ~w12825;
assign w12827 = ~w12824 & w12825;
assign w12828 = ~w12826 & ~w12827;
assign w12829 = ~w12754 & w12828;
assign w12830 = w12828 & ~w12829;
assign w12831 = ~w12828 & ~w12754;
assign w12832 = ~w12830 & ~w12831;
assign w12833 = ~w12440 & ~w12446;
assign w12834 = w12832 & w12833;
assign w12835 = ~w12832 & ~w12833;
assign w12836 = ~w12834 & ~w12835;
assign w12837 = b_19 & w6761;
assign w12838 = w7075 & w29852;
assign w12839 = b_18 & w6756;
assign w12840 = ~w12838 & ~w12839;
assign w12841 = ~w12837 & w12840;
assign w12842 = (w12841 & ~w1372) | (w12841 & w29853) | (~w1372 & w29853);
assign w12843 = (w1372 & w40141) | (w1372 & w40142) | (w40141 & w40142);
assign w12844 = (~w1372 & w40143) | (~w1372 & w40144) | (w40143 & w40144);
assign w12845 = ~w12842 & ~w12843;
assign w12846 = ~w12844 & ~w12845;
assign w12847 = ~w12836 & w12846;
assign w12848 = w12836 & ~w12846;
assign w12849 = ~w12847 & ~w12848;
assign w12850 = (~w12459 & w12355) | (~w12459 & w27193) | (w12355 & w27193);
assign w12851 = w12849 & ~w12850;
assign w12852 = ~w12849 & w12850;
assign w12853 = ~w12851 & ~w12852;
assign w12854 = ~w12744 & w12853;
assign w12855 = w12853 & ~w12854;
assign w12856 = ~w12853 & ~w12744;
assign w12857 = ~w12855 & ~w12856;
assign w12858 = (~w12464 & w12344) | (~w12464 & w27194) | (w12344 & w27194);
assign w12859 = w12857 & w12858;
assign w12860 = ~w12857 & ~w12858;
assign w12861 = ~w12859 & ~w12860;
assign w12862 = b_25 & w5196;
assign w12863 = w5459 & w29854;
assign w12864 = b_24 & w5191;
assign w12865 = ~w12863 & ~w12864;
assign w12866 = ~w12862 & w12865;
assign w12867 = (w12866 & ~w2108) | (w12866 & w29855) | (~w2108 & w29855);
assign w12868 = (w2108 & w40145) | (w2108 & w40146) | (w40145 & w40146);
assign w12869 = (~w2108 & w40147) | (~w2108 & w40148) | (w40147 & w40148);
assign w12870 = ~w12867 & ~w12868;
assign w12871 = ~w12869 & ~w12870;
assign w12872 = w12861 & ~w12871;
assign w12873 = w12861 & ~w12872;
assign w12874 = ~w12861 & ~w12871;
assign w12875 = ~w12873 & ~w12874;
assign w12876 = (~w12480 & w12483) | (~w12480 & w27195) | (w12483 & w27195);
assign w12877 = w12875 & w12876;
assign w12878 = ~w12875 & ~w12876;
assign w12879 = ~w12877 & ~w12878;
assign w12880 = b_28 & w4499;
assign w12881 = w4723 & w29856;
assign w12882 = b_27 & w4494;
assign w12883 = ~w12881 & ~w12882;
assign w12884 = ~w12880 & w12883;
assign w12885 = (w12884 & ~w2771) | (w12884 & w26303) | (~w2771 & w26303);
assign w12886 = (w2771 & w29857) | (w2771 & w29858) | (w29857 & w29858);
assign w12887 = (~w2771 & w29859) | (~w2771 & w29860) | (w29859 & w29860);
assign w12888 = ~w12885 & ~w12886;
assign w12889 = ~w12887 & ~w12888;
assign w12890 = w12879 & ~w12889;
assign w12891 = w12879 & ~w12890;
assign w12892 = ~w12879 & ~w12889;
assign w12893 = ~w12891 & ~w12892;
assign w12894 = (~w12498 & w12501) | (~w12498 & w27368) | (w12501 & w27368);
assign w12895 = w12893 & w12894;
assign w12896 = ~w12893 & ~w12894;
assign w12897 = ~w12895 & ~w12896;
assign w12898 = b_31 & w3803;
assign w12899 = w4027 & w29861;
assign w12900 = b_30 & w3798;
assign w12901 = ~w12899 & ~w12900;
assign w12902 = ~w12898 & w12901;
assign w12903 = (w12902 & ~w3345) | (w12902 & w25942) | (~w3345 & w25942);
assign w12904 = (w3345 & w26304) | (w3345 & w26305) | (w26304 & w26305);
assign w12905 = (~w3345 & w29862) | (~w3345 & w29863) | (w29862 & w29863);
assign w12906 = ~w12903 & ~w12904;
assign w12907 = ~w12905 & ~w12906;
assign w12908 = ~w12897 & w12907;
assign w12909 = w12897 & ~w12907;
assign w12910 = ~w12908 & ~w12909;
assign w12911 = (~w12517 & w12519) | (~w12517 & w25450) | (w12519 & w25450);
assign w12912 = w12910 & ~w12911;
assign w12913 = ~w12910 & w12911;
assign w12914 = ~w12912 & ~w12913;
assign w12915 = ~w12734 & w12914;
assign w12916 = w12914 & ~w12915;
assign w12917 = ~w12914 & ~w12734;
assign w12918 = ~w12916 & ~w12917;
assign w12919 = (~w12523 & w12526) | (~w12523 & w27555) | (w12526 & w27555);
assign w12920 = w12918 & w12919;
assign w12921 = ~w12918 & ~w12919;
assign w12922 = ~w12920 & ~w12921;
assign w12923 = b_37 & w2639;
assign w12924 = w2820 & w29864;
assign w12925 = b_36 & w2634;
assign w12926 = ~w12924 & ~w12925;
assign w12927 = ~w12923 & w12926;
assign w12928 = (w12927 & ~w4636) | (w12927 & w25648) | (~w4636 & w25648);
assign w12929 = (w4636 & w25943) | (w4636 & w25944) | (w25943 & w25944);
assign w12930 = (~w4636 & w29865) | (~w4636 & w29866) | (w29865 & w29866);
assign w12931 = ~w12928 & ~w12929;
assign w12932 = ~w12930 & ~w12931;
assign w12933 = w12922 & ~w12932;
assign w12934 = w12922 & ~w12933;
assign w12935 = ~w12922 & ~w12932;
assign w12936 = ~w12934 & ~w12935;
assign w12937 = (~w12540 & w12333) | (~w12540 & w25137) | (w12333 & w25137);
assign w12938 = w12936 & w12937;
assign w12939 = ~w12936 & ~w12937;
assign w12940 = ~w12938 & ~w12939;
assign w12941 = b_40 & w2158;
assign w12942 = w2294 & w29867;
assign w12943 = b_39 & w2153;
assign w12944 = ~w12942 & ~w12943;
assign w12945 = ~w12941 & w12944;
assign w12946 = (w12945 & ~w5363) | (w12945 & w25451) | (~w5363 & w25451);
assign w12947 = (w5363 & w25649) | (w5363 & w25650) | (w25649 & w25650);
assign w12948 = (~w5363 & w25945) | (~w5363 & w25946) | (w25945 & w25946);
assign w12949 = ~w12946 & ~w12947;
assign w12950 = ~w12948 & ~w12949;
assign w12951 = w12940 & ~w12950;
assign w12952 = w12950 & w12940;
assign w12953 = ~w12940 & ~w12950;
assign w12954 = ~w12952 & ~w12953;
assign w12955 = (~w12557 & w12332) | (~w12557 & w25138) | (w12332 & w25138);
assign w12956 = ~w12954 & ~w12955;
assign w12957 = ~w12954 & ~w12956;
assign w12958 = b_43 & w1694;
assign w12959 = w1834 & w29868;
assign w12960 = b_42 & w1689;
assign w12961 = ~w12959 & ~w12960;
assign w12962 = ~w12958 & w12961;
assign w12963 = (w12962 & ~w5888) | (w12962 & w26306) | (~w5888 & w26306);
assign w12964 = (w5888 & w29869) | (w5888 & w29870) | (w29869 & w29870);
assign w12965 = (~w5888 & w29871) | (~w5888 & w29872) | (w29871 & w29872);
assign w12966 = ~w12963 & ~w12964;
assign w12967 = ~w12965 & ~w12966;
assign w12968 = (w12967 & w12957) | (w12967 & w27768) | (w12957 & w27768);
assign w12969 = ~w12957 & w27769;
assign w12970 = ~w12968 & ~w12969;
assign w12971 = ~w12724 & ~w12970;
assign w12972 = w12724 & w12970;
assign w12973 = ~w12971 & ~w12972;
assign w12974 = ~w12723 & w12973;
assign w12975 = ~w12973 & ~w12723;
assign w12976 = w12723 & w12973;
assign w12977 = ~w12975 & ~w12976;
assign w12978 = ~w12713 & ~w12977;
assign w12979 = w12713 & w12977;
assign w12980 = ~w12978 & ~w12979;
assign w12981 = ~w12712 & w12980;
assign w12982 = ~w12980 & ~w12712;
assign w12983 = w12980 & ~w12981;
assign w12984 = ~w12982 & ~w12983;
assign w12985 = ~w12702 & ~w12984;
assign w12986 = w12702 & w12984;
assign w12987 = ~w12985 & ~w12986;
assign w12988 = ~w12701 & w12987;
assign w12989 = w12701 & ~w12987;
assign w12990 = ~w12988 & ~w12989;
assign w12991 = ~w12691 & w12990;
assign w12992 = w12691 & ~w12990;
assign w12993 = ~w12991 & ~w12992;
assign w12994 = ~w12690 & w12993;
assign w12995 = w12690 & ~w12993;
assign w12996 = ~w12994 & ~w12995;
assign w12997 = ~w12680 & w12996;
assign w12998 = w12680 & ~w12996;
assign w12999 = ~w12997 & ~w12998;
assign w13000 = b_58 & w239;
assign w13001 = w266 & w29873;
assign w13002 = b_57 & w234;
assign w13003 = ~w13001 & ~w13002;
assign w13004 = ~w13000 & w13003;
assign w13005 = (w13004 & ~w10476) | (w13004 & w29874) | (~w10476 & w29874);
assign w13006 = (w10476 & w40149) | (w10476 & w40150) | (w40149 & w40150);
assign w13007 = (~w10476 & w40151) | (~w10476 & w40152) | (w40151 & w40152);
assign w13008 = ~w13005 & ~w13006;
assign w13009 = ~w13007 & ~w13008;
assign w13010 = w12999 & ~w13009;
assign w13011 = w12999 & ~w13010;
assign w13012 = b_61 & w99;
assign w13013 = w136 & w29875;
assign w13014 = b_60 & w94;
assign w13015 = ~w13013 & ~w13014;
assign w13016 = ~w13012 & w13015;
assign w13017 = (w13016 & ~w11901) | (w13016 & w27556) | (~w11901 & w27556);
assign w13018 = (w11901 & w29876) | (w11901 & w29877) | (w29876 & w29877);
assign w13019 = (~w11901 & w29878) | (~w11901 & w29879) | (w29878 & w29879);
assign w13020 = ~w13017 & ~w13018;
assign w13021 = ~w13019 & ~w13020;
assign w13022 = (w13021 & w13011) | (w13021 & w26659) | (w13011 & w26659);
assign w13023 = ~w13011 & w26660;
assign w13024 = ~w13022 & ~w13023;
assign w13025 = ~w12679 & ~w13024;
assign w13026 = w12679 & w13024;
assign w13027 = ~w13025 & ~w13026;
assign w13028 = ~w12677 & w13027;
assign w13029 = w12677 & ~w13027;
assign w13030 = ~w13028 & ~w13029;
assign w13031 = ~w12666 & w13030;
assign w13032 = w12666 & ~w13030;
assign w13033 = ~w13031 & ~w13032;
assign w13034 = ~w12665 & w13033;
assign w13035 = w12665 & ~w13033;
assign w13036 = ~w13034 & ~w13035;
assign w13037 = b_53 & w657;
assign w13038 = w754 & w29880;
assign w13039 = b_52 & w652;
assign w13040 = ~w13038 & ~w13039;
assign w13041 = ~w13037 & w13040;
assign w13042 = (w9109 & w40153) | (w9109 & w40154) | (w40153 & w40154);
assign w13043 = a_14 & ~w13042;
assign w13044 = w13042 & a_14;
assign w13045 = ~w13042 & ~w13043;
assign w13046 = ~w13044 & ~w13045;
assign w13047 = ~w12981 & ~w12985;
assign w13048 = (~w12974 & w12977) | (~w12974 & w26307) | (w12977 & w26307);
assign w13049 = b_47 & w1295;
assign w13050 = w1422 & w29882;
assign w13051 = b_46 & w1290;
assign w13052 = ~w13050 & ~w13051;
assign w13053 = ~w13049 & w13052;
assign w13054 = (w13053 & ~w6998) | (w13053 & w25651) | (~w6998 & w25651);
assign w13055 = (w6998 & w25947) | (w6998 & w25948) | (w25947 & w25948);
assign w13056 = (~w6998 & w26308) | (~w6998 & w26309) | (w26308 & w26309);
assign w13057 = ~w13054 & ~w13055;
assign w13058 = ~w13056 & ~w13057;
assign w13059 = (~w12951 & w12954) | (~w12951 & w25949) | (w12954 & w25949);
assign w13060 = (~w12909 & w12911) | (~w12909 & w26928) | (w12911 & w26928);
assign w13061 = ~w12854 & ~w12860;
assign w13062 = ~w12848 & ~w12851;
assign w13063 = (~w12829 & w12833) | (~w12829 & w27369) | (w12833 & w27369);
assign w13064 = (~w12823 & w12825) | (~w12823 & w29883) | (w12825 & w29883);
assign w13065 = b_14 & w8526;
assign w13066 = w8886 & w29884;
assign w13067 = b_13 & w8521;
assign w13068 = ~w13066 & ~w13067;
assign w13069 = ~w13065 & w13068;
assign w13070 = (w13069 & ~w735) | (w13069 & w29885) | (~w735 & w29885);
assign w13071 = (w735 & w40155) | (w735 & w40156) | (w40155 & w40156);
assign w13072 = (~w735 & w40157) | (~w735 & w40158) | (w40157 & w40158);
assign w13073 = ~w13070 & ~w13071;
assign w13074 = ~w13072 & ~w13073;
assign w13075 = ~w12804 & ~w12810;
assign w13076 = ~w12799 & ~w12801;
assign w13077 = w12380 & w29886;
assign w13078 = b_2 & ~w12380;
assign w13079 = ~w13077 & ~w13078;
assign w13080 = b_5 & w11620;
assign w13081 = w11969 & w29887;
assign w13082 = b_4 & w11615;
assign w13083 = ~w13081 & ~w13082;
assign w13084 = ~w13080 & w13083;
assign w13085 = w129 & w11623;
assign w13086 = w13084 & ~w13085;
assign w13087 = (a_62 & w13085) | (a_62 & w29888) | (w13085 & w29888);
assign w13088 = ~w13085 & w40159;
assign w13089 = ~w13086 & ~w13087;
assign w13090 = ~w13088 & ~w13089;
assign w13091 = (~w13079 & w13089) | (~w13079 & w40160) | (w13089 & w40160);
assign w13092 = ~w13089 & w40161;
assign w13093 = ~w13090 & ~w13091;
assign w13094 = ~w13092 & ~w13093;
assign w13095 = (w12784 & w40162) | (w12784 & w40163) | (w40162 & w40163);
assign w13096 = (~w12784 & w40164) | (~w12784 & w40165) | (w40164 & w40165);
assign w13097 = ~w13095 & ~w13096;
assign w13098 = b_8 & w10562;
assign w13099 = w10902 & w29891;
assign w13100 = b_7 & w10557;
assign w13101 = ~w13099 & ~w13100;
assign w13102 = ~w13098 & w13101;
assign w13103 = ~w308 & w29892;
assign w13104 = (w13102 & ~w29892) | (w13102 & w40166) | (~w29892 & w40166);
assign w13105 = (w29892 & w40167) | (w29892 & w40168) | (w40167 & w40168);
assign w13106 = ~w13103 & w29894;
assign w13107 = ~w13104 & ~w13105;
assign w13108 = ~w13106 & ~w13107;
assign w13109 = w13097 & ~w13108;
assign w13110 = ~w13097 & w13108;
assign w13111 = (w27252 & w12801) | (w27252 & w40169) | (w12801 & w40169);
assign w13112 = ~w13076 & ~w13111;
assign w13113 = (~w13109 & w13076) | (~w13109 & w27371) | (w13076 & w27371);
assign w13114 = (w13076 & w27252) | (w13076 & w40170) | (w27252 & w40170);
assign w13115 = ~w13112 & ~w13114;
assign w13116 = b_11 & w9534;
assign w13117 = w9876 & w29895;
assign w13118 = b_10 & w9529;
assign w13119 = ~w13117 & ~w13118;
assign w13120 = ~w13116 & w13119;
assign w13121 = (w13120 & ~w530) | (w13120 & w29896) | (~w530 & w29896);
assign w13122 = (w530 & w40171) | (w530 & w40172) | (w40171 & w40172);
assign w13123 = (~w530 & w40173) | (~w530 & w40174) | (w40173 & w40174);
assign w13124 = ~w13121 & ~w13122;
assign w13125 = ~w13123 & ~w13124;
assign w13126 = w13115 & w13125;
assign w13127 = ~w13115 & ~w13125;
assign w13128 = ~w13126 & ~w13127;
assign w13129 = ~w13075 & w13128;
assign w13130 = w13075 & ~w13128;
assign w13131 = ~w13129 & ~w13130;
assign w13132 = ~w13074 & w13131;
assign w13133 = w13131 & ~w13132;
assign w13134 = ~w13131 & ~w13074;
assign w13135 = ~w13133 & ~w13134;
assign w13136 = ~w13064 & w13135;
assign w13137 = w13064 & ~w13135;
assign w13138 = ~w13136 & ~w13137;
assign w13139 = b_17 & w7613;
assign w13140 = w7941 & w29897;
assign w13141 = b_16 & w7608;
assign w13142 = ~w13140 & ~w13141;
assign w13143 = ~w13139 & w13142;
assign w13144 = (w13143 & ~w1038) | (w13143 & w29898) | (~w1038 & w29898);
assign w13145 = (w1038 & w40175) | (w1038 & w40176) | (w40175 & w40176);
assign w13146 = (~w1038 & w40177) | (~w1038 & w40178) | (w40177 & w40178);
assign w13147 = ~w13144 & ~w13145;
assign w13148 = ~w13146 & ~w13147;
assign w13149 = ~w13138 & ~w13148;
assign w13150 = w13138 & w13148;
assign w13151 = ~w13149 & ~w13150;
assign w13152 = w13063 & ~w13151;
assign w13153 = ~w13063 & w13151;
assign w13154 = ~w13152 & ~w13153;
assign w13155 = b_20 & w6761;
assign w13156 = w7075 & w29899;
assign w13157 = b_19 & w6756;
assign w13158 = ~w13156 & ~w13157;
assign w13159 = ~w13155 & w13158;
assign w13160 = (w13159 & ~w1503) | (w13159 & w29900) | (~w1503 & w29900);
assign w13161 = (w1503 & w40179) | (w1503 & w40180) | (w40179 & w40180);
assign w13162 = (~w1503 & w40181) | (~w1503 & w40182) | (w40181 & w40182);
assign w13163 = ~w13160 & ~w13161;
assign w13164 = ~w13162 & ~w13163;
assign w13165 = w13154 & ~w13164;
assign w13166 = w13154 & ~w13165;
assign w13167 = ~w13154 & ~w13164;
assign w13168 = ~w13166 & ~w13167;
assign w13169 = ~w13062 & w13168;
assign w13170 = w13062 & ~w13168;
assign w13171 = ~w13169 & ~w13170;
assign w13172 = b_23 & w5962;
assign w13173 = w6246 & w29901;
assign w13174 = b_22 & w5957;
assign w13175 = ~w13173 & ~w13174;
assign w13176 = ~w13172 & w13175;
assign w13177 = (w13176 & ~w1933) | (w13176 & w29902) | (~w1933 & w29902);
assign w13178 = (w1933 & w40183) | (w1933 & w40184) | (w40183 & w40184);
assign w13179 = (~w1933 & w40185) | (~w1933 & w40186) | (w40185 & w40186);
assign w13180 = ~w13177 & ~w13178;
assign w13181 = ~w13179 & ~w13180;
assign w13182 = ~w13171 & ~w13181;
assign w13183 = w13171 & w13181;
assign w13184 = ~w13182 & ~w13183;
assign w13185 = w13061 & ~w13184;
assign w13186 = ~w13061 & w13184;
assign w13187 = ~w13185 & ~w13186;
assign w13188 = b_26 & w5196;
assign w13189 = w5459 & w29903;
assign w13190 = b_25 & w5191;
assign w13191 = ~w13189 & ~w13190;
assign w13192 = ~w13188 & w13191;
assign w13193 = (w13192 & ~w2416) | (w13192 & w29904) | (~w2416 & w29904);
assign w13194 = (w2416 & w40187) | (w2416 & w40188) | (w40187 & w40188);
assign w13195 = (~w2416 & w40189) | (~w2416 & w40190) | (w40189 & w40190);
assign w13196 = ~w13193 & ~w13194;
assign w13197 = ~w13195 & ~w13196;
assign w13198 = w13187 & ~w13197;
assign w13199 = w13187 & ~w13198;
assign w13200 = ~w13187 & ~w13197;
assign w13201 = ~w13199 & ~w13200;
assign w13202 = ~w12872 & ~w12878;
assign w13203 = w13201 & w13202;
assign w13204 = ~w13201 & ~w13202;
assign w13205 = ~w13203 & ~w13204;
assign w13206 = b_29 & w4499;
assign w13207 = w4723 & w29905;
assign w13208 = b_28 & w4494;
assign w13209 = ~w13207 & ~w13208;
assign w13210 = ~w13206 & w13209;
assign w13211 = (w13210 & ~w2954) | (w13210 & w29906) | (~w2954 & w29906);
assign w13212 = (w2954 & w40191) | (w2954 & w40192) | (w40191 & w40192);
assign w13213 = (~w2954 & w40193) | (~w2954 & w40194) | (w40193 & w40194);
assign w13214 = ~w13211 & ~w13212;
assign w13215 = ~w13213 & ~w13214;
assign w13216 = w13205 & ~w13215;
assign w13217 = w13205 & ~w13216;
assign w13218 = ~w13205 & ~w13215;
assign w13219 = ~w13217 & ~w13218;
assign w13220 = (~w12890 & w12894) | (~w12890 & w27253) | (w12894 & w27253);
assign w13221 = w13219 & w13220;
assign w13222 = ~w13219 & ~w13220;
assign w13223 = ~w13221 & ~w13222;
assign w13224 = b_32 & w3803;
assign w13225 = w4027 & w29907;
assign w13226 = b_31 & w3798;
assign w13227 = ~w13225 & ~w13226;
assign w13228 = ~w13224 & w13227;
assign w13229 = (w13228 & ~w3545) | (w13228 & w26310) | (~w3545 & w26310);
assign w13230 = (w3545 & w29908) | (w3545 & w29909) | (w29908 & w29909);
assign w13231 = (~w3545 & w29910) | (~w3545 & w29911) | (w29910 & w29911);
assign w13232 = ~w13229 & ~w13230;
assign w13233 = ~w13231 & ~w13232;
assign w13234 = w13223 & ~w13233;
assign w13235 = ~w13223 & w13233;
assign w13236 = ~w13060 & w27196;
assign w13237 = ~w13060 & ~w13236;
assign w13238 = (~w13234 & w13060) | (~w13234 & w27254) | (w13060 & w27254);
assign w13239 = (w27254 & w27196) | (w27254 & w27372) | (w27196 & w27372);
assign w13240 = ~w13237 & ~w13239;
assign w13241 = b_35 & w3195;
assign w13242 = w3388 & w29912;
assign w13243 = b_34 & w3190;
assign w13244 = ~w13242 & ~w13243;
assign w13245 = ~w13241 & w13244;
assign w13246 = (w13245 & ~w4181) | (w13245 & w29913) | (~w4181 & w29913);
assign w13247 = (w4181 & w40195) | (w4181 & w40196) | (w40195 & w40196);
assign w13248 = (~w4181 & w40197) | (~w4181 & w40198) | (w40197 & w40198);
assign w13249 = ~w13246 & ~w13247;
assign w13250 = ~w13248 & ~w13249;
assign w13251 = ~w13240 & ~w13250;
assign w13252 = ~w13240 & ~w13251;
assign w13253 = w13240 & ~w13250;
assign w13254 = ~w13252 & ~w13253;
assign w13255 = (~w12915 & w12918) | (~w12915 & w29914) | (w12918 & w29914);
assign w13256 = w13254 & w13255;
assign w13257 = ~w13254 & ~w13255;
assign w13258 = ~w13256 & ~w13257;
assign w13259 = b_38 & w2639;
assign w13260 = w2820 & w29915;
assign w13261 = b_37 & w2634;
assign w13262 = ~w13260 & ~w13261;
assign w13263 = ~w13259 & w13262;
assign w13264 = (w13263 & ~w4658) | (w13263 & w26311) | (~w4658 & w26311);
assign w13265 = (w4658 & w29916) | (w4658 & w29917) | (w29916 & w29917);
assign w13266 = (~w4658 & w29918) | (~w4658 & w29919) | (w29918 & w29919);
assign w13267 = ~w13264 & ~w13265;
assign w13268 = ~w13266 & ~w13267;
assign w13269 = w13258 & ~w13268;
assign w13270 = w13258 & ~w13269;
assign w13271 = ~w13258 & ~w13268;
assign w13272 = (~w12933 & w12936) | (~w12933 & w27255) | (w12936 & w27255);
assign w13273 = ~w13270 & w27478;
assign w13274 = (~w13272 & w13270) | (~w13272 & w27479) | (w13270 & w27479);
assign w13275 = ~w13273 & ~w13274;
assign w13276 = b_41 & w2158;
assign w13277 = w2294 & w29920;
assign w13278 = b_40 & w2153;
assign w13279 = ~w13277 & ~w13278;
assign w13280 = ~w13276 & w13279;
assign w13281 = (w13280 & ~w5609) | (w13280 & w25950) | (~w5609 & w25950);
assign w13282 = (w5609 & w26312) | (w5609 & w26313) | (w26312 & w26313);
assign w13283 = (~w5609 & w29921) | (~w5609 & w29922) | (w29921 & w29922);
assign w13284 = ~w13281 & ~w13282;
assign w13285 = ~w13283 & ~w13284;
assign w13286 = w13275 & ~w13285;
assign w13287 = ~w13275 & w13285;
assign w13288 = ~w13059 & w26314;
assign w13289 = ~w26314 & ~w13059;
assign w13290 = (~w13286 & ~w26314) | (~w13286 & w29923) | (~w26314 & w29923);
assign w13291 = ~w13288 & w26314;
assign w13292 = ~w13289 & ~w13291;
assign w13293 = b_44 & w1694;
assign w13294 = w1834 & w29924;
assign w13295 = b_43 & w1689;
assign w13296 = ~w13294 & ~w13295;
assign w13297 = ~w13293 & w13296;
assign w13298 = (w13297 & ~w6408) | (w13297 & w25951) | (~w6408 & w25951);
assign w13299 = (w6408 & w26315) | (w6408 & w26316) | (w26315 & w26316);
assign w13300 = (~w6408 & w29925) | (~w6408 & w29926) | (w29925 & w29926);
assign w13301 = ~w13298 & ~w13299;
assign w13302 = ~w13300 & ~w13301;
assign w13303 = (~w13302 & w13291) | (~w13302 & w27770) | (w13291 & w27770);
assign w13304 = ~w13292 & ~w13303;
assign w13305 = ~w13291 & w27782;
assign w13306 = ~w13304 & ~w13305;
assign w13307 = (~w12967 & w12957) | (~w12967 & w29927) | (w12957 & w29927);
assign w13308 = (~w13307 & w12724) | (~w13307 & w27783) | (w12724 & w27783);
assign w13309 = ~w13306 & ~w13308;
assign w13310 = w13306 & w13308;
assign w13311 = ~w13309 & ~w13310;
assign w13312 = ~w13058 & w13311;
assign w13313 = ~w13311 & ~w13058;
assign w13314 = w13058 & w13311;
assign w13315 = ~w13313 & ~w13314;
assign w13316 = ~w13048 & ~w13315;
assign w13317 = ~w13315 & ~w13316;
assign w13318 = b_50 & w986;
assign w13319 = w1069 & w29928;
assign w13320 = b_49 & w981;
assign w13321 = ~w13319 & ~w13320;
assign w13322 = ~w13318 & w13321;
assign w13323 = (w13322 & ~w8162) | (w13322 & w27557) | (~w8162 & w27557);
assign w13324 = (w8162 & w29929) | (w8162 & w29930) | (w29929 & w29930);
assign w13325 = (~w8162 & w29931) | (~w8162 & w29932) | (w29931 & w29932);
assign w13326 = ~w13323 & ~w13324;
assign w13327 = ~w13325 & ~w13326;
assign w13328 = ~w13317 & w26661;
assign w13329 = (~w13327 & w13317) | (~w13327 & w26662) | (w13317 & w26662);
assign w13330 = ~w13328 & ~w13329;
assign w13331 = ~w13047 & w13330;
assign w13332 = w13047 & ~w13330;
assign w13333 = ~w13331 & ~w13332;
assign w13334 = ~w13046 & w13333;
assign w13335 = w13333 & ~w13334;
assign w13336 = ~w13333 & ~w13046;
assign w13337 = ~w13335 & ~w13336;
assign w13338 = ~w12988 & ~w12991;
assign w13339 = w13337 & w13338;
assign w13340 = ~w13337 & ~w13338;
assign w13341 = ~w13339 & ~w13340;
assign w13342 = b_56 & w418;
assign w13343 = w481 & w29933;
assign w13344 = b_55 & w413;
assign w13345 = ~w13343 & ~w13344;
assign w13346 = ~w13342 & w13345;
assign w13347 = (w13346 & ~w9798) | (w13346 & w29934) | (~w9798 & w29934);
assign w13348 = (w9798 & w40199) | (w9798 & w40200) | (w40199 & w40200);
assign w13349 = (~w9798 & w40201) | (~w9798 & w40202) | (w40201 & w40202);
assign w13350 = ~w13347 & ~w13348;
assign w13351 = ~w13349 & ~w13350;
assign w13352 = ~w13341 & w13351;
assign w13353 = w13341 & ~w13351;
assign w13354 = ~w13352 & ~w13353;
assign w13355 = b_59 & w239;
assign w13356 = w266 & w29935;
assign w13357 = b_58 & w234;
assign w13358 = ~w13356 & ~w13357;
assign w13359 = ~w13355 & w13358;
assign w13360 = (w13359 & ~w11169) | (w13359 & w29936) | (~w11169 & w29936);
assign w13361 = (w11169 & w40203) | (w11169 & w40204) | (w40203 & w40204);
assign w13362 = (~w11169 & w40205) | (~w11169 & w40206) | (w40205 & w40206);
assign w13363 = ~w13360 & ~w13361;
assign w13364 = ~w13362 & ~w13363;
assign w13365 = w13354 & ~w13364;
assign w13366 = w13354 & ~w13365;
assign w13367 = (~w12994 & w12680) | (~w12994 & w29937) | (w12680 & w29937);
assign w13368 = ~w13366 & w26317;
assign w13369 = (~w13367 & w13366) | (~w13367 & w26318) | (w13366 & w26318);
assign w13370 = ~w13368 & ~w13369;
assign w13371 = b_62 & w99;
assign w13372 = w136 & w29938;
assign w13373 = b_61 & w94;
assign w13374 = ~w13372 & ~w13373;
assign w13375 = ~w13371 & w13374;
assign w13376 = (w13375 & ~w12273) | (w13375 & w29939) | (~w12273 & w29939);
assign w13377 = (w12273 & w40207) | (w12273 & w40208) | (w40207 & w40208);
assign w13378 = (~w12273 & w40209) | (~w12273 & w40210) | (w40209 & w40210);
assign w13379 = ~w13376 & ~w13377;
assign w13380 = ~w13378 & ~w13379;
assign w13381 = w13370 & ~w13380;
assign w13382 = w13370 & ~w13381;
assign w13383 = ~w13370 & ~w13380;
assign w13384 = ~w13382 & ~w13383;
assign w13385 = (w6406 & w40211) | (w6406 & w40212) | (w40211 & w40212);
assign w13386 = ~a_2 & ~w13385;
assign w13387 = ~w8 & w29942;
assign w13388 = (a_2 & w13385) | (a_2 & w29943) | (w13385 & w29943);
assign w13389 = ~w13386 & ~w13388;
assign w13390 = (w13011 & w37620) | (w13011 & w37621) | (w37620 & w37621);
assign w13391 = (~w13011 & w37622) | (~w13011 & w37623) | (w37622 & w37623);
assign w13392 = ~w13390 & ~w13391;
assign w13393 = (w13392 & w13382) | (w13392 & w26839) | (w13382 & w26839);
assign w13394 = ~w13384 & ~w13393;
assign w13395 = ~w13382 & w27256;
assign w13396 = (~w13025 & ~w13027) | (~w13025 & w26840) | (~w13027 & w26840);
assign w13397 = ~w13394 & w26664;
assign w13398 = (~w13396 & w13394) | (~w13396 & w26665) | (w13394 & w26665);
assign w13399 = ~w13397 & ~w13398;
assign w13400 = (~w13031 & w12665) | (~w13031 & w25139) | (w12665 & w25139);
assign w13401 = w13399 & ~w13400;
assign w13402 = ~w13399 & w13400;
assign w13403 = ~w13401 & ~w13402;
assign w13404 = (~w13369 & ~w13370) | (~w13369 & w25140) | (~w13370 & w25140);
assign w13405 = b_63 & w99;
assign w13406 = w136 & w29944;
assign w13407 = b_62 & w94;
assign w13408 = ~w13406 & ~w13407;
assign w13409 = ~w13405 & w13408;
assign w13410 = (w13409 & ~w12646) | (w13409 & w29945) | (~w12646 & w29945);
assign w13411 = (w12646 & w40213) | (w12646 & w40214) | (w40213 & w40214);
assign w13412 = (~w12646 & w40215) | (~w12646 & w40216) | (w40215 & w40216);
assign w13413 = ~w13410 & ~w13411;
assign w13414 = ~w13412 & ~w13413;
assign w13415 = (w13370 & w37660) | (w13370 & w37661) | (w37660 & w37661);
assign w13416 = ~w13404 & ~w13415;
assign w13417 = (~w13370 & w38054) | (~w13370 & w38055) | (w38054 & w38055);
assign w13418 = ~w13416 & ~w13417;
assign w13419 = b_57 & w418;
assign w13420 = w481 & w29946;
assign w13421 = b_56 & w413;
assign w13422 = ~w13420 & ~w13421;
assign w13423 = ~w13419 & w13422;
assign w13424 = (w13423 & ~w10452) | (w13423 & w29947) | (~w10452 & w29947);
assign w13425 = (w10452 & w40217) | (w10452 & w40218) | (w40217 & w40218);
assign w13426 = (~w10452 & w40219) | (~w10452 & w40220) | (w40219 & w40220);
assign w13427 = ~w13424 & ~w13425;
assign w13428 = ~w13426 & ~w13427;
assign w13429 = (~w13334 & w13337) | (~w13334 & w26319) | (w13337 & w26319);
assign w13430 = (w13337 & w37662) | (w13337 & w37663) | (w37662 & w37663);
assign w13431 = (~w13337 & w37664) | (~w13337 & w37665) | (w37664 & w37665);
assign w13432 = ~w13430 & ~w13431;
assign w13433 = b_51 & w986;
assign w13434 = w1069 & w29948;
assign w13435 = b_50 & w981;
assign w13436 = ~w13434 & ~w13435;
assign w13437 = ~w13433 & w13436;
assign w13438 = (w13437 & ~w8186) | (w13437 & w26320) | (~w8186 & w26320);
assign w13439 = (w8186 & w27558) | (w8186 & w27559) | (w27558 & w27559);
assign w13440 = (~w8186 & w29949) | (~w8186 & w29950) | (w29949 & w29950);
assign w13441 = ~w13438 & ~w13439;
assign w13442 = ~w13440 & ~w13441;
assign w13443 = (w27560 & w27771) | (w27560 & w27772) | (w27771 & w27772);
assign w13444 = (~w27560 & w27773) | (~w27560 & w27774) | (w27773 & w27774);
assign w13445 = ~w13443 & ~w13444;
assign w13446 = b_48 & w1295;
assign w13447 = w1422 & w29951;
assign w13448 = b_47 & w1290;
assign w13449 = ~w13447 & ~w13448;
assign w13450 = ~w13446 & w13449;
assign w13451 = (w13450 & ~w7284) | (w13450 & w27561) | (~w7284 & w27561);
assign w13452 = (w7284 & w29952) | (w7284 & w29953) | (w29952 & w29953);
assign w13453 = (~w7284 & w29954) | (~w7284 & w29955) | (w29954 & w29955);
assign w13454 = ~w13451 & ~w13452;
assign w13455 = ~w13453 & ~w13454;
assign w13456 = (~w13303 & w13306) | (~w13303 & w29956) | (w13306 & w29956);
assign w13457 = w13455 & w13456;
assign w13458 = ~w13455 & ~w13456;
assign w13459 = ~w13457 & ~w13458;
assign w13460 = b_45 & w1694;
assign w13461 = w1834 & w29957;
assign w13462 = b_44 & w1689;
assign w13463 = ~w13461 & ~w13462;
assign w13464 = ~w13460 & w13463;
assign w13465 = (w13464 & ~w6682) | (w13464 & w26666) | (~w6682 & w26666);
assign w13466 = (w6682 & w27480) | (w6682 & w27481) | (w27480 & w27481);
assign w13467 = (~w6682 & w29958) | (~w6682 & w29959) | (w29958 & w29959);
assign w13468 = ~w13465 & ~w13466;
assign w13469 = ~w13467 & ~w13468;
assign w13470 = ~w13290 & w13469;
assign w13471 = w13290 & ~w13469;
assign w13472 = ~w13470 & ~w13471;
assign w13473 = b_42 & w2158;
assign w13474 = w2294 & w29960;
assign w13475 = b_41 & w2153;
assign w13476 = ~w13474 & ~w13475;
assign w13477 = ~w13473 & w13476;
assign w13478 = (w13477 & ~w5864) | (w13477 & w29961) | (~w5864 & w29961);
assign w13479 = (w5864 & w40221) | (w5864 & w40222) | (w40221 & w40222);
assign w13480 = (~w5864 & w40223) | (~w5864 & w40224) | (w40223 & w40224);
assign w13481 = ~w13478 & ~w13479;
assign w13482 = ~w13480 & ~w13481;
assign w13483 = (~w27479 & w29962) | (~w27479 & w29963) | (w29962 & w29963);
assign w13484 = w13482 & w13483;
assign w13485 = ~w13482 & ~w13483;
assign w13486 = ~w13484 & ~w13485;
assign w13487 = (~w13251 & w13254) | (~w13251 & w29964) | (w13254 & w29964);
assign w13488 = b_39 & w2639;
assign w13489 = w2820 & w29965;
assign w13490 = b_38 & w2634;
assign w13491 = ~w13489 & ~w13490;
assign w13492 = ~w13488 & w13491;
assign w13493 = w13491 & w29966;
assign w13494 = (~w4888 & w40225) | (~w4888 & w40226) | (w40225 & w40226);
assign w13495 = (w4888 & w29968) | (w4888 & w29969) | (w29968 & w29969);
assign w13496 = ~w13494 & ~w13495;
assign w13497 = ~w13487 & ~w13496;
assign w13498 = w13487 & w13496;
assign w13499 = ~w13497 & ~w13498;
assign w13500 = b_33 & w3803;
assign w13501 = w4027 & w29970;
assign w13502 = b_32 & w3798;
assign w13503 = ~w13501 & ~w13502;
assign w13504 = ~w13500 & w13503;
assign w13505 = (w13504 & ~w3744) | (w13504 & w29971) | (~w3744 & w29971);
assign w13506 = (w3744 & w40227) | (w3744 & w40228) | (w40227 & w40228);
assign w13507 = (~w3744 & w40229) | (~w3744 & w40230) | (w40229 & w40230);
assign w13508 = ~w13505 & ~w13506;
assign w13509 = ~w13507 & ~w13508;
assign w13510 = b_24 & w5962;
assign w13511 = w6246 & w29972;
assign w13512 = b_23 & w5957;
assign w13513 = ~w13511 & ~w13512;
assign w13514 = ~w13510 & w13513;
assign w13515 = (w13514 & ~w2083) | (w13514 & w29973) | (~w2083 & w29973);
assign w13516 = (w2083 & w40231) | (w2083 & w40232) | (w40231 & w40232);
assign w13517 = (~w2083 & w40233) | (~w2083 & w40234) | (w40233 & w40234);
assign w13518 = ~w13515 & ~w13516;
assign w13519 = ~w13517 & ~w13518;
assign w13520 = b_15 & w8526;
assign w13521 = w8886 & w29974;
assign w13522 = b_14 & w8521;
assign w13523 = ~w13521 & ~w13522;
assign w13524 = ~w13520 & w13523;
assign w13525 = (w13524 & ~w827) | (w13524 & w29975) | (~w827 & w29975);
assign w13526 = (w827 & w40235) | (w827 & w40236) | (w40235 & w40236);
assign w13527 = (~w827 & w40237) | (~w827 & w40238) | (w40237 & w40238);
assign w13528 = ~w13525 & ~w13526;
assign w13529 = ~w13527 & ~w13528;
assign w13530 = w12380 & w29976;
assign w13531 = b_3 & ~w12380;
assign w13532 = ~w13530 & ~w13531;
assign w13533 = a_2 & ~w13532;
assign w13534 = ~a_2 & w13532;
assign w13535 = ~w13533 & ~w13534;
assign w13536 = b_6 & w11620;
assign w13537 = w11969 & w29977;
assign w13538 = b_5 & w11615;
assign w13539 = ~w13537 & ~w13538;
assign w13540 = ~w13536 & w13539;
assign w13541 = w13539 & w29978;
assign w13542 = (~w13541 & w190) | (~w13541 & w29979) | (w190 & w29979);
assign w13543 = a_62 & ~w13542;
assign w13544 = ~a_62 & w13542;
assign w13545 = ~w13543 & ~w13544;
assign w13546 = w13535 & ~w13545;
assign w13547 = ~w13535 & w13545;
assign w13548 = ~w13546 & ~w13547;
assign w13549 = (w13548 & w13096) | (w13548 & w29980) | (w13096 & w29980);
assign w13550 = ~w13096 & w29981;
assign w13551 = ~w13549 & ~w13550;
assign w13552 = b_9 & w10562;
assign w13553 = w10902 & w29982;
assign w13554 = b_8 & w10557;
assign w13555 = ~w13553 & ~w13554;
assign w13556 = ~w13552 & w13555;
assign w13557 = (w13556 & ~w371) | (w13556 & w29983) | (~w371 & w29983);
assign w13558 = (w371 & w40239) | (w371 & w40240) | (w40239 & w40240);
assign w13559 = (~w371 & w40241) | (~w371 & w40242) | (w40241 & w40242);
assign w13560 = ~w13557 & ~w13558;
assign w13561 = ~w13559 & ~w13560;
assign w13562 = w13551 & ~w13561;
assign w13563 = w13551 & ~w13562;
assign w13564 = ~w13551 & ~w13561;
assign w13565 = ~w13563 & ~w13564;
assign w13566 = ~w13113 & w13565;
assign w13567 = w13113 & ~w13565;
assign w13568 = ~w13566 & ~w13567;
assign w13569 = b_12 & w9534;
assign w13570 = w9876 & w29984;
assign w13571 = b_11 & w9529;
assign w13572 = ~w13570 & ~w13571;
assign w13573 = ~w13569 & w13572;
assign w13574 = (w13573 & ~w552) | (w13573 & w29985) | (~w552 & w29985);
assign w13575 = (w552 & w40243) | (w552 & w40244) | (w40243 & w40244);
assign w13576 = (~w552 & w40245) | (~w552 & w40246) | (w40245 & w40246);
assign w13577 = ~w13574 & ~w13575;
assign w13578 = ~w13576 & ~w13577;
assign w13579 = w13568 & w13578;
assign w13580 = ~w13568 & ~w13578;
assign w13581 = ~w13579 & ~w13580;
assign w13582 = (w13581 & w13129) | (w13581 & w29986) | (w13129 & w29986);
assign w13583 = ~w13129 & w29987;
assign w13584 = ~w13582 & ~w13583;
assign w13585 = ~w13529 & w13584;
assign w13586 = w13584 & ~w13585;
assign w13587 = ~w13584 & ~w13529;
assign w13588 = ~w13586 & ~w13587;
assign w13589 = (~w13132 & w13135) | (~w13132 & w29988) | (w13135 & w29988);
assign w13590 = w13588 & w13589;
assign w13591 = ~w13588 & ~w13589;
assign w13592 = ~w13590 & ~w13591;
assign w13593 = b_18 & w7613;
assign w13594 = w7941 & w29989;
assign w13595 = b_17 & w7608;
assign w13596 = ~w13594 & ~w13595;
assign w13597 = ~w13593 & w13596;
assign w13598 = (w13597 & ~w1238) | (w13597 & w29990) | (~w1238 & w29990);
assign w13599 = (w1238 & w40247) | (w1238 & w40248) | (w40247 & w40248);
assign w13600 = (~w1238 & w40249) | (~w1238 & w40250) | (w40249 & w40250);
assign w13601 = ~w13598 & ~w13599;
assign w13602 = ~w13600 & ~w13601;
assign w13603 = w13592 & ~w13602;
assign w13604 = w13592 & ~w13603;
assign w13605 = ~w13592 & ~w13602;
assign w13606 = ~w13604 & ~w13605;
assign w13607 = (~w13149 & w13063) | (~w13149 & w29991) | (w13063 & w29991);
assign w13608 = w13606 & w13607;
assign w13609 = ~w13606 & ~w13607;
assign w13610 = ~w13608 & ~w13609;
assign w13611 = b_21 & w6761;
assign w13612 = w7075 & w29992;
assign w13613 = b_20 & w6756;
assign w13614 = ~w13612 & ~w13613;
assign w13615 = ~w13611 & w13614;
assign w13616 = (w13615 & ~w1634) | (w13615 & w29993) | (~w1634 & w29993);
assign w13617 = (w1634 & w40251) | (w1634 & w40252) | (w40251 & w40252);
assign w13618 = (~w1634 & w40253) | (~w1634 & w40254) | (w40253 & w40254);
assign w13619 = ~w13616 & ~w13617;
assign w13620 = ~w13618 & ~w13619;
assign w13621 = ~w13610 & w13620;
assign w13622 = w13610 & ~w13620;
assign w13623 = ~w13621 & ~w13622;
assign w13624 = (~w13165 & w13168) | (~w13165 & w29994) | (w13168 & w29994);
assign w13625 = w13623 & ~w13624;
assign w13626 = ~w13623 & w13624;
assign w13627 = ~w13625 & ~w13626;
assign w13628 = ~w13519 & w13627;
assign w13629 = w13627 & ~w13628;
assign w13630 = ~w13627 & ~w13519;
assign w13631 = ~w13629 & ~w13630;
assign w13632 = (~w13182 & w13061) | (~w13182 & w40255) | (w13061 & w40255);
assign w13633 = w13631 & w13632;
assign w13634 = ~w13631 & ~w13632;
assign w13635 = ~w13633 & ~w13634;
assign w13636 = b_27 & w5196;
assign w13637 = w5459 & w29995;
assign w13638 = b_26 & w5191;
assign w13639 = ~w13637 & ~w13638;
assign w13640 = ~w13636 & w13639;
assign w13641 = (w13640 & ~w2582) | (w13640 & w29996) | (~w2582 & w29996);
assign w13642 = (w2582 & w40256) | (w2582 & w40257) | (w40256 & w40257);
assign w13643 = (~w2582 & w40258) | (~w2582 & w40259) | (w40258 & w40259);
assign w13644 = ~w13641 & ~w13642;
assign w13645 = ~w13643 & ~w13644;
assign w13646 = w13635 & ~w13645;
assign w13647 = w13635 & ~w13646;
assign w13648 = ~w13635 & ~w13645;
assign w13649 = ~w13647 & ~w13648;
assign w13650 = ~w13198 & ~w13204;
assign w13651 = w13649 & w13650;
assign w13652 = ~w13649 & ~w13650;
assign w13653 = ~w13651 & ~w13652;
assign w13654 = b_30 & w4499;
assign w13655 = w4723 & w29997;
assign w13656 = b_29 & w4494;
assign w13657 = ~w13655 & ~w13656;
assign w13658 = ~w13654 & w13657;
assign w13659 = (w13658 & ~w3138) | (w13658 & w29998) | (~w3138 & w29998);
assign w13660 = (w3138 & w40260) | (w3138 & w40261) | (w40260 & w40261);
assign w13661 = (~w3138 & w40262) | (~w3138 & w40263) | (w40262 & w40263);
assign w13662 = ~w13659 & ~w13660;
assign w13663 = ~w13661 & ~w13662;
assign w13664 = ~w13653 & w13663;
assign w13665 = w13653 & ~w13663;
assign w13666 = ~w13664 & ~w13665;
assign w13667 = (~w13216 & w13219) | (~w13216 & w29999) | (w13219 & w29999);
assign w13668 = w13666 & ~w13667;
assign w13669 = ~w13666 & w13667;
assign w13670 = ~w13668 & ~w13669;
assign w13671 = ~w13509 & w13670;
assign w13672 = w13670 & ~w13671;
assign w13673 = ~w13670 & ~w13509;
assign w13674 = ~w13672 & ~w13673;
assign w13675 = b_36 & w3195;
assign w13676 = w3388 & w30000;
assign w13677 = b_35 & w3190;
assign w13678 = ~w13676 & ~w13677;
assign w13679 = ~w13675 & w13678;
assign w13680 = w13678 & w30001;
assign w13681 = (~w4395 & w40264) | (~w4395 & w40265) | (w40264 & w40265);
assign w13682 = (w4395 & w30003) | (w4395 & w30004) | (w30003 & w30004);
assign w13683 = ~w13681 & ~w13682;
assign w13684 = (~w27254 & w30005) | (~w27254 & w30006) | (w30005 & w30006);
assign w13685 = ~w13238 & ~w13684;
assign w13686 = ~w13683 & ~w13684;
assign w13687 = ~w13685 & ~w13686;
assign w13688 = ~w13674 & ~w13687;
assign w13689 = w13687 & ~w13674;
assign w13690 = ~w13687 & ~w13688;
assign w13691 = ~w13689 & ~w13690;
assign w13692 = w13499 & ~w13691;
assign w13693 = w13499 & ~w13692;
assign w13694 = ~w13499 & ~w13691;
assign w13695 = ~w13693 & ~w13694;
assign w13696 = w13486 & ~w13695;
assign w13697 = ~w13486 & w13695;
assign w13698 = ~w13472 & ~w13697;
assign w13699 = ~w13472 & w30007;
assign w13700 = ~w13472 & ~w13699;
assign w13701 = w30007 & w13472;
assign w13702 = ~w13700 & ~w13701;
assign w13703 = w13459 & ~w13702;
assign w13704 = ~w13459 & w13702;
assign w13705 = w13445 & w27784;
assign w13706 = w13445 & ~w13705;
assign w13707 = w27784 & ~w13445;
assign w13708 = ~w13706 & ~w13707;
assign w13709 = (~w13329 & w13047) | (~w13329 & w26667) | (w13047 & w26667);
assign w13710 = b_54 & w657;
assign w13711 = w754 & w30008;
assign w13712 = b_53 & w652;
assign w13713 = ~w13711 & ~w13712;
assign w13714 = ~w13710 & w13713;
assign w13715 = w13713 & w30009;
assign w13716 = (~w9134 & w30010) | (~w9134 & w30011) | (w30010 & w30011);
assign w13717 = (w9134 & w30012) | (w9134 & w30013) | (w30012 & w30013);
assign w13718 = ~w13716 & ~w13717;
assign w13719 = (~w13047 & w27482) | (~w13047 & w27483) | (w27482 & w27483);
assign w13720 = ~w13709 & ~w13719;
assign w13721 = (~w27483 & w27563) | (~w27483 & w27564) | (w27563 & w27564);
assign w13722 = ~w13720 & ~w13721;
assign w13723 = (~w13708 & w13720) | (~w13708 & w30014) | (w13720 & w30014);
assign w13724 = ~w13708 & ~w13723;
assign w13725 = ~w13722 & ~w13723;
assign w13726 = ~w13724 & ~w13725;
assign w13727 = w13432 & ~w13726;
assign w13728 = w13432 & ~w13727;
assign w13729 = ~w13432 & ~w13726;
assign w13730 = ~w13728 & ~w13729;
assign w13731 = b_60 & w239;
assign w13732 = w266 & w30015;
assign w13733 = b_59 & w234;
assign w13734 = ~w13732 & ~w13733;
assign w13735 = ~w13731 & w13734;
assign w13736 = (w13735 & ~w11196) | (w13735 & w30016) | (~w11196 & w30016);
assign w13737 = (w11196 & w40266) | (w11196 & w40267) | (w40266 & w40267);
assign w13738 = (~w11196 & w40268) | (~w11196 & w40269) | (w40268 & w40269);
assign w13739 = ~w13736 & ~w13737;
assign w13740 = ~w13738 & ~w13739;
assign w13741 = (~w13353 & ~w13354) | (~w13353 & w26321) | (~w13354 & w26321);
assign w13742 = (w13354 & w37666) | (w13354 & w37667) | (w37666 & w37667);
assign w13743 = (~w13354 & w37668) | (~w13354 & w37669) | (w37668 & w37669);
assign w13744 = ~w13741 & ~w13742;
assign w13745 = ~w13743 & ~w13744;
assign w13746 = (~w13730 & w13744) | (~w13730 & w26322) | (w13744 & w26322);
assign w13747 = ~w13730 & ~w13746;
assign w13748 = ~w13745 & ~w13746;
assign w13749 = ~w13747 & ~w13748;
assign w13750 = (~w13749 & w13416) | (~w13749 & w26668) | (w13416 & w26668);
assign w13751 = ~w13418 & ~w13750;
assign w13752 = ~w13416 & w26669;
assign w13753 = (~w13382 & w38056) | (~w13382 & w38057) | (w38056 & w38057);
assign w13754 = ~w13751 & w26323;
assign w13755 = (~w13753 & w13751) | (~w13753 & w26324) | (w13751 & w26324);
assign w13756 = ~w13754 & ~w13755;
assign w13757 = (w12665 & w27785) | (w12665 & w27786) | (w27785 & w27786);
assign w13758 = (~w27786 & w30017) | (~w27786 & w30018) | (w30017 & w30018);
assign w13759 = (w27786 & w30019) | (w27786 & w30020) | (w30019 & w30020);
assign w13760 = ~w13758 & ~w13759;
assign w13761 = (w27786 & w38058) | (w27786 & w38059) | (w38058 & w38059);
assign w13762 = (~w26668 & w27787) | (~w26668 & w27788) | (w27787 & w27788);
assign w13763 = b_55 & w657;
assign w13764 = w754 & w30021;
assign w13765 = b_54 & w652;
assign w13766 = ~w13764 & ~w13765;
assign w13767 = ~w13763 & w13766;
assign w13768 = (w13767 & ~w9776) | (w13767 & w26325) | (~w9776 & w26325);
assign w13769 = (w9776 & w30022) | (w9776 & w30023) | (w30022 & w30023);
assign w13770 = (~w9776 & w30024) | (~w9776 & w30025) | (w30024 & w30025);
assign w13771 = ~w13768 & ~w13769;
assign w13772 = ~w13770 & ~w13771;
assign w13773 = (~w13444 & ~w13445) | (~w13444 & w27789) | (~w13445 & w27789);
assign w13774 = w13772 & w13773;
assign w13775 = ~w13772 & ~w13773;
assign w13776 = ~w13774 & ~w13775;
assign w13777 = b_49 & w1295;
assign w13778 = w1422 & w30026;
assign w13779 = b_48 & w1290;
assign w13780 = ~w13778 & ~w13779;
assign w13781 = ~w13777 & w13780;
assign w13782 = (w13781 & ~w7859) | (w13781 & w25952) | (~w7859 & w25952);
assign w13783 = (w7859 & w26326) | (w7859 & w26327) | (w26326 & w26327);
assign w13784 = (~w7859 & w27484) | (~w7859 & w27485) | (w27484 & w27485);
assign w13785 = ~w13782 & ~w13783;
assign w13786 = ~w13784 & ~w13785;
assign w13787 = (~w13698 & w30027) | (~w13698 & w30028) | (w30027 & w30028);
assign w13788 = (w13698 & w30029) | (w13698 & w30030) | (w30029 & w30030);
assign w13789 = ~w13787 & ~w13788;
assign w13790 = b_43 & w2158;
assign w13791 = w2294 & w30031;
assign w13792 = b_42 & w2153;
assign w13793 = ~w13791 & ~w13792;
assign w13794 = ~w13790 & w13793;
assign w13795 = (w13794 & ~w5888) | (w13794 & w27565) | (~w5888 & w27565);
assign w13796 = (w5888 & w30032) | (w5888 & w30033) | (w30032 & w30033);
assign w13797 = (~w5888 & w30034) | (~w5888 & w30035) | (w30034 & w30035);
assign w13798 = ~w13795 & ~w13796;
assign w13799 = ~w13797 & ~w13798;
assign w13800 = (~w13497 & ~w13499) | (~w13497 & w30036) | (~w13499 & w30036);
assign w13801 = w13799 & w13800;
assign w13802 = ~w13799 & ~w13800;
assign w13803 = ~w13801 & ~w13802;
assign w13804 = (~w13668 & ~w13670) | (~w13668 & w30037) | (~w13670 & w30037);
assign w13805 = b_37 & w3195;
assign w13806 = w3388 & w30038;
assign w13807 = b_36 & w3190;
assign w13808 = ~w13806 & ~w13807;
assign w13809 = ~w13805 & w13808;
assign w13810 = w13808 & w30039;
assign w13811 = (~w4636 & w40270) | (~w4636 & w40271) | (w40270 & w40271);
assign w13812 = (w4636 & w30041) | (w4636 & w30042) | (w30041 & w30042);
assign w13813 = ~w13811 & ~w13812;
assign w13814 = ~w13804 & ~w13813;
assign w13815 = w13804 & w13813;
assign w13816 = ~w13814 & ~w13815;
assign w13817 = b_34 & w3803;
assign w13818 = w4027 & w30043;
assign w13819 = b_33 & w3798;
assign w13820 = ~w13818 & ~w13819;
assign w13821 = ~w13817 & w13820;
assign w13822 = (w13821 & ~w3967) | (w13821 & w30044) | (~w3967 & w30044);
assign w13823 = (w3967 & w40272) | (w3967 & w40273) | (w40272 & w40273);
assign w13824 = (~w3967 & w40274) | (~w3967 & w40275) | (w40274 & w40275);
assign w13825 = ~w13822 & ~w13823;
assign w13826 = ~w13824 & ~w13825;
assign w13827 = (~w13652 & ~w13653) | (~w13652 & w30045) | (~w13653 & w30045);
assign w13828 = b_16 & w8526;
assign w13829 = w8886 & w30046;
assign w13830 = b_15 & w8521;
assign w13831 = ~w13829 & ~w13830;
assign w13832 = ~w13828 & w13831;
assign w13833 = (w13832 & ~w926) | (w13832 & w30047) | (~w926 & w30047);
assign w13834 = (w926 & w40276) | (w926 & w40277) | (w40276 & w40277);
assign w13835 = (~w926 & w40278) | (~w926 & w40279) | (w40278 & w40279);
assign w13836 = ~w13833 & ~w13834;
assign w13837 = ~w13835 & ~w13836;
assign w13838 = b_7 & w11620;
assign w13839 = w11969 & w30048;
assign w13840 = b_6 & w11615;
assign w13841 = ~w13839 & ~w13840;
assign w13842 = ~w13838 & w13841;
assign w13843 = (w13842 & ~w213) | (w13842 & w30049) | (~w213 & w30049);
assign w13844 = (w213 & w40280) | (w213 & w40281) | (w40280 & w40281);
assign w13845 = (~w213 & w40282) | (~w213 & w40283) | (w40282 & w40283);
assign w13846 = ~w13843 & ~w13844;
assign w13847 = ~w13845 & ~w13846;
assign w13848 = w12380 & w30050;
assign w13849 = b_4 & ~w12380;
assign w13850 = ~w13848 & ~w13849;
assign w13851 = a_2 & ~w13850;
assign w13852 = w13850 & a_2;
assign w13853 = ~w13850 & ~w13851;
assign w13854 = ~w13852 & ~w13853;
assign w13855 = (~w13854 & w13846) | (~w13854 & w30051) | (w13846 & w30051);
assign w13856 = ~w13847 & ~w13855;
assign w13857 = ~w13854 & ~w13855;
assign w13858 = ~w13856 & ~w13857;
assign w13859 = (~w13533 & w13545) | (~w13533 & w30052) | (w13545 & w30052);
assign w13860 = w13858 & w13859;
assign w13861 = ~w13858 & ~w13859;
assign w13862 = ~w13860 & ~w13861;
assign w13863 = b_10 & w10562;
assign w13864 = w10902 & w30053;
assign w13865 = b_9 & w10557;
assign w13866 = ~w13864 & ~w13865;
assign w13867 = ~w13863 & w13866;
assign w13868 = (w13867 & ~w454) | (w13867 & w30054) | (~w454 & w30054);
assign w13869 = (w454 & w40284) | (w454 & w40285) | (w40284 & w40285);
assign w13870 = (~w454 & w40286) | (~w454 & w40287) | (w40286 & w40287);
assign w13871 = ~w13868 & ~w13869;
assign w13872 = ~w13870 & ~w13871;
assign w13873 = w13862 & ~w13872;
assign w13874 = w13862 & ~w13873;
assign w13875 = ~w13862 & ~w13872;
assign w13876 = ~w13874 & ~w13875;
assign w13877 = (~w13549 & ~w13551) | (~w13549 & w30055) | (~w13551 & w30055);
assign w13878 = w13876 & w13877;
assign w13879 = ~w13876 & ~w13877;
assign w13880 = ~w13878 & ~w13879;
assign w13881 = b_13 & w9534;
assign w13882 = w9876 & w30056;
assign w13883 = b_12 & w9529;
assign w13884 = ~w13882 & ~w13883;
assign w13885 = ~w13881 & w13884;
assign w13886 = (w13885 & ~w711) | (w13885 & w30057) | (~w711 & w30057);
assign w13887 = (w711 & w40288) | (w711 & w40289) | (w40288 & w40289);
assign w13888 = (~w711 & w40290) | (~w711 & w40291) | (w40290 & w40291);
assign w13889 = ~w13886 & ~w13887;
assign w13890 = ~w13888 & ~w13889;
assign w13891 = ~w13880 & w13890;
assign w13892 = w13880 & ~w13890;
assign w13893 = ~w13891 & ~w13892;
assign w13894 = ~w13113 & ~w13565;
assign w13895 = (~w13894 & w13568) | (~w13894 & w30058) | (w13568 & w30058);
assign w13896 = w13893 & ~w13895;
assign w13897 = ~w13893 & w13895;
assign w13898 = ~w13896 & ~w13897;
assign w13899 = ~w13837 & w13898;
assign w13900 = w13898 & ~w13899;
assign w13901 = ~w13898 & ~w13837;
assign w13902 = ~w13900 & ~w13901;
assign w13903 = (~w13582 & ~w13584) | (~w13582 & w30059) | (~w13584 & w30059);
assign w13904 = w13902 & w13903;
assign w13905 = ~w13902 & ~w13903;
assign w13906 = ~w13904 & ~w13905;
assign w13907 = b_19 & w7613;
assign w13908 = w7941 & w30060;
assign w13909 = b_18 & w7608;
assign w13910 = ~w13908 & ~w13909;
assign w13911 = ~w13907 & w13910;
assign w13912 = (w13911 & ~w1372) | (w13911 & w30061) | (~w1372 & w30061);
assign w13913 = (w1372 & w40292) | (w1372 & w40293) | (w40292 & w40293);
assign w13914 = (~w1372 & w40294) | (~w1372 & w40295) | (w40294 & w40295);
assign w13915 = ~w13912 & ~w13913;
assign w13916 = ~w13914 & ~w13915;
assign w13917 = w13906 & ~w13916;
assign w13918 = w13906 & ~w13917;
assign w13919 = ~w13906 & ~w13916;
assign w13920 = ~w13918 & ~w13919;
assign w13921 = (~w13591 & ~w13592) | (~w13591 & w30062) | (~w13592 & w30062);
assign w13922 = w13920 & w13921;
assign w13923 = ~w13920 & ~w13921;
assign w13924 = ~w13922 & ~w13923;
assign w13925 = b_22 & w6761;
assign w13926 = w7075 & w30063;
assign w13927 = b_21 & w6756;
assign w13928 = ~w13926 & ~w13927;
assign w13929 = ~w13925 & w13928;
assign w13930 = (w13929 & ~w1786) | (w13929 & w30064) | (~w1786 & w30064);
assign w13931 = (w1786 & w40296) | (w1786 & w40297) | (w40296 & w40297);
assign w13932 = (~w1786 & w40298) | (~w1786 & w40299) | (w40298 & w40299);
assign w13933 = ~w13930 & ~w13931;
assign w13934 = ~w13932 & ~w13933;
assign w13935 = w13924 & ~w13934;
assign w13936 = w13924 & ~w13935;
assign w13937 = ~w13924 & ~w13934;
assign w13938 = ~w13936 & ~w13937;
assign w13939 = (~w13609 & ~w13610) | (~w13609 & w30065) | (~w13610 & w30065);
assign w13940 = ~w13938 & ~w13939;
assign w13941 = ~w13938 & ~w13940;
assign w13942 = ~w13939 & ~w13940;
assign w13943 = ~w13941 & ~w13942;
assign w13944 = b_25 & w5962;
assign w13945 = w6246 & w30066;
assign w13946 = b_24 & w5957;
assign w13947 = ~w13945 & ~w13946;
assign w13948 = ~w13944 & w13947;
assign w13949 = (w13948 & ~w2108) | (w13948 & w30067) | (~w2108 & w30067);
assign w13950 = (w2108 & w40300) | (w2108 & w40301) | (w40300 & w40301);
assign w13951 = (~w2108 & w40302) | (~w2108 & w40303) | (w40302 & w40303);
assign w13952 = ~w13949 & ~w13950;
assign w13953 = ~w13951 & ~w13952;
assign w13954 = ~w13943 & ~w13953;
assign w13955 = ~w13943 & ~w13954;
assign w13956 = w13943 & ~w13953;
assign w13957 = ~w13955 & ~w13956;
assign w13958 = (~w13625 & ~w13627) | (~w13625 & w30068) | (~w13627 & w30068);
assign w13959 = ~w13955 & w40304;
assign w13960 = (~w13958 & w13955) | (~w13958 & w40305) | (w13955 & w40305);
assign w13961 = ~w13959 & ~w13960;
assign w13962 = b_28 & w5196;
assign w13963 = w5459 & w30069;
assign w13964 = b_27 & w5191;
assign w13965 = ~w13963 & ~w13964;
assign w13966 = ~w13962 & w13965;
assign w13967 = (w13966 & ~w2771) | (w13966 & w30070) | (~w2771 & w30070);
assign w13968 = (w2771 & w40306) | (w2771 & w40307) | (w40306 & w40307);
assign w13969 = (~w2771 & w40308) | (~w2771 & w40309) | (w40308 & w40309);
assign w13970 = ~w13967 & ~w13968;
assign w13971 = ~w13969 & ~w13970;
assign w13972 = w13961 & ~w13971;
assign w13973 = w13961 & ~w13972;
assign w13974 = ~w13961 & ~w13971;
assign w13975 = ~w13973 & ~w13974;
assign w13976 = (~w13634 & ~w13635) | (~w13634 & w30071) | (~w13635 & w30071);
assign w13977 = w13975 & w13976;
assign w13978 = ~w13975 & ~w13976;
assign w13979 = ~w13977 & ~w13978;
assign w13980 = b_31 & w4499;
assign w13981 = w4723 & w30072;
assign w13982 = b_30 & w4494;
assign w13983 = ~w13981 & ~w13982;
assign w13984 = ~w13980 & w13983;
assign w13985 = (w13984 & ~w3345) | (w13984 & w30073) | (~w3345 & w30073);
assign w13986 = (w3345 & w40310) | (w3345 & w40311) | (w40310 & w40311);
assign w13987 = (~w3345 & w40312) | (~w3345 & w40313) | (w40312 & w40313);
assign w13988 = ~w13985 & ~w13986;
assign w13989 = ~w13987 & ~w13988;
assign w13990 = ~w13979 & w13989;
assign w13991 = w13979 & ~w13989;
assign w13992 = ~w13990 & ~w13991;
assign w13993 = ~w13827 & w13992;
assign w13994 = ~w13827 & ~w13993;
assign w13995 = w13827 & w13992;
assign w13996 = ~w13994 & ~w13995;
assign w13997 = (~w13826 & w13994) | (~w13826 & w40314) | (w13994 & w40314);
assign w13998 = ~w13994 & w40315;
assign w13999 = ~w13996 & ~w13997;
assign w14000 = ~w13998 & ~w13999;
assign w14001 = ~w13816 & w14000;
assign w14002 = w13816 & ~w14000;
assign w14003 = ~w14001 & ~w14002;
assign w14004 = (~w13684 & w13687) | (~w13684 & w30074) | (w13687 & w30074);
assign w14005 = b_40 & w2639;
assign w14006 = w2820 & w30075;
assign w14007 = b_39 & w2634;
assign w14008 = ~w14006 & ~w14007;
assign w14009 = ~w14005 & w14008;
assign w14010 = w14008 & w30076;
assign w14011 = (~w5363 & w40316) | (~w5363 & w40317) | (w40316 & w40317);
assign w14012 = (w5363 & w30078) | (w5363 & w30079) | (w30078 & w30079);
assign w14013 = ~w14011 & ~w14012;
assign w14014 = (~w13687 & w30080) | (~w13687 & w30081) | (w30080 & w30081);
assign w14015 = ~w14004 & ~w14014;
assign w14016 = ~w14013 & ~w14014;
assign w14017 = ~w14015 & ~w14016;
assign w14018 = w14003 & ~w14017;
assign w14019 = w14017 & w14003;
assign w14020 = ~w14017 & ~w14018;
assign w14021 = ~w14019 & ~w14020;
assign w14022 = w13803 & ~w14021;
assign w14023 = w13803 & ~w14022;
assign w14024 = ~w13803 & ~w14021;
assign w14025 = ~w14023 & ~w14024;
assign w14026 = b_46 & w1694;
assign w14027 = w1834 & w30082;
assign w14028 = b_45 & w1689;
assign w14029 = ~w14027 & ~w14028;
assign w14030 = ~w14026 & w14029;
assign w14031 = (w14030 & ~w6974) | (w14030 & w26328) | (~w6974 & w26328);
assign w14032 = (w6974 & w26671) | (w6974 & w26672) | (w26671 & w26672);
assign w14033 = (~w6974 & w27486) | (~w6974 & w27487) | (w27486 & w27487);
assign w14034 = ~w14031 & ~w14032;
assign w14035 = ~w14033 & ~w14034;
assign w14036 = (~w13485 & ~w13486) | (~w13485 & w27791) | (~w13486 & w27791);
assign w14037 = (~w14036 & w14034) | (~w14036 & w27488) | (w14034 & w27488);
assign w14038 = (~w27488 & w30083) | (~w27488 & w30084) | (w30083 & w30084);
assign w14039 = ~w27488 & w30085;
assign w14040 = ~w14038 & ~w14039;
assign w14041 = ~w14025 & w14040;
assign w14042 = w14025 & ~w14040;
assign w14043 = ~w14041 & ~w14042;
assign w14044 = w13789 & ~w14043;
assign w14045 = w13789 & ~w14044;
assign w14046 = ~w13789 & ~w14043;
assign w14047 = ~w14045 & ~w14046;
assign w14048 = b_52 & w986;
assign w14049 = w1069 & w30086;
assign w14050 = b_51 & w981;
assign w14051 = ~w14049 & ~w14050;
assign w14052 = ~w14048 & w14051;
assign w14053 = (w14052 & ~w8793) | (w14052 & w25652) | (~w8793 & w25652);
assign w14054 = (w8793 & w25953) | (w8793 & w25954) | (w25953 & w25954);
assign w14055 = (~w8793 & w26329) | (~w8793 & w26330) | (w26329 & w26330);
assign w14056 = ~w14053 & ~w14054;
assign w14057 = ~w14055 & ~w14056;
assign w14058 = (~w13458 & ~w13459) | (~w13458 & w30087) | (~w13459 & w30087);
assign w14059 = (w13459 & w40318) | (w13459 & w40319) | (w40318 & w40319);
assign w14060 = (w30088 & ~w13459) | (w30088 & w40320) | (~w13459 & w40320);
assign w14061 = ~w14058 & ~w14059;
assign w14062 = ~w14060 & ~w14061;
assign w14063 = ~w14061 & w30089;
assign w14064 = (w14047 & w14061) | (w14047 & w30090) | (w14061 & w30090);
assign w14065 = ~w14063 & ~w14064;
assign w14066 = w13776 & ~w14065;
assign w14067 = w13776 & ~w14066;
assign w14068 = ~w13776 & ~w14065;
assign w14069 = ~w14067 & ~w14068;
assign w14070 = (~w13719 & w13722) | (~w13719 & w27566) | (w13722 & w27566);
assign w14071 = b_58 & w418;
assign w14072 = w481 & w30091;
assign w14073 = b_57 & w413;
assign w14074 = ~w14072 & ~w14073;
assign w14075 = ~w14071 & w14074;
assign w14076 = w14074 & w30092;
assign w14077 = (~w10476 & w30093) | (~w10476 & w30094) | (w30093 & w30094);
assign w14078 = (w10476 & w30095) | (w10476 & w30096) | (w30095 & w30096);
assign w14079 = ~w14077 & ~w14078;
assign w14080 = (~w13722 & w38060) | (~w13722 & w38061) | (w38060 & w38061);
assign w14081 = ~w14070 & ~w14080;
assign w14082 = (w13722 & w38062) | (w13722 & w38063) | (w38062 & w38063);
assign w14083 = ~w14081 & ~w14082;
assign w14084 = (~w14069 & w14081) | (~w14069 & w26332) | (w14081 & w26332);
assign w14085 = ~w14069 & ~w14084;
assign w14086 = ~w14083 & ~w14084;
assign w14087 = ~w14085 & ~w14086;
assign w14088 = (~w13431 & ~w13432) | (~w13431 & w26673) | (~w13432 & w26673);
assign w14089 = b_61 & w239;
assign w14090 = w266 & w30097;
assign w14091 = b_60 & w234;
assign w14092 = ~w14090 & ~w14091;
assign w14093 = ~w14089 & w14092;
assign w14094 = w14092 & w30098;
assign w14095 = (~w11901 & w30099) | (~w11901 & w30100) | (w30099 & w30100);
assign w14096 = (w11901 & w30101) | (w11901 & w30102) | (w30101 & w30102);
assign w14097 = ~w14095 & ~w14096;
assign w14098 = ~w14088 & ~w14097;
assign w14099 = ~w14088 & ~w14098;
assign w14100 = w14088 & ~w14097;
assign w14101 = ~w14099 & ~w14100;
assign w14102 = (~w14087 & w14099) | (~w14087 & w27793) | (w14099 & w27793);
assign w14103 = ~w14087 & ~w14102;
assign w14104 = ~w14101 & ~w14102;
assign w14105 = ~w14103 & ~w14104;
assign w14106 = (~w26322 & w27794) | (~w26322 & w27795) | (w27794 & w27795);
assign w14107 = w136 & w30103;
assign w14108 = b_63 & w94;
assign w14109 = ~w14107 & ~w14108;
assign w14110 = ~w12671 & w30104;
assign w14111 = (a_5 & w14110) | (a_5 & w30105) | (w14110 & w30105);
assign w14112 = ~w14110 & w30106;
assign w14113 = ~w14111 & ~w14112;
assign w14114 = (~w27795 & w30107) | (~w27795 & w30108) | (w30107 & w30108);
assign w14115 = ~w14106 & ~w14114;
assign w14116 = (w27795 & w30109) | (w27795 & w30110) | (w30109 & w30110);
assign w14117 = (~w14105 & w14115) | (~w14105 & w26674) | (w14115 & w26674);
assign w14118 = w14105 & ~w14116;
assign w14119 = ~w14115 & w14118;
assign w14120 = ~w14117 & ~w14119;
assign w14121 = ~w13762 & w14120;
assign w14122 = ~w13762 & ~w14121;
assign w14123 = w13762 & w14120;
assign w14124 = ~w14122 & ~w14123;
assign w14125 = (~w13757 & w30111) | (~w13757 & w30112) | (w30111 & w30112);
assign w14126 = (w27786 & w38064) | (w27786 & w38065) | (w38064 & w38065);
assign w14127 = ~w14122 & w14126;
assign w14128 = ~w14125 & ~w14127;
assign w14129 = ~w14114 & ~w14117;
assign w14130 = (~w14098 & w14101) | (~w14098 & w26334) | (w14101 & w26334);
assign w14131 = w136 & w30115;
assign w14132 = (~w14131 & ~w12670) | (~w14131 & w30116) | (~w12670 & w30116);
assign w14133 = (w12670 & w40321) | (w12670 & w40322) | (w40321 & w40322);
assign w14134 = (~w12670 & w40323) | (~w12670 & w40324) | (w40323 & w40324);
assign w14135 = ~w14132 & ~w14133;
assign w14136 = ~w14134 & ~w14135;
assign w14137 = (~w14101 & w27796) | (~w14101 & w27797) | (w27796 & w27797);
assign w14138 = ~w14130 & ~w14137;
assign w14139 = (w14101 & w38066) | (w14101 & w38067) | (w38066 & w38067);
assign w14140 = ~w14138 & ~w14139;
assign w14141 = b_59 & w418;
assign w14142 = w481 & w30117;
assign w14143 = b_58 & w413;
assign w14144 = ~w14142 & ~w14143;
assign w14145 = ~w14141 & w14144;
assign w14146 = (w14145 & ~w25453) | (w14145 & w30118) | (~w25453 & w30118);
assign w14147 = a_11 & ~w14146;
assign w14148 = w14146 & a_11;
assign w14149 = ~w14146 & ~w14147;
assign w14150 = ~w14148 & ~w14149;
assign w14151 = (~w13775 & ~w13776) | (~w13775 & w30119) | (~w13776 & w30119);
assign w14152 = w14150 & w14151;
assign w14153 = ~w14150 & ~w14151;
assign w14154 = ~w14152 & ~w14153;
assign w14155 = b_56 & w657;
assign w14156 = w754 & w30120;
assign w14157 = b_55 & w652;
assign w14158 = ~w14156 & ~w14157;
assign w14159 = ~w14155 & w14158;
assign w14160 = (w14159 & ~w9798) | (w14159 & w25454) | (~w9798 & w25454);
assign w14161 = (w9798 & w25955) | (w9798 & w25956) | (w25955 & w25956);
assign w14162 = (~w9798 & w25957) | (~w9798 & w25958) | (w25957 & w25958);
assign w14163 = ~w14160 & ~w14161;
assign w14164 = ~w14162 & ~w14163;
assign w14165 = (~w14062 & w30121) | (~w14062 & w30122) | (w30121 & w30122);
assign w14166 = (w14062 & w40325) | (w14062 & w40326) | (w40325 & w40326);
assign w14167 = (~w14062 & w30123) | (~w14062 & w30124) | (w30123 & w30124);
assign w14168 = (~w13788 & ~w13789) | (~w13788 & w25959) | (~w13789 & w25959);
assign w14169 = b_53 & w986;
assign w14170 = w1069 & w30125;
assign w14171 = b_52 & w981;
assign w14172 = ~w14170 & ~w14171;
assign w14173 = ~w14169 & w14172;
assign w14174 = w14172 & w30126;
assign w14175 = (w9109 & w40327) | (w9109 & w40328) | (w40327 & w40328);
assign w14176 = (~w9109 & w40329) | (~w9109 & w40330) | (w40329 & w40330);
assign w14177 = ~w14175 & ~w14176;
assign w14178 = ~w14168 & ~w14177;
assign w14179 = w14168 & w14177;
assign w14180 = ~w14178 & ~w14179;
assign w14181 = b_50 & w1295;
assign w14182 = w1422 & w30127;
assign w14183 = b_49 & w1290;
assign w14184 = ~w14182 & ~w14183;
assign w14185 = ~w14181 & w14184;
assign w14186 = (w14185 & ~w8162) | (w14185 & w25961) | (~w8162 & w25961);
assign w14187 = (w8162 & w26339) | (w8162 & w26340) | (w26339 & w26340);
assign w14188 = (~w8162 & w27489) | (~w8162 & w27490) | (w27489 & w27490);
assign w14189 = ~w14186 & ~w14187;
assign w14190 = ~w14188 & ~w14189;
assign w14191 = (~w14037 & w14040) | (~w14037 & w25962) | (w14040 & w25962);
assign w14192 = (~w14040 & w40331) | (~w14040 & w40332) | (w40331 & w40332);
assign w14193 = (w14040 & w40333) | (w14040 & w40334) | (w40333 & w40334);
assign w14194 = (~w14040 & w40335) | (~w14040 & w40336) | (w40335 & w40336);
assign w14195 = ~w14193 & ~w14194;
assign w14196 = b_47 & w1694;
assign w14197 = w1834 & w30128;
assign w14198 = b_46 & w1689;
assign w14199 = ~w14197 & ~w14198;
assign w14200 = ~w14196 & w14199;
assign w14201 = (w14200 & ~w6998) | (w14200 & w25963) | (~w6998 & w25963);
assign w14202 = (w6998 & w26341) | (w6998 & w26342) | (w26341 & w26342);
assign w14203 = (~w6998 & w26675) | (~w6998 & w26676) | (w26675 & w26676);
assign w14204 = ~w14201 & ~w14202;
assign w14205 = (~w13802 & ~w13803) | (~w13802 & w30129) | (~w13803 & w30129);
assign w14206 = w14205 & w30130;
assign w14207 = (~w14205 & w14204) | (~w14205 & w26677) | (w14204 & w26677);
assign w14208 = ~w14206 & ~w14207;
assign w14209 = b_41 & w2639;
assign w14210 = w2820 & w30131;
assign w14211 = b_40 & w2634;
assign w14212 = ~w14210 & ~w14211;
assign w14213 = ~w14209 & w14212;
assign w14214 = (w14213 & ~w5609) | (w14213 & w27567) | (~w5609 & w27567);
assign w14215 = (w5609 & w30132) | (w5609 & w30133) | (w30132 & w30133);
assign w14216 = (~w5609 & w30134) | (~w5609 & w30135) | (w30134 & w30135);
assign w14217 = ~w14214 & ~w14215;
assign w14218 = ~w14216 & ~w14217;
assign w14219 = (w30136 & ~w13816) | (w30136 & w40337) | (~w13816 & w40337);
assign w14220 = (w13816 & w40338) | (w13816 & w40339) | (w40338 & w40339);
assign w14221 = ~w14219 & ~w14220;
assign w14222 = b_35 & w3803;
assign w14223 = w4027 & w30138;
assign w14224 = b_34 & w3798;
assign w14225 = ~w14223 & ~w14224;
assign w14226 = ~w14222 & w14225;
assign w14227 = (w14226 & ~w4181) | (w14226 & w30139) | (~w4181 & w30139);
assign w14228 = (w4181 & w40340) | (w4181 & w40341) | (w40340 & w40341);
assign w14229 = (~w4181 & w40342) | (~w4181 & w40343) | (w40342 & w40343);
assign w14230 = ~w14227 & ~w14228;
assign w14231 = ~w14229 & ~w14230;
assign w14232 = b_23 & w6761;
assign w14233 = w7075 & w30140;
assign w14234 = b_22 & w6756;
assign w14235 = ~w14233 & ~w14234;
assign w14236 = ~w14232 & w14235;
assign w14237 = (w14236 & ~w1933) | (w14236 & w30141) | (~w1933 & w30141);
assign w14238 = (w1933 & w40344) | (w1933 & w40345) | (w40344 & w40345);
assign w14239 = (~w1933 & w40346) | (~w1933 & w40347) | (w40346 & w40347);
assign w14240 = ~w14237 & ~w14238;
assign w14241 = ~w14239 & ~w14240;
assign w14242 = b_14 & w9534;
assign w14243 = w9876 & w30142;
assign w14244 = b_13 & w9529;
assign w14245 = ~w14243 & ~w14244;
assign w14246 = ~w14242 & w14245;
assign w14247 = (w14246 & ~w735) | (w14246 & w30143) | (~w735 & w30143);
assign w14248 = (w735 & w40348) | (w735 & w40349) | (w40348 & w40349);
assign w14249 = (~w735 & w40350) | (~w735 & w40351) | (w40350 & w40351);
assign w14250 = ~w14247 & ~w14248;
assign w14251 = ~w14249 & ~w14250;
assign w14252 = b_8 & w11620;
assign w14253 = w11969 & w30144;
assign w14254 = b_7 & w11615;
assign w14255 = ~w14253 & ~w14254;
assign w14256 = ~w14252 & w14255;
assign w14257 = ~w308 & w27798;
assign w14258 = (w14256 & ~w27798) | (w14256 & w40352) | (~w27798 & w40352);
assign w14259 = (w27798 & w40353) | (w27798 & w40354) | (w40353 & w40354);
assign w14260 = ~w14257 & w30146;
assign w14261 = ~w14258 & ~w14259;
assign w14262 = ~w14260 & ~w14261;
assign w14263 = w12380 & w30147;
assign w14264 = b_5 & ~w12380;
assign w14265 = ~w14263 & ~w14264;
assign w14266 = a_2 & ~w14265;
assign w14267 = w14265 & a_2;
assign w14268 = ~w14265 & ~w14266;
assign w14269 = ~w14267 & ~w14268;
assign w14270 = (~w14269 & w14261) | (~w14269 & w30148) | (w14261 & w30148);
assign w14271 = ~w14262 & ~w14270;
assign w14272 = ~w14269 & ~w14270;
assign w14273 = ~w14271 & ~w14272;
assign w14274 = ~w13851 & ~w13855;
assign w14275 = w14273 & w14274;
assign w14276 = ~w14273 & ~w14274;
assign w14277 = ~w14275 & ~w14276;
assign w14278 = b_11 & w10562;
assign w14279 = w10902 & w30149;
assign w14280 = b_10 & w10557;
assign w14281 = ~w14279 & ~w14280;
assign w14282 = ~w14278 & w14281;
assign w14283 = (w14282 & ~w530) | (w14282 & w30150) | (~w530 & w30150);
assign w14284 = (w530 & w40355) | (w530 & w40356) | (w40355 & w40356);
assign w14285 = (~w530 & w40357) | (~w530 & w40358) | (w40357 & w40358);
assign w14286 = ~w14283 & ~w14284;
assign w14287 = ~w14285 & ~w14286;
assign w14288 = ~w14277 & w14287;
assign w14289 = w14277 & ~w14287;
assign w14290 = ~w14288 & ~w14289;
assign w14291 = (~w13861 & ~w13862) | (~w13861 & w30151) | (~w13862 & w30151);
assign w14292 = w14290 & ~w14291;
assign w14293 = ~w14290 & w14291;
assign w14294 = ~w14292 & ~w14293;
assign w14295 = ~w14251 & w14294;
assign w14296 = w14294 & ~w14295;
assign w14297 = ~w14294 & ~w14251;
assign w14298 = ~w14296 & ~w14297;
assign w14299 = (~w13879 & ~w13880) | (~w13879 & w30152) | (~w13880 & w30152);
assign w14300 = ~w14298 & ~w14299;
assign w14301 = ~w14298 & ~w14300;
assign w14302 = w14298 & ~w14299;
assign w14303 = ~w14301 & ~w14302;
assign w14304 = b_17 & w8526;
assign w14305 = w8886 & w30153;
assign w14306 = b_16 & w8521;
assign w14307 = ~w14305 & ~w14306;
assign w14308 = ~w14304 & w14307;
assign w14309 = (w14308 & ~w1038) | (w14308 & w30154) | (~w1038 & w30154);
assign w14310 = (w1038 & w40359) | (w1038 & w40360) | (w40359 & w40360);
assign w14311 = (~w1038 & w40361) | (~w1038 & w40362) | (w40361 & w40362);
assign w14312 = ~w14309 & ~w14310;
assign w14313 = ~w14311 & ~w14312;
assign w14314 = (~w14313 & w14301) | (~w14313 & w30155) | (w14301 & w30155);
assign w14315 = ~w14303 & ~w14314;
assign w14316 = ~w14313 & ~w14314;
assign w14317 = ~w14315 & ~w14316;
assign w14318 = (~w13896 & ~w13898) | (~w13896 & w30156) | (~w13898 & w30156);
assign w14319 = w14317 & w14318;
assign w14320 = ~w14317 & ~w14318;
assign w14321 = ~w14319 & ~w14320;
assign w14322 = b_20 & w7613;
assign w14323 = w7941 & w30157;
assign w14324 = b_19 & w7608;
assign w14325 = ~w14323 & ~w14324;
assign w14326 = ~w14322 & w14325;
assign w14327 = (w14326 & ~w1503) | (w14326 & w30158) | (~w1503 & w30158);
assign w14328 = (w1503 & w40363) | (w1503 & w40364) | (w40363 & w40364);
assign w14329 = (~w1503 & w40365) | (~w1503 & w40366) | (w40365 & w40366);
assign w14330 = ~w14327 & ~w14328;
assign w14331 = ~w14329 & ~w14330;
assign w14332 = ~w14321 & w14331;
assign w14333 = w14321 & ~w14331;
assign w14334 = ~w14332 & ~w14333;
assign w14335 = (~w13905 & ~w13906) | (~w13905 & w30159) | (~w13906 & w30159);
assign w14336 = w14334 & ~w14335;
assign w14337 = ~w14334 & w14335;
assign w14338 = ~w14336 & ~w14337;
assign w14339 = ~w14241 & w14338;
assign w14340 = w14338 & ~w14339;
assign w14341 = ~w14338 & ~w14241;
assign w14342 = ~w14340 & ~w14341;
assign w14343 = (~w13923 & ~w13924) | (~w13923 & w30160) | (~w13924 & w30160);
assign w14344 = w14342 & w14343;
assign w14345 = ~w14342 & ~w14343;
assign w14346 = ~w14344 & ~w14345;
assign w14347 = b_26 & w5962;
assign w14348 = w6246 & w30161;
assign w14349 = b_25 & w5957;
assign w14350 = ~w14348 & ~w14349;
assign w14351 = ~w14347 & w14350;
assign w14352 = (w14351 & ~w2416) | (w14351 & w30162) | (~w2416 & w30162);
assign w14353 = (w2416 & w40367) | (w2416 & w40368) | (w40367 & w40368);
assign w14354 = (~w2416 & w40369) | (~w2416 & w40370) | (w40369 & w40370);
assign w14355 = ~w14352 & ~w14353;
assign w14356 = ~w14354 & ~w14355;
assign w14357 = w14346 & ~w14356;
assign w14358 = w14346 & ~w14357;
assign w14359 = ~w14346 & ~w14356;
assign w14360 = ~w14358 & ~w14359;
assign w14361 = (~w13940 & w13943) | (~w13940 & w30163) | (w13943 & w30163);
assign w14362 = w14360 & w14361;
assign w14363 = ~w14360 & ~w14361;
assign w14364 = ~w14362 & ~w14363;
assign w14365 = b_29 & w5196;
assign w14366 = w5459 & w30164;
assign w14367 = b_28 & w5191;
assign w14368 = ~w14366 & ~w14367;
assign w14369 = ~w14365 & w14368;
assign w14370 = (w14369 & ~w2954) | (w14369 & w30165) | (~w2954 & w30165);
assign w14371 = (w2954 & w40371) | (w2954 & w40372) | (w40371 & w40372);
assign w14372 = (~w2954 & w40373) | (~w2954 & w40374) | (w40373 & w40374);
assign w14373 = ~w14370 & ~w14371;
assign w14374 = ~w14372 & ~w14373;
assign w14375 = w14364 & ~w14374;
assign w14376 = w14364 & ~w14375;
assign w14377 = ~w14364 & ~w14374;
assign w14378 = ~w14376 & ~w14377;
assign w14379 = (~w13960 & ~w13961) | (~w13960 & w30166) | (~w13961 & w30166);
assign w14380 = w14378 & w14379;
assign w14381 = ~w14378 & ~w14379;
assign w14382 = ~w14380 & ~w14381;
assign w14383 = b_32 & w4499;
assign w14384 = w4723 & w30167;
assign w14385 = b_31 & w4494;
assign w14386 = ~w14384 & ~w14385;
assign w14387 = ~w14383 & w14386;
assign w14388 = (w14387 & ~w3545) | (w14387 & w30168) | (~w3545 & w30168);
assign w14389 = (w3545 & w40375) | (w3545 & w40376) | (w40375 & w40376);
assign w14390 = (~w3545 & w40377) | (~w3545 & w40378) | (w40377 & w40378);
assign w14391 = ~w14388 & ~w14389;
assign w14392 = ~w14390 & ~w14391;
assign w14393 = ~w14382 & w14392;
assign w14394 = w14382 & ~w14392;
assign w14395 = ~w14393 & ~w14394;
assign w14396 = (~w13978 & ~w13979) | (~w13978 & w30169) | (~w13979 & w30169);
assign w14397 = w14395 & ~w14396;
assign w14398 = ~w14395 & w14396;
assign w14399 = ~w14397 & ~w14398;
assign w14400 = ~w14231 & w14399;
assign w14401 = w14399 & ~w14400;
assign w14402 = ~w14399 & ~w14231;
assign w14403 = ~w14401 & ~w14402;
assign w14404 = b_38 & w3195;
assign w14405 = w3388 & w30170;
assign w14406 = b_37 & w3190;
assign w14407 = ~w14405 & ~w14406;
assign w14408 = ~w14404 & w14407;
assign w14409 = w14407 & w30171;
assign w14410 = (~w4658 & w40379) | (~w4658 & w40380) | (w40379 & w40380);
assign w14411 = (w4658 & w30173) | (w4658 & w30174) | (w30173 & w30174);
assign w14412 = ~w14410 & ~w14411;
assign w14413 = (~w13996 & w30175) | (~w13996 & w30176) | (w30175 & w30176);
assign w14414 = (w13996 & w30177) | (w13996 & w30178) | (w30177 & w30178);
assign w14415 = ~w14413 & ~w14414;
assign w14416 = ~w14403 & w14415;
assign w14417 = ~w14415 & ~w14403;
assign w14418 = w14415 & ~w14416;
assign w14419 = ~w14417 & ~w14418;
assign w14420 = w14221 & ~w14419;
assign w14421 = w14221 & ~w14420;
assign w14422 = ~w14221 & ~w14419;
assign w14423 = ~w14421 & ~w14422;
assign w14424 = b_44 & w2158;
assign w14425 = w2294 & w30179;
assign w14426 = b_43 & w2153;
assign w14427 = ~w14425 & ~w14426;
assign w14428 = ~w14424 & w14427;
assign w14429 = w14427 & w30180;
assign w14430 = (~w6408 & w25964) | (~w6408 & w25965) | (w25964 & w25965);
assign w14431 = (w6408 & w25966) | (w6408 & w25967) | (w25966 & w25967);
assign w14432 = ~w14430 & ~w14431;
assign w14433 = (~w14017 & w30181) | (~w14017 & w30182) | (w30181 & w30182);
assign w14434 = (~w14017 & w30183) | (~w14017 & w30184) | (w30183 & w30184);
assign w14435 = (w14017 & w40381) | (w14017 & w40382) | (w40381 & w40382);
assign w14436 = ~w14434 & ~w14435;
assign w14437 = (~w14423 & w14435) | (~w14423 & w30185) | (w14435 & w30185);
assign w14438 = ~w30185 & w40383;
assign w14439 = ~w14436 & ~w14437;
assign w14440 = ~w14438 & ~w14439;
assign w14441 = ~w14207 & w30186;
assign w14442 = w14208 & ~w14441;
assign w14443 = (~w14440 & w14207) | (~w14440 & w30187) | (w14207 & w30187);
assign w14444 = ~w14442 & ~w14443;
assign w14445 = ~w14195 & w14444;
assign w14446 = w14195 & ~w14444;
assign w14447 = ~w14445 & ~w14446;
assign w14448 = w14180 & ~w14447;
assign w14449 = w14180 & ~w14448;
assign w14450 = ~w14180 & ~w14447;
assign w14451 = ~w14449 & ~w14450;
assign w14452 = (w14451 & w14166) | (w14451 & w26343) | (w14166 & w26343);
assign w14453 = ~w14166 & w26344;
assign w14454 = ~w14452 & ~w14453;
assign w14455 = w14154 & ~w14454;
assign w14456 = w14154 & ~w14455;
assign w14457 = ~w14154 & ~w14454;
assign w14458 = ~w14456 & ~w14457;
assign w14459 = (~w14080 & w14083) | (~w14080 & w25968) | (w14083 & w25968);
assign w14460 = b_62 & w239;
assign w14461 = w266 & w30188;
assign w14462 = b_61 & w234;
assign w14463 = ~w14461 & ~w14462;
assign w14464 = ~w14460 & w14463;
assign w14465 = w14463 & w30189;
assign w14466 = (~w12273 & w40384) | (~w12273 & w40385) | (w40384 & w40385);
assign w14467 = (w12273 & w30191) | (w12273 & w30192) | (w30191 & w30192);
assign w14468 = ~w14466 & ~w14467;
assign w14469 = (~w14083 & w27799) | (~w14083 & w27800) | (w27799 & w27800);
assign w14470 = ~w14459 & ~w14469;
assign w14471 = (w14083 & w40386) | (w14083 & w40387) | (w40386 & w40387);
assign w14472 = ~w14470 & ~w14471;
assign w14473 = (~w14458 & w14470) | (~w14458 & w40388) | (w14470 & w40388);
assign w14474 = (w14458 & w14469) | (w14458 & w30193) | (w14469 & w30193);
assign w14475 = ~w14470 & w14474;
assign w14476 = ~w14473 & ~w14475;
assign w14477 = (w14476 & w14138) | (w14476 & w38068) | (w14138 & w38068);
assign w14478 = ~w14138 & w38069;
assign w14479 = ~w14477 & ~w14478;
assign w14480 = ~w14129 & w14479;
assign w14481 = ~w14129 & ~w14480;
assign w14482 = w14129 & w14479;
assign w14483 = ~w14481 & ~w14482;
assign w14484 = (~w13761 & w30194) | (~w13761 & w30195) | (w30194 & w30195);
assign w14485 = (w13757 & w37670) | (w13757 & w37671) | (w37670 & w37671);
assign w14486 = ~w14481 & w14485;
assign w14487 = ~w14484 & ~w14486;
assign w14488 = (w13757 & w37672) | (w13757 & w37673) | (w37672 & w37673);
assign w14489 = (~w14469 & w14472) | (~w14469 & w30201) | (w14472 & w30201);
assign w14490 = b_63 & w239;
assign w14491 = w266 & w30202;
assign w14492 = b_62 & w234;
assign w14493 = ~w14491 & ~w14492;
assign w14494 = ~w14490 & w14493;
assign w14495 = (w14494 & ~w12646) | (w14494 & w30203) | (~w12646 & w30203);
assign w14496 = (w12646 & w40389) | (w12646 & w40390) | (w40389 & w40390);
assign w14497 = (~w12646 & w40391) | (~w12646 & w40392) | (w40391 & w40392);
assign w14498 = ~w14495 & ~w14496;
assign w14499 = ~w14497 & ~w14498;
assign w14500 = (~w14472 & w30204) | (~w14472 & w30205) | (w30204 & w30205);
assign w14501 = ~w14489 & ~w14500;
assign w14502 = (w14472 & w40393) | (w14472 & w40394) | (w40393 & w40394);
assign w14503 = ~w14501 & ~w14502;
assign w14504 = b_60 & w418;
assign w14505 = w481 & w30206;
assign w14506 = b_59 & w413;
assign w14507 = ~w14505 & ~w14506;
assign w14508 = ~w14504 & w14507;
assign w14509 = (w14508 & ~w11196) | (w14508 & w30207) | (~w11196 & w30207);
assign w14510 = (w11196 & w40395) | (w11196 & w40396) | (w40395 & w40396);
assign w14511 = (~w11196 & w40397) | (~w11196 & w40398) | (w40397 & w40398);
assign w14512 = ~w14509 & ~w14510;
assign w14513 = ~w14511 & ~w14512;
assign w14514 = (~w14153 & ~w14154) | (~w14153 & w25969) | (~w14154 & w25969);
assign w14515 = w14513 & w14514;
assign w14516 = ~w14513 & ~w14514;
assign w14517 = ~w14515 & ~w14516;
assign w14518 = (~w14178 & ~w14180) | (~w14178 & w30208) | (~w14180 & w30208);
assign w14519 = b_54 & w986;
assign w14520 = w1069 & w30209;
assign w14521 = b_53 & w981;
assign w14522 = ~w14520 & ~w14521;
assign w14523 = ~w14519 & w14522;
assign w14524 = (w14523 & ~w9134) | (w14523 & w26345) | (~w9134 & w26345);
assign w14525 = (w9134 & w30210) | (w9134 & w30211) | (w30210 & w30211);
assign w14526 = (~w9134 & w30212) | (~w9134 & w30213) | (w30212 & w30213);
assign w14527 = ~w14524 & ~w14525;
assign w14528 = ~w14526 & ~w14527;
assign w14529 = ~w14518 & ~w14528;
assign w14530 = ~w14518 & ~w14529;
assign w14531 = w14518 & ~w14528;
assign w14532 = ~w14530 & ~w14531;
assign w14533 = b_48 & w1694;
assign w14534 = w1834 & w30214;
assign w14535 = b_47 & w1689;
assign w14536 = ~w14534 & ~w14535;
assign w14537 = ~w14533 & w14536;
assign w14538 = (w14537 & ~w7284) | (w14537 & w27568) | (~w7284 & w27568);
assign w14539 = (w7284 & w27801) | (w7284 & w27802) | (w27801 & w27802);
assign w14540 = (~w7284 & w30215) | (~w7284 & w30216) | (w30215 & w30216);
assign w14541 = ~w14538 & ~w14539;
assign w14542 = ~w14540 & ~w14541;
assign w14543 = (~w14207 & ~w14208) | (~w14207 & w27569) | (~w14208 & w27569);
assign w14544 = (~w14208 & w40399) | (~w14208 & w40400) | (w40399 & w40400);
assign w14545 = (w14208 & w40401) | (w14208 & w40402) | (w40401 & w40402);
assign w14546 = ~w14544 & ~w14545;
assign w14547 = (~w14433 & w14436) | (~w14433 & w26346) | (w14436 & w26346);
assign w14548 = b_45 & w2158;
assign w14549 = w2294 & w30217;
assign w14550 = b_44 & w2153;
assign w14551 = ~w14549 & ~w14550;
assign w14552 = ~w14548 & w14551;
assign w14553 = (w14552 & ~w6682) | (w14552 & w26347) | (~w6682 & w26347);
assign w14554 = (w6682 & w27570) | (w6682 & w27571) | (w27570 & w27571);
assign w14555 = (~w6682 & w30218) | (~w6682 & w30219) | (w30218 & w30219);
assign w14556 = ~w14553 & ~w14554;
assign w14557 = ~w14555 & ~w14556;
assign w14558 = (~w14436 & w30220) | (~w14436 & w30221) | (w30220 & w30221);
assign w14559 = ~w14547 & ~w14558;
assign w14560 = (w14436 & w30222) | (w14436 & w30223) | (w30222 & w30223);
assign w14561 = b_42 & w2639;
assign w14562 = w2820 & w30224;
assign w14563 = b_41 & w2634;
assign w14564 = ~w14562 & ~w14563;
assign w14565 = ~w14561 & w14564;
assign w14566 = (w14565 & ~w5864) | (w14565 & w30225) | (~w5864 & w30225);
assign w14567 = (w5864 & w40403) | (w5864 & w40404) | (w40403 & w40404);
assign w14568 = (~w5864 & w40405) | (~w5864 & w40406) | (w40405 & w40406);
assign w14569 = ~w14566 & ~w14567;
assign w14570 = ~w14568 & ~w14569;
assign w14571 = (w30226 & w40407) | (w30226 & w40408) | (w40407 & w40408);
assign w14572 = (~w30226 & w40409) | (~w30226 & w40410) | (w40409 & w40410);
assign w14573 = ~w14571 & ~w14572;
assign w14574 = (~w14397 & ~w14399) | (~w14397 & w30227) | (~w14399 & w30227);
assign w14575 = (~w14381 & ~w14382) | (~w14381 & w30228) | (~w14382 & w30228);
assign w14576 = (~w14363 & ~w14364) | (~w14363 & w30229) | (~w14364 & w30229);
assign w14577 = (~w14336 & ~w14338) | (~w14336 & w30230) | (~w14338 & w30230);
assign w14578 = (~w14320 & ~w14321) | (~w14320 & w30231) | (~w14321 & w30231);
assign w14579 = (~w14276 & ~w14277) | (~w14276 & w30232) | (~w14277 & w30232);
assign w14580 = b_12 & w10562;
assign w14581 = w10902 & w30233;
assign w14582 = b_11 & w10557;
assign w14583 = ~w14581 & ~w14582;
assign w14584 = ~w14580 & w14583;
assign w14585 = (w14584 & ~w552) | (w14584 & w30234) | (~w552 & w30234);
assign w14586 = (w552 & w40411) | (w552 & w40412) | (w40411 & w40412);
assign w14587 = (~w552 & w40413) | (~w552 & w40414) | (w40413 & w40414);
assign w14588 = ~w14585 & ~w14586;
assign w14589 = ~w14587 & ~w14588;
assign w14590 = w12380 & w30235;
assign w14591 = b_6 & ~w12380;
assign w14592 = ~w14590 & ~w14591;
assign w14593 = a_2 & ~a_5;
assign w14594 = ~a_2 & a_5;
assign w14595 = ~w14593 & ~w14594;
assign w14596 = ~w14592 & ~w14595;
assign w14597 = w14592 & w14595;
assign w14598 = ~w14596 & ~w14597;
assign w14599 = ~w14270 & w30236;
assign w14600 = (w14598 & w14270) | (w14598 & w30237) | (w14270 & w30237);
assign w14601 = ~w14599 & ~w14600;
assign w14602 = b_9 & w11620;
assign w14603 = w11969 & w30238;
assign w14604 = b_8 & w11615;
assign w14605 = ~w14603 & ~w14604;
assign w14606 = ~w14602 & w14605;
assign w14607 = (w14606 & ~w371) | (w14606 & w30239) | (~w371 & w30239);
assign w14608 = (w371 & w40415) | (w371 & w40416) | (w40415 & w40416);
assign w14609 = (~w371 & w40417) | (~w371 & w40418) | (w40417 & w40418);
assign w14610 = ~w14607 & ~w14608;
assign w14611 = ~w14609 & ~w14610;
assign w14612 = ~w14601 & w14611;
assign w14613 = w14601 & ~w14611;
assign w14614 = ~w14612 & ~w14613;
assign w14615 = ~w14589 & w14614;
assign w14616 = ~w14614 & ~w14589;
assign w14617 = w14614 & ~w14615;
assign w14618 = ~w14616 & ~w14617;
assign w14619 = (~w14579 & w14617) | (~w14579 & w30240) | (w14617 & w30240);
assign w14620 = ~w14579 & ~w14619;
assign w14621 = ~w14618 & ~w14619;
assign w14622 = ~w14620 & ~w14621;
assign w14623 = b_15 & w9534;
assign w14624 = w9876 & w30241;
assign w14625 = b_14 & w9529;
assign w14626 = ~w14624 & ~w14625;
assign w14627 = ~w14623 & w14626;
assign w14628 = (w14627 & ~w827) | (w14627 & w30242) | (~w827 & w30242);
assign w14629 = (w827 & w40419) | (w827 & w40420) | (w40419 & w40420);
assign w14630 = (~w827 & w40421) | (~w827 & w40422) | (w40421 & w40422);
assign w14631 = ~w14628 & ~w14629;
assign w14632 = ~w14630 & ~w14631;
assign w14633 = ~w14622 & ~w14632;
assign w14634 = ~w14622 & ~w14633;
assign w14635 = w14622 & ~w14632;
assign w14636 = (~w14292 & ~w14294) | (~w14292 & w30243) | (~w14294 & w30243);
assign w14637 = ~w14634 & w30244;
assign w14638 = (~w14636 & w14634) | (~w14636 & w30245) | (w14634 & w30245);
assign w14639 = ~w14637 & ~w14638;
assign w14640 = b_18 & w8526;
assign w14641 = w8886 & w30246;
assign w14642 = b_17 & w8521;
assign w14643 = ~w14641 & ~w14642;
assign w14644 = ~w14640 & w14643;
assign w14645 = (w14644 & ~w1238) | (w14644 & w30247) | (~w1238 & w30247);
assign w14646 = (w1238 & w40423) | (w1238 & w40424) | (w40423 & w40424);
assign w14647 = (~w1238 & w40425) | (~w1238 & w40426) | (w40425 & w40426);
assign w14648 = ~w14645 & ~w14646;
assign w14649 = ~w14647 & ~w14648;
assign w14650 = w14639 & ~w14649;
assign w14651 = w14639 & ~w14650;
assign w14652 = ~w14639 & ~w14649;
assign w14653 = ~w14651 & ~w14652;
assign w14654 = ~w14300 & ~w14314;
assign w14655 = w14653 & w14654;
assign w14656 = ~w14653 & ~w14654;
assign w14657 = ~w14655 & ~w14656;
assign w14658 = b_21 & w7613;
assign w14659 = w7941 & w30248;
assign w14660 = b_20 & w7608;
assign w14661 = ~w14659 & ~w14660;
assign w14662 = ~w14658 & w14661;
assign w14663 = (w14662 & ~w1634) | (w14662 & w30249) | (~w1634 & w30249);
assign w14664 = (w1634 & w40427) | (w1634 & w40428) | (w40427 & w40428);
assign w14665 = (~w1634 & w40429) | (~w1634 & w40430) | (w40429 & w40430);
assign w14666 = ~w14663 & ~w14664;
assign w14667 = ~w14665 & ~w14666;
assign w14668 = w14657 & ~w14667;
assign w14669 = w14657 & ~w14668;
assign w14670 = ~w14657 & ~w14667;
assign w14671 = ~w14669 & w30250;
assign w14672 = (w14578 & w14669) | (w14578 & w30251) | (w14669 & w30251);
assign w14673 = ~w14671 & ~w14672;
assign w14674 = b_24 & w6761;
assign w14675 = w7075 & w30252;
assign w14676 = b_23 & w6756;
assign w14677 = ~w14675 & ~w14676;
assign w14678 = ~w14674 & w14677;
assign w14679 = (w14678 & ~w2083) | (w14678 & w30253) | (~w2083 & w30253);
assign w14680 = (w2083 & w40431) | (w2083 & w40432) | (w40431 & w40432);
assign w14681 = (~w2083 & w40433) | (~w2083 & w40434) | (w40433 & w40434);
assign w14682 = ~w14679 & ~w14680;
assign w14683 = ~w14681 & ~w14682;
assign w14684 = ~w14673 & ~w14683;
assign w14685 = w14673 & w14683;
assign w14686 = ~w14684 & ~w14685;
assign w14687 = w14577 & ~w14686;
assign w14688 = ~w14577 & w14686;
assign w14689 = ~w14687 & ~w14688;
assign w14690 = b_27 & w5962;
assign w14691 = w6246 & w30254;
assign w14692 = b_26 & w5957;
assign w14693 = ~w14691 & ~w14692;
assign w14694 = ~w14690 & w14693;
assign w14695 = (w14694 & ~w2582) | (w14694 & w30255) | (~w2582 & w30255);
assign w14696 = (w2582 & w40435) | (w2582 & w40436) | (w40435 & w40436);
assign w14697 = (~w2582 & w40437) | (~w2582 & w40438) | (w40437 & w40438);
assign w14698 = ~w14695 & ~w14696;
assign w14699 = ~w14697 & ~w14698;
assign w14700 = w14689 & ~w14699;
assign w14701 = w14689 & ~w14700;
assign w14702 = ~w14689 & ~w14699;
assign w14703 = ~w14701 & ~w14702;
assign w14704 = (~w14345 & ~w14346) | (~w14345 & w30256) | (~w14346 & w30256);
assign w14705 = w14703 & w14704;
assign w14706 = ~w14703 & ~w14704;
assign w14707 = ~w14705 & ~w14706;
assign w14708 = b_30 & w5196;
assign w14709 = w5459 & w30257;
assign w14710 = b_29 & w5191;
assign w14711 = ~w14709 & ~w14710;
assign w14712 = ~w14708 & w14711;
assign w14713 = (w14712 & ~w3138) | (w14712 & w30258) | (~w3138 & w30258);
assign w14714 = (w3138 & w40439) | (w3138 & w40440) | (w40439 & w40440);
assign w14715 = (~w3138 & w40441) | (~w3138 & w40442) | (w40441 & w40442);
assign w14716 = ~w14713 & ~w14714;
assign w14717 = ~w14715 & ~w14716;
assign w14718 = w14707 & ~w14717;
assign w14719 = ~w14707 & w14717;
assign w14720 = (w14364 & w40443) | (w14364 & w40444) | (w40443 & w40444);
assign w14721 = ~w14576 & ~w14720;
assign w14722 = (~w14718 & w14576) | (~w14718 & w30260) | (w14576 & w30260);
assign w14723 = (w14576 & w30259) | (w14576 & w40445) | (w30259 & w40445);
assign w14724 = ~w14721 & ~w14723;
assign w14725 = b_33 & w4499;
assign w14726 = w4723 & w30261;
assign w14727 = b_32 & w4494;
assign w14728 = ~w14726 & ~w14727;
assign w14729 = ~w14725 & w14728;
assign w14730 = (w14729 & ~w3744) | (w14729 & w30262) | (~w3744 & w30262);
assign w14731 = (w3744 & w40446) | (w3744 & w40447) | (w40446 & w40447);
assign w14732 = (~w3744 & w40448) | (~w3744 & w40449) | (w40448 & w40449);
assign w14733 = ~w14730 & ~w14731;
assign w14734 = ~w14732 & ~w14733;
assign w14735 = ~w14724 & ~w14734;
assign w14736 = ~w14724 & ~w14735;
assign w14737 = w14724 & ~w14734;
assign w14738 = ~w14736 & ~w14737;
assign w14739 = ~w14575 & w14738;
assign w14740 = w14575 & ~w14738;
assign w14741 = ~w14739 & ~w14740;
assign w14742 = b_36 & w3803;
assign w14743 = w4027 & w30263;
assign w14744 = b_35 & w3798;
assign w14745 = ~w14743 & ~w14744;
assign w14746 = ~w14742 & w14745;
assign w14747 = (w14746 & ~w4395) | (w14746 & w30264) | (~w4395 & w30264);
assign w14748 = (w4395 & w40450) | (w4395 & w40451) | (w40450 & w40451);
assign w14749 = (~w4395 & w40452) | (~w4395 & w40453) | (w40452 & w40453);
assign w14750 = ~w14747 & ~w14748;
assign w14751 = ~w14749 & ~w14750;
assign w14752 = ~w14741 & ~w14751;
assign w14753 = w14741 & w14751;
assign w14754 = ~w14752 & ~w14753;
assign w14755 = w14574 & ~w14754;
assign w14756 = ~w14574 & w14754;
assign w14757 = ~w14755 & ~w14756;
assign w14758 = b_39 & w3195;
assign w14759 = w3388 & w30265;
assign w14760 = b_38 & w3190;
assign w14761 = ~w14759 & ~w14760;
assign w14762 = ~w14758 & w14761;
assign w14763 = (w14762 & ~w4888) | (w14762 & w30266) | (~w4888 & w30266);
assign w14764 = (w4888 & w40454) | (w4888 & w40455) | (w40454 & w40455);
assign w14765 = (~w4888 & w40456) | (~w4888 & w40457) | (w40456 & w40457);
assign w14766 = ~w14763 & ~w14764;
assign w14767 = ~w14765 & ~w14766;
assign w14768 = (~w14413 & ~w14415) | (~w14413 & w30267) | (~w14415 & w30267);
assign w14769 = w14767 & w14768;
assign w14770 = ~w14767 & ~w14768;
assign w14771 = ~w14769 & ~w14770;
assign w14772 = w14757 & w14771;
assign w14773 = ~w14757 & ~w14771;
assign w14774 = ~w14772 & ~w14773;
assign w14775 = w14573 & w14774;
assign w14776 = ~w14573 & ~w14774;
assign w14777 = ~w14775 & ~w14776;
assign w14778 = (~w14777 & w14559) | (~w14777 & w30268) | (w14559 & w30268);
assign w14779 = ~w14559 & w30269;
assign w14780 = ~w14778 & ~w14779;
assign w14781 = w14546 & ~w14780;
assign w14782 = w14546 & ~w14781;
assign w14783 = ~w14546 & ~w14780;
assign w14784 = ~w14782 & ~w14783;
assign w14785 = b_51 & w1295;
assign w14786 = w1422 & w30270;
assign w14787 = b_50 & w1290;
assign w14788 = ~w14786 & ~w14787;
assign w14789 = ~w14785 & w14788;
assign w14790 = (w14789 & ~w8186) | (w14789 & w27572) | (~w8186 & w27572);
assign w14791 = (w8186 & w30271) | (w8186 & w30272) | (w30271 & w30272);
assign w14792 = (~w8186 & w30273) | (~w8186 & w30274) | (w30273 & w30274);
assign w14793 = ~w14790 & ~w14791;
assign w14794 = ~w14792 & ~w14793;
assign w14795 = (~w14192 & w14195) | (~w14192 & w27491) | (w14195 & w27491);
assign w14796 = ~w14794 & ~w14795;
assign w14797 = w14794 & w14795;
assign w14798 = ~w14796 & ~w14797;
assign w14799 = ~w14784 & w14798;
assign w14800 = ~w14798 & ~w14784;
assign w14801 = w14798 & ~w14799;
assign w14802 = ~w14800 & ~w14801;
assign w14803 = (~w14802 & w14530) | (~w14802 & w40458) | (w14530 & w40458);
assign w14804 = ~w14532 & ~w14803;
assign w14805 = ~w14530 & w40459;
assign w14806 = ~w14804 & ~w14805;
assign w14807 = b_57 & w657;
assign w14808 = w754 & w30275;
assign w14809 = b_56 & w652;
assign w14810 = ~w14808 & ~w14809;
assign w14811 = ~w14807 & w14810;
assign w14812 = (w14811 & ~w10452) | (w14811 & w30276) | (~w10452 & w30276);
assign w14813 = (w10452 & w40460) | (w10452 & w40461) | (w40460 & w40461);
assign w14814 = (~w10452 & w40462) | (~w10452 & w40463) | (w40462 & w40463);
assign w14815 = ~w14812 & ~w14813;
assign w14816 = ~w14814 & ~w14815;
assign w14817 = (~w14451 & w14166) | (~w14451 & w25970) | (w14166 & w25970);
assign w14818 = (~w14816 & w14817) | (~w14816 & w26348) | (w14817 & w26348);
assign w14819 = ~w14817 & w26349;
assign w14820 = ~w14818 & ~w14819;
assign w14821 = ~w14806 & w14820;
assign w14822 = ~w14820 & ~w14806;
assign w14823 = w14820 & ~w14821;
assign w14824 = ~w14822 & ~w14823;
assign w14825 = w14517 & ~w14824;
assign w14826 = w14517 & ~w14825;
assign w14827 = ~w14517 & ~w14824;
assign w14828 = ~w14826 & ~w14827;
assign w14829 = (w14828 & w14501) | (w14828 & w40464) | (w14501 & w40464);
assign w14830 = ~w14501 & w40465;
assign w14831 = ~w14829 & ~w14830;
assign w14832 = (~w14140 & w40466) | (~w14140 & w40467) | (w40466 & w40467);
assign w14833 = (w14140 & w40468) | (w14140 & w40469) | (w40468 & w40469);
assign w14834 = ~w14832 & ~w14833;
assign w14835 = (~w13757 & w37674) | (~w13757 & w37675) | (w37674 & w37675);
assign w14836 = w14488 & ~w14834;
assign w14837 = ~w14835 & ~w14836;
assign w14838 = (~w14516 & ~w14517) | (~w14516 & w30279) | (~w14517 & w30279);
assign w14839 = w266 & w30280;
assign w14840 = b_63 & w234;
assign w14841 = ~w14839 & ~w14840;
assign w14842 = ~w12671 & w30281;
assign w14843 = (a_8 & w14842) | (a_8 & w30282) | (w14842 & w30282);
assign w14844 = ~w14842 & w30283;
assign w14845 = ~w14843 & ~w14844;
assign w14846 = ~w14838 & ~w14845;
assign w14847 = w14838 & w14845;
assign w14848 = ~w14846 & ~w14847;
assign w14849 = b_61 & w418;
assign w14850 = w481 & w30284;
assign w14851 = b_60 & w413;
assign w14852 = ~w14850 & ~w14851;
assign w14853 = ~w14849 & w14852;
assign w14854 = (w14853 & ~w11901) | (w14853 & w30285) | (~w11901 & w30285);
assign w14855 = (w11901 & w40470) | (w11901 & w40471) | (w40470 & w40471);
assign w14856 = (~w11901 & w40472) | (~w11901 & w40473) | (w40472 & w40473);
assign w14857 = ~w14854 & ~w14855;
assign w14858 = ~w14856 & ~w14857;
assign w14859 = (~w14818 & ~w14820) | (~w14818 & w30286) | (~w14820 & w30286);
assign w14860 = w14858 & w14859;
assign w14861 = ~w14858 & ~w14859;
assign w14862 = ~w14860 & ~w14861;
assign w14863 = b_58 & w657;
assign w14864 = w754 & w30287;
assign w14865 = b_57 & w652;
assign w14866 = ~w14864 & ~w14865;
assign w14867 = ~w14863 & w14866;
assign w14868 = w14866 & w30288;
assign w14869 = (~w10476 & w30289) | (~w10476 & w30290) | (w30289 & w30290);
assign w14870 = (w10476 & w30291) | (w10476 & w30292) | (w30291 & w30292);
assign w14871 = ~w14869 & ~w14870;
assign w14872 = (~w14532 & w40474) | (~w14532 & w40475) | (w40474 & w40475);
assign w14873 = (w14532 & w40476) | (w14532 & w40477) | (w40476 & w40477);
assign w14874 = ~w14872 & ~w14873;
assign w14875 = b_55 & w986;
assign w14876 = w1069 & w30293;
assign w14877 = b_54 & w981;
assign w14878 = ~w14876 & ~w14877;
assign w14879 = ~w14875 & w14878;
assign w14880 = (w14879 & ~w9776) | (w14879 & w27574) | (~w9776 & w27574);
assign w14881 = (w9776 & w30294) | (w9776 & w30295) | (w30294 & w30295);
assign w14882 = (~w9776 & w30296) | (~w9776 & w30297) | (w30296 & w30297);
assign w14883 = ~w14880 & ~w14881;
assign w14884 = ~w14882 & ~w14883;
assign w14885 = (~w14796 & ~w14798) | (~w14796 & w27575) | (~w14798 & w27575);
assign w14886 = w14884 & w14885;
assign w14887 = ~w14884 & ~w14885;
assign w14888 = ~w14886 & ~w14887;
assign w14889 = b_52 & w1295;
assign w14890 = w1422 & w30298;
assign w14891 = b_51 & w1290;
assign w14892 = ~w14890 & ~w14891;
assign w14893 = ~w14889 & w14892;
assign w14894 = (w14893 & ~w8793) | (w14893 & w26350) | (~w8793 & w26350);
assign w14895 = (w8793 & w27803) | (w8793 & w27804) | (w27803 & w27804);
assign w14896 = (~w8793 & w30299) | (~w8793 & w30300) | (w30299 & w30300);
assign w14897 = ~w14894 & ~w14895;
assign w14898 = ~w14896 & ~w14897;
assign w14899 = (~w14545 & ~w14546) | (~w14545 & w27805) | (~w14546 & w27805);
assign w14900 = w14898 & w14899;
assign w14901 = ~w14898 & ~w14899;
assign w14902 = ~w14900 & ~w14901;
assign w14903 = b_49 & w1694;
assign w14904 = w1834 & w30301;
assign w14905 = b_48 & w1689;
assign w14906 = ~w14904 & ~w14905;
assign w14907 = ~w14903 & w14906;
assign w14908 = (w14907 & ~w7859) | (w14907 & w25456) | (~w7859 & w25456);
assign w14909 = (w7859 & w25971) | (w7859 & w25972) | (w25971 & w25972);
assign w14910 = (~w7859 & w26351) | (~w7859 & w26352) | (w26351 & w26352);
assign w14911 = ~w14908 & ~w14909;
assign w14912 = ~w14910 & ~w14911;
assign w14913 = (w14777 & w14559) | (w14777 & w27576) | (w14559 & w27576);
assign w14914 = (~w14912 & w14913) | (~w14912 & w30302) | (w14913 & w30302);
assign w14915 = ~w14913 & w30303;
assign w14916 = (w14912 & w14913) | (w14912 & w30304) | (w14913 & w30304);
assign w14917 = ~w14915 & ~w14916;
assign w14918 = (~w14572 & ~w14573) | (~w14572 & w30305) | (~w14573 & w30305);
assign w14919 = b_46 & w2158;
assign w14920 = w2294 & w30306;
assign w14921 = b_45 & w2153;
assign w14922 = ~w14920 & ~w14921;
assign w14923 = ~w14919 & w14922;
assign w14924 = w14922 & w30307;
assign w14925 = (~w6974 & w27577) | (~w6974 & w27578) | (w27577 & w27578);
assign w14926 = (w6974 & w27579) | (w6974 & w27580) | (w27579 & w27580);
assign w14927 = ~w14925 & ~w14926;
assign w14928 = ~w14918 & ~w14927;
assign w14929 = w14918 & w14927;
assign w14930 = ~w14928 & ~w14929;
assign w14931 = b_43 & w2639;
assign w14932 = w2820 & w30308;
assign w14933 = b_42 & w2634;
assign w14934 = ~w14932 & ~w14933;
assign w14935 = ~w14931 & w14934;
assign w14936 = (w14935 & ~w5888) | (w14935 & w30309) | (~w5888 & w30309);
assign w14937 = (w5888 & w40478) | (w5888 & w40479) | (w40478 & w40479);
assign w14938 = (~w5888 & w40480) | (~w5888 & w40481) | (w40480 & w40481);
assign w14939 = ~w14936 & ~w14937;
assign w14940 = ~w14938 & ~w14939;
assign w14941 = (~w14770 & ~w14771) | (~w14770 & w30310) | (~w14771 & w30310);
assign w14942 = (w14771 & w40482) | (w14771 & w40483) | (w40482 & w40483);
assign w14943 = ~w14941 & ~w14942;
assign w14944 = b_40 & w3195;
assign w14945 = w3388 & w30311;
assign w14946 = b_39 & w3190;
assign w14947 = ~w14945 & ~w14946;
assign w14948 = ~w14944 & w14947;
assign w14949 = (w14948 & ~w5363) | (w14948 & w30312) | (~w5363 & w30312);
assign w14950 = (w5363 & w40484) | (w5363 & w40485) | (w40484 & w40485);
assign w14951 = (~w5363 & w40486) | (~w5363 & w40487) | (w40486 & w40487);
assign w14952 = ~w14949 & ~w14950;
assign w14953 = ~w14951 & ~w14952;
assign w14954 = ~w14756 & w30313;
assign w14955 = (~w14953 & w14756) | (~w14953 & w30314) | (w14756 & w30314);
assign w14956 = ~w14954 & ~w14955;
assign w14957 = b_37 & w3803;
assign w14958 = w4027 & w30315;
assign w14959 = b_36 & w3798;
assign w14960 = ~w14958 & ~w14959;
assign w14961 = ~w14957 & w14960;
assign w14962 = (w14961 & ~w4636) | (w14961 & w30316) | (~w4636 & w30316);
assign w14963 = (w4636 & w40488) | (w4636 & w40489) | (w40488 & w40489);
assign w14964 = (~w4636 & w40490) | (~w4636 & w40491) | (w40490 & w40491);
assign w14965 = ~w14962 & ~w14963;
assign w14966 = ~w14964 & ~w14965;
assign w14967 = (~w14735 & w14738) | (~w14735 & w30317) | (w14738 & w30317);
assign w14968 = b_34 & w4499;
assign w14969 = w4723 & w30318;
assign w14970 = b_33 & w4494;
assign w14971 = ~w14969 & ~w14970;
assign w14972 = ~w14968 & w14971;
assign w14973 = (w14972 & ~w3967) | (w14972 & w30319) | (~w3967 & w30319);
assign w14974 = (w3967 & w40492) | (w3967 & w40493) | (w40492 & w40493);
assign w14975 = (~w3967 & w40494) | (~w3967 & w40495) | (w40494 & w40495);
assign w14976 = ~w14973 & ~w14974;
assign w14977 = ~w14975 & ~w14976;
assign w14978 = (~w14600 & ~w14601) | (~w14600 & w30320) | (~w14601 & w30320);
assign w14979 = ~a_2 & ~a_5;
assign w14980 = (~w14979 & w14592) | (~w14979 & w30321) | (w14592 & w30321);
assign w14981 = w12380 & w30322;
assign w14982 = b_7 & ~w12380;
assign w14983 = ~w14981 & ~w14982;
assign w14984 = ~w14980 & w14983;
assign w14985 = w14980 & ~w14983;
assign w14986 = ~w14984 & ~w14985;
assign w14987 = b_10 & w11620;
assign w14988 = w11969 & w30323;
assign w14989 = b_9 & w11615;
assign w14990 = ~w14988 & ~w14989;
assign w14991 = ~w14987 & w14990;
assign w14992 = w14990 & w30324;
assign w14993 = (~w454 & w40496) | (~w454 & w40497) | (w40496 & w40497);
assign w14994 = (w454 & w30326) | (w454 & w30327) | (w30326 & w30327);
assign w14995 = (w14986 & w14993) | (w14986 & w30328) | (w14993 & w30328);
assign w14996 = ~w14993 & w30329;
assign w14997 = ~w14995 & ~w14996;
assign w14998 = ~w14978 & w14997;
assign w14999 = w14978 & ~w14997;
assign w15000 = ~w14998 & ~w14999;
assign w15001 = b_13 & w10562;
assign w15002 = w10902 & w30330;
assign w15003 = b_12 & w10557;
assign w15004 = ~w15002 & ~w15003;
assign w15005 = ~w15001 & w15004;
assign w15006 = (w15005 & ~w711) | (w15005 & w30331) | (~w711 & w30331);
assign w15007 = (w711 & w40498) | (w711 & w40499) | (w40498 & w40499);
assign w15008 = (~w711 & w40500) | (~w711 & w40501) | (w40500 & w40501);
assign w15009 = ~w15006 & ~w15007;
assign w15010 = ~w15008 & ~w15009;
assign w15011 = w15000 & ~w15010;
assign w15012 = w15000 & ~w15011;
assign w15013 = ~w15000 & ~w15010;
assign w15014 = ~w15012 & ~w15013;
assign w15015 = ~w14615 & ~w14619;
assign w15016 = w15014 & w15015;
assign w15017 = ~w15014 & ~w15015;
assign w15018 = ~w15016 & ~w15017;
assign w15019 = b_16 & w9534;
assign w15020 = w9876 & w30332;
assign w15021 = b_15 & w9529;
assign w15022 = ~w15020 & ~w15021;
assign w15023 = ~w15019 & w15022;
assign w15024 = (w15023 & ~w926) | (w15023 & w30333) | (~w926 & w30333);
assign w15025 = (w926 & w40502) | (w926 & w40503) | (w40502 & w40503);
assign w15026 = (~w926 & w40504) | (~w926 & w40505) | (w40504 & w40505);
assign w15027 = ~w15024 & ~w15025;
assign w15028 = ~w15026 & ~w15027;
assign w15029 = w15018 & ~w15028;
assign w15030 = w15018 & ~w15029;
assign w15031 = ~w15018 & ~w15028;
assign w15032 = ~w15030 & ~w15031;
assign w15033 = ~w14633 & ~w14638;
assign w15034 = w15032 & w15033;
assign w15035 = ~w15032 & ~w15033;
assign w15036 = ~w15034 & ~w15035;
assign w15037 = b_19 & w8526;
assign w15038 = w8886 & w30334;
assign w15039 = b_18 & w8521;
assign w15040 = ~w15038 & ~w15039;
assign w15041 = ~w15037 & w15040;
assign w15042 = (w15041 & ~w1372) | (w15041 & w30335) | (~w1372 & w30335);
assign w15043 = (w1372 & w40506) | (w1372 & w40507) | (w40506 & w40507);
assign w15044 = (~w1372 & w40508) | (~w1372 & w40509) | (w40508 & w40509);
assign w15045 = ~w15042 & ~w15043;
assign w15046 = ~w15044 & ~w15045;
assign w15047 = w15036 & ~w15046;
assign w15048 = w15036 & ~w15047;
assign w15049 = ~w15036 & ~w15046;
assign w15050 = ~w15048 & ~w15049;
assign w15051 = (~w14650 & w14653) | (~w14650 & w30336) | (w14653 & w30336);
assign w15052 = w15050 & w15051;
assign w15053 = ~w15050 & ~w15051;
assign w15054 = ~w15052 & ~w15053;
assign w15055 = b_22 & w7613;
assign w15056 = w7941 & w30337;
assign w15057 = b_21 & w7608;
assign w15058 = ~w15056 & ~w15057;
assign w15059 = ~w15055 & w15058;
assign w15060 = (w15059 & ~w1786) | (w15059 & w30338) | (~w1786 & w30338);
assign w15061 = (w1786 & w40510) | (w1786 & w40511) | (w40510 & w40511);
assign w15062 = (~w1786 & w40512) | (~w1786 & w40513) | (w40512 & w40513);
assign w15063 = ~w15060 & ~w15061;
assign w15064 = ~w15062 & ~w15063;
assign w15065 = w15054 & ~w15064;
assign w15066 = w15054 & ~w15065;
assign w15067 = ~w15054 & ~w15064;
assign w15068 = ~w15066 & ~w15067;
assign w15069 = (~w14578 & w14669) | (~w14578 & w30339) | (w14669 & w30339);
assign w15070 = ~w14668 & ~w15069;
assign w15071 = w15068 & w15070;
assign w15072 = ~w15068 & ~w15070;
assign w15073 = ~w15071 & ~w15072;
assign w15074 = b_25 & w6761;
assign w15075 = w7075 & w30340;
assign w15076 = b_24 & w6756;
assign w15077 = ~w15075 & ~w15076;
assign w15078 = ~w15074 & w15077;
assign w15079 = (w15078 & ~w2108) | (w15078 & w30341) | (~w2108 & w30341);
assign w15080 = (w2108 & w40514) | (w2108 & w40515) | (w40514 & w40515);
assign w15081 = (~w2108 & w40516) | (~w2108 & w40517) | (w40516 & w40517);
assign w15082 = ~w15079 & ~w15080;
assign w15083 = ~w15081 & ~w15082;
assign w15084 = w15073 & ~w15083;
assign w15085 = w15073 & ~w15084;
assign w15086 = ~w15073 & ~w15083;
assign w15087 = (~w14684 & ~w14686) | (~w14684 & w30342) | (~w14686 & w30342);
assign w15088 = ~w15085 & w30343;
assign w15089 = (~w15087 & w15085) | (~w15087 & w30344) | (w15085 & w30344);
assign w15090 = ~w15088 & ~w15089;
assign w15091 = b_28 & w5962;
assign w15092 = w6246 & w30345;
assign w15093 = b_27 & w5957;
assign w15094 = ~w15092 & ~w15093;
assign w15095 = ~w15091 & w15094;
assign w15096 = (w15095 & ~w2771) | (w15095 & w30346) | (~w2771 & w30346);
assign w15097 = (w2771 & w40518) | (w2771 & w40519) | (w40518 & w40519);
assign w15098 = (~w2771 & w40520) | (~w2771 & w40521) | (w40520 & w40521);
assign w15099 = ~w15096 & ~w15097;
assign w15100 = ~w15098 & ~w15099;
assign w15101 = w15090 & ~w15100;
assign w15102 = w15090 & ~w15101;
assign w15103 = ~w15090 & ~w15100;
assign w15104 = (~w14700 & w14703) | (~w14700 & w30347) | (w14703 & w30347);
assign w15105 = ~w15102 & w30348;
assign w15106 = (~w15104 & w15102) | (~w15104 & w30349) | (w15102 & w30349);
assign w15107 = ~w15105 & ~w15106;
assign w15108 = b_31 & w5196;
assign w15109 = w5459 & w30350;
assign w15110 = b_30 & w5191;
assign w15111 = ~w15109 & ~w15110;
assign w15112 = ~w15108 & w15111;
assign w15113 = (w15112 & ~w3345) | (w15112 & w30351) | (~w3345 & w30351);
assign w15114 = (w3345 & w40522) | (w3345 & w40523) | (w40522 & w40523);
assign w15115 = (~w3345 & w40524) | (~w3345 & w40525) | (w40524 & w40525);
assign w15116 = ~w15113 & ~w15114;
assign w15117 = ~w15115 & ~w15116;
assign w15118 = ~w15107 & w15117;
assign w15119 = w15107 & ~w15117;
assign w15120 = ~w15118 & ~w15119;
assign w15121 = ~w14722 & w15120;
assign w15122 = w14722 & ~w15120;
assign w15123 = ~w15121 & ~w15122;
assign w15124 = ~w14977 & w15123;
assign w15125 = w14977 & ~w15123;
assign w15126 = ~w15124 & ~w15125;
assign w15127 = (~w30317 & w40526) | (~w30317 & w40527) | (w40526 & w40527);
assign w15128 = (w30317 & w40528) | (w30317 & w40529) | (w40528 & w40529);
assign w15129 = ~w15127 & ~w15128;
assign w15130 = ~w14966 & w15129;
assign w15131 = ~w15129 & ~w14966;
assign w15132 = w15129 & ~w15130;
assign w15133 = ~w15131 & ~w15132;
assign w15134 = w14956 & ~w15133;
assign w15135 = w14956 & ~w15134;
assign w15136 = ~w14956 & ~w15133;
assign w15137 = ~w15135 & ~w15136;
assign w15138 = (w15137 & w14943) | (w15137 & w30352) | (w14943 & w30352);
assign w15139 = ~w14943 & w30353;
assign w15140 = ~w15138 & ~w15139;
assign w15141 = w14930 & ~w15140;
assign w15142 = w14930 & ~w15141;
assign w15143 = ~w14930 & ~w15140;
assign w15144 = ~w15142 & ~w15143;
assign w15145 = ~w14917 & w15144;
assign w15146 = w14917 & ~w15144;
assign w15147 = ~w15145 & ~w15146;
assign w15148 = w14902 & ~w15147;
assign w15149 = w14902 & ~w15148;
assign w15150 = ~w14902 & ~w15147;
assign w15151 = ~w15149 & ~w15150;
assign w15152 = w14888 & ~w15151;
assign w15153 = ~w14888 & w15151;
assign w15154 = w14874 & w27581;
assign w15155 = w14874 & ~w15154;
assign w15156 = w27581 & ~w14874;
assign w15157 = ~w15155 & ~w15156;
assign w15158 = w14862 & ~w15157;
assign w15159 = ~w14862 & w15157;
assign w15160 = w14848 & w30354;
assign w15161 = w14848 & ~w15160;
assign w15162 = w30354 & ~w14848;
assign w15163 = ~w15161 & ~w15162;
assign w15164 = (~w14500 & w14503) | (~w14500 & w30355) | (w14503 & w30355);
assign w15165 = ~w15163 & ~w15164;
assign w15166 = w15164 & ~w15163;
assign w15167 = ~w15164 & ~w15165;
assign w15168 = ~w15166 & ~w15167;
assign w15169 = (~w15168 & w14835) | (~w15168 & w25146) | (w14835 & w25146);
assign w15170 = ~w14835 & w30356;
assign w15171 = ~w15169 & ~w15170;
assign w15172 = (~w14846 & ~w14848) | (~w14846 & w30358) | (~w14848 & w30358);
assign w15173 = (~w14861 & ~w14862) | (~w14861 & w30359) | (~w14862 & w30359);
assign w15174 = w266 & w30360;
assign w15175 = (~w15174 & ~w12670) | (~w15174 & w30361) | (~w12670 & w30361);
assign w15176 = (w12670 & w40530) | (w12670 & w40531) | (w40530 & w40531);
assign w15177 = (~w12670 & w40532) | (~w12670 & w40533) | (w40532 & w40533);
assign w15178 = ~w15175 & ~w15176;
assign w15179 = ~w15177 & ~w15178;
assign w15180 = ~w15173 & ~w15179;
assign w15181 = ~w15173 & ~w15180;
assign w15182 = w15173 & ~w15179;
assign w15183 = b_56 & w986;
assign w15184 = w1069 & w30362;
assign w15185 = b_55 & w981;
assign w15186 = ~w15184 & ~w15185;
assign w15187 = ~w15183 & w15186;
assign w15188 = (w15187 & ~w9798) | (w15187 & w25973) | (~w9798 & w25973);
assign w15189 = (w9798 & w26353) | (w9798 & w26354) | (w26353 & w26354);
assign w15190 = (~w9798 & w27806) | (~w9798 & w27807) | (w27806 & w27807);
assign w15191 = ~w15188 & ~w15189;
assign w15192 = ~w15190 & ~w15191;
assign w15193 = (~w14901 & ~w14902) | (~w14901 & w30363) | (~w14902 & w30363);
assign w15194 = (~w14902 & w40534) | (~w14902 & w40535) | (w40534 & w40535);
assign w15195 = (w14902 & w40536) | (w14902 & w40537) | (w40536 & w40537);
assign w15196 = ~w15194 & ~w15195;
assign w15197 = b_50 & w1694;
assign w15198 = w1834 & w30364;
assign w15199 = b_49 & w1689;
assign w15200 = ~w15198 & ~w15199;
assign w15201 = ~w15197 & w15200;
assign w15202 = (w15201 & ~w8162) | (w15201 & w26355) | (~w8162 & w26355);
assign w15203 = (w8162 & w27582) | (w8162 & w27583) | (w27582 & w27583);
assign w15204 = (~w8162 & w27808) | (~w8162 & w27809) | (w27808 & w27809);
assign w15205 = ~w15202 & ~w15203;
assign w15206 = ~w15204 & ~w15205;
assign w15207 = (~w14928 & ~w14930) | (~w14928 & w30365) | (~w14930 & w30365);
assign w15208 = w15206 & w15207;
assign w15209 = ~w15206 & ~w15207;
assign w15210 = ~w15208 & ~w15209;
assign w15211 = b_47 & w2158;
assign w15212 = w2294 & w30366;
assign w15213 = b_46 & w2153;
assign w15214 = ~w15212 & ~w15213;
assign w15215 = ~w15211 & w15214;
assign w15216 = (w15215 & ~w6998) | (w15215 & w25974) | (~w6998 & w25974);
assign w15217 = (w6998 & w26356) | (w6998 & w26357) | (w26356 & w26357);
assign w15218 = (~w6998 & w26679) | (~w6998 & w26680) | (w26679 & w26680);
assign w15219 = ~w15216 & ~w15217;
assign w15220 = ~w15218 & ~w15219;
assign w15221 = (~w15137 & w14943) | (~w15137 & w30367) | (w14943 & w30367);
assign w15222 = ~w14942 & ~w15221;
assign w15223 = (~w15220 & w15221) | (~w15220 & w30368) | (w15221 & w30368);
assign w15224 = ~w15221 & w30369;
assign w15225 = (w15220 & w15221) | (w15220 & w30370) | (w15221 & w30370);
assign w15226 = ~w15224 & ~w15225;
assign w15227 = b_41 & w3195;
assign w15228 = w3388 & w30371;
assign w15229 = b_40 & w3190;
assign w15230 = ~w15228 & ~w15229;
assign w15231 = ~w15227 & w15230;
assign w15232 = (w15231 & ~w5609) | (w15231 & w25653) | (~w5609 & w25653);
assign w15233 = (w5609 & w25975) | (w5609 & w25976) | (w25975 & w25976);
assign w15234 = (~w5609 & w26358) | (~w5609 & w26359) | (w26358 & w26359);
assign w15235 = ~w15232 & ~w15233;
assign w15236 = (~w15127 & ~w15129) | (~w15127 & w30372) | (~w15129 & w30372);
assign w15237 = w15236 & w30373;
assign w15238 = (~w15236 & w15235) | (~w15236 & w26360) | (w15235 & w26360);
assign w15239 = ~w15237 & ~w15238;
assign w15240 = b_35 & w4499;
assign w15241 = w4723 & w30374;
assign w15242 = b_34 & w4494;
assign w15243 = ~w15241 & ~w15242;
assign w15244 = ~w15240 & w15243;
assign w15245 = (w15244 & ~w4181) | (w15244 & w30375) | (~w4181 & w30375);
assign w15246 = (w4181 & w40538) | (w4181 & w40539) | (w40538 & w40539);
assign w15247 = (~w4181 & w40540) | (~w4181 & w40541) | (w40540 & w40541);
assign w15248 = ~w15245 & ~w15246;
assign w15249 = ~w15247 & ~w15248;
assign w15250 = b_26 & w6761;
assign w15251 = w7075 & w30376;
assign w15252 = b_25 & w6756;
assign w15253 = ~w15251 & ~w15252;
assign w15254 = ~w15250 & w15253;
assign w15255 = (w15254 & ~w2416) | (w15254 & w30377) | (~w2416 & w30377);
assign w15256 = (w2416 & w40542) | (w2416 & w40543) | (w40542 & w40543);
assign w15257 = (~w2416 & w40544) | (~w2416 & w40545) | (w40544 & w40545);
assign w15258 = ~w15255 & ~w15256;
assign w15259 = ~w15257 & ~w15258;
assign w15260 = (~w15053 & ~w15054) | (~w15053 & w30378) | (~w15054 & w30378);
assign w15261 = b_23 & w7613;
assign w15262 = w7941 & w30379;
assign w15263 = b_22 & w7608;
assign w15264 = ~w15262 & ~w15263;
assign w15265 = ~w15261 & w15264;
assign w15266 = (w15265 & ~w1933) | (w15265 & w30380) | (~w1933 & w30380);
assign w15267 = (w1933 & w40546) | (w1933 & w40547) | (w40546 & w40547);
assign w15268 = (~w1933 & w40548) | (~w1933 & w40549) | (w40548 & w40549);
assign w15269 = ~w15266 & ~w15267;
assign w15270 = ~w15268 & ~w15269;
assign w15271 = (~w15035 & ~w15036) | (~w15035 & w30381) | (~w15036 & w30381);
assign w15272 = (~w14998 & ~w15000) | (~w14998 & w30382) | (~w15000 & w30382);
assign w15273 = (~w30328 & w40550) | (~w30328 & w40551) | (w40550 & w40551);
assign w15274 = w12380 & w30383;
assign w15275 = b_8 & ~w12380;
assign w15276 = ~w15274 & ~w15275;
assign w15277 = w14983 & ~w15276;
assign w15278 = ~w14983 & w15276;
assign w15279 = (w30328 & w40552) | (w30328 & w40553) | (w40552 & w40553);
assign w15280 = ~w15273 & ~w15279;
assign w15281 = (~w30328 & w40554) | (~w30328 & w40555) | (w40554 & w40555);
assign w15282 = b_11 & w11620;
assign w15283 = w11969 & w30389;
assign w15284 = b_10 & w11615;
assign w15285 = ~w15283 & ~w15284;
assign w15286 = ~w15282 & w15285;
assign w15287 = (w15286 & ~w530) | (w15286 & w30390) | (~w530 & w30390);
assign w15288 = (w530 & w40556) | (w530 & w40557) | (w40556 & w40557);
assign w15289 = (~w530 & w40558) | (~w530 & w40559) | (w40558 & w40559);
assign w15290 = ~w15287 & ~w15288;
assign w15291 = ~w15289 & ~w15290;
assign w15292 = (w15291 & w15280) | (w15291 & w30391) | (w15280 & w30391);
assign w15293 = ~w15280 & w30392;
assign w15294 = ~w15292 & ~w15293;
assign w15295 = b_14 & w10562;
assign w15296 = w10902 & w30393;
assign w15297 = b_13 & w10557;
assign w15298 = ~w15296 & ~w15297;
assign w15299 = ~w15295 & w15298;
assign w15300 = (w15299 & ~w735) | (w15299 & w30394) | (~w735 & w30394);
assign w15301 = (w735 & w40560) | (w735 & w40561) | (w40560 & w40561);
assign w15302 = (~w735 & w40562) | (~w735 & w40563) | (w40562 & w40563);
assign w15303 = ~w15300 & ~w15301;
assign w15304 = ~w15302 & ~w15303;
assign w15305 = ~w15294 & ~w15304;
assign w15306 = w15294 & w15304;
assign w15307 = ~w15305 & ~w15306;
assign w15308 = w15272 & ~w15307;
assign w15309 = ~w15272 & w15307;
assign w15310 = ~w15308 & ~w15309;
assign w15311 = b_17 & w9534;
assign w15312 = w9876 & w30395;
assign w15313 = b_16 & w9529;
assign w15314 = ~w15312 & ~w15313;
assign w15315 = ~w15311 & w15314;
assign w15316 = (w15315 & ~w1038) | (w15315 & w30396) | (~w1038 & w30396);
assign w15317 = (w1038 & w40564) | (w1038 & w40565) | (w40564 & w40565);
assign w15318 = (~w1038 & w40566) | (~w1038 & w40567) | (w40566 & w40567);
assign w15319 = ~w15316 & ~w15317;
assign w15320 = ~w15318 & ~w15319;
assign w15321 = w15310 & ~w15320;
assign w15322 = w15310 & ~w15321;
assign w15323 = ~w15310 & ~w15320;
assign w15324 = ~w15322 & ~w15323;
assign w15325 = (~w15017 & ~w15018) | (~w15017 & w30397) | (~w15018 & w30397);
assign w15326 = w15324 & w15325;
assign w15327 = ~w15324 & ~w15325;
assign w15328 = ~w15326 & ~w15327;
assign w15329 = b_20 & w8526;
assign w15330 = w8886 & w30398;
assign w15331 = b_19 & w8521;
assign w15332 = ~w15330 & ~w15331;
assign w15333 = ~w15329 & w15332;
assign w15334 = (w15333 & ~w1503) | (w15333 & w30399) | (~w1503 & w30399);
assign w15335 = (w1503 & w40568) | (w1503 & w40569) | (w40568 & w40569);
assign w15336 = (~w1503 & w40570) | (~w1503 & w40571) | (w40570 & w40571);
assign w15337 = ~w15334 & ~w15335;
assign w15338 = ~w15336 & ~w15337;
assign w15339 = ~w15328 & w15338;
assign w15340 = w15328 & ~w15338;
assign w15341 = ~w15339 & ~w15340;
assign w15342 = ~w15271 & w15341;
assign w15343 = ~w15271 & ~w15342;
assign w15344 = w15271 & w15341;
assign w15345 = (~w15270 & w15343) | (~w15270 & w30400) | (w15343 & w30400);
assign w15346 = (w15270 & ~w15271) | (w15270 & w40572) | (~w15271 & w40572);
assign w15347 = ~w15343 & w15346;
assign w15348 = ~w15345 & ~w15347;
assign w15349 = ~w15260 & w15348;
assign w15350 = w15260 & ~w15348;
assign w15351 = ~w15349 & ~w15350;
assign w15352 = ~w15259 & w15351;
assign w15353 = w15351 & ~w15352;
assign w15354 = ~w15351 & ~w15259;
assign w15355 = ~w15353 & ~w15354;
assign w15356 = (~w15072 & ~w15073) | (~w15072 & w30401) | (~w15073 & w30401);
assign w15357 = w15355 & w15356;
assign w15358 = ~w15355 & ~w15356;
assign w15359 = ~w15357 & ~w15358;
assign w15360 = b_29 & w5962;
assign w15361 = w6246 & w30402;
assign w15362 = b_28 & w5957;
assign w15363 = ~w15361 & ~w15362;
assign w15364 = ~w15360 & w15363;
assign w15365 = (w15364 & ~w2954) | (w15364 & w30403) | (~w2954 & w30403);
assign w15366 = (w2954 & w40573) | (w2954 & w40574) | (w40573 & w40574);
assign w15367 = (~w2954 & w40575) | (~w2954 & w40576) | (w40575 & w40576);
assign w15368 = ~w15365 & ~w15366;
assign w15369 = ~w15367 & ~w15368;
assign w15370 = w15359 & ~w15369;
assign w15371 = w15359 & ~w15370;
assign w15372 = ~w15359 & ~w15369;
assign w15373 = ~w15371 & ~w15372;
assign w15374 = (~w15089 & ~w15090) | (~w15089 & w30404) | (~w15090 & w30404);
assign w15375 = w15373 & w15374;
assign w15376 = ~w15373 & ~w15374;
assign w15377 = ~w15375 & ~w15376;
assign w15378 = b_32 & w5196;
assign w15379 = w5459 & w30405;
assign w15380 = b_31 & w5191;
assign w15381 = ~w15379 & ~w15380;
assign w15382 = ~w15378 & w15381;
assign w15383 = (w15382 & ~w3545) | (w15382 & w30406) | (~w3545 & w30406);
assign w15384 = (w3545 & w40577) | (w3545 & w40578) | (w40577 & w40578);
assign w15385 = (~w3545 & w40579) | (~w3545 & w40580) | (w40579 & w40580);
assign w15386 = ~w15383 & ~w15384;
assign w15387 = ~w15385 & ~w15386;
assign w15388 = ~w15377 & w15387;
assign w15389 = w15377 & ~w15387;
assign w15390 = ~w15388 & ~w15389;
assign w15391 = (~w15106 & ~w15107) | (~w15106 & w30407) | (~w15107 & w30407);
assign w15392 = w15390 & ~w15391;
assign w15393 = ~w15390 & w15391;
assign w15394 = ~w15392 & ~w15393;
assign w15395 = ~w15249 & w15394;
assign w15396 = w15394 & ~w15395;
assign w15397 = ~w15394 & ~w15249;
assign w15398 = (~w15121 & ~w15123) | (~w15121 & w30408) | (~w15123 & w30408);
assign w15399 = ~w15396 & w30409;
assign w15400 = (~w15398 & w15396) | (~w15398 & w30410) | (w15396 & w30410);
assign w15401 = ~w15399 & ~w15400;
assign w15402 = b_38 & w3803;
assign w15403 = w4027 & w30411;
assign w15404 = b_37 & w3798;
assign w15405 = ~w15403 & ~w15404;
assign w15406 = ~w15402 & w15405;
assign w15407 = (w15406 & ~w4658) | (w15406 & w30412) | (~w4658 & w30412);
assign w15408 = (w4658 & w40581) | (w4658 & w40582) | (w40581 & w40582);
assign w15409 = (~w4658 & w40583) | (~w4658 & w40584) | (w40583 & w40584);
assign w15410 = ~w15407 & ~w15408;
assign w15411 = ~w15409 & ~w15410;
assign w15412 = w15401 & ~w15411;
assign w15413 = ~w15401 & w15411;
assign w15414 = ~w15238 & w30413;
assign w15415 = ~w15238 & w40585;
assign w15416 = w15239 & ~w15415;
assign w15417 = (w15238 & w40586) | (w15238 & w40587) | (w40586 & w40587);
assign w15418 = ~w15416 & ~w15417;
assign w15419 = (~w14955 & ~w14956) | (~w14955 & w30417) | (~w14956 & w30417);
assign w15420 = b_44 & w2639;
assign w15421 = w2820 & w30418;
assign w15422 = b_43 & w2634;
assign w15423 = ~w15421 & ~w15422;
assign w15424 = ~w15420 & w15423;
assign w15425 = w15423 & w30419;
assign w15426 = (~w6408 & w25654) | (~w6408 & w25655) | (w25654 & w25655);
assign w15427 = (w6408 & w25656) | (w6408 & w25657) | (w25656 & w25657);
assign w15428 = ~w15426 & ~w15427;
assign w15429 = ~w15419 & ~w15428;
assign w15430 = w15428 & ~w15419;
assign w15431 = w15419 & ~w15428;
assign w15432 = ~w15430 & ~w15431;
assign w15433 = ~w15418 & ~w15432;
assign w15434 = w15432 & ~w15418;
assign w15435 = ~w15432 & ~w15433;
assign w15436 = ~w15434 & ~w15435;
assign w15437 = (w27763 & w30420) | (w27763 & w30421) | (w30420 & w30421);
assign w15438 = ~w15226 & ~w15437;
assign w15439 = ~w26681 & w30422;
assign w15440 = ~w15438 & ~w15439;
assign w15441 = ~w15210 & w15440;
assign w15442 = w15210 & ~w15440;
assign w15443 = ~w15441 & ~w15442;
assign w15444 = (~w26361 & w30423) | (~w26361 & w30424) | (w30423 & w30424);
assign w15445 = b_53 & w1295;
assign w15446 = w1422 & w30425;
assign w15447 = b_52 & w1290;
assign w15448 = ~w15446 & ~w15447;
assign w15449 = ~w15445 & w15448;
assign w15450 = w15448 & w30426;
assign w15451 = (w9109 & w40588) | (w9109 & w40589) | (w40588 & w40589);
assign w15452 = (~w9109 & w40590) | (~w9109 & w40591) | (w40590 & w40591);
assign w15453 = ~w15451 & ~w15452;
assign w15454 = ~w15444 & ~w15453;
assign w15455 = ~w15444 & ~w15454;
assign w15456 = w15444 & ~w15453;
assign w15457 = ~w15455 & ~w15456;
assign w15458 = (w15443 & w15455) | (w15443 & w27584) | (w15455 & w27584);
assign w15459 = w15443 & ~w15458;
assign w15460 = ~w15457 & ~w15458;
assign w15461 = ~w15459 & ~w15460;
assign w15462 = w15196 & ~w15461;
assign w15463 = w15196 & ~w15462;
assign w15464 = ~w15196 & ~w15461;
assign w15465 = ~w15463 & ~w15464;
assign w15466 = b_59 & w657;
assign w15467 = w754 & w30431;
assign w15468 = b_58 & w652;
assign w15469 = ~w15467 & ~w15468;
assign w15470 = ~w15466 & w15469;
assign w15471 = (w15470 & ~w27585) | (w15470 & w30432) | (~w27585 & w30432);
assign w15472 = a_14 & ~w15471;
assign w15473 = w15471 & a_14;
assign w15474 = ~w15471 & ~w15472;
assign w15475 = ~w15473 & ~w15474;
assign w15476 = (~w14887 & ~w14888) | (~w14887 & w30433) | (~w14888 & w30433);
assign w15477 = ~w15475 & ~w15476;
assign w15478 = w15476 & ~w15475;
assign w15479 = ~w15476 & ~w15477;
assign w15480 = ~w15479 & w30434;
assign w15481 = (w15465 & w15479) | (w15465 & w30435) | (w15479 & w30435);
assign w15482 = ~w15480 & ~w15481;
assign w15483 = (~w14872 & ~w14874) | (~w14872 & w30436) | (~w14874 & w30436);
assign w15484 = b_62 & w418;
assign w15485 = w481 & w30437;
assign w15486 = b_61 & w413;
assign w15487 = ~w15485 & ~w15486;
assign w15488 = ~w15484 & w15487;
assign w15489 = w15487 & w30438;
assign w15490 = (~w12273 & w40592) | (~w12273 & w40593) | (w40592 & w40593);
assign w15491 = (w12273 & w30440) | (w12273 & w30441) | (w30440 & w30441);
assign w15492 = ~w15490 & ~w15491;
assign w15493 = ~w15483 & ~w15492;
assign w15494 = ~w15483 & ~w15493;
assign w15495 = w15483 & ~w15492;
assign w15496 = (~w15482 & w15494) | (~w15482 & w30442) | (w15494 & w30442);
assign w15497 = w15482 & ~w15495;
assign w15498 = ~w15494 & w15497;
assign w15499 = ~w15496 & ~w15498;
assign w15500 = (w15499 & w15181) | (w15499 & w30443) | (w15181 & w30443);
assign w15501 = ~w15181 & w30444;
assign w15502 = ~w15500 & ~w15501;
assign w15503 = ~w15172 & w15502;
assign w15504 = ~w15172 & ~w15503;
assign w15505 = w15172 & w15502;
assign w15506 = ~w15504 & ~w15505;
assign w15507 = (w14835 & w30445) | (w14835 & w30446) | (w30445 & w30446);
assign w15508 = (w13761 & w37676) | (w13761 & w37677) | (w37676 & w37677);
assign w15509 = ~w15507 & ~w15508;
assign w15510 = ~w15180 & ~w15500;
assign w15511 = ~w15493 & ~w15496;
assign w15512 = b_63 & w418;
assign w15513 = w481 & w30450;
assign w15514 = b_62 & w413;
assign w15515 = ~w15513 & ~w15514;
assign w15516 = ~w15512 & w15515;
assign w15517 = (w15516 & ~w12646) | (w15516 & w30451) | (~w12646 & w30451);
assign w15518 = (w12646 & w40594) | (w12646 & w40595) | (w40594 & w40595);
assign w15519 = (~w12646 & w40596) | (~w12646 & w40597) | (w40596 & w40597);
assign w15520 = ~w15517 & ~w15518;
assign w15521 = ~w15519 & ~w15520;
assign w15522 = (~w15521 & w15496) | (~w15521 & w30452) | (w15496 & w30452);
assign w15523 = ~w15511 & ~w15522;
assign w15524 = ~w15496 & w30453;
assign w15525 = (~w15465 & w15479) | (~w15465 & w30454) | (w15479 & w30454);
assign w15526 = b_60 & w657;
assign w15527 = w754 & w30455;
assign w15528 = b_59 & w652;
assign w15529 = ~w15527 & ~w15528;
assign w15530 = ~w15526 & w15529;
assign w15531 = (w15530 & ~w11196) | (w15530 & w30456) | (~w11196 & w30456);
assign w15532 = (w11196 & w40598) | (w11196 & w40599) | (w40598 & w40599);
assign w15533 = (~w11196 & w40600) | (~w11196 & w40601) | (w40600 & w40601);
assign w15534 = ~w15531 & ~w15532;
assign w15535 = ~w15533 & ~w15534;
assign w15536 = (w15535 & w15525) | (w15535 & w30457) | (w15525 & w30457);
assign w15537 = ~w15525 & w30458;
assign w15538 = ~w15536 & ~w15537;
assign w15539 = b_57 & w986;
assign w15540 = w1069 & w30459;
assign w15541 = b_56 & w981;
assign w15542 = ~w15540 & ~w15541;
assign w15543 = ~w15539 & w15542;
assign w15544 = (w15543 & ~w10452) | (w15543 & w30460) | (~w10452 & w30460);
assign w15545 = (w10452 & w40602) | (w10452 & w40603) | (w40602 & w40603);
assign w15546 = (~w10452 & w40604) | (~w10452 & w40605) | (w40604 & w40605);
assign w15547 = ~w15544 & ~w15545;
assign w15548 = ~w15546 & ~w15547;
assign w15549 = (~w15195 & ~w15196) | (~w15195 & w27810) | (~w15196 & w27810);
assign w15550 = w15548 & w15549;
assign w15551 = ~w15548 & ~w15549;
assign w15552 = ~w15550 & ~w15551;
assign w15553 = ~w15454 & ~w15458;
assign w15554 = b_54 & w1295;
assign w15555 = w1422 & w30461;
assign w15556 = b_53 & w1290;
assign w15557 = ~w15555 & ~w15556;
assign w15558 = ~w15554 & w15557;
assign w15559 = (w15558 & ~w9134) | (w15558 & w30462) | (~w9134 & w30462);
assign w15560 = (w9134 & w40606) | (w9134 & w40607) | (w40606 & w40607);
assign w15561 = (~w9134 & w40608) | (~w9134 & w40609) | (w40608 & w40609);
assign w15562 = ~w15559 & ~w15560;
assign w15563 = ~w15561 & ~w15562;
assign w15564 = (~w15563 & w15458) | (~w15563 & w30463) | (w15458 & w30463);
assign w15565 = ~w15553 & ~w15564;
assign w15566 = ~w15458 & w30464;
assign w15567 = ~w15565 & ~w15566;
assign w15568 = b_48 & w2158;
assign w15569 = w2294 & w30465;
assign w15570 = b_47 & w2153;
assign w15571 = ~w15569 & ~w15570;
assign w15572 = ~w15568 & w15571;
assign w15573 = (w15572 & ~w7284) | (w15572 & w30466) | (~w7284 & w30466);
assign w15574 = (w7284 & w40610) | (w7284 & w40611) | (w40610 & w40611);
assign w15575 = (~w7284 & w40612) | (~w7284 & w40613) | (w40612 & w40613);
assign w15576 = ~w15573 & ~w15574;
assign w15577 = ~w15575 & ~w15576;
assign w15578 = (~w26681 & w30467) | (~w26681 & w30468) | (w30467 & w30468);
assign w15579 = w15577 & w15578;
assign w15580 = ~w15577 & ~w15578;
assign w15581 = ~w15579 & ~w15580;
assign w15582 = (~w15429 & w15432) | (~w15429 & w25977) | (w15432 & w25977);
assign w15583 = b_45 & w2639;
assign w15584 = w2820 & w30469;
assign w15585 = b_44 & w2634;
assign w15586 = ~w15584 & ~w15585;
assign w15587 = ~w15583 & w15586;
assign w15588 = (w15587 & ~w6682) | (w15587 & w25978) | (~w6682 & w25978);
assign w15589 = (w6682 & w26363) | (w6682 & w26364) | (w26363 & w26364);
assign w15590 = (~w6682 & w30470) | (~w6682 & w30471) | (w30470 & w30471);
assign w15591 = ~w15588 & ~w15589;
assign w15592 = ~w15590 & ~w15591;
assign w15593 = (~w25977 & w30472) | (~w25977 & w30473) | (w30472 & w30473);
assign w15594 = ~w15582 & ~w15593;
assign w15595 = (w25977 & w30474) | (w25977 & w30475) | (w30474 & w30475);
assign w15596 = ~w15594 & ~w15595;
assign w15597 = (~w15238 & ~w15414) | (~w15238 & w30476) | (~w15414 & w30476);
assign w15598 = b_42 & w3195;
assign w15599 = w3388 & w30477;
assign w15600 = b_41 & w3190;
assign w15601 = ~w15599 & ~w15600;
assign w15602 = ~w15598 & w15601;
assign w15603 = (w15602 & ~w5864) | (w15602 & w30478) | (~w5864 & w30478);
assign w15604 = (w5864 & w40614) | (w5864 & w40615) | (w40614 & w40615);
assign w15605 = (~w5864 & w40616) | (~w5864 & w40617) | (w40616 & w40617);
assign w15606 = ~w15603 & ~w15604;
assign w15607 = ~w15605 & ~w15606;
assign w15608 = (w15414 & w40618) | (w15414 & w40619) | (w40618 & w40619);
assign w15609 = ~w15597 & ~w15608;
assign w15610 = (~w15414 & w40620) | (~w15414 & w40621) | (w40620 & w40621);
assign w15611 = ~w15609 & ~w15610;
assign w15612 = (~w15392 & ~w15394) | (~w15392 & w30479) | (~w15394 & w30479);
assign w15613 = (~w15376 & ~w15377) | (~w15376 & w30480) | (~w15377 & w30480);
assign w15614 = (~w15358 & ~w15359) | (~w15358 & w30481) | (~w15359 & w30481);
assign w15615 = ~w15342 & ~w15345;
assign w15616 = b_24 & w7613;
assign w15617 = w7941 & w30482;
assign w15618 = b_23 & w7608;
assign w15619 = ~w15617 & ~w15618;
assign w15620 = ~w15616 & w15619;
assign w15621 = (w15620 & ~w2083) | (w15620 & w30483) | (~w2083 & w30483);
assign w15622 = (w2083 & w40622) | (w2083 & w40623) | (w40622 & w40623);
assign w15623 = (~w2083 & w40624) | (~w2083 & w40625) | (w40624 & w40625);
assign w15624 = ~w15621 & ~w15622;
assign w15625 = ~w15623 & ~w15624;
assign w15626 = b_18 & w9534;
assign w15627 = w9876 & w30484;
assign w15628 = b_17 & w9529;
assign w15629 = ~w15627 & ~w15628;
assign w15630 = ~w15626 & w15629;
assign w15631 = (w15630 & ~w1238) | (w15630 & w30485) | (~w1238 & w30485);
assign w15632 = (w1238 & w40626) | (w1238 & w40627) | (w40626 & w40627);
assign w15633 = (~w1238 & w40628) | (~w1238 & w40629) | (w40628 & w40629);
assign w15634 = ~w15631 & ~w15632;
assign w15635 = ~w15633 & ~w15634;
assign w15636 = (~w15291 & w15280) | (~w15291 & w30486) | (w15280 & w30486);
assign w15637 = (~w15636 & w15294) | (~w15636 & w40630) | (w15294 & w40630);
assign w15638 = b_12 & w11620;
assign w15639 = w11969 & w30487;
assign w15640 = b_11 & w11615;
assign w15641 = ~w15639 & ~w15640;
assign w15642 = ~w15638 & w15641;
assign w15643 = (w15642 & ~w552) | (w15642 & w30488) | (~w552 & w30488);
assign w15644 = (w552 & w40631) | (w552 & w40632) | (w40631 & w40632);
assign w15645 = (~w552 & w40633) | (~w552 & w40634) | (w40633 & w40634);
assign w15646 = ~w15643 & ~w15644;
assign w15647 = ~w15645 & ~w15646;
assign w15648 = w12380 & w30489;
assign w15649 = b_9 & ~w12380;
assign w15650 = ~w15648 & ~w15649;
assign w15651 = a_8 & ~w15276;
assign w15652 = ~a_8 & w15276;
assign w15653 = ~w15651 & ~w15652;
assign w15654 = ~w15650 & ~w15653;
assign w15655 = w15650 & w15653;
assign w15656 = ~w15654 & ~w15655;
assign w15657 = (w30328 & w40635) | (w30328 & w40636) | (w40635 & w40636);
assign w15658 = (~w30328 & w40637) | (~w30328 & w40638) | (w40637 & w40638);
assign w15659 = ~w15657 & ~w15658;
assign w15660 = w15647 & w15659;
assign w15661 = ~w15647 & ~w15659;
assign w15662 = ~w15660 & ~w15661;
assign w15663 = b_15 & w10562;
assign w15664 = w10902 & w30494;
assign w15665 = b_14 & w10557;
assign w15666 = ~w15664 & ~w15665;
assign w15667 = ~w15663 & w15666;
assign w15668 = (w15667 & ~w827) | (w15667 & w30495) | (~w827 & w30495);
assign w15669 = (w827 & w40639) | (w827 & w40640) | (w40639 & w40640);
assign w15670 = (~w827 & w40641) | (~w827 & w40642) | (w40641 & w40642);
assign w15671 = ~w15668 & ~w15669;
assign w15672 = ~w15670 & ~w15671;
assign w15673 = ~w15662 & ~w15672;
assign w15674 = w15662 & w15672;
assign w15675 = ~w15673 & ~w15674;
assign w15676 = ~w15637 & w15675;
assign w15677 = w15637 & ~w15675;
assign w15678 = ~w15676 & ~w15677;
assign w15679 = ~w15635 & w15678;
assign w15680 = w15678 & ~w15679;
assign w15681 = ~w15678 & ~w15635;
assign w15682 = (~w15309 & ~w15310) | (~w15309 & w30496) | (~w15310 & w30496);
assign w15683 = ~w15680 & w30497;
assign w15684 = (~w15682 & w15680) | (~w15682 & w30498) | (w15680 & w30498);
assign w15685 = ~w15683 & ~w15684;
assign w15686 = b_21 & w8526;
assign w15687 = w8886 & w30499;
assign w15688 = b_20 & w8521;
assign w15689 = ~w15687 & ~w15688;
assign w15690 = ~w15686 & w15689;
assign w15691 = (w15690 & ~w1634) | (w15690 & w30500) | (~w1634 & w30500);
assign w15692 = (w1634 & w40643) | (w1634 & w40644) | (w40643 & w40644);
assign w15693 = (~w1634 & w40645) | (~w1634 & w40646) | (w40645 & w40646);
assign w15694 = ~w15691 & ~w15692;
assign w15695 = ~w15693 & ~w15694;
assign w15696 = w15685 & ~w15695;
assign w15697 = w15685 & ~w15696;
assign w15698 = ~w15685 & ~w15695;
assign w15699 = ~w15697 & ~w15698;
assign w15700 = (~w15327 & ~w15328) | (~w15327 & w30501) | (~w15328 & w30501);
assign w15701 = ~w15699 & ~w15700;
assign w15702 = w15699 & w15700;
assign w15703 = ~w15701 & ~w15702;
assign w15704 = ~w15625 & w15703;
assign w15705 = ~w15703 & ~w15625;
assign w15706 = w15703 & ~w15704;
assign w15707 = ~w15705 & ~w15706;
assign w15708 = ~w15615 & ~w15707;
assign w15709 = ~w15615 & ~w15708;
assign w15710 = ~w15707 & ~w15708;
assign w15711 = ~w15709 & ~w15710;
assign w15712 = b_27 & w6761;
assign w15713 = w7075 & w30502;
assign w15714 = b_26 & w6756;
assign w15715 = ~w15713 & ~w15714;
assign w15716 = ~w15712 & w15715;
assign w15717 = (w15716 & ~w2582) | (w15716 & w30503) | (~w2582 & w30503);
assign w15718 = (w2582 & w40647) | (w2582 & w40648) | (w40647 & w40648);
assign w15719 = (~w2582 & w40649) | (~w2582 & w40650) | (w40649 & w40650);
assign w15720 = ~w15717 & ~w15718;
assign w15721 = ~w15719 & ~w15720;
assign w15722 = ~w15711 & ~w15721;
assign w15723 = ~w15711 & ~w15722;
assign w15724 = w15711 & ~w15721;
assign w15725 = (~w15349 & ~w15351) | (~w15349 & w30504) | (~w15351 & w30504);
assign w15726 = ~w15723 & w30505;
assign w15727 = (~w15725 & w15723) | (~w15725 & w30506) | (w15723 & w30506);
assign w15728 = ~w15726 & ~w15727;
assign w15729 = b_30 & w5962;
assign w15730 = w6246 & w30507;
assign w15731 = b_29 & w5957;
assign w15732 = ~w15730 & ~w15731;
assign w15733 = ~w15729 & w15732;
assign w15734 = (w15733 & ~w3138) | (w15733 & w30508) | (~w3138 & w30508);
assign w15735 = (w3138 & w40651) | (w3138 & w40652) | (w40651 & w40652);
assign w15736 = (~w3138 & w40653) | (~w3138 & w40654) | (w40653 & w40654);
assign w15737 = ~w15734 & ~w15735;
assign w15738 = ~w15736 & ~w15737;
assign w15739 = w15728 & ~w15738;
assign w15740 = ~w15728 & w15738;
assign w15741 = ~w15614 & w30509;
assign w15742 = ~w15614 & ~w15741;
assign w15743 = ~w15739 & ~w15741;
assign w15744 = ~w15741 & w30509;
assign w15745 = ~w15742 & ~w15744;
assign w15746 = b_33 & w5196;
assign w15747 = w5459 & w30510;
assign w15748 = b_32 & w5191;
assign w15749 = ~w15747 & ~w15748;
assign w15750 = ~w15746 & w15749;
assign w15751 = (w15750 & ~w3744) | (w15750 & w30511) | (~w3744 & w30511);
assign w15752 = (w3744 & w40655) | (w3744 & w40656) | (w40655 & w40656);
assign w15753 = (~w3744 & w40657) | (~w3744 & w40658) | (w40657 & w40658);
assign w15754 = ~w15751 & ~w15752;
assign w15755 = ~w15753 & ~w15754;
assign w15756 = ~w15745 & ~w15755;
assign w15757 = ~w15745 & ~w15756;
assign w15758 = w15745 & ~w15755;
assign w15759 = ~w15757 & ~w15758;
assign w15760 = ~w15613 & w15759;
assign w15761 = w15613 & ~w15759;
assign w15762 = ~w15760 & ~w15761;
assign w15763 = b_36 & w4499;
assign w15764 = w4723 & w30512;
assign w15765 = b_35 & w4494;
assign w15766 = ~w15764 & ~w15765;
assign w15767 = ~w15763 & w15766;
assign w15768 = (w15767 & ~w4395) | (w15767 & w30513) | (~w4395 & w30513);
assign w15769 = (w4395 & w40659) | (w4395 & w40660) | (w40659 & w40660);
assign w15770 = (~w4395 & w40661) | (~w4395 & w40662) | (w40661 & w40662);
assign w15771 = ~w15768 & ~w15769;
assign w15772 = ~w15770 & ~w15771;
assign w15773 = ~w15762 & ~w15772;
assign w15774 = w15762 & w15772;
assign w15775 = ~w15773 & ~w15774;
assign w15776 = w15612 & ~w15775;
assign w15777 = ~w15612 & w15775;
assign w15778 = ~w15776 & ~w15777;
assign w15779 = b_39 & w3803;
assign w15780 = w4027 & w30514;
assign w15781 = b_38 & w3798;
assign w15782 = ~w15780 & ~w15781;
assign w15783 = ~w15779 & w15782;
assign w15784 = (w15783 & ~w4888) | (w15783 & w30515) | (~w4888 & w30515);
assign w15785 = (w4888 & w40663) | (w4888 & w40664) | (w40663 & w40664);
assign w15786 = (~w4888 & w40665) | (~w4888 & w40666) | (w40665 & w40666);
assign w15787 = ~w15784 & ~w15785;
assign w15788 = ~w15786 & ~w15787;
assign w15789 = w15778 & ~w15788;
assign w15790 = w15778 & ~w15789;
assign w15791 = ~w15778 & ~w15788;
assign w15792 = ~w15790 & ~w15791;
assign w15793 = (~w15400 & ~w15401) | (~w15400 & w30516) | (~w15401 & w30516);
assign w15794 = (~w15793 & w15790) | (~w15793 & w30517) | (w15790 & w30517);
assign w15795 = ~w15792 & ~w15794;
assign w15796 = ~w30517 & w40667;
assign w15797 = ~w15795 & ~w15796;
assign w15798 = (~w15797 & w15609) | (~w15797 & w30518) | (w15609 & w30518);
assign w15799 = ~w15611 & ~w15798;
assign w15800 = ~w15797 & ~w15798;
assign w15801 = ~w15799 & ~w15800;
assign w15802 = (w15801 & w15594) | (w15801 & w40668) | (w15594 & w40668);
assign w15803 = ~w15594 & w40669;
assign w15804 = ~w15802 & ~w15803;
assign w15805 = w15581 & ~w15804;
assign w15806 = w15581 & ~w15805;
assign w15807 = ~w15581 & ~w15804;
assign w15808 = ~w15806 & ~w15807;
assign w15809 = b_51 & w1694;
assign w15810 = w1834 & w30519;
assign w15811 = b_50 & w1689;
assign w15812 = ~w15810 & ~w15811;
assign w15813 = ~w15809 & w15812;
assign w15814 = (w15813 & ~w8186) | (w15813 & w27812) | (~w8186 & w27812);
assign w15815 = (w8186 & w30520) | (w8186 & w30521) | (w30520 & w30521);
assign w15816 = (~w8186 & w30522) | (~w8186 & w30523) | (w30522 & w30523);
assign w15817 = ~w15814 & ~w15815;
assign w15818 = ~w15816 & ~w15817;
assign w15819 = (~w15209 & ~w15210) | (~w15209 & w30524) | (~w15210 & w30524);
assign w15820 = ~w15818 & ~w15819;
assign w15821 = w15818 & w15819;
assign w15822 = ~w15820 & ~w15821;
assign w15823 = ~w15808 & w15822;
assign w15824 = ~w15822 & ~w15808;
assign w15825 = w15822 & ~w15823;
assign w15826 = ~w15824 & ~w15825;
assign w15827 = (~w15826 & w15565) | (~w15826 & w27813) | (w15565 & w27813);
assign w15828 = ~w15567 & ~w15827;
assign w15829 = ~w15826 & ~w15827;
assign w15830 = ~w15828 & ~w15829;
assign w15831 = w15552 & ~w15830;
assign w15832 = ~w15552 & w15830;
assign w15833 = ~w15538 & ~w15832;
assign w15834 = ~w15538 & w30525;
assign w15835 = ~w15538 & ~w15834;
assign w15836 = w30525 & w15538;
assign w15837 = ~w15835 & ~w15836;
assign w15838 = (w15837 & w15523) | (w15837 & w30526) | (w15523 & w30526);
assign w15839 = ~w15523 & w30527;
assign w15840 = ~w15838 & ~w15839;
assign w15841 = ~w15510 & ~w15840;
assign w15842 = ~w15510 & ~w15841;
assign w15843 = w15510 & ~w15840;
assign w15844 = ~w15842 & ~w15843;
assign w15845 = (w14835 & w27438) | (w14835 & w27439) | (w27438 & w27439);
assign w15846 = (w13761 & w37678) | (w13761 & w37679) | (w37678 & w37679);
assign w15847 = ~w15845 & ~w15846;
assign w15848 = (~w15837 & w15523) | (~w15837 & w30531) | (w15523 & w30531);
assign w15849 = ~w15522 & ~w15848;
assign w15850 = b_61 & w657;
assign w15851 = w754 & w30532;
assign w15852 = b_60 & w652;
assign w15853 = ~w15851 & ~w15852;
assign w15854 = ~w15850 & w15853;
assign w15855 = (w15854 & ~w11901) | (w15854 & w30533) | (~w11901 & w30533);
assign w15856 = (w11901 & w40670) | (w11901 & w40671) | (w40670 & w40671);
assign w15857 = (~w11901 & w40672) | (~w11901 & w40673) | (w40672 & w40673);
assign w15858 = ~w15855 & ~w15856;
assign w15859 = ~w15857 & ~w15858;
assign w15860 = (~w15551 & ~w15552) | (~w15551 & w30534) | (~w15552 & w30534);
assign w15861 = ~w15859 & ~w15860;
assign w15862 = w15860 & ~w15859;
assign w15863 = ~w15860 & ~w15861;
assign w15864 = ~w15862 & ~w15863;
assign w15865 = b_55 & w1295;
assign w15866 = w1422 & w30535;
assign w15867 = b_54 & w1290;
assign w15868 = ~w15866 & ~w15867;
assign w15869 = ~w15865 & w15868;
assign w15870 = (w15869 & ~w9776) | (w15869 & w27814) | (~w9776 & w27814);
assign w15871 = (w9776 & w30536) | (w9776 & w30537) | (w30536 & w30537);
assign w15872 = (~w9776 & w30538) | (~w9776 & w30539) | (w30538 & w30539);
assign w15873 = ~w15870 & ~w15871;
assign w15874 = ~w15872 & ~w15873;
assign w15875 = (~w15822 & w40674) | (~w15822 & w40675) | (w40674 & w40675);
assign w15876 = (w15822 & w40676) | (w15822 & w40677) | (w40676 & w40677);
assign w15877 = ~w15875 & ~w15876;
assign w15878 = b_52 & w1694;
assign w15879 = w1834 & w30544;
assign w15880 = b_51 & w1689;
assign w15881 = ~w15879 & ~w15880;
assign w15882 = ~w15878 & w15881;
assign w15883 = (w15882 & ~w8793) | (w15882 & w30545) | (~w8793 & w30545);
assign w15884 = (w8793 & w40678) | (w8793 & w40679) | (w40678 & w40679);
assign w15885 = (~w8793 & w40680) | (~w8793 & w40681) | (w40680 & w40681);
assign w15886 = ~w15883 & ~w15884;
assign w15887 = ~w15885 & ~w15886;
assign w15888 = (~w15580 & ~w15581) | (~w15580 & w27586) | (~w15581 & w27586);
assign w15889 = (~w15581 & w40682) | (~w15581 & w40683) | (w40682 & w40683);
assign w15890 = (w15581 & w40684) | (w15581 & w40685) | (w40684 & w40685);
assign w15891 = ~w15889 & ~w15890;
assign w15892 = b_49 & w2158;
assign w15893 = w2294 & w30546;
assign w15894 = b_48 & w2153;
assign w15895 = ~w15893 & ~w15894;
assign w15896 = ~w15892 & w15895;
assign w15897 = (w15896 & ~w7859) | (w15896 & w25458) | (~w7859 & w25458);
assign w15898 = (w7859 & w25658) | (w7859 & w25659) | (w25658 & w25659);
assign w15899 = (~w7859 & w25660) | (~w7859 & w25661) | (w25660 & w25661);
assign w15900 = ~w15897 & ~w15898;
assign w15901 = ~w15899 & ~w15900;
assign w15902 = (~w15593 & w15596) | (~w15593 & w25662) | (w15596 & w25662);
assign w15903 = (~w15902 & w15900) | (~w15902 & w25979) | (w15900 & w25979);
assign w15904 = (~w25979 & w30547) | (~w25979 & w30548) | (w30547 & w30548);
assign w15905 = (~w15596 & w40686) | (~w15596 & w40687) | (w40686 & w40687);
assign w15906 = ~w15904 & ~w15905;
assign w15907 = b_43 & w3195;
assign w15908 = w3388 & w30549;
assign w15909 = b_42 & w3190;
assign w15910 = ~w15908 & ~w15909;
assign w15911 = ~w15907 & w15910;
assign w15912 = (w15911 & ~w5888) | (w15911 & w26682) | (~w5888 & w26682);
assign w15913 = (w5888 & w30550) | (w5888 & w30551) | (w30550 & w30551);
assign w15914 = (~w5888 & w30552) | (~w5888 & w30553) | (w30552 & w30553);
assign w15915 = ~w15912 & ~w15913;
assign w15916 = ~w15914 & ~w15915;
assign w15917 = (~w30517 & w40688) | (~w30517 & w40689) | (w40688 & w40689);
assign w15918 = (w30517 & w40690) | (w30517 & w40691) | (w40690 & w40691);
assign w15919 = ~w15917 & ~w15918;
assign w15920 = b_40 & w3803;
assign w15921 = w4027 & w30556;
assign w15922 = b_39 & w3798;
assign w15923 = ~w15921 & ~w15922;
assign w15924 = ~w15920 & w15923;
assign w15925 = (w15924 & ~w5363) | (w15924 & w30557) | (~w5363 & w30557);
assign w15926 = (w5363 & w40692) | (w5363 & w40693) | (w40692 & w40693);
assign w15927 = (~w5363 & w40694) | (~w5363 & w40695) | (w40694 & w40695);
assign w15928 = ~w15925 & ~w15926;
assign w15929 = ~w15927 & ~w15928;
assign w15930 = (~w15773 & ~w15775) | (~w15773 & w30558) | (~w15775 & w30558);
assign w15931 = b_37 & w4499;
assign w15932 = w4723 & w30559;
assign w15933 = b_36 & w4494;
assign w15934 = ~w15932 & ~w15933;
assign w15935 = ~w15931 & w15934;
assign w15936 = (w15935 & ~w4636) | (w15935 & w30560) | (~w4636 & w30560);
assign w15937 = (w4636 & w40696) | (w4636 & w40697) | (w40696 & w40697);
assign w15938 = (~w4636 & w40698) | (~w4636 & w40699) | (w40698 & w40699);
assign w15939 = ~w15936 & ~w15937;
assign w15940 = ~w15938 & ~w15939;
assign w15941 = (~w15756 & w15759) | (~w15756 & w30561) | (w15759 & w30561);
assign w15942 = b_34 & w5196;
assign w15943 = w5459 & w30562;
assign w15944 = b_33 & w5191;
assign w15945 = ~w15943 & ~w15944;
assign w15946 = ~w15942 & w15945;
assign w15947 = (w15946 & ~w3967) | (w15946 & w30563) | (~w3967 & w30563);
assign w15948 = (w3967 & w40700) | (w3967 & w40701) | (w40700 & w40701);
assign w15949 = (~w3967 & w40702) | (~w3967 & w40703) | (w40702 & w40703);
assign w15950 = ~w15947 & ~w15948;
assign w15951 = ~w15949 & ~w15950;
assign w15952 = b_13 & w11620;
assign w15953 = w11969 & w30564;
assign w15954 = b_12 & w11615;
assign w15955 = ~w15953 & ~w15954;
assign w15956 = ~w15952 & w15955;
assign w15957 = (w15956 & ~w711) | (w15956 & w30565) | (~w711 & w30565);
assign w15958 = (w711 & w40704) | (w711 & w40705) | (w40704 & w40705);
assign w15959 = (~w711 & w40706) | (~w711 & w40707) | (w40706 & w40707);
assign w15960 = ~w15957 & ~w15958;
assign w15961 = ~w15959 & ~w15960;
assign w15962 = w12380 & w30566;
assign w15963 = b_10 & ~w12380;
assign w15964 = ~w15962 & ~w15963;
assign w15965 = ~a_8 & ~w15276;
assign w15966 = (~w15965 & w15653) | (~w15965 & w30567) | (w15653 & w30567);
assign w15967 = w15964 & ~w15966;
assign w15968 = w15966 & w15964;
assign w15969 = ~w15966 & ~w15967;
assign w15970 = ~w15968 & ~w15969;
assign w15971 = (~w15970 & w15960) | (~w15970 & w30568) | (w15960 & w30568);
assign w15972 = ~w15961 & ~w15971;
assign w15973 = ~w15970 & ~w15971;
assign w15974 = ~w15972 & ~w15973;
assign w15975 = (~w15657 & ~w15659) | (~w15657 & w30569) | (~w15659 & w30569);
assign w15976 = ~w15974 & ~w15975;
assign w15977 = ~w15974 & ~w15976;
assign w15978 = w15974 & ~w15975;
assign w15979 = ~w15977 & ~w15978;
assign w15980 = b_16 & w10562;
assign w15981 = w10902 & w30570;
assign w15982 = b_15 & w10557;
assign w15983 = ~w15981 & ~w15982;
assign w15984 = ~w15980 & w15983;
assign w15985 = (w15984 & ~w926) | (w15984 & w30571) | (~w926 & w30571);
assign w15986 = (w926 & w40708) | (w926 & w40709) | (w40708 & w40709);
assign w15987 = (~w926 & w40710) | (~w926 & w40711) | (w40710 & w40711);
assign w15988 = ~w15985 & ~w15986;
assign w15989 = ~w15987 & ~w15988;
assign w15990 = (~w15989 & w15977) | (~w15989 & w30572) | (w15977 & w30572);
assign w15991 = ~w15979 & ~w15990;
assign w15992 = ~w15989 & ~w15990;
assign w15993 = ~w15991 & ~w15992;
assign w15994 = (~w15673 & ~w15675) | (~w15673 & w40712) | (~w15675 & w40712);
assign w15995 = w15993 & w15994;
assign w15996 = ~w15993 & ~w15994;
assign w15997 = ~w15995 & ~w15996;
assign w15998 = b_19 & w9534;
assign w15999 = w9876 & w30573;
assign w16000 = b_18 & w9529;
assign w16001 = ~w15999 & ~w16000;
assign w16002 = ~w15998 & w16001;
assign w16003 = (w16002 & ~w1372) | (w16002 & w30574) | (~w1372 & w30574);
assign w16004 = (w1372 & w40713) | (w1372 & w40714) | (w40713 & w40714);
assign w16005 = (~w1372 & w40715) | (~w1372 & w40716) | (w40715 & w40716);
assign w16006 = ~w16003 & ~w16004;
assign w16007 = ~w16005 & ~w16006;
assign w16008 = w15997 & ~w16007;
assign w16009 = w15997 & ~w16008;
assign w16010 = ~w15997 & ~w16007;
assign w16011 = ~w15679 & ~w15684;
assign w16012 = ~w16009 & w30575;
assign w16013 = (~w16011 & w16009) | (~w16011 & w30576) | (w16009 & w30576);
assign w16014 = ~w16012 & ~w16013;
assign w16015 = b_22 & w8526;
assign w16016 = w8886 & w30577;
assign w16017 = b_21 & w8521;
assign w16018 = ~w16016 & ~w16017;
assign w16019 = ~w16015 & w16018;
assign w16020 = (w16019 & ~w1786) | (w16019 & w30578) | (~w1786 & w30578);
assign w16021 = (w1786 & w40717) | (w1786 & w40718) | (w40717 & w40718);
assign w16022 = (~w1786 & w40719) | (~w1786 & w40720) | (w40719 & w40720);
assign w16023 = ~w16020 & ~w16021;
assign w16024 = ~w16022 & ~w16023;
assign w16025 = w16014 & ~w16024;
assign w16026 = w16014 & ~w16025;
assign w16027 = ~w16014 & ~w16024;
assign w16028 = (~w15696 & w15699) | (~w15696 & w30579) | (w15699 & w30579);
assign w16029 = ~w16026 & w30580;
assign w16030 = (~w16028 & w16026) | (~w16028 & w30581) | (w16026 & w30581);
assign w16031 = ~w16029 & ~w16030;
assign w16032 = b_25 & w7613;
assign w16033 = w7941 & w30582;
assign w16034 = b_24 & w7608;
assign w16035 = ~w16033 & ~w16034;
assign w16036 = ~w16032 & w16035;
assign w16037 = (w16036 & ~w2108) | (w16036 & w30583) | (~w2108 & w30583);
assign w16038 = (w2108 & w40721) | (w2108 & w40722) | (w40721 & w40722);
assign w16039 = (~w2108 & w40723) | (~w2108 & w40724) | (w40723 & w40724);
assign w16040 = ~w16037 & ~w16038;
assign w16041 = ~w16039 & ~w16040;
assign w16042 = w16031 & ~w16041;
assign w16043 = w16031 & ~w16042;
assign w16044 = ~w16031 & ~w16041;
assign w16045 = ~w16043 & ~w16044;
assign w16046 = ~w15704 & ~w15708;
assign w16047 = w16045 & w16046;
assign w16048 = ~w16045 & ~w16046;
assign w16049 = ~w16047 & ~w16048;
assign w16050 = b_28 & w6761;
assign w16051 = w7075 & w30584;
assign w16052 = b_27 & w6756;
assign w16053 = ~w16051 & ~w16052;
assign w16054 = ~w16050 & w16053;
assign w16055 = (w16054 & ~w2771) | (w16054 & w30585) | (~w2771 & w30585);
assign w16056 = (w2771 & w40725) | (w2771 & w40726) | (w40725 & w40726);
assign w16057 = (~w2771 & w40727) | (~w2771 & w40728) | (w40727 & w40728);
assign w16058 = ~w16055 & ~w16056;
assign w16059 = ~w16057 & ~w16058;
assign w16060 = w16049 & ~w16059;
assign w16061 = w16049 & ~w16060;
assign w16062 = ~w16049 & ~w16059;
assign w16063 = ~w16061 & ~w16062;
assign w16064 = ~w15722 & ~w15727;
assign w16065 = w16063 & w16064;
assign w16066 = ~w16063 & ~w16064;
assign w16067 = ~w16065 & ~w16066;
assign w16068 = b_31 & w5962;
assign w16069 = w6246 & w30586;
assign w16070 = b_30 & w5957;
assign w16071 = ~w16069 & ~w16070;
assign w16072 = ~w16068 & w16071;
assign w16073 = (w16072 & ~w3345) | (w16072 & w30587) | (~w3345 & w30587);
assign w16074 = (w3345 & w40729) | (w3345 & w40730) | (w40729 & w40730);
assign w16075 = (~w3345 & w40731) | (~w3345 & w40732) | (w40731 & w40732);
assign w16076 = ~w16073 & ~w16074;
assign w16077 = ~w16075 & ~w16076;
assign w16078 = ~w16067 & w16077;
assign w16079 = w16067 & ~w16077;
assign w16080 = ~w16078 & ~w16079;
assign w16081 = ~w15743 & w16080;
assign w16082 = w15743 & ~w16080;
assign w16083 = ~w16081 & ~w16082;
assign w16084 = ~w15951 & w16083;
assign w16085 = w15951 & ~w16083;
assign w16086 = ~w16084 & ~w16085;
assign w16087 = ~w15941 & w16086;
assign w16088 = ~w15941 & ~w16087;
assign w16089 = w15941 & w16086;
assign w16090 = (~w15940 & w16088) | (~w15940 & w30588) | (w16088 & w30588);
assign w16091 = (w15940 & ~w15941) | (w15940 & w40733) | (~w15941 & w40733);
assign w16092 = ~w16088 & w16091;
assign w16093 = ~w16090 & ~w16092;
assign w16094 = ~w15930 & w16093;
assign w16095 = ~w15930 & ~w16094;
assign w16096 = w16093 & ~w16094;
assign w16097 = ~w16095 & ~w16096;
assign w16098 = ~w15929 & ~w16097;
assign w16099 = w16097 & ~w15929;
assign w16100 = ~w16097 & ~w16098;
assign w16101 = ~w16099 & ~w16100;
assign w16102 = w15919 & ~w16101;
assign w16103 = w15919 & ~w16102;
assign w16104 = ~w16101 & ~w16102;
assign w16105 = ~w16103 & ~w16104;
assign w16106 = b_46 & w2639;
assign w16107 = w2820 & w30589;
assign w16108 = b_45 & w2634;
assign w16109 = ~w16107 & ~w16108;
assign w16110 = ~w16106 & w16109;
assign w16111 = w16109 & w30590;
assign w16112 = (~w6974 & w25980) | (~w6974 & w25981) | (w25980 & w25981);
assign w16113 = (w6974 & w25982) | (w6974 & w25983) | (w25982 & w25983);
assign w16114 = ~w16112 & ~w16113;
assign w16115 = (~w15611 & w30593) | (~w15611 & w30594) | (w30593 & w30594);
assign w16116 = (w15611 & w40734) | (w15611 & w40735) | (w40734 & w40735);
assign w16117 = ~w16115 & ~w16116;
assign w16118 = (~w16105 & w16116) | (~w16105 & w30595) | (w16116 & w30595);
assign w16119 = ~w30595 & w40736;
assign w16120 = ~w16117 & ~w16118;
assign w16121 = ~w16119 & ~w16120;
assign w16122 = (~w16121 & w15904) | (~w16121 & w25664) | (w15904 & w25664);
assign w16123 = ~w15906 & ~w16122;
assign w16124 = ~w15904 & w40737;
assign w16125 = ~w16123 & ~w16124;
assign w16126 = w15891 & ~w16125;
assign w16127 = ~w15891 & w16125;
assign w16128 = w15877 & w27815;
assign w16129 = w15877 & ~w16128;
assign w16130 = (~w15877 & w27815) | (~w15877 & w40738) | (w27815 & w40738);
assign w16131 = ~w16129 & ~w16130;
assign w16132 = (~w15564 & w15567) | (~w15564 & w25665) | (w15567 & w25665);
assign w16133 = b_58 & w986;
assign w16134 = w1069 & w30597;
assign w16135 = b_57 & w981;
assign w16136 = ~w16134 & ~w16135;
assign w16137 = ~w16133 & w16136;
assign w16138 = w16136 & w30598;
assign w16139 = (~w10476 & w40739) | (~w10476 & w40740) | (w40739 & w40740);
assign w16140 = (w10476 & w30600) | (w10476 & w30601) | (w30600 & w30601);
assign w16141 = ~w16139 & ~w16140;
assign w16142 = (~w15567 & w30602) | (~w15567 & w30603) | (w30602 & w30603);
assign w16143 = ~w16132 & ~w16142;
assign w16144 = (w15567 & w30604) | (w15567 & w30605) | (w30604 & w30605);
assign w16145 = ~w16143 & ~w16144;
assign w16146 = (~w16131 & w16143) | (~w16131 & w30606) | (w16143 & w30606);
assign w16147 = ~w16131 & ~w16146;
assign w16148 = ~w16145 & ~w16146;
assign w16149 = ~w16147 & ~w16148;
assign w16150 = (~w16149 & w15863) | (~w16149 & w30607) | (w15863 & w30607);
assign w16151 = ~w15864 & ~w16150;
assign w16152 = ~w16149 & ~w16150;
assign w16153 = ~w16151 & ~w16152;
assign w16154 = (~w15535 & w15525) | (~w15535 & w30608) | (w15525 & w30608);
assign w16155 = (w15538 & w40741) | (w15538 & w40742) | (w40741 & w40742);
assign w16156 = w481 & w30609;
assign w16157 = b_63 & w413;
assign w16158 = ~w16156 & ~w16157;
assign w16159 = ~w12671 & w30610;
assign w16160 = (a_11 & w16159) | (a_11 & w30611) | (w16159 & w30611);
assign w16161 = ~w16159 & w30612;
assign w16162 = ~w16160 & ~w16161;
assign w16163 = (w15833 & w30613) | (w15833 & w30614) | (w30613 & w30614);
assign w16164 = ~w16155 & ~w16163;
assign w16165 = (~w15833 & w40743) | (~w15833 & w40744) | (w40743 & w40744);
assign w16166 = ~w16164 & ~w16165;
assign w16167 = (~w16153 & w16164) | (~w16153 & w40745) | (w16164 & w40745);
assign w16168 = (w16153 & w16163) | (w16153 & w30615) | (w16163 & w30615);
assign w16169 = ~w16164 & w16168;
assign w16170 = ~w16167 & ~w16169;
assign w16171 = ~w15849 & w16170;
assign w16172 = ~w15849 & ~w16171;
assign w16173 = w15849 & w16170;
assign w16174 = ~w16172 & ~w16173;
assign w16175 = (w14835 & w30616) | (w14835 & w30617) | (w30616 & w30617);
assign w16176 = (w13761 & w37680) | (w13761 & w37681) | (w37680 & w37681);
assign w16177 = ~w16175 & ~w16176;
assign w16178 = (~w16163 & w16166) | (~w16163 & w30621) | (w16166 & w30621);
assign w16179 = ~w15861 & ~w16150;
assign w16180 = w481 & w30622;
assign w16181 = (~w16180 & ~w12670) | (~w16180 & w30623) | (~w12670 & w30623);
assign w16182 = (w12670 & w40746) | (w12670 & w40747) | (w40746 & w40747);
assign w16183 = (~w12670 & w40748) | (~w12670 & w40749) | (w40748 & w40749);
assign w16184 = ~w16181 & ~w16182;
assign w16185 = ~w16183 & ~w16184;
assign w16186 = (~w16185 & w16150) | (~w16185 & w30624) | (w16150 & w30624);
assign w16187 = ~w16179 & ~w16186;
assign w16188 = ~w16150 & w30625;
assign w16189 = b_62 & w657;
assign w16190 = w754 & w30626;
assign w16191 = b_61 & w652;
assign w16192 = ~w16190 & ~w16191;
assign w16193 = ~w16189 & w16192;
assign w16194 = w16192 & w30627;
assign w16195 = (~w12273 & w40750) | (~w12273 & w40751) | (w40750 & w40751);
assign w16196 = (w12273 & w30629) | (w12273 & w30630) | (w30629 & w30630);
assign w16197 = ~w16195 & ~w16196;
assign w16198 = (~w16145 & w30631) | (~w16145 & w30632) | (w30631 & w30632);
assign w16199 = (w16145 & w30633) | (w16145 & w30634) | (w30633 & w30634);
assign w16200 = ~w16198 & ~w16199;
assign w16201 = b_59 & w986;
assign w16202 = w1069 & w30635;
assign w16203 = b_58 & w981;
assign w16204 = ~w16202 & ~w16203;
assign w16205 = ~w16201 & w16204;
assign w16206 = (w16205 & ~w11169) | (w16205 & w30636) | (~w11169 & w30636);
assign w16207 = (w11169 & w40752) | (w11169 & w40753) | (w40752 & w40753);
assign w16208 = (~w11169 & w40754) | (~w11169 & w40755) | (w40754 & w40755);
assign w16209 = ~w16206 & ~w16207;
assign w16210 = ~w16208 & ~w16209;
assign w16211 = (~w15876 & ~w15877) | (~w15876 & w30637) | (~w15877 & w30637);
assign w16212 = w16210 & w16211;
assign w16213 = ~w16210 & ~w16211;
assign w16214 = ~w16212 & ~w16213;
assign w16215 = b_56 & w1295;
assign w16216 = w1422 & w30638;
assign w16217 = b_55 & w1290;
assign w16218 = ~w16216 & ~w16217;
assign w16219 = ~w16215 & w16218;
assign w16220 = (w16219 & ~w9798) | (w16219 & w25984) | (~w9798 & w25984);
assign w16221 = (w9798 & w26365) | (w9798 & w26366) | (w26365 & w26366);
assign w16222 = (~w9798 & w30639) | (~w9798 & w30640) | (w30639 & w30640);
assign w16223 = ~w16220 & ~w16221;
assign w16224 = ~w16222 & ~w16223;
assign w16225 = (~w15890 & ~w15891) | (~w15890 & w25667) | (~w15891 & w25667);
assign w16226 = (~w25667 & w40756) | (~w25667 & w40757) | (w40756 & w40757);
assign w16227 = (w25667 & w40758) | (w25667 & w40759) | (w40758 & w40759);
assign w16228 = ~w16225 & ~w16226;
assign w16229 = ~w16227 & ~w16228;
assign w16230 = b_50 & w2158;
assign w16231 = w2294 & w30641;
assign w16232 = b_49 & w2153;
assign w16233 = ~w16231 & ~w16232;
assign w16234 = ~w16230 & w16233;
assign w16235 = w16233 & w30642;
assign w16236 = (~w8162 & w25985) | (~w8162 & w25986) | (w25985 & w25986);
assign w16237 = (w8162 & w25987) | (w8162 & w25988) | (w25987 & w25988);
assign w16238 = ~w16236 & ~w16237;
assign w16239 = (~w16117 & w30643) | (~w16117 & w30644) | (w30643 & w30644);
assign w16240 = (w16117 & w30645) | (w16117 & w30646) | (w30645 & w30646);
assign w16241 = ~w16239 & ~w16240;
assign w16242 = b_47 & w2639;
assign w16243 = w2820 & w30647;
assign w16244 = b_46 & w2634;
assign w16245 = ~w16243 & ~w16244;
assign w16246 = ~w16242 & w16245;
assign w16247 = (w16246 & ~w6998) | (w16246 & w25669) | (~w6998 & w25669);
assign w16248 = (w6998 & w25989) | (w6998 & w25990) | (w25989 & w25990);
assign w16249 = (~w6998 & w26367) | (~w6998 & w26368) | (w26367 & w26368);
assign w16250 = ~w16247 & ~w16248;
assign w16251 = ~w15918 & ~w16102;
assign w16252 = ~w16102 & w40760;
assign w16253 = (~w16251 & w16250) | (~w16251 & w26369) | (w16250 & w26369);
assign w16254 = ~w16252 & ~w16253;
assign w16255 = b_44 & w3195;
assign w16256 = w3388 & w30649;
assign w16257 = b_43 & w3190;
assign w16258 = ~w16256 & ~w16257;
assign w16259 = ~w16255 & w16258;
assign w16260 = w16258 & w30650;
assign w16261 = (~w6408 & w27587) | (~w6408 & w27588) | (w27587 & w27588);
assign w16262 = (w6408 & w27589) | (w6408 & w27590) | (w27589 & w27590);
assign w16263 = ~w16261 & ~w16262;
assign w16264 = (~w16097 & w30651) | (~w16097 & w30652) | (w30651 & w30652);
assign w16265 = (w16097 & w30653) | (w16097 & w30654) | (w30653 & w30654);
assign w16266 = ~w16264 & ~w16265;
assign w16267 = b_41 & w3803;
assign w16268 = w4027 & w30655;
assign w16269 = b_40 & w3798;
assign w16270 = ~w16268 & ~w16269;
assign w16271 = ~w16267 & w16270;
assign w16272 = (w16271 & ~w5609) | (w16271 & w30656) | (~w5609 & w30656);
assign w16273 = (w5609 & w40761) | (w5609 & w40762) | (w40761 & w40762);
assign w16274 = (~w5609 & w40763) | (~w5609 & w40764) | (w40763 & w40764);
assign w16275 = ~w16272 & ~w16273;
assign w16276 = ~w16274 & ~w16275;
assign w16277 = ~w16087 & ~w16090;
assign w16278 = b_35 & w5196;
assign w16279 = w5459 & w30657;
assign w16280 = b_34 & w5191;
assign w16281 = ~w16279 & ~w16280;
assign w16282 = ~w16278 & w16281;
assign w16283 = (w16282 & ~w4181) | (w16282 & w30658) | (~w4181 & w30658);
assign w16284 = (w4181 & w40765) | (w4181 & w40766) | (w40765 & w40766);
assign w16285 = (~w4181 & w40767) | (~w4181 & w40768) | (w40767 & w40768);
assign w16286 = ~w16283 & ~w16284;
assign w16287 = ~w16285 & ~w16286;
assign w16288 = (~w16030 & ~w16031) | (~w16030 & w30659) | (~w16031 & w30659);
assign w16289 = b_26 & w7613;
assign w16290 = w7941 & w30660;
assign w16291 = b_25 & w7608;
assign w16292 = ~w16290 & ~w16291;
assign w16293 = ~w16289 & w16292;
assign w16294 = (w16293 & ~w2416) | (w16293 & w30661) | (~w2416 & w30661);
assign w16295 = (w2416 & w40769) | (w2416 & w40770) | (w40769 & w40770);
assign w16296 = (~w2416 & w40771) | (~w2416 & w40772) | (w40771 & w40772);
assign w16297 = ~w16294 & ~w16295;
assign w16298 = ~w16296 & ~w16297;
assign w16299 = (~w16013 & ~w16014) | (~w16013 & w30662) | (~w16014 & w30662);
assign w16300 = b_23 & w8526;
assign w16301 = w8886 & w30663;
assign w16302 = b_22 & w8521;
assign w16303 = ~w16301 & ~w16302;
assign w16304 = ~w16300 & w16303;
assign w16305 = (w16304 & ~w1933) | (w16304 & w30664) | (~w1933 & w30664);
assign w16306 = (w1933 & w40773) | (w1933 & w40774) | (w40773 & w40774);
assign w16307 = (~w1933 & w40775) | (~w1933 & w40776) | (w40775 & w40776);
assign w16308 = ~w16305 & ~w16306;
assign w16309 = ~w16307 & ~w16308;
assign w16310 = (~w15996 & ~w15997) | (~w15996 & w30665) | (~w15997 & w30665);
assign w16311 = ~w15967 & ~w15971;
assign w16312 = w12380 & w30666;
assign w16313 = b_11 & ~w12380;
assign w16314 = ~w16312 & ~w16313;
assign w16315 = w15964 & ~w16314;
assign w16316 = w15964 & ~w16315;
assign w16317 = ~w16314 & ~w16315;
assign w16318 = ~w16316 & ~w16317;
assign w16319 = (~w16318 & w15971) | (~w16318 & w30667) | (w15971 & w30667);
assign w16320 = ~w16311 & ~w16319;
assign w16321 = ~w15971 & w30668;
assign w16322 = ~w16320 & ~w16321;
assign w16323 = b_14 & w11620;
assign w16324 = w11969 & w30669;
assign w16325 = b_13 & w11615;
assign w16326 = ~w16324 & ~w16325;
assign w16327 = ~w16323 & w16326;
assign w16328 = (w16327 & ~w735) | (w16327 & w30670) | (~w735 & w30670);
assign w16329 = (w735 & w40777) | (w735 & w40778) | (w40777 & w40778);
assign w16330 = (~w735 & w40779) | (~w735 & w40780) | (w40779 & w40780);
assign w16331 = ~w16328 & ~w16329;
assign w16332 = ~w16330 & ~w16331;
assign w16333 = (~w16332 & w16320) | (~w16332 & w30671) | (w16320 & w30671);
assign w16334 = ~w16322 & ~w16333;
assign w16335 = ~w16332 & ~w16333;
assign w16336 = ~w16334 & ~w16335;
assign w16337 = b_17 & w10562;
assign w16338 = w10902 & w30672;
assign w16339 = b_16 & w10557;
assign w16340 = ~w16338 & ~w16339;
assign w16341 = ~w16337 & w16340;
assign w16342 = (w16341 & ~w1038) | (w16341 & w30673) | (~w1038 & w30673);
assign w16343 = (w1038 & w40781) | (w1038 & w40782) | (w40781 & w40782);
assign w16344 = (~w1038 & w40783) | (~w1038 & w40784) | (w40783 & w40784);
assign w16345 = ~w16342 & ~w16343;
assign w16346 = ~w16344 & ~w16345;
assign w16347 = ~w16336 & ~w16346;
assign w16348 = ~w16336 & ~w16347;
assign w16349 = w16336 & ~w16346;
assign w16350 = ~w15976 & ~w15990;
assign w16351 = ~w16348 & w30674;
assign w16352 = (~w16350 & w16348) | (~w16350 & w30675) | (w16348 & w30675);
assign w16353 = ~w16351 & ~w16352;
assign w16354 = b_20 & w9534;
assign w16355 = w9876 & w30676;
assign w16356 = b_19 & w9529;
assign w16357 = ~w16355 & ~w16356;
assign w16358 = ~w16354 & w16357;
assign w16359 = (w16358 & ~w1503) | (w16358 & w30677) | (~w1503 & w30677);
assign w16360 = (w1503 & w40785) | (w1503 & w40786) | (w40785 & w40786);
assign w16361 = (~w1503 & w40787) | (~w1503 & w40788) | (w40787 & w40788);
assign w16362 = ~w16359 & ~w16360;
assign w16363 = ~w16361 & ~w16362;
assign w16364 = ~w16353 & w16363;
assign w16365 = w16353 & ~w16363;
assign w16366 = ~w16364 & ~w16365;
assign w16367 = ~w16310 & w16366;
assign w16368 = ~w16366 & ~w16310;
assign w16369 = w16366 & ~w16367;
assign w16370 = (~w16309 & w16369) | (~w16309 & w30678) | (w16369 & w30678);
assign w16371 = ~w16369 & w30679;
assign w16372 = ~w16370 & ~w16371;
assign w16373 = ~w16299 & w16372;
assign w16374 = w16299 & ~w16372;
assign w16375 = ~w16373 & ~w16374;
assign w16376 = ~w16298 & w16375;
assign w16377 = w16298 & ~w16375;
assign w16378 = ~w16376 & ~w16377;
assign w16379 = ~w16288 & w16378;
assign w16380 = w16288 & ~w16378;
assign w16381 = ~w16379 & ~w16380;
assign w16382 = b_29 & w6761;
assign w16383 = w7075 & w30680;
assign w16384 = b_28 & w6756;
assign w16385 = ~w16383 & ~w16384;
assign w16386 = ~w16382 & w16385;
assign w16387 = (w16386 & ~w2954) | (w16386 & w30681) | (~w2954 & w30681);
assign w16388 = (w2954 & w40789) | (w2954 & w40790) | (w40789 & w40790);
assign w16389 = (~w2954 & w40791) | (~w2954 & w40792) | (w40791 & w40792);
assign w16390 = ~w16387 & ~w16388;
assign w16391 = ~w16389 & ~w16390;
assign w16392 = w16381 & ~w16391;
assign w16393 = w16381 & ~w16392;
assign w16394 = ~w16381 & ~w16391;
assign w16395 = ~w16393 & ~w16394;
assign w16396 = (~w16048 & ~w16049) | (~w16048 & w30682) | (~w16049 & w30682);
assign w16397 = w16395 & w16396;
assign w16398 = ~w16395 & ~w16396;
assign w16399 = ~w16397 & ~w16398;
assign w16400 = b_32 & w5962;
assign w16401 = w6246 & w30683;
assign w16402 = b_31 & w5957;
assign w16403 = ~w16401 & ~w16402;
assign w16404 = ~w16400 & w16403;
assign w16405 = (w16404 & ~w3545) | (w16404 & w30684) | (~w3545 & w30684);
assign w16406 = (w3545 & w40793) | (w3545 & w40794) | (w40793 & w40794);
assign w16407 = (~w3545 & w40795) | (~w3545 & w40796) | (w40795 & w40796);
assign w16408 = ~w16405 & ~w16406;
assign w16409 = ~w16407 & ~w16408;
assign w16410 = ~w16399 & w16409;
assign w16411 = w16399 & ~w16409;
assign w16412 = ~w16410 & ~w16411;
assign w16413 = (~w16066 & ~w16067) | (~w16066 & w30685) | (~w16067 & w30685);
assign w16414 = w16412 & ~w16413;
assign w16415 = ~w16412 & w16413;
assign w16416 = ~w16414 & ~w16415;
assign w16417 = ~w16287 & w16416;
assign w16418 = w16416 & ~w16417;
assign w16419 = ~w16416 & ~w16287;
assign w16420 = ~w16418 & ~w16419;
assign w16421 = (~w16081 & ~w16083) | (~w16081 & w30686) | (~w16083 & w30686);
assign w16422 = w16420 & w16421;
assign w16423 = ~w16420 & ~w16421;
assign w16424 = ~w16422 & ~w16423;
assign w16425 = b_38 & w4499;
assign w16426 = w4723 & w30687;
assign w16427 = b_37 & w4494;
assign w16428 = ~w16426 & ~w16427;
assign w16429 = ~w16425 & w16428;
assign w16430 = (w16429 & ~w4658) | (w16429 & w30688) | (~w4658 & w30688);
assign w16431 = (w4658 & w40797) | (w4658 & w40798) | (w40797 & w40798);
assign w16432 = (~w4658 & w40799) | (~w4658 & w40800) | (w40799 & w40800);
assign w16433 = ~w16430 & ~w16431;
assign w16434 = ~w16432 & ~w16433;
assign w16435 = ~w16424 & w16434;
assign w16436 = w16424 & ~w16434;
assign w16437 = ~w16435 & ~w16436;
assign w16438 = ~w16277 & w16437;
assign w16439 = w16277 & ~w16437;
assign w16440 = ~w16438 & ~w16439;
assign w16441 = ~w16276 & w16440;
assign w16442 = ~w16440 & ~w16276;
assign w16443 = w16440 & ~w16441;
assign w16444 = ~w16442 & ~w16443;
assign w16445 = w16266 & ~w16444;
assign w16446 = w16266 & ~w16445;
assign w16447 = ~w16444 & ~w16445;
assign w16448 = ~w16446 & ~w16447;
assign w16449 = ~w16253 & w30689;
assign w16450 = (w16448 & w16253) | (w16448 & w30690) | (w16253 & w30690);
assign w16451 = w16241 & w26370;
assign w16452 = w16241 & ~w16451;
assign w16453 = w26370 & ~w16241;
assign w16454 = ~w16452 & ~w16453;
assign w16455 = (~w25664 & w25991) | (~w25664 & w25992) | (w25991 & w25992);
assign w16456 = b_53 & w1694;
assign w16457 = w1834 & w30691;
assign w16458 = b_52 & w1689;
assign w16459 = ~w16457 & ~w16458;
assign w16460 = ~w16456 & w16459;
assign w16461 = w16459 & w30692;
assign w16462 = (w9109 & w40801) | (w9109 & w40802) | (w40801 & w40802);
assign w16463 = (~w9109 & w40803) | (~w9109 & w40804) | (w40803 & w40804);
assign w16464 = ~w16462 & ~w16463;
assign w16465 = (~w25992 & w27591) | (~w25992 & w27592) | (w27591 & w27592);
assign w16466 = ~w16455 & ~w16465;
assign w16467 = w16455 & ~w16464;
assign w16468 = ~w16466 & ~w16467;
assign w16469 = (~w16454 & w16466) | (~w16454 & w30693) | (w16466 & w30693);
assign w16470 = ~w30693 & w40805;
assign w16471 = ~w16468 & ~w16469;
assign w16472 = ~w16470 & ~w16471;
assign w16473 = (~w16472 & w16228) | (~w16472 & w30694) | (w16228 & w30694);
assign w16474 = ~w16229 & ~w16473;
assign w16475 = ~w30694 & w40806;
assign w16476 = ~w16474 & ~w16475;
assign w16477 = w16214 & ~w16476;
assign w16478 = ~w16214 & w16476;
assign w16479 = w16200 & w30695;
assign w16480 = w16200 & ~w16479;
assign w16481 = w30695 & ~w16200;
assign w16482 = ~w16480 & ~w16481;
assign w16483 = (w16482 & w16187) | (w16482 & w30696) | (w16187 & w30696);
assign w16484 = ~w16187 & w30697;
assign w16485 = ~w16483 & ~w16484;
assign w16486 = (~w16166 & w30698) | (~w16166 & w30699) | (w30698 & w30699);
assign w16487 = ~w16178 & ~w16486;
assign w16488 = ~w16485 & ~w16486;
assign w16489 = ~w16487 & ~w16488;
assign w16490 = (w14835 & w27757) | (w14835 & w27758) | (w27757 & w27758);
assign w16491 = (w13761 & w37682) | (w13761 & w37683) | (w37682 & w37683);
assign w16492 = ~w16490 & ~w16491;
assign w16493 = (~w16482 & w16187) | (~w16482 & w30703) | (w16187 & w30703);
assign w16494 = ~w16186 & ~w16493;
assign w16495 = (~w16198 & ~w16200) | (~w16198 & w30704) | (~w16200 & w30704);
assign w16496 = b_63 & w657;
assign w16497 = w754 & w30705;
assign w16498 = b_62 & w652;
assign w16499 = ~w16497 & ~w16498;
assign w16500 = ~w16496 & w16499;
assign w16501 = (w16500 & ~w12646) | (w16500 & w30706) | (~w12646 & w30706);
assign w16502 = (w12646 & w40807) | (w12646 & w40808) | (w40807 & w40808);
assign w16503 = (~w12646 & w40809) | (~w12646 & w40810) | (w40809 & w40810);
assign w16504 = ~w16501 & ~w16502;
assign w16505 = ~w16503 & ~w16504;
assign w16506 = ~w16495 & ~w16505;
assign w16507 = ~w16495 & ~w16506;
assign w16508 = w16495 & ~w16505;
assign w16509 = b_60 & w986;
assign w16510 = w1069 & w30707;
assign w16511 = b_59 & w981;
assign w16512 = ~w16510 & ~w16511;
assign w16513 = ~w16509 & w16512;
assign w16514 = (w16513 & ~w11196) | (w16513 & w30708) | (~w11196 & w30708);
assign w16515 = (w11196 & w40811) | (w11196 & w40812) | (w40811 & w40812);
assign w16516 = (~w11196 & w40813) | (~w11196 & w40814) | (w40813 & w40814);
assign w16517 = ~w16514 & ~w16515;
assign w16518 = ~w16516 & ~w16517;
assign w16519 = (w16518 & w16477) | (w16518 & w30709) | (w16477 & w30709);
assign w16520 = ~w16477 & w30710;
assign w16521 = ~w16519 & ~w16520;
assign w16522 = b_57 & w1295;
assign w16523 = w1422 & w30711;
assign w16524 = b_56 & w1290;
assign w16525 = ~w16523 & ~w16524;
assign w16526 = ~w16522 & w16525;
assign w16527 = (w16526 & ~w10452) | (w16526 & w30712) | (~w10452 & w30712);
assign w16528 = (w10452 & w40815) | (w10452 & w40816) | (w40815 & w40816);
assign w16529 = (~w10452 & w40817) | (~w10452 & w40818) | (w40817 & w40818);
assign w16530 = ~w16527 & ~w16528;
assign w16531 = ~w16529 & ~w16530;
assign w16532 = (~w30694 & w40819) | (~w30694 & w40820) | (w40819 & w40820);
assign w16533 = (w30694 & w40821) | (w30694 & w40822) | (w40821 & w40822);
assign w16534 = ~w16532 & ~w16533;
assign w16535 = (~w16465 & w16468) | (~w16465 & w26371) | (w16468 & w26371);
assign w16536 = b_54 & w1694;
assign w16537 = w1834 & w30715;
assign w16538 = b_53 & w1689;
assign w16539 = ~w16537 & ~w16538;
assign w16540 = ~w16536 & w16539;
assign w16541 = (w16540 & ~w9134) | (w16540 & w26372) | (~w9134 & w26372);
assign w16542 = (w9134 & w30716) | (w9134 & w30717) | (w30716 & w30717);
assign w16543 = (~w9134 & w30718) | (~w9134 & w30719) | (w30718 & w30719);
assign w16544 = ~w16541 & ~w16542;
assign w16545 = ~w16543 & ~w16544;
assign w16546 = (~w16468 & w30720) | (~w16468 & w30721) | (w30720 & w30721);
assign w16547 = ~w16535 & ~w16546;
assign w16548 = (w16468 & w30722) | (w16468 & w30723) | (w30722 & w30723);
assign w16549 = ~w16547 & ~w16548;
assign w16550 = b_51 & w2158;
assign w16551 = w2294 & w30724;
assign w16552 = b_50 & w2153;
assign w16553 = ~w16551 & ~w16552;
assign w16554 = ~w16550 & w16553;
assign w16555 = (w16554 & ~w8186) | (w16554 & w30725) | (~w8186 & w30725);
assign w16556 = (w8186 & w40823) | (w8186 & w40824) | (w40823 & w40824);
assign w16557 = (~w8186 & w40825) | (~w8186 & w40826) | (w40825 & w40826);
assign w16558 = ~w16555 & ~w16556;
assign w16559 = ~w16557 & ~w16558;
assign w16560 = (~w16239 & ~w16241) | (~w16239 & w30726) | (~w16241 & w30726);
assign w16561 = w16559 & w16560;
assign w16562 = ~w16559 & ~w16560;
assign w16563 = ~w16561 & ~w16562;
assign w16564 = (~w16253 & ~w16254) | (~w16253 & w26684) | (~w16254 & w26684);
assign w16565 = b_48 & w2639;
assign w16566 = w2820 & w30727;
assign w16567 = b_47 & w2634;
assign w16568 = ~w16566 & ~w16567;
assign w16569 = ~w16565 & w16568;
assign w16570 = (w16569 & ~w7284) | (w16569 & w26685) | (~w7284 & w26685);
assign w16571 = (w7284 & w27593) | (w7284 & w27594) | (w27593 & w27594);
assign w16572 = (~w7284 & w30728) | (~w7284 & w30729) | (w30728 & w30729);
assign w16573 = ~w16570 & ~w16571;
assign w16574 = ~w16572 & ~w16573;
assign w16575 = ~w16564 & w16574;
assign w16576 = w16564 & ~w16574;
assign w16577 = ~w16575 & ~w16576;
assign w16578 = (~w16438 & ~w16440) | (~w16438 & w30730) | (~w16440 & w30730);
assign w16579 = (~w16423 & ~w16424) | (~w16423 & w30731) | (~w16424 & w30731);
assign w16580 = (~w16414 & ~w16416) | (~w16414 & w30732) | (~w16416 & w30732);
assign w16581 = (~w16398 & ~w16399) | (~w16398 & w30733) | (~w16399 & w30733);
assign w16582 = (~w16379 & ~w16381) | (~w16379 & w30734) | (~w16381 & w30734);
assign w16583 = ~w16367 & ~w16370;
assign w16584 = b_24 & w8526;
assign w16585 = w8886 & w30735;
assign w16586 = b_23 & w8521;
assign w16587 = ~w16585 & ~w16586;
assign w16588 = ~w16584 & w16587;
assign w16589 = (w16588 & ~w2083) | (w16588 & w30736) | (~w2083 & w30736);
assign w16590 = (w2083 & w40827) | (w2083 & w40828) | (w40827 & w40828);
assign w16591 = (~w2083 & w40829) | (~w2083 & w40830) | (w40829 & w40830);
assign w16592 = ~w16589 & ~w16590;
assign w16593 = ~w16591 & ~w16592;
assign w16594 = (~w15971 & w30737) | (~w15971 & w30738) | (w30737 & w30738);
assign w16595 = b_15 & w11620;
assign w16596 = w11969 & w30739;
assign w16597 = b_14 & w11615;
assign w16598 = ~w16596 & ~w16597;
assign w16599 = ~w16595 & w16598;
assign w16600 = (w16599 & ~w827) | (w16599 & w30740) | (~w827 & w30740);
assign w16601 = (w827 & w40831) | (w827 & w40832) | (w40831 & w40832);
assign w16602 = (~w827 & w40833) | (~w827 & w40834) | (w40833 & w40834);
assign w16603 = ~w16600 & ~w16601;
assign w16604 = ~w16602 & ~w16603;
assign w16605 = w12380 & w30741;
assign w16606 = b_12 & ~w12380;
assign w16607 = ~w16605 & ~w16606;
assign w16608 = a_11 & ~w15964;
assign w16609 = ~a_11 & w15964;
assign w16610 = ~w16608 & ~w16609;
assign w16611 = ~w16607 & ~w16610;
assign w16612 = w16607 & w16610;
assign w16613 = ~w16611 & ~w16612;
assign w16614 = (w16613 & w16603) | (w16613 & w30742) | (w16603 & w30742);
assign w16615 = ~w16604 & ~w16614;
assign w16616 = w16613 & ~w16614;
assign w16617 = ~w16615 & ~w16616;
assign w16618 = ~w16594 & ~w16617;
assign w16619 = w16617 & ~w16594;
assign w16620 = ~w16617 & ~w16618;
assign w16621 = ~w16619 & ~w16620;
assign w16622 = b_18 & w10562;
assign w16623 = w10902 & w30743;
assign w16624 = b_17 & w10557;
assign w16625 = ~w16623 & ~w16624;
assign w16626 = ~w16622 & w16625;
assign w16627 = (w16626 & ~w1238) | (w16626 & w30744) | (~w1238 & w30744);
assign w16628 = (w1238 & w40835) | (w1238 & w40836) | (w40835 & w40836);
assign w16629 = (~w1238 & w40837) | (~w1238 & w40838) | (w40837 & w40838);
assign w16630 = ~w16627 & ~w16628;
assign w16631 = ~w16629 & ~w16630;
assign w16632 = (~w16631 & w16620) | (~w16631 & w30745) | (w16620 & w30745);
assign w16633 = ~w16621 & ~w16632;
assign w16634 = ~w16631 & ~w16632;
assign w16635 = ~w16633 & ~w16634;
assign w16636 = (~w16333 & w16336) | (~w16333 & w30746) | (w16336 & w30746);
assign w16637 = w16635 & w16636;
assign w16638 = ~w16635 & ~w16636;
assign w16639 = ~w16637 & ~w16638;
assign w16640 = b_21 & w9534;
assign w16641 = w9876 & w30747;
assign w16642 = b_20 & w9529;
assign w16643 = ~w16641 & ~w16642;
assign w16644 = ~w16640 & w16643;
assign w16645 = (w16644 & ~w1634) | (w16644 & w30748) | (~w1634 & w30748);
assign w16646 = (w1634 & w40839) | (w1634 & w40840) | (w40839 & w40840);
assign w16647 = (~w1634 & w40841) | (~w1634 & w40842) | (w40841 & w40842);
assign w16648 = ~w16645 & ~w16646;
assign w16649 = ~w16647 & ~w16648;
assign w16650 = w16639 & ~w16649;
assign w16651 = w16639 & ~w16650;
assign w16652 = ~w16639 & ~w16649;
assign w16653 = (~w16352 & ~w16353) | (~w16352 & w30749) | (~w16353 & w30749);
assign w16654 = (~w16653 & w16651) | (~w16653 & w30750) | (w16651 & w30750);
assign w16655 = ~w16651 & w30751;
assign w16656 = ~w16654 & ~w16655;
assign w16657 = ~w16593 & w16656;
assign w16658 = ~w16656 & ~w16593;
assign w16659 = w16656 & ~w16657;
assign w16660 = ~w16658 & ~w16659;
assign w16661 = ~w16583 & ~w16660;
assign w16662 = w16660 & ~w16583;
assign w16663 = ~w16660 & ~w16661;
assign w16664 = ~w16662 & ~w16663;
assign w16665 = b_27 & w7613;
assign w16666 = w7941 & w30752;
assign w16667 = b_26 & w7608;
assign w16668 = ~w16666 & ~w16667;
assign w16669 = ~w16665 & w16668;
assign w16670 = (w16669 & ~w2582) | (w16669 & w30753) | (~w2582 & w30753);
assign w16671 = (w2582 & w40843) | (w2582 & w40844) | (w40843 & w40844);
assign w16672 = (~w2582 & w40845) | (~w2582 & w40846) | (w40845 & w40846);
assign w16673 = ~w16670 & ~w16671;
assign w16674 = ~w16672 & ~w16673;
assign w16675 = (~w16674 & w16663) | (~w16674 & w30754) | (w16663 & w30754);
assign w16676 = ~w16664 & ~w16675;
assign w16677 = ~w16674 & ~w16675;
assign w16678 = ~w16676 & ~w16677;
assign w16679 = (~w16373 & ~w16375) | (~w16373 & w30755) | (~w16375 & w30755);
assign w16680 = w16678 & w16679;
assign w16681 = ~w16678 & ~w16679;
assign w16682 = ~w16680 & ~w16681;
assign w16683 = b_30 & w6761;
assign w16684 = w7075 & w30756;
assign w16685 = b_29 & w6756;
assign w16686 = ~w16684 & ~w16685;
assign w16687 = ~w16683 & w16686;
assign w16688 = (w16687 & ~w3138) | (w16687 & w30757) | (~w3138 & w30757);
assign w16689 = (w3138 & w40847) | (w3138 & w40848) | (w40847 & w40848);
assign w16690 = (~w3138 & w40849) | (~w3138 & w40850) | (w40849 & w40850);
assign w16691 = ~w16688 & ~w16689;
assign w16692 = ~w16690 & ~w16691;
assign w16693 = w16682 & ~w16692;
assign w16694 = ~w16682 & w16692;
assign w16695 = (~w16582 & w16682) | (~w16582 & w30758) | (w16682 & w30758);
assign w16696 = ~w16693 & w16695;
assign w16697 = ~w16582 & ~w16696;
assign w16698 = ~w16693 & ~w16696;
assign w16699 = ~w16696 & w30759;
assign w16700 = ~w16697 & ~w16699;
assign w16701 = b_33 & w5962;
assign w16702 = w6246 & w30760;
assign w16703 = b_32 & w5957;
assign w16704 = ~w16702 & ~w16703;
assign w16705 = ~w16701 & w16704;
assign w16706 = (w16705 & ~w3744) | (w16705 & w30761) | (~w3744 & w30761);
assign w16707 = (w3744 & w40851) | (w3744 & w40852) | (w40851 & w40852);
assign w16708 = (~w3744 & w40853) | (~w3744 & w40854) | (w40853 & w40854);
assign w16709 = ~w16706 & ~w16707;
assign w16710 = ~w16708 & ~w16709;
assign w16711 = ~w16700 & ~w16710;
assign w16712 = ~w16700 & ~w16711;
assign w16713 = w16700 & ~w16710;
assign w16714 = ~w16712 & w30762;
assign w16715 = (w16581 & w16712) | (w16581 & w30763) | (w16712 & w30763);
assign w16716 = ~w16714 & ~w16715;
assign w16717 = b_36 & w5196;
assign w16718 = w5459 & w30764;
assign w16719 = b_35 & w5191;
assign w16720 = ~w16718 & ~w16719;
assign w16721 = ~w16717 & w16720;
assign w16722 = (w16721 & ~w4395) | (w16721 & w30765) | (~w4395 & w30765);
assign w16723 = (w4395 & w40855) | (w4395 & w40856) | (w40855 & w40856);
assign w16724 = (~w4395 & w40857) | (~w4395 & w40858) | (w40857 & w40858);
assign w16725 = ~w16722 & ~w16723;
assign w16726 = ~w16724 & ~w16725;
assign w16727 = ~w16716 & ~w16726;
assign w16728 = w16716 & w16726;
assign w16729 = ~w16727 & ~w16728;
assign w16730 = w16580 & ~w16729;
assign w16731 = ~w16580 & w16729;
assign w16732 = ~w16730 & ~w16731;
assign w16733 = b_39 & w4499;
assign w16734 = w4723 & w30766;
assign w16735 = b_38 & w4494;
assign w16736 = ~w16734 & ~w16735;
assign w16737 = ~w16733 & w16736;
assign w16738 = (w16737 & ~w4888) | (w16737 & w30767) | (~w4888 & w30767);
assign w16739 = (w4888 & w40859) | (w4888 & w40860) | (w40859 & w40860);
assign w16740 = (~w4888 & w40861) | (~w4888 & w40862) | (w40861 & w40862);
assign w16741 = ~w16738 & ~w16739;
assign w16742 = ~w16740 & ~w16741;
assign w16743 = w16732 & ~w16742;
assign w16744 = w16732 & ~w16743;
assign w16745 = ~w16732 & ~w16742;
assign w16746 = ~w16744 & w30768;
assign w16747 = (w16579 & w16744) | (w16579 & w30769) | (w16744 & w30769);
assign w16748 = ~w16746 & ~w16747;
assign w16749 = b_42 & w3803;
assign w16750 = w4027 & w30770;
assign w16751 = b_41 & w3798;
assign w16752 = ~w16750 & ~w16751;
assign w16753 = ~w16749 & w16752;
assign w16754 = (w16753 & ~w5864) | (w16753 & w30771) | (~w5864 & w30771);
assign w16755 = (w5864 & w40863) | (w5864 & w40864) | (w40863 & w40864);
assign w16756 = (~w5864 & w40865) | (~w5864 & w40866) | (w40865 & w40866);
assign w16757 = ~w16754 & ~w16755;
assign w16758 = ~w16756 & ~w16757;
assign w16759 = ~w16748 & ~w16758;
assign w16760 = w16748 & w16758;
assign w16761 = ~w16759 & ~w16760;
assign w16762 = w16578 & ~w16761;
assign w16763 = ~w16578 & w16761;
assign w16764 = ~w16762 & ~w16763;
assign w16765 = ~w16264 & ~w16445;
assign w16766 = b_45 & w3195;
assign w16767 = w3388 & w30772;
assign w16768 = b_44 & w3190;
assign w16769 = ~w16767 & ~w16768;
assign w16770 = ~w16766 & w16769;
assign w16771 = (w16770 & ~w6682) | (w16770 & w27595) | (~w6682 & w27595);
assign w16772 = (w6682 & w30773) | (w6682 & w30774) | (w30773 & w30774);
assign w16773 = (~w6682 & w30775) | (~w6682 & w30776) | (w30775 & w30776);
assign w16774 = ~w16771 & ~w16772;
assign w16775 = ~w16773 & ~w16774;
assign w16776 = (~w16775 & w16445) | (~w16775 & w30777) | (w16445 & w30777);
assign w16777 = ~w16765 & ~w16776;
assign w16778 = (w16764 & w16777) | (w16764 & w30779) | (w16777 & w30779);
assign w16779 = ~w16777 & w30780;
assign w16780 = ~w16577 & w27596;
assign w16781 = ~w16577 & ~w16780;
assign w16782 = w27596 & w16577;
assign w16783 = ~w16781 & ~w16782;
assign w16784 = w16563 & ~w16783;
assign w16785 = ~w16563 & w16783;
assign w16786 = (~w16785 & w16547) | (~w16785 & w26686) | (w16547 & w26686);
assign w16787 = ~w16784 & w16786;
assign w16788 = ~w16549 & ~w16787;
assign w16789 = (~w16786 & w30782) | (~w16786 & w30783) | (w30782 & w30783);
assign w16790 = ~w16788 & ~w16789;
assign w16791 = w16534 & ~w16790;
assign w16792 = ~w16534 & w16790;
assign w16793 = ~w16521 & w30784;
assign w16794 = ~w16521 & ~w16793;
assign w16795 = (w16521 & w30784) | (w16521 & w40867) | (w30784 & w40867);
assign w16796 = ~w16794 & ~w16795;
assign w16797 = (w16796 & w16507) | (w16796 & w30786) | (w16507 & w30786);
assign w16798 = ~w16507 & w30787;
assign w16799 = ~w16797 & ~w16798;
assign w16800 = (~w16799 & w16493) | (~w16799 & w30788) | (w16493 & w30788);
assign w16801 = ~w16494 & ~w16800;
assign w16802 = ~w16493 & w30789;
assign w16803 = ~w16801 & ~w16802;
assign w16804 = (w14835 & w30790) | (w14835 & w30791) | (w30790 & w30791);
assign w16805 = (w13761 & w37684) | (w13761 & w37685) | (w37684 & w37685);
assign w16806 = ~w16804 & ~w16805;
assign w16807 = (~w16796 & w16507) | (~w16796 & w30795) | (w16507 & w30795);
assign w16808 = ~w16506 & ~w16807;
assign w16809 = b_61 & w986;
assign w16810 = w1069 & w30796;
assign w16811 = b_60 & w981;
assign w16812 = ~w16810 & ~w16811;
assign w16813 = ~w16809 & w16812;
assign w16814 = (w16813 & ~w11901) | (w16813 & w30797) | (~w11901 & w30797);
assign w16815 = (w11901 & w40868) | (w11901 & w40869) | (w40868 & w40869);
assign w16816 = (~w11901 & w40870) | (~w11901 & w40871) | (w40870 & w40871);
assign w16817 = ~w16814 & ~w16815;
assign w16818 = ~w16816 & ~w16817;
assign w16819 = (~w16533 & ~w16534) | (~w16533 & w30798) | (~w16534 & w30798);
assign w16820 = (~w30798 & w40872) | (~w30798 & w40873) | (w40872 & w40873);
assign w16821 = (w30798 & w40874) | (w30798 & w40875) | (w40874 & w40875);
assign w16822 = ~w16819 & ~w16820;
assign w16823 = ~w16821 & ~w16822;
assign w16824 = b_55 & w1694;
assign w16825 = w1834 & w30799;
assign w16826 = b_54 & w1689;
assign w16827 = ~w16825 & ~w16826;
assign w16828 = ~w16824 & w16827;
assign w16829 = (w16828 & ~w9776) | (w16828 & w30800) | (~w9776 & w30800);
assign w16830 = (w9776 & w40876) | (w9776 & w40877) | (w40876 & w40877);
assign w16831 = (~w9776 & w40878) | (~w9776 & w40879) | (w40878 & w40879);
assign w16832 = ~w16829 & ~w16830;
assign w16833 = ~w16831 & ~w16832;
assign w16834 = (~w16562 & ~w16563) | (~w16562 & w30801) | (~w16563 & w30801);
assign w16835 = ~w16833 & ~w16834;
assign w16836 = w16834 & ~w16833;
assign w16837 = ~w16834 & ~w16835;
assign w16838 = ~w16836 & ~w16837;
assign w16839 = b_49 & w2639;
assign w16840 = w2820 & w30802;
assign w16841 = b_48 & w2634;
assign w16842 = ~w16840 & ~w16841;
assign w16843 = ~w16839 & w16842;
assign w16844 = (w16843 & ~w7859) | (w16843 & w26373) | (~w7859 & w26373);
assign w16845 = (w7859 & w27597) | (w7859 & w27598) | (w27597 & w27598);
assign w16846 = (~w7859 & w30803) | (~w7859 & w30804) | (w30803 & w30804);
assign w16847 = ~w16844 & ~w16845;
assign w16848 = ~w16846 & ~w16847;
assign w16849 = (~w16777 & w40880) | (~w16777 & w40881) | (w40880 & w40881);
assign w16850 = (w16777 & w40882) | (w16777 & w40883) | (w40882 & w40883);
assign w16851 = (~w16777 & w40884) | (~w16777 & w40885) | (w40884 & w40885);
assign w16852 = ~w16849 & ~w16850;
assign w16853 = ~w16851 & ~w16852;
assign w16854 = b_43 & w3803;
assign w16855 = w4027 & w30807;
assign w16856 = b_42 & w3798;
assign w16857 = ~w16855 & ~w16856;
assign w16858 = ~w16854 & w16857;
assign w16859 = (w16858 & ~w5888) | (w16858 & w30808) | (~w5888 & w30808);
assign w16860 = (w5888 & w40886) | (w5888 & w40887) | (w40886 & w40887);
assign w16861 = (~w5888 & w40888) | (~w5888 & w40889) | (w40888 & w40889);
assign w16862 = ~w16859 & ~w16860;
assign w16863 = ~w16861 & ~w16862;
assign w16864 = (~w16579 & w16744) | (~w16579 & w30809) | (w16744 & w30809);
assign w16865 = ~w16743 & ~w16864;
assign w16866 = b_40 & w4499;
assign w16867 = w4723 & w30810;
assign w16868 = b_39 & w4494;
assign w16869 = ~w16867 & ~w16868;
assign w16870 = ~w16866 & w16869;
assign w16871 = (w16870 & ~w5363) | (w16870 & w30811) | (~w5363 & w30811);
assign w16872 = (w5363 & w40890) | (w5363 & w40891) | (w40890 & w40891);
assign w16873 = (~w5363 & w40892) | (~w5363 & w40893) | (w40892 & w40893);
assign w16874 = ~w16871 & ~w16872;
assign w16875 = ~w16873 & ~w16874;
assign w16876 = (~w16727 & ~w16729) | (~w16727 & w30812) | (~w16729 & w30812);
assign w16877 = b_37 & w5196;
assign w16878 = w5459 & w30813;
assign w16879 = b_36 & w5191;
assign w16880 = ~w16878 & ~w16879;
assign w16881 = ~w16877 & w16880;
assign w16882 = (w16881 & ~w4636) | (w16881 & w30814) | (~w4636 & w30814);
assign w16883 = (w4636 & w40894) | (w4636 & w40895) | (w40894 & w40895);
assign w16884 = (~w4636 & w40896) | (~w4636 & w40897) | (w40896 & w40897);
assign w16885 = ~w16882 & ~w16883;
assign w16886 = ~w16884 & ~w16885;
assign w16887 = (~w16581 & w16712) | (~w16581 & w30815) | (w16712 & w30815);
assign w16888 = ~w16711 & ~w16887;
assign w16889 = b_34 & w5962;
assign w16890 = w6246 & w30816;
assign w16891 = b_33 & w5957;
assign w16892 = ~w16890 & ~w16891;
assign w16893 = ~w16889 & w16892;
assign w16894 = (w16893 & ~w3967) | (w16893 & w30817) | (~w3967 & w30817);
assign w16895 = (w3967 & w40898) | (w3967 & w40899) | (w40898 & w40899);
assign w16896 = (~w3967 & w40900) | (~w3967 & w40901) | (w40900 & w40901);
assign w16897 = ~w16894 & ~w16895;
assign w16898 = ~w16896 & ~w16897;
assign w16899 = b_31 & w6761;
assign w16900 = w7075 & w30818;
assign w16901 = b_30 & w6756;
assign w16902 = ~w16900 & ~w16901;
assign w16903 = ~w16899 & w16902;
assign w16904 = (w16903 & ~w3345) | (w16903 & w30819) | (~w3345 & w30819);
assign w16905 = (w3345 & w40902) | (w3345 & w40903) | (w40902 & w40903);
assign w16906 = (~w3345 & w40904) | (~w3345 & w40905) | (w40904 & w40905);
assign w16907 = ~w16904 & ~w16905;
assign w16908 = ~w16906 & ~w16907;
assign w16909 = (~w16675 & w16678) | (~w16675 & w30820) | (w16678 & w30820);
assign w16910 = w12380 & w30821;
assign w16911 = b_13 & ~w12380;
assign w16912 = ~w16910 & ~w16911;
assign w16913 = ~a_11 & ~w15964;
assign w16914 = (~w16913 & w16610) | (~w16913 & w30822) | (w16610 & w30822);
assign w16915 = w16912 & ~w16914;
assign w16916 = w16914 & w16912;
assign w16917 = ~w16914 & ~w16915;
assign w16918 = ~w16916 & ~w16917;
assign w16919 = b_16 & w11620;
assign w16920 = w11969 & w30823;
assign w16921 = b_15 & w11615;
assign w16922 = ~w16920 & ~w16921;
assign w16923 = ~w16919 & w16922;
assign w16924 = (w16923 & ~w926) | (w16923 & w30824) | (~w926 & w30824);
assign w16925 = (w926 & w40906) | (w926 & w40907) | (w40906 & w40907);
assign w16926 = ~w16924 & ~w16925;
assign w16927 = ~w16926 & w30825;
assign w16928 = (w16918 & w16926) | (w16918 & w30826) | (w16926 & w30826);
assign w16929 = ~w16927 & ~w16928;
assign w16930 = (~w16614 & w16617) | (~w16614 & w30827) | (w16617 & w30827);
assign w16931 = w16929 & w16930;
assign w16932 = ~w16929 & ~w16930;
assign w16933 = ~w16931 & ~w16932;
assign w16934 = b_19 & w10562;
assign w16935 = w10902 & w30828;
assign w16936 = b_18 & w10557;
assign w16937 = ~w16935 & ~w16936;
assign w16938 = ~w16934 & w16937;
assign w16939 = (w16938 & ~w1372) | (w16938 & w30829) | (~w1372 & w30829);
assign w16940 = (w1372 & w40908) | (w1372 & w40909) | (w40908 & w40909);
assign w16941 = (~w1372 & w40910) | (~w1372 & w40911) | (w40910 & w40911);
assign w16942 = ~w16939 & ~w16940;
assign w16943 = ~w16941 & ~w16942;
assign w16944 = w16933 & ~w16943;
assign w16945 = w16933 & ~w16944;
assign w16946 = ~w16933 & ~w16943;
assign w16947 = ~w16945 & ~w16946;
assign w16948 = (~w16632 & w16635) | (~w16632 & w30830) | (w16635 & w30830);
assign w16949 = w16947 & w16948;
assign w16950 = ~w16947 & ~w16948;
assign w16951 = ~w16949 & ~w16950;
assign w16952 = b_22 & w9534;
assign w16953 = w9876 & w30831;
assign w16954 = b_21 & w9529;
assign w16955 = ~w16953 & ~w16954;
assign w16956 = ~w16952 & w16955;
assign w16957 = (w16956 & ~w1786) | (w16956 & w30832) | (~w1786 & w30832);
assign w16958 = (w1786 & w40912) | (w1786 & w40913) | (w40912 & w40913);
assign w16959 = (~w1786 & w40914) | (~w1786 & w40915) | (w40914 & w40915);
assign w16960 = ~w16957 & ~w16958;
assign w16961 = ~w16959 & ~w16960;
assign w16962 = w16951 & ~w16961;
assign w16963 = w16951 & ~w16962;
assign w16964 = ~w16951 & ~w16961;
assign w16965 = ~w16963 & ~w16964;
assign w16966 = ~w16650 & ~w16654;
assign w16967 = w16965 & w16966;
assign w16968 = ~w16965 & ~w16966;
assign w16969 = ~w16967 & ~w16968;
assign w16970 = b_25 & w8526;
assign w16971 = w8886 & w30833;
assign w16972 = b_24 & w8521;
assign w16973 = ~w16971 & ~w16972;
assign w16974 = ~w16970 & w16973;
assign w16975 = (w16974 & ~w2108) | (w16974 & w30834) | (~w2108 & w30834);
assign w16976 = (w2108 & w40916) | (w2108 & w40917) | (w40916 & w40917);
assign w16977 = (~w2108 & w40918) | (~w2108 & w40919) | (w40918 & w40919);
assign w16978 = ~w16975 & ~w16976;
assign w16979 = ~w16977 & ~w16978;
assign w16980 = w16969 & ~w16979;
assign w16981 = w16969 & ~w16980;
assign w16982 = ~w16969 & ~w16979;
assign w16983 = ~w16981 & ~w16982;
assign w16984 = (~w16657 & w16660) | (~w16657 & w30835) | (w16660 & w30835);
assign w16985 = w16983 & w16984;
assign w16986 = ~w16983 & ~w16984;
assign w16987 = ~w16985 & ~w16986;
assign w16988 = b_28 & w7613;
assign w16989 = w7941 & w30836;
assign w16990 = b_27 & w7608;
assign w16991 = ~w16989 & ~w16990;
assign w16992 = ~w16988 & w16991;
assign w16993 = (w16992 & ~w2771) | (w16992 & w30837) | (~w2771 & w30837);
assign w16994 = (w2771 & w40920) | (w2771 & w40921) | (w40920 & w40921);
assign w16995 = (~w2771 & w40922) | (~w2771 & w40923) | (w40922 & w40923);
assign w16996 = ~w16993 & ~w16994;
assign w16997 = ~w16995 & ~w16996;
assign w16998 = ~w16987 & w16997;
assign w16999 = w16987 & ~w16997;
assign w17000 = ~w16998 & ~w16999;
assign w17001 = ~w16909 & w17000;
assign w17002 = ~w16909 & ~w17001;
assign w17003 = w17000 & ~w17001;
assign w17004 = ~w17002 & ~w17003;
assign w17005 = ~w16908 & ~w17004;
assign w17006 = (w16908 & w17001) | (w16908 & w30838) | (w17001 & w30838);
assign w17007 = ~w17002 & w17006;
assign w17008 = ~w17005 & ~w17007;
assign w17009 = ~w16698 & w17008;
assign w17010 = w16698 & ~w17008;
assign w17011 = ~w17009 & ~w17010;
assign w17012 = ~w16898 & w17011;
assign w17013 = w16898 & ~w17011;
assign w17014 = ~w17012 & ~w17013;
assign w17015 = ~w16888 & w17014;
assign w17016 = ~w16888 & ~w17015;
assign w17017 = w17014 & ~w17015;
assign w17018 = ~w17016 & ~w17017;
assign w17019 = ~w16886 & ~w17018;
assign w17020 = (w16886 & w17015) | (w16886 & w30839) | (w17015 & w30839);
assign w17021 = ~w17016 & w17020;
assign w17022 = ~w17019 & ~w17021;
assign w17023 = ~w17019 & w30840;
assign w17024 = ~w16876 & ~w17023;
assign w17025 = w17022 & ~w17023;
assign w17026 = ~w17024 & ~w17025;
assign w17027 = ~w16875 & ~w17026;
assign w17028 = w16875 & ~w17025;
assign w17029 = ~w17024 & w17028;
assign w17030 = ~w17027 & ~w17029;
assign w17031 = ~w16865 & w17030;
assign w17032 = w16865 & ~w17030;
assign w17033 = ~w17031 & ~w17032;
assign w17034 = ~w16863 & w17033;
assign w17035 = w17033 & ~w17034;
assign w17036 = ~w17033 & ~w16863;
assign w17037 = ~w17035 & ~w17036;
assign w17038 = b_46 & w3195;
assign w17039 = w3388 & w30841;
assign w17040 = b_45 & w3190;
assign w17041 = ~w17039 & ~w17040;
assign w17042 = ~w17038 & w17041;
assign w17043 = w17041 & w30842;
assign w17044 = (~w6974 & w26687) | (~w6974 & w26688) | (w26687 & w26688);
assign w17045 = (w6974 & w26689) | (w6974 & w26690) | (w26689 & w26690);
assign w17046 = ~w17044 & ~w17045;
assign w17047 = (~w17046 & w16763) | (~w17046 & w30843) | (w16763 & w30843);
assign w17048 = (w17046 & w16763) | (w17046 & w30844) | (w16763 & w30844);
assign w17049 = ~w16763 & w40924;
assign w17050 = ~w17048 & ~w17049;
assign w17051 = ~w27599 & w30845;
assign w17052 = (~w27599 & w30846) | (~w27599 & w30847) | (w30846 & w30847);
assign w17053 = ~w17051 & ~w17052;
assign w17054 = (~w17053 & w16852) | (~w17053 & w30848) | (w16852 & w30848);
assign w17055 = ~w16853 & ~w17054;
assign w17056 = ~w30848 & w40925;
assign w17057 = ~w17055 & ~w17056;
assign w17058 = ~w16564 & ~w16574;
assign w17059 = b_52 & w2158;
assign w17060 = w2294 & w30850;
assign w17061 = b_51 & w2153;
assign w17062 = ~w17060 & ~w17061;
assign w17063 = ~w17059 & w17062;
assign w17064 = w17062 & w30851;
assign w17065 = (~w8793 & w40926) | (~w8793 & w40927) | (w40926 & w40927);
assign w17066 = (w8793 & w30853) | (w8793 & w30854) | (w30853 & w30854);
assign w17067 = ~w17065 & ~w17066;
assign w17068 = (~w16577 & w40928) | (~w16577 & w40929) | (w40928 & w40929);
assign w17069 = (w16577 & w40930) | (w16577 & w40931) | (w40930 & w40931);
assign w17070 = ~w17068 & ~w17069;
assign w17071 = ~w17057 & w17070;
assign w17072 = ~w17070 & ~w17057;
assign w17073 = w17070 & ~w17071;
assign w17074 = ~w17072 & ~w17073;
assign w17075 = (~w17074 & w16837) | (~w17074 & w30855) | (w16837 & w30855);
assign w17076 = ~w16838 & ~w17075;
assign w17077 = ~w16837 & w40932;
assign w17078 = ~w17076 & ~w17077;
assign w17079 = (~w16546 & ~w16786) | (~w16546 & w30856) | (~w16786 & w30856);
assign w17080 = b_58 & w1295;
assign w17081 = w1422 & w30857;
assign w17082 = b_57 & w1290;
assign w17083 = ~w17081 & ~w17082;
assign w17084 = ~w17080 & w17083;
assign w17085 = w17083 & w30858;
assign w17086 = (~w10476 & w40933) | (~w10476 & w40934) | (w40933 & w40934);
assign w17087 = (w10476 & w30860) | (w10476 & w30861) | (w30860 & w30861);
assign w17088 = ~w17086 & ~w17087;
assign w17089 = (w16786 & w30862) | (w16786 & w30863) | (w30862 & w30863);
assign w17090 = ~w17079 & ~w17089;
assign w17091 = (~w16786 & w40935) | (~w16786 & w40936) | (w40935 & w40936);
assign w17092 = ~w17090 & ~w17091;
assign w17093 = (~w17078 & w17090) | (~w17078 & w40937) | (w17090 & w40937);
assign w17094 = ~w17090 & w40938;
assign w17095 = ~w17092 & ~w17093;
assign w17096 = ~w17094 & ~w17095;
assign w17097 = (~w17096 & w16822) | (~w17096 & w30864) | (w16822 & w30864);
assign w17098 = ~w16823 & ~w17097;
assign w17099 = ~w17096 & ~w17097;
assign w17100 = ~w17098 & ~w17099;
assign w17101 = (~w16518 & w16477) | (~w16518 & w30865) | (w16477 & w30865);
assign w17102 = (~w17101 & w16521) | (~w17101 & w40939) | (w16521 & w40939);
assign w17103 = w754 & w30866;
assign w17104 = b_63 & w652;
assign w17105 = ~w17103 & ~w17104;
assign w17106 = ~w12671 & w30867;
assign w17107 = (a_14 & w17106) | (a_14 & w30868) | (w17106 & w30868);
assign w17108 = ~w17106 & w30869;
assign w17109 = ~w17107 & ~w17108;
assign w17110 = (~w17109 & w16793) | (~w17109 & w30870) | (w16793 & w30870);
assign w17111 = ~w17102 & ~w17110;
assign w17112 = ~w16793 & w30871;
assign w17113 = ~w17111 & ~w17112;
assign w17114 = (~w17100 & w17111) | (~w17100 & w40940) | (w17111 & w40940);
assign w17115 = w17100 & ~w17112;
assign w17116 = ~w17111 & w17115;
assign w17117 = ~w17114 & ~w17116;
assign w17118 = (w17117 & w16807) | (w17117 & w40941) | (w16807 & w40941);
assign w17119 = ~w16808 & ~w17118;
assign w17120 = ~w16807 & w40942;
assign w17121 = ~w17119 & ~w17120;
assign w17122 = (w14835 & w30872) | (w14835 & w30873) | (w30872 & w30873);
assign w17123 = (w13761 & w37686) | (w13761 & w37687) | (w37686 & w37687);
assign w17124 = ~w17122 & ~w17123;
assign w17125 = (~w17110 & w17113) | (~w17110 & w30876) | (w17113 & w30876);
assign w17126 = ~w16820 & ~w17097;
assign w17127 = w754 & w30877;
assign w17128 = (~w17127 & ~w12670) | (~w17127 & w30878) | (~w12670 & w30878);
assign w17129 = (w12670 & w40943) | (w12670 & w40944) | (w40943 & w40944);
assign w17130 = (~w12670 & w40945) | (~w12670 & w40946) | (w40945 & w40946);
assign w17131 = ~w17128 & ~w17129;
assign w17132 = ~w17130 & ~w17131;
assign w17133 = (~w17132 & w17097) | (~w17132 & w30879) | (w17097 & w30879);
assign w17134 = ~w17126 & ~w17133;
assign w17135 = ~w17097 & w30880;
assign w17136 = b_59 & w1295;
assign w17137 = w1422 & w30881;
assign w17138 = b_58 & w1290;
assign w17139 = ~w17137 & ~w17138;
assign w17140 = ~w17136 & w17139;
assign w17141 = (w17140 & ~w11169) | (w17140 & w30882) | (~w11169 & w30882);
assign w17142 = (w11169 & w40947) | (w11169 & w40948) | (w40947 & w40948);
assign w17143 = (~w11169 & w40949) | (~w11169 & w40950) | (w40949 & w40950);
assign w17144 = ~w17141 & ~w17142;
assign w17145 = ~w17143 & ~w17144;
assign w17146 = (~w16837 & w40951) | (~w16837 & w40952) | (w40951 & w40952);
assign w17147 = (w16837 & w40953) | (w16837 & w40954) | (w40953 & w40954);
assign w17148 = ~w17146 & ~w17147;
assign w17149 = b_56 & w1694;
assign w17150 = w1834 & w30885;
assign w17151 = b_55 & w1689;
assign w17152 = ~w17150 & ~w17151;
assign w17153 = ~w17149 & w17152;
assign w17154 = (w17153 & ~w9798) | (w17153 & w26375) | (~w9798 & w26375);
assign w17155 = (w9798 & w30886) | (w9798 & w30887) | (w30886 & w30887);
assign w17156 = (~w9798 & w30888) | (~w9798 & w30889) | (w30888 & w30889);
assign w17157 = ~w17154 & ~w17155;
assign w17158 = ~w17156 & ~w17157;
assign w17159 = (~w17068 & ~w17070) | (~w17068 & w30890) | (~w17070 & w30890);
assign w17160 = w17158 & w17159;
assign w17161 = ~w17158 & ~w17159;
assign w17162 = ~w17160 & ~w17161;
assign w17163 = b_53 & w2158;
assign w17164 = w2294 & w30891;
assign w17165 = b_52 & w2153;
assign w17166 = ~w17164 & ~w17165;
assign w17167 = ~w17163 & w17166;
assign w17168 = (w9109 & w40955) | (w9109 & w40956) | (w40955 & w40956);
assign w17169 = a_26 & ~w17168;
assign w17170 = w17168 & a_26;
assign w17171 = ~w17168 & ~w17169;
assign w17172 = ~w17170 & ~w17171;
assign w17173 = (~w30848 & w40957) | (~w30848 & w40958) | (w40957 & w40958);
assign w17174 = (w30848 & w40959) | (w30848 & w40960) | (w40959 & w40960);
assign w17175 = ~w17173 & ~w17174;
assign w17176 = b_47 & w3195;
assign w17177 = w3388 & w30896;
assign w17178 = b_46 & w3190;
assign w17179 = ~w17177 & ~w17178;
assign w17180 = ~w17176 & w17179;
assign w17181 = w17179 & w30897;
assign w17182 = (~w6998 & w25671) | (~w6998 & w25672) | (w25671 & w25672);
assign w17183 = (w6998 & w25673) | (w6998 & w25674) | (w25673 & w25674);
assign w17184 = ~w17182 & ~w17183;
assign w17185 = (w17033 & w40961) | (w17033 & w40962) | (w40961 & w40962);
assign w17186 = (~w17033 & w40963) | (~w17033 & w40964) | (w40963 & w40964);
assign w17187 = ~w17185 & ~w17186;
assign w17188 = b_44 & w3803;
assign w17189 = w4027 & w30898;
assign w17190 = b_43 & w3798;
assign w17191 = ~w17189 & ~w17190;
assign w17192 = ~w17188 & w17191;
assign w17193 = (w17192 & ~w6408) | (w17192 & w30899) | (~w6408 & w30899);
assign w17194 = (w6408 & w40965) | (w6408 & w40966) | (w40965 & w40966);
assign w17195 = (~w6408 & w40967) | (~w6408 & w40968) | (w40967 & w40968);
assign w17196 = ~w17193 & ~w17194;
assign w17197 = ~w17195 & ~w17196;
assign w17198 = (~w17023 & w17026) | (~w17023 & w30900) | (w17026 & w30900);
assign w17199 = b_41 & w4499;
assign w17200 = w4723 & w30901;
assign w17201 = b_40 & w4494;
assign w17202 = ~w17200 & ~w17201;
assign w17203 = ~w17199 & w17202;
assign w17204 = (w17203 & ~w5609) | (w17203 & w30902) | (~w5609 & w30902);
assign w17205 = (w5609 & w40969) | (w5609 & w40970) | (w40969 & w40970);
assign w17206 = (~w5609 & w40971) | (~w5609 & w40972) | (w40971 & w40972);
assign w17207 = ~w17204 & ~w17205;
assign w17208 = ~w17206 & ~w17207;
assign w17209 = (~w17015 & w17018) | (~w17015 & w30903) | (w17018 & w30903);
assign w17210 = (~w17001 & w17004) | (~w17001 & w30904) | (w17004 & w30904);
assign w17211 = (~w16968 & ~w16969) | (~w16968 & w30905) | (~w16969 & w30905);
assign w17212 = b_26 & w8526;
assign w17213 = w8886 & w30906;
assign w17214 = b_25 & w8521;
assign w17215 = ~w17213 & ~w17214;
assign w17216 = ~w17212 & w17215;
assign w17217 = (w17216 & ~w2416) | (w17216 & w30907) | (~w2416 & w30907);
assign w17218 = (w2416 & w40973) | (w2416 & w40974) | (w40973 & w40974);
assign w17219 = (~w2416 & w40975) | (~w2416 & w40976) | (w40975 & w40976);
assign w17220 = ~w17217 & ~w17218;
assign w17221 = ~w17219 & ~w17220;
assign w17222 = (~w16950 & ~w16951) | (~w16950 & w30908) | (~w16951 & w30908);
assign w17223 = (~w16918 & w16926) | (~w16918 & w30909) | (w16926 & w30909);
assign w17224 = ~w16915 & ~w17223;
assign w17225 = w12380 & w30910;
assign w17226 = b_14 & ~w12380;
assign w17227 = ~w17225 & ~w17226;
assign w17228 = w16912 & ~w17227;
assign w17229 = ~w16912 & w17227;
assign w17230 = ~w17228 & ~w17229;
assign w17231 = b_17 & w11620;
assign w17232 = w11969 & w30911;
assign w17233 = b_16 & w11615;
assign w17234 = ~w17232 & ~w17233;
assign w17235 = ~w17231 & w17234;
assign w17236 = w17234 & w30912;
assign w17237 = (~w1038 & w40977) | (~w1038 & w40978) | (w40977 & w40978);
assign w17238 = (w17230 & w17237) | (w17230 & w30915) | (w17237 & w30915);
assign w17239 = ~w17237 & w30916;
assign w17240 = ~w17238 & ~w17239;
assign w17241 = ~w17224 & w17240;
assign w17242 = w17224 & ~w17240;
assign w17243 = ~w17241 & ~w17242;
assign w17244 = b_20 & w10562;
assign w17245 = w10902 & w30917;
assign w17246 = b_19 & w10557;
assign w17247 = ~w17245 & ~w17246;
assign w17248 = ~w17244 & w17247;
assign w17249 = (w17248 & ~w1503) | (w17248 & w30918) | (~w1503 & w30918);
assign w17250 = (w1503 & w40979) | (w1503 & w40980) | (w40979 & w40980);
assign w17251 = (~w1503 & w40981) | (~w1503 & w40982) | (w40981 & w40982);
assign w17252 = ~w17249 & ~w17250;
assign w17253 = ~w17251 & ~w17252;
assign w17254 = w17243 & ~w17253;
assign w17255 = w17243 & ~w17254;
assign w17256 = ~w17243 & ~w17253;
assign w17257 = ~w17255 & ~w17256;
assign w17258 = (~w16932 & ~w16933) | (~w16932 & w30919) | (~w16933 & w30919);
assign w17259 = w17257 & w17258;
assign w17260 = ~w17257 & ~w17258;
assign w17261 = ~w17259 & ~w17260;
assign w17262 = b_23 & w9534;
assign w17263 = w9876 & w30920;
assign w17264 = b_22 & w9529;
assign w17265 = ~w17263 & ~w17264;
assign w17266 = ~w17262 & w17265;
assign w17267 = (w17266 & ~w1933) | (w17266 & w30921) | (~w1933 & w30921);
assign w17268 = (w1933 & w40983) | (w1933 & w40984) | (w40983 & w40984);
assign w17269 = (~w1933 & w40985) | (~w1933 & w40986) | (w40985 & w40986);
assign w17270 = ~w17267 & ~w17268;
assign w17271 = ~w17269 & ~w17270;
assign w17272 = ~w17261 & w17271;
assign w17273 = w17261 & ~w17271;
assign w17274 = ~w17272 & ~w17273;
assign w17275 = ~w17222 & w17274;
assign w17276 = w17222 & ~w17274;
assign w17277 = ~w17275 & ~w17276;
assign w17278 = ~w17221 & w17277;
assign w17279 = w17221 & ~w17277;
assign w17280 = ~w17278 & ~w17279;
assign w17281 = ~w17211 & w17280;
assign w17282 = w17211 & ~w17280;
assign w17283 = ~w17281 & ~w17282;
assign w17284 = b_29 & w7613;
assign w17285 = w7941 & w30922;
assign w17286 = b_28 & w7608;
assign w17287 = ~w17285 & ~w17286;
assign w17288 = ~w17284 & w17287;
assign w17289 = (w17288 & ~w2954) | (w17288 & w30923) | (~w2954 & w30923);
assign w17290 = (w2954 & w40987) | (w2954 & w40988) | (w40987 & w40988);
assign w17291 = (~w2954 & w40989) | (~w2954 & w40990) | (w40989 & w40990);
assign w17292 = ~w17289 & ~w17290;
assign w17293 = ~w17291 & ~w17292;
assign w17294 = w17283 & ~w17293;
assign w17295 = w17283 & ~w17294;
assign w17296 = ~w17283 & ~w17293;
assign w17297 = ~w17295 & ~w17296;
assign w17298 = (~w16986 & ~w16987) | (~w16986 & w30924) | (~w16987 & w30924);
assign w17299 = ~w17297 & ~w17298;
assign w17300 = ~w17297 & ~w17299;
assign w17301 = ~w17298 & ~w17299;
assign w17302 = ~w17300 & ~w17301;
assign w17303 = b_32 & w6761;
assign w17304 = w7075 & w30925;
assign w17305 = b_31 & w6756;
assign w17306 = ~w17304 & ~w17305;
assign w17307 = ~w17303 & w17306;
assign w17308 = (w17307 & ~w3545) | (w17307 & w30926) | (~w3545 & w30926);
assign w17309 = (w3545 & w40991) | (w3545 & w40992) | (w40991 & w40992);
assign w17310 = (~w3545 & w40993) | (~w3545 & w40994) | (w40993 & w40994);
assign w17311 = ~w17308 & ~w17309;
assign w17312 = ~w17310 & ~w17311;
assign w17313 = ~w17302 & w17312;
assign w17314 = w17302 & ~w17312;
assign w17315 = ~w17313 & ~w17314;
assign w17316 = w17210 & w17315;
assign w17317 = ~w17210 & ~w17315;
assign w17318 = ~w17316 & ~w17317;
assign w17319 = b_35 & w5962;
assign w17320 = w6246 & w30927;
assign w17321 = b_34 & w5957;
assign w17322 = ~w17320 & ~w17321;
assign w17323 = ~w17319 & w17322;
assign w17324 = (w17323 & ~w4181) | (w17323 & w30928) | (~w4181 & w30928);
assign w17325 = (w4181 & w40995) | (w4181 & w40996) | (w40995 & w40996);
assign w17326 = (~w4181 & w40997) | (~w4181 & w40998) | (w40997 & w40998);
assign w17327 = ~w17324 & ~w17325;
assign w17328 = ~w17326 & ~w17327;
assign w17329 = w17318 & ~w17328;
assign w17330 = w17318 & ~w17329;
assign w17331 = ~w17318 & ~w17328;
assign w17332 = ~w17330 & ~w17331;
assign w17333 = (~w17009 & ~w17011) | (~w17009 & w30929) | (~w17011 & w30929);
assign w17334 = w17332 & w17333;
assign w17335 = ~w17332 & ~w17333;
assign w17336 = ~w17334 & ~w17335;
assign w17337 = b_38 & w5196;
assign w17338 = w5459 & w30930;
assign w17339 = b_37 & w5191;
assign w17340 = ~w17338 & ~w17339;
assign w17341 = ~w17337 & w17340;
assign w17342 = (w17341 & ~w4658) | (w17341 & w30931) | (~w4658 & w30931);
assign w17343 = (w4658 & w40999) | (w4658 & w41000) | (w40999 & w41000);
assign w17344 = (~w4658 & w41001) | (~w4658 & w41002) | (w41001 & w41002);
assign w17345 = ~w17342 & ~w17343;
assign w17346 = ~w17344 & ~w17345;
assign w17347 = ~w17336 & w17346;
assign w17348 = w17336 & ~w17346;
assign w17349 = ~w17347 & ~w17348;
assign w17350 = ~w17209 & w17349;
assign w17351 = w17209 & ~w17349;
assign w17352 = ~w17350 & ~w17351;
assign w17353 = ~w17208 & w17352;
assign w17354 = w17208 & ~w17352;
assign w17355 = ~w17353 & ~w17354;
assign w17356 = ~w17198 & w17355;
assign w17357 = w17198 & ~w17355;
assign w17358 = ~w17356 & ~w17357;
assign w17359 = ~w17197 & w17358;
assign w17360 = ~w17358 & ~w17197;
assign w17361 = w17358 & ~w17359;
assign w17362 = ~w17360 & ~w17361;
assign w17363 = w17187 & ~w17362;
assign w17364 = w17187 & ~w17363;
assign w17365 = ~w17187 & ~w17362;
assign w17366 = ~w17364 & ~w17365;
assign w17367 = (~w27599 & w30932) | (~w27599 & w30933) | (w30932 & w30933);
assign w17368 = b_50 & w2639;
assign w17369 = w2820 & w30934;
assign w17370 = b_49 & w2634;
assign w17371 = ~w17369 & ~w17370;
assign w17372 = ~w17368 & w17371;
assign w17373 = w17371 & w30935;
assign w17374 = (~w8162 & w27600) | (~w8162 & w27601) | (w27600 & w27601);
assign w17375 = (w8162 & w27602) | (w8162 & w27603) | (w27602 & w27603);
assign w17376 = ~w17374 & ~w17375;
assign w17377 = ~w17367 & ~w17376;
assign w17378 = w17367 & w17376;
assign w17379 = ~w17377 & ~w17378;
assign w17380 = ~w17366 & w17379;
assign w17381 = ~w17379 & ~w17366;
assign w17382 = w17379 & ~w17380;
assign w17383 = ~w17381 & ~w17382;
assign w17384 = w17175 & ~w17383;
assign w17385 = w17175 & ~w17384;
assign w17386 = ~w17383 & ~w17384;
assign w17387 = ~w17385 & ~w17386;
assign w17388 = w17162 & ~w17387;
assign w17389 = ~w17162 & w17387;
assign w17390 = w17148 & w30936;
assign w17391 = w17148 & ~w17390;
assign w17392 = w30936 & ~w17148;
assign w17393 = ~w17391 & ~w17392;
assign w17394 = (~w17089 & w17092) | (~w17089 & w27776) | (w17092 & w27776);
assign w17395 = b_62 & w986;
assign w17396 = w1069 & w30937;
assign w17397 = b_61 & w981;
assign w17398 = ~w17396 & ~w17397;
assign w17399 = ~w17395 & w17398;
assign w17400 = w17398 & w30938;
assign w17401 = (~w12273 & w41003) | (~w12273 & w41004) | (w41003 & w41004);
assign w17402 = (w12273 & w30940) | (w12273 & w30941) | (w30940 & w30941);
assign w17403 = ~w17401 & ~w17402;
assign w17404 = (~w17092 & w30942) | (~w17092 & w30943) | (w30942 & w30943);
assign w17405 = ~w17394 & ~w17404;
assign w17406 = ~w17403 & ~w17404;
assign w17407 = ~w17405 & ~w17406;
assign w17408 = ~w17393 & ~w17407;
assign w17409 = (w17393 & w17404) | (w17393 & w30944) | (w17404 & w30944);
assign w17410 = ~w17405 & w17409;
assign w17411 = ~w17408 & ~w17410;
assign w17412 = (w17411 & w17134) | (w17411 & w30945) | (w17134 & w30945);
assign w17413 = ~w17134 & w30946;
assign w17414 = ~w17412 & ~w17413;
assign w17415 = ~w17125 & w17414;
assign w17416 = w17125 & ~w17414;
assign w17417 = ~w17415 & ~w17416;
assign w17418 = (w14835 & w30947) | (w14835 & w30948) | (w30947 & w30948);
assign w17419 = (~w14835 & w30949) | (~w14835 & w30950) | (w30949 & w30950);
assign w17420 = ~w17418 & ~w17419;
assign w17421 = (~w17404 & w17407) | (~w17404 & w30951) | (w17407 & w30951);
assign w17422 = b_63 & w986;
assign w17423 = w1069 & w30952;
assign w17424 = b_62 & w981;
assign w17425 = ~w17423 & ~w17424;
assign w17426 = ~w17422 & w17425;
assign w17427 = (w17426 & ~w12646) | (w17426 & w30953) | (~w12646 & w30953);
assign w17428 = (w12646 & w41005) | (w12646 & w41006) | (w41005 & w41006);
assign w17429 = (~w12646 & w41007) | (~w12646 & w41008) | (w41007 & w41008);
assign w17430 = ~w17427 & ~w17428;
assign w17431 = ~w17429 & ~w17430;
assign w17432 = (~w17407 & w30954) | (~w17407 & w30955) | (w30954 & w30955);
assign w17433 = ~w17421 & ~w17432;
assign w17434 = ~w17431 & ~w17432;
assign w17435 = ~w17433 & ~w17434;
assign w17436 = b_60 & w1295;
assign w17437 = w1422 & w30956;
assign w17438 = b_59 & w1290;
assign w17439 = ~w17437 & ~w17438;
assign w17440 = ~w17436 & w17439;
assign w17441 = (w17440 & ~w11196) | (w17440 & w30957) | (~w11196 & w30957);
assign w17442 = (w11196 & w41009) | (w11196 & w41010) | (w41009 & w41010);
assign w17443 = (~w11196 & w41011) | (~w11196 & w41012) | (w41011 & w41012);
assign w17444 = ~w17441 & ~w17442;
assign w17445 = ~w17443 & ~w17444;
assign w17446 = (~w17147 & ~w17148) | (~w17147 & w30958) | (~w17148 & w30958);
assign w17447 = w17445 & w17446;
assign w17448 = ~w17445 & ~w17446;
assign w17449 = ~w17447 & ~w17448;
assign w17450 = (~w17161 & ~w17162) | (~w17161 & w30959) | (~w17162 & w30959);
assign w17451 = b_57 & w1694;
assign w17452 = w1834 & w30960;
assign w17453 = b_56 & w1689;
assign w17454 = ~w17452 & ~w17453;
assign w17455 = ~w17451 & w17454;
assign w17456 = (w17455 & ~w10452) | (w17455 & w30961) | (~w10452 & w30961);
assign w17457 = (w10452 & w41013) | (w10452 & w41014) | (w41013 & w41014);
assign w17458 = (~w10452 & w41015) | (~w10452 & w41016) | (w41015 & w41016);
assign w17459 = ~w17456 & ~w17457;
assign w17460 = ~w17458 & ~w17459;
assign w17461 = ~w17450 & w17460;
assign w17462 = w17450 & ~w17460;
assign w17463 = ~w17461 & ~w17462;
assign w17464 = b_54 & w2158;
assign w17465 = w2294 & w30962;
assign w17466 = b_53 & w2153;
assign w17467 = ~w17465 & ~w17466;
assign w17468 = ~w17464 & w17467;
assign w17469 = (w17468 & ~w9134) | (w17468 & w30963) | (~w9134 & w30963);
assign w17470 = (w9134 & w41017) | (w9134 & w41018) | (w41017 & w41018);
assign w17471 = (~w9134 & w41019) | (~w9134 & w41020) | (w41019 & w41020);
assign w17472 = ~w17469 & ~w17470;
assign w17473 = ~w17471 & ~w17472;
assign w17474 = ~w17384 & w30964;
assign w17475 = (~w17473 & w17384) | (~w17473 & w30965) | (w17384 & w30965);
assign w17476 = ~w17474 & ~w17475;
assign w17477 = b_51 & w2639;
assign w17478 = w2820 & w30966;
assign w17479 = b_50 & w2634;
assign w17480 = ~w17478 & ~w17479;
assign w17481 = ~w17477 & w17480;
assign w17482 = (w17481 & ~w8186) | (w17481 & w27604) | (~w8186 & w27604);
assign w17483 = (w8186 & w30967) | (w8186 & w30968) | (w30967 & w30968);
assign w17484 = (~w8186 & w30969) | (~w8186 & w30970) | (w30969 & w30970);
assign w17485 = ~w17482 & ~w17483;
assign w17486 = ~w17484 & ~w17485;
assign w17487 = (~w17377 & ~w17379) | (~w17377 & w30971) | (~w17379 & w30971);
assign w17488 = w17486 & w17487;
assign w17489 = ~w17486 & ~w17487;
assign w17490 = ~w17488 & ~w17489;
assign w17491 = (~w17350 & ~w17352) | (~w17350 & w30972) | (~w17352 & w30972);
assign w17492 = (~w17335 & ~w17336) | (~w17335 & w30973) | (~w17336 & w30973);
assign w17493 = (~w17317 & ~w17318) | (~w17317 & w30974) | (~w17318 & w30974);
assign w17494 = (~w17299 & w17302) | (~w17299 & w30975) | (w17302 & w30975);
assign w17495 = (~w17260 & ~w17261) | (~w17260 & w41021) | (~w17261 & w41021);
assign w17496 = w12380 & w30976;
assign w17497 = b_15 & ~w12380;
assign w17498 = ~w17496 & ~w17497;
assign w17499 = ~a_14 & ~w17498;
assign w17500 = w17498 & ~a_14;
assign w17501 = ~w17498 & ~w17499;
assign w17502 = ~w17500 & ~w17501;
assign w17503 = (~w16912 & w17501) | (~w16912 & w30977) | (w17501 & w30977);
assign w17504 = ~w16912 & ~w17503;
assign w17505 = ~w17502 & ~w17503;
assign w17506 = ~w17504 & ~w17505;
assign w17507 = b_18 & w11620;
assign w17508 = w11969 & w30978;
assign w17509 = b_17 & w11615;
assign w17510 = ~w17508 & ~w17509;
assign w17511 = ~w17507 & w17510;
assign w17512 = (w17511 & ~w1238) | (w17511 & w30979) | (~w1238 & w30979);
assign w17513 = (w1238 & w41022) | (w1238 & w41023) | (w41022 & w41023);
assign w17514 = (~w1238 & w41024) | (~w1238 & w41025) | (w41024 & w41025);
assign w17515 = ~w17512 & ~w17513;
assign w17516 = ~w17514 & ~w17515;
assign w17517 = (~w17506 & w17515) | (~w17506 & w30980) | (w17515 & w30980);
assign w17518 = ~w17506 & ~w17517;
assign w17519 = ~w17516 & ~w17517;
assign w17520 = ~w17518 & ~w17519;
assign w17521 = ~w17228 & ~w17238;
assign w17522 = w17520 & w17521;
assign w17523 = ~w17520 & ~w17521;
assign w17524 = ~w17522 & ~w17523;
assign w17525 = b_21 & w10562;
assign w17526 = w10902 & w30981;
assign w17527 = b_20 & w10557;
assign w17528 = ~w17526 & ~w17527;
assign w17529 = ~w17525 & w17528;
assign w17530 = (w17529 & ~w1634) | (w17529 & w30982) | (~w1634 & w30982);
assign w17531 = (w1634 & w41026) | (w1634 & w41027) | (w41026 & w41027);
assign w17532 = (~w1634 & w41028) | (~w1634 & w41029) | (w41028 & w41029);
assign w17533 = ~w17530 & ~w17531;
assign w17534 = ~w17532 & ~w17533;
assign w17535 = w17524 & ~w17534;
assign w17536 = w17524 & ~w17535;
assign w17537 = ~w17524 & ~w17534;
assign w17538 = (~w17241 & ~w17243) | (~w17241 & w30983) | (~w17243 & w30983);
assign w17539 = ~w17536 & w30984;
assign w17540 = (~w17538 & w17536) | (~w17538 & w30985) | (w17536 & w30985);
assign w17541 = ~w17539 & ~w17540;
assign w17542 = b_24 & w9534;
assign w17543 = w9876 & w30986;
assign w17544 = b_23 & w9529;
assign w17545 = ~w17543 & ~w17544;
assign w17546 = ~w17542 & w17545;
assign w17547 = (w17546 & ~w2083) | (w17546 & w30987) | (~w2083 & w30987);
assign w17548 = (w2083 & w41030) | (w2083 & w41031) | (w41030 & w41031);
assign w17549 = (~w2083 & w41032) | (~w2083 & w41033) | (w41032 & w41033);
assign w17550 = ~w17547 & ~w17548;
assign w17551 = ~w17549 & ~w17550;
assign w17552 = w17541 & ~w17551;
assign w17553 = ~w17541 & w17551;
assign w17554 = ~w17495 & w30988;
assign w17555 = ~w30988 & ~w17495;
assign w17556 = (~w17552 & ~w30988) | (~w17552 & w41034) | (~w30988 & w41034);
assign w17557 = ~w17554 & w30988;
assign w17558 = ~w17555 & ~w17557;
assign w17559 = b_27 & w8526;
assign w17560 = w8886 & w30989;
assign w17561 = b_26 & w8521;
assign w17562 = ~w17560 & ~w17561;
assign w17563 = ~w17559 & w17562;
assign w17564 = (w17563 & ~w2582) | (w17563 & w30990) | (~w2582 & w30990);
assign w17565 = (w2582 & w41035) | (w2582 & w41036) | (w41035 & w41036);
assign w17566 = (~w2582 & w41037) | (~w2582 & w41038) | (w41037 & w41038);
assign w17567 = ~w17564 & ~w17565;
assign w17568 = ~w17566 & ~w17567;
assign w17569 = (~w17568 & w17557) | (~w17568 & w41039) | (w17557 & w41039);
assign w17570 = ~w17558 & ~w17569;
assign w17571 = ~w17557 & w41040;
assign w17572 = (~w17275 & ~w17277) | (~w17275 & w30991) | (~w17277 & w30991);
assign w17573 = ~w17570 & w30992;
assign w17574 = (~w17572 & w17570) | (~w17572 & w30993) | (w17570 & w30993);
assign w17575 = ~w17573 & ~w17574;
assign w17576 = b_30 & w7613;
assign w17577 = w7941 & w30994;
assign w17578 = b_29 & w7608;
assign w17579 = ~w17577 & ~w17578;
assign w17580 = ~w17576 & w17579;
assign w17581 = (w17580 & ~w3138) | (w17580 & w30995) | (~w3138 & w30995);
assign w17582 = (w3138 & w41041) | (w3138 & w41042) | (w41041 & w41042);
assign w17583 = (~w3138 & w41043) | (~w3138 & w41044) | (w41043 & w41044);
assign w17584 = ~w17581 & ~w17582;
assign w17585 = ~w17583 & ~w17584;
assign w17586 = w17575 & ~w17585;
assign w17587 = w17575 & ~w17586;
assign w17588 = ~w17575 & ~w17585;
assign w17589 = (~w17281 & ~w17283) | (~w17281 & w30996) | (~w17283 & w30996);
assign w17590 = ~w17587 & w30997;
assign w17591 = (~w17589 & w17587) | (~w17589 & w30998) | (w17587 & w30998);
assign w17592 = ~w17590 & ~w17591;
assign w17593 = b_33 & w6761;
assign w17594 = w7075 & w30999;
assign w17595 = b_32 & w6756;
assign w17596 = ~w17594 & ~w17595;
assign w17597 = ~w17593 & w17596;
assign w17598 = (w17597 & ~w3744) | (w17597 & w31000) | (~w3744 & w31000);
assign w17599 = (w3744 & w41045) | (w3744 & w41046) | (w41045 & w41046);
assign w17600 = (~w3744 & w41047) | (~w3744 & w41048) | (w41047 & w41048);
assign w17601 = ~w17598 & ~w17599;
assign w17602 = ~w17600 & ~w17601;
assign w17603 = w17592 & ~w17602;
assign w17604 = w17592 & ~w17603;
assign w17605 = ~w17592 & ~w17602;
assign w17606 = ~w17604 & ~w17605;
assign w17607 = ~w17494 & w17606;
assign w17608 = w17494 & ~w17606;
assign w17609 = ~w17607 & ~w17608;
assign w17610 = b_36 & w5962;
assign w17611 = w6246 & w31001;
assign w17612 = b_35 & w5957;
assign w17613 = ~w17611 & ~w17612;
assign w17614 = ~w17610 & w17613;
assign w17615 = (w17614 & ~w4395) | (w17614 & w31002) | (~w4395 & w31002);
assign w17616 = (w4395 & w41049) | (w4395 & w41050) | (w41049 & w41050);
assign w17617 = (~w4395 & w41051) | (~w4395 & w41052) | (w41051 & w41052);
assign w17618 = ~w17615 & ~w17616;
assign w17619 = ~w17617 & ~w17618;
assign w17620 = ~w17609 & ~w17619;
assign w17621 = w17609 & w17619;
assign w17622 = ~w17620 & ~w17621;
assign w17623 = w17493 & ~w17622;
assign w17624 = ~w17493 & w17622;
assign w17625 = ~w17623 & ~w17624;
assign w17626 = b_39 & w5196;
assign w17627 = w5459 & w31003;
assign w17628 = b_38 & w5191;
assign w17629 = ~w17627 & ~w17628;
assign w17630 = ~w17626 & w17629;
assign w17631 = (w17630 & ~w4888) | (w17630 & w31004) | (~w4888 & w31004);
assign w17632 = (w4888 & w41053) | (w4888 & w41054) | (w41053 & w41054);
assign w17633 = (~w4888 & w41055) | (~w4888 & w41056) | (w41055 & w41056);
assign w17634 = ~w17631 & ~w17632;
assign w17635 = ~w17633 & ~w17634;
assign w17636 = w17625 & ~w17635;
assign w17637 = w17625 & ~w17636;
assign w17638 = ~w17625 & ~w17635;
assign w17639 = ~w17637 & ~w17638;
assign w17640 = ~w17492 & w17639;
assign w17641 = w17492 & ~w17639;
assign w17642 = ~w17640 & ~w17641;
assign w17643 = b_42 & w4499;
assign w17644 = w4723 & w31005;
assign w17645 = b_41 & w4494;
assign w17646 = ~w17644 & ~w17645;
assign w17647 = ~w17643 & w17646;
assign w17648 = (w17647 & ~w5864) | (w17647 & w31006) | (~w5864 & w31006);
assign w17649 = (w5864 & w41057) | (w5864 & w41058) | (w41057 & w41058);
assign w17650 = (~w5864 & w41059) | (~w5864 & w41060) | (w41059 & w41060);
assign w17651 = ~w17648 & ~w17649;
assign w17652 = ~w17650 & ~w17651;
assign w17653 = ~w17642 & ~w17652;
assign w17654 = w17642 & w17652;
assign w17655 = ~w17653 & ~w17654;
assign w17656 = w17491 & ~w17655;
assign w17657 = ~w17491 & w17655;
assign w17658 = ~w17656 & ~w17657;
assign w17659 = b_45 & w3803;
assign w17660 = w4027 & w31007;
assign w17661 = b_44 & w3798;
assign w17662 = ~w17660 & ~w17661;
assign w17663 = ~w17659 & w17662;
assign w17664 = (w17663 & ~w6682) | (w17663 & w26691) | (~w6682 & w26691);
assign w17665 = (w6682 & w27605) | (w6682 & w27606) | (w27605 & w27606);
assign w17666 = (~w6682 & w31008) | (~w6682 & w31009) | (w31008 & w31009);
assign w17667 = ~w17664 & ~w17665;
assign w17668 = ~w17666 & ~w17667;
assign w17669 = w17658 & ~w17668;
assign w17670 = w17658 & ~w17669;
assign w17671 = ~w17658 & ~w17668;
assign w17672 = ~w17670 & ~w17671;
assign w17673 = (~w17356 & ~w17358) | (~w17356 & w31010) | (~w17358 & w31010);
assign w17674 = w17672 & w17673;
assign w17675 = ~w17672 & ~w17673;
assign w17676 = ~w17674 & ~w17675;
assign w17677 = (~w17185 & ~w17187) | (~w17185 & w25997) | (~w17187 & w25997);
assign w17678 = b_48 & w3195;
assign w17679 = w3388 & w31011;
assign w17680 = b_47 & w3190;
assign w17681 = ~w17679 & ~w17680;
assign w17682 = ~w17678 & w17681;
assign w17683 = (w17682 & ~w7284) | (w17682 & w25998) | (~w7284 & w25998);
assign w17684 = (w7284 & w26377) | (w7284 & w26378) | (w26377 & w26378);
assign w17685 = (~w7284 & w31012) | (~w7284 & w31013) | (w31012 & w31013);
assign w17686 = ~w17683 & ~w17684;
assign w17687 = ~w17685 & ~w17686;
assign w17688 = (~w25997 & w41061) | (~w25997 & w41062) | (w41061 & w41062);
assign w17689 = ~w17677 & ~w17688;
assign w17690 = (w17676 & w17689) | (w17676 & w26379) | (w17689 & w26379);
assign w17691 = ~w17689 & w31014;
assign w17692 = w17490 & w31015;
assign w17693 = w17490 & ~w17692;
assign w17694 = w31015 & ~w17490;
assign w17695 = ~w17693 & ~w17694;
assign w17696 = w17476 & ~w17695;
assign w17697 = ~w17476 & w17695;
assign w17698 = ~w17463 & w31016;
assign w17699 = ~w17463 & ~w17698;
assign w17700 = w31016 & w17463;
assign w17701 = ~w17699 & ~w17700;
assign w17702 = w17449 & ~w17701;
assign w17703 = ~w17449 & w17701;
assign w17704 = ~w17435 & w31017;
assign w17705 = ~w17435 & ~w17704;
assign w17706 = w31017 & w17435;
assign w17707 = ~w17705 & ~w17706;
assign w17708 = ~w17133 & ~w17412;
assign w17709 = w17707 & w17708;
assign w17710 = ~w17707 & ~w17708;
assign w17711 = ~w17709 & ~w17710;
assign w17712 = (w14835 & w31019) | (w14835 & w31020) | (w31019 & w31020);
assign w17713 = (~w14835 & w31021) | (~w14835 & w31022) | (w31021 & w31022);
assign w17714 = ~w17712 & ~w17713;
assign w17715 = (~w17448 & ~w17449) | (~w17448 & w31023) | (~w17449 & w31023);
assign w17716 = w1069 & w31024;
assign w17717 = b_63 & w981;
assign w17718 = ~w17716 & ~w17717;
assign w17719 = ~w12671 & w31025;
assign w17720 = (a_17 & w17719) | (a_17 & w31026) | (w17719 & w31026);
assign w17721 = ~w17719 & w31027;
assign w17722 = ~w17720 & ~w17721;
assign w17723 = (~w31023 & w41063) | (~w31023 & w41064) | (w41063 & w41064);
assign w17724 = (w31023 & w41065) | (w31023 & w41066) | (w41065 & w41066);
assign w17725 = ~w17723 & ~w17724;
assign w17726 = b_61 & w1295;
assign w17727 = w1422 & w31028;
assign w17728 = b_60 & w1290;
assign w17729 = ~w17727 & ~w17728;
assign w17730 = ~w17726 & w17729;
assign w17731 = (w17730 & ~w11901) | (w17730 & w31029) | (~w11901 & w31029);
assign w17732 = (w11901 & w41067) | (w11901 & w41068) | (w41067 & w41068);
assign w17733 = (~w11901 & w41069) | (~w11901 & w41070) | (w41069 & w41070);
assign w17734 = ~w17731 & ~w17732;
assign w17735 = ~w17733 & ~w17734;
assign w17736 = ~w17450 & ~w17460;
assign w17737 = (w17463 & w41071) | (w17463 & w41072) | (w41071 & w41072);
assign w17738 = (~w17463 & w41073) | (~w17463 & w41074) | (w41073 & w41074);
assign w17739 = ~w17737 & ~w17738;
assign w17740 = b_58 & w1694;
assign w17741 = w1834 & w31031;
assign w17742 = b_57 & w1689;
assign w17743 = ~w17741 & ~w17742;
assign w17744 = ~w17740 & w17743;
assign w17745 = w17743 & w31032;
assign w17746 = (~w10476 & w41075) | (~w10476 & w41076) | (w41075 & w41076);
assign w17747 = (w10476 & w31034) | (w10476 & w31035) | (w31034 & w31035);
assign w17748 = ~w17746 & ~w17747;
assign w17749 = (~w17748 & w17696) | (~w17748 & w31036) | (w17696 & w31036);
assign w17750 = ~w17696 & w31037;
assign w17751 = ~w17749 & ~w17750;
assign w17752 = b_55 & w2158;
assign w17753 = w2294 & w31038;
assign w17754 = b_54 & w2153;
assign w17755 = ~w17753 & ~w17754;
assign w17756 = ~w17752 & w17755;
assign w17757 = (w17756 & ~w9776) | (w17756 & w31039) | (~w9776 & w31039);
assign w17758 = (w9776 & w41077) | (w9776 & w41078) | (w41077 & w41078);
assign w17759 = (~w9776 & w41079) | (~w9776 & w41080) | (w41079 & w41080);
assign w17760 = ~w17757 & ~w17758;
assign w17761 = ~w17759 & ~w17760;
assign w17762 = (~w17489 & ~w17490) | (~w17489 & w31040) | (~w17490 & w31040);
assign w17763 = w17761 & w17762;
assign w17764 = ~w17761 & ~w17762;
assign w17765 = ~w17763 & ~w17764;
assign w17766 = b_52 & w2639;
assign w17767 = w2820 & w31041;
assign w17768 = b_51 & w2634;
assign w17769 = ~w17767 & ~w17768;
assign w17770 = ~w17766 & w17769;
assign w17771 = (w17770 & ~w8793) | (w17770 & w25675) | (~w8793 & w25675);
assign w17772 = (w8793 & w25999) | (w8793 & w26000) | (w25999 & w26000);
assign w17773 = (~w8793 & w26380) | (~w8793 & w26381) | (w26380 & w26381);
assign w17774 = ~w17771 & ~w17772;
assign w17775 = ~w17773 & ~w17774;
assign w17776 = ~w17690 & w31042;
assign w17777 = (w17775 & w17690) | (w17775 & w31043) | (w17690 & w31043);
assign w17778 = ~w17776 & ~w17777;
assign w17779 = b_49 & w3195;
assign w17780 = w3388 & w31044;
assign w17781 = b_48 & w3190;
assign w17782 = ~w17780 & ~w17781;
assign w17783 = ~w17779 & w17782;
assign w17784 = (w17783 & ~w7859) | (w17783 & w26001) | (~w7859 & w26001);
assign w17785 = (w7859 & w26382) | (w7859 & w26383) | (w26382 & w26383);
assign w17786 = (~w7859 & w27607) | (~w7859 & w27608) | (w27607 & w27608);
assign w17787 = ~w17784 & ~w17785;
assign w17788 = ~w17786 & ~w17787;
assign w17789 = (~w17669 & w17672) | (~w17669 & w31045) | (w17672 & w31045);
assign w17790 = w17788 & w17789;
assign w17791 = ~w17788 & ~w17789;
assign w17792 = ~w17790 & ~w17791;
assign w17793 = b_43 & w4499;
assign w17794 = w4723 & w31046;
assign w17795 = b_42 & w4494;
assign w17796 = ~w17794 & ~w17795;
assign w17797 = ~w17793 & w17796;
assign w17798 = (w17797 & ~w5888) | (w17797 & w31047) | (~w5888 & w31047);
assign w17799 = (w5888 & w41081) | (w5888 & w41082) | (w41081 & w41082);
assign w17800 = (~w5888 & w41083) | (~w5888 & w41084) | (w41083 & w41084);
assign w17801 = ~w17798 & ~w17799;
assign w17802 = ~w17800 & ~w17801;
assign w17803 = ~w17492 & ~w17639;
assign w17804 = ~w17636 & ~w17803;
assign w17805 = b_40 & w5196;
assign w17806 = w5459 & w31048;
assign w17807 = b_39 & w5191;
assign w17808 = ~w17806 & ~w17807;
assign w17809 = ~w17805 & w17808;
assign w17810 = (w17809 & ~w5363) | (w17809 & w31049) | (~w5363 & w31049);
assign w17811 = (w5363 & w41085) | (w5363 & w41086) | (w41085 & w41086);
assign w17812 = (~w5363 & w41087) | (~w5363 & w41088) | (w41087 & w41088);
assign w17813 = ~w17810 & ~w17811;
assign w17814 = ~w17812 & ~w17813;
assign w17815 = ~w17620 & ~w17624;
assign w17816 = b_37 & w5962;
assign w17817 = w6246 & w31050;
assign w17818 = b_36 & w5957;
assign w17819 = ~w17817 & ~w17818;
assign w17820 = ~w17816 & w17819;
assign w17821 = (w17820 & ~w4636) | (w17820 & w31051) | (~w4636 & w31051);
assign w17822 = (w4636 & w41089) | (w4636 & w41090) | (w41089 & w41090);
assign w17823 = (~w4636 & w41091) | (~w4636 & w41092) | (w41091 & w41092);
assign w17824 = ~w17821 & ~w17822;
assign w17825 = ~w17823 & ~w17824;
assign w17826 = ~w17494 & ~w17606;
assign w17827 = ~w17603 & ~w17826;
assign w17828 = b_31 & w7613;
assign w17829 = w7941 & w31052;
assign w17830 = b_30 & w7608;
assign w17831 = ~w17829 & ~w17830;
assign w17832 = ~w17828 & w17831;
assign w17833 = (w17832 & ~w3345) | (w17832 & w31053) | (~w3345 & w31053);
assign w17834 = (w3345 & w41093) | (w3345 & w41094) | (w41093 & w41094);
assign w17835 = (~w3345 & w41095) | (~w3345 & w41096) | (w41095 & w41096);
assign w17836 = ~w17833 & ~w17834;
assign w17837 = ~w17835 & ~w17836;
assign w17838 = w12380 & w31055;
assign w17839 = b_16 & ~w12380;
assign w17840 = ~w17838 & ~w17839;
assign w17841 = ~w17503 & w31056;
assign w17842 = (w17840 & w17503) | (w17840 & w31057) | (w17503 & w31057);
assign w17843 = ~w17841 & ~w17842;
assign w17844 = b_19 & w11620;
assign w17845 = w11969 & w31058;
assign w17846 = b_18 & w11615;
assign w17847 = ~w17845 & ~w17846;
assign w17848 = ~w17844 & w17847;
assign w17849 = w17847 & w31059;
assign w17850 = (~w1372 & w41097) | (~w1372 & w41098) | (w41097 & w41098);
assign w17851 = (w17843 & w17850) | (w17843 & w31063) | (w17850 & w31063);
assign w17852 = ~w17850 & w31064;
assign w17853 = ~w17851 & ~w17852;
assign w17854 = (~w17520 & w31065) | (~w17520 & w31066) | (w31065 & w31066);
assign w17855 = (w17520 & w31067) | (w17520 & w31068) | (w31067 & w31068);
assign w17856 = ~w17854 & ~w17855;
assign w17857 = b_22 & w10562;
assign w17858 = w10902 & w31069;
assign w17859 = b_21 & w10557;
assign w17860 = ~w17858 & ~w17859;
assign w17861 = ~w17857 & w17860;
assign w17862 = (w17861 & ~w1786) | (w17861 & w31070) | (~w1786 & w31070);
assign w17863 = (w1786 & w41099) | (w1786 & w41100) | (w41099 & w41100);
assign w17864 = (~w1786 & w41101) | (~w1786 & w41102) | (w41101 & w41102);
assign w17865 = ~w17862 & ~w17863;
assign w17866 = ~w17864 & ~w17865;
assign w17867 = w17856 & ~w17866;
assign w17868 = w17856 & ~w17867;
assign w17869 = ~w17856 & ~w17866;
assign w17870 = ~w17868 & ~w17869;
assign w17871 = ~w17535 & ~w17540;
assign w17872 = w17870 & w17871;
assign w17873 = ~w17870 & ~w17871;
assign w17874 = ~w17872 & ~w17873;
assign w17875 = b_25 & w9534;
assign w17876 = w9876 & w31071;
assign w17877 = b_24 & w9529;
assign w17878 = ~w17876 & ~w17877;
assign w17879 = ~w17875 & w17878;
assign w17880 = (w17879 & ~w2108) | (w17879 & w31072) | (~w2108 & w31072);
assign w17881 = (w2108 & w41103) | (w2108 & w41104) | (w41103 & w41104);
assign w17882 = (~w2108 & w41105) | (~w2108 & w41106) | (w41105 & w41106);
assign w17883 = ~w17880 & ~w17881;
assign w17884 = ~w17882 & ~w17883;
assign w17885 = w17874 & ~w17884;
assign w17886 = w17874 & ~w17885;
assign w17887 = ~w17874 & ~w17884;
assign w17888 = ~w17886 & ~w17887;
assign w17889 = ~w17886 & w41107;
assign w17890 = (w17556 & w17886) | (w17556 & w41108) | (w17886 & w41108);
assign w17891 = ~w17889 & ~w17890;
assign w17892 = b_28 & w8526;
assign w17893 = w8886 & w31073;
assign w17894 = b_27 & w8521;
assign w17895 = ~w17893 & ~w17894;
assign w17896 = ~w17892 & w17895;
assign w17897 = (w17896 & ~w2771) | (w17896 & w31074) | (~w2771 & w31074);
assign w17898 = (w2771 & w41109) | (w2771 & w41110) | (w41109 & w41110);
assign w17899 = (~w2771 & w41111) | (~w2771 & w41112) | (w41111 & w41112);
assign w17900 = ~w17897 & ~w17898;
assign w17901 = ~w17899 & ~w17900;
assign w17902 = w17891 & w17901;
assign w17903 = ~w17891 & ~w17901;
assign w17904 = ~w17902 & ~w17903;
assign w17905 = (~w30993 & w41113) | (~w30993 & w41114) | (w41113 & w41114);
assign w17906 = w17904 & ~w17905;
assign w17907 = ~w17904 & w17905;
assign w17908 = ~w17906 & ~w17907;
assign w17909 = ~w17837 & w17908;
assign w17910 = w17908 & ~w17909;
assign w17911 = ~w17908 & ~w17837;
assign w17912 = ~w17910 & ~w17911;
assign w17913 = (~w30998 & w41115) | (~w30998 & w41116) | (w41115 & w41116);
assign w17914 = w17912 & w17913;
assign w17915 = ~w17912 & ~w17913;
assign w17916 = ~w17914 & ~w17915;
assign w17917 = b_34 & w6761;
assign w17918 = w7075 & w31075;
assign w17919 = b_33 & w6756;
assign w17920 = ~w17918 & ~w17919;
assign w17921 = ~w17917 & w17920;
assign w17922 = (w17921 & ~w3967) | (w17921 & w31076) | (~w3967 & w31076);
assign w17923 = (w3967 & w41117) | (w3967 & w41118) | (w41117 & w41118);
assign w17924 = (~w3967 & w41119) | (~w3967 & w41120) | (w41119 & w41120);
assign w17925 = ~w17922 & ~w17923;
assign w17926 = ~w17924 & ~w17925;
assign w17927 = ~w17916 & w17926;
assign w17928 = w17916 & ~w17926;
assign w17929 = ~w17927 & ~w17928;
assign w17930 = (w17929 & w17826) | (w17929 & w41121) | (w17826 & w41121);
assign w17931 = ~w17827 & ~w17930;
assign w17932 = w17929 & ~w17930;
assign w17933 = ~w17931 & ~w17932;
assign w17934 = ~w17825 & ~w17933;
assign w17935 = (w17825 & w17930) | (w17825 & w31077) | (w17930 & w31077);
assign w17936 = ~w17931 & w17935;
assign w17937 = ~w17934 & ~w17936;
assign w17938 = ~w17815 & w17937;
assign w17939 = ~w17937 & ~w17815;
assign w17940 = w17937 & ~w17938;
assign w17941 = (~w17814 & w17940) | (~w17814 & w31078) | (w17940 & w31078);
assign w17942 = ~w17940 & w31079;
assign w17943 = ~w17941 & ~w17942;
assign w17944 = ~w17804 & w17943;
assign w17945 = w17804 & ~w17943;
assign w17946 = ~w17944 & ~w17945;
assign w17947 = ~w17802 & w17946;
assign w17948 = w17946 & ~w17947;
assign w17949 = ~w17946 & ~w17802;
assign w17950 = ~w17948 & ~w17949;
assign w17951 = ~w17653 & ~w17657;
assign w17952 = w17950 & w17951;
assign w17953 = ~w17950 & ~w17951;
assign w17954 = ~w17952 & ~w17953;
assign w17955 = b_46 & w3803;
assign w17956 = w4027 & w31080;
assign w17957 = b_45 & w3798;
assign w17958 = ~w17956 & ~w17957;
assign w17959 = ~w17955 & w17958;
assign w17960 = (w17959 & ~w6974) | (w17959 & w31081) | (~w6974 & w31081);
assign w17961 = (w6974 & w41122) | (w6974 & w41123) | (w41122 & w41123);
assign w17962 = (~w6974 & w41124) | (~w6974 & w41125) | (w41124 & w41125);
assign w17963 = ~w17960 & ~w17961;
assign w17964 = ~w17962 & ~w17963;
assign w17965 = w17954 & ~w17964;
assign w17966 = w17954 & ~w17965;
assign w17967 = ~w17954 & ~w17964;
assign w17968 = ~w17966 & ~w17967;
assign w17969 = w17792 & ~w17968;
assign w17970 = ~w17792 & w17968;
assign w17971 = (w26384 & w27609) | (w26384 & w27610) | (w27609 & w27610);
assign w17972 = ~w17778 & ~w17971;
assign w17973 = ~w17971 & w27609;
assign w17974 = ~w17972 & ~w17973;
assign w17975 = w17765 & ~w17974;
assign w17976 = ~w17765 & w17974;
assign w17977 = w17751 & w31082;
assign w17978 = w17751 & ~w17977;
assign w17979 = (~w17976 & ~w17751) | (~w17976 & w31083) | (~w17751 & w31083);
assign w17980 = ~w17975 & w17979;
assign w17981 = ~w17978 & ~w17980;
assign w17982 = w17739 & ~w17981;
assign w17983 = ~w17739 & w17981;
assign w17984 = w17725 & w31084;
assign w17985 = w17725 & ~w17984;
assign w17986 = w31084 & ~w17725;
assign w17987 = ~w17985 & ~w17986;
assign w17988 = (w17435 & w41126) | (w17435 & w41127) | (w41126 & w41127);
assign w17989 = (~w17435 & w41128) | (~w17435 & w41129) | (w41128 & w41129);
assign w17990 = ~w17988 & ~w17989;
assign w17991 = (~w13761 & w37688) | (~w13761 & w37689) | (w37688 & w37689);
assign w17992 = (~w14835 & w31088) | (~w14835 & w31089) | (w31088 & w31089);
assign w17993 = ~w17991 & ~w17992;
assign w17994 = (~w17723 & ~w17725) | (~w17723 & w31091) | (~w17725 & w31091);
assign w17995 = (~w17738 & ~w17739) | (~w17738 & w31092) | (~w17739 & w31092);
assign w17996 = w1069 & w31093;
assign w17997 = (~w17996 & ~w12670) | (~w17996 & w31094) | (~w12670 & w31094);
assign w17998 = (w12670 & w41130) | (w12670 & w41131) | (w41130 & w41131);
assign w17999 = (~w12670 & w41132) | (~w12670 & w41133) | (w41132 & w41133);
assign w18000 = ~w17997 & ~w17998;
assign w18001 = ~w17999 & ~w18000;
assign w18002 = ~w17995 & ~w18001;
assign w18003 = ~w17995 & ~w18002;
assign w18004 = w17995 & ~w18001;
assign w18005 = b_62 & w1295;
assign w18006 = w1422 & w31095;
assign w18007 = b_61 & w1290;
assign w18008 = ~w18006 & ~w18007;
assign w18009 = ~w18005 & w18008;
assign w18010 = (w18009 & ~w12273) | (w18009 & w31096) | (~w12273 & w31096);
assign w18011 = (w12273 & w41134) | (w12273 & w41135) | (w41134 & w41135);
assign w18012 = (~w12273 & w41136) | (~w12273 & w41137) | (w41136 & w41137);
assign w18013 = ~w18010 & ~w18011;
assign w18014 = ~w18012 & ~w18013;
assign w18015 = (~w17749 & ~w17751) | (~w17749 & w31097) | (~w17751 & w31097);
assign w18016 = w18014 & w18015;
assign w18017 = ~w18014 & ~w18015;
assign w18018 = ~w18016 & ~w18017;
assign w18019 = b_59 & w1694;
assign w18020 = w1834 & w31098;
assign w18021 = b_58 & w1689;
assign w18022 = ~w18020 & ~w18021;
assign w18023 = ~w18019 & w18022;
assign w18024 = (w18023 & ~w11169) | (w18023 & w31099) | (~w11169 & w31099);
assign w18025 = (w11169 & w41138) | (w11169 & w41139) | (w41138 & w41139);
assign w18026 = (~w11169 & w41140) | (~w11169 & w41141) | (w41140 & w41141);
assign w18027 = ~w18024 & ~w18025;
assign w18028 = ~w18026 & ~w18027;
assign w18029 = (~w17764 & ~w17765) | (~w17764 & w31100) | (~w17765 & w31100);
assign w18030 = ~w18028 & ~w18029;
assign w18031 = w18029 & ~w18028;
assign w18032 = ~w18029 & ~w18030;
assign w18033 = ~w18031 & ~w18032;
assign w18034 = b_56 & w2158;
assign w18035 = w2294 & w31101;
assign w18036 = b_55 & w2153;
assign w18037 = ~w18035 & ~w18036;
assign w18038 = ~w18034 & w18037;
assign w18039 = (w18038 & ~w9798) | (w18038 & w26385) | (~w9798 & w26385);
assign w18040 = (w9798 & w31102) | (w9798 & w31103) | (w31102 & w31103);
assign w18041 = (~w9798 & w31104) | (~w9798 & w31105) | (w31104 & w31105);
assign w18042 = ~w18039 & ~w18040;
assign w18043 = ~w18041 & ~w18042;
assign w18044 = ~w17971 & w31106;
assign w18045 = (~w18043 & w17971) | (~w18043 & w31107) | (w17971 & w31107);
assign w18046 = ~w18044 & ~w18045;
assign w18047 = b_53 & w2639;
assign w18048 = w2820 & w31108;
assign w18049 = b_52 & w2634;
assign w18050 = ~w18048 & ~w18049;
assign w18051 = ~w18047 & w18050;
assign w18052 = (w9109 & w41142) | (w9109 & w41143) | (w41142 & w41143);
assign w18053 = (~w9109 & w41144) | (~w9109 & w41145) | (w41144 & w41145);
assign w18054 = (w9109 & w41146) | (w9109 & w41147) | (w41146 & w41147);
assign w18055 = ~w18052 & ~w18053;
assign w18056 = ~w18054 & ~w18055;
assign w18057 = (~w17791 & ~w17792) | (~w17791 & w27611) | (~w17792 & w27611);
assign w18058 = (~w27611 & w31111) | (~w27611 & w31112) | (w31111 & w31112);
assign w18059 = ~w18056 & ~w18058;
assign w18060 = ~w18057 & ~w18058;
assign w18061 = ~w18059 & ~w18060;
assign w18062 = b_50 & w3195;
assign w18063 = w3388 & w31113;
assign w18064 = b_49 & w3190;
assign w18065 = ~w18063 & ~w18064;
assign w18066 = ~w18062 & w18065;
assign w18067 = (w18066 & ~w8162) | (w18066 & w26388) | (~w8162 & w26388);
assign w18068 = (w8162 & w27612) | (w8162 & w27613) | (w27612 & w27613);
assign w18069 = (~w8162 & w31114) | (~w8162 & w31115) | (w31114 & w31115);
assign w18070 = ~w18067 & ~w18068;
assign w18071 = ~w18069 & ~w18070;
assign w18072 = (~w17954 & w41148) | (~w17954 & w41149) | (w41148 & w41149);
assign w18073 = (w17954 & w41150) | (w17954 & w41151) | (w41150 & w41151);
assign w18074 = ~w18072 & ~w18073;
assign w18075 = (~w17944 & ~w17946) | (~w17944 & w31117) | (~w17946 & w31117);
assign w18076 = b_44 & w4499;
assign w18077 = w4723 & w31118;
assign w18078 = b_43 & w4494;
assign w18079 = ~w18077 & ~w18078;
assign w18080 = ~w18076 & w18079;
assign w18081 = (w18080 & ~w6408) | (w18080 & w31119) | (~w6408 & w31119);
assign w18082 = (w6408 & w41152) | (w6408 & w41153) | (w41152 & w41153);
assign w18083 = (~w6408 & w41154) | (~w6408 & w41155) | (w41154 & w41155);
assign w18084 = ~w18081 & ~w18082;
assign w18085 = ~w18083 & ~w18084;
assign w18086 = ~w17938 & ~w17941;
assign w18087 = b_41 & w5196;
assign w18088 = w5459 & w31120;
assign w18089 = b_40 & w5191;
assign w18090 = ~w18088 & ~w18089;
assign w18091 = ~w18087 & w18090;
assign w18092 = (w18091 & ~w5609) | (w18091 & w31121) | (~w5609 & w31121);
assign w18093 = (w5609 & w41156) | (w5609 & w41157) | (w41156 & w41157);
assign w18094 = (~w5609 & w41158) | (~w5609 & w41159) | (w41158 & w41159);
assign w18095 = ~w18092 & ~w18093;
assign w18096 = ~w18094 & ~w18095;
assign w18097 = (~w17930 & w17933) | (~w17930 & w31122) | (w17933 & w31122);
assign w18098 = (~w17873 & ~w17874) | (~w17873 & w31123) | (~w17874 & w31123);
assign w18099 = b_26 & w9534;
assign w18100 = w9876 & w31124;
assign w18101 = b_25 & w9529;
assign w18102 = ~w18100 & ~w18101;
assign w18103 = ~w18099 & w18102;
assign w18104 = (w18103 & ~w2416) | (w18103 & w31125) | (~w2416 & w31125);
assign w18105 = (w2416 & w41160) | (w2416 & w41161) | (w41160 & w41161);
assign w18106 = (~w2416 & w41162) | (~w2416 & w41163) | (w41162 & w41163);
assign w18107 = ~w18104 & ~w18105;
assign w18108 = ~w18106 & ~w18107;
assign w18109 = (~w17854 & ~w17856) | (~w17854 & w31126) | (~w17856 & w31126);
assign w18110 = b_20 & w11620;
assign w18111 = w11969 & w31127;
assign w18112 = b_19 & w11615;
assign w18113 = ~w18111 & ~w18112;
assign w18114 = ~w18110 & w18113;
assign w18115 = (w18114 & ~w1503) | (w18114 & w31128) | (~w1503 & w31128);
assign w18116 = (w1503 & w41164) | (w1503 & w41165) | (w41164 & w41165);
assign w18117 = (~w1503 & w41166) | (~w1503 & w41167) | (w41166 & w41167);
assign w18118 = ~w18115 & ~w18116;
assign w18119 = ~w18117 & ~w18118;
assign w18120 = w12380 & w31129;
assign w18121 = b_17 & ~w12380;
assign w18122 = ~w18120 & ~w18121;
assign w18123 = w17840 & ~w18122;
assign w18124 = ~w17840 & w18122;
assign w18125 = (~w18124 & w18118) | (~w18124 & w31130) | (w18118 & w31130);
assign w18126 = ~w18123 & w18125;
assign w18127 = ~w18119 & ~w18126;
assign w18128 = (~w18124 & ~w18125) | (~w18124 & w31131) | (~w18125 & w31131);
assign w18129 = (~w31063 & w41168) | (~w31063 & w41169) | (w41168 & w41169);
assign w18130 = ~w18127 & w31134;
assign w18131 = (~w18129 & w18127) | (~w18129 & w31135) | (w18127 & w31135);
assign w18132 = ~w18130 & ~w18131;
assign w18133 = b_23 & w10562;
assign w18134 = w10902 & w31136;
assign w18135 = b_22 & w10557;
assign w18136 = ~w18134 & ~w18135;
assign w18137 = ~w18133 & w18136;
assign w18138 = (w18137 & ~w1933) | (w18137 & w31137) | (~w1933 & w31137);
assign w18139 = (w1933 & w41170) | (w1933 & w41171) | (w41170 & w41171);
assign w18140 = (~w1933 & w41172) | (~w1933 & w41173) | (w41172 & w41173);
assign w18141 = ~w18138 & ~w18139;
assign w18142 = ~w18140 & ~w18141;
assign w18143 = ~w18132 & w18142;
assign w18144 = w18132 & ~w18142;
assign w18145 = ~w18143 & ~w18144;
assign w18146 = ~w18109 & w18145;
assign w18147 = w18109 & ~w18145;
assign w18148 = ~w18146 & ~w18147;
assign w18149 = ~w18108 & w18148;
assign w18150 = w18108 & ~w18148;
assign w18151 = ~w18149 & ~w18150;
assign w18152 = ~w18098 & w18151;
assign w18153 = w18098 & ~w18151;
assign w18154 = ~w18152 & ~w18153;
assign w18155 = b_29 & w8526;
assign w18156 = w8886 & w31138;
assign w18157 = b_28 & w8521;
assign w18158 = ~w18156 & ~w18157;
assign w18159 = ~w18155 & w18158;
assign w18160 = (w18159 & ~w2954) | (w18159 & w31139) | (~w2954 & w31139);
assign w18161 = (w2954 & w41174) | (w2954 & w41175) | (w41174 & w41175);
assign w18162 = (~w2954 & w41176) | (~w2954 & w41177) | (w41176 & w41177);
assign w18163 = ~w18160 & ~w18161;
assign w18164 = ~w18162 & ~w18163;
assign w18165 = w18154 & ~w18164;
assign w18166 = w18154 & ~w18165;
assign w18167 = ~w18154 & ~w18164;
assign w18168 = ~w18166 & ~w18167;
assign w18169 = (~w17556 & w17886) | (~w17556 & w41178) | (w17886 & w41178);
assign w18170 = (~w18169 & w17891) | (~w18169 & w31140) | (w17891 & w31140);
assign w18171 = ~w18168 & ~w18170;
assign w18172 = ~w18168 & ~w18171;
assign w18173 = w18168 & ~w18170;
assign w18174 = ~w18172 & ~w18173;
assign w18175 = b_32 & w7613;
assign w18176 = w7941 & w31141;
assign w18177 = b_31 & w7608;
assign w18178 = ~w18176 & ~w18177;
assign w18179 = ~w18175 & w18178;
assign w18180 = (w18179 & ~w3545) | (w18179 & w31142) | (~w3545 & w31142);
assign w18181 = (w3545 & w41179) | (w3545 & w41180) | (w41179 & w41180);
assign w18182 = (~w3545 & w41181) | (~w3545 & w41182) | (w41181 & w41182);
assign w18183 = ~w18180 & ~w18181;
assign w18184 = ~w18182 & ~w18183;
assign w18185 = (w18184 & w18172) | (w18184 & w41183) | (w18172 & w41183);
assign w18186 = ~w18172 & w41184;
assign w18187 = ~w18185 & ~w18186;
assign w18188 = (~w17906 & ~w17908) | (~w17906 & w31143) | (~w17908 & w31143);
assign w18189 = w18187 & w18188;
assign w18190 = ~w18187 & ~w18188;
assign w18191 = ~w18189 & ~w18190;
assign w18192 = b_35 & w6761;
assign w18193 = w7075 & w31144;
assign w18194 = b_34 & w6756;
assign w18195 = ~w18193 & ~w18194;
assign w18196 = ~w18192 & w18195;
assign w18197 = (w18196 & ~w4181) | (w18196 & w31145) | (~w4181 & w31145);
assign w18198 = (w4181 & w41185) | (w4181 & w41186) | (w41185 & w41186);
assign w18199 = (~w4181 & w41187) | (~w4181 & w41188) | (w41187 & w41188);
assign w18200 = ~w18197 & ~w18198;
assign w18201 = ~w18199 & ~w18200;
assign w18202 = w18191 & ~w18201;
assign w18203 = w18191 & ~w18202;
assign w18204 = ~w18191 & ~w18201;
assign w18205 = ~w18203 & ~w18204;
assign w18206 = (~w17915 & ~w17916) | (~w17915 & w31146) | (~w17916 & w31146);
assign w18207 = ~w18205 & ~w18206;
assign w18208 = ~w18205 & ~w18207;
assign w18209 = w18205 & ~w18206;
assign w18210 = b_38 & w5962;
assign w18211 = w6246 & w31147;
assign w18212 = b_37 & w5957;
assign w18213 = ~w18211 & ~w18212;
assign w18214 = ~w18210 & w18213;
assign w18215 = (w18214 & ~w4658) | (w18214 & w31148) | (~w4658 & w31148);
assign w18216 = (w4658 & w41189) | (w4658 & w41190) | (w41189 & w41190);
assign w18217 = (~w4658 & w41191) | (~w4658 & w41192) | (w41191 & w41192);
assign w18218 = ~w18215 & ~w18216;
assign w18219 = ~w18217 & ~w18218;
assign w18220 = (w18219 & w18208) | (w18219 & w31149) | (w18208 & w31149);
assign w18221 = ~w18208 & w31150;
assign w18222 = ~w18220 & ~w18221;
assign w18223 = ~w18097 & ~w18222;
assign w18224 = w18097 & w18222;
assign w18225 = ~w18223 & ~w18224;
assign w18226 = ~w18096 & w18225;
assign w18227 = w18096 & ~w18225;
assign w18228 = ~w18226 & ~w18227;
assign w18229 = ~w18086 & w18228;
assign w18230 = w18086 & ~w18228;
assign w18231 = ~w18229 & ~w18230;
assign w18232 = ~w18085 & w18231;
assign w18233 = w18085 & ~w18231;
assign w18234 = ~w18232 & ~w18233;
assign w18235 = ~w18075 & w18234;
assign w18236 = w18075 & ~w18234;
assign w18237 = ~w18235 & ~w18236;
assign w18238 = b_47 & w3803;
assign w18239 = w4027 & w31151;
assign w18240 = b_46 & w3798;
assign w18241 = ~w18239 & ~w18240;
assign w18242 = ~w18238 & w18241;
assign w18243 = (w18242 & ~w6998) | (w18242 & w27614) | (~w6998 & w27614);
assign w18244 = (w6998 & w31152) | (w6998 & w31153) | (w31152 & w31153);
assign w18245 = (~w6998 & w31154) | (~w6998 & w31155) | (w31154 & w31155);
assign w18246 = ~w18243 & ~w18244;
assign w18247 = ~w18245 & ~w18246;
assign w18248 = w18237 & ~w18247;
assign w18249 = w18237 & ~w18248;
assign w18250 = ~w18237 & ~w18247;
assign w18251 = ~w18249 & ~w18250;
assign w18252 = w18074 & ~w18251;
assign w18253 = ~w18074 & w18251;
assign w18254 = ~w18061 & w31156;
assign w18255 = ~w18061 & ~w18254;
assign w18256 = w31156 & w18061;
assign w18257 = ~w18255 & ~w18256;
assign w18258 = w18046 & ~w18257;
assign w18259 = ~w18046 & w18257;
assign w18260 = (~w18259 & w18032) | (~w18259 & w31157) | (w18032 & w31157);
assign w18261 = ~w18258 & w18260;
assign w18262 = ~w18033 & ~w18261;
assign w18263 = (~w18260 & w31159) | (~w18260 & w31160) | (w31159 & w31160);
assign w18264 = ~w18262 & ~w18263;
assign w18265 = ~w18018 & w18264;
assign w18266 = w18018 & ~w18264;
assign w18267 = ~w18265 & ~w18266;
assign w18268 = (w18267 & w18003) | (w18267 & w31161) | (w18003 & w31161);
assign w18269 = ~w18003 & w31162;
assign w18270 = ~w18268 & ~w18269;
assign w18271 = ~w17994 & w18270;
assign w18272 = ~w17994 & ~w18271;
assign w18273 = w17994 & w18270;
assign w18274 = ~w18272 & ~w18273;
assign w18275 = (w14835 & w31163) | (w14835 & w31164) | (w31163 & w31164);
assign w18276 = (w13761 & w37690) | (w13761 & w37691) | (w37690 & w37691);
assign w18277 = ~w18275 & ~w18276;
assign w18278 = ~w18002 & ~w18268;
assign w18279 = (~w18017 & w18264) | (~w18017 & w31168) | (w18264 & w31168);
assign w18280 = b_63 & w1295;
assign w18281 = w1422 & w31169;
assign w18282 = b_62 & w1290;
assign w18283 = ~w18281 & ~w18282;
assign w18284 = ~w18280 & w18283;
assign w18285 = (w18284 & ~w12646) | (w18284 & w31170) | (~w12646 & w31170);
assign w18286 = (w12646 & w41193) | (w12646 & w41194) | (w41193 & w41194);
assign w18287 = (~w12646 & w41195) | (~w12646 & w41196) | (w41195 & w41196);
assign w18288 = ~w18285 & ~w18286;
assign w18289 = ~w18287 & ~w18288;
assign w18290 = ~w18279 & ~w18289;
assign w18291 = ~w18279 & ~w18290;
assign w18292 = w18279 & ~w18289;
assign w18293 = b_60 & w1694;
assign w18294 = w1834 & w31171;
assign w18295 = b_59 & w1689;
assign w18296 = ~w18294 & ~w18295;
assign w18297 = ~w18293 & w18296;
assign w18298 = (w18297 & ~w11196) | (w18297 & w31172) | (~w11196 & w31172);
assign w18299 = (w11196 & w41197) | (w11196 & w41198) | (w41197 & w41198);
assign w18300 = (~w11196 & w41199) | (~w11196 & w41200) | (w41199 & w41200);
assign w18301 = ~w18298 & ~w18299;
assign w18302 = ~w18300 & ~w18301;
assign w18303 = (~w18260 & w31173) | (~w18260 & w31174) | (w31173 & w31174);
assign w18304 = (w18260 & w31175) | (w18260 & w31176) | (w31175 & w31176);
assign w18305 = ~w18303 & ~w18304;
assign w18306 = b_54 & w2639;
assign w18307 = w2820 & w31177;
assign w18308 = b_53 & w2634;
assign w18309 = ~w18307 & ~w18308;
assign w18310 = ~w18306 & w18309;
assign w18311 = (w18310 & ~w9134) | (w18310 & w31178) | (~w9134 & w31178);
assign w18312 = (w9134 & w41201) | (w9134 & w41202) | (w41201 & w41202);
assign w18313 = (~w9134 & w41203) | (~w9134 & w41204) | (w41203 & w41204);
assign w18314 = ~w18311 & ~w18312;
assign w18315 = ~w18313 & ~w18314;
assign w18316 = (w18061 & w31180) | (w18061 & w31181) | (w31180 & w31181);
assign w18317 = (~w18061 & w31182) | (~w18061 & w31183) | (w31182 & w31183);
assign w18318 = ~w18316 & ~w18317;
assign w18319 = (~w18223 & ~w18225) | (~w18223 & w31184) | (~w18225 & w31184);
assign w18320 = (~w18219 & w18208) | (~w18219 & w31185) | (w18208 & w31185);
assign w18321 = ~w18207 & ~w18320;
assign w18322 = (~w18190 & ~w18191) | (~w18190 & w31186) | (~w18191 & w31186);
assign w18323 = b_27 & w9534;
assign w18324 = w9876 & w31187;
assign w18325 = b_26 & w9529;
assign w18326 = ~w18324 & ~w18325;
assign w18327 = ~w18323 & w18326;
assign w18328 = (w18327 & ~w2582) | (w18327 & w31188) | (~w2582 & w31188);
assign w18329 = (w2582 & w41205) | (w2582 & w41206) | (w41205 & w41206);
assign w18330 = (~w2582 & w41207) | (~w2582 & w41208) | (w41207 & w41208);
assign w18331 = ~w18328 & ~w18329;
assign w18332 = ~w18330 & ~w18331;
assign w18333 = (~w18131 & ~w18132) | (~w18131 & w31189) | (~w18132 & w31189);
assign w18334 = b_21 & w11620;
assign w18335 = w11969 & w31190;
assign w18336 = b_20 & w11615;
assign w18337 = ~w18335 & ~w18336;
assign w18338 = ~w18334 & w18337;
assign w18339 = (w18338 & ~w1634) | (w18338 & w31191) | (~w1634 & w31191);
assign w18340 = (w1634 & w41209) | (w1634 & w41210) | (w41209 & w41210);
assign w18341 = (~w1634 & w41211) | (~w1634 & w41212) | (w41211 & w41212);
assign w18342 = ~w18339 & ~w18340;
assign w18343 = ~w18341 & ~w18342;
assign w18344 = w12380 & w31192;
assign w18345 = b_18 & ~w12380;
assign w18346 = ~w18344 & ~w18345;
assign w18347 = ~a_17 & ~w18346;
assign w18348 = a_17 & w18346;
assign w18349 = ~w18347 & ~w18348;
assign w18350 = ~w18122 & w18349;
assign w18351 = w18122 & ~w18349;
assign w18352 = ~w18350 & ~w18351;
assign w18353 = (w18352 & w18342) | (w18352 & w31193) | (w18342 & w31193);
assign w18354 = ~w18343 & ~w18353;
assign w18355 = w18352 & ~w18353;
assign w18356 = ~w18354 & ~w18355;
assign w18357 = ~w18128 & ~w18356;
assign w18358 = w18356 & ~w18128;
assign w18359 = ~w18356 & ~w18357;
assign w18360 = b_24 & w10562;
assign w18361 = w10902 & w31194;
assign w18362 = b_23 & w10557;
assign w18363 = ~w18361 & ~w18362;
assign w18364 = ~w18360 & w18363;
assign w18365 = (w18364 & ~w2083) | (w18364 & w31195) | (~w2083 & w31195);
assign w18366 = (w2083 & w41213) | (w2083 & w41214) | (w41213 & w41214);
assign w18367 = (~w2083 & w41215) | (~w2083 & w41216) | (w41215 & w41216);
assign w18368 = ~w18365 & ~w18366;
assign w18369 = ~w18367 & ~w18368;
assign w18370 = ~w18359 & w31196;
assign w18371 = (~w18369 & w18359) | (~w18369 & w31197) | (w18359 & w31197);
assign w18372 = ~w18370 & ~w18371;
assign w18373 = ~w18333 & w18372;
assign w18374 = w18333 & ~w18372;
assign w18375 = ~w18373 & ~w18374;
assign w18376 = ~w18332 & w18375;
assign w18377 = w18375 & ~w18376;
assign w18378 = ~w18375 & ~w18332;
assign w18379 = (~w18146 & ~w18148) | (~w18146 & w31198) | (~w18148 & w31198);
assign w18380 = ~w18377 & w31199;
assign w18381 = (~w18379 & w18377) | (~w18379 & w31200) | (w18377 & w31200);
assign w18382 = ~w18380 & ~w18381;
assign w18383 = b_30 & w8526;
assign w18384 = w8886 & w31201;
assign w18385 = b_29 & w8521;
assign w18386 = ~w18384 & ~w18385;
assign w18387 = ~w18383 & w18386;
assign w18388 = (w18387 & ~w3138) | (w18387 & w31202) | (~w3138 & w31202);
assign w18389 = (w3138 & w41217) | (w3138 & w41218) | (w41217 & w41218);
assign w18390 = (~w3138 & w41219) | (~w3138 & w41220) | (w41219 & w41220);
assign w18391 = ~w18388 & ~w18389;
assign w18392 = ~w18390 & ~w18391;
assign w18393 = w18382 & ~w18392;
assign w18394 = w18382 & ~w18393;
assign w18395 = ~w18382 & ~w18392;
assign w18396 = (~w18152 & ~w18154) | (~w18152 & w31203) | (~w18154 & w31203);
assign w18397 = ~w18394 & w31204;
assign w18398 = (~w18396 & w18394) | (~w18396 & w31205) | (w18394 & w31205);
assign w18399 = ~w18397 & ~w18398;
assign w18400 = b_33 & w7613;
assign w18401 = w7941 & w31206;
assign w18402 = b_32 & w7608;
assign w18403 = ~w18401 & ~w18402;
assign w18404 = ~w18400 & w18403;
assign w18405 = (w18404 & ~w3744) | (w18404 & w31207) | (~w3744 & w31207);
assign w18406 = (w3744 & w41221) | (w3744 & w41222) | (w41221 & w41222);
assign w18407 = (~w3744 & w41223) | (~w3744 & w41224) | (w41223 & w41224);
assign w18408 = ~w18405 & ~w18406;
assign w18409 = ~w18407 & ~w18408;
assign w18410 = (~w18174 & w41225) | (~w18174 & w41226) | (w41225 & w41226);
assign w18411 = ~w18410 & w31211;
assign w18412 = (w18399 & w18410) | (w18399 & w31212) | (w18410 & w31212);
assign w18413 = ~w18411 & ~w18412;
assign w18414 = b_36 & w6761;
assign w18415 = w7075 & w31213;
assign w18416 = b_35 & w6756;
assign w18417 = ~w18415 & ~w18416;
assign w18418 = ~w18414 & w18417;
assign w18419 = (w18418 & ~w4395) | (w18418 & w31214) | (~w4395 & w31214);
assign w18420 = (w4395 & w41227) | (w4395 & w41228) | (w41227 & w41228);
assign w18421 = (~w4395 & w41229) | (~w4395 & w41230) | (w41229 & w41230);
assign w18422 = ~w18419 & ~w18420;
assign w18423 = ~w18421 & ~w18422;
assign w18424 = ~w18413 & ~w18423;
assign w18425 = w18413 & w18423;
assign w18426 = ~w18424 & ~w18425;
assign w18427 = w18322 & ~w18426;
assign w18428 = ~w18322 & w18426;
assign w18429 = ~w18427 & ~w18428;
assign w18430 = b_39 & w5962;
assign w18431 = w6246 & w31215;
assign w18432 = b_38 & w5957;
assign w18433 = ~w18431 & ~w18432;
assign w18434 = ~w18430 & w18433;
assign w18435 = (w18434 & ~w4888) | (w18434 & w31216) | (~w4888 & w31216);
assign w18436 = (w4888 & w41231) | (w4888 & w41232) | (w41231 & w41232);
assign w18437 = (~w4888 & w41233) | (~w4888 & w41234) | (w41233 & w41234);
assign w18438 = ~w18435 & ~w18436;
assign w18439 = ~w18437 & ~w18438;
assign w18440 = w18429 & ~w18439;
assign w18441 = w18429 & ~w18440;
assign w18442 = ~w18429 & ~w18439;
assign w18443 = ~w18441 & ~w18442;
assign w18444 = ~w18321 & w18443;
assign w18445 = w18321 & ~w18443;
assign w18446 = ~w18444 & ~w18445;
assign w18447 = b_42 & w5196;
assign w18448 = w5459 & w31217;
assign w18449 = b_41 & w5191;
assign w18450 = ~w18448 & ~w18449;
assign w18451 = ~w18447 & w18450;
assign w18452 = (w18451 & ~w5864) | (w18451 & w31218) | (~w5864 & w31218);
assign w18453 = (w5864 & w41235) | (w5864 & w41236) | (w41235 & w41236);
assign w18454 = (~w5864 & w41237) | (~w5864 & w41238) | (w41237 & w41238);
assign w18455 = ~w18452 & ~w18453;
assign w18456 = ~w18454 & ~w18455;
assign w18457 = ~w18446 & ~w18456;
assign w18458 = w18446 & w18456;
assign w18459 = ~w18457 & ~w18458;
assign w18460 = w18319 & ~w18459;
assign w18461 = ~w18319 & w18459;
assign w18462 = ~w18460 & ~w18461;
assign w18463 = b_45 & w4499;
assign w18464 = w4723 & w31219;
assign w18465 = b_44 & w4494;
assign w18466 = ~w18464 & ~w18465;
assign w18467 = ~w18463 & w18466;
assign w18468 = (w18467 & ~w6682) | (w18467 & w26692) | (~w6682 & w26692);
assign w18469 = (w6682 & w27615) | (w6682 & w27616) | (w27615 & w27616);
assign w18470 = (~w6682 & w31220) | (~w6682 & w31221) | (w31220 & w31221);
assign w18471 = ~w18468 & ~w18469;
assign w18472 = ~w18470 & ~w18471;
assign w18473 = w18462 & ~w18472;
assign w18474 = w18462 & ~w18473;
assign w18475 = ~w18462 & ~w18472;
assign w18476 = ~w18474 & ~w18475;
assign w18477 = (~w18229 & ~w18231) | (~w18229 & w31222) | (~w18231 & w31222);
assign w18478 = w18476 & w18477;
assign w18479 = ~w18476 & ~w18477;
assign w18480 = ~w18478 & ~w18479;
assign w18481 = b_48 & w3803;
assign w18482 = w4027 & w31223;
assign w18483 = b_47 & w3798;
assign w18484 = ~w18482 & ~w18483;
assign w18485 = ~w18481 & w18484;
assign w18486 = (w18485 & ~w7284) | (w18485 & w26693) | (~w7284 & w26693);
assign w18487 = (w7284 & w27617) | (w7284 & w27618) | (w27617 & w27618);
assign w18488 = (~w7284 & w31224) | (~w7284 & w31225) | (w31224 & w31225);
assign w18489 = ~w18486 & ~w18487;
assign w18490 = ~w18488 & ~w18489;
assign w18491 = w18480 & ~w18490;
assign w18492 = w18480 & ~w18491;
assign w18493 = ~w18480 & ~w18490;
assign w18494 = (~w18235 & ~w18237) | (~w18235 & w31226) | (~w18237 & w31226);
assign w18495 = ~w18492 & w31227;
assign w18496 = (~w18494 & w18492) | (~w18494 & w31228) | (w18492 & w31228);
assign w18497 = ~w18495 & ~w18496;
assign w18498 = b_51 & w3195;
assign w18499 = w3388 & w31229;
assign w18500 = b_50 & w3190;
assign w18501 = ~w18499 & ~w18500;
assign w18502 = ~w18498 & w18501;
assign w18503 = (w18502 & ~w8186) | (w18502 & w31230) | (~w8186 & w31230);
assign w18504 = (w8186 & w41239) | (w8186 & w41240) | (w41239 & w41240);
assign w18505 = (~w8186 & w41241) | (~w8186 & w41242) | (w41241 & w41242);
assign w18506 = ~w18503 & ~w18504;
assign w18507 = ~w18505 & ~w18506;
assign w18508 = (~w18073 & ~w18074) | (~w18073 & w31231) | (~w18074 & w31231);
assign w18509 = ~w18507 & ~w18508;
assign w18510 = w18507 & w18508;
assign w18511 = ~w18509 & ~w18510;
assign w18512 = w18497 & w18511;
assign w18513 = ~w18511 & w18497;
assign w18514 = w18511 & ~w18512;
assign w18515 = ~w18513 & ~w18514;
assign w18516 = w18318 & ~w18515;
assign w18517 = w18318 & ~w18516;
assign w18518 = ~w18318 & ~w18515;
assign w18519 = ~w18517 & ~w18518;
assign w18520 = b_57 & w2158;
assign w18521 = w2294 & w31232;
assign w18522 = b_56 & w2153;
assign w18523 = ~w18521 & ~w18522;
assign w18524 = ~w18520 & w18523;
assign w18525 = (w18524 & ~w10452) | (w18524 & w31233) | (~w10452 & w31233);
assign w18526 = (w10452 & w41243) | (w10452 & w41244) | (w41243 & w41244);
assign w18527 = (~w10452 & w41245) | (~w10452 & w41246) | (w41245 & w41246);
assign w18528 = ~w18525 & ~w18526;
assign w18529 = ~w18527 & ~w18528;
assign w18530 = (~w18045 & w18257) | (~w18045 & w41247) | (w18257 & w41247);
assign w18531 = ~w18529 & ~w18530;
assign w18532 = w18529 & w18530;
assign w18533 = ~w18531 & ~w18532;
assign w18534 = ~w18519 & w18533;
assign w18535 = ~w18533 & ~w18519;
assign w18536 = w18533 & ~w18534;
assign w18537 = ~w18535 & ~w18536;
assign w18538 = w18305 & ~w18537;
assign w18539 = w18305 & ~w18538;
assign w18540 = ~w18305 & ~w18537;
assign w18541 = ~w18539 & ~w18540;
assign w18542 = (w18541 & w18291) | (w18541 & w31234) | (w18291 & w31234);
assign w18543 = ~w18291 & w31235;
assign w18544 = ~w18542 & ~w18543;
assign w18545 = (~w18544 & w18268) | (~w18544 & w31236) | (w18268 & w31236);
assign w18546 = (~w31236 & w41248) | (~w31236 & w41249) | (w41248 & w41249);
assign w18547 = ~w31236 & w41250;
assign w18548 = ~w18546 & ~w18547;
assign w18549 = (w14835 & w31237) | (w14835 & w31238) | (w31237 & w31238);
assign w18550 = (w13761 & w37692) | (w13761 & w37693) | (w37692 & w37693);
assign w18551 = ~w18549 & ~w18550;
assign w18552 = (~w18541 & w18291) | (~w18541 & w31242) | (w18291 & w31242);
assign w18553 = ~w18290 & ~w18552;
assign w18554 = b_61 & w1694;
assign w18555 = w1834 & w31243;
assign w18556 = b_60 & w1689;
assign w18557 = ~w18555 & ~w18556;
assign w18558 = ~w18554 & w18557;
assign w18559 = (w18558 & ~w11901) | (w18558 & w31244) | (~w11901 & w31244);
assign w18560 = (w11901 & w41251) | (w11901 & w41252) | (w41251 & w41252);
assign w18561 = (~w11901 & w41253) | (~w11901 & w41254) | (w41253 & w41254);
assign w18562 = ~w18559 & ~w18560;
assign w18563 = ~w18561 & ~w18562;
assign w18564 = (~w18531 & ~w18533) | (~w18531 & w31245) | (~w18533 & w31245);
assign w18565 = w18563 & w18564;
assign w18566 = ~w18563 & ~w18564;
assign w18567 = ~w18565 & ~w18566;
assign w18568 = b_58 & w2158;
assign w18569 = w2294 & w31246;
assign w18570 = b_57 & w2153;
assign w18571 = ~w18569 & ~w18570;
assign w18572 = ~w18568 & w18571;
assign w18573 = (w18572 & ~w10476) | (w18572 & w31247) | (~w10476 & w31247);
assign w18574 = (w10476 & w41255) | (w10476 & w41256) | (w41255 & w41256);
assign w18575 = (~w10476 & w41257) | (~w10476 & w41258) | (w41257 & w41258);
assign w18576 = ~w18573 & ~w18574;
assign w18577 = ~w18575 & ~w18576;
assign w18578 = ~w18516 & w31248;
assign w18579 = (~w18577 & w18516) | (~w18577 & w31249) | (w18516 & w31249);
assign w18580 = ~w18578 & ~w18579;
assign w18581 = b_55 & w2639;
assign w18582 = w2820 & w31250;
assign w18583 = b_54 & w2634;
assign w18584 = ~w18582 & ~w18583;
assign w18585 = ~w18581 & w18584;
assign w18586 = (w18585 & ~w9776) | (w18585 & w31251) | (~w9776 & w31251);
assign w18587 = (w9776 & w41259) | (w9776 & w41260) | (w41259 & w41260);
assign w18588 = (~w9776 & w41261) | (~w9776 & w41262) | (w41261 & w41262);
assign w18589 = ~w18586 & ~w18587;
assign w18590 = ~w18588 & ~w18589;
assign w18591 = (~w18509 & ~w18511) | (~w18509 & w31252) | (~w18511 & w31252);
assign w18592 = (~w18511 & w41263) | (~w18511 & w41264) | (w41263 & w41264);
assign w18593 = (w18511 & w41265) | (w18511 & w41266) | (w41265 & w41266);
assign w18594 = ~w18592 & ~w18593;
assign w18595 = b_52 & w3195;
assign w18596 = w3388 & w31253;
assign w18597 = b_51 & w3190;
assign w18598 = ~w18596 & ~w18597;
assign w18599 = ~w18595 & w18598;
assign w18600 = (w18599 & ~w8793) | (w18599 & w26389) | (~w8793 & w26389);
assign w18601 = (w8793 & w31254) | (w8793 & w31255) | (w31254 & w31255);
assign w18602 = (~w8793 & w31256) | (~w8793 & w31257) | (w31256 & w31257);
assign w18603 = ~w18600 & ~w18601;
assign w18604 = ~w18602 & ~w18603;
assign w18605 = (~w31228 & w41267) | (~w31228 & w41268) | (w41267 & w41268);
assign w18606 = (w31228 & w41269) | (w31228 & w41270) | (w41269 & w41270);
assign w18607 = ~w18605 & ~w18606;
assign w18608 = b_43 & w5196;
assign w18609 = w5459 & w31260;
assign w18610 = b_42 & w5191;
assign w18611 = ~w18609 & ~w18610;
assign w18612 = ~w18608 & w18611;
assign w18613 = (w18612 & ~w5888) | (w18612 & w31261) | (~w5888 & w31261);
assign w18614 = (w5888 & w41271) | (w5888 & w41272) | (w41271 & w41272);
assign w18615 = (~w5888 & w41273) | (~w5888 & w41274) | (w41273 & w41274);
assign w18616 = ~w18613 & ~w18614;
assign w18617 = ~w18615 & ~w18616;
assign w18618 = ~w18321 & ~w18443;
assign w18619 = ~w18440 & ~w18618;
assign w18620 = b_40 & w5962;
assign w18621 = w6246 & w31262;
assign w18622 = b_39 & w5957;
assign w18623 = ~w18621 & ~w18622;
assign w18624 = ~w18620 & w18623;
assign w18625 = (w18624 & ~w5363) | (w18624 & w31263) | (~w5363 & w31263);
assign w18626 = (w5363 & w41275) | (w5363 & w41276) | (w41275 & w41276);
assign w18627 = (~w5363 & w41277) | (~w5363 & w41278) | (w41277 & w41278);
assign w18628 = ~w18625 & ~w18626;
assign w18629 = ~w18627 & ~w18628;
assign w18630 = (~w18424 & ~w18426) | (~w18424 & w31264) | (~w18426 & w31264);
assign w18631 = b_31 & w8526;
assign w18632 = w8886 & w31265;
assign w18633 = b_30 & w8521;
assign w18634 = ~w18632 & ~w18633;
assign w18635 = ~w18631 & w18634;
assign w18636 = (w18635 & ~w3345) | (w18635 & w31266) | (~w3345 & w31266);
assign w18637 = (w3345 & w41279) | (w3345 & w41280) | (w41279 & w41280);
assign w18638 = (~w3345 & w41281) | (~w3345 & w41282) | (w41281 & w41282);
assign w18639 = ~w18636 & ~w18637;
assign w18640 = ~w18638 & ~w18639;
assign w18641 = (~w18371 & ~w18372) | (~w18371 & w31267) | (~w18372 & w31267);
assign w18642 = b_25 & w10562;
assign w18643 = w10902 & w31268;
assign w18644 = b_24 & w10557;
assign w18645 = ~w18643 & ~w18644;
assign w18646 = ~w18642 & w18645;
assign w18647 = (w18646 & ~w2108) | (w18646 & w31269) | (~w2108 & w31269);
assign w18648 = (w2108 & w41283) | (w2108 & w41284) | (w41283 & w41284);
assign w18649 = (~w2108 & w41285) | (~w2108 & w41286) | (w41285 & w41286);
assign w18650 = ~w18647 & ~w18648;
assign w18651 = ~w18649 & ~w18650;
assign w18652 = w12380 & w31270;
assign w18653 = b_19 & ~w12380;
assign w18654 = ~w18652 & ~w18653;
assign w18655 = (~w18347 & ~w18349) | (~w18347 & w31271) | (~w18349 & w31271);
assign w18656 = ~w18654 & w18655;
assign w18657 = w18654 & ~w18655;
assign w18658 = ~w18656 & ~w18657;
assign w18659 = b_22 & w11620;
assign w18660 = w11969 & w31272;
assign w18661 = b_21 & w11615;
assign w18662 = ~w18660 & ~w18661;
assign w18663 = ~w18659 & w18662;
assign w18664 = (w18663 & ~w1786) | (w18663 & w31273) | (~w1786 & w31273);
assign w18665 = (w1786 & w41287) | (w1786 & w41288) | (w41287 & w41288);
assign w18666 = ~w18664 & ~w18665;
assign w18667 = ~w18666 & w31274;
assign w18668 = (w18658 & w18666) | (w18658 & w31275) | (w18666 & w31275);
assign w18669 = ~w18667 & ~w18668;
assign w18670 = (~w18353 & w18356) | (~w18353 & w31276) | (w18356 & w31276);
assign w18671 = w18669 & ~w18670;
assign w18672 = ~w18669 & w18670;
assign w18673 = ~w18671 & ~w18672;
assign w18674 = ~w18651 & w18673;
assign w18675 = w18673 & ~w18674;
assign w18676 = ~w18673 & ~w18651;
assign w18677 = ~w18675 & ~w18676;
assign w18678 = ~w18641 & w18677;
assign w18679 = w18641 & ~w18677;
assign w18680 = ~w18678 & ~w18679;
assign w18681 = b_28 & w9534;
assign w18682 = w9876 & w31277;
assign w18683 = b_27 & w9529;
assign w18684 = ~w18682 & ~w18683;
assign w18685 = ~w18681 & w18684;
assign w18686 = (w18685 & ~w2771) | (w18685 & w31278) | (~w2771 & w31278);
assign w18687 = (w2771 & w41289) | (w2771 & w41290) | (w41289 & w41290);
assign w18688 = (~w2771 & w41291) | (~w2771 & w41292) | (w41291 & w41292);
assign w18689 = ~w18686 & ~w18687;
assign w18690 = ~w18688 & ~w18689;
assign w18691 = w18680 & w18690;
assign w18692 = ~w18680 & ~w18690;
assign w18693 = ~w18691 & ~w18692;
assign w18694 = ~w18376 & ~w18381;
assign w18695 = w18693 & ~w18694;
assign w18696 = ~w18693 & w18694;
assign w18697 = ~w18695 & ~w18696;
assign w18698 = ~w18640 & w18697;
assign w18699 = w18697 & ~w18698;
assign w18700 = ~w18697 & ~w18640;
assign w18701 = ~w18699 & ~w18700;
assign w18702 = (~w31205 & w41293) | (~w31205 & w41294) | (w41293 & w41294);
assign w18703 = w18701 & w18702;
assign w18704 = ~w18701 & ~w18702;
assign w18705 = ~w18703 & ~w18704;
assign w18706 = b_34 & w7613;
assign w18707 = w7941 & w31279;
assign w18708 = b_33 & w7608;
assign w18709 = ~w18707 & ~w18708;
assign w18710 = ~w18706 & w18709;
assign w18711 = (w18710 & ~w3967) | (w18710 & w31280) | (~w3967 & w31280);
assign w18712 = (w3967 & w41295) | (w3967 & w41296) | (w41295 & w41296);
assign w18713 = (~w3967 & w41297) | (~w3967 & w41298) | (w41297 & w41298);
assign w18714 = ~w18711 & ~w18712;
assign w18715 = ~w18713 & ~w18714;
assign w18716 = w18705 & ~w18715;
assign w18717 = w18705 & ~w18716;
assign w18718 = ~w18705 & ~w18715;
assign w18719 = ~w18717 & ~w18718;
assign w18720 = ~w18410 & w31281;
assign w18721 = ~w18410 & ~w18720;
assign w18722 = w18719 & w18721;
assign w18723 = ~w18719 & ~w18721;
assign w18724 = ~w18722 & ~w18723;
assign w18725 = b_37 & w6761;
assign w18726 = w7075 & w31282;
assign w18727 = b_36 & w6756;
assign w18728 = ~w18726 & ~w18727;
assign w18729 = ~w18725 & w18728;
assign w18730 = (w18729 & ~w4636) | (w18729 & w31283) | (~w4636 & w31283);
assign w18731 = (w4636 & w41299) | (w4636 & w41300) | (w41299 & w41300);
assign w18732 = (~w4636 & w41301) | (~w4636 & w41302) | (w41301 & w41302);
assign w18733 = ~w18730 & ~w18731;
assign w18734 = ~w18732 & ~w18733;
assign w18735 = ~w18724 & w18734;
assign w18736 = w18724 & ~w18734;
assign w18737 = ~w18735 & ~w18736;
assign w18738 = ~w18630 & w18737;
assign w18739 = ~w18737 & ~w18630;
assign w18740 = w18737 & ~w18738;
assign w18741 = (~w18629 & w18740) | (~w18629 & w31284) | (w18740 & w31284);
assign w18742 = ~w18740 & w31285;
assign w18743 = ~w18741 & ~w18742;
assign w18744 = ~w18619 & w18743;
assign w18745 = w18619 & ~w18743;
assign w18746 = ~w18744 & ~w18745;
assign w18747 = ~w18617 & w18746;
assign w18748 = w18746 & ~w18747;
assign w18749 = ~w18746 & ~w18617;
assign w18750 = (~w18457 & ~w18459) | (~w18457 & w31286) | (~w18459 & w31286);
assign w18751 = ~w18748 & w31287;
assign w18752 = (~w18750 & w18748) | (~w18750 & w31288) | (w18748 & w31288);
assign w18753 = ~w18751 & ~w18752;
assign w18754 = b_46 & w4499;
assign w18755 = w4723 & w31289;
assign w18756 = b_45 & w4494;
assign w18757 = ~w18755 & ~w18756;
assign w18758 = ~w18754 & w18757;
assign w18759 = (w18758 & ~w6974) | (w18758 & w27619) | (~w6974 & w27619);
assign w18760 = (w6974 & w31290) | (w6974 & w31291) | (w31290 & w31291);
assign w18761 = (~w6974 & w31292) | (~w6974 & w31293) | (w31292 & w31293);
assign w18762 = ~w18759 & ~w18760;
assign w18763 = ~w18761 & ~w18762;
assign w18764 = w18753 & ~w18763;
assign w18765 = w18753 & ~w18764;
assign w18766 = ~w18753 & ~w18763;
assign w18767 = ~w18765 & ~w18766;
assign w18768 = (~w18473 & w18476) | (~w18473 & w31294) | (w18476 & w31294);
assign w18769 = w18767 & w18768;
assign w18770 = ~w18767 & ~w18768;
assign w18771 = ~w18769 & ~w18770;
assign w18772 = b_49 & w3803;
assign w18773 = w4027 & w31295;
assign w18774 = b_48 & w3798;
assign w18775 = ~w18773 & ~w18774;
assign w18776 = ~w18772 & w18775;
assign w18777 = (w18776 & ~w7859) | (w18776 & w31296) | (~w7859 & w31296);
assign w18778 = (w7859 & w41303) | (w7859 & w41304) | (w41303 & w41304);
assign w18779 = (~w7859 & w41305) | (~w7859 & w41306) | (w41305 & w41306);
assign w18780 = ~w18777 & ~w18778;
assign w18781 = ~w18779 & ~w18780;
assign w18782 = w18771 & ~w18781;
assign w18783 = w18771 & ~w18782;
assign w18784 = ~w18771 & ~w18781;
assign w18785 = ~w18783 & ~w18784;
assign w18786 = w18607 & ~w18785;
assign w18787 = ~w18607 & w18785;
assign w18788 = w18594 & w31297;
assign w18789 = w18594 & ~w18788;
assign w18790 = w31297 & ~w18594;
assign w18791 = ~w18789 & ~w18790;
assign w18792 = w18580 & ~w18791;
assign w18793 = ~w18580 & w18791;
assign w18794 = w18567 & w31298;
assign w18795 = w18567 & ~w18794;
assign w18796 = w31298 & ~w18567;
assign w18797 = ~w18795 & ~w18796;
assign w18798 = (~w18304 & ~w18305) | (~w18304 & w31299) | (~w18305 & w31299);
assign w18799 = w1422 & w31300;
assign w18800 = b_63 & w1290;
assign w18801 = ~w18799 & ~w18800;
assign w18802 = ~w12671 & w31301;
assign w18803 = (a_20 & w18802) | (a_20 & w31302) | (w18802 & w31302);
assign w18804 = ~w18802 & w31303;
assign w18805 = ~w18803 & ~w18804;
assign w18806 = ~w18798 & ~w18805;
assign w18807 = ~w18798 & ~w18806;
assign w18808 = w18798 & ~w18805;
assign w18809 = (~w18797 & w18807) | (~w18797 & w31304) | (w18807 & w31304);
assign w18810 = w18797 & ~w18808;
assign w18811 = ~w18807 & w18810;
assign w18812 = ~w18809 & ~w18811;
assign w18813 = ~w18553 & w18812;
assign w18814 = ~w18553 & ~w18813;
assign w18815 = w18553 & w18812;
assign w18816 = ~w18814 & ~w18815;
assign w18817 = (w14835 & w31305) | (w14835 & w31306) | (w31305 & w31306);
assign w18818 = (w13761 & w37694) | (w13761 & w37695) | (w37694 & w37695);
assign w18819 = ~w18817 & ~w18818;
assign w18820 = ~w18806 & ~w18809;
assign w18821 = (~w18566 & ~w18567) | (~w18566 & w31311) | (~w18567 & w31311);
assign w18822 = w1422 & w31312;
assign w18823 = (~w18822 & ~w12670) | (~w18822 & w31313) | (~w12670 & w31313);
assign w18824 = (w12670 & w41307) | (w12670 & w41308) | (w41307 & w41308);
assign w18825 = (~w12670 & w41309) | (~w12670 & w41310) | (w41309 & w41310);
assign w18826 = ~w18823 & ~w18824;
assign w18827 = ~w18825 & ~w18826;
assign w18828 = ~w18821 & ~w18827;
assign w18829 = ~w18821 & ~w18828;
assign w18830 = w18821 & ~w18827;
assign w18831 = b_62 & w1694;
assign w18832 = w1834 & w31314;
assign w18833 = b_61 & w1689;
assign w18834 = ~w18832 & ~w18833;
assign w18835 = ~w18831 & w18834;
assign w18836 = (w18835 & ~w12273) | (w18835 & w31315) | (~w12273 & w31315);
assign w18837 = (w12273 & w41311) | (w12273 & w41312) | (w41311 & w41312);
assign w18838 = (~w12273 & w41313) | (~w12273 & w41314) | (w41313 & w41314);
assign w18839 = ~w18836 & ~w18837;
assign w18840 = ~w18838 & ~w18839;
assign w18841 = (~w18579 & ~w18580) | (~w18579 & w41315) | (~w18580 & w41315);
assign w18842 = (w18580 & w41316) | (w18580 & w41317) | (w41316 & w41317);
assign w18843 = ~w18792 & w31317;
assign w18844 = ~w18841 & ~w18842;
assign w18845 = ~w18843 & ~w18844;
assign w18846 = b_59 & w2158;
assign w18847 = w2294 & w31318;
assign w18848 = b_58 & w2153;
assign w18849 = ~w18847 & ~w18848;
assign w18850 = ~w18846 & w18849;
assign w18851 = (w18850 & ~w11169) | (w18850 & w31319) | (~w11169 & w31319);
assign w18852 = (w11169 & w41318) | (w11169 & w41319) | (w41318 & w41319);
assign w18853 = (~w11169 & w41320) | (~w11169 & w41321) | (w41320 & w41321);
assign w18854 = ~w18851 & ~w18852;
assign w18855 = ~w18853 & ~w18854;
assign w18856 = (~w18593 & ~w18594) | (~w18593 & w31320) | (~w18594 & w31320);
assign w18857 = w18855 & w18856;
assign w18858 = ~w18855 & ~w18856;
assign w18859 = ~w18857 & ~w18858;
assign w18860 = b_56 & w2639;
assign w18861 = w2820 & w31321;
assign w18862 = b_55 & w2634;
assign w18863 = ~w18861 & ~w18862;
assign w18864 = ~w18860 & w18863;
assign w18865 = (w18864 & ~w9798) | (w18864 & w26003) | (~w9798 & w26003);
assign w18866 = (w9798 & w26390) | (w9798 & w26391) | (w26390 & w26391);
assign w18867 = (~w9798 & w31322) | (~w9798 & w31323) | (w31322 & w31323);
assign w18868 = ~w18865 & ~w18866;
assign w18869 = ~w18867 & ~w18868;
assign w18870 = (~w18606 & w18785) | (~w18606 & w41322) | (w18785 & w41322);
assign w18871 = (~w18785 & w41323) | (~w18785 & w41324) | (w41323 & w41324);
assign w18872 = (w31325 & w18785) | (w31325 & w41325) | (w18785 & w41325);
assign w18873 = ~w18870 & ~w18871;
assign w18874 = ~w18872 & ~w18873;
assign w18875 = b_53 & w3195;
assign w18876 = w3388 & w31326;
assign w18877 = b_52 & w3190;
assign w18878 = ~w18876 & ~w18877;
assign w18879 = ~w18875 & w18878;
assign w18880 = (w9109 & w41326) | (w9109 & w41327) | (w41326 & w41327);
assign w18881 = (~w9109 & w41328) | (~w9109 & w41329) | (w41328 & w41329);
assign w18882 = (w9109 & w41330) | (w9109 & w41331) | (w41330 & w41331);
assign w18883 = ~w18880 & ~w18881;
assign w18884 = ~w18882 & ~w18883;
assign w18885 = (~w18771 & w41332) | (~w18771 & w41333) | (w41332 & w41333);
assign w18886 = (w18771 & w41334) | (w18771 & w41335) | (w41334 & w41335);
assign w18887 = ~w18885 & ~w18886;
assign w18888 = (~w18744 & ~w18746) | (~w18744 & w31332) | (~w18746 & w31332);
assign w18889 = b_44 & w5196;
assign w18890 = w5459 & w31333;
assign w18891 = b_43 & w5191;
assign w18892 = ~w18890 & ~w18891;
assign w18893 = ~w18889 & w18892;
assign w18894 = (w18893 & ~w6408) | (w18893 & w31334) | (~w6408 & w31334);
assign w18895 = (w6408 & w41336) | (w6408 & w41337) | (w41336 & w41337);
assign w18896 = (~w6408 & w41338) | (~w6408 & w41339) | (w41338 & w41339);
assign w18897 = ~w18894 & ~w18895;
assign w18898 = ~w18896 & ~w18897;
assign w18899 = ~w18738 & ~w18741;
assign w18900 = b_41 & w5962;
assign w18901 = w6246 & w31335;
assign w18902 = b_40 & w5957;
assign w18903 = ~w18901 & ~w18902;
assign w18904 = ~w18900 & w18903;
assign w18905 = (w18904 & ~w5609) | (w18904 & w31336) | (~w5609 & w31336);
assign w18906 = (w5609 & w41340) | (w5609 & w41341) | (w41340 & w41341);
assign w18907 = (~w5609 & w41342) | (~w5609 & w41343) | (w41342 & w41343);
assign w18908 = ~w18905 & ~w18906;
assign w18909 = ~w18907 & ~w18908;
assign w18910 = (~w18723 & ~w18724) | (~w18723 & w31337) | (~w18724 & w31337);
assign w18911 = b_38 & w6761;
assign w18912 = w7075 & w31338;
assign w18913 = b_37 & w6756;
assign w18914 = ~w18912 & ~w18913;
assign w18915 = ~w18911 & w18914;
assign w18916 = (w18915 & ~w4658) | (w18915 & w31339) | (~w4658 & w31339);
assign w18917 = (w4658 & w41344) | (w4658 & w41345) | (w41344 & w41345);
assign w18918 = (~w4658 & w41346) | (~w4658 & w41347) | (w41346 & w41347);
assign w18919 = ~w18916 & ~w18917;
assign w18920 = ~w18918 & ~w18919;
assign w18921 = (~w18704 & ~w18705) | (~w18704 & w31340) | (~w18705 & w31340);
assign w18922 = b_35 & w7613;
assign w18923 = w7941 & w31341;
assign w18924 = b_34 & w7608;
assign w18925 = ~w18923 & ~w18924;
assign w18926 = ~w18922 & w18925;
assign w18927 = (w18926 & ~w4181) | (w18926 & w31342) | (~w4181 & w31342);
assign w18928 = (w4181 & w41348) | (w4181 & w41349) | (w41348 & w41349);
assign w18929 = (~w4181 & w41350) | (~w4181 & w41351) | (w41350 & w41351);
assign w18930 = ~w18927 & ~w18928;
assign w18931 = ~w18929 & ~w18930;
assign w18932 = (~w18695 & ~w18697) | (~w18695 & w31343) | (~w18697 & w31343);
assign w18933 = (~w18671 & ~w18673) | (~w18671 & w31344) | (~w18673 & w31344);
assign w18934 = b_26 & w10562;
assign w18935 = w10902 & w31345;
assign w18936 = b_25 & w10557;
assign w18937 = ~w18935 & ~w18936;
assign w18938 = ~w18934 & w18937;
assign w18939 = (w18938 & ~w2416) | (w18938 & w31346) | (~w2416 & w31346);
assign w18940 = (w2416 & w41352) | (w2416 & w41353) | (w41352 & w41353);
assign w18941 = (~w2416 & w41354) | (~w2416 & w41355) | (w41354 & w41355);
assign w18942 = ~w18939 & ~w18940;
assign w18943 = ~w18941 & ~w18942;
assign w18944 = ~w18657 & ~w18668;
assign w18945 = w12380 & w31347;
assign w18946 = b_20 & ~w12380;
assign w18947 = ~w18945 & ~w18946;
assign w18948 = ~w18654 & w18947;
assign w18949 = w18654 & ~w18947;
assign w18950 = ~w18948 & ~w18949;
assign w18951 = b_23 & w11620;
assign w18952 = w11969 & w31348;
assign w18953 = b_22 & w11615;
assign w18954 = ~w18952 & ~w18953;
assign w18955 = ~w18951 & w18954;
assign w18956 = w18954 & w31349;
assign w18957 = (~w1933 & w41356) | (~w1933 & w41357) | (w41356 & w41357);
assign w18958 = (w18950 & w18957) | (w18950 & w31352) | (w18957 & w31352);
assign w18959 = ~w18957 & w31353;
assign w18960 = ~w18958 & ~w18959;
assign w18961 = ~w18944 & w18960;
assign w18962 = w18944 & ~w18960;
assign w18963 = ~w18961 & ~w18962;
assign w18964 = ~w18943 & w18963;
assign w18965 = w18943 & ~w18963;
assign w18966 = ~w18964 & ~w18965;
assign w18967 = ~w18933 & w18966;
assign w18968 = w18933 & ~w18966;
assign w18969 = ~w18967 & ~w18968;
assign w18970 = b_29 & w9534;
assign w18971 = w9876 & w31354;
assign w18972 = b_28 & w9529;
assign w18973 = ~w18971 & ~w18972;
assign w18974 = ~w18970 & w18973;
assign w18975 = (w18974 & ~w2954) | (w18974 & w31355) | (~w2954 & w31355);
assign w18976 = (w2954 & w41358) | (w2954 & w41359) | (w41358 & w41359);
assign w18977 = (~w2954 & w41360) | (~w2954 & w41361) | (w41360 & w41361);
assign w18978 = ~w18975 & ~w18976;
assign w18979 = ~w18977 & ~w18978;
assign w18980 = w18969 & ~w18979;
assign w18981 = w18969 & ~w18980;
assign w18982 = ~w18969 & ~w18979;
assign w18983 = ~w18981 & ~w18982;
assign w18984 = ~w18641 & ~w18677;
assign w18985 = (~w18984 & w18680) | (~w18984 & w31356) | (w18680 & w31356);
assign w18986 = ~w18983 & ~w18985;
assign w18987 = ~w18983 & ~w18986;
assign w18988 = ~w18985 & ~w18986;
assign w18989 = ~w18987 & ~w18988;
assign w18990 = b_32 & w8526;
assign w18991 = w8886 & w31357;
assign w18992 = b_31 & w8521;
assign w18993 = ~w18991 & ~w18992;
assign w18994 = ~w18990 & w18993;
assign w18995 = (w18994 & ~w3545) | (w18994 & w31358) | (~w3545 & w31358);
assign w18996 = (w3545 & w41362) | (w3545 & w41363) | (w41362 & w41363);
assign w18997 = (~w3545 & w41364) | (~w3545 & w41365) | (w41364 & w41365);
assign w18998 = ~w18995 & ~w18996;
assign w18999 = ~w18997 & ~w18998;
assign w19000 = ~w18989 & w18999;
assign w19001 = w18989 & ~w18999;
assign w19002 = ~w19000 & ~w19001;
assign w19003 = ~w18932 & ~w19002;
assign w19004 = w18932 & w19002;
assign w19005 = ~w19003 & ~w19004;
assign w19006 = ~w18931 & w19005;
assign w19007 = w18931 & ~w19005;
assign w19008 = ~w19006 & ~w19007;
assign w19009 = ~w18921 & w19008;
assign w19010 = w18921 & ~w19008;
assign w19011 = ~w19009 & ~w19010;
assign w19012 = ~w18920 & w19011;
assign w19013 = w18920 & ~w19011;
assign w19014 = ~w19012 & ~w19013;
assign w19015 = ~w18910 & w19014;
assign w19016 = w18910 & ~w19014;
assign w19017 = ~w19015 & ~w19016;
assign w19018 = ~w18909 & w19017;
assign w19019 = w18909 & ~w19017;
assign w19020 = ~w19018 & ~w19019;
assign w19021 = ~w18899 & w19020;
assign w19022 = w18899 & ~w19020;
assign w19023 = ~w19021 & ~w19022;
assign w19024 = ~w18898 & w19023;
assign w19025 = w18898 & ~w19023;
assign w19026 = ~w19024 & ~w19025;
assign w19027 = ~w18888 & w19026;
assign w19028 = w18888 & ~w19026;
assign w19029 = ~w19027 & ~w19028;
assign w19030 = b_47 & w4499;
assign w19031 = w4723 & w31359;
assign w19032 = b_46 & w4494;
assign w19033 = ~w19031 & ~w19032;
assign w19034 = ~w19030 & w19033;
assign w19035 = (w19034 & ~w6998) | (w19034 & w27620) | (~w6998 & w27620);
assign w19036 = (w6998 & w31360) | (w6998 & w31361) | (w31360 & w31361);
assign w19037 = (~w6998 & w31362) | (~w6998 & w31363) | (w31362 & w31363);
assign w19038 = ~w19035 & ~w19036;
assign w19039 = ~w19037 & ~w19038;
assign w19040 = w19029 & ~w19039;
assign w19041 = w19029 & ~w19040;
assign w19042 = ~w19029 & ~w19039;
assign w19043 = ~w19041 & ~w19042;
assign w19044 = (~w18752 & ~w18753) | (~w18752 & w31364) | (~w18753 & w31364);
assign w19045 = w19043 & w19044;
assign w19046 = ~w19043 & ~w19044;
assign w19047 = ~w19045 & ~w19046;
assign w19048 = b_50 & w3803;
assign w19049 = w4027 & w31365;
assign w19050 = b_49 & w3798;
assign w19051 = ~w19049 & ~w19050;
assign w19052 = ~w19048 & w19051;
assign w19053 = (w19052 & ~w8162) | (w19052 & w31366) | (~w8162 & w31366);
assign w19054 = (w8162 & w41366) | (w8162 & w41367) | (w41366 & w41367);
assign w19055 = (~w8162 & w41368) | (~w8162 & w41369) | (w41368 & w41369);
assign w19056 = ~w19053 & ~w19054;
assign w19057 = ~w19055 & ~w19056;
assign w19058 = w19047 & ~w19057;
assign w19059 = ~w19047 & w19057;
assign w19060 = w18887 & w31367;
assign w19061 = w18887 & ~w19060;
assign w19062 = w31367 & ~w18887;
assign w19063 = ~w19061 & ~w19062;
assign w19064 = ~w18874 & w19063;
assign w19065 = w18874 & ~w19063;
assign w19066 = ~w19064 & ~w19065;
assign w19067 = w18859 & ~w19066;
assign w19068 = w18859 & ~w19067;
assign w19069 = ~w18859 & ~w19066;
assign w19070 = ~w19068 & ~w19069;
assign w19071 = ~w18845 & w19070;
assign w19072 = w18845 & ~w19070;
assign w19073 = ~w19071 & ~w19072;
assign w19074 = (~w19073 & w18829) | (~w19073 & w31368) | (w18829 & w31368);
assign w19075 = ~w18829 & w31369;
assign w19076 = ~w19074 & ~w19075;
assign w19077 = ~w18820 & w19076;
assign w19078 = w18820 & ~w19076;
assign w19079 = ~w19077 & ~w19078;
assign w19080 = (w14835 & w31370) | (w14835 & w31371) | (w31370 & w31371);
assign w19081 = (w13761 & w37696) | (w13761 & w37697) | (w37696 & w37697);
assign w19082 = ~w19080 & ~w19081;
assign w19083 = (~w18842 & w18845) | (~w18842 & w31372) | (w18845 & w31372);
assign w19084 = b_63 & w1694;
assign w19085 = w1834 & w31373;
assign w19086 = b_62 & w1689;
assign w19087 = ~w19085 & ~w19086;
assign w19088 = ~w19084 & w19087;
assign w19089 = (w19088 & ~w12646) | (w19088 & w31374) | (~w12646 & w31374);
assign w19090 = (w12646 & w41370) | (w12646 & w41371) | (w41370 & w41371);
assign w19091 = (~w12646 & w41372) | (~w12646 & w41373) | (w41372 & w41373);
assign w19092 = ~w19089 & ~w19090;
assign w19093 = ~w19091 & ~w19092;
assign w19094 = (~w18845 & w41374) | (~w18845 & w41375) | (w41374 & w41375);
assign w19095 = ~w19083 & ~w19094;
assign w19096 = (w18845 & w41376) | (w18845 & w41377) | (w41376 & w41377);
assign w19097 = ~w19095 & ~w19096;
assign w19098 = b_60 & w2158;
assign w19099 = w2294 & w31375;
assign w19100 = b_59 & w2153;
assign w19101 = ~w19099 & ~w19100;
assign w19102 = ~w19098 & w19101;
assign w19103 = (w19102 & ~w11196) | (w19102 & w31376) | (~w11196 & w31376);
assign w19104 = (w11196 & w41378) | (w11196 & w41379) | (w41378 & w41379);
assign w19105 = (~w11196 & w41380) | (~w11196 & w41381) | (w41380 & w41381);
assign w19106 = ~w19103 & ~w19104;
assign w19107 = ~w19105 & ~w19106;
assign w19108 = (~w18858 & ~w18859) | (~w18858 & w31377) | (~w18859 & w31377);
assign w19109 = w19107 & w19108;
assign w19110 = ~w19107 & ~w19108;
assign w19111 = ~w19109 & ~w19110;
assign w19112 = (~w18871 & w18874) | (~w18871 & w31378) | (w18874 & w31378);
assign w19113 = b_57 & w2639;
assign w19114 = w2820 & w31379;
assign w19115 = b_56 & w2634;
assign w19116 = ~w19114 & ~w19115;
assign w19117 = ~w19113 & w19116;
assign w19118 = (w19117 & ~w10452) | (w19117 & w31380) | (~w10452 & w31380);
assign w19119 = (w10452 & w41382) | (w10452 & w41383) | (w41382 & w41383);
assign w19120 = (~w10452 & w41384) | (~w10452 & w41385) | (w41384 & w41385);
assign w19121 = ~w19118 & ~w19119;
assign w19122 = ~w19120 & ~w19121;
assign w19123 = ~w19112 & w19122;
assign w19124 = w19112 & ~w19122;
assign w19125 = ~w19123 & ~w19124;
assign w19126 = b_54 & w3195;
assign w19127 = w3388 & w31381;
assign w19128 = b_53 & w3190;
assign w19129 = ~w19127 & ~w19128;
assign w19130 = ~w19126 & w19129;
assign w19131 = (w19130 & ~w9134) | (w19130 & w31382) | (~w9134 & w31382);
assign w19132 = (w9134 & w41386) | (w9134 & w41387) | (w41386 & w41387);
assign w19133 = (~w9134 & w41388) | (~w9134 & w41389) | (w41388 & w41389);
assign w19134 = ~w19131 & ~w19132;
assign w19135 = ~w19133 & ~w19134;
assign w19136 = (~w18886 & ~w18887) | (~w18886 & w31383) | (~w18887 & w31383);
assign w19137 = w19135 & w19136;
assign w19138 = ~w19135 & ~w19136;
assign w19139 = ~w19137 & ~w19138;
assign w19140 = (~w19046 & ~w19047) | (~w19046 & w31384) | (~w19047 & w31384);
assign w19141 = (~w19003 & ~w19005) | (~w19003 & w31385) | (~w19005 & w31385);
assign w19142 = w12380 & w31386;
assign w19143 = b_21 & ~w12380;
assign w19144 = ~w19142 & ~w19143;
assign w19145 = ~a_20 & ~w19144;
assign w19146 = a_20 & w19144;
assign w19147 = ~w19145 & ~w19146;
assign w19148 = ~w18947 & w19147;
assign w19149 = w18947 & ~w19147;
assign w19150 = ~w19148 & ~w19149;
assign w19151 = b_24 & w11620;
assign w19152 = w11969 & w31387;
assign w19153 = b_23 & w11615;
assign w19154 = ~w19152 & ~w19153;
assign w19155 = ~w19151 & w19154;
assign w19156 = (w19155 & ~w2083) | (w19155 & w31388) | (~w2083 & w31388);
assign w19157 = (w2083 & w41390) | (w2083 & w41391) | (w41390 & w41391);
assign w19158 = (~w2083 & w41392) | (~w2083 & w41393) | (w41392 & w41393);
assign w19159 = ~w19156 & ~w19157;
assign w19160 = ~w19158 & ~w19159;
assign w19161 = (w19150 & w19159) | (w19150 & w31389) | (w19159 & w31389);
assign w19162 = w19150 & ~w19161;
assign w19163 = ~w19160 & ~w19161;
assign w19164 = ~w19162 & ~w19163;
assign w19165 = ~w18948 & ~w18958;
assign w19166 = ~w19164 & ~w19165;
assign w19167 = ~w19164 & ~w19166;
assign w19168 = w19164 & ~w19165;
assign w19169 = ~w19167 & ~w19168;
assign w19170 = b_27 & w10562;
assign w19171 = w10902 & w31390;
assign w19172 = b_26 & w10557;
assign w19173 = ~w19171 & ~w19172;
assign w19174 = ~w19170 & w19173;
assign w19175 = (w19174 & ~w2582) | (w19174 & w31391) | (~w2582 & w31391);
assign w19176 = (w2582 & w41394) | (w2582 & w41395) | (w41394 & w41395);
assign w19177 = (~w2582 & w41396) | (~w2582 & w41397) | (w41396 & w41397);
assign w19178 = ~w19175 & ~w19176;
assign w19179 = ~w19177 & ~w19178;
assign w19180 = (~w19179 & w19167) | (~w19179 & w31392) | (w19167 & w31392);
assign w19181 = ~w19169 & ~w19180;
assign w19182 = ~w19167 & w41398;
assign w19183 = ~w19181 & ~w19182;
assign w19184 = (~w18961 & ~w18963) | (~w18961 & w31393) | (~w18963 & w31393);
assign w19185 = ~w19181 & w41399;
assign w19186 = (~w19184 & w19181) | (~w19184 & w41400) | (w19181 & w41400);
assign w19187 = ~w19185 & ~w19186;
assign w19188 = b_30 & w9534;
assign w19189 = w9876 & w31394;
assign w19190 = b_29 & w9529;
assign w19191 = ~w19189 & ~w19190;
assign w19192 = ~w19188 & w19191;
assign w19193 = (w19192 & ~w3138) | (w19192 & w31395) | (~w3138 & w31395);
assign w19194 = (w3138 & w41401) | (w3138 & w41402) | (w41401 & w41402);
assign w19195 = (~w3138 & w41403) | (~w3138 & w41404) | (w41403 & w41404);
assign w19196 = ~w19193 & ~w19194;
assign w19197 = ~w19195 & ~w19196;
assign w19198 = w19187 & ~w19197;
assign w19199 = w19187 & ~w19198;
assign w19200 = (~w18967 & ~w18969) | (~w18967 & w31396) | (~w18969 & w31396);
assign w19201 = ~w19199 & w31397;
assign w19202 = (~w19200 & w19199) | (~w19200 & w31398) | (w19199 & w31398);
assign w19203 = ~w19201 & ~w19202;
assign w19204 = b_33 & w8526;
assign w19205 = w8886 & w31399;
assign w19206 = b_32 & w8521;
assign w19207 = ~w19205 & ~w19206;
assign w19208 = ~w19204 & w19207;
assign w19209 = (w19208 & ~w3744) | (w19208 & w31400) | (~w3744 & w31400);
assign w19210 = (w3744 & w41405) | (w3744 & w41406) | (w41405 & w41406);
assign w19211 = (~w3744 & w41407) | (~w3744 & w41408) | (w41407 & w41408);
assign w19212 = ~w19209 & ~w19210;
assign w19213 = ~w19211 & ~w19212;
assign w19214 = (~w18986 & w18989) | (~w18986 & w31401) | (w18989 & w31401);
assign w19215 = (~w18989 & w41409) | (~w18989 & w41410) | (w41409 & w41410);
assign w19216 = (w18989 & w31402) | (w18989 & w31403) | (w31402 & w31403);
assign w19217 = ~w19215 & w31404;
assign w19218 = (w19203 & w19215) | (w19203 & w31405) | (w19215 & w31405);
assign w19219 = ~w19217 & ~w19218;
assign w19220 = b_36 & w7613;
assign w19221 = w7941 & w31406;
assign w19222 = b_35 & w7608;
assign w19223 = ~w19221 & ~w19222;
assign w19224 = ~w19220 & w19223;
assign w19225 = (w19224 & ~w4395) | (w19224 & w31407) | (~w4395 & w31407);
assign w19226 = (w4395 & w41411) | (w4395 & w41412) | (w41411 & w41412);
assign w19227 = (~w4395 & w41413) | (~w4395 & w41414) | (w41413 & w41414);
assign w19228 = ~w19225 & ~w19226;
assign w19229 = ~w19227 & ~w19228;
assign w19230 = ~w19219 & ~w19229;
assign w19231 = w19219 & w19229;
assign w19232 = ~w19230 & ~w19231;
assign w19233 = w19141 & ~w19232;
assign w19234 = ~w19141 & w19232;
assign w19235 = ~w19233 & ~w19234;
assign w19236 = b_39 & w6761;
assign w19237 = w7075 & w31408;
assign w19238 = b_38 & w6756;
assign w19239 = ~w19237 & ~w19238;
assign w19240 = ~w19236 & w19239;
assign w19241 = (w19240 & ~w4888) | (w19240 & w31409) | (~w4888 & w31409);
assign w19242 = (w4888 & w41415) | (w4888 & w41416) | (w41415 & w41416);
assign w19243 = (~w4888 & w41417) | (~w4888 & w41418) | (w41417 & w41418);
assign w19244 = ~w19241 & ~w19242;
assign w19245 = ~w19243 & ~w19244;
assign w19246 = w19235 & ~w19245;
assign w19247 = w19235 & ~w19246;
assign w19248 = ~w19235 & ~w19245;
assign w19249 = (~w19009 & ~w19011) | (~w19009 & w31410) | (~w19011 & w31410);
assign w19250 = ~w19247 & w31411;
assign w19251 = (~w19249 & w19247) | (~w19249 & w31412) | (w19247 & w31412);
assign w19252 = ~w19250 & ~w19251;
assign w19253 = b_42 & w5962;
assign w19254 = w6246 & w31413;
assign w19255 = b_41 & w5957;
assign w19256 = ~w19254 & ~w19255;
assign w19257 = ~w19253 & w19256;
assign w19258 = (w19257 & ~w5864) | (w19257 & w31414) | (~w5864 & w31414);
assign w19259 = (w5864 & w41419) | (w5864 & w41420) | (w41419 & w41420);
assign w19260 = (~w5864 & w41421) | (~w5864 & w41422) | (w41421 & w41422);
assign w19261 = ~w19258 & ~w19259;
assign w19262 = ~w19260 & ~w19261;
assign w19263 = w19252 & ~w19262;
assign w19264 = w19252 & ~w19263;
assign w19265 = ~w19252 & ~w19262;
assign w19266 = ~w19264 & ~w19265;
assign w19267 = (~w19015 & ~w19017) | (~w19015 & w31415) | (~w19017 & w31415);
assign w19268 = w19266 & w19267;
assign w19269 = ~w19266 & ~w19267;
assign w19270 = ~w19268 & ~w19269;
assign w19271 = b_45 & w5196;
assign w19272 = w5459 & w31416;
assign w19273 = b_44 & w5191;
assign w19274 = ~w19272 & ~w19273;
assign w19275 = ~w19271 & w19274;
assign w19276 = (w19275 & ~w6682) | (w19275 & w27621) | (~w6682 & w27621);
assign w19277 = (w6682 & w31417) | (w6682 & w31418) | (w31417 & w31418);
assign w19278 = (~w6682 & w31419) | (~w6682 & w31420) | (w31419 & w31420);
assign w19279 = ~w19276 & ~w19277;
assign w19280 = ~w19278 & ~w19279;
assign w19281 = w19270 & ~w19280;
assign w19282 = w19270 & ~w19281;
assign w19283 = ~w19270 & ~w19280;
assign w19284 = ~w19282 & ~w19283;
assign w19285 = (~w19021 & ~w19023) | (~w19021 & w31421) | (~w19023 & w31421);
assign w19286 = w19284 & w19285;
assign w19287 = ~w19284 & ~w19285;
assign w19288 = ~w19286 & ~w19287;
assign w19289 = b_48 & w4499;
assign w19290 = w4723 & w31422;
assign w19291 = b_47 & w4494;
assign w19292 = ~w19290 & ~w19291;
assign w19293 = ~w19289 & w19292;
assign w19294 = (w19293 & ~w7284) | (w19293 & w27622) | (~w7284 & w27622);
assign w19295 = (w7284 & w31423) | (w7284 & w31424) | (w31423 & w31424);
assign w19296 = (~w7284 & w31425) | (~w7284 & w31426) | (w31425 & w31426);
assign w19297 = ~w19294 & ~w19295;
assign w19298 = ~w19296 & ~w19297;
assign w19299 = w19288 & ~w19298;
assign w19300 = w19288 & ~w19299;
assign w19301 = ~w19288 & ~w19298;
assign w19302 = (~w19027 & ~w19029) | (~w19027 & w31427) | (~w19029 & w31427);
assign w19303 = ~w19300 & w31428;
assign w19304 = (~w19302 & w19300) | (~w19302 & w31429) | (w19300 & w31429);
assign w19305 = ~w19303 & ~w19304;
assign w19306 = b_51 & w3803;
assign w19307 = w4027 & w31430;
assign w19308 = b_50 & w3798;
assign w19309 = ~w19307 & ~w19308;
assign w19310 = ~w19306 & w19309;
assign w19311 = (w19310 & ~w8186) | (w19310 & w31431) | (~w8186 & w31431);
assign w19312 = (w8186 & w41423) | (w8186 & w41424) | (w41423 & w41424);
assign w19313 = (~w8186 & w41425) | (~w8186 & w41426) | (w41425 & w41426);
assign w19314 = ~w19311 & ~w19312;
assign w19315 = ~w19313 & ~w19314;
assign w19316 = w19305 & ~w19315;
assign w19317 = ~w19305 & w19315;
assign w19318 = ~w19140 & w31432;
assign w19319 = ~w19140 & ~w19318;
assign w19320 = ~w19318 & w31432;
assign w19321 = ~w19319 & ~w19320;
assign w19322 = w19139 & ~w19321;
assign w19323 = ~w19139 & w19321;
assign w19324 = ~w19125 & w31433;
assign w19325 = ~w19125 & ~w19324;
assign w19326 = w31433 & w19125;
assign w19327 = ~w19325 & ~w19326;
assign w19328 = w19111 & ~w19327;
assign w19329 = ~w19111 & w19327;
assign w19330 = (~w19329 & w19095) | (~w19329 & w31434) | (w19095 & w31434);
assign w19331 = ~w19328 & w19330;
assign w19332 = ~w19097 & ~w19331;
assign w19333 = (~w19330 & w31436) | (~w19330 & w31437) | (w31436 & w31437);
assign w19334 = ~w19332 & ~w19333;
assign w19335 = ~w18828 & ~w19074;
assign w19336 = w19334 & w19335;
assign w19337 = ~w19334 & ~w19335;
assign w19338 = ~w19336 & ~w19337;
assign w19339 = (w14835 & w31440) | (w14835 & w31441) | (w31440 & w31441);
assign w19340 = (w13761 & w37698) | (w13761 & w37699) | (w37698 & w37699);
assign w19341 = ~w19339 & ~w19340;
assign w19342 = (~w19110 & ~w19111) | (~w19110 & w31442) | (~w19111 & w31442);
assign w19343 = w1834 & w31443;
assign w19344 = b_63 & w1689;
assign w19345 = ~w19343 & ~w19344;
assign w19346 = ~w12671 & w31444;
assign w19347 = (a_23 & w19346) | (a_23 & w31445) | (w19346 & w31445);
assign w19348 = ~w19346 & w31446;
assign w19349 = ~w19347 & ~w19348;
assign w19350 = ~w19342 & ~w19349;
assign w19351 = w19342 & w19349;
assign w19352 = ~w19350 & ~w19351;
assign w19353 = b_61 & w2158;
assign w19354 = w2294 & w31447;
assign w19355 = b_60 & w2153;
assign w19356 = ~w19354 & ~w19355;
assign w19357 = ~w19353 & w19356;
assign w19358 = (w19357 & ~w11901) | (w19357 & w31448) | (~w11901 & w31448);
assign w19359 = (w11901 & w41427) | (w11901 & w41428) | (w41427 & w41428);
assign w19360 = (~w11901 & w41429) | (~w11901 & w41430) | (w41429 & w41430);
assign w19361 = ~w19358 & ~w19359;
assign w19362 = ~w19360 & ~w19361;
assign w19363 = ~w19112 & ~w19122;
assign w19364 = (~w19363 & w19125) | (~w19363 & w31449) | (w19125 & w31449);
assign w19365 = w19362 & w19364;
assign w19366 = ~w19362 & ~w19364;
assign w19367 = ~w19365 & ~w19366;
assign w19368 = (~w19138 & ~w19139) | (~w19138 & w31450) | (~w19139 & w31450);
assign w19369 = b_58 & w2639;
assign w19370 = w2820 & w31451;
assign w19371 = b_57 & w2634;
assign w19372 = ~w19370 & ~w19371;
assign w19373 = ~w19369 & w19372;
assign w19374 = w19372 & w31452;
assign w19375 = (~w10476 & w41431) | (~w10476 & w41432) | (w41431 & w41432);
assign w19376 = (w10476 & w31454) | (w10476 & w31455) | (w31454 & w31455);
assign w19377 = ~w19375 & ~w19376;
assign w19378 = (w19139 & w41433) | (w19139 & w41434) | (w41433 & w41434);
assign w19379 = (~w19139 & w41435) | (~w19139 & w41436) | (w41435 & w41436);
assign w19380 = ~w19378 & ~w19379;
assign w19381 = b_55 & w3195;
assign w19382 = w3388 & w31456;
assign w19383 = b_54 & w3190;
assign w19384 = ~w19382 & ~w19383;
assign w19385 = ~w19381 & w19384;
assign w19386 = (w19385 & ~w9776) | (w19385 & w31457) | (~w9776 & w31457);
assign w19387 = (w9776 & w41437) | (w9776 & w41438) | (w41437 & w41438);
assign w19388 = (~w9776 & w41439) | (~w9776 & w41440) | (w41439 & w41440);
assign w19389 = ~w19386 & ~w19387;
assign w19390 = ~w19388 & ~w19389;
assign w19391 = (w19390 & w19318) | (w19390 & w31458) | (w19318 & w31458);
assign w19392 = ~w19318 & w31459;
assign w19393 = ~w19391 & ~w19392;
assign w19394 = b_43 & w5962;
assign w19395 = w6246 & w31460;
assign w19396 = b_42 & w5957;
assign w19397 = ~w19395 & ~w19396;
assign w19398 = ~w19394 & w19397;
assign w19399 = (w19398 & ~w5888) | (w19398 & w31461) | (~w5888 & w31461);
assign w19400 = (w5888 & w41441) | (w5888 & w41442) | (w41441 & w41442);
assign w19401 = (~w5888 & w41443) | (~w5888 & w41444) | (w41443 & w41444);
assign w19402 = ~w19399 & ~w19400;
assign w19403 = ~w19401 & ~w19402;
assign w19404 = ~w19246 & ~w19251;
assign w19405 = b_40 & w6761;
assign w19406 = w7075 & w31462;
assign w19407 = b_39 & w6756;
assign w19408 = ~w19406 & ~w19407;
assign w19409 = ~w19405 & w19408;
assign w19410 = (w19409 & ~w5363) | (w19409 & w31463) | (~w5363 & w31463);
assign w19411 = (w5363 & w41445) | (w5363 & w41446) | (w41445 & w41446);
assign w19412 = (~w5363 & w41447) | (~w5363 & w41448) | (w41447 & w41448);
assign w19413 = ~w19410 & ~w19411;
assign w19414 = ~w19412 & ~w19413;
assign w19415 = (~w19230 & ~w19232) | (~w19230 & w31464) | (~w19232 & w31464);
assign w19416 = b_28 & w10562;
assign w19417 = w10902 & w31466;
assign w19418 = b_27 & w10557;
assign w19419 = ~w19417 & ~w19418;
assign w19420 = ~w19416 & w19419;
assign w19421 = (w19420 & ~w2771) | (w19420 & w31467) | (~w2771 & w31467);
assign w19422 = (w2771 & w41449) | (w2771 & w41450) | (w41449 & w41450);
assign w19423 = (~w2771 & w41451) | (~w2771 & w41452) | (w41451 & w41452);
assign w19424 = ~w19421 & ~w19422;
assign w19425 = ~w19423 & ~w19424;
assign w19426 = w12380 & w31469;
assign w19427 = b_22 & ~w12380;
assign w19428 = ~w19426 & ~w19427;
assign w19429 = (~w19145 & ~w19147) | (~w19145 & w31470) | (~w19147 & w31470);
assign w19430 = ~w19428 & w19429;
assign w19431 = w19428 & ~w19429;
assign w19432 = ~w19430 & ~w19431;
assign w19433 = b_25 & w11620;
assign w19434 = w11969 & w31471;
assign w19435 = b_24 & w11615;
assign w19436 = ~w19434 & ~w19435;
assign w19437 = ~w19433 & w19436;
assign w19438 = w19436 & w31472;
assign w19439 = (~w2108 & w41453) | (~w2108 & w41454) | (w41453 & w41454);
assign w19440 = (w19432 & w19439) | (w19432 & w31476) | (w19439 & w31476);
assign w19441 = ~w19439 & w31477;
assign w19442 = ~w19440 & ~w19441;
assign w19443 = (~w19164 & w31478) | (~w19164 & w31479) | (w31478 & w31479);
assign w19444 = (w19164 & w31480) | (w19164 & w31481) | (w31480 & w31481);
assign w19445 = ~w19443 & ~w19444;
assign w19446 = ~w19425 & w19445;
assign w19447 = w19425 & ~w19445;
assign w19448 = ~w19446 & ~w19447;
assign w19449 = (~w19183 & w31482) | (~w19183 & w31483) | (w31482 & w31483);
assign w19450 = (w19183 & w31484) | (w19183 & w31485) | (w31484 & w31485);
assign w19451 = ~w19449 & ~w19450;
assign w19452 = b_31 & w9534;
assign w19453 = w9876 & w31486;
assign w19454 = b_30 & w9529;
assign w19455 = ~w19453 & ~w19454;
assign w19456 = ~w19452 & w19455;
assign w19457 = (w19456 & ~w3345) | (w19456 & w31487) | (~w3345 & w31487);
assign w19458 = (w3345 & w41455) | (w3345 & w41456) | (w41455 & w41456);
assign w19459 = (~w3345 & w41457) | (~w3345 & w41458) | (w41457 & w41458);
assign w19460 = ~w19457 & ~w19458;
assign w19461 = ~w19459 & ~w19460;
assign w19462 = w19451 & ~w19461;
assign w19463 = w19451 & ~w19462;
assign w19464 = ~w19451 & ~w19461;
assign w19465 = ~w19463 & ~w19464;
assign w19466 = (~w19199 & w41459) | (~w19199 & w41460) | (w41459 & w41460);
assign w19467 = w19465 & w19466;
assign w19468 = ~w19465 & ~w19466;
assign w19469 = ~w19467 & ~w19468;
assign w19470 = b_34 & w8526;
assign w19471 = w8886 & w31488;
assign w19472 = b_33 & w8521;
assign w19473 = ~w19471 & ~w19472;
assign w19474 = ~w19470 & w19473;
assign w19475 = (w19474 & ~w3967) | (w19474 & w31489) | (~w3967 & w31489);
assign w19476 = (w3967 & w41461) | (w3967 & w41462) | (w41461 & w41462);
assign w19477 = (~w3967 & w41463) | (~w3967 & w41464) | (w41463 & w41464);
assign w19478 = ~w19475 & ~w19476;
assign w19479 = ~w19477 & ~w19478;
assign w19480 = w19469 & ~w19479;
assign w19481 = w19469 & ~w19480;
assign w19482 = ~w19469 & ~w19479;
assign w19483 = ~w19481 & ~w19482;
assign w19484 = ~w19215 & w31490;
assign w19485 = ~w31490 & ~w19215;
assign w19486 = w19483 & w19485;
assign w19487 = ~w19483 & ~w19485;
assign w19488 = ~w19486 & ~w19487;
assign w19489 = b_37 & w7613;
assign w19490 = w7941 & w31491;
assign w19491 = b_36 & w7608;
assign w19492 = ~w19490 & ~w19491;
assign w19493 = ~w19489 & w19492;
assign w19494 = (w19493 & ~w4636) | (w19493 & w31492) | (~w4636 & w31492);
assign w19495 = (w4636 & w41465) | (w4636 & w41466) | (w41465 & w41466);
assign w19496 = (~w4636 & w41467) | (~w4636 & w41468) | (w41467 & w41468);
assign w19497 = ~w19494 & ~w19495;
assign w19498 = ~w19496 & ~w19497;
assign w19499 = ~w19488 & w19498;
assign w19500 = w19488 & ~w19498;
assign w19501 = ~w19499 & ~w19500;
assign w19502 = ~w19415 & w19501;
assign w19503 = w19501 & ~w19502;
assign w19504 = (~w19414 & w19503) | (~w19414 & w31493) | (w19503 & w31493);
assign w19505 = ~w19503 & w31494;
assign w19506 = ~w19504 & ~w19505;
assign w19507 = ~w19404 & w19506;
assign w19508 = w19404 & ~w19506;
assign w19509 = ~w19507 & ~w19508;
assign w19510 = ~w19403 & w19509;
assign w19511 = w19509 & ~w19510;
assign w19512 = ~w19509 & ~w19403;
assign w19513 = (~w19263 & w19266) | (~w19263 & w31495) | (w19266 & w31495);
assign w19514 = ~w19511 & w31496;
assign w19515 = (~w19513 & w19511) | (~w19513 & w31497) | (w19511 & w31497);
assign w19516 = ~w19514 & ~w19515;
assign w19517 = b_46 & w5196;
assign w19518 = w5459 & w31498;
assign w19519 = b_45 & w5191;
assign w19520 = ~w19518 & ~w19519;
assign w19521 = ~w19517 & w19520;
assign w19522 = (w19521 & ~w6974) | (w19521 & w27623) | (~w6974 & w27623);
assign w19523 = (w6974 & w31499) | (w6974 & w31500) | (w31499 & w31500);
assign w19524 = (~w6974 & w31501) | (~w6974 & w31502) | (w31501 & w31502);
assign w19525 = ~w19522 & ~w19523;
assign w19526 = ~w19524 & ~w19525;
assign w19527 = w19516 & ~w19526;
assign w19528 = w19516 & ~w19527;
assign w19529 = ~w19516 & ~w19526;
assign w19530 = ~w19528 & ~w19529;
assign w19531 = (~w19281 & w19284) | (~w19281 & w31503) | (w19284 & w31503);
assign w19532 = w19530 & w19531;
assign w19533 = ~w19530 & ~w19531;
assign w19534 = ~w19532 & ~w19533;
assign w19535 = b_49 & w4499;
assign w19536 = w4723 & w31504;
assign w19537 = b_48 & w4494;
assign w19538 = ~w19536 & ~w19537;
assign w19539 = ~w19535 & w19538;
assign w19540 = (w19539 & ~w7859) | (w19539 & w31505) | (~w7859 & w31505);
assign w19541 = (w7859 & w41469) | (w7859 & w41470) | (w41469 & w41470);
assign w19542 = (~w7859 & w41471) | (~w7859 & w41472) | (w41471 & w41472);
assign w19543 = ~w19540 & ~w19541;
assign w19544 = ~w19542 & ~w19543;
assign w19545 = w19534 & ~w19544;
assign w19546 = w19534 & ~w19545;
assign w19547 = ~w19534 & ~w19544;
assign w19548 = ~w19546 & ~w19547;
assign w19549 = ~w19299 & ~w19304;
assign w19550 = w19548 & w19549;
assign w19551 = ~w19548 & ~w19549;
assign w19552 = ~w19550 & ~w19551;
assign w19553 = b_52 & w3803;
assign w19554 = w4027 & w31506;
assign w19555 = b_51 & w3798;
assign w19556 = ~w19554 & ~w19555;
assign w19557 = ~w19553 & w19556;
assign w19558 = (w19557 & ~w8793) | (w19557 & w31507) | (~w8793 & w31507);
assign w19559 = (w8793 & w41473) | (w8793 & w41474) | (w41473 & w41474);
assign w19560 = (~w8793 & w41475) | (~w8793 & w41476) | (w41475 & w41476);
assign w19561 = ~w19558 & ~w19559;
assign w19562 = ~w19560 & ~w19561;
assign w19563 = w19552 & ~w19562;
assign w19564 = w19552 & ~w19563;
assign w19565 = ~w19552 & ~w19562;
assign w19566 = ~w19564 & ~w19565;
assign w19567 = ~w19393 & ~w19566;
assign w19568 = w19393 & w19566;
assign w19569 = w19380 & w31508;
assign w19570 = w19380 & ~w19569;
assign w19571 = w31508 & ~w19380;
assign w19572 = ~w19570 & ~w19571;
assign w19573 = w19367 & ~w19572;
assign w19574 = ~w19367 & w19572;
assign w19575 = w19352 & w31509;
assign w19576 = w19352 & ~w19575;
assign w19577 = w31509 & ~w19352;
assign w19578 = ~w19576 & ~w19577;
assign w19579 = (~w19094 & ~w19330) | (~w19094 & w31510) | (~w19330 & w31510);
assign w19580 = w19578 & w19579;
assign w19581 = ~w19578 & ~w19579;
assign w19582 = ~w19580 & ~w19581;
assign w19583 = (w14835 & w31513) | (w14835 & w31514) | (w31513 & w31514);
assign w19584 = (w13761 & w37700) | (w13761 & w37701) | (w37700 & w37701);
assign w19585 = ~w19583 & ~w19584;
assign w19586 = (~w19350 & ~w19352) | (~w19350 & w31516) | (~w19352 & w31516);
assign w19587 = (~w19366 & ~w19367) | (~w19366 & w31517) | (~w19367 & w31517);
assign w19588 = w1834 & w31518;
assign w19589 = (~w19588 & ~w12670) | (~w19588 & w31519) | (~w12670 & w31519);
assign w19590 = (w12670 & w41477) | (w12670 & w41478) | (w41477 & w41478);
assign w19591 = (~w12670 & w41479) | (~w12670 & w41480) | (w41479 & w41480);
assign w19592 = ~w19589 & ~w19590;
assign w19593 = ~w19591 & ~w19592;
assign w19594 = ~w19587 & ~w19593;
assign w19595 = ~w19587 & ~w19594;
assign w19596 = w19587 & ~w19593;
assign w19597 = b_62 & w2158;
assign w19598 = w2294 & w31520;
assign w19599 = b_61 & w2153;
assign w19600 = ~w19598 & ~w19599;
assign w19601 = ~w19597 & w19600;
assign w19602 = (w19601 & ~w12273) | (w19601 & w31521) | (~w12273 & w31521);
assign w19603 = (w12273 & w41481) | (w12273 & w41482) | (w41481 & w41482);
assign w19604 = (~w12273 & w41483) | (~w12273 & w41484) | (w41483 & w41484);
assign w19605 = ~w19602 & ~w19603;
assign w19606 = ~w19604 & ~w19605;
assign w19607 = (~w19378 & ~w19380) | (~w19378 & w31522) | (~w19380 & w31522);
assign w19608 = w19606 & w19607;
assign w19609 = ~w19606 & ~w19607;
assign w19610 = ~w19608 & ~w19609;
assign w19611 = b_59 & w2639;
assign w19612 = w2820 & w31523;
assign w19613 = b_58 & w2634;
assign w19614 = ~w19612 & ~w19613;
assign w19615 = ~w19611 & w19614;
assign w19616 = (w19615 & ~w11169) | (w19615 & w31524) | (~w11169 & w31524);
assign w19617 = (w11169 & w41485) | (w11169 & w41486) | (w41485 & w41486);
assign w19618 = (~w11169 & w41487) | (~w11169 & w41488) | (w41487 & w41488);
assign w19619 = ~w19616 & ~w19617;
assign w19620 = ~w19618 & ~w19619;
assign w19621 = (~w19390 & w19318) | (~w19390 & w31525) | (w19318 & w31525);
assign w19622 = (~w19621 & w19566) | (~w19621 & w41489) | (w19566 & w41489);
assign w19623 = (~w19566 & w41490) | (~w19566 & w41491) | (w41490 & w41491);
assign w19624 = (w31527 & w19566) | (w31527 & w41492) | (w19566 & w41492);
assign w19625 = ~w19622 & ~w19623;
assign w19626 = ~w19624 & ~w19625;
assign w19627 = b_56 & w3195;
assign w19628 = w3388 & w31528;
assign w19629 = b_55 & w3190;
assign w19630 = ~w19628 & ~w19629;
assign w19631 = ~w19627 & w19630;
assign w19632 = (w19631 & ~w9798) | (w19631 & w26393) | (~w9798 & w26393);
assign w19633 = (w9798 & w31529) | (w9798 & w31530) | (w31529 & w31530);
assign w19634 = (~w9798 & w31531) | (~w9798 & w31532) | (w31531 & w31532);
assign w19635 = ~w19632 & ~w19633;
assign w19636 = ~w19634 & ~w19635;
assign w19637 = (~w19552 & w41493) | (~w19552 & w41494) | (w41493 & w41494);
assign w19638 = (w19552 & w41495) | (w19552 & w41496) | (w41495 & w41496);
assign w19639 = ~w19637 & ~w19638;
assign w19640 = b_53 & w3803;
assign w19641 = w4027 & w31534;
assign w19642 = b_52 & w3798;
assign w19643 = ~w19641 & ~w19642;
assign w19644 = ~w19640 & w19643;
assign w19645 = (w9109 & w41497) | (w9109 & w41498) | (w41497 & w41498);
assign w19646 = a_35 & ~w19645;
assign w19647 = w19645 & a_35;
assign w19648 = ~w19645 & ~w19646;
assign w19649 = ~w19647 & ~w19648;
assign w19650 = (~w19533 & ~w19534) | (~w19533 & w31536) | (~w19534 & w31536);
assign w19651 = (~w19507 & ~w19509) | (~w19507 & w31537) | (~w19509 & w31537);
assign w19652 = b_44 & w5962;
assign w19653 = w6246 & w31538;
assign w19654 = b_43 & w5957;
assign w19655 = ~w19653 & ~w19654;
assign w19656 = ~w19652 & w19655;
assign w19657 = (w19656 & ~w6408) | (w19656 & w31539) | (~w6408 & w31539);
assign w19658 = (w6408 & w41499) | (w6408 & w41500) | (w41499 & w41500);
assign w19659 = (~w6408 & w41501) | (~w6408 & w41502) | (w41501 & w41502);
assign w19660 = ~w19657 & ~w19658;
assign w19661 = ~w19659 & ~w19660;
assign w19662 = (~w19503 & w41503) | (~w19503 & w41504) | (w41503 & w41504);
assign w19663 = (~w19468 & ~w19469) | (~w19468 & w31540) | (~w19469 & w31540);
assign w19664 = b_35 & w8526;
assign w19665 = w8886 & w31541;
assign w19666 = b_34 & w8521;
assign w19667 = ~w19665 & ~w19666;
assign w19668 = ~w19664 & w19667;
assign w19669 = (w19668 & ~w4181) | (w19668 & w31542) | (~w4181 & w31542);
assign w19670 = (w4181 & w41505) | (w4181 & w41506) | (w41505 & w41506);
assign w19671 = (~w4181 & w41507) | (~w4181 & w41508) | (w41507 & w41508);
assign w19672 = ~w19669 & ~w19670;
assign w19673 = ~w19671 & ~w19672;
assign w19674 = (~w19449 & ~w19451) | (~w19449 & w31543) | (~w19451 & w31543);
assign w19675 = ~w19431 & ~w19440;
assign w19676 = w12380 & w31544;
assign w19677 = b_23 & ~w12380;
assign w19678 = ~w19676 & ~w19677;
assign w19679 = ~w19428 & w19678;
assign w19680 = w19428 & ~w19678;
assign w19681 = ~w19679 & ~w19680;
assign w19682 = b_26 & w11620;
assign w19683 = w11969 & w31545;
assign w19684 = b_25 & w11615;
assign w19685 = ~w19683 & ~w19684;
assign w19686 = ~w19682 & w19685;
assign w19687 = w19685 & w31546;
assign w19688 = (~w2416 & w41509) | (~w2416 & w41510) | (w41509 & w41510);
assign w19689 = (w19681 & w19688) | (w19681 & w31549) | (w19688 & w31549);
assign w19690 = ~w19688 & w31550;
assign w19691 = ~w19689 & ~w19690;
assign w19692 = ~w19675 & w19691;
assign w19693 = w19675 & ~w19691;
assign w19694 = ~w19692 & ~w19693;
assign w19695 = b_29 & w10562;
assign w19696 = w10902 & w31551;
assign w19697 = b_28 & w10557;
assign w19698 = ~w19696 & ~w19697;
assign w19699 = ~w19695 & w19698;
assign w19700 = (w19699 & ~w2954) | (w19699 & w31552) | (~w2954 & w31552);
assign w19701 = (w2954 & w41511) | (w2954 & w41512) | (w41511 & w41512);
assign w19702 = (~w2954 & w41513) | (~w2954 & w41514) | (w41513 & w41514);
assign w19703 = ~w19700 & ~w19701;
assign w19704 = ~w19702 & ~w19703;
assign w19705 = w19694 & ~w19704;
assign w19706 = w19694 & ~w19705;
assign w19707 = ~w19694 & ~w19704;
assign w19708 = ~w19706 & ~w19707;
assign w19709 = (~w19443 & ~w19445) | (~w19443 & w31553) | (~w19445 & w31553);
assign w19710 = w19708 & w19709;
assign w19711 = ~w19708 & ~w19709;
assign w19712 = ~w19710 & ~w19711;
assign w19713 = b_32 & w9534;
assign w19714 = w9876 & w31554;
assign w19715 = b_31 & w9529;
assign w19716 = ~w19714 & ~w19715;
assign w19717 = ~w19713 & w19716;
assign w19718 = (w19717 & ~w3545) | (w19717 & w31555) | (~w3545 & w31555);
assign w19719 = (w3545 & w41515) | (w3545 & w41516) | (w41515 & w41516);
assign w19720 = (~w3545 & w41517) | (~w3545 & w41518) | (w41517 & w41518);
assign w19721 = ~w19718 & ~w19719;
assign w19722 = ~w19720 & ~w19721;
assign w19723 = ~w19712 & w19722;
assign w19724 = w19712 & ~w19722;
assign w19725 = ~w19723 & ~w19724;
assign w19726 = ~w19674 & w19725;
assign w19727 = w19674 & ~w19725;
assign w19728 = ~w19726 & ~w19727;
assign w19729 = ~w19673 & w19728;
assign w19730 = w19673 & ~w19728;
assign w19731 = ~w19729 & ~w19730;
assign w19732 = ~w19663 & w19731;
assign w19733 = w19663 & ~w19731;
assign w19734 = ~w19732 & ~w19733;
assign w19735 = b_38 & w7613;
assign w19736 = w7941 & w31556;
assign w19737 = b_37 & w7608;
assign w19738 = ~w19736 & ~w19737;
assign w19739 = ~w19735 & w19738;
assign w19740 = (w19739 & ~w4658) | (w19739 & w31557) | (~w4658 & w31557);
assign w19741 = (w4658 & w41519) | (w4658 & w41520) | (w41519 & w41520);
assign w19742 = (~w4658 & w41521) | (~w4658 & w41522) | (w41521 & w41522);
assign w19743 = ~w19740 & ~w19741;
assign w19744 = ~w19742 & ~w19743;
assign w19745 = w19734 & ~w19744;
assign w19746 = w19734 & ~w19745;
assign w19747 = ~w19734 & ~w19744;
assign w19748 = ~w19746 & ~w19747;
assign w19749 = (~w19487 & ~w19488) | (~w19487 & w31558) | (~w19488 & w31558);
assign w19750 = ~w19748 & ~w19749;
assign w19751 = ~w19748 & ~w19750;
assign w19752 = ~w19749 & ~w19750;
assign w19753 = ~w19751 & ~w19752;
assign w19754 = b_41 & w6761;
assign w19755 = w7075 & w31559;
assign w19756 = b_40 & w6756;
assign w19757 = ~w19755 & ~w19756;
assign w19758 = ~w19754 & w19757;
assign w19759 = (w19758 & ~w5609) | (w19758 & w31560) | (~w5609 & w31560);
assign w19760 = (w5609 & w41523) | (w5609 & w41524) | (w41523 & w41524);
assign w19761 = (~w5609 & w41525) | (~w5609 & w41526) | (w41525 & w41526);
assign w19762 = ~w19759 & ~w19760;
assign w19763 = ~w19761 & ~w19762;
assign w19764 = ~w19753 & w19763;
assign w19765 = w19753 & ~w19763;
assign w19766 = ~w19764 & ~w19765;
assign w19767 = ~w19662 & ~w19766;
assign w19768 = w19662 & w19766;
assign w19769 = ~w19767 & ~w19768;
assign w19770 = ~w19661 & w19769;
assign w19771 = w19661 & ~w19769;
assign w19772 = ~w19770 & ~w19771;
assign w19773 = ~w19651 & w19772;
assign w19774 = w19651 & ~w19772;
assign w19775 = ~w19773 & ~w19774;
assign w19776 = b_47 & w5196;
assign w19777 = w5459 & w31561;
assign w19778 = b_46 & w5191;
assign w19779 = ~w19777 & ~w19778;
assign w19780 = ~w19776 & w19779;
assign w19781 = (w19780 & ~w6998) | (w19780 & w26694) | (~w6998 & w26694);
assign w19782 = (w6998 & w27624) | (w6998 & w27625) | (w27624 & w27625);
assign w19783 = (~w6998 & w31562) | (~w6998 & w31563) | (w31562 & w31563);
assign w19784 = ~w19781 & ~w19782;
assign w19785 = ~w19783 & ~w19784;
assign w19786 = w19775 & ~w19785;
assign w19787 = w19775 & ~w19786;
assign w19788 = ~w19775 & ~w19785;
assign w19789 = (~w19515 & ~w19516) | (~w19515 & w31564) | (~w19516 & w31564);
assign w19790 = ~w19787 & w31565;
assign w19791 = (~w19789 & w19787) | (~w19789 & w31566) | (w19787 & w31566);
assign w19792 = ~w19790 & ~w19791;
assign w19793 = b_50 & w4499;
assign w19794 = w4723 & w31567;
assign w19795 = b_49 & w4494;
assign w19796 = ~w19794 & ~w19795;
assign w19797 = ~w19793 & w19796;
assign w19798 = (w19797 & ~w8162) | (w19797 & w31568) | (~w8162 & w31568);
assign w19799 = (w8162 & w41527) | (w8162 & w41528) | (w41527 & w41528);
assign w19800 = (~w8162 & w41529) | (~w8162 & w41530) | (w41529 & w41530);
assign w19801 = ~w19798 & ~w19799;
assign w19802 = ~w19800 & ~w19801;
assign w19803 = ~w19792 & w19802;
assign w19804 = w19792 & ~w19802;
assign w19805 = ~w19803 & ~w19804;
assign w19806 = ~w19650 & w19805;
assign w19807 = ~w19650 & ~w19806;
assign w19808 = w19805 & ~w19806;
assign w19809 = ~w19807 & ~w19808;
assign w19810 = ~w19649 & ~w19809;
assign w19811 = w19809 & ~w19649;
assign w19812 = ~w19809 & ~w19810;
assign w19813 = ~w19811 & ~w19812;
assign w19814 = w19639 & ~w19813;
assign w19815 = w19639 & ~w19814;
assign w19816 = ~w19639 & ~w19813;
assign w19817 = ~w19815 & ~w19816;
assign w19818 = ~w19626 & w19817;
assign w19819 = w19626 & ~w19817;
assign w19820 = ~w19818 & ~w19819;
assign w19821 = w19610 & ~w19820;
assign w19822 = w19610 & ~w19821;
assign w19823 = ~w19610 & ~w19820;
assign w19824 = ~w19822 & ~w19823;
assign w19825 = (w19824 & w19595) | (w19824 & w31569) | (w19595 & w31569);
assign w19826 = ~w19595 & w31570;
assign w19827 = ~w19825 & ~w19826;
assign w19828 = ~w19586 & ~w19827;
assign w19829 = ~w19586 & ~w19828;
assign w19830 = ~w19827 & ~w19828;
assign w19831 = ~w19829 & ~w19830;
assign w19832 = (w14835 & w31571) | (w14835 & w31572) | (w31571 & w31572);
assign w19833 = (w13761 & w37702) | (w13761 & w37703) | (w37702 & w37703);
assign w19834 = ~w19832 & ~w19833;
assign w19835 = (~w19824 & w19595) | (~w19824 & w31575) | (w19595 & w31575);
assign w19836 = ~w19594 & ~w19835;
assign w19837 = (~w19609 & ~w19610) | (~w19609 & w31576) | (~w19610 & w31576);
assign w19838 = b_63 & w2158;
assign w19839 = w2294 & w31577;
assign w19840 = b_62 & w2153;
assign w19841 = ~w19839 & ~w19840;
assign w19842 = ~w19838 & w19841;
assign w19843 = (w19842 & ~w12646) | (w19842 & w31578) | (~w12646 & w31578);
assign w19844 = (w12646 & w41531) | (w12646 & w41532) | (w41531 & w41532);
assign w19845 = (~w12646 & w41533) | (~w12646 & w41534) | (w41533 & w41534);
assign w19846 = ~w19843 & ~w19844;
assign w19847 = ~w19845 & ~w19846;
assign w19848 = ~w19837 & ~w19847;
assign w19849 = ~w19837 & ~w19848;
assign w19850 = w19837 & ~w19847;
assign w19851 = (~w19623 & w19626) | (~w19623 & w31579) | (w19626 & w31579);
assign w19852 = b_60 & w2639;
assign w19853 = w2820 & w31580;
assign w19854 = b_59 & w2634;
assign w19855 = ~w19853 & ~w19854;
assign w19856 = ~w19852 & w19855;
assign w19857 = (w19856 & ~w11196) | (w19856 & w31581) | (~w11196 & w31581);
assign w19858 = (w11196 & w41535) | (w11196 & w41536) | (w41535 & w41536);
assign w19859 = (~w11196 & w41537) | (~w11196 & w41538) | (w41537 & w41538);
assign w19860 = ~w19857 & ~w19858;
assign w19861 = ~w19859 & ~w19860;
assign w19862 = ~w19851 & w19861;
assign w19863 = w19851 & ~w19861;
assign w19864 = ~w19862 & ~w19863;
assign w19865 = b_57 & w3195;
assign w19866 = w3388 & w31582;
assign w19867 = b_56 & w3190;
assign w19868 = ~w19866 & ~w19867;
assign w19869 = ~w19865 & w19868;
assign w19870 = (w19869 & ~w10452) | (w19869 & w31583) | (~w10452 & w31583);
assign w19871 = (w10452 & w41539) | (w10452 & w41540) | (w41539 & w41540);
assign w19872 = (~w10452 & w41541) | (~w10452 & w41542) | (w41541 & w41542);
assign w19873 = ~w19870 & ~w19871;
assign w19874 = ~w19872 & ~w19873;
assign w19875 = (~w19638 & ~w19639) | (~w19638 & w31584) | (~w19639 & w31584);
assign w19876 = (w31584 & w41543) | (w31584 & w41544) | (w41543 & w41544);
assign w19877 = (~w31584 & w41545) | (~w31584 & w41546) | (w41545 & w41546);
assign w19878 = ~w19876 & ~w19877;
assign w19879 = (~w19806 & w19809) | (~w19806 & w31585) | (w19809 & w31585);
assign w19880 = (~w19791 & ~w19792) | (~w19791 & w31586) | (~w19792 & w31586);
assign w19881 = (~w19767 & ~w19769) | (~w19767 & w31587) | (~w19769 & w31587);
assign w19882 = (~w19750 & w19753) | (~w19750 & w31588) | (w19753 & w31588);
assign w19883 = b_36 & w8526;
assign w19884 = w8886 & w31589;
assign w19885 = b_35 & w8521;
assign w19886 = ~w19884 & ~w19885;
assign w19887 = ~w19883 & w19886;
assign w19888 = (w19887 & ~w4395) | (w19887 & w31590) | (~w4395 & w31590);
assign w19889 = (w4395 & w41547) | (w4395 & w41548) | (w41547 & w41548);
assign w19890 = (~w4395 & w41549) | (~w4395 & w41550) | (w41549 & w41550);
assign w19891 = ~w19888 & ~w19889;
assign w19892 = ~w19890 & ~w19891;
assign w19893 = (~w19692 & ~w19694) | (~w19692 & w31591) | (~w19694 & w31591);
assign w19894 = ~w19679 & ~w19689;
assign w19895 = w12380 & w31592;
assign w19896 = b_24 & ~w12380;
assign w19897 = ~w19895 & ~w19896;
assign w19898 = ~a_23 & ~w19897;
assign w19899 = a_23 & w19897;
assign w19900 = ~w19898 & ~w19899;
assign w19901 = ~w19678 & w19900;
assign w19902 = w19678 & ~w19900;
assign w19903 = ~w19901 & ~w19902;
assign w19904 = b_27 & w11620;
assign w19905 = w11969 & w31593;
assign w19906 = b_26 & w11615;
assign w19907 = ~w19905 & ~w19906;
assign w19908 = ~w19904 & w19907;
assign w19909 = (w19908 & ~w2582) | (w19908 & w31594) | (~w2582 & w31594);
assign w19910 = (w2582 & w41551) | (w2582 & w41552) | (w41551 & w41552);
assign w19911 = (~w2582 & w41553) | (~w2582 & w41554) | (w41553 & w41554);
assign w19912 = ~w19909 & ~w19910;
assign w19913 = ~w19911 & ~w19912;
assign w19914 = (w19903 & w19912) | (w19903 & w31595) | (w19912 & w31595);
assign w19915 = w19903 & ~w19914;
assign w19916 = ~w19913 & ~w19914;
assign w19917 = ~w19915 & ~w19916;
assign w19918 = ~w19894 & w19917;
assign w19919 = w19894 & ~w19917;
assign w19920 = ~w19918 & ~w19919;
assign w19921 = b_30 & w10562;
assign w19922 = w10902 & w31596;
assign w19923 = b_29 & w10557;
assign w19924 = ~w19922 & ~w19923;
assign w19925 = ~w19921 & w19924;
assign w19926 = (w19925 & ~w3138) | (w19925 & w31597) | (~w3138 & w31597);
assign w19927 = (w3138 & w41555) | (w3138 & w41556) | (w41555 & w41556);
assign w19928 = (~w3138 & w41557) | (~w3138 & w41558) | (w41557 & w41558);
assign w19929 = ~w19926 & ~w19927;
assign w19930 = ~w19928 & ~w19929;
assign w19931 = ~w19920 & ~w19930;
assign w19932 = w19920 & w19930;
assign w19933 = ~w19931 & ~w19932;
assign w19934 = w19893 & ~w19933;
assign w19935 = ~w19893 & w19933;
assign w19936 = ~w19934 & ~w19935;
assign w19937 = b_33 & w9534;
assign w19938 = w9876 & w31598;
assign w19939 = b_32 & w9529;
assign w19940 = ~w19938 & ~w19939;
assign w19941 = ~w19937 & w19940;
assign w19942 = (w19941 & ~w3744) | (w19941 & w31599) | (~w3744 & w31599);
assign w19943 = (w3744 & w41559) | (w3744 & w41560) | (w41559 & w41560);
assign w19944 = (~w3744 & w41561) | (~w3744 & w41562) | (w41561 & w41562);
assign w19945 = ~w19942 & ~w19943;
assign w19946 = ~w19944 & ~w19945;
assign w19947 = (~w19711 & ~w19712) | (~w19711 & w31600) | (~w19712 & w31600);
assign w19948 = ~w19946 & ~w19947;
assign w19949 = w19946 & w19947;
assign w19950 = ~w19948 & ~w19949;
assign w19951 = w19936 & w19950;
assign w19952 = ~w19936 & ~w19950;
assign w19953 = ~w19951 & ~w19952;
assign w19954 = ~w19892 & w19953;
assign w19955 = w19953 & ~w19954;
assign w19956 = ~w19953 & ~w19892;
assign w19957 = (~w19726 & ~w19728) | (~w19726 & w31601) | (~w19728 & w31601);
assign w19958 = ~w19955 & w31602;
assign w19959 = (~w19957 & w19955) | (~w19957 & w31603) | (w19955 & w31603);
assign w19960 = ~w19958 & ~w19959;
assign w19961 = b_39 & w7613;
assign w19962 = w7941 & w31604;
assign w19963 = b_38 & w7608;
assign w19964 = ~w19962 & ~w19963;
assign w19965 = ~w19961 & w19964;
assign w19966 = (w19965 & ~w4888) | (w19965 & w27626) | (~w4888 & w27626);
assign w19967 = (w4888 & w31605) | (w4888 & w31606) | (w31605 & w31606);
assign w19968 = (~w4888 & w31607) | (~w4888 & w31608) | (w31607 & w31608);
assign w19969 = ~w19966 & ~w19967;
assign w19970 = ~w19968 & ~w19969;
assign w19971 = w19960 & ~w19970;
assign w19972 = w19960 & ~w19971;
assign w19973 = ~w19960 & ~w19970;
assign w19974 = ~w19972 & ~w19973;
assign w19975 = (~w19732 & ~w19734) | (~w19732 & w31609) | (~w19734 & w31609);
assign w19976 = w19974 & w19975;
assign w19977 = ~w19974 & ~w19975;
assign w19978 = ~w19976 & ~w19977;
assign w19979 = b_42 & w6761;
assign w19980 = w7075 & w31610;
assign w19981 = b_41 & w6756;
assign w19982 = ~w19980 & ~w19981;
assign w19983 = ~w19979 & w19982;
assign w19984 = (w19983 & ~w5864) | (w19983 & w26695) | (~w5864 & w26695);
assign w19985 = (w5864 & w27627) | (w5864 & w27628) | (w27627 & w27628);
assign w19986 = (~w5864 & w31611) | (~w5864 & w31612) | (w31611 & w31612);
assign w19987 = ~w19984 & ~w19985;
assign w19988 = ~w19986 & ~w19987;
assign w19989 = w19978 & ~w19988;
assign w19990 = w19978 & ~w19989;
assign w19991 = ~w19978 & ~w19988;
assign w19992 = ~w19990 & ~w19991;
assign w19993 = ~w19882 & w19992;
assign w19994 = w19882 & ~w19992;
assign w19995 = ~w19993 & ~w19994;
assign w19996 = b_45 & w5962;
assign w19997 = w6246 & w31613;
assign w19998 = b_44 & w5957;
assign w19999 = ~w19997 & ~w19998;
assign w20000 = ~w19996 & w19999;
assign w20001 = (w20000 & ~w6682) | (w20000 & w26696) | (~w6682 & w26696);
assign w20002 = (w6682 & w27629) | (w6682 & w27630) | (w27629 & w27630);
assign w20003 = (~w6682 & w31614) | (~w6682 & w31615) | (w31614 & w31615);
assign w20004 = ~w20001 & ~w20002;
assign w20005 = ~w20003 & ~w20004;
assign w20006 = ~w19995 & ~w20005;
assign w20007 = w19995 & w20005;
assign w20008 = ~w20006 & ~w20007;
assign w20009 = w19881 & ~w20008;
assign w20010 = ~w19881 & w20008;
assign w20011 = ~w20009 & ~w20010;
assign w20012 = b_48 & w5196;
assign w20013 = w5459 & w31616;
assign w20014 = b_47 & w5191;
assign w20015 = ~w20013 & ~w20014;
assign w20016 = ~w20012 & w20015;
assign w20017 = (w20016 & ~w7284) | (w20016 & w26394) | (~w7284 & w26394);
assign w20018 = (w7284 & w26697) | (w7284 & w26698) | (w26697 & w26698);
assign w20019 = (~w7284 & w27631) | (~w7284 & w27632) | (w27631 & w27632);
assign w20020 = ~w20017 & ~w20018;
assign w20021 = ~w20019 & ~w20020;
assign w20022 = w20011 & ~w20021;
assign w20023 = w20021 & w20011;
assign w20024 = ~w20011 & ~w20021;
assign w20025 = ~w20023 & ~w20024;
assign w20026 = (~w19773 & ~w19775) | (~w19773 & w31617) | (~w19775 & w31617);
assign w20027 = w20025 & w20026;
assign w20028 = (~w20026 & w20024) | (~w20026 & w27633) | (w20024 & w27633);
assign w20029 = b_51 & w4499;
assign w20030 = w4723 & w31618;
assign w20031 = b_50 & w4494;
assign w20032 = ~w20030 & ~w20031;
assign w20033 = ~w20029 & w20032;
assign w20034 = (w20033 & ~w8186) | (w20033 & w31619) | (~w8186 & w31619);
assign w20035 = (w8186 & w41563) | (w8186 & w41564) | (w41563 & w41564);
assign w20036 = (~w8186 & w41565) | (~w8186 & w41566) | (w41565 & w41566);
assign w20037 = ~w20034 & ~w20035;
assign w20038 = ~w20036 & ~w20037;
assign w20039 = ~w20028 & w31620;
assign w20040 = (w20038 & w20028) | (w20038 & w31621) | (w20028 & w31621);
assign w20041 = ~w19880 & w31622;
assign w20042 = ~w19880 & ~w20041;
assign w20043 = (~w20039 & w19880) | (~w20039 & w41567) | (w19880 & w41567);
assign w20044 = w19880 & w31622;
assign w20045 = ~w20042 & ~w20044;
assign w20046 = b_54 & w3803;
assign w20047 = w4027 & w31623;
assign w20048 = b_53 & w3798;
assign w20049 = ~w20047 & ~w20048;
assign w20050 = ~w20046 & w20049;
assign w20051 = (w20050 & ~w9134) | (w20050 & w31624) | (~w9134 & w31624);
assign w20052 = (w9134 & w41568) | (w9134 & w41569) | (w41568 & w41569);
assign w20053 = (~w9134 & w41570) | (~w9134 & w41571) | (w41570 & w41571);
assign w20054 = ~w20051 & ~w20052;
assign w20055 = ~w20053 & ~w20054;
assign w20056 = ~w20042 & w41572;
assign w20057 = (~w20055 & w20042) | (~w20055 & w41573) | (w20042 & w41573);
assign w20058 = ~w20056 & ~w20057;
assign w20059 = ~w19879 & w20058;
assign w20060 = w19879 & ~w20058;
assign w20061 = ~w20059 & ~w20060;
assign w20062 = w19878 & w20061;
assign w20063 = ~w19878 & ~w20061;
assign w20064 = ~w19864 & w31625;
assign w20065 = ~w19864 & ~w20064;
assign w20066 = w31625 & w19864;
assign w20067 = ~w20065 & ~w20066;
assign w20068 = (w20067 & w19849) | (w20067 & w31626) | (w19849 & w31626);
assign w20069 = ~w19849 & w31627;
assign w20070 = ~w20068 & ~w20069;
assign w20071 = (~w20070 & w19835) | (~w20070 & w41574) | (w19835 & w41574);
assign w20072 = ~w19836 & ~w20071;
assign w20073 = ~w19835 & w41575;
assign w20074 = ~w20072 & ~w20073;
assign w20075 = (w14835 & w31628) | (w14835 & w31629) | (w31628 & w31629);
assign w20076 = (w13761 & w37704) | (w13761 & w37705) | (w37704 & w37705);
assign w20077 = ~w20075 & ~w20076;
assign w20078 = (~w20067 & w19849) | (~w20067 & w31632) | (w19849 & w31632);
assign w20079 = ~w19848 & ~w20078;
assign w20080 = b_61 & w2639;
assign w20081 = w2820 & w31633;
assign w20082 = b_60 & w2634;
assign w20083 = ~w20081 & ~w20082;
assign w20084 = ~w20080 & w20083;
assign w20085 = (w20084 & ~w11901) | (w20084 & w31634) | (~w11901 & w31634);
assign w20086 = (w11901 & w41576) | (w11901 & w41577) | (w41576 & w41577);
assign w20087 = (~w11901 & w41578) | (~w11901 & w41579) | (w41578 & w41579);
assign w20088 = ~w20085 & ~w20086;
assign w20089 = ~w20087 & ~w20088;
assign w20090 = (~w19877 & ~w19878) | (~w19877 & w31635) | (~w19878 & w31635);
assign w20091 = ~w20089 & ~w20090;
assign w20092 = w20090 & ~w20089;
assign w20093 = ~w20090 & ~w20091;
assign w20094 = ~w20092 & ~w20093;
assign w20095 = b_58 & w3195;
assign w20096 = w3388 & w31636;
assign w20097 = b_57 & w3190;
assign w20098 = ~w20096 & ~w20097;
assign w20099 = ~w20095 & w20098;
assign w20100 = w20098 & w31637;
assign w20101 = (~w10476 & w41580) | (~w10476 & w41581) | (w41580 & w41581);
assign w20102 = (w10476 & w31639) | (w10476 & w31640) | (w31639 & w31640);
assign w20103 = ~w20101 & ~w20102;
assign w20104 = (~w19879 & w41582) | (~w19879 & w41583) | (w41582 & w41583);
assign w20105 = (w31642 & w19879) | (w31642 & w41584) | (w19879 & w41584);
assign w20106 = ~w20104 & ~w20105;
assign w20107 = b_43 & w6761;
assign w20108 = w7075 & w31643;
assign w20109 = b_42 & w6756;
assign w20110 = ~w20108 & ~w20109;
assign w20111 = ~w20107 & w20110;
assign w20112 = (w20111 & ~w5888) | (w20111 & w26699) | (~w5888 & w26699);
assign w20113 = (w5888 & w27634) | (w5888 & w27635) | (w27634 & w27635);
assign w20114 = (~w5888 & w31644) | (~w5888 & w31645) | (w31644 & w31645);
assign w20115 = ~w20112 & ~w20113;
assign w20116 = ~w20114 & ~w20115;
assign w20117 = (~w19971 & w19974) | (~w19971 & w41585) | (w19974 & w41585);
assign w20118 = b_40 & w7613;
assign w20119 = w7941 & w31646;
assign w20120 = b_39 & w7608;
assign w20121 = ~w20119 & ~w20120;
assign w20122 = ~w20118 & w20121;
assign w20123 = (w20122 & ~w5363) | (w20122 & w27636) | (~w5363 & w27636);
assign w20124 = (w5363 & w31647) | (w5363 & w31648) | (w31647 & w31648);
assign w20125 = (~w5363 & w31649) | (~w5363 & w31650) | (w31649 & w31650);
assign w20126 = ~w20123 & ~w20124;
assign w20127 = ~w20125 & ~w20126;
assign w20128 = ~w19954 & ~w19959;
assign w20129 = w12380 & w41586;
assign w20130 = b_25 & ~w12380;
assign w20131 = ~w20129 & ~w20130;
assign w20132 = (~w19898 & ~w19900) | (~w19898 & w31652) | (~w19900 & w31652);
assign w20133 = ~w20131 & w20132;
assign w20134 = w20131 & ~w20132;
assign w20135 = ~w20133 & ~w20134;
assign w20136 = b_28 & w11620;
assign w20137 = w11969 & w31653;
assign w20138 = b_27 & w11615;
assign w20139 = ~w20137 & ~w20138;
assign w20140 = ~w20136 & w20139;
assign w20141 = w20139 & w31654;
assign w20142 = (~w2771 & w41587) | (~w2771 & w41588) | (w41587 & w41588);
assign w20143 = (w20135 & w20142) | (w20135 & w31658) | (w20142 & w31658);
assign w20144 = ~w20142 & w31659;
assign w20145 = ~w20143 & ~w20144;
assign w20146 = (~w19917 & w31660) | (~w19917 & w31661) | (w31660 & w31661);
assign w20147 = (w19917 & w31662) | (w19917 & w31663) | (w31662 & w31663);
assign w20148 = ~w20146 & ~w20147;
assign w20149 = b_31 & w10562;
assign w20150 = w10902 & w31664;
assign w20151 = b_30 & w10557;
assign w20152 = ~w20150 & ~w20151;
assign w20153 = ~w20149 & w20152;
assign w20154 = (w20153 & ~w3345) | (w20153 & w31665) | (~w3345 & w31665);
assign w20155 = (w3345 & w41589) | (w3345 & w41590) | (w41589 & w41590);
assign w20156 = (~w3345 & w41591) | (~w3345 & w41592) | (w41591 & w41592);
assign w20157 = ~w20154 & ~w20155;
assign w20158 = ~w20156 & ~w20157;
assign w20159 = w20148 & ~w20158;
assign w20160 = w20148 & ~w20159;
assign w20161 = ~w20148 & ~w20158;
assign w20162 = ~w20160 & ~w20161;
assign w20163 = (~w19931 & ~w19933) | (~w19931 & w31666) | (~w19933 & w31666);
assign w20164 = w20162 & w20163;
assign w20165 = ~w20162 & ~w20163;
assign w20166 = ~w20164 & ~w20165;
assign w20167 = b_34 & w9534;
assign w20168 = w9876 & w31667;
assign w20169 = b_33 & w9529;
assign w20170 = ~w20168 & ~w20169;
assign w20171 = ~w20167 & w20170;
assign w20172 = (w20171 & ~w3967) | (w20171 & w31668) | (~w3967 & w31668);
assign w20173 = (w3967 & w41593) | (w3967 & w41594) | (w41593 & w41594);
assign w20174 = (~w3967 & w41595) | (~w3967 & w41596) | (w41595 & w41596);
assign w20175 = ~w20172 & ~w20173;
assign w20176 = ~w20174 & ~w20175;
assign w20177 = w20166 & ~w20176;
assign w20178 = w20166 & ~w20177;
assign w20179 = ~w20166 & ~w20176;
assign w20180 = ~w20178 & ~w20179;
assign w20181 = (~w19948 & ~w19950) | (~w19948 & w31669) | (~w19950 & w31669);
assign w20182 = w20180 & w20181;
assign w20183 = ~w20180 & ~w20181;
assign w20184 = ~w20182 & ~w20183;
assign w20185 = b_37 & w8526;
assign w20186 = w8886 & w31670;
assign w20187 = b_36 & w8521;
assign w20188 = ~w20186 & ~w20187;
assign w20189 = ~w20185 & w20188;
assign w20190 = (w20189 & ~w4636) | (w20189 & w31671) | (~w4636 & w31671);
assign w20191 = (w4636 & w41597) | (w4636 & w41598) | (w41597 & w41598);
assign w20192 = (~w4636 & w41599) | (~w4636 & w41600) | (w41599 & w41600);
assign w20193 = ~w20190 & ~w20191;
assign w20194 = ~w20192 & ~w20193;
assign w20195 = ~w20184 & w20194;
assign w20196 = w20184 & ~w20194;
assign w20197 = ~w20195 & ~w20196;
assign w20198 = ~w20128 & w20197;
assign w20199 = ~w20128 & ~w20198;
assign w20200 = w20197 & ~w20198;
assign w20201 = ~w20199 & ~w20200;
assign w20202 = ~w20127 & ~w20201;
assign w20203 = (w20127 & w20198) | (w20127 & w31672) | (w20198 & w31672);
assign w20204 = ~w20199 & w20203;
assign w20205 = ~w20202 & ~w20204;
assign w20206 = ~w20117 & w20205;
assign w20207 = w20117 & ~w20205;
assign w20208 = ~w20206 & ~w20207;
assign w20209 = ~w20116 & w20208;
assign w20210 = w20208 & ~w20209;
assign w20211 = ~w20208 & ~w20116;
assign w20212 = ~w20210 & ~w20211;
assign w20213 = (~w19989 & w19882) | (~w19989 & w31673) | (w19882 & w31673);
assign w20214 = w20212 & w20213;
assign w20215 = ~w20212 & ~w20213;
assign w20216 = ~w20214 & ~w20215;
assign w20217 = b_46 & w5962;
assign w20218 = w6246 & w31674;
assign w20219 = b_45 & w5957;
assign w20220 = ~w20218 & ~w20219;
assign w20221 = ~w20217 & w20220;
assign w20222 = (w20221 & ~w6974) | (w20221 & w26395) | (~w6974 & w26395);
assign w20223 = (w6974 & w26700) | (w6974 & w26701) | (w26700 & w26701);
assign w20224 = (~w6974 & w27637) | (~w6974 & w27638) | (w27637 & w27638);
assign w20225 = ~w20222 & ~w20223;
assign w20226 = ~w20224 & ~w20225;
assign w20227 = w20216 & ~w20226;
assign w20228 = w20226 & w20216;
assign w20229 = ~w20216 & ~w20226;
assign w20230 = ~w20228 & ~w20229;
assign w20231 = ~w20006 & ~w20010;
assign w20232 = w20230 & w20231;
assign w20233 = ~w20230 & ~w20231;
assign w20234 = ~w20232 & ~w20233;
assign w20235 = b_49 & w5196;
assign w20236 = w5459 & w31675;
assign w20237 = b_48 & w5191;
assign w20238 = ~w20236 & ~w20237;
assign w20239 = ~w20235 & w20238;
assign w20240 = (w20239 & ~w7859) | (w20239 & w26396) | (~w7859 & w26396);
assign w20241 = (w7859 & w27639) | (w7859 & w27640) | (w27639 & w27640);
assign w20242 = (~w7859 & w31676) | (~w7859 & w31677) | (w31676 & w31677);
assign w20243 = ~w20240 & ~w20241;
assign w20244 = ~w20242 & ~w20243;
assign w20245 = w20234 & ~w20244;
assign w20246 = w20234 & ~w20245;
assign w20247 = ~w20234 & ~w20244;
assign w20248 = ~w20246 & ~w20247;
assign w20249 = (~w27633 & w31678) | (~w27633 & w31679) | (w31678 & w31679);
assign w20250 = w20248 & w20249;
assign w20251 = ~w20248 & ~w20249;
assign w20252 = ~w20250 & ~w20251;
assign w20253 = b_52 & w4499;
assign w20254 = w4723 & w31680;
assign w20255 = b_51 & w4494;
assign w20256 = ~w20254 & ~w20255;
assign w20257 = ~w20253 & w20256;
assign w20258 = (w20257 & ~w8793) | (w20257 & w31681) | (~w8793 & w31681);
assign w20259 = (w8793 & w41601) | (w8793 & w41602) | (w41601 & w41602);
assign w20260 = (~w8793 & w41603) | (~w8793 & w41604) | (w41603 & w41604);
assign w20261 = ~w20258 & ~w20259;
assign w20262 = ~w20260 & ~w20261;
assign w20263 = w20252 & ~w20262;
assign w20264 = w20252 & ~w20263;
assign w20265 = ~w20252 & ~w20262;
assign w20266 = ~w20264 & w31682;
assign w20267 = (w20043 & w20264) | (w20043 & w31683) | (w20264 & w31683);
assign w20268 = ~w20266 & ~w20267;
assign w20269 = b_55 & w3803;
assign w20270 = w4027 & w31684;
assign w20271 = b_54 & w3798;
assign w20272 = ~w20270 & ~w20271;
assign w20273 = ~w20269 & w20272;
assign w20274 = (w20273 & ~w9776) | (w20273 & w31685) | (~w9776 & w31685);
assign w20275 = (w9776 & w41605) | (w9776 & w41606) | (w41605 & w41606);
assign w20276 = (~w9776 & w41607) | (~w9776 & w41608) | (w41607 & w41608);
assign w20277 = ~w20274 & ~w20275;
assign w20278 = ~w20276 & ~w20277;
assign w20279 = ~w20268 & ~w20278;
assign w20280 = w20268 & w20278;
assign w20281 = ~w20279 & ~w20280;
assign w20282 = w20106 & w20281;
assign w20283 = ~w20106 & ~w20281;
assign w20284 = ~w20282 & ~w20283;
assign w20285 = (w20284 & w20093) | (w20284 & w31686) | (w20093 & w31686);
assign w20286 = ~w20094 & ~w20285;
assign w20287 = ~w20093 & w41609;
assign w20288 = ~w20286 & ~w20287;
assign w20289 = ~w19851 & ~w19861;
assign w20290 = (~w20289 & w19864) | (~w20289 & w31687) | (w19864 & w31687);
assign w20291 = w2294 & w31688;
assign w20292 = b_63 & w2153;
assign w20293 = ~w20291 & ~w20292;
assign w20294 = ~w12671 & w31689;
assign w20295 = (a_26 & w20294) | (a_26 & w31690) | (w20294 & w31690);
assign w20296 = ~w20294 & w31691;
assign w20297 = ~w20295 & ~w20296;
assign w20298 = ~w20290 & ~w20297;
assign w20299 = ~w20290 & ~w20298;
assign w20300 = w20290 & ~w20297;
assign w20301 = (~w20288 & w20299) | (~w20288 & w31692) | (w20299 & w31692);
assign w20302 = w20288 & ~w20300;
assign w20303 = ~w20299 & w20302;
assign w20304 = ~w20301 & ~w20303;
assign w20305 = ~w20079 & w20304;
assign w20306 = ~w20079 & ~w20305;
assign w20307 = w20079 & w20304;
assign w20308 = ~w20306 & ~w20307;
assign w20309 = (w14835 & w31693) | (w14835 & w31694) | (w31693 & w31694);
assign w20310 = (w13761 & w37706) | (w13761 & w37707) | (w37706 & w37707);
assign w20311 = ~w20309 & ~w20310;
assign w20312 = (~w20093 & w41610) | (~w20093 & w41611) | (w41610 & w41611);
assign w20313 = w2294 & w31699;
assign w20314 = (~w20313 & ~w12670) | (~w20313 & w31700) | (~w12670 & w31700);
assign w20315 = (w12670 & w41612) | (w12670 & w41613) | (w41612 & w41613);
assign w20316 = (~w12670 & w41614) | (~w12670 & w41615) | (w41614 & w41615);
assign w20317 = ~w20314 & ~w20315;
assign w20318 = ~w20316 & ~w20317;
assign w20319 = (w20093 & w41616) | (w20093 & w41617) | (w41616 & w41617);
assign w20320 = ~w20312 & ~w20319;
assign w20321 = b_62 & w2639;
assign w20322 = w2820 & w31703;
assign w20323 = b_61 & w2634;
assign w20324 = ~w20322 & ~w20323;
assign w20325 = ~w20321 & w20324;
assign w20326 = (w20325 & ~w12273) | (w20325 & w31704) | (~w12273 & w31704);
assign w20327 = (w12273 & w41618) | (w12273 & w41619) | (w41618 & w41619);
assign w20328 = (~w12273 & w41620) | (~w12273 & w41621) | (w41620 & w41621);
assign w20329 = ~w20326 & ~w20327;
assign w20330 = ~w20328 & ~w20329;
assign w20331 = (~w20104 & ~w20106) | (~w20104 & w31705) | (~w20106 & w31705);
assign w20332 = w20330 & w20331;
assign w20333 = ~w20330 & ~w20331;
assign w20334 = ~w20332 & ~w20333;
assign w20335 = b_59 & w3195;
assign w20336 = w3388 & w31706;
assign w20337 = b_58 & w3190;
assign w20338 = ~w20336 & ~w20337;
assign w20339 = ~w20335 & w20338;
assign w20340 = (w20339 & ~w11169) | (w20339 & w31707) | (~w11169 & w31707);
assign w20341 = (w11169 & w41622) | (w11169 & w41623) | (w41622 & w41623);
assign w20342 = (~w11169 & w41624) | (~w11169 & w41625) | (w41624 & w41625);
assign w20343 = ~w20340 & ~w20341;
assign w20344 = ~w20342 & ~w20343;
assign w20345 = (~w20043 & w20264) | (~w20043 & w31708) | (w20264 & w31708);
assign w20346 = (~w20345 & w20268) | (~w20345 & w27641) | (w20268 & w27641);
assign w20347 = w20344 & w20346;
assign w20348 = ~w20344 & ~w20346;
assign w20349 = ~w20347 & ~w20348;
assign w20350 = b_56 & w3803;
assign w20351 = w4027 & w31709;
assign w20352 = b_55 & w3798;
assign w20353 = ~w20351 & ~w20352;
assign w20354 = ~w20350 & w20353;
assign w20355 = (w20354 & ~w9798) | (w20354 & w31710) | (~w9798 & w31710);
assign w20356 = (w9798 & w41626) | (w9798 & w41627) | (w41626 & w41627);
assign w20357 = (~w9798 & w41628) | (~w9798 & w41629) | (w41628 & w41629);
assign w20358 = ~w20355 & ~w20356;
assign w20359 = ~w20357 & ~w20358;
assign w20360 = (~w20251 & ~w20252) | (~w20251 & w31711) | (~w20252 & w31711);
assign w20361 = b_53 & w4499;
assign w20362 = w4723 & w31712;
assign w20363 = b_52 & w4494;
assign w20364 = ~w20362 & ~w20363;
assign w20365 = ~w20361 & w20364;
assign w20366 = (w9109 & w41630) | (w9109 & w41631) | (w41630 & w41631);
assign w20367 = a_38 & ~w20366;
assign w20368 = w20366 & a_38;
assign w20369 = ~w20366 & ~w20367;
assign w20370 = ~w20368 & ~w20369;
assign w20371 = (~w20233 & ~w20234) | (~w20233 & w31714) | (~w20234 & w31714);
assign w20372 = (~w20206 & ~w20208) | (~w20206 & w31715) | (~w20208 & w31715);
assign w20373 = b_44 & w6761;
assign w20374 = w7075 & w31716;
assign w20375 = b_43 & w6756;
assign w20376 = ~w20374 & ~w20375;
assign w20377 = ~w20373 & w20376;
assign w20378 = (w20377 & ~w6408) | (w20377 & w26397) | (~w6408 & w26397);
assign w20379 = (w6408 & w31717) | (w6408 & w31718) | (w31717 & w31718);
assign w20380 = (~w6408 & w31719) | (~w6408 & w31720) | (w31719 & w31720);
assign w20381 = ~w20378 & ~w20379;
assign w20382 = ~w20380 & ~w20381;
assign w20383 = (~w20198 & w20201) | (~w20198 & w31721) | (w20201 & w31721);
assign w20384 = (~w20165 & ~w20166) | (~w20165 & w31722) | (~w20166 & w31722);
assign w20385 = b_35 & w9534;
assign w20386 = w9876 & w31723;
assign w20387 = b_34 & w9529;
assign w20388 = ~w20386 & ~w20387;
assign w20389 = ~w20385 & w20388;
assign w20390 = (w20389 & ~w4181) | (w20389 & w31724) | (~w4181 & w31724);
assign w20391 = (w4181 & w41632) | (w4181 & w41633) | (w41632 & w41633);
assign w20392 = (~w4181 & w41634) | (~w4181 & w41635) | (w41634 & w41635);
assign w20393 = ~w20390 & ~w20391;
assign w20394 = ~w20392 & ~w20393;
assign w20395 = (~w20146 & ~w20148) | (~w20146 & w31725) | (~w20148 & w31725);
assign w20396 = b_32 & w10562;
assign w20397 = w10902 & w31726;
assign w20398 = b_31 & w10557;
assign w20399 = ~w20397 & ~w20398;
assign w20400 = ~w20396 & w20399;
assign w20401 = (w20400 & ~w3545) | (w20400 & w31727) | (~w3545 & w31727);
assign w20402 = (w3545 & w41636) | (w3545 & w41637) | (w41636 & w41637);
assign w20403 = (~w3545 & w41638) | (~w3545 & w41639) | (w41638 & w41639);
assign w20404 = ~w20401 & ~w20402;
assign w20405 = ~w20403 & ~w20404;
assign w20406 = ~w20134 & ~w20143;
assign w20407 = w12380 & w31728;
assign w20408 = b_26 & ~w12380;
assign w20409 = ~w20407 & ~w20408;
assign w20410 = ~w20131 & w20409;
assign w20411 = w20131 & ~w20409;
assign w20412 = ~w20410 & ~w20411;
assign w20413 = b_29 & w11620;
assign w20414 = w11969 & w31729;
assign w20415 = b_28 & w11615;
assign w20416 = ~w20414 & ~w20415;
assign w20417 = ~w20413 & w20416;
assign w20418 = w20416 & w31730;
assign w20419 = (~w2954 & w41640) | (~w2954 & w41641) | (w41640 & w41641);
assign w20420 = (w20412 & w20419) | (w20412 & w31734) | (w20419 & w31734);
assign w20421 = ~w20419 & w31735;
assign w20422 = ~w20420 & ~w20421;
assign w20423 = ~w20406 & w20422;
assign w20424 = w20406 & ~w20422;
assign w20425 = ~w20423 & ~w20424;
assign w20426 = ~w20405 & w20425;
assign w20427 = w20405 & ~w20425;
assign w20428 = ~w20426 & ~w20427;
assign w20429 = ~w20395 & w20428;
assign w20430 = w20395 & ~w20428;
assign w20431 = ~w20429 & ~w20430;
assign w20432 = ~w20394 & w20431;
assign w20433 = w20394 & ~w20431;
assign w20434 = ~w20432 & ~w20433;
assign w20435 = ~w20384 & w20434;
assign w20436 = w20384 & ~w20434;
assign w20437 = ~w20435 & ~w20436;
assign w20438 = b_38 & w8526;
assign w20439 = w8886 & w31736;
assign w20440 = b_37 & w8521;
assign w20441 = ~w20439 & ~w20440;
assign w20442 = ~w20438 & w20441;
assign w20443 = (w20442 & ~w4658) | (w20442 & w31737) | (~w4658 & w31737);
assign w20444 = (w4658 & w41642) | (w4658 & w41643) | (w41642 & w41643);
assign w20445 = (~w4658 & w41644) | (~w4658 & w41645) | (w41644 & w41645);
assign w20446 = ~w20443 & ~w20444;
assign w20447 = ~w20445 & ~w20446;
assign w20448 = w20437 & ~w20447;
assign w20449 = w20437 & ~w20448;
assign w20450 = ~w20437 & ~w20447;
assign w20451 = ~w20449 & ~w20450;
assign w20452 = (~w20183 & ~w20184) | (~w20183 & w31738) | (~w20184 & w31738);
assign w20453 = ~w20451 & ~w20452;
assign w20454 = ~w20451 & ~w20453;
assign w20455 = ~w20452 & ~w20453;
assign w20456 = ~w20454 & ~w20455;
assign w20457 = b_41 & w7613;
assign w20458 = w7941 & w31739;
assign w20459 = b_40 & w7608;
assign w20460 = ~w20458 & ~w20459;
assign w20461 = ~w20457 & w20460;
assign w20462 = (w20461 & ~w5609) | (w20461 & w31740) | (~w5609 & w31740);
assign w20463 = (w5609 & w41646) | (w5609 & w41647) | (w41646 & w41647);
assign w20464 = (~w5609 & w41648) | (~w5609 & w41649) | (w41648 & w41649);
assign w20465 = ~w20462 & ~w20463;
assign w20466 = ~w20464 & ~w20465;
assign w20467 = ~w20456 & w20466;
assign w20468 = w20456 & ~w20466;
assign w20469 = ~w20467 & ~w20468;
assign w20470 = ~w20383 & ~w20469;
assign w20471 = w20383 & w20469;
assign w20472 = ~w20470 & ~w20471;
assign w20473 = ~w20382 & w20472;
assign w20474 = w20382 & ~w20472;
assign w20475 = ~w20473 & ~w20474;
assign w20476 = ~w20372 & w20475;
assign w20477 = w20372 & ~w20475;
assign w20478 = ~w20476 & ~w20477;
assign w20479 = b_47 & w5962;
assign w20480 = w6246 & w31741;
assign w20481 = b_46 & w5957;
assign w20482 = ~w20480 & ~w20481;
assign w20483 = ~w20479 & w20482;
assign w20484 = (w20483 & ~w6998) | (w20483 & w25676) | (~w6998 & w25676);
assign w20485 = (w6998 & w26004) | (w6998 & w26005) | (w26004 & w26005);
assign w20486 = (~w6998 & w26398) | (~w6998 & w26399) | (w26398 & w26399);
assign w20487 = ~w20484 & ~w20485;
assign w20488 = ~w20486 & ~w20487;
assign w20489 = w20488 & w20478;
assign w20490 = ~w20478 & ~w20488;
assign w20491 = (~w20215 & ~w20216) | (~w20215 & w41650) | (~w20216 & w41650);
assign w20492 = w20491 & w31742;
assign w20493 = (~w20491 & w20490) | (~w20491 & w26400) | (w20490 & w26400);
assign w20494 = ~w20492 & ~w20493;
assign w20495 = b_50 & w5196;
assign w20496 = w5459 & w31743;
assign w20497 = b_49 & w5191;
assign w20498 = ~w20496 & ~w20497;
assign w20499 = ~w20495 & w20498;
assign w20500 = (w20499 & ~w8162) | (w20499 & w26401) | (~w8162 & w26401);
assign w20501 = (w8162 & w31744) | (w8162 & w31745) | (w31744 & w31745);
assign w20502 = (~w8162 & w31746) | (~w8162 & w31747) | (w31746 & w31747);
assign w20503 = ~w20500 & ~w20501;
assign w20504 = ~w20502 & ~w20503;
assign w20505 = (w20504 & w20493) | (w20504 & w31748) | (w20493 & w31748);
assign w20506 = ~w20493 & w31749;
assign w20507 = ~w20505 & ~w20506;
assign w20508 = ~w20371 & w20507;
assign w20509 = ~w20371 & ~w20508;
assign w20510 = w20507 & ~w20508;
assign w20511 = ~w20509 & ~w20510;
assign w20512 = ~w20370 & ~w20511;
assign w20513 = (w20370 & w20508) | (w20370 & w31750) | (w20508 & w31750);
assign w20514 = ~w20509 & w20513;
assign w20515 = ~w20512 & ~w20514;
assign w20516 = ~w20360 & w20515;
assign w20517 = w20360 & ~w20515;
assign w20518 = ~w20516 & ~w20517;
assign w20519 = ~w20359 & w20518;
assign w20520 = ~w20518 & ~w20359;
assign w20521 = w20518 & ~w20519;
assign w20522 = ~w20520 & ~w20521;
assign w20523 = w20349 & ~w20522;
assign w20524 = w20349 & ~w20523;
assign w20525 = ~w20349 & ~w20522;
assign w20526 = ~w20524 & ~w20525;
assign w20527 = ~w20334 & w20526;
assign w20528 = w20334 & ~w20526;
assign w20529 = ~w20527 & ~w20528;
assign w20530 = (w20529 & w20320) | (w20529 & w31751) | (w20320 & w31751);
assign w20531 = ~w20320 & w31752;
assign w20532 = ~w20530 & ~w20531;
assign w20533 = (w20532 & w20301) | (w20532 & w41651) | (w20301 & w41651);
assign w20534 = ~w20301 & w41652;
assign w20535 = ~w20533 & ~w20534;
assign w20536 = (w14835 & w31753) | (w14835 & w31754) | (w31753 & w31754);
assign w20537 = (w13761 & w37708) | (w13761 & w37709) | (w37708 & w37709);
assign w20538 = ~w20536 & ~w20537;
assign w20539 = ~w20333 & ~w20528;
assign w20540 = b_63 & w2639;
assign w20541 = w2820 & w31755;
assign w20542 = b_62 & w2634;
assign w20543 = ~w20541 & ~w20542;
assign w20544 = ~w20540 & w20543;
assign w20545 = (w20544 & ~w12646) | (w20544 & w31756) | (~w12646 & w31756);
assign w20546 = (w12646 & w41653) | (w12646 & w41654) | (w41653 & w41654);
assign w20547 = (~w12646 & w41655) | (~w12646 & w41656) | (w41655 & w41656);
assign w20548 = ~w20545 & ~w20546;
assign w20549 = ~w20547 & ~w20548;
assign w20550 = (~w20549 & w20528) | (~w20549 & w31757) | (w20528 & w31757);
assign w20551 = ~w20539 & ~w20550;
assign w20552 = ~w20528 & w31758;
assign w20553 = b_57 & w3803;
assign w20554 = w4027 & w31759;
assign w20555 = b_56 & w3798;
assign w20556 = ~w20554 & ~w20555;
assign w20557 = ~w20553 & w20556;
assign w20558 = (w20557 & ~w10452) | (w20557 & w31760) | (~w10452 & w31760);
assign w20559 = (w10452 & w41657) | (w10452 & w41658) | (w41657 & w41658);
assign w20560 = (~w10452 & w41659) | (~w10452 & w41660) | (w41659 & w41660);
assign w20561 = ~w20558 & ~w20559;
assign w20562 = ~w20560 & ~w20561;
assign w20563 = (~w20508 & w20511) | (~w20508 & w31761) | (w20511 & w31761);
assign w20564 = (~w20493 & ~w20494) | (~w20493 & w26702) | (~w20494 & w26702);
assign w20565 = (~w20470 & ~w20472) | (~w20470 & w31762) | (~w20472 & w31762);
assign w20566 = (~w20453 & w20456) | (~w20453 & w31763) | (w20456 & w31763);
assign w20567 = b_33 & w10562;
assign w20568 = w10902 & w31764;
assign w20569 = b_32 & w10557;
assign w20570 = ~w20568 & ~w20569;
assign w20571 = ~w20567 & w20570;
assign w20572 = (w20571 & ~w3744) | (w20571 & w31765) | (~w3744 & w31765);
assign w20573 = (w3744 & w41661) | (w3744 & w41662) | (w41661 & w41662);
assign w20574 = (~w3744 & w41663) | (~w3744 & w41664) | (w41663 & w41664);
assign w20575 = ~w20572 & ~w20573;
assign w20576 = ~w20574 & ~w20575;
assign w20577 = (~w20423 & ~w20425) | (~w20423 & w31766) | (~w20425 & w31766);
assign w20578 = w20576 & w20577;
assign w20579 = ~w20576 & ~w20577;
assign w20580 = ~w20578 & ~w20579;
assign w20581 = w12380 & w31767;
assign w20582 = b_27 & ~w12380;
assign w20583 = ~w20581 & ~w20582;
assign w20584 = ~a_26 & ~w20583;
assign w20585 = a_26 & w20583;
assign w20586 = ~w20584 & ~w20585;
assign w20587 = ~w20409 & w20586;
assign w20588 = w20409 & ~w20586;
assign w20589 = ~w20587 & ~w20588;
assign w20590 = (w20589 & w20420) | (w20589 & w31768) | (w20420 & w31768);
assign w20591 = ~w20420 & w31769;
assign w20592 = ~w20590 & ~w20591;
assign w20593 = b_30 & w11620;
assign w20594 = w11969 & w31770;
assign w20595 = b_29 & w11615;
assign w20596 = ~w20594 & ~w20595;
assign w20597 = ~w20593 & w20596;
assign w20598 = (w20597 & ~w3138) | (w20597 & w31771) | (~w3138 & w31771);
assign w20599 = (w3138 & w41665) | (w3138 & w41666) | (w41665 & w41666);
assign w20600 = (~w3138 & w41667) | (~w3138 & w41668) | (w41667 & w41668);
assign w20601 = ~w20598 & ~w20599;
assign w20602 = ~w20600 & ~w20601;
assign w20603 = w20592 & ~w20602;
assign w20604 = w20592 & ~w20603;
assign w20605 = ~w20592 & ~w20602;
assign w20606 = ~w20604 & ~w20605;
assign w20607 = ~w20580 & w20606;
assign w20608 = w20580 & ~w20606;
assign w20609 = ~w20607 & ~w20608;
assign w20610 = b_36 & w9534;
assign w20611 = w9876 & w31772;
assign w20612 = b_35 & w9529;
assign w20613 = ~w20611 & ~w20612;
assign w20614 = ~w20610 & w20613;
assign w20615 = (w20614 & ~w4395) | (w20614 & w31773) | (~w4395 & w31773);
assign w20616 = (w4395 & w41669) | (w4395 & w41670) | (w41669 & w41670);
assign w20617 = (~w4395 & w41671) | (~w4395 & w41672) | (w41671 & w41672);
assign w20618 = ~w20615 & ~w20616;
assign w20619 = ~w20617 & ~w20618;
assign w20620 = w20609 & ~w20619;
assign w20621 = w20609 & ~w20620;
assign w20622 = ~w20609 & ~w20619;
assign w20623 = (~w20429 & ~w20431) | (~w20429 & w31774) | (~w20431 & w31774);
assign w20624 = ~w20621 & w31775;
assign w20625 = (~w20623 & w20621) | (~w20623 & w31776) | (w20621 & w31776);
assign w20626 = ~w20624 & ~w20625;
assign w20627 = b_39 & w8526;
assign w20628 = w8886 & w31777;
assign w20629 = b_38 & w8521;
assign w20630 = ~w20628 & ~w20629;
assign w20631 = ~w20627 & w20630;
assign w20632 = (w20631 & ~w4888) | (w20631 & w31778) | (~w4888 & w31778);
assign w20633 = (w4888 & w41673) | (w4888 & w41674) | (w41673 & w41674);
assign w20634 = (~w4888 & w41675) | (~w4888 & w41676) | (w41675 & w41676);
assign w20635 = ~w20632 & ~w20633;
assign w20636 = ~w20634 & ~w20635;
assign w20637 = w20626 & ~w20636;
assign w20638 = w20626 & ~w20637;
assign w20639 = ~w20626 & ~w20636;
assign w20640 = (~w20435 & ~w20437) | (~w20435 & w31779) | (~w20437 & w31779);
assign w20641 = ~w20638 & w31780;
assign w20642 = (~w20640 & w20638) | (~w20640 & w31781) | (w20638 & w31781);
assign w20643 = ~w20641 & ~w20642;
assign w20644 = b_42 & w7613;
assign w20645 = w7941 & w31782;
assign w20646 = b_41 & w7608;
assign w20647 = ~w20645 & ~w20646;
assign w20648 = ~w20644 & w20647;
assign w20649 = (w20648 & ~w5864) | (w20648 & w26402) | (~w5864 & w26402);
assign w20650 = (w5864 & w31783) | (w5864 & w31784) | (w31783 & w31784);
assign w20651 = (~w5864 & w31785) | (~w5864 & w31786) | (w31785 & w31786);
assign w20652 = ~w20649 & ~w20650;
assign w20653 = ~w20651 & ~w20652;
assign w20654 = w20643 & ~w20653;
assign w20655 = w20643 & ~w20654;
assign w20656 = ~w20643 & ~w20653;
assign w20657 = ~w20655 & ~w20656;
assign w20658 = ~w20566 & w20657;
assign w20659 = w20566 & ~w20657;
assign w20660 = ~w20658 & ~w20659;
assign w20661 = b_45 & w6761;
assign w20662 = w7075 & w31787;
assign w20663 = b_44 & w6756;
assign w20664 = ~w20662 & ~w20663;
assign w20665 = ~w20661 & w20664;
assign w20666 = (w20665 & ~w6682) | (w20665 & w26006) | (~w6682 & w26006);
assign w20667 = (w6682 & w26403) | (w6682 & w26404) | (w26403 & w26404);
assign w20668 = (~w6682 & w31788) | (~w6682 & w31789) | (w31788 & w31789);
assign w20669 = ~w20666 & ~w20667;
assign w20670 = ~w20668 & ~w20669;
assign w20671 = ~w20660 & ~w20670;
assign w20672 = w20660 & w20670;
assign w20673 = ~w20671 & ~w20672;
assign w20674 = w20565 & ~w20673;
assign w20675 = ~w20565 & w20673;
assign w20676 = ~w20674 & ~w20675;
assign w20677 = b_48 & w5962;
assign w20678 = w6246 & w31790;
assign w20679 = b_47 & w5957;
assign w20680 = ~w20678 & ~w20679;
assign w20681 = ~w20677 & w20680;
assign w20682 = (w20681 & ~w7284) | (w20681 & w25677) | (~w7284 & w25677);
assign w20683 = (w7284 & w26007) | (w7284 & w26008) | (w26007 & w26008);
assign w20684 = (~w7284 & w26405) | (~w7284 & w26406) | (w26405 & w26406);
assign w20685 = ~w20682 & ~w20683;
assign w20686 = ~w20684 & ~w20685;
assign w20687 = w20676 & ~w20686;
assign w20688 = w20686 & w20676;
assign w20689 = ~w20676 & ~w20686;
assign w20690 = (~w20476 & ~w20478) | (~w20476 & w31791) | (~w20478 & w31791);
assign w20691 = w20690 & w31792;
assign w20692 = (~w20690 & w20689) | (~w20690 & w26407) | (w20689 & w26407);
assign w20693 = b_51 & w5196;
assign w20694 = w5459 & w31793;
assign w20695 = b_50 & w5191;
assign w20696 = ~w20694 & ~w20695;
assign w20697 = ~w20693 & w20696;
assign w20698 = (w20697 & ~w8186) | (w20697 & w26009) | (~w8186 & w26009);
assign w20699 = (w8186 & w26408) | (w8186 & w26409) | (w26408 & w26409);
assign w20700 = (~w8186 & w31794) | (~w8186 & w31795) | (w31794 & w31795);
assign w20701 = ~w20698 & ~w20699;
assign w20702 = ~w20700 & ~w20701;
assign w20703 = ~w20692 & w31796;
assign w20704 = (w20702 & w20692) | (w20702 & w31797) | (w20692 & w31797);
assign w20705 = ~w20564 & ~w20704;
assign w20706 = (~w20564 & ~w20705) | (~w20564 & w27642) | (~w20705 & w27642);
assign w20707 = (~w20703 & w20564) | (~w20703 & w31798) | (w20564 & w31798);
assign w20708 = b_54 & w4499;
assign w20709 = w4723 & w31799;
assign w20710 = b_53 & w4494;
assign w20711 = ~w20709 & ~w20710;
assign w20712 = ~w20708 & w20711;
assign w20713 = (w20712 & ~w9134) | (w20712 & w31800) | (~w9134 & w31800);
assign w20714 = (w9134 & w41677) | (w9134 & w41678) | (w41677 & w41678);
assign w20715 = (~w9134 & w41679) | (~w9134 & w41680) | (w41679 & w41680);
assign w20716 = ~w20713 & ~w20714;
assign w20717 = ~w20715 & ~w20716;
assign w20718 = ~w20706 & w31801;
assign w20719 = (~w20717 & w20706) | (~w20717 & w31802) | (w20706 & w31802);
assign w20720 = ~w20718 & ~w20719;
assign w20721 = ~w20563 & w20720;
assign w20722 = w20563 & ~w20720;
assign w20723 = ~w20721 & ~w20722;
assign w20724 = ~w20562 & w20723;
assign w20725 = w20723 & ~w20724;
assign w20726 = ~w20723 & ~w20562;
assign w20727 = ~w20725 & ~w20726;
assign w20728 = (~w20516 & ~w20518) | (~w20516 & w31803) | (~w20518 & w31803);
assign w20729 = w20727 & w20728;
assign w20730 = ~w20727 & ~w20728;
assign w20731 = ~w20729 & ~w20730;
assign w20732 = b_60 & w3195;
assign w20733 = w3388 & w31804;
assign w20734 = b_59 & w3190;
assign w20735 = ~w20733 & ~w20734;
assign w20736 = ~w20732 & w20735;
assign w20737 = (w20736 & ~w11196) | (w20736 & w31805) | (~w11196 & w31805);
assign w20738 = (w11196 & w41681) | (w11196 & w41682) | (w41681 & w41682);
assign w20739 = (~w11196 & w41683) | (~w11196 & w41684) | (w41683 & w41684);
assign w20740 = ~w20737 & ~w20738;
assign w20741 = ~w20739 & ~w20740;
assign w20742 = (~w20348 & ~w20349) | (~w20348 & w31806) | (~w20349 & w31806);
assign w20743 = w20741 & w20742;
assign w20744 = ~w20741 & ~w20742;
assign w20745 = ~w20743 & ~w20744;
assign w20746 = w20731 & ~w20745;
assign w20747 = ~w20731 & w20745;
assign w20748 = ~w20746 & ~w20747;
assign w20749 = (~w20748 & w20551) | (~w20748 & w31807) | (w20551 & w31807);
assign w20750 = ~w20551 & w31808;
assign w20751 = ~w20749 & ~w20750;
assign w20752 = ~w20530 & w31809;
assign w20753 = (w20751 & w20530) | (w20751 & w31810) | (w20530 & w31810);
assign w20754 = ~w20752 & ~w20753;
assign w20755 = (~w13761 & w37642) | (~w13761 & w37643) | (w37642 & w37643);
assign w20756 = (w13761 & w37710) | (w13761 & w37711) | (w37710 & w37711);
assign w20757 = ~w20755 & ~w20756;
assign w20758 = (~w20744 & ~w20745) | (~w20744 & w31815) | (~w20745 & w31815);
assign w20759 = w2820 & w41685;
assign w20760 = b_63 & w2634;
assign w20761 = ~w20759 & ~w20760;
assign w20762 = ~w20759 & w31816;
assign w20763 = ~w12671 & w31817;
assign w20764 = (a_29 & w20763) | (a_29 & w31818) | (w20763 & w31818);
assign w20765 = ~w20763 & w31819;
assign w20766 = ~w20764 & ~w20765;
assign w20767 = (w20745 & w41686) | (w20745 & w41687) | (w41686 & w41687);
assign w20768 = (~w20745 & w41688) | (~w20745 & w41689) | (w41688 & w41689);
assign w20769 = ~w20767 & ~w20768;
assign w20770 = b_61 & w3195;
assign w20771 = w3388 & w31820;
assign w20772 = b_60 & w3190;
assign w20773 = ~w20771 & ~w20772;
assign w20774 = ~w20770 & w20773;
assign w20775 = (w20774 & ~w11901) | (w20774 & w31821) | (~w11901 & w31821);
assign w20776 = (w11901 & w41690) | (w11901 & w41691) | (w41690 & w41691);
assign w20777 = (~w11901 & w41692) | (~w11901 & w41693) | (w41692 & w41693);
assign w20778 = ~w20775 & ~w20776;
assign w20779 = ~w20777 & ~w20778;
assign w20780 = (~w20724 & w20727) | (~w20724 & w31822) | (w20727 & w31822);
assign w20781 = w20779 & w20780;
assign w20782 = ~w20779 & ~w20780;
assign w20783 = ~w20781 & ~w20782;
assign w20784 = b_58 & w3803;
assign w20785 = w4027 & w31823;
assign w20786 = b_57 & w3798;
assign w20787 = ~w20785 & ~w20786;
assign w20788 = ~w20784 & w20787;
assign w20789 = (w20788 & ~w10476) | (w20788 & w31824) | (~w10476 & w31824);
assign w20790 = (w10476 & w41694) | (w10476 & w41695) | (w41694 & w41695);
assign w20791 = (~w10476 & w41696) | (~w10476 & w41697) | (w41696 & w41697);
assign w20792 = ~w20789 & ~w20790;
assign w20793 = ~w20791 & ~w20792;
assign w20794 = ~w20719 & ~w20721;
assign w20795 = b_43 & w7613;
assign w20796 = w7941 & w31825;
assign w20797 = b_42 & w7608;
assign w20798 = ~w20796 & ~w20797;
assign w20799 = ~w20795 & w20798;
assign w20800 = (w20799 & ~w5888) | (w20799 & w27644) | (~w5888 & w27644);
assign w20801 = (w5888 & w31826) | (w5888 & w31827) | (w31826 & w31827);
assign w20802 = (~w5888 & w31828) | (~w5888 & w31829) | (w31828 & w31829);
assign w20803 = ~w20800 & ~w20801;
assign w20804 = ~w20802 & ~w20803;
assign w20805 = (~w31781 & w41698) | (~w31781 & w41699) | (w41698 & w41699);
assign w20806 = b_40 & w8526;
assign w20807 = w8886 & w31830;
assign w20808 = b_39 & w8521;
assign w20809 = ~w20807 & ~w20808;
assign w20810 = ~w20806 & w20809;
assign w20811 = (w20810 & ~w5363) | (w20810 & w31831) | (~w5363 & w31831);
assign w20812 = (w5363 & w41700) | (w5363 & w41701) | (w41700 & w41701);
assign w20813 = (~w5363 & w41702) | (~w5363 & w41703) | (w41702 & w41703);
assign w20814 = ~w20811 & ~w20812;
assign w20815 = ~w20813 & ~w20814;
assign w20816 = ~w20620 & ~w20625;
assign w20817 = b_34 & w10562;
assign w20818 = w10902 & w31832;
assign w20819 = b_33 & w10557;
assign w20820 = ~w20818 & ~w20819;
assign w20821 = ~w20817 & w20820;
assign w20822 = (w20821 & ~w3967) | (w20821 & w31833) | (~w3967 & w31833);
assign w20823 = (w3967 & w41704) | (w3967 & w41705) | (w41704 & w41705);
assign w20824 = (~w3967 & w41706) | (~w3967 & w41707) | (w41706 & w41707);
assign w20825 = ~w20822 & ~w20823;
assign w20826 = ~w20824 & ~w20825;
assign w20827 = w12380 & w31834;
assign w20828 = b_28 & ~w12380;
assign w20829 = ~w20827 & ~w20828;
assign w20830 = (~w20584 & ~w20586) | (~w20584 & w31835) | (~w20586 & w31835);
assign w20831 = ~w20829 & w20830;
assign w20832 = w20829 & ~w20830;
assign w20833 = ~w20831 & ~w20832;
assign w20834 = b_31 & w11620;
assign w20835 = w11969 & w31836;
assign w20836 = b_30 & w11615;
assign w20837 = ~w20835 & ~w20836;
assign w20838 = ~w20834 & w20837;
assign w20839 = (w20838 & ~w3345) | (w20838 & w26703) | (~w3345 & w26703);
assign w20840 = (w3345 & w31837) | (w3345 & w31838) | (w31837 & w31838);
assign w20841 = ~w20839 & ~w20840;
assign w20842 = ~w20841 & w31841;
assign w20843 = (w20833 & w20841) | (w20833 & w31842) | (w20841 & w31842);
assign w20844 = ~w20842 & ~w20843;
assign w20845 = (~w20590 & ~w20592) | (~w20590 & w31843) | (~w20592 & w31843);
assign w20846 = w20844 & ~w20845;
assign w20847 = ~w20844 & w20845;
assign w20848 = ~w20846 & ~w20847;
assign w20849 = ~w20826 & w20848;
assign w20850 = w20848 & ~w20849;
assign w20851 = ~w20848 & ~w20826;
assign w20852 = ~w20850 & ~w20851;
assign w20853 = (~w20579 & ~w20580) | (~w20579 & w31844) | (~w20580 & w31844);
assign w20854 = ~w20852 & ~w20853;
assign w20855 = ~w20852 & ~w20854;
assign w20856 = w20852 & ~w20853;
assign w20857 = b_37 & w9534;
assign w20858 = w9876 & w31845;
assign w20859 = b_36 & w9529;
assign w20860 = ~w20858 & ~w20859;
assign w20861 = ~w20857 & w20860;
assign w20862 = (w20861 & ~w4636) | (w20861 & w31846) | (~w4636 & w31846);
assign w20863 = (w4636 & w41708) | (w4636 & w41709) | (w41708 & w41709);
assign w20864 = (~w4636 & w41710) | (~w4636 & w41711) | (w41710 & w41711);
assign w20865 = ~w20862 & ~w20863;
assign w20866 = ~w20864 & ~w20865;
assign w20867 = (w20866 & w20855) | (w20866 & w31847) | (w20855 & w31847);
assign w20868 = ~w20855 & w31848;
assign w20869 = ~w20867 & ~w20868;
assign w20870 = ~w20816 & ~w20869;
assign w20871 = ~w20816 & ~w20870;
assign w20872 = ~w20869 & ~w20870;
assign w20873 = ~w20871 & ~w20872;
assign w20874 = ~w20815 & ~w20873;
assign w20875 = (w20815 & w20870) | (w20815 & w31849) | (w20870 & w31849);
assign w20876 = ~w20871 & w20875;
assign w20877 = ~w20874 & ~w20876;
assign w20878 = ~w20805 & w20877;
assign w20879 = w20805 & ~w20877;
assign w20880 = ~w20878 & ~w20879;
assign w20881 = ~w20804 & w20880;
assign w20882 = w20880 & ~w20881;
assign w20883 = ~w20880 & ~w20804;
assign w20884 = ~w20882 & ~w20883;
assign w20885 = ~w20566 & ~w20657;
assign w20886 = ~w20654 & ~w20885;
assign w20887 = w20884 & w20886;
assign w20888 = ~w20884 & ~w20886;
assign w20889 = ~w20887 & ~w20888;
assign w20890 = b_46 & w6761;
assign w20891 = w7075 & w31850;
assign w20892 = b_45 & w6756;
assign w20893 = ~w20891 & ~w20892;
assign w20894 = ~w20890 & w20893;
assign w20895 = (w20894 & ~w6974) | (w20894 & w26704) | (~w6974 & w26704);
assign w20896 = (w6974 & w27645) | (w6974 & w27646) | (w27645 & w27646);
assign w20897 = (~w6974 & w31851) | (~w6974 & w31852) | (w31851 & w31852);
assign w20898 = ~w20895 & ~w20896;
assign w20899 = ~w20897 & ~w20898;
assign w20900 = w20889 & ~w20899;
assign w20901 = w20889 & ~w20900;
assign w20902 = ~w20889 & ~w20899;
assign w20903 = ~w20671 & ~w20675;
assign w20904 = ~w20901 & w31853;
assign w20905 = (~w20903 & w20901) | (~w20903 & w31854) | (w20901 & w31854);
assign w20906 = ~w20904 & ~w20905;
assign w20907 = b_49 & w5962;
assign w20908 = w6246 & w31855;
assign w20909 = b_48 & w5957;
assign w20910 = ~w20908 & ~w20909;
assign w20911 = ~w20907 & w20910;
assign w20912 = (w20911 & ~w7859) | (w20911 & w27647) | (~w7859 & w27647);
assign w20913 = (w7859 & w31856) | (w7859 & w31857) | (w31856 & w31857);
assign w20914 = (~w7859 & w31858) | (~w7859 & w31859) | (w31858 & w31859);
assign w20915 = ~w20912 & ~w20913;
assign w20916 = ~w20914 & ~w20915;
assign w20917 = w20906 & ~w20916;
assign w20918 = w20906 & ~w20917;
assign w20919 = ~w20906 & ~w20916;
assign w20920 = (~w26407 & w31860) | (~w26407 & w31861) | (w31860 & w31861);
assign w20921 = ~w20918 & w31862;
assign w20922 = (~w20920 & w20918) | (~w20920 & w31863) | (w20918 & w31863);
assign w20923 = ~w20921 & ~w20922;
assign w20924 = b_52 & w5196;
assign w20925 = w5459 & w31864;
assign w20926 = b_51 & w5191;
assign w20927 = ~w20925 & ~w20926;
assign w20928 = ~w20924 & w20927;
assign w20929 = (w20928 & ~w8793) | (w20928 & w31865) | (~w8793 & w31865);
assign w20930 = (w8793 & w41712) | (w8793 & w41713) | (w41712 & w41713);
assign w20931 = (~w8793 & w41714) | (~w8793 & w41715) | (w41714 & w41715);
assign w20932 = ~w20929 & ~w20930;
assign w20933 = ~w20931 & ~w20932;
assign w20934 = w20923 & ~w20933;
assign w20935 = w20923 & ~w20934;
assign w20936 = ~w20923 & ~w20933;
assign w20937 = ~w20935 & ~w20936;
assign w20938 = ~w20707 & w20937;
assign w20939 = w20707 & ~w20937;
assign w20940 = ~w20938 & ~w20939;
assign w20941 = b_55 & w4499;
assign w20942 = w4723 & w31866;
assign w20943 = b_54 & w4494;
assign w20944 = ~w20942 & ~w20943;
assign w20945 = ~w20941 & w20944;
assign w20946 = (w20945 & ~w9776) | (w20945 & w31867) | (~w9776 & w31867);
assign w20947 = (w9776 & w41716) | (w9776 & w41717) | (w41716 & w41717);
assign w20948 = (~w9776 & w41718) | (~w9776 & w41719) | (w41718 & w41719);
assign w20949 = ~w20946 & ~w20947;
assign w20950 = ~w20948 & ~w20949;
assign w20951 = ~w20940 & ~w20950;
assign w20952 = w20940 & w20950;
assign w20953 = ~w20951 & ~w20952;
assign w20954 = ~w20794 & w20953;
assign w20955 = w20794 & ~w20953;
assign w20956 = ~w20954 & ~w20955;
assign w20957 = ~w20793 & w20956;
assign w20958 = w20956 & ~w20957;
assign w20959 = ~w20956 & ~w20793;
assign w20960 = ~w20958 & ~w20959;
assign w20961 = w20783 & ~w20960;
assign w20962 = ~w20783 & w20960;
assign w20963 = w20769 & w31868;
assign w20964 = w20769 & ~w20963;
assign w20965 = w31868 & ~w20769;
assign w20966 = ~w20964 & ~w20965;
assign w20967 = ~w20550 & ~w20749;
assign w20968 = w20966 & w20967;
assign w20969 = ~w20966 & ~w20967;
assign w20970 = ~w20968 & ~w20969;
assign w20971 = (~w13761 & w37712) | (~w13761 & w37713) | (w37712 & w37713);
assign w20972 = (w13761 & w37714) | (w13761 & w37715) | (w37714 & w37715);
assign w20973 = ~w20971 & ~w20972;
assign w20974 = (~w20767 & ~w20769) | (~w20767 & w31871) | (~w20769 & w31871);
assign w20975 = (~w20782 & ~w20783) | (~w20782 & w31872) | (~w20783 & w31872);
assign w20976 = w2820 & w31873;
assign w20977 = (w6406 & w41720) | (w6406 & w41721) | (w41720 & w41721);
assign w20978 = ~w20976 & ~w20977;
assign w20979 = (a_29 & w20977) | (a_29 & w31876) | (w20977 & w31876);
assign w20980 = ~w20977 & w31877;
assign w20981 = ~w20978 & ~w20979;
assign w20982 = ~w20980 & ~w20981;
assign w20983 = ~w20975 & ~w20982;
assign w20984 = ~w20975 & ~w20983;
assign w20985 = w20975 & ~w20982;
assign w20986 = b_62 & w3195;
assign w20987 = w3388 & w31878;
assign w20988 = b_61 & w3190;
assign w20989 = ~w20987 & ~w20988;
assign w20990 = ~w20986 & w20989;
assign w20991 = (w20990 & ~w12273) | (w20990 & w31879) | (~w12273 & w31879);
assign w20992 = (w12273 & w41722) | (w12273 & w41723) | (w41722 & w41723);
assign w20993 = (~w12273 & w41724) | (~w12273 & w41725) | (w41724 & w41725);
assign w20994 = ~w20991 & ~w20992;
assign w20995 = ~w20993 & ~w20994;
assign w20996 = (~w20954 & ~w20956) | (~w20954 & w31880) | (~w20956 & w31880);
assign w20997 = w20995 & w20996;
assign w20998 = ~w20995 & ~w20996;
assign w20999 = ~w20997 & ~w20998;
assign w21000 = ~w20707 & ~w20937;
assign w21001 = (~w21000 & w20940) | (~w21000 & w31881) | (w20940 & w31881);
assign w21002 = b_56 & w4499;
assign w21003 = w4723 & w31882;
assign w21004 = b_55 & w4494;
assign w21005 = ~w21003 & ~w21004;
assign w21006 = ~w21002 & w21005;
assign w21007 = (w21006 & ~w9798) | (w21006 & w31883) | (~w9798 & w31883);
assign w21008 = (w9798 & w41726) | (w9798 & w41727) | (w41726 & w41727);
assign w21009 = (~w9798 & w41728) | (~w9798 & w41729) | (w41728 & w41729);
assign w21010 = ~w21007 & ~w21008;
assign w21011 = ~w21009 & ~w21010;
assign w21012 = (~w20922 & ~w20923) | (~w20922 & w31884) | (~w20923 & w31884);
assign w21013 = b_53 & w5196;
assign w21014 = w5459 & w31885;
assign w21015 = b_52 & w5191;
assign w21016 = ~w21014 & ~w21015;
assign w21017 = ~w21013 & w21016;
assign w21018 = (w9109 & w41730) | (w9109 & w41731) | (w41730 & w41731);
assign w21019 = a_41 & ~w21018;
assign w21020 = w21018 & a_41;
assign w21021 = ~w21018 & ~w21019;
assign w21022 = ~w21020 & ~w21021;
assign w21023 = (~w20905 & ~w20906) | (~w20905 & w31887) | (~w20906 & w31887);
assign w21024 = (~w20878 & ~w20880) | (~w20878 & w31888) | (~w20880 & w31888);
assign w21025 = b_44 & w7613;
assign w21026 = w7941 & w31889;
assign w21027 = b_43 & w7608;
assign w21028 = ~w21026 & ~w21027;
assign w21029 = ~w21025 & w21028;
assign w21030 = (w21029 & ~w6408) | (w21029 & w26410) | (~w6408 & w26410);
assign w21031 = (w6408 & w31890) | (w6408 & w31891) | (w31890 & w31891);
assign w21032 = (~w6408 & w31892) | (~w6408 & w31893) | (w31892 & w31893);
assign w21033 = ~w21030 & ~w21031;
assign w21034 = ~w21032 & ~w21033;
assign w21035 = (~w20870 & w20873) | (~w20870 & w31894) | (w20873 & w31894);
assign w21036 = (~w20846 & ~w20848) | (~w20846 & w31895) | (~w20848 & w31895);
assign w21037 = b_35 & w10562;
assign w21038 = w10902 & w31896;
assign w21039 = b_34 & w10557;
assign w21040 = ~w21038 & ~w21039;
assign w21041 = ~w21037 & w21040;
assign w21042 = (w21041 & ~w4181) | (w21041 & w31897) | (~w4181 & w31897);
assign w21043 = (w4181 & w41732) | (w4181 & w41733) | (w41732 & w41733);
assign w21044 = (~w4181 & w41734) | (~w4181 & w41735) | (w41734 & w41735);
assign w21045 = ~w21042 & ~w21043;
assign w21046 = ~w21044 & ~w21045;
assign w21047 = (~w20841 & w41736) | (~w20841 & w41737) | (w41736 & w41737);
assign w21048 = w12380 & w31898;
assign w21049 = b_29 & ~w12380;
assign w21050 = ~w21048 & ~w21049;
assign w21051 = w20829 & ~w21050;
assign w21052 = ~w20829 & w21050;
assign w21053 = (w20841 & w41738) | (w20841 & w41739) | (w41738 & w41739);
assign w21054 = ~w21047 & ~w21053;
assign w21055 = (~w20841 & w41740) | (~w20841 & w41741) | (w41740 & w41741);
assign w21056 = (~w20841 & w41742) | (~w20841 & w41743) | (w41742 & w41743);
assign w21057 = b_32 & w11620;
assign w21058 = w11969 & w31904;
assign w21059 = b_31 & w11615;
assign w21060 = ~w21058 & ~w21059;
assign w21061 = ~w21057 & w21060;
assign w21062 = (w21061 & ~w3545) | (w21061 & w31905) | (~w3545 & w31905);
assign w21063 = (w3545 & w41744) | (w3545 & w41745) | (w41744 & w41745);
assign w21064 = (~w3545 & w41746) | (~w3545 & w41747) | (w41746 & w41747);
assign w21065 = ~w21062 & ~w21063;
assign w21066 = ~w21064 & ~w21065;
assign w21067 = (w21066 & w21054) | (w21066 & w31906) | (w21054 & w31906);
assign w21068 = ~w21054 & w31907;
assign w21069 = ~w21067 & ~w21068;
assign w21070 = ~w21046 & ~w21069;
assign w21071 = w21046 & w21069;
assign w21072 = ~w21070 & ~w21071;
assign w21073 = ~w21036 & w21072;
assign w21074 = w21036 & ~w21072;
assign w21075 = ~w21073 & ~w21074;
assign w21076 = b_38 & w9534;
assign w21077 = w9876 & w31908;
assign w21078 = b_37 & w9529;
assign w21079 = ~w21077 & ~w21078;
assign w21080 = ~w21076 & w21079;
assign w21081 = (w21080 & ~w4658) | (w21080 & w31909) | (~w4658 & w31909);
assign w21082 = (w4658 & w41748) | (w4658 & w41749) | (w41748 & w41749);
assign w21083 = (~w4658 & w41750) | (~w4658 & w41751) | (w41750 & w41751);
assign w21084 = ~w21081 & ~w21082;
assign w21085 = ~w21083 & ~w21084;
assign w21086 = w21075 & ~w21085;
assign w21087 = w21075 & ~w21086;
assign w21088 = ~w21075 & ~w21085;
assign w21089 = ~w21087 & ~w21088;
assign w21090 = (~w20866 & w20855) | (~w20866 & w31910) | (w20855 & w31910);
assign w21091 = ~w20854 & ~w21090;
assign w21092 = ~w21089 & ~w21091;
assign w21093 = w21091 & ~w21089;
assign w21094 = ~w21091 & ~w21092;
assign w21095 = b_41 & w8526;
assign w21096 = w8886 & w31911;
assign w21097 = b_40 & w8521;
assign w21098 = ~w21096 & ~w21097;
assign w21099 = ~w21095 & w21098;
assign w21100 = (w21099 & ~w5609) | (w21099 & w31912) | (~w5609 & w31912);
assign w21101 = (w5609 & w41752) | (w5609 & w41753) | (w41752 & w41753);
assign w21102 = (~w5609 & w41754) | (~w5609 & w41755) | (w41754 & w41755);
assign w21103 = ~w21100 & ~w21101;
assign w21104 = ~w21102 & ~w21103;
assign w21105 = (w21104 & w21094) | (w21104 & w31913) | (w21094 & w31913);
assign w21106 = ~w21094 & w31914;
assign w21107 = ~w21105 & ~w21106;
assign w21108 = ~w21035 & ~w21107;
assign w21109 = w21035 & w21107;
assign w21110 = ~w21108 & ~w21109;
assign w21111 = ~w21034 & w21110;
assign w21112 = w21034 & ~w21110;
assign w21113 = ~w21111 & ~w21112;
assign w21114 = ~w21024 & w21113;
assign w21115 = w21024 & ~w21113;
assign w21116 = ~w21114 & ~w21115;
assign w21117 = b_47 & w6761;
assign w21118 = w7075 & w31915;
assign w21119 = b_46 & w6756;
assign w21120 = ~w21118 & ~w21119;
assign w21121 = ~w21117 & w21120;
assign w21122 = (w21121 & ~w6998) | (w21121 & w25678) | (~w6998 & w25678);
assign w21123 = (w6998 & w26010) | (w6998 & w26011) | (w26010 & w26011);
assign w21124 = (~w6998 & w26411) | (~w6998 & w26412) | (w26411 & w26412);
assign w21125 = ~w21122 & ~w21123;
assign w21126 = ~w21124 & ~w21125;
assign w21127 = w21126 & w21116;
assign w21128 = ~w21116 & ~w21126;
assign w21129 = (~w20888 & ~w20889) | (~w20888 & w41756) | (~w20889 & w41756);
assign w21130 = w21129 & w31916;
assign w21131 = (~w21129 & w21128) | (~w21129 & w26705) | (w21128 & w26705);
assign w21132 = ~w21130 & ~w21131;
assign w21133 = b_50 & w5962;
assign w21134 = w6246 & w31917;
assign w21135 = b_49 & w5957;
assign w21136 = ~w21134 & ~w21135;
assign w21137 = ~w21133 & w21136;
assign w21138 = (w21137 & ~w8162) | (w21137 & w26413) | (~w8162 & w26413);
assign w21139 = (w8162 & w31918) | (w8162 & w31919) | (w31918 & w31919);
assign w21140 = (~w8162 & w31920) | (~w8162 & w31921) | (w31920 & w31921);
assign w21141 = ~w21138 & ~w21139;
assign w21142 = ~w21140 & ~w21141;
assign w21143 = (w21142 & w21131) | (w21142 & w31922) | (w21131 & w31922);
assign w21144 = ~w21131 & w31923;
assign w21145 = ~w21143 & ~w21144;
assign w21146 = ~w21023 & w21145;
assign w21147 = w21023 & w21145;
assign w21148 = (~w21022 & w21147) | (~w21022 & w31924) | (w21147 & w31924);
assign w21149 = ~w21147 & w31925;
assign w21150 = ~w21148 & ~w21149;
assign w21151 = ~w21012 & w21150;
assign w21152 = w21012 & ~w21150;
assign w21153 = ~w21151 & ~w21152;
assign w21154 = ~w21011 & w21153;
assign w21155 = w21011 & ~w21153;
assign w21156 = ~w21154 & ~w21155;
assign w21157 = ~w21001 & w21156;
assign w21158 = w21001 & ~w21156;
assign w21159 = ~w21157 & ~w21158;
assign w21160 = b_59 & w3803;
assign w21161 = w4027 & w31926;
assign w21162 = b_58 & w3798;
assign w21163 = ~w21161 & ~w21162;
assign w21164 = ~w21160 & w21163;
assign w21165 = (w21164 & ~w11169) | (w21164 & w31927) | (~w11169 & w31927);
assign w21166 = (w11169 & w41757) | (w11169 & w41758) | (w41757 & w41758);
assign w21167 = (~w11169 & w41759) | (~w11169 & w41760) | (w41759 & w41760);
assign w21168 = ~w21165 & ~w21166;
assign w21169 = ~w21167 & ~w21168;
assign w21170 = w21159 & ~w21169;
assign w21171 = w21159 & ~w21170;
assign w21172 = ~w21159 & ~w21169;
assign w21173 = ~w21171 & ~w21172;
assign w21174 = ~w20999 & w21173;
assign w21175 = w20999 & ~w21173;
assign w21176 = ~w21174 & ~w21175;
assign w21177 = (w21176 & w20984) | (w21176 & w31928) | (w20984 & w31928);
assign w21178 = ~w20984 & w31929;
assign w21179 = ~w21177 & ~w21178;
assign w21180 = ~w20974 & w21179;
assign w21181 = ~w20974 & ~w21180;
assign w21182 = w20974 & w21179;
assign w21183 = ~w21181 & ~w21182;
assign w21184 = (~w13761 & w37716) | (~w13761 & w37717) | (w37716 & w37717);
assign w21185 = (w13761 & w37718) | (w13761 & w37719) | (w37718 & w37719);
assign w21186 = ~w21184 & ~w21185;
assign w21187 = ~w20983 & ~w21177;
assign w21188 = b_57 & w4499;
assign w21189 = w4723 & w31934;
assign w21190 = b_56 & w4494;
assign w21191 = ~w21189 & ~w21190;
assign w21192 = ~w21188 & w21191;
assign w21193 = (w21192 & ~w10452) | (w21192 & w31935) | (~w10452 & w31935);
assign w21194 = (w10452 & w41761) | (w10452 & w41762) | (w41761 & w41762);
assign w21195 = (~w10452 & w41763) | (~w10452 & w41764) | (w41763 & w41764);
assign w21196 = ~w21193 & ~w21194;
assign w21197 = ~w21195 & ~w21196;
assign w21198 = (~w31924 & w41765) | (~w31924 & w41766) | (w41765 & w41766);
assign w21199 = (~w21131 & ~w21132) | (~w21131 & w26414) | (~w21132 & w26414);
assign w21200 = (~w21108 & ~w21110) | (~w21108 & w31936) | (~w21110 & w31936);
assign w21201 = (~w21104 & w21094) | (~w21104 & w31937) | (w21094 & w31937);
assign w21202 = ~w21092 & ~w21201;
assign w21203 = b_39 & w9534;
assign w21204 = w9876 & w31938;
assign w21205 = b_38 & w9529;
assign w21206 = ~w21204 & ~w21205;
assign w21207 = ~w21203 & w21206;
assign w21208 = (w21207 & ~w4888) | (w21207 & w26706) | (~w4888 & w26706);
assign w21209 = (w4888 & w31939) | (w4888 & w31940) | (w31939 & w31940);
assign w21210 = (~w4888 & w31941) | (~w4888 & w31942) | (w31941 & w31942);
assign w21211 = ~w21208 & ~w21209;
assign w21212 = ~w21210 & ~w21211;
assign w21213 = (~w21066 & w21054) | (~w21066 & w31943) | (w21054 & w31943);
assign w21214 = (~w21213 & w21069) | (~w21213 & w41767) | (w21069 & w41767);
assign w21215 = w12380 & w31944;
assign w21216 = b_30 & ~w12380;
assign w21217 = ~w21215 & ~w21216;
assign w21218 = ~a_29 & ~w21217;
assign w21219 = a_29 & w21217;
assign w21220 = ~w21218 & ~w21219;
assign w21221 = ~w21050 & w21220;
assign w21222 = ~w21220 & ~w21050;
assign w21223 = w21220 & ~w21221;
assign w21224 = ~w21222 & ~w21223;
assign w21225 = (w20841 & w41768) | (w20841 & w41769) | (w41768 & w41769);
assign w21226 = ~w21055 & ~w21225;
assign w21227 = (~w20841 & w41770) | (~w20841 & w41771) | (w41770 & w41771);
assign w21228 = ~w21226 & ~w21227;
assign w21229 = b_33 & w11620;
assign w21230 = w11969 & w31949;
assign w21231 = b_32 & w11615;
assign w21232 = ~w21230 & ~w21231;
assign w21233 = ~w21229 & w21232;
assign w21234 = (w21233 & ~w3744) | (w21233 & w31950) | (~w3744 & w31950);
assign w21235 = (w3744 & w41772) | (w3744 & w41773) | (w41772 & w41773);
assign w21236 = (~w3744 & w41774) | (~w3744 & w41775) | (w41774 & w41775);
assign w21237 = ~w21234 & ~w21235;
assign w21238 = ~w21236 & ~w21237;
assign w21239 = (w21238 & w21226) | (w21238 & w41776) | (w21226 & w41776);
assign w21240 = ~w21226 & w41777;
assign w21241 = ~w21239 & ~w21240;
assign w21242 = b_36 & w10562;
assign w21243 = w10902 & w31951;
assign w21244 = b_35 & w10557;
assign w21245 = ~w21243 & ~w21244;
assign w21246 = ~w21242 & w21245;
assign w21247 = (w21246 & ~w4395) | (w21246 & w31952) | (~w4395 & w31952);
assign w21248 = (w4395 & w41778) | (w4395 & w41779) | (w41778 & w41779);
assign w21249 = (~w4395 & w41780) | (~w4395 & w41781) | (w41780 & w41781);
assign w21250 = ~w21247 & ~w21248;
assign w21251 = ~w21249 & ~w21250;
assign w21252 = ~w21241 & ~w21251;
assign w21253 = w21241 & w21251;
assign w21254 = ~w21252 & ~w21253;
assign w21255 = ~w21214 & w21254;
assign w21256 = w21214 & ~w21254;
assign w21257 = ~w21255 & ~w21256;
assign w21258 = ~w21212 & w21257;
assign w21259 = w21257 & ~w21258;
assign w21260 = ~w21257 & ~w21212;
assign w21261 = (~w21073 & ~w21075) | (~w21073 & w31953) | (~w21075 & w31953);
assign w21262 = ~w21259 & w31954;
assign w21263 = (~w21261 & w21259) | (~w21261 & w31955) | (w21259 & w31955);
assign w21264 = ~w21262 & ~w21263;
assign w21265 = b_42 & w8526;
assign w21266 = w8886 & w31956;
assign w21267 = b_41 & w8521;
assign w21268 = ~w21266 & ~w21267;
assign w21269 = ~w21265 & w21268;
assign w21270 = (w21269 & ~w5864) | (w21269 & w26415) | (~w5864 & w26415);
assign w21271 = (w5864 & w26707) | (w5864 & w26708) | (w26707 & w26708);
assign w21272 = (~w5864 & w31957) | (~w5864 & w31958) | (w31957 & w31958);
assign w21273 = ~w21270 & ~w21271;
assign w21274 = ~w21272 & ~w21273;
assign w21275 = w21264 & ~w21274;
assign w21276 = w21264 & ~w21275;
assign w21277 = ~w21264 & ~w21274;
assign w21278 = ~w21276 & ~w21277;
assign w21279 = ~w21202 & w21278;
assign w21280 = w21202 & ~w21278;
assign w21281 = ~w21279 & ~w21280;
assign w21282 = b_45 & w7613;
assign w21283 = w7941 & w31959;
assign w21284 = b_44 & w7608;
assign w21285 = ~w21283 & ~w21284;
assign w21286 = ~w21282 & w21285;
assign w21287 = (w21286 & ~w6682) | (w21286 & w26012) | (~w6682 & w26012);
assign w21288 = (w6682 & w26416) | (w6682 & w26417) | (w26416 & w26417);
assign w21289 = (~w6682 & w31960) | (~w6682 & w31961) | (w31960 & w31961);
assign w21290 = ~w21287 & ~w21288;
assign w21291 = ~w21289 & ~w21290;
assign w21292 = ~w21281 & ~w21291;
assign w21293 = w21281 & w21291;
assign w21294 = ~w21292 & ~w21293;
assign w21295 = w21200 & ~w21294;
assign w21296 = ~w21200 & w21294;
assign w21297 = ~w21295 & ~w21296;
assign w21298 = b_48 & w6761;
assign w21299 = w7075 & w31962;
assign w21300 = b_47 & w6756;
assign w21301 = ~w21299 & ~w21300;
assign w21302 = ~w21298 & w21301;
assign w21303 = (w21302 & ~w7284) | (w21302 & w25679) | (~w7284 & w25679);
assign w21304 = (w7284 & w26013) | (w7284 & w26014) | (w26013 & w26014);
assign w21305 = (~w7284 & w26418) | (~w7284 & w26419) | (w26418 & w26419);
assign w21306 = ~w21303 & ~w21304;
assign w21307 = ~w21305 & ~w21306;
assign w21308 = w21297 & ~w21307;
assign w21309 = w21307 & w21297;
assign w21310 = ~w21297 & ~w21307;
assign w21311 = (~w21114 & ~w21116) | (~w21114 & w31963) | (~w21116 & w31963);
assign w21312 = ~w21310 & w26420;
assign w21313 = (~w21311 & w21310) | (~w21311 & w26421) | (w21310 & w26421);
assign w21314 = ~w21312 & ~w21313;
assign w21315 = b_51 & w5962;
assign w21316 = w6246 & w31964;
assign w21317 = b_50 & w5957;
assign w21318 = ~w21316 & ~w21317;
assign w21319 = ~w21315 & w21318;
assign w21320 = (w21319 & ~w8186) | (w21319 & w26015) | (~w8186 & w26015);
assign w21321 = (w8186 & w26422) | (w8186 & w26423) | (w26422 & w26423);
assign w21322 = (~w8186 & w31965) | (~w8186 & w31966) | (w31965 & w31966);
assign w21323 = ~w21320 & ~w21321;
assign w21324 = ~w21322 & ~w21323;
assign w21325 = w21314 & ~w21324;
assign w21326 = ~w21314 & w21324;
assign w21327 = (w21132 & w41782) | (w21132 & w41783) | (w41782 & w41783);
assign w21328 = (~w21199 & ~w21327) | (~w21199 & w27648) | (~w21327 & w27648);
assign w21329 = (~w21325 & w21199) | (~w21325 & w31967) | (w21199 & w31967);
assign w21330 = (w27649 & w21199) | (w27649 & w31968) | (w21199 & w31968);
assign w21331 = b_54 & w5196;
assign w21332 = w5459 & w31969;
assign w21333 = b_53 & w5191;
assign w21334 = ~w21332 & ~w21333;
assign w21335 = ~w21331 & w21334;
assign w21336 = (w21335 & ~w9134) | (w21335 & w31970) | (~w9134 & w31970);
assign w21337 = (w9134 & w41784) | (w9134 & w41785) | (w41784 & w41785);
assign w21338 = (~w9134 & w41786) | (~w9134 & w41787) | (w41786 & w41787);
assign w21339 = ~w21336 & ~w21337;
assign w21340 = ~w21338 & ~w21339;
assign w21341 = ~w21328 & w31971;
assign w21342 = (~w21340 & w21328) | (~w21340 & w31972) | (w21328 & w31972);
assign w21343 = ~w21341 & ~w21342;
assign w21344 = ~w21198 & w21343;
assign w21345 = w21198 & ~w21343;
assign w21346 = ~w21344 & ~w21345;
assign w21347 = ~w21197 & w21346;
assign w21348 = w21346 & ~w21347;
assign w21349 = ~w21346 & ~w21197;
assign w21350 = (~w21151 & ~w21153) | (~w21151 & w31973) | (~w21153 & w31973);
assign w21351 = ~w21348 & w31974;
assign w21352 = (~w21350 & w21348) | (~w21350 & w31975) | (w21348 & w31975);
assign w21353 = ~w21351 & ~w21352;
assign w21354 = b_60 & w3803;
assign w21355 = w4027 & w31976;
assign w21356 = b_59 & w3798;
assign w21357 = ~w21355 & ~w21356;
assign w21358 = ~w21354 & w21357;
assign w21359 = (w21358 & ~w11196) | (w21358 & w31977) | (~w11196 & w31977);
assign w21360 = (w11196 & w41788) | (w11196 & w41789) | (w41788 & w41789);
assign w21361 = (~w11196 & w41790) | (~w11196 & w41791) | (w41790 & w41791);
assign w21362 = ~w21359 & ~w21360;
assign w21363 = ~w21361 & ~w21362;
assign w21364 = w21353 & ~w21363;
assign w21365 = w21353 & ~w21364;
assign w21366 = ~w21353 & ~w21363;
assign w21367 = (~w21157 & ~w21159) | (~w21157 & w31978) | (~w21159 & w31978);
assign w21368 = ~w21365 & w31979;
assign w21369 = (~w21367 & w21365) | (~w21367 & w31980) | (w21365 & w31980);
assign w21370 = ~w21368 & ~w21369;
assign w21371 = (~w20998 & ~w20999) | (~w20998 & w31981) | (~w20999 & w31981);
assign w21372 = b_63 & w3195;
assign w21373 = w3388 & w31982;
assign w21374 = b_62 & w3190;
assign w21375 = ~w21373 & ~w21374;
assign w21376 = ~w21372 & w21375;
assign w21377 = (w21376 & ~w12646) | (w21376 & w31983) | (~w12646 & w31983);
assign w21378 = (w12646 & w41792) | (w12646 & w41793) | (w41792 & w41793);
assign w21379 = (~w12646 & w41794) | (~w12646 & w41795) | (w41794 & w41795);
assign w21380 = ~w21377 & ~w21378;
assign w21381 = ~w21379 & ~w21380;
assign w21382 = ~w21371 & ~w21381;
assign w21383 = ~w21371 & ~w21382;
assign w21384 = ~w21383 & w31984;
assign w21385 = (w21370 & w21383) | (w21370 & w31985) | (w21383 & w31985);
assign w21386 = ~w21384 & ~w21385;
assign w21387 = ~w21187 & w21386;
assign w21388 = w21187 & ~w21386;
assign w21389 = ~w21387 & ~w21388;
assign w21390 = (~w13761 & w37720) | (~w13761 & w37721) | (w37720 & w37721);
assign w21391 = (w13761 & w37722) | (w13761 & w37723) | (w37722 & w37723);
assign w21392 = ~w21390 & ~w21391;
assign w21393 = w3388 & w31986;
assign w21394 = b_63 & w3190;
assign w21395 = ~w21393 & ~w21394;
assign w21396 = ~w12671 & w31987;
assign w21397 = (a_32 & w21396) | (a_32 & w31988) | (w21396 & w31988);
assign w21398 = ~w21396 & w31989;
assign w21399 = ~w21397 & ~w21398;
assign w21400 = (w31980 & w41796) | (w31980 & w41797) | (w41796 & w41797);
assign w21401 = (~w31980 & w41798) | (~w31980 & w41799) | (w41798 & w41799);
assign w21402 = ~w21400 & ~w21401;
assign w21403 = b_58 & w4499;
assign w21404 = w4723 & w31992;
assign w21405 = b_57 & w4494;
assign w21406 = ~w21404 & ~w21405;
assign w21407 = ~w21403 & w21406;
assign w21408 = (w21407 & ~w10476) | (w21407 & w31993) | (~w10476 & w31993);
assign w21409 = (w10476 & w41800) | (w10476 & w41801) | (w41800 & w41801);
assign w21410 = (~w10476 & w41802) | (~w10476 & w41803) | (w41802 & w41803);
assign w21411 = ~w21408 & ~w21409;
assign w21412 = ~w21410 & ~w21411;
assign w21413 = ~w21342 & ~w21344;
assign w21414 = b_43 & w8526;
assign w21415 = w8886 & w31994;
assign w21416 = b_42 & w8521;
assign w21417 = ~w21415 & ~w21416;
assign w21418 = ~w21414 & w21417;
assign w21419 = (w21418 & ~w5888) | (w21418 & w26424) | (~w5888 & w26424);
assign w21420 = (w5888 & w26709) | (w5888 & w26710) | (w26709 & w26710);
assign w21421 = (~w5888 & w31995) | (~w5888 & w31996) | (w31995 & w31996);
assign w21422 = ~w21419 & ~w21420;
assign w21423 = ~w21421 & ~w21422;
assign w21424 = ~w21258 & ~w21263;
assign w21425 = b_40 & w9534;
assign w21426 = w9876 & w31997;
assign w21427 = b_39 & w9529;
assign w21428 = ~w21426 & ~w21427;
assign w21429 = ~w21425 & w21428;
assign w21430 = (w21429 & ~w5363) | (w21429 & w26711) | (~w5363 & w26711);
assign w21431 = (w5363 & w31998) | (w5363 & w31999) | (w31998 & w31999);
assign w21432 = (~w5363 & w32000) | (~w5363 & w32001) | (w32000 & w32001);
assign w21433 = ~w21430 & ~w21431;
assign w21434 = ~w21432 & ~w21433;
assign w21435 = (~w21252 & ~w21254) | (~w21252 & w32002) | (~w21254 & w32002);
assign w21436 = b_37 & w10562;
assign w21437 = w10902 & w32003;
assign w21438 = b_36 & w10557;
assign w21439 = ~w21437 & ~w21438;
assign w21440 = ~w21436 & w21439;
assign w21441 = (w21440 & ~w4636) | (w21440 & w32004) | (~w4636 & w32004);
assign w21442 = (w4636 & w41804) | (w4636 & w41805) | (w41804 & w41805);
assign w21443 = (~w4636 & w41806) | (~w4636 & w41807) | (w41806 & w41807);
assign w21444 = ~w21441 & ~w21442;
assign w21445 = ~w21443 & ~w21444;
assign w21446 = (~w21225 & w21228) | (~w21225 & w32005) | (w21228 & w32005);
assign w21447 = w12380 & w41808;
assign w21448 = b_31 & ~w12380;
assign w21449 = ~w21447 & ~w21448;
assign w21450 = (~w21218 & ~w21220) | (~w21218 & w32006) | (~w21220 & w32006);
assign w21451 = ~w21449 & w21450;
assign w21452 = w21449 & ~w21450;
assign w21453 = ~w21451 & ~w21452;
assign w21454 = b_34 & w11620;
assign w21455 = w11969 & w32007;
assign w21456 = b_33 & w11615;
assign w21457 = ~w21455 & ~w21456;
assign w21458 = ~w21454 & w21457;
assign w21459 = (w21458 & ~w3967) | (w21458 & w26425) | (~w3967 & w26425);
assign w21460 = (w3967 & w32008) | (w3967 & w32009) | (w32008 & w32009);
assign w21461 = ~w21459 & ~w21460;
assign w21462 = ~w21461 & w32012;
assign w21463 = (w21453 & w21461) | (w21453 & w32013) | (w21461 & w32013);
assign w21464 = ~w21462 & ~w21463;
assign w21465 = (~w21228 & w41809) | (~w21228 & w41810) | (w41809 & w41810);
assign w21466 = ~w21446 & ~w21465;
assign w21467 = (w21228 & w41811) | (w21228 & w41812) | (w41811 & w41812);
assign w21468 = (~w21445 & w21466) | (~w21445 & w32014) | (w21466 & w32014);
assign w21469 = w21445 & ~w21467;
assign w21470 = ~w21466 & w21469;
assign w21471 = ~w21468 & ~w21470;
assign w21472 = ~w21435 & w21471;
assign w21473 = ~w21435 & ~w21472;
assign w21474 = w21471 & ~w21472;
assign w21475 = ~w21473 & ~w21474;
assign w21476 = ~w21434 & ~w21475;
assign w21477 = (w21434 & w21472) | (w21434 & w32015) | (w21472 & w32015);
assign w21478 = ~w21473 & w21477;
assign w21479 = ~w21476 & ~w21478;
assign w21480 = ~w21424 & w21479;
assign w21481 = w21424 & ~w21479;
assign w21482 = ~w21480 & ~w21481;
assign w21483 = ~w21423 & w21482;
assign w21484 = w21482 & ~w21483;
assign w21485 = ~w21482 & ~w21423;
assign w21486 = ~w21484 & ~w21485;
assign w21487 = (~w21275 & w21202) | (~w21275 & w41813) | (w21202 & w41813);
assign w21488 = w21486 & w21487;
assign w21489 = ~w21486 & ~w21487;
assign w21490 = ~w21488 & ~w21489;
assign w21491 = b_46 & w7613;
assign w21492 = w7941 & w32016;
assign w21493 = b_45 & w7608;
assign w21494 = ~w21492 & ~w21493;
assign w21495 = ~w21491 & w21494;
assign w21496 = (w21495 & ~w6974) | (w21495 & w26016) | (~w6974 & w26016);
assign w21497 = (w6974 & w26426) | (w6974 & w26427) | (w26426 & w26427);
assign w21498 = (~w6974 & w26712) | (~w6974 & w26713) | (w26712 & w26713);
assign w21499 = ~w21496 & ~w21497;
assign w21500 = ~w21498 & ~w21499;
assign w21501 = w21500 & w21490;
assign w21502 = ~w21490 & ~w21500;
assign w21503 = ~w21501 & ~w21502;
assign w21504 = (~w21292 & ~w21294) | (~w21292 & w32017) | (~w21294 & w32017);
assign w21505 = w21503 & w21504;
assign w21506 = ~w21503 & ~w21504;
assign w21507 = ~w21505 & ~w21506;
assign w21508 = b_49 & w6761;
assign w21509 = w7075 & w32018;
assign w21510 = b_48 & w6756;
assign w21511 = ~w21509 & ~w21510;
assign w21512 = ~w21508 & w21511;
assign w21513 = (w21512 & ~w7859) | (w21512 & w26017) | (~w7859 & w26017);
assign w21514 = (w7859 & w26428) | (w7859 & w26429) | (w26428 & w26429);
assign w21515 = (~w7859 & w32019) | (~w7859 & w32020) | (w32019 & w32020);
assign w21516 = ~w21513 & ~w21514;
assign w21517 = ~w21515 & ~w21516;
assign w21518 = w21507 & ~w21517;
assign w21519 = w21507 & ~w21518;
assign w21520 = ~w21507 & ~w21517;
assign w21521 = (~w26421 & w32021) | (~w26421 & w32022) | (w32021 & w32022);
assign w21522 = ~w21519 & w32023;
assign w21523 = (~w21521 & w21519) | (~w21521 & w32024) | (w21519 & w32024);
assign w21524 = ~w21522 & ~w21523;
assign w21525 = b_52 & w5962;
assign w21526 = w6246 & w32025;
assign w21527 = b_51 & w5957;
assign w21528 = ~w21526 & ~w21527;
assign w21529 = ~w21525 & w21528;
assign w21530 = (w21529 & ~w8793) | (w21529 & w26430) | (~w8793 & w26430);
assign w21531 = (w8793 & w32026) | (w8793 & w32027) | (w32026 & w32027);
assign w21532 = (~w8793 & w32028) | (~w8793 & w32029) | (w32028 & w32029);
assign w21533 = ~w21530 & ~w21531;
assign w21534 = ~w21532 & ~w21533;
assign w21535 = w21524 & ~w21534;
assign w21536 = w21524 & ~w21535;
assign w21537 = ~w21524 & ~w21534;
assign w21538 = ~w21536 & ~w21537;
assign w21539 = (w21329 & w21536) | (w21329 & w26714) | (w21536 & w26714);
assign w21540 = b_55 & w5196;
assign w21541 = w5459 & w32030;
assign w21542 = b_54 & w5191;
assign w21543 = ~w21541 & ~w21542;
assign w21544 = ~w21540 & w21543;
assign w21545 = (w21544 & ~w9776) | (w21544 & w32031) | (~w9776 & w32031);
assign w21546 = (w9776 & w41814) | (w9776 & w41815) | (w41814 & w41815);
assign w21547 = (~w9776 & w41816) | (~w9776 & w41817) | (w41816 & w41817);
assign w21548 = ~w21545 & ~w21546;
assign w21549 = ~w21547 & ~w21548;
assign w21550 = (~w21549 & w21539) | (~w21549 & w32032) | (w21539 & w32032);
assign w21551 = ~w21539 & w32033;
assign w21552 = ~w21550 & ~w21551;
assign w21553 = ~w21413 & w21552;
assign w21554 = w21413 & ~w21552;
assign w21555 = ~w21553 & ~w21554;
assign w21556 = ~w21412 & w21555;
assign w21557 = w21555 & ~w21556;
assign w21558 = ~w21555 & ~w21412;
assign w21559 = ~w21557 & ~w21558;
assign w21560 = (~w31975 & w41818) | (~w31975 & w41819) | (w41818 & w41819);
assign w21561 = w21559 & w21560;
assign w21562 = ~w21559 & ~w21560;
assign w21563 = ~w21561 & ~w21562;
assign w21564 = b_61 & w3803;
assign w21565 = w4027 & w32034;
assign w21566 = b_60 & w3798;
assign w21567 = ~w21565 & ~w21566;
assign w21568 = ~w21564 & w21567;
assign w21569 = (w21568 & ~w11901) | (w21568 & w32035) | (~w11901 & w32035);
assign w21570 = (w11901 & w41820) | (w11901 & w41821) | (w41820 & w41821);
assign w21571 = (~w11901 & w41822) | (~w11901 & w41823) | (w41822 & w41823);
assign w21572 = ~w21569 & ~w21570;
assign w21573 = ~w21571 & ~w21572;
assign w21574 = w21563 & ~w21573;
assign w21575 = ~w21563 & w21573;
assign w21576 = w21402 & w32036;
assign w21577 = w21402 & ~w21576;
assign w21578 = ~w21402 & w32036;
assign w21579 = ~w21577 & ~w21578;
assign w21580 = (~w21383 & w41824) | (~w21383 & w41825) | (w41824 & w41825);
assign w21581 = (~w21579 & w21385) | (~w21579 & w32037) | (w21385 & w32037);
assign w21582 = ~w21579 & ~w21581;
assign w21583 = ~w21580 & ~w21581;
assign w21584 = ~w21582 & ~w21583;
assign w21585 = (~w13761 & w37724) | (~w13761 & w37725) | (w37724 & w37725);
assign w21586 = (w13761 & w37726) | (w13761 & w37727) | (w37726 & w37727);
assign w21587 = ~w21585 & ~w21586;
assign w21588 = (~w21400 & ~w21402) | (~w21400 & w41826) | (~w21402 & w41826);
assign w21589 = (~w21562 & ~w21563) | (~w21562 & w27650) | (~w21563 & w27650);
assign w21590 = w3388 & w32040;
assign w21591 = (~w21590 & ~w12670) | (~w21590 & w32041) | (~w12670 & w32041);
assign w21592 = (w12670 & w41827) | (w12670 & w41828) | (w41827 & w41828);
assign w21593 = (~w12670 & w41829) | (~w12670 & w41830) | (w41829 & w41830);
assign w21594 = ~w21591 & ~w21592;
assign w21595 = ~w21593 & ~w21594;
assign w21596 = (w21563 & w41831) | (w21563 & w41832) | (w41831 & w41832);
assign w21597 = ~w21589 & ~w21596;
assign w21598 = (~w21563 & w41833) | (~w21563 & w41834) | (w41833 & w41834);
assign w21599 = ~w21329 & ~w21538;
assign w21600 = b_56 & w5196;
assign w21601 = w5459 & w32042;
assign w21602 = b_55 & w5191;
assign w21603 = ~w21601 & ~w21602;
assign w21604 = ~w21600 & w21603;
assign w21605 = (w21604 & ~w9798) | (w21604 & w26431) | (~w9798 & w26431);
assign w21606 = (w9798 & w32043) | (w9798 & w32044) | (w32043 & w32044);
assign w21607 = (~w9798 & w32045) | (~w9798 & w32046) | (w32045 & w32046);
assign w21608 = ~w21605 & ~w21606;
assign w21609 = ~w21607 & ~w21608;
assign w21610 = (~w21523 & ~w21524) | (~w21523 & w27651) | (~w21524 & w27651);
assign w21611 = b_53 & w5962;
assign w21612 = w6246 & w32047;
assign w21613 = b_52 & w5957;
assign w21614 = ~w21612 & ~w21613;
assign w21615 = ~w21611 & w21614;
assign w21616 = (w9109 & w41835) | (w9109 & w41836) | (w41835 & w41836);
assign w21617 = (~w9109 & w41837) | (~w9109 & w41838) | (w41837 & w41838);
assign w21618 = (w9109 & w41839) | (w9109 & w41840) | (w41839 & w41840);
assign w21619 = ~w21616 & ~w21617;
assign w21620 = ~w21618 & ~w21619;
assign w21621 = (~w21506 & ~w21507) | (~w21506 & w27652) | (~w21507 & w27652);
assign w21622 = (~w21480 & ~w21482) | (~w21480 & w32052) | (~w21482 & w32052);
assign w21623 = b_44 & w8526;
assign w21624 = w8886 & w32053;
assign w21625 = b_43 & w8521;
assign w21626 = ~w21624 & ~w21625;
assign w21627 = ~w21623 & w21626;
assign w21628 = (w21627 & ~w6408) | (w21627 & w26018) | (~w6408 & w26018);
assign w21629 = (w6408 & w26433) | (w6408 & w26434) | (w26433 & w26434);
assign w21630 = (~w6408 & w27653) | (~w6408 & w27654) | (w27653 & w27654);
assign w21631 = ~w21628 & ~w21629;
assign w21632 = ~w21630 & ~w21631;
assign w21633 = (~w21472 & w21475) | (~w21472 & w32054) | (w21475 & w32054);
assign w21634 = b_41 & w9534;
assign w21635 = w9876 & w32055;
assign w21636 = b_40 & w9529;
assign w21637 = ~w21635 & ~w21636;
assign w21638 = ~w21634 & w21637;
assign w21639 = (w21638 & ~w5609) | (w21638 & w27655) | (~w5609 & w27655);
assign w21640 = (w5609 & w32056) | (w5609 & w32057) | (w32056 & w32057);
assign w21641 = (~w5609 & w32058) | (~w5609 & w32059) | (w32058 & w32059);
assign w21642 = ~w21639 & ~w21640;
assign w21643 = ~w21641 & ~w21642;
assign w21644 = ~w21465 & ~w21468;
assign w21645 = (~w21461 & w41841) | (~w21461 & w41842) | (w41841 & w41842);
assign w21646 = w12380 & w32060;
assign w21647 = b_32 & ~w12380;
assign w21648 = ~w21646 & ~w21647;
assign w21649 = ~w21449 & w21648;
assign w21650 = w21449 & ~w21648;
assign w21651 = (w21461 & w41843) | (w21461 & w41844) | (w41843 & w41844);
assign w21652 = ~w21645 & ~w21651;
assign w21653 = (~w21461 & w41845) | (~w21461 & w41846) | (w41845 & w41846);
assign w21654 = (~w21461 & w41847) | (~w21461 & w41848) | (w41847 & w41848);
assign w21655 = ~w21652 & ~w21654;
assign w21656 = b_35 & w11620;
assign w21657 = w11969 & w32067;
assign w21658 = b_34 & w11615;
assign w21659 = ~w21657 & ~w21658;
assign w21660 = ~w21656 & w21659;
assign w21661 = (w21660 & ~w4181) | (w21660 & w32068) | (~w4181 & w32068);
assign w21662 = (w4181 & w41849) | (w4181 & w41850) | (w41849 & w41850);
assign w21663 = (~w4181 & w41851) | (~w4181 & w41852) | (w41851 & w41852);
assign w21664 = ~w21661 & ~w21662;
assign w21665 = ~w21663 & ~w21664;
assign w21666 = (~w21665 & w21652) | (~w21665 & w32069) | (w21652 & w32069);
assign w21667 = ~w21655 & ~w21666;
assign w21668 = ~w21665 & ~w21666;
assign w21669 = ~w21667 & ~w21668;
assign w21670 = b_38 & w10562;
assign w21671 = w10902 & w32070;
assign w21672 = b_37 & w10557;
assign w21673 = ~w21671 & ~w21672;
assign w21674 = ~w21670 & w21673;
assign w21675 = (w21674 & ~w4658) | (w21674 & w32071) | (~w4658 & w32071);
assign w21676 = (w4658 & w41853) | (w4658 & w41854) | (w41853 & w41854);
assign w21677 = (~w4658 & w41855) | (~w4658 & w41856) | (w41855 & w41856);
assign w21678 = ~w21675 & ~w21676;
assign w21679 = ~w21677 & ~w21678;
assign w21680 = ~w21669 & w21679;
assign w21681 = w21669 & ~w21679;
assign w21682 = ~w21680 & ~w21681;
assign w21683 = ~w21644 & ~w21682;
assign w21684 = w21644 & w21682;
assign w21685 = ~w21683 & ~w21684;
assign w21686 = ~w21643 & w21685;
assign w21687 = w21643 & ~w21685;
assign w21688 = ~w21686 & ~w21687;
assign w21689 = ~w21633 & w21688;
assign w21690 = w21633 & ~w21688;
assign w21691 = ~w21689 & ~w21690;
assign w21692 = ~w21632 & w21691;
assign w21693 = w21632 & ~w21691;
assign w21694 = ~w21692 & ~w21693;
assign w21695 = ~w21622 & w21694;
assign w21696 = w21622 & ~w21694;
assign w21697 = ~w21695 & ~w21696;
assign w21698 = b_47 & w7613;
assign w21699 = w7941 & w32072;
assign w21700 = b_46 & w7608;
assign w21701 = ~w21699 & ~w21700;
assign w21702 = ~w21698 & w21701;
assign w21703 = (w21702 & ~w6998) | (w21702 & w25460) | (~w6998 & w25460);
assign w21704 = (w6998 & w25680) | (w6998 & w25681) | (w25680 & w25681);
assign w21705 = (~w6998 & w26019) | (~w6998 & w26020) | (w26019 & w26020);
assign w21706 = ~w21703 & ~w21704;
assign w21707 = ~w21705 & ~w21706;
assign w21708 = w21697 & w21707;
assign w21709 = (~w26435 & w32073) | (~w26435 & w32074) | (w32073 & w32074);
assign w21710 = (~w21489 & ~w21490) | (~w21489 & w32075) | (~w21490 & w32075);
assign w21711 = w21710 & w32076;
assign w21712 = (~w21710 & w21709) | (~w21710 & w26021) | (w21709 & w26021);
assign w21713 = ~w21711 & ~w21712;
assign w21714 = b_50 & w6761;
assign w21715 = w7075 & w32077;
assign w21716 = b_49 & w6756;
assign w21717 = ~w21715 & ~w21716;
assign w21718 = ~w21714 & w21717;
assign w21719 = (w21718 & ~w8162) | (w21718 & w26022) | (~w8162 & w26022);
assign w21720 = (w8162 & w26436) | (w8162 & w26437) | (w26436 & w26437);
assign w21721 = (~w8162 & w27656) | (~w8162 & w27657) | (w27656 & w27657);
assign w21722 = ~w21719 & ~w21720;
assign w21723 = ~w21721 & ~w21722;
assign w21724 = (w21723 & w21712) | (w21723 & w32078) | (w21712 & w32078);
assign w21725 = ~w21712 & w32079;
assign w21726 = ~w21724 & ~w21725;
assign w21727 = ~w21621 & w21726;
assign w21728 = ~w21726 & ~w21621;
assign w21729 = w21726 & ~w21727;
assign w21730 = (~w21620 & w21729) | (~w21620 & w27658) | (w21729 & w27658);
assign w21731 = ~w21729 & w27659;
assign w21732 = ~w21730 & ~w21731;
assign w21733 = ~w21610 & w21732;
assign w21734 = w21610 & ~w21732;
assign w21735 = ~w21733 & ~w21734;
assign w21736 = ~w21609 & w21735;
assign w21737 = w21609 & ~w21735;
assign w21738 = ~w21736 & ~w21737;
assign w21739 = (w21738 & w21550) | (w21738 & w32080) | (w21550 & w32080);
assign w21740 = ~w21550 & w32081;
assign w21741 = ~w21739 & ~w21740;
assign w21742 = b_59 & w4499;
assign w21743 = w4723 & w32082;
assign w21744 = b_58 & w4494;
assign w21745 = ~w21743 & ~w21744;
assign w21746 = ~w21742 & w21745;
assign w21747 = (w21746 & ~w11169) | (w21746 & w32083) | (~w11169 & w32083);
assign w21748 = (w11169 & w41857) | (w11169 & w41858) | (w41857 & w41858);
assign w21749 = (~w11169 & w41859) | (~w11169 & w41860) | (w41859 & w41860);
assign w21750 = ~w21747 & ~w21748;
assign w21751 = ~w21749 & ~w21750;
assign w21752 = w21741 & ~w21751;
assign w21753 = w21741 & ~w21752;
assign w21754 = ~w21741 & ~w21751;
assign w21755 = ~w21753 & ~w21754;
assign w21756 = (~w21553 & ~w21555) | (~w21553 & w32084) | (~w21555 & w32084);
assign w21757 = w21755 & w21756;
assign w21758 = ~w21755 & ~w21756;
assign w21759 = ~w21757 & ~w21758;
assign w21760 = b_62 & w3803;
assign w21761 = w4027 & w32085;
assign w21762 = b_61 & w3798;
assign w21763 = ~w21761 & ~w21762;
assign w21764 = ~w21760 & w21763;
assign w21765 = (w21764 & ~w12273) | (w21764 & w32086) | (~w12273 & w32086);
assign w21766 = (w12273 & w41861) | (w12273 & w41862) | (w41861 & w41862);
assign w21767 = (~w12273 & w41863) | (~w12273 & w41864) | (w41863 & w41864);
assign w21768 = ~w21765 & ~w21766;
assign w21769 = ~w21767 & ~w21768;
assign w21770 = w21759 & ~w21769;
assign w21771 = w21759 & ~w21770;
assign w21772 = ~w21759 & ~w21769;
assign w21773 = ~w21771 & ~w21772;
assign w21774 = (w21773 & w21597) | (w21773 & w32087) | (w21597 & w32087);
assign w21775 = ~w21597 & w32088;
assign w21776 = ~w21774 & ~w21775;
assign w21777 = ~w21588 & ~w21776;
assign w21778 = w21776 & ~w21588;
assign w21779 = ~w21776 & ~w21777;
assign w21780 = ~w21778 & ~w21779;
assign w21781 = (~w13761 & w37728) | (~w13761 & w37729) | (w37728 & w37729);
assign w21782 = (w13761 & w37730) | (w13761 & w37731) | (w37730 & w37731);
assign w21783 = ~w21781 & ~w21782;
assign w21784 = (~w21773 & w21597) | (~w21773 & w32093) | (w21597 & w32093);
assign w21785 = b_57 & w5196;
assign w21786 = w5459 & w32094;
assign w21787 = b_56 & w5191;
assign w21788 = ~w21786 & ~w21787;
assign w21789 = ~w21785 & w21788;
assign w21790 = (w21789 & ~w10452) | (w21789 & w32095) | (~w10452 & w32095);
assign w21791 = (w10452 & w41865) | (w10452 & w41866) | (w41865 & w41866);
assign w21792 = (~w10452 & w41867) | (~w10452 & w41868) | (w41867 & w41868);
assign w21793 = ~w21790 & ~w21791;
assign w21794 = ~w21792 & ~w21793;
assign w21795 = ~w21727 & ~w21730;
assign w21796 = (~w21712 & ~w21713) | (~w21712 & w26438) | (~w21713 & w26438);
assign w21797 = b_42 & w9534;
assign w21798 = w9876 & w32096;
assign w21799 = b_41 & w9529;
assign w21800 = ~w21798 & ~w21799;
assign w21801 = ~w21797 & w21800;
assign w21802 = (w21801 & ~w5864) | (w21801 & w25682) | (~w5864 & w25682);
assign w21803 = (w5864 & w26023) | (w5864 & w26024) | (w26023 & w26024);
assign w21804 = (~w5864 & w26439) | (~w5864 & w26440) | (w26439 & w26440);
assign w21805 = ~w21802 & ~w21803;
assign w21806 = ~w21804 & ~w21805;
assign w21807 = (~w21666 & w21669) | (~w21666 & w32097) | (w21669 & w32097);
assign w21808 = w12380 & w41869;
assign w21809 = (~a_32 & w21808) | (~a_32 & w32098) | (w21808 & w32098);
assign w21810 = ~w21808 & w32099;
assign w21811 = ~w21809 & ~w21810;
assign w21812 = ~w21648 & w21811;
assign w21813 = ~w21811 & ~w21648;
assign w21814 = w21811 & ~w21812;
assign w21815 = ~w21813 & ~w21814;
assign w21816 = (w21461 & w41870) | (w21461 & w41871) | (w41870 & w41871);
assign w21817 = ~w21653 & ~w21816;
assign w21818 = (~w21461 & w41872) | (~w21461 & w41873) | (w41872 & w41873);
assign w21819 = b_36 & w11620;
assign w21820 = w11969 & w32104;
assign w21821 = b_35 & w11615;
assign w21822 = ~w21820 & ~w21821;
assign w21823 = ~w21819 & w21822;
assign w21824 = (w21823 & ~w4395) | (w21823 & w32105) | (~w4395 & w32105);
assign w21825 = (w4395 & w41874) | (w4395 & w41875) | (w41874 & w41875);
assign w21826 = (~w4395 & w41876) | (~w4395 & w41877) | (w41876 & w41877);
assign w21827 = ~w21824 & ~w21825;
assign w21828 = ~w21826 & ~w21827;
assign w21829 = (w21828 & w21817) | (w21828 & w32106) | (w21817 & w32106);
assign w21830 = ~w21817 & w32107;
assign w21831 = ~w21829 & ~w21830;
assign w21832 = b_39 & w10562;
assign w21833 = w10902 & w32108;
assign w21834 = b_38 & w10557;
assign w21835 = ~w21833 & ~w21834;
assign w21836 = ~w21832 & w21835;
assign w21837 = (w21836 & ~w4888) | (w21836 & w26441) | (~w4888 & w26441);
assign w21838 = (w4888 & w32109) | (w4888 & w32110) | (w32109 & w32110);
assign w21839 = (~w4888 & w32111) | (~w4888 & w32112) | (w32111 & w32112);
assign w21840 = ~w21837 & ~w21838;
assign w21841 = ~w21839 & ~w21840;
assign w21842 = ~w21831 & ~w21841;
assign w21843 = w21831 & w21841;
assign w21844 = ~w21842 & ~w21843;
assign w21845 = ~w21807 & w21844;
assign w21846 = w21807 & ~w21844;
assign w21847 = ~w21845 & ~w21846;
assign w21848 = ~w21806 & w21847;
assign w21849 = w21806 & w21847;
assign w21850 = ~w21847 & ~w21806;
assign w21851 = ~w21849 & ~w21850;
assign w21852 = (~w21683 & ~w21685) | (~w21683 & w32113) | (~w21685 & w32113);
assign w21853 = w21851 & w21852;
assign w21854 = ~w21851 & ~w21852;
assign w21855 = ~w21853 & ~w21854;
assign w21856 = b_45 & w8526;
assign w21857 = w8886 & w32114;
assign w21858 = b_44 & w8521;
assign w21859 = ~w21857 & ~w21858;
assign w21860 = ~w21856 & w21859;
assign w21861 = (w21860 & ~w6682) | (w21860 & w25461) | (~w6682 & w25461);
assign w21862 = (w6682 & w25683) | (w6682 & w25684) | (w25683 & w25684);
assign w21863 = (~w6682 & w26025) | (~w6682 & w26026) | (w26025 & w26026);
assign w21864 = ~w21861 & ~w21862;
assign w21865 = ~w21863 & ~w21864;
assign w21866 = w21855 & ~w21865;
assign w21867 = w21865 & w21855;
assign w21868 = ~w21855 & ~w21865;
assign w21869 = (~w21689 & ~w21691) | (~w21689 & w32115) | (~w21691 & w32115);
assign w21870 = w21869 & w32116;
assign w21871 = (~w21869 & w21868) | (~w21869 & w26027) | (w21868 & w26027);
assign w21872 = b_48 & w7613;
assign w21873 = w7941 & w32117;
assign w21874 = b_47 & w7608;
assign w21875 = ~w21873 & ~w21874;
assign w21876 = ~w21872 & w21875;
assign w21877 = (w21876 & ~w7284) | (w21876 & w25462) | (~w7284 & w25462);
assign w21878 = (w7284 & w25685) | (w7284 & w25686) | (w25685 & w25686);
assign w21879 = (~w7284 & w26028) | (~w7284 & w26029) | (w26028 & w26029);
assign w21880 = ~w21877 & ~w21878;
assign w21881 = ~w21879 & ~w21880;
assign w21882 = ~w21871 & w32118;
assign w21883 = ~w21871 & w32119;
assign w21884 = ~w21881 & ~w21882;
assign w21885 = (~w26435 & w32120) | (~w26435 & w32121) | (w32120 & w32121);
assign w21886 = w21885 & w41878;
assign w21887 = (~w21885 & w21884) | (~w21885 & w26030) | (w21884 & w26030);
assign w21888 = ~w21886 & ~w21887;
assign w21889 = b_51 & w6761;
assign w21890 = w7075 & w32122;
assign w21891 = b_50 & w6756;
assign w21892 = ~w21890 & ~w21891;
assign w21893 = ~w21889 & w21892;
assign w21894 = (w21893 & ~w8186) | (w21893 & w25687) | (~w8186 & w25687);
assign w21895 = (w8186 & w26031) | (w8186 & w26032) | (w26031 & w26032);
assign w21896 = (~w8186 & w26442) | (~w8186 & w26443) | (w26442 & w26443);
assign w21897 = ~w21894 & ~w21895;
assign w21898 = ~w21896 & ~w21897;
assign w21899 = ~w21887 & w41879;
assign w21900 = (w21898 & w21887) | (w21898 & w41880) | (w21887 & w41880);
assign w21901 = (~w32124 & w41881) | (~w32124 & w41882) | (w41881 & w41882);
assign w21902 = (~w26715 & w32125) | (~w26715 & w32126) | (w32125 & w32126);
assign w21903 = (w32126 & w41883) | (w32126 & w41884) | (w41883 & w41884);
assign w21904 = ~w21901 & ~w21903;
assign w21905 = b_54 & w5962;
assign w21906 = w6246 & w32127;
assign w21907 = b_53 & w5957;
assign w21908 = ~w21906 & ~w21907;
assign w21909 = ~w21905 & w21908;
assign w21910 = (w21909 & ~w9134) | (w21909 & w26444) | (~w9134 & w26444);
assign w21911 = (w9134 & w32128) | (w9134 & w32129) | (w32128 & w32129);
assign w21912 = (~w9134 & w32130) | (~w9134 & w32131) | (w32130 & w32131);
assign w21913 = ~w21910 & ~w21911;
assign w21914 = ~w21912 & ~w21913;
assign w21915 = w21904 & w21914;
assign w21916 = ~w21904 & ~w21914;
assign w21917 = ~w21915 & ~w21916;
assign w21918 = ~w21795 & w21917;
assign w21919 = w21795 & ~w21917;
assign w21920 = ~w21918 & ~w21919;
assign w21921 = ~w21794 & w21920;
assign w21922 = w21920 & ~w21921;
assign w21923 = (~w21733 & ~w21735) | (~w21733 & w32132) | (~w21735 & w32132);
assign w21924 = ~w21922 & w27660;
assign w21925 = (~w21923 & w21922) | (~w21923 & w27661) | (w21922 & w27661);
assign w21926 = ~w21924 & ~w21925;
assign w21927 = b_60 & w4499;
assign w21928 = w4723 & w32133;
assign w21929 = b_59 & w4494;
assign w21930 = ~w21928 & ~w21929;
assign w21931 = ~w21927 & w21930;
assign w21932 = (w21931 & ~w11196) | (w21931 & w32134) | (~w11196 & w32134);
assign w21933 = (w11196 & w41885) | (w11196 & w41886) | (w41885 & w41886);
assign w21934 = (~w11196 & w41887) | (~w11196 & w41888) | (w41887 & w41888);
assign w21935 = ~w21932 & ~w21933;
assign w21936 = ~w21934 & ~w21935;
assign w21937 = w21926 & ~w21936;
assign w21938 = w21926 & ~w21937;
assign w21939 = ~w21926 & ~w21936;
assign w21940 = (~w21739 & ~w21741) | (~w21739 & w32135) | (~w21741 & w32135);
assign w21941 = ~w21938 & w32136;
assign w21942 = (~w21940 & w21938) | (~w21940 & w32137) | (w21938 & w32137);
assign w21943 = ~w21941 & ~w21942;
assign w21944 = (~w21758 & ~w21759) | (~w21758 & w27662) | (~w21759 & w27662);
assign w21945 = b_63 & w3803;
assign w21946 = w4027 & w32138;
assign w21947 = b_62 & w3798;
assign w21948 = ~w21946 & ~w21947;
assign w21949 = ~w21945 & w21948;
assign w21950 = (w21949 & ~w12646) | (w21949 & w32139) | (~w12646 & w32139);
assign w21951 = (w12646 & w41889) | (w12646 & w41890) | (w41889 & w41890);
assign w21952 = (~w12646 & w41891) | (~w12646 & w41892) | (w41891 & w41892);
assign w21953 = ~w21950 & ~w21951;
assign w21954 = ~w21952 & ~w21953;
assign w21955 = ~w21944 & ~w21954;
assign w21956 = ~w21944 & ~w21955;
assign w21957 = ~w21956 & w32140;
assign w21958 = (w21943 & w21956) | (w21943 & w32141) | (w21956 & w32141);
assign w21959 = ~w21957 & ~w21958;
assign w21960 = (w21959 & w21784) | (w21959 & w32142) | (w21784 & w32142);
assign w21961 = ~w21784 & w32143;
assign w21962 = ~w21960 & ~w21961;
assign w21963 = (~w13761 & w37732) | (~w13761 & w37733) | (w37732 & w37733);
assign w21964 = (w13761 & w37734) | (w13761 & w37735) | (w37734 & w37735);
assign w21965 = ~w21963 & ~w21964;
assign w21966 = w4027 & w32144;
assign w21967 = b_63 & w3798;
assign w21968 = ~w21966 & ~w21967;
assign w21969 = ~w12671 & w32145;
assign w21970 = (a_35 & w21969) | (a_35 & w32146) | (w21969 & w32146);
assign w21971 = ~w21969 & w32147;
assign w21972 = ~w21970 & ~w21971;
assign w21973 = (~w21972 & w21942) | (~w21972 & w32148) | (w21942 & w32148);
assign w21974 = ~w21942 & w32149;
assign w21975 = ~w21973 & ~w21974;
assign w21976 = b_58 & w5196;
assign w21977 = w5459 & w32150;
assign w21978 = b_57 & w5191;
assign w21979 = ~w21977 & ~w21978;
assign w21980 = ~w21976 & w21979;
assign w21981 = (w21980 & ~w10476) | (w21980 & w32151) | (~w10476 & w32151);
assign w21982 = (w10476 & w41893) | (w10476 & w41894) | (w41893 & w41894);
assign w21983 = (~w10476 & w41895) | (~w10476 & w41896) | (w41895 & w41896);
assign w21984 = ~w21981 & ~w21982;
assign w21985 = ~w21983 & ~w21984;
assign w21986 = (~w21916 & ~w21917) | (~w21916 & w32152) | (~w21917 & w32152);
assign w21987 = b_43 & w9534;
assign w21988 = w9876 & w32153;
assign w21989 = b_42 & w9529;
assign w21990 = ~w21988 & ~w21989;
assign w21991 = ~w21987 & w21990;
assign w21992 = (w21991 & ~w5888) | (w21991 & w27663) | (~w5888 & w27663);
assign w21993 = (w5888 & w32154) | (w5888 & w32155) | (w32154 & w32155);
assign w21994 = (~w5888 & w32156) | (~w5888 & w32157) | (w32156 & w32157);
assign w21995 = ~w21992 & ~w21993;
assign w21996 = ~w21994 & ~w21995;
assign w21997 = ~w21842 & ~w21845;
assign w21998 = b_40 & w10562;
assign w21999 = w10902 & w32158;
assign w22000 = b_39 & w10557;
assign w22001 = ~w21999 & ~w22000;
assign w22002 = ~w21998 & w22001;
assign w22003 = (w22002 & ~w5363) | (w22002 & w32159) | (~w5363 & w32159);
assign w22004 = (w5363 & w41897) | (w5363 & w41898) | (w41897 & w41898);
assign w22005 = (~w5363 & w41899) | (~w5363 & w41900) | (w41899 & w41900);
assign w22006 = ~w22003 & ~w22004;
assign w22007 = ~w22005 & ~w22006;
assign w22008 = (~w21828 & w21817) | (~w21828 & w32160) | (w21817 & w32160);
assign w22009 = ~w21816 & ~w22008;
assign w22010 = w12380 & w32161;
assign w22011 = b_34 & ~w12380;
assign w22012 = ~w22010 & ~w22011;
assign w22013 = (~w21809 & ~w21811) | (~w21809 & w32162) | (~w21811 & w32162);
assign w22014 = ~w22012 & w22013;
assign w22015 = w22012 & ~w22013;
assign w22016 = ~w22014 & ~w22015;
assign w22017 = b_37 & w11620;
assign w22018 = w11969 & w32163;
assign w22019 = b_36 & w11615;
assign w22020 = ~w22018 & ~w22019;
assign w22021 = ~w22017 & w22020;
assign w22022 = (w22021 & ~w4636) | (w22021 & w25688) | (~w4636 & w25688);
assign w22023 = (w4636 & w26033) | (w4636 & w26034) | (w26033 & w26034);
assign w22024 = ~w22022 & ~w22023;
assign w22025 = ~w22024 & w32166;
assign w22026 = (w22016 & w22024) | (w22016 & w32167) | (w22024 & w32167);
assign w22027 = ~w22025 & ~w22026;
assign w22028 = (w22027 & w22008) | (w22027 & w32168) | (w22008 & w32168);
assign w22029 = ~w22009 & ~w22028;
assign w22030 = ~w22008 & w32169;
assign w22031 = (~w22007 & w22029) | (~w22007 & w32170) | (w22029 & w32170);
assign w22032 = (w22007 & ~w32169) | (w22007 & w41901) | (~w32169 & w41901);
assign w22033 = ~w22029 & w22032;
assign w22034 = ~w22031 & ~w22033;
assign w22035 = ~w21997 & w22034;
assign w22036 = w21997 & ~w22034;
assign w22037 = ~w22035 & ~w22036;
assign w22038 = ~w21996 & w22037;
assign w22039 = w22037 & ~w22038;
assign w22040 = ~w22037 & ~w21996;
assign w22041 = ~w22039 & ~w22040;
assign w22042 = ~w21848 & ~w21854;
assign w22043 = w22041 & w22042;
assign w22044 = ~w22041 & ~w22042;
assign w22045 = ~w22043 & ~w22044;
assign w22046 = b_46 & w8526;
assign w22047 = w8886 & w32171;
assign w22048 = b_45 & w8521;
assign w22049 = ~w22047 & ~w22048;
assign w22050 = ~w22046 & w22049;
assign w22051 = (w22050 & ~w6974) | (w22050 & w26716) | (~w6974 & w26716);
assign w22052 = (w6974 & w27664) | (w6974 & w27665) | (w27664 & w27665);
assign w22053 = (~w6974 & w32172) | (~w6974 & w32173) | (w32172 & w32173);
assign w22054 = ~w22051 & ~w22052;
assign w22055 = ~w22053 & ~w22054;
assign w22056 = w22045 & ~w22055;
assign w22057 = w22045 & ~w22056;
assign w22058 = ~w22045 & ~w22055;
assign w22059 = (~w26027 & w32174) | (~w26027 & w32175) | (w32174 & w32175);
assign w22060 = ~w22057 & w32176;
assign w22061 = (~w22059 & w22057) | (~w22059 & w32177) | (w22057 & w32177);
assign w22062 = ~w22060 & ~w22061;
assign w22063 = b_49 & w7613;
assign w22064 = w7941 & w32178;
assign w22065 = b_48 & w7608;
assign w22066 = ~w22064 & ~w22065;
assign w22067 = ~w22063 & w22066;
assign w22068 = (w22067 & ~w7859) | (w22067 & w27666) | (~w7859 & w27666);
assign w22069 = (w7859 & w32179) | (w7859 & w32180) | (w32179 & w32180);
assign w22070 = (~w7859 & w32181) | (~w7859 & w32182) | (w32181 & w32182);
assign w22071 = ~w22068 & ~w22069;
assign w22072 = ~w22070 & ~w22071;
assign w22073 = w22062 & ~w22072;
assign w22074 = w22062 & ~w22073;
assign w22075 = ~w22062 & ~w22072;
assign w22076 = ~w22074 & ~w22075;
assign w22077 = (~w26030 & w32183) | (~w26030 & w32184) | (w32183 & w32184);
assign w22078 = w22076 & w22077;
assign w22079 = ~w22076 & ~w22077;
assign w22080 = ~w22078 & ~w22079;
assign w22081 = b_52 & w6761;
assign w22082 = w7075 & w32185;
assign w22083 = b_51 & w6756;
assign w22084 = ~w22082 & ~w22083;
assign w22085 = ~w22081 & w22084;
assign w22086 = (w22085 & ~w8793) | (w22085 & w32186) | (~w8793 & w32186);
assign w22087 = (w8793 & w41902) | (w8793 & w41903) | (w41902 & w41903);
assign w22088 = (~w8793 & w41904) | (~w8793 & w41905) | (w41904 & w41905);
assign w22089 = ~w22086 & ~w22087;
assign w22090 = ~w22088 & ~w22089;
assign w22091 = w22080 & ~w22090;
assign w22092 = w22080 & ~w22091;
assign w22093 = ~w22080 & ~w22090;
assign w22094 = ~w22092 & ~w22093;
assign w22095 = ~w21902 & w22094;
assign w22096 = w21902 & ~w22094;
assign w22097 = ~w22095 & ~w22096;
assign w22098 = b_55 & w5962;
assign w22099 = w6246 & w32187;
assign w22100 = b_54 & w5957;
assign w22101 = ~w22099 & ~w22100;
assign w22102 = ~w22098 & w22101;
assign w22103 = (w22102 & ~w9776) | (w22102 & w32188) | (~w9776 & w32188);
assign w22104 = (w9776 & w41906) | (w9776 & w41907) | (w41906 & w41907);
assign w22105 = (~w9776 & w41908) | (~w9776 & w41909) | (w41908 & w41909);
assign w22106 = ~w22103 & ~w22104;
assign w22107 = ~w22105 & ~w22106;
assign w22108 = ~w22097 & ~w22107;
assign w22109 = w22097 & w22107;
assign w22110 = ~w22108 & ~w22109;
assign w22111 = ~w21986 & w22110;
assign w22112 = w21986 & ~w22110;
assign w22113 = ~w22111 & ~w22112;
assign w22114 = ~w21985 & w22113;
assign w22115 = w22113 & ~w22114;
assign w22116 = ~w22113 & ~w21985;
assign w22117 = ~w22115 & ~w22116;
assign w22118 = (~w27661 & w41910) | (~w27661 & w41911) | (w41910 & w41911);
assign w22119 = w22117 & w22118;
assign w22120 = ~w22117 & ~w22118;
assign w22121 = ~w22119 & ~w22120;
assign w22122 = b_61 & w4499;
assign w22123 = w4723 & w32189;
assign w22124 = b_60 & w4494;
assign w22125 = ~w22123 & ~w22124;
assign w22126 = ~w22122 & w22125;
assign w22127 = (w22126 & ~w11901) | (w22126 & w32190) | (~w11901 & w32190);
assign w22128 = (w11901 & w41912) | (w11901 & w41913) | (w41912 & w41913);
assign w22129 = (~w11901 & w41914) | (~w11901 & w41915) | (w41914 & w41915);
assign w22130 = ~w22127 & ~w22128;
assign w22131 = ~w22129 & ~w22130;
assign w22132 = w22121 & ~w22131;
assign w22133 = ~w22121 & w22131;
assign w22134 = w21975 & w32191;
assign w22135 = w21975 & ~w22134;
assign w22136 = (~w22133 & ~w21975) | (~w22133 & w32192) | (~w21975 & w32192);
assign w22137 = ~w22132 & w22136;
assign w22138 = ~w22135 & ~w22137;
assign w22139 = (~w21956 & w41916) | (~w21956 & w41917) | (w41916 & w41917);
assign w22140 = ~w22138 & ~w22139;
assign w22141 = w22139 & ~w22138;
assign w22142 = ~w22139 & ~w22140;
assign w22143 = ~w22141 & ~w22142;
assign w22144 = (~w13761 & w37736) | (~w13761 & w37737) | (w37736 & w37737);
assign w22145 = (w13761 & w37738) | (w13761 & w37739) | (w37738 & w37739);
assign w22146 = ~w22144 & ~w22145;
assign w22147 = (~w21973 & ~w21975) | (~w21973 & w32197) | (~w21975 & w32197);
assign w22148 = (~w22120 & ~w22121) | (~w22120 & w32198) | (~w22121 & w32198);
assign w22149 = w4027 & w32199;
assign w22150 = (~w22149 & ~w12670) | (~w22149 & w32200) | (~w12670 & w32200);
assign w22151 = (w12670 & w41918) | (w12670 & w41919) | (w41918 & w41919);
assign w22152 = (~w12670 & w41920) | (~w12670 & w41921) | (w41920 & w41921);
assign w22153 = ~w22150 & ~w22151;
assign w22154 = ~w22152 & ~w22153;
assign w22155 = ~w22148 & ~w22154;
assign w22156 = ~w22148 & ~w22155;
assign w22157 = w22148 & ~w22154;
assign w22158 = ~w21902 & ~w22094;
assign w22159 = (~w22158 & w22097) | (~w22158 & w32201) | (w22097 & w32201);
assign w22160 = b_56 & w5962;
assign w22161 = w6246 & w32202;
assign w22162 = b_55 & w5957;
assign w22163 = ~w22161 & ~w22162;
assign w22164 = ~w22160 & w22163;
assign w22165 = (w22164 & ~w9798) | (w22164 & w32203) | (~w9798 & w32203);
assign w22166 = (w9798 & w41922) | (w9798 & w41923) | (w41922 & w41923);
assign w22167 = (~w9798 & w41924) | (~w9798 & w41925) | (w41924 & w41925);
assign w22168 = ~w22165 & ~w22166;
assign w22169 = ~w22167 & ~w22168;
assign w22170 = (~w22079 & ~w22080) | (~w22079 & w32204) | (~w22080 & w32204);
assign w22171 = b_53 & w6761;
assign w22172 = w7075 & w32205;
assign w22173 = b_52 & w6756;
assign w22174 = ~w22172 & ~w22173;
assign w22175 = ~w22171 & w22174;
assign w22176 = (w9109 & w41926) | (w9109 & w41927) | (w41926 & w41927);
assign w22177 = a_47 & ~w22176;
assign w22178 = w22176 & a_47;
assign w22179 = ~w22176 & ~w22177;
assign w22180 = ~w22178 & ~w22179;
assign w22181 = (~w22061 & ~w22062) | (~w22061 & w32207) | (~w22062 & w32207);
assign w22182 = (~w22035 & ~w22037) | (~w22035 & w32208) | (~w22037 & w32208);
assign w22183 = b_44 & w9534;
assign w22184 = w9876 & w32209;
assign w22185 = b_43 & w9529;
assign w22186 = ~w22184 & ~w22185;
assign w22187 = ~w22183 & w22186;
assign w22188 = (w22187 & ~w6408) | (w22187 & w27667) | (~w6408 & w27667);
assign w22189 = (w6408 & w32210) | (w6408 & w32211) | (w32210 & w32211);
assign w22190 = (~w6408 & w32212) | (~w6408 & w32213) | (w32212 & w32213);
assign w22191 = ~w22188 & ~w22189;
assign w22192 = ~w22190 & ~w22191;
assign w22193 = (~w32170 & w41928) | (~w32170 & w41929) | (w41928 & w41929);
assign w22194 = (~w22024 & w41930) | (~w22024 & w41931) | (w41930 & w41931);
assign w22195 = w12380 & w32214;
assign w22196 = b_35 & ~w12380;
assign w22197 = ~w22195 & ~w22196;
assign w22198 = ~w22012 & w22197;
assign w22199 = w22012 & ~w22197;
assign w22200 = (w22024 & w41932) | (w22024 & w41933) | (w41932 & w41933);
assign w22201 = ~w22194 & ~w22200;
assign w22202 = (~w22024 & w41934) | (~w22024 & w41935) | (w41934 & w41935);
assign w22203 = ~w22201 & ~w22202;
assign w22204 = b_38 & w11620;
assign w22205 = w11969 & w32220;
assign w22206 = b_37 & w11615;
assign w22207 = ~w22205 & ~w22206;
assign w22208 = ~w22204 & w22207;
assign w22209 = (w22208 & ~w4658) | (w22208 & w32221) | (~w4658 & w32221);
assign w22210 = a_62 & ~w22209;
assign w22211 = w22209 & a_62;
assign w22212 = ~w22209 & ~w22210;
assign w22213 = ~w22211 & ~w22212;
assign w22214 = (~w22213 & w22201) | (~w22213 & w32222) | (w22201 & w32222);
assign w22215 = ~w22203 & ~w22214;
assign w22216 = ~w22213 & ~w22214;
assign w22217 = ~w22215 & ~w22216;
assign w22218 = b_41 & w10562;
assign w22219 = w10902 & w32223;
assign w22220 = b_40 & w10557;
assign w22221 = ~w22219 & ~w22220;
assign w22222 = ~w22218 & w22221;
assign w22223 = (w22222 & ~w5609) | (w22222 & w32224) | (~w5609 & w32224);
assign w22224 = a_59 & ~w22223;
assign w22225 = w22223 & a_59;
assign w22226 = ~w22223 & ~w22224;
assign w22227 = ~w22225 & ~w22226;
assign w22228 = ~w22217 & w22227;
assign w22229 = w22217 & ~w22227;
assign w22230 = ~w22228 & ~w22229;
assign w22231 = ~w22193 & ~w22230;
assign w22232 = w22193 & w22230;
assign w22233 = ~w22231 & ~w22232;
assign w22234 = ~w22192 & w22233;
assign w22235 = w22192 & ~w22233;
assign w22236 = ~w22234 & ~w22235;
assign w22237 = ~w22182 & w22236;
assign w22238 = w22182 & ~w22236;
assign w22239 = ~w22237 & ~w22238;
assign w22240 = b_47 & w8526;
assign w22241 = w8886 & w32225;
assign w22242 = b_46 & w8521;
assign w22243 = ~w22241 & ~w22242;
assign w22244 = ~w22240 & w22243;
assign w22245 = (w22244 & ~w6998) | (w22244 & w26035) | (~w6998 & w26035);
assign w22246 = (w6998 & w26445) | (w6998 & w26446) | (w26445 & w26446);
assign w22247 = (~w6998 & w27668) | (~w6998 & w27669) | (w27668 & w27669);
assign w22248 = ~w22245 & ~w22246;
assign w22249 = ~w22247 & ~w22248;
assign w22250 = w22249 & w22239;
assign w22251 = ~w22239 & ~w22249;
assign w22252 = (~w22044 & ~w22045) | (~w22044 & w32226) | (~w22045 & w32226);
assign w22253 = (~w22252 & w22251) | (~w22252 & w27670) | (w22251 & w27670);
assign w22254 = b_50 & w7613;
assign w22255 = w7941 & w32228;
assign w22256 = b_49 & w7608;
assign w22257 = ~w22255 & ~w22256;
assign w22258 = ~w22254 & w22257;
assign w22259 = (w22258 & ~w8162) | (w22258 & w32229) | (~w8162 & w32229);
assign w22260 = a_50 & ~w22259;
assign w22261 = w22259 & a_50;
assign w22262 = ~w22259 & ~w22260;
assign w22263 = ~w22261 & ~w22262;
assign w22264 = (w22263 & w22253) | (w22263 & w32230) | (w22253 & w32230);
assign w22265 = ~w22253 & w32231;
assign w22266 = ~w22264 & ~w22265;
assign w22267 = ~w22181 & w22266;
assign w22268 = ~w22181 & ~w22267;
assign w22269 = w22266 & ~w22267;
assign w22270 = ~w22268 & ~w22269;
assign w22271 = ~w22180 & ~w22270;
assign w22272 = (w22180 & w22267) | (w22180 & w32232) | (w22267 & w32232);
assign w22273 = ~w22268 & w22272;
assign w22274 = ~w22271 & ~w22273;
assign w22275 = ~w22170 & w22274;
assign w22276 = w22170 & ~w22274;
assign w22277 = ~w22275 & ~w22276;
assign w22278 = ~w22169 & w22277;
assign w22279 = w22169 & ~w22277;
assign w22280 = ~w22278 & ~w22279;
assign w22281 = ~w22159 & w22280;
assign w22282 = w22159 & ~w22280;
assign w22283 = ~w22281 & ~w22282;
assign w22284 = b_59 & w5196;
assign w22285 = w5459 & w32233;
assign w22286 = b_58 & w5191;
assign w22287 = ~w22285 & ~w22286;
assign w22288 = ~w22284 & w22287;
assign w22289 = (w22288 & ~w11169) | (w22288 & w32234) | (~w11169 & w32234);
assign w22290 = a_41 & ~w22289;
assign w22291 = w22289 & a_41;
assign w22292 = ~w22289 & ~w22290;
assign w22293 = ~w22291 & ~w22292;
assign w22294 = w22283 & ~w22293;
assign w22295 = w22283 & ~w22294;
assign w22296 = ~w22283 & ~w22293;
assign w22297 = ~w22295 & ~w22296;
assign w22298 = (~w22111 & ~w22113) | (~w22111 & w32235) | (~w22113 & w32235);
assign w22299 = w22297 & w22298;
assign w22300 = ~w22297 & ~w22298;
assign w22301 = ~w22299 & ~w22300;
assign w22302 = b_62 & w4499;
assign w22303 = w4723 & w32236;
assign w22304 = b_61 & w4494;
assign w22305 = ~w22303 & ~w22304;
assign w22306 = ~w22302 & w22305;
assign w22307 = (w22306 & ~w12273) | (w22306 & w32237) | (~w12273 & w32237);
assign w22308 = a_38 & ~w22307;
assign w22309 = w22307 & a_38;
assign w22310 = ~w22307 & ~w22308;
assign w22311 = ~w22309 & ~w22310;
assign w22312 = w22301 & ~w22311;
assign w22313 = w22301 & ~w22312;
assign w22314 = ~w22301 & ~w22311;
assign w22315 = ~w22313 & ~w22314;
assign w22316 = (w22315 & w22156) | (w22315 & w32238) | (w22156 & w32238);
assign w22317 = ~w22156 & w32239;
assign w22318 = ~w22316 & ~w22317;
assign w22319 = ~w22147 & ~w22318;
assign w22320 = w22147 & w22318;
assign w22321 = ~w22319 & ~w22320;
assign w22322 = (~w13761 & w37740) | (~w13761 & w37741) | (w37740 & w37741);
assign w22323 = (w13761 & w37742) | (w13761 & w37743) | (w37742 & w37743);
assign w22324 = ~w22322 & ~w22323;
assign w22325 = (~w22267 & w22270) | (~w22267 & w32242) | (w22270 & w32242);
assign w22326 = b_54 & w6761;
assign w22327 = w7075 & w32243;
assign w22328 = b_53 & w6756;
assign w22329 = ~w22327 & ~w22328;
assign w22330 = ~w22326 & w22329;
assign w22331 = (w22330 & ~w9134) | (w22330 & w32244) | (~w9134 & w32244);
assign w22332 = a_47 & ~w22331;
assign w22333 = w22331 & a_47;
assign w22334 = ~w22331 & ~w22332;
assign w22335 = ~w22333 & ~w22334;
assign w22336 = ~w22253 & ~w22265;
assign w22337 = w12380 & w32245;
assign w22338 = b_36 & ~w12380;
assign w22339 = ~w22337 & ~w22338;
assign w22340 = a_35 & ~w22197;
assign w22341 = ~a_35 & w22197;
assign w22342 = ~w22340 & ~w22341;
assign w22343 = ~w22339 & ~w22342;
assign w22344 = w22339 & w22342;
assign w22345 = ~w22343 & ~w22344;
assign w22346 = (w22026 & w32246) | (w22026 & w32247) | (w32246 & w32247);
assign w22347 = (~w22026 & w32248) | (~w22026 & w32249) | (w32248 & w32249);
assign w22348 = ~w22346 & ~w22347;
assign w22349 = b_39 & w11620;
assign w22350 = w11969 & w32250;
assign w22351 = b_38 & w11615;
assign w22352 = ~w22350 & ~w22351;
assign w22353 = ~w22349 & w22352;
assign w22354 = (w22353 & ~w4888) | (w22353 & w32251) | (~w4888 & w32251);
assign w22355 = a_62 & ~w22354;
assign w22356 = w22354 & a_62;
assign w22357 = ~w22354 & ~w22355;
assign w22358 = ~w22356 & ~w22357;
assign w22359 = ~w22348 & w22358;
assign w22360 = w22348 & ~w22358;
assign w22361 = ~w22359 & ~w22360;
assign w22362 = b_42 & w10562;
assign w22363 = w10902 & w32252;
assign w22364 = b_41 & w10557;
assign w22365 = ~w22363 & ~w22364;
assign w22366 = ~w22362 & w22365;
assign w22367 = (w22366 & ~w5864) | (w22366 & w25463) | (~w5864 & w25463);
assign w22368 = (w5864 & w25689) | (w5864 & w25690) | (w25689 & w25690);
assign w22369 = (~w5864 & w26036) | (~w5864 & w26037) | (w26036 & w26037);
assign w22370 = ~w22367 & ~w22368;
assign w22371 = ~w22369 & ~w22370;
assign w22372 = w22361 & ~w22371;
assign w22373 = w22371 & w22361;
assign w22374 = ~w22361 & ~w22371;
assign w22375 = ~w22373 & ~w22374;
assign w22376 = (~w22214 & w22217) | (~w22214 & w32253) | (w22217 & w32253);
assign w22377 = ~w22375 & ~w22376;
assign w22378 = ~w22375 & ~w22377;
assign w22379 = w22375 & ~w22376;
assign w22380 = ~w22378 & ~w22379;
assign w22381 = b_45 & w9534;
assign w22382 = w9876 & w32254;
assign w22383 = b_44 & w9529;
assign w22384 = ~w22382 & ~w22383;
assign w22385 = ~w22381 & w22384;
assign w22386 = (w22385 & ~w6682) | (w22385 & w25464) | (~w6682 & w25464);
assign w22387 = (w6682 & w25691) | (w6682 & w25692) | (w25691 & w25692);
assign w22388 = (~w6682 & w26038) | (~w6682 & w26039) | (w26038 & w26039);
assign w22389 = ~w22386 & ~w22387;
assign w22390 = ~w22388 & ~w22389;
assign w22391 = (~w22390 & w22378) | (~w22390 & w32255) | (w22378 & w32255);
assign w22392 = ~w22380 & ~w22391;
assign w22393 = ~w22390 & ~w22391;
assign w22394 = ~w22392 & ~w22393;
assign w22395 = (~w22231 & ~w22233) | (~w22231 & w32256) | (~w22233 & w32256);
assign w22396 = w22394 & w22395;
assign w22397 = ~w22394 & ~w22395;
assign w22398 = ~w22396 & ~w22397;
assign w22399 = b_48 & w8526;
assign w22400 = w8886 & w32257;
assign w22401 = b_47 & w8521;
assign w22402 = ~w22400 & ~w22401;
assign w22403 = ~w22399 & w22402;
assign w22404 = (w22403 & ~w7284) | (w22403 & w25465) | (~w7284 & w25465);
assign w22405 = (w7284 & w25693) | (w7284 & w25694) | (w25693 & w25694);
assign w22406 = (~w7284 & w26040) | (~w7284 & w26041) | (w26040 & w26041);
assign w22407 = ~w22404 & ~w22405;
assign w22408 = ~w22406 & ~w22407;
assign w22409 = w22398 & ~w22408;
assign w22410 = w22398 & ~w22409;
assign w22411 = ~w22398 & ~w22408;
assign w22412 = ~w22410 & ~w22411;
assign w22413 = (~w22237 & ~w22239) | (~w22237 & w32258) | (~w22239 & w32258);
assign w22414 = w22412 & w22413;
assign w22415 = (~w22413 & w22410) | (~w22413 & w32259) | (w22410 & w32259);
assign w22416 = b_51 & w7613;
assign w22417 = w7941 & w32260;
assign w22418 = b_50 & w7608;
assign w22419 = ~w22417 & ~w22418;
assign w22420 = ~w22416 & w22419;
assign w22421 = (w22420 & ~w8186) | (w22420 & w26042) | (~w8186 & w26042);
assign w22422 = (w8186 & w26447) | (w8186 & w26448) | (w26447 & w26448);
assign w22423 = (~w8186 & w32261) | (~w8186 & w32262) | (w32261 & w32262);
assign w22424 = ~w22421 & ~w22422;
assign w22425 = ~w22423 & ~w22424;
assign w22426 = (w22425 & w22414) | (w22425 & w32263) | (w22414 & w32263);
assign w22427 = ~w22414 & w32264;
assign w22428 = ~w22426 & ~w22427;
assign w22429 = ~w22336 & w22428;
assign w22430 = w22336 & ~w22428;
assign w22431 = ~w22429 & ~w22430;
assign w22432 = ~w22335 & w22431;
assign w22433 = w22335 & ~w22431;
assign w22434 = ~w22432 & ~w22433;
assign w22435 = ~w22325 & w22434;
assign w22436 = w22325 & ~w22434;
assign w22437 = ~w22435 & ~w22436;
assign w22438 = b_57 & w5962;
assign w22439 = w6246 & w32265;
assign w22440 = b_56 & w5957;
assign w22441 = ~w22439 & ~w22440;
assign w22442 = ~w22438 & w22441;
assign w22443 = (w22442 & ~w10452) | (w22442 & w32266) | (~w10452 & w32266);
assign w22444 = a_44 & ~w22443;
assign w22445 = w22443 & a_44;
assign w22446 = ~w22443 & ~w22444;
assign w22447 = ~w22445 & ~w22446;
assign w22448 = w22437 & ~w22447;
assign w22449 = w22437 & ~w22448;
assign w22450 = ~w22437 & ~w22447;
assign w22451 = (~w22275 & ~w22277) | (~w22275 & w32267) | (~w22277 & w32267);
assign w22452 = ~w22449 & w27671;
assign w22453 = (~w22451 & w22449) | (~w22451 & w27672) | (w22449 & w27672);
assign w22454 = ~w22452 & ~w22453;
assign w22455 = b_60 & w5196;
assign w22456 = w5459 & w32268;
assign w22457 = b_59 & w5191;
assign w22458 = ~w22456 & ~w22457;
assign w22459 = ~w22455 & w22458;
assign w22460 = (w22459 & ~w11196) | (w22459 & w32269) | (~w11196 & w32269);
assign w22461 = a_41 & ~w22460;
assign w22462 = w22460 & a_41;
assign w22463 = ~w22460 & ~w22461;
assign w22464 = ~w22462 & ~w22463;
assign w22465 = w22454 & ~w22464;
assign w22466 = w22454 & ~w22465;
assign w22467 = ~w22454 & ~w22464;
assign w22468 = ~w22466 & ~w22467;
assign w22469 = (~w22281 & ~w22283) | (~w22281 & w32270) | (~w22283 & w32270);
assign w22470 = w22468 & w22469;
assign w22471 = ~w22468 & ~w22469;
assign w22472 = ~w22470 & ~w22471;
assign w22473 = b_63 & w4499;
assign w22474 = w4723 & w32271;
assign w22475 = b_62 & w4494;
assign w22476 = ~w22474 & ~w22475;
assign w22477 = ~w22473 & w22476;
assign w22478 = (w22477 & ~w12646) | (w22477 & w32272) | (~w12646 & w32272);
assign w22479 = a_38 & ~w22478;
assign w22480 = w22478 & a_38;
assign w22481 = ~w22478 & ~w22479;
assign w22482 = ~w22480 & ~w22481;
assign w22483 = w22472 & ~w22482;
assign w22484 = w22472 & ~w22483;
assign w22485 = ~w22472 & ~w22482;
assign w22486 = ~w22484 & ~w22485;
assign w22487 = (~w22300 & ~w22301) | (~w22300 & w32273) | (~w22301 & w32273);
assign w22488 = w22486 & w22487;
assign w22489 = ~w22486 & ~w22487;
assign w22490 = ~w22488 & ~w22489;
assign w22491 = (~w22315 & w22156) | (~w22315 & w32274) | (w22156 & w32274);
assign w22492 = (w22490 & w22491) | (w22490 & w32275) | (w22491 & w32275);
assign w22493 = ~w22491 & w32276;
assign w22494 = ~w22492 & ~w22493;
assign w22495 = (~w13761 & w37744) | (~w13761 & w37745) | (w37744 & w37745);
assign w22496 = (w13761 & w37746) | (w13761 & w37747) | (w37746 & w37747);
assign w22497 = ~w22495 & ~w22496;
assign w22498 = (~w22465 & w22468) | (~w22465 & w32277) | (w22468 & w32277);
assign w22499 = w4723 & w32278;
assign w22500 = b_63 & w4494;
assign w22501 = ~w22499 & ~w22500;
assign w22502 = ~w12671 & w32279;
assign w22503 = (a_38 & w22502) | (a_38 & w32280) | (w22502 & w32280);
assign w22504 = ~w22502 & w32281;
assign w22505 = ~w22503 & ~w22504;
assign w22506 = ~w22498 & ~w22505;
assign w22507 = w22498 & w22505;
assign w22508 = ~w22506 & ~w22507;
assign w22509 = b_40 & w11620;
assign w22510 = w11969 & w32282;
assign w22511 = b_39 & w11615;
assign w22512 = ~w22510 & ~w22511;
assign w22513 = ~w22509 & w22512;
assign w22514 = (w22513 & ~w5363) | (w22513 & w25695) | (~w5363 & w25695);
assign w22515 = (w5363 & w26043) | (w5363 & w26044) | (w26043 & w26044);
assign w22516 = (~w5363 & w32283) | (~w5363 & w32284) | (w32283 & w32284);
assign w22517 = ~w22514 & ~w22515;
assign w22518 = ~w22516 & ~w22517;
assign w22519 = w12380 & w32285;
assign w22520 = b_37 & ~w12380;
assign w22521 = ~w22519 & ~w22520;
assign w22522 = ~a_35 & ~w22197;
assign w22523 = (~w22522 & w22342) | (~w22522 & w32286) | (w22342 & w32286);
assign w22524 = w22521 & ~w22523;
assign w22525 = w22523 & w22521;
assign w22526 = ~w22523 & ~w22524;
assign w22527 = ~w22525 & ~w22526;
assign w22528 = (~w22527 & w22517) | (~w22527 & w32287) | (w22517 & w32287);
assign w22529 = ~w22518 & ~w22528;
assign w22530 = ~w22527 & ~w22528;
assign w22531 = ~w22529 & ~w22530;
assign w22532 = ~w22346 & ~w22360;
assign w22533 = w22531 & w22532;
assign w22534 = ~w22531 & ~w22532;
assign w22535 = ~w22533 & ~w22534;
assign w22536 = b_43 & w10562;
assign w22537 = w10902 & w32288;
assign w22538 = b_42 & w10557;
assign w22539 = ~w22537 & ~w22538;
assign w22540 = ~w22536 & w22539;
assign w22541 = (w22540 & ~w5888) | (w22540 & w25696) | (~w5888 & w25696);
assign w22542 = (w5888 & w26045) | (w5888 & w26046) | (w26045 & w26046);
assign w22543 = (~w5888 & w32289) | (~w5888 & w32290) | (w32289 & w32290);
assign w22544 = ~w22541 & ~w22542;
assign w22545 = ~w22543 & ~w22544;
assign w22546 = w22535 & ~w22545;
assign w22547 = w22535 & ~w22546;
assign w22548 = ~w22535 & ~w22545;
assign w22549 = ~w22547 & ~w22548;
assign w22550 = ~w22372 & ~w22377;
assign w22551 = w22549 & w22550;
assign w22552 = ~w22549 & ~w22550;
assign w22553 = ~w22551 & ~w22552;
assign w22554 = b_46 & w9534;
assign w22555 = w9876 & w32291;
assign w22556 = b_45 & w9529;
assign w22557 = ~w22555 & ~w22556;
assign w22558 = ~w22554 & w22557;
assign w22559 = (w22558 & ~w6974) | (w22558 & w25466) | (~w6974 & w25466);
assign w22560 = (w6974 & w25697) | (w6974 & w25698) | (w25697 & w25698);
assign w22561 = (~w6974 & w26047) | (~w6974 & w26048) | (w26047 & w26048);
assign w22562 = ~w22559 & ~w22560;
assign w22563 = ~w22561 & ~w22562;
assign w22564 = w22563 & w22553;
assign w22565 = ~w22553 & ~w22563;
assign w22566 = ~w22564 & ~w22565;
assign w22567 = (~w22391 & w22394) | (~w22391 & w26049) | (w22394 & w26049);
assign w22568 = w22566 & w22567;
assign w22569 = ~w22566 & ~w22567;
assign w22570 = ~w22568 & ~w22569;
assign w22571 = b_49 & w8526;
assign w22572 = w8886 & w32292;
assign w22573 = b_48 & w8521;
assign w22574 = ~w22572 & ~w22573;
assign w22575 = ~w22571 & w22574;
assign w22576 = (w22575 & ~w7859) | (w22575 & w25467) | (~w7859 & w25467);
assign w22577 = (w7859 & w25699) | (w7859 & w25700) | (w25699 & w25700);
assign w22578 = (~w7859 & w26050) | (~w7859 & w26051) | (w26050 & w26051);
assign w22579 = ~w22576 & ~w22577;
assign w22580 = ~w22578 & ~w22579;
assign w22581 = w22570 & ~w22580;
assign w22582 = w22570 & ~w22581;
assign w22583 = ~w22570 & ~w22580;
assign w22584 = ~w22582 & ~w22583;
assign w22585 = (~w22409 & w22412) | (~w22409 & w26052) | (w22412 & w26052);
assign w22586 = w22584 & w22585;
assign w22587 = ~w22584 & ~w22585;
assign w22588 = ~w22586 & ~w22587;
assign w22589 = b_52 & w7613;
assign w22590 = w7941 & w32293;
assign w22591 = b_51 & w7608;
assign w22592 = ~w22590 & ~w22591;
assign w22593 = ~w22589 & w22592;
assign w22594 = (w22593 & ~w8793) | (w22593 & w25701) | (~w8793 & w25701);
assign w22595 = (w8793 & w26053) | (w8793 & w26054) | (w26053 & w26054);
assign w22596 = (~w8793 & w32294) | (~w8793 & w32295) | (w32294 & w32295);
assign w22597 = ~w22594 & ~w22595;
assign w22598 = ~w22596 & ~w22597;
assign w22599 = w22588 & ~w22598;
assign w22600 = w22588 & ~w22599;
assign w22601 = ~w22588 & ~w22598;
assign w22602 = ~w22600 & ~w22601;
assign w22603 = (~w22427 & w22336) | (~w22427 & w32296) | (w22336 & w32296);
assign w22604 = (~w22603 & w22600) | (~w22603 & w26449) | (w22600 & w26449);
assign w22605 = ~w22602 & ~w22604;
assign w22606 = ~w22600 & w26717;
assign w22607 = ~w22605 & ~w22606;
assign w22608 = b_55 & w6761;
assign w22609 = w7075 & w32297;
assign w22610 = b_54 & w6756;
assign w22611 = ~w22609 & ~w22610;
assign w22612 = ~w22608 & w22611;
assign w22613 = (w22612 & ~w9776) | (w22612 & w26450) | (~w9776 & w26450);
assign w22614 = (w9776 & w32298) | (w9776 & w32299) | (w32298 & w32299);
assign w22615 = (~w9776 & w32300) | (~w9776 & w32301) | (w32300 & w32301);
assign w22616 = ~w22613 & ~w22614;
assign w22617 = ~w22615 & ~w22616;
assign w22618 = (~w22617 & w22605) | (~w22617 & w26055) | (w22605 & w26055);
assign w22619 = ~w22607 & ~w22618;
assign w22620 = ~w26055 & w26451;
assign w22621 = ~w22619 & ~w22620;
assign w22622 = ~w22432 & ~w22435;
assign w22623 = w22621 & w22622;
assign w22624 = ~w22621 & ~w22622;
assign w22625 = ~w22623 & ~w22624;
assign w22626 = b_58 & w5962;
assign w22627 = w6246 & w32302;
assign w22628 = b_57 & w5957;
assign w22629 = ~w22627 & ~w22628;
assign w22630 = ~w22626 & w22629;
assign w22631 = (w22630 & ~w10476) | (w22630 & w32303) | (~w10476 & w32303);
assign w22632 = a_44 & ~w22631;
assign w22633 = w22631 & a_44;
assign w22634 = ~w22631 & ~w22632;
assign w22635 = ~w22633 & ~w22634;
assign w22636 = w22625 & ~w22635;
assign w22637 = w22625 & ~w22636;
assign w22638 = ~w22625 & ~w22635;
assign w22639 = (~w27672 & w32304) | (~w27672 & w32305) | (w32304 & w32305);
assign w22640 = ~w22637 & w27673;
assign w22641 = (~w22639 & w22637) | (~w22639 & w27674) | (w22637 & w27674);
assign w22642 = ~w22640 & ~w22641;
assign w22643 = b_61 & w5196;
assign w22644 = w5459 & w32306;
assign w22645 = b_60 & w5191;
assign w22646 = ~w22644 & ~w22645;
assign w22647 = ~w22643 & w22646;
assign w22648 = (w22647 & ~w11901) | (w22647 & w32307) | (~w11901 & w32307);
assign w22649 = a_41 & ~w22648;
assign w22650 = w22648 & a_41;
assign w22651 = ~w22648 & ~w22649;
assign w22652 = ~w22650 & ~w22651;
assign w22653 = w22642 & ~w22652;
assign w22654 = ~w22642 & w22652;
assign w22655 = w22508 & w32308;
assign w22656 = w22508 & ~w22655;
assign w22657 = w32308 & ~w22508;
assign w22658 = ~w22656 & ~w22657;
assign w22659 = (~w22483 & w22486) | (~w22483 & w32309) | (w22486 & w32309);
assign w22660 = w22658 & w22659;
assign w22661 = ~w22658 & ~w22659;
assign w22662 = ~w22660 & ~w22661;
assign w22663 = (~w13761 & w37748) | (~w13761 & w37749) | (w37748 & w37749);
assign w22664 = (w13761 & w37750) | (w13761 & w37751) | (w37750 & w37751);
assign w22665 = ~w22663 & ~w22664;
assign w22666 = (~w22506 & ~w22508) | (~w22506 & w32314) | (~w22508 & w32314);
assign w22667 = (~w22641 & ~w22642) | (~w22641 & w26452) | (~w22642 & w26452);
assign w22668 = w4723 & w32315;
assign w22669 = (~w22668 & ~w12670) | (~w22668 & w32316) | (~w12670 & w32316);
assign w22670 = a_38 & ~w22669;
assign w22671 = w22669 & a_38;
assign w22672 = ~w22669 & ~w22670;
assign w22673 = ~w22671 & ~w22672;
assign w22674 = ~w22667 & ~w22673;
assign w22675 = ~w22667 & ~w22674;
assign w22676 = w22667 & ~w22673;
assign w22677 = ~w22675 & ~w22676;
assign w22678 = ~w22604 & ~w22618;
assign w22679 = b_56 & w6761;
assign w22680 = w7075 & w32317;
assign w22681 = b_55 & w6756;
assign w22682 = ~w22680 & ~w22681;
assign w22683 = ~w22679 & w22682;
assign w22684 = (w22683 & ~w9798) | (w22683 & w32318) | (~w9798 & w32318);
assign w22685 = a_47 & ~w22684;
assign w22686 = w22684 & a_47;
assign w22687 = ~w22684 & ~w22685;
assign w22688 = ~w22686 & ~w22687;
assign w22689 = (~w22587 & ~w22588) | (~w22587 & w32319) | (~w22588 & w32319);
assign w22690 = b_53 & w7613;
assign w22691 = w7941 & w32320;
assign w22692 = b_52 & w7608;
assign w22693 = ~w22691 & ~w22692;
assign w22694 = ~w22690 & w22693;
assign w22695 = (w22694 & ~w9110) | (w22694 & w32321) | (~w9110 & w32321);
assign w22696 = a_50 & ~w22695;
assign w22697 = w22695 & a_50;
assign w22698 = ~w22695 & ~w22696;
assign w22699 = ~w22697 & ~w22698;
assign w22700 = (~w22569 & ~w22570) | (~w22569 & w32322) | (~w22570 & w32322);
assign w22701 = ~w22524 & ~w22528;
assign w22702 = w12380 & w32323;
assign w22703 = b_38 & ~w12380;
assign w22704 = ~w22702 & ~w22703;
assign w22705 = w22521 & ~w22704;
assign w22706 = w22521 & ~w22705;
assign w22707 = ~w22704 & ~w22705;
assign w22708 = ~w22706 & ~w22707;
assign w22709 = (~w22708 & w22528) | (~w22708 & w32324) | (w22528 & w32324);
assign w22710 = ~w22701 & ~w22709;
assign w22711 = ~w22528 & w32325;
assign w22712 = ~w22710 & ~w22711;
assign w22713 = b_41 & w11620;
assign w22714 = w11969 & w32326;
assign w22715 = b_40 & w11615;
assign w22716 = ~w22714 & ~w22715;
assign w22717 = ~w22713 & w22716;
assign w22718 = (w22717 & ~w5609) | (w22717 & w32327) | (~w5609 & w32327);
assign w22719 = a_62 & ~w22718;
assign w22720 = w22718 & a_62;
assign w22721 = ~w22718 & ~w22719;
assign w22722 = ~w22720 & ~w22721;
assign w22723 = (~w22722 & w22710) | (~w22722 & w32328) | (w22710 & w32328);
assign w22724 = ~w22712 & ~w22723;
assign w22725 = ~w22722 & ~w22723;
assign w22726 = ~w22724 & ~w22725;
assign w22727 = b_44 & w10562;
assign w22728 = w10902 & w32329;
assign w22729 = b_43 & w10557;
assign w22730 = ~w22728 & ~w22729;
assign w22731 = ~w22727 & w22730;
assign w22732 = (w22731 & ~w6408) | (w22731 & w26453) | (~w6408 & w26453);
assign w22733 = (w6408 & w27675) | (w6408 & w27676) | (w27675 & w27676);
assign w22734 = (~w6408 & w32330) | (~w6408 & w32331) | (w32330 & w32331);
assign w22735 = ~w22732 & ~w22733;
assign w22736 = ~w22734 & ~w22735;
assign w22737 = ~w22726 & w22736;
assign w22738 = w22726 & ~w22736;
assign w22739 = ~w22737 & ~w22738;
assign w22740 = (~w22534 & ~w22535) | (~w22534 & w32332) | (~w22535 & w32332);
assign w22741 = w22739 & w22740;
assign w22742 = ~w22739 & ~w22740;
assign w22743 = ~w22741 & ~w22742;
assign w22744 = b_47 & w9534;
assign w22745 = w9876 & w32333;
assign w22746 = b_46 & w9529;
assign w22747 = ~w22745 & ~w22746;
assign w22748 = ~w22744 & w22747;
assign w22749 = (w22748 & ~w6998) | (w22748 & w25702) | (~w6998 & w25702);
assign w22750 = (w6998 & w26056) | (w6998 & w26057) | (w26056 & w26057);
assign w22751 = (~w6998 & w26454) | (~w6998 & w26455) | (w26454 & w26455);
assign w22752 = ~w22749 & ~w22750;
assign w22753 = ~w22751 & ~w22752;
assign w22754 = w22743 & w22753;
assign w22755 = (~w27677 & w32334) | (~w27677 & w32335) | (w32334 & w32335);
assign w22756 = (~w22552 & ~w22553) | (~w22552 & w32336) | (~w22553 & w32336);
assign w22757 = ~w22755 & w26456;
assign w22758 = (~w22756 & w22755) | (~w22756 & w26457) | (w22755 & w26457);
assign w22759 = ~w22757 & ~w22758;
assign w22760 = b_50 & w8526;
assign w22761 = w8886 & w32337;
assign w22762 = b_49 & w8521;
assign w22763 = ~w22761 & ~w22762;
assign w22764 = ~w22760 & w22763;
assign w22765 = (w22764 & ~w8162) | (w22764 & w26458) | (~w8162 & w26458);
assign w22766 = (w8162 & w32338) | (w8162 & w32339) | (w32338 & w32339);
assign w22767 = (~w8162 & w32340) | (~w8162 & w32341) | (w32340 & w32341);
assign w22768 = ~w22765 & ~w22766;
assign w22769 = ~w22767 & ~w22768;
assign w22770 = ~w22759 & w22769;
assign w22771 = w22759 & ~w22769;
assign w22772 = ~w22770 & ~w22771;
assign w22773 = ~w22700 & w22772;
assign w22774 = ~w22772 & ~w22700;
assign w22775 = w22772 & ~w22773;
assign w22776 = (~w22699 & w22775) | (~w22699 & w32342) | (w22775 & w32342);
assign w22777 = ~w22775 & w32343;
assign w22778 = ~w22776 & ~w22777;
assign w22779 = ~w22689 & w22778;
assign w22780 = w22689 & ~w22778;
assign w22781 = ~w22779 & ~w22780;
assign w22782 = ~w22688 & w22781;
assign w22783 = w22688 & ~w22781;
assign w22784 = ~w22782 & ~w22783;
assign w22785 = ~w22678 & w22784;
assign w22786 = w22678 & ~w22784;
assign w22787 = ~w22785 & ~w22786;
assign w22788 = b_59 & w5962;
assign w22789 = w6246 & w32344;
assign w22790 = b_58 & w5957;
assign w22791 = ~w22789 & ~w22790;
assign w22792 = ~w22788 & w22791;
assign w22793 = (w22792 & ~w11169) | (w22792 & w32345) | (~w11169 & w32345);
assign w22794 = a_44 & ~w22793;
assign w22795 = w22793 & a_44;
assign w22796 = ~w22793 & ~w22794;
assign w22797 = ~w22795 & ~w22796;
assign w22798 = w22787 & ~w22797;
assign w22799 = w22787 & ~w22798;
assign w22800 = ~w22787 & ~w22797;
assign w22801 = ~w22799 & ~w22800;
assign w22802 = (~w22624 & ~w22625) | (~w22624 & w32346) | (~w22625 & w32346);
assign w22803 = w22801 & w22802;
assign w22804 = ~w22801 & ~w22802;
assign w22805 = ~w22803 & ~w22804;
assign w22806 = b_62 & w5196;
assign w22807 = w5459 & w32347;
assign w22808 = b_61 & w5191;
assign w22809 = ~w22807 & ~w22808;
assign w22810 = ~w22806 & w22809;
assign w22811 = (w22810 & ~w12273) | (w22810 & w32348) | (~w12273 & w32348);
assign w22812 = a_41 & ~w22811;
assign w22813 = w22811 & a_41;
assign w22814 = ~w22811 & ~w22812;
assign w22815 = ~w22813 & ~w22814;
assign w22816 = w22805 & ~w22815;
assign w22817 = w22805 & ~w22816;
assign w22818 = ~w22805 & ~w22815;
assign w22819 = ~w22817 & ~w22818;
assign w22820 = ~w22677 & w22819;
assign w22821 = w22677 & ~w22819;
assign w22822 = ~w22820 & ~w22821;
assign w22823 = ~w22666 & ~w22822;
assign w22824 = w22666 & w22822;
assign w22825 = ~w22823 & ~w22824;
assign w22826 = (~w13761 & w37752) | (~w13761 & w37753) | (w37752 & w37753);
assign w22827 = (w13761 & w37754) | (w13761 & w37755) | (w37754 & w37755);
assign w22828 = ~w22826 & ~w22827;
assign w22829 = ~w22773 & ~w22776;
assign w22830 = b_54 & w7613;
assign w22831 = w7941 & w32351;
assign w22832 = b_53 & w7608;
assign w22833 = ~w22831 & ~w22832;
assign w22834 = ~w22830 & w22833;
assign w22835 = (w22834 & ~w9134) | (w22834 & w26058) | (~w9134 & w26058);
assign w22836 = (w9134 & w26459) | (w9134 & w26460) | (w26459 & w26460);
assign w22837 = (~w9134 & w32352) | (~w9134 & w32353) | (w32352 & w32353);
assign w22838 = ~w22835 & ~w22836;
assign w22839 = ~w22837 & ~w22838;
assign w22840 = (~w22758 & ~w22759) | (~w22758 & w32354) | (~w22759 & w32354);
assign w22841 = w12380 & w32357;
assign w22842 = b_39 & ~w12380;
assign w22843 = ~w22841 & ~w22842;
assign w22844 = a_38 & ~w22521;
assign w22845 = ~a_38 & w22521;
assign w22846 = ~w22844 & ~w22845;
assign w22847 = ~w22843 & ~w22846;
assign w22848 = w22843 & w22846;
assign w22849 = ~w22847 & ~w22848;
assign w22850 = (w22528 & w32358) | (w22528 & w32359) | (w32358 & w32359);
assign w22851 = (~w22528 & w32360) | (~w22528 & w32361) | (w32360 & w32361);
assign w22852 = ~w22850 & ~w22851;
assign w22853 = b_42 & w11620;
assign w22854 = w11969 & w32362;
assign w22855 = b_41 & w11615;
assign w22856 = ~w22854 & ~w22855;
assign w22857 = ~w22853 & w22856;
assign w22858 = (w22857 & ~w5864) | (w22857 & w32363) | (~w5864 & w32363);
assign w22859 = a_62 & ~w22858;
assign w22860 = w22858 & a_62;
assign w22861 = ~w22858 & ~w22859;
assign w22862 = ~w22860 & ~w22861;
assign w22863 = w22852 & ~w22862;
assign w22864 = w22852 & ~w22863;
assign w22865 = ~w22852 & ~w22862;
assign w22866 = b_45 & w10562;
assign w22867 = w10902 & w32364;
assign w22868 = b_44 & w10557;
assign w22869 = ~w22867 & ~w22868;
assign w22870 = ~w22866 & w22869;
assign w22871 = (w22870 & ~w6682) | (w22870 & w25468) | (~w6682 & w25468);
assign w22872 = (w6682 & w25703) | (w6682 & w25704) | (w25703 & w25704);
assign w22873 = (~w6682 & w26059) | (~w6682 & w26060) | (w26059 & w26060);
assign w22874 = ~w22871 & ~w22872;
assign w22875 = ~w22873 & ~w22874;
assign w22876 = (~w22875 & w22864) | (~w22875 & w32365) | (w22864 & w32365);
assign w22877 = (w22875 & w22864) | (w22875 & w32366) | (w22864 & w32366);
assign w22878 = ~w22875 & ~w22876;
assign w22879 = ~w22877 & ~w22878;
assign w22880 = (~w22723 & w22726) | (~w22723 & w32367) | (w22726 & w32367);
assign w22881 = (~w22880 & w22878) | (~w22880 & w26461) | (w22878 & w26461);
assign w22882 = ~w22879 & ~w22881;
assign w22883 = ~w22878 & w27678;
assign w22884 = ~w22882 & ~w22883;
assign w22885 = b_48 & w9534;
assign w22886 = w9876 & w32368;
assign w22887 = b_47 & w9529;
assign w22888 = ~w22886 & ~w22887;
assign w22889 = ~w22885 & w22888;
assign w22890 = (w22889 & ~w7284) | (w22889 & w25705) | (~w7284 & w25705);
assign w22891 = (w7284 & w26061) | (w7284 & w26062) | (w26061 & w26062);
assign w22892 = (~w7284 & w26462) | (~w7284 & w26463) | (w26462 & w26463);
assign w22893 = ~w22890 & ~w22891;
assign w22894 = ~w22892 & ~w22893;
assign w22895 = (~w22894 & w22882) | (~w22894 & w32369) | (w22882 & w32369);
assign w22896 = ~w22884 & ~w22895;
assign w22897 = ~w22882 & w32370;
assign w22898 = (~w27677 & w32371) | (~w27677 & w32372) | (w32371 & w32372);
assign w22899 = ~w22896 & w26063;
assign w22900 = (~w22898 & w22896) | (~w22898 & w26064) | (w22896 & w26064);
assign w22901 = ~w22899 & ~w22900;
assign w22902 = b_51 & w8526;
assign w22903 = w8886 & w32373;
assign w22904 = b_50 & w8521;
assign w22905 = ~w22903 & ~w22904;
assign w22906 = ~w22902 & w22905;
assign w22907 = (w22906 & ~w8186) | (w22906 & w26065) | (~w8186 & w26065);
assign w22908 = (w8186 & w26464) | (w8186 & w26465) | (w26464 & w26465);
assign w22909 = (~w8186 & w32374) | (~w8186 & w32375) | (w32374 & w32375);
assign w22910 = ~w22907 & ~w22908;
assign w22911 = ~w22909 & ~w22910;
assign w22912 = ~w22901 & w22911;
assign w22913 = w22901 & ~w22911;
assign w22914 = ~w22912 & ~w22913;
assign w22915 = ~w22840 & w22914;
assign w22916 = w22840 & ~w22914;
assign w22917 = ~w22915 & ~w22916;
assign w22918 = ~w22839 & w22917;
assign w22919 = w22839 & ~w22917;
assign w22920 = ~w22918 & ~w22919;
assign w22921 = ~w22829 & w22920;
assign w22922 = w22829 & ~w22920;
assign w22923 = ~w22921 & ~w22922;
assign w22924 = b_57 & w6761;
assign w22925 = w7075 & w32376;
assign w22926 = b_56 & w6756;
assign w22927 = ~w22925 & ~w22926;
assign w22928 = ~w22924 & w22927;
assign w22929 = (w22928 & ~w10452) | (w22928 & w26466) | (~w10452 & w26466);
assign w22930 = (w10452 & w32377) | (w10452 & w32378) | (w32377 & w32378);
assign w22931 = (~w10452 & w32379) | (~w10452 & w32380) | (w32379 & w32380);
assign w22932 = ~w22929 & ~w22930;
assign w22933 = ~w22931 & ~w22932;
assign w22934 = w22923 & ~w22933;
assign w22935 = w22923 & ~w22934;
assign w22936 = ~w22923 & ~w22933;
assign w22937 = (~w22779 & ~w22781) | (~w22779 & w32381) | (~w22781 & w32381);
assign w22938 = ~w22935 & w27679;
assign w22939 = (~w22937 & w22935) | (~w22937 & w27680) | (w22935 & w27680);
assign w22940 = ~w22938 & ~w22939;
assign w22941 = b_60 & w5962;
assign w22942 = w6246 & w32382;
assign w22943 = b_59 & w5957;
assign w22944 = ~w22942 & ~w22943;
assign w22945 = ~w22941 & w22944;
assign w22946 = (w22945 & ~w11196) | (w22945 & w32383) | (~w11196 & w32383);
assign w22947 = a_44 & ~w22946;
assign w22948 = w22946 & a_44;
assign w22949 = ~w22946 & ~w22947;
assign w22950 = ~w22948 & ~w22949;
assign w22951 = w22940 & ~w22950;
assign w22952 = w22940 & ~w22951;
assign w22953 = ~w22940 & ~w22950;
assign w22954 = ~w22952 & ~w22953;
assign w22955 = (~w22785 & ~w22787) | (~w22785 & w32384) | (~w22787 & w32384);
assign w22956 = w22954 & w22955;
assign w22957 = (~w22955 & w22952) | (~w22955 & w26467) | (w22952 & w26467);
assign w22958 = ~w22956 & ~w22957;
assign w22959 = b_63 & w5196;
assign w22960 = w5459 & w32385;
assign w22961 = b_62 & w5191;
assign w22962 = ~w22960 & ~w22961;
assign w22963 = ~w22959 & w22962;
assign w22964 = (w22963 & ~w12646) | (w22963 & w32386) | (~w12646 & w32386);
assign w22965 = a_41 & ~w22964;
assign w22966 = w22964 & a_41;
assign w22967 = ~w22964 & ~w22965;
assign w22968 = ~w22966 & ~w22967;
assign w22969 = w22958 & ~w22968;
assign w22970 = w22958 & ~w22969;
assign w22971 = ~w22958 & ~w22968;
assign w22972 = ~w22970 & ~w22971;
assign w22973 = (~w22804 & ~w22805) | (~w22804 & w32387) | (~w22805 & w32387);
assign w22974 = w22972 & w22973;
assign w22975 = ~w22972 & ~w22973;
assign w22976 = ~w22974 & ~w22975;
assign w22977 = (~w22674 & w22677) | (~w22674 & w32388) | (w22677 & w32388);
assign w22978 = w22976 & ~w22977;
assign w22979 = ~w22976 & w22977;
assign w22980 = ~w22978 & ~w22979;
assign w22981 = (~w13761 & w37756) | (~w13761 & w37757) | (w37756 & w37757);
assign w22982 = (w13761 & w37758) | (w13761 & w37759) | (w37758 & w37759);
assign w22983 = ~w22981 & ~w22982;
assign w22984 = (~w26467 & w32389) | (~w26467 & w32390) | (w32389 & w32390);
assign w22985 = w5459 & w32391;
assign w22986 = b_63 & w5191;
assign w22987 = ~w22985 & ~w22986;
assign w22988 = ~w12671 & w32392;
assign w22989 = (a_41 & w22988) | (a_41 & w32393) | (w22988 & w32393);
assign w22990 = ~w22988 & w32394;
assign w22991 = ~w22989 & ~w22990;
assign w22992 = ~w22984 & ~w22991;
assign w22993 = w22984 & w22991;
assign w22994 = ~w22992 & ~w22993;
assign w22995 = (~w22850 & ~w22852) | (~w22850 & w32395) | (~w22852 & w32395);
assign w22996 = w12380 & w32396;
assign w22997 = b_40 & ~w12380;
assign w22998 = ~w22996 & ~w22997;
assign w22999 = ~a_38 & ~w22521;
assign w23000 = (~w22999 & w22846) | (~w22999 & w32397) | (w22846 & w32397);
assign w23001 = w22998 & ~w23000;
assign w23002 = ~w22998 & w23000;
assign w23003 = ~w23001 & ~w23002;
assign w23004 = b_43 & w11620;
assign w23005 = w11969 & w32398;
assign w23006 = b_42 & w11615;
assign w23007 = ~w23005 & ~w23006;
assign w23008 = ~w23004 & w23007;
assign w23009 = w23007 & w32399;
assign w23010 = (~w23009 & w5888) | (~w23009 & w32400) | (w5888 & w32400);
assign w23011 = a_62 & ~w23010;
assign w23012 = (w23003 & w23011) | (w23003 & w32403) | (w23011 & w32403);
assign w23013 = ~w23011 & w32404;
assign w23014 = ~w23012 & ~w23013;
assign w23015 = ~w22995 & w23014;
assign w23016 = w22995 & ~w23014;
assign w23017 = ~w23015 & ~w23016;
assign w23018 = b_46 & w10562;
assign w23019 = w10902 & w32405;
assign w23020 = b_45 & w10557;
assign w23021 = ~w23019 & ~w23020;
assign w23022 = ~w23018 & w23021;
assign w23023 = (w23022 & ~w6974) | (w23022 & w25706) | (~w6974 & w25706);
assign w23024 = (w6974 & w26066) | (w6974 & w26067) | (w26066 & w26067);
assign w23025 = (~w6974 & w26468) | (~w6974 & w26469) | (w26468 & w26469);
assign w23026 = ~w23023 & ~w23024;
assign w23027 = ~w23025 & ~w23026;
assign w23028 = w23027 & w23017;
assign w23029 = ~w23017 & ~w23027;
assign w23030 = ~w23028 & ~w23029;
assign w23031 = (~w26461 & w32406) | (~w26461 & w32407) | (w32406 & w32407);
assign w23032 = w23030 & w23031;
assign w23033 = ~w23030 & ~w23031;
assign w23034 = ~w23032 & ~w23033;
assign w23035 = b_49 & w9534;
assign w23036 = w9876 & w32408;
assign w23037 = b_48 & w9529;
assign w23038 = ~w23036 & ~w23037;
assign w23039 = ~w23035 & w23038;
assign w23040 = (w23039 & ~w7859) | (w23039 & w25707) | (~w7859 & w25707);
assign w23041 = (w7859 & w26068) | (w7859 & w26069) | (w26068 & w26069);
assign w23042 = (~w7859 & w26470) | (~w7859 & w26471) | (w26470 & w26471);
assign w23043 = ~w23040 & ~w23041;
assign w23044 = ~w23042 & ~w23043;
assign w23045 = w23034 & ~w23044;
assign w23046 = w23034 & ~w23045;
assign w23047 = ~w23034 & ~w23044;
assign w23048 = ~w23046 & ~w23047;
assign w23049 = (~w26064 & w26472) | (~w26064 & w26473) | (w26472 & w26473);
assign w23050 = w23048 & w23049;
assign w23051 = ~w23048 & ~w23049;
assign w23052 = ~w23050 & ~w23051;
assign w23053 = b_52 & w8526;
assign w23054 = w8886 & w32409;
assign w23055 = b_51 & w8521;
assign w23056 = ~w23054 & ~w23055;
assign w23057 = ~w23053 & w23056;
assign w23058 = (w23057 & ~w8793) | (w23057 & w26070) | (~w8793 & w26070);
assign w23059 = (w8793 & w26474) | (w8793 & w26475) | (w26474 & w26475);
assign w23060 = (~w8793 & w32410) | (~w8793 & w32411) | (w32410 & w32411);
assign w23061 = ~w23058 & ~w23059;
assign w23062 = ~w23060 & ~w23061;
assign w23063 = w23052 & ~w23062;
assign w23064 = w23052 & ~w23063;
assign w23065 = ~w23052 & ~w23062;
assign w23066 = ~w23064 & ~w23065;
assign w23067 = (~w22913 & ~w22914) | (~w22913 & w27681) | (~w22914 & w27681);
assign w23068 = (~w23067 & w23064) | (~w23067 & w26720) | (w23064 & w26720);
assign w23069 = ~w23066 & ~w23068;
assign w23070 = ~w23064 & w26721;
assign w23071 = ~w23069 & ~w23070;
assign w23072 = b_55 & w7613;
assign w23073 = w7941 & w32412;
assign w23074 = b_54 & w7608;
assign w23075 = ~w23073 & ~w23074;
assign w23076 = ~w23072 & w23075;
assign w23077 = (w23076 & ~w9776) | (w23076 & w32413) | (~w9776 & w32413);
assign w23078 = a_50 & ~w23077;
assign w23079 = w23077 & a_50;
assign w23080 = ~w23077 & ~w23078;
assign w23081 = ~w23079 & ~w23080;
assign w23082 = (~w23081 & w23069) | (~w23081 & w26476) | (w23069 & w26476);
assign w23083 = ~w23071 & ~w23082;
assign w23084 = ~w23081 & ~w23082;
assign w23085 = ~w23083 & ~w23084;
assign w23086 = ~w22918 & ~w22921;
assign w23087 = w23085 & w23086;
assign w23088 = ~w23085 & ~w23086;
assign w23089 = ~w23087 & ~w23088;
assign w23090 = b_58 & w6761;
assign w23091 = w7075 & w32414;
assign w23092 = b_57 & w6756;
assign w23093 = ~w23091 & ~w23092;
assign w23094 = ~w23090 & w23093;
assign w23095 = (w23094 & ~w10476) | (w23094 & w32415) | (~w10476 & w32415);
assign w23096 = a_47 & ~w23095;
assign w23097 = w23095 & a_47;
assign w23098 = ~w23095 & ~w23096;
assign w23099 = ~w23097 & ~w23098;
assign w23100 = w23089 & ~w23099;
assign w23101 = w23089 & ~w23100;
assign w23102 = ~w23089 & ~w23099;
assign w23103 = ~w22934 & ~w22939;
assign w23104 = ~w23101 & w27682;
assign w23105 = (~w23103 & w23101) | (~w23103 & w27683) | (w23101 & w27683);
assign w23106 = ~w23104 & ~w23105;
assign w23107 = b_61 & w5962;
assign w23108 = w6246 & w32416;
assign w23109 = b_60 & w5957;
assign w23110 = ~w23108 & ~w23109;
assign w23111 = ~w23107 & w23110;
assign w23112 = (w23111 & ~w11901) | (w23111 & w32417) | (~w11901 & w32417);
assign w23113 = a_44 & ~w23112;
assign w23114 = w23112 & a_44;
assign w23115 = ~w23112 & ~w23113;
assign w23116 = ~w23114 & ~w23115;
assign w23117 = w23106 & ~w23116;
assign w23118 = ~w23106 & w23116;
assign w23119 = w22994 & w32418;
assign w23120 = w22994 & ~w23119;
assign w23121 = (~w23118 & ~w22994) | (~w23118 & w32419) | (~w22994 & w32419);
assign w23122 = ~w23117 & w23121;
assign w23123 = ~w23120 & ~w23122;
assign w23124 = (~w22969 & w22972) | (~w22969 & w32420) | (w22972 & w32420);
assign w23125 = w23123 & w23124;
assign w23126 = ~w23123 & ~w23124;
assign w23127 = ~w23125 & ~w23126;
assign w23128 = (~w13761 & w37760) | (~w13761 & w37761) | (w37760 & w37761);
assign w23129 = (w13761 & w37762) | (w13761 & w37763) | (w37762 & w37763);
assign w23130 = ~w23128 & ~w23129;
assign w23131 = (~w22992 & ~w22994) | (~w22992 & w32421) | (~w22994 & w32421);
assign w23132 = (~w23105 & ~w23106) | (~w23105 & w32422) | (~w23106 & w32422);
assign w23133 = w5459 & w32423;
assign w23134 = (~w23133 & ~w12670) | (~w23133 & w32424) | (~w12670 & w32424);
assign w23135 = a_41 & ~w23134;
assign w23136 = w23134 & a_41;
assign w23137 = ~w23134 & ~w23135;
assign w23138 = ~w23136 & ~w23137;
assign w23139 = ~w23132 & ~w23138;
assign w23140 = ~w23132 & ~w23139;
assign w23141 = w23132 & ~w23138;
assign w23142 = b_59 & w6761;
assign w23143 = w7075 & w32425;
assign w23144 = b_58 & w6756;
assign w23145 = ~w23143 & ~w23144;
assign w23146 = ~w23142 & w23145;
assign w23147 = (w23146 & ~w11169) | (w23146 & w32426) | (~w11169 & w32426);
assign w23148 = a_47 & ~w23147;
assign w23149 = w23147 & a_47;
assign w23150 = ~w23147 & ~w23148;
assign w23151 = ~w23149 & ~w23150;
assign w23152 = b_56 & w7613;
assign w23153 = w7941 & w32427;
assign w23154 = b_55 & w7608;
assign w23155 = ~w23153 & ~w23154;
assign w23156 = ~w23152 & w23155;
assign w23157 = (w23156 & ~w9798) | (w23156 & w32428) | (~w9798 & w32428);
assign w23158 = a_50 & ~w23157;
assign w23159 = w23157 & a_50;
assign w23160 = ~w23157 & ~w23158;
assign w23161 = ~w23159 & ~w23160;
assign w23162 = (~w23051 & ~w23052) | (~w23051 & w32429) | (~w23052 & w32429);
assign w23163 = b_53 & w8526;
assign w23164 = w8886 & w32430;
assign w23165 = b_52 & w8521;
assign w23166 = ~w23164 & ~w23165;
assign w23167 = ~w23163 & w23166;
assign w23168 = (w23167 & ~w9110) | (w23167 & w32431) | (~w9110 & w32431);
assign w23169 = a_53 & ~w23168;
assign w23170 = w23168 & a_53;
assign w23171 = ~w23168 & ~w23169;
assign w23172 = ~w23170 & ~w23171;
assign w23173 = (~w23033 & ~w23034) | (~w23033 & w32432) | (~w23034 & w32432);
assign w23174 = (~w23015 & ~w23017) | (~w23015 & w32433) | (~w23017 & w32433);
assign w23175 = ~w23001 & ~w23012;
assign w23176 = w12380 & w32434;
assign w23177 = b_41 & ~w12380;
assign w23178 = ~w23176 & ~w23177;
assign w23179 = w22998 & ~w23178;
assign w23180 = w22998 & ~w23179;
assign w23181 = ~w23178 & ~w23179;
assign w23182 = ~w23180 & ~w23181;
assign w23183 = (~w23182 & w23012) | (~w23182 & w32435) | (w23012 & w32435);
assign w23184 = ~w23175 & ~w23183;
assign w23185 = ~w23012 & w32436;
assign w23186 = b_44 & w11620;
assign w23187 = w11969 & w32437;
assign w23188 = b_43 & w11615;
assign w23189 = ~w23187 & ~w23188;
assign w23190 = ~w23186 & w23189;
assign w23191 = (w23190 & ~w6408) | (w23190 & w32438) | (~w6408 & w32438);
assign w23192 = a_62 & ~w23191;
assign w23193 = w23191 & a_62;
assign w23194 = ~w23191 & ~w23192;
assign w23195 = ~w23193 & ~w23194;
assign w23196 = (w23195 & w23184) | (w23195 & w32439) | (w23184 & w32439);
assign w23197 = ~w23184 & w32440;
assign w23198 = ~w23196 & ~w23197;
assign w23199 = b_47 & w10562;
assign w23200 = w10902 & w32441;
assign w23201 = b_46 & w10557;
assign w23202 = ~w23200 & ~w23201;
assign w23203 = ~w23199 & w23202;
assign w23204 = (w23203 & ~w6998) | (w23203 & w26722) | (~w6998 & w26722);
assign w23205 = (w6998 & w27684) | (w6998 & w27685) | (w27684 & w27685);
assign w23206 = (~w6998 & w32442) | (~w6998 & w32443) | (w32442 & w32443);
assign w23207 = ~w23204 & ~w23205;
assign w23208 = ~w23206 & ~w23207;
assign w23209 = ~w23198 & ~w23208;
assign w23210 = w23198 & w23208;
assign w23211 = ~w23209 & ~w23210;
assign w23212 = w23174 & ~w23211;
assign w23213 = ~w23174 & w23211;
assign w23214 = ~w23212 & ~w23213;
assign w23215 = b_50 & w9534;
assign w23216 = w9876 & w32444;
assign w23217 = b_49 & w9529;
assign w23218 = ~w23216 & ~w23217;
assign w23219 = ~w23215 & w23218;
assign w23220 = (w23219 & ~w8162) | (w23219 & w32445) | (~w8162 & w32445);
assign w23221 = a_56 & ~w23220;
assign w23222 = w23220 & a_56;
assign w23223 = ~w23220 & ~w23221;
assign w23224 = ~w23222 & ~w23223;
assign w23225 = ~w23214 & w23224;
assign w23226 = w23214 & ~w23224;
assign w23227 = ~w23225 & ~w23226;
assign w23228 = ~w23173 & w23227;
assign w23229 = ~w23173 & ~w23228;
assign w23230 = w23173 & w23227;
assign w23231 = (~w23172 & w23229) | (~w23172 & w32446) | (w23229 & w32446);
assign w23232 = w23172 & ~w23230;
assign w23233 = ~w23229 & w23232;
assign w23234 = ~w23231 & ~w23233;
assign w23235 = ~w23162 & w23234;
assign w23236 = ~w23162 & ~w23235;
assign w23237 = w23162 & w23234;
assign w23238 = (~w23161 & w23236) | (~w23161 & w32447) | (w23236 & w32447);
assign w23239 = w23161 & ~w23237;
assign w23240 = ~w23236 & w23239;
assign w23241 = ~w23238 & ~w23240;
assign w23242 = (w23241 & w23082) | (w23241 & w32448) | (w23082 & w32448);
assign w23243 = ~w23082 & w32449;
assign w23244 = ~w23242 & ~w23243;
assign w23245 = ~w23151 & w23244;
assign w23246 = w23244 & ~w23245;
assign w23247 = ~w23244 & ~w23151;
assign w23248 = ~w23246 & ~w23247;
assign w23249 = (~w23088 & ~w23089) | (~w23088 & w32450) | (~w23089 & w32450);
assign w23250 = w23248 & w23249;
assign w23251 = ~w23248 & ~w23249;
assign w23252 = ~w23250 & ~w23251;
assign w23253 = b_62 & w5962;
assign w23254 = w6246 & w32451;
assign w23255 = b_61 & w5957;
assign w23256 = ~w23254 & ~w23255;
assign w23257 = ~w23253 & w23256;
assign w23258 = (w23257 & ~w12273) | (w23257 & w32452) | (~w12273 & w32452);
assign w23259 = a_44 & ~w23258;
assign w23260 = w23258 & a_44;
assign w23261 = ~w23258 & ~w23259;
assign w23262 = ~w23260 & ~w23261;
assign w23263 = w23252 & ~w23262;
assign w23264 = w23252 & ~w23263;
assign w23265 = ~w23252 & ~w23262;
assign w23266 = ~w23264 & ~w23265;
assign w23267 = (w23266 & w23140) | (w23266 & w32453) | (w23140 & w32453);
assign w23268 = ~w23140 & w32454;
assign w23269 = ~w23267 & ~w23268;
assign w23270 = ~w23131 & ~w23269;
assign w23271 = w23131 & w23269;
assign w23272 = ~w23270 & ~w23271;
assign w23273 = (~w13761 & w37764) | (~w13761 & w37765) | (w37764 & w37765);
assign w23274 = (w13761 & w37766) | (w13761 & w37767) | (w37766 & w37767);
assign w23275 = ~w23273 & ~w23274;
assign w23276 = b_60 & w6761;
assign w23277 = w7075 & w32455;
assign w23278 = b_59 & w6756;
assign w23279 = ~w23277 & ~w23278;
assign w23280 = ~w23276 & w23279;
assign w23281 = (w23280 & ~w11196) | (w23280 & w32456) | (~w11196 & w32456);
assign w23282 = a_47 & ~w23281;
assign w23283 = w23281 & a_47;
assign w23284 = ~w23281 & ~w23282;
assign w23285 = ~w23283 & ~w23284;
assign w23286 = ~w23235 & ~w23238;
assign w23287 = b_57 & w7613;
assign w23288 = w7941 & w32457;
assign w23289 = b_56 & w7608;
assign w23290 = ~w23288 & ~w23289;
assign w23291 = ~w23287 & w23290;
assign w23292 = (w23291 & ~w10452) | (w23291 & w32458) | (~w10452 & w32458);
assign w23293 = a_50 & ~w23292;
assign w23294 = w23292 & a_50;
assign w23295 = ~w23292 & ~w23293;
assign w23296 = ~w23294 & ~w23295;
assign w23297 = ~w23228 & ~w23231;
assign w23298 = (~w23213 & ~w23214) | (~w23213 & w32459) | (~w23214 & w32459);
assign w23299 = b_51 & w9534;
assign w23300 = w9876 & w32460;
assign w23301 = b_50 & w9529;
assign w23302 = ~w23300 & ~w23301;
assign w23303 = ~w23299 & w23302;
assign w23304 = (w23303 & ~w8186) | (w23303 & w27686) | (~w8186 & w27686);
assign w23305 = (w8186 & w32461) | (w8186 & w32462) | (w32461 & w32462);
assign w23306 = (~w8186 & w32463) | (~w8186 & w32464) | (w32463 & w32464);
assign w23307 = ~w23304 & ~w23305;
assign w23308 = ~w23306 & ~w23307;
assign w23309 = a_41 & ~w22998;
assign w23310 = ~a_41 & w22998;
assign w23311 = ~w23309 & ~w23310;
assign w23312 = w12380 & w32465;
assign w23313 = b_42 & ~w12380;
assign w23314 = ~w23312 & ~w23313;
assign w23315 = w23311 & w23314;
assign w23316 = ~w23311 & ~w23314;
assign w23317 = ~w23315 & ~w23316;
assign w23318 = b_45 & w11620;
assign w23319 = w11969 & w32466;
assign w23320 = b_44 & w11615;
assign w23321 = ~w23319 & ~w23320;
assign w23322 = ~w23318 & w23321;
assign w23323 = (w23322 & ~w6682) | (w23322 & w26477) | (~w6682 & w26477);
assign w23324 = (w6682 & w26723) | (w6682 & w26724) | (w26723 & w26724);
assign w23325 = (~w6682 & w27687) | (~w6682 & w27688) | (w27687 & w27688);
assign w23326 = ~w23323 & ~w23324;
assign w23327 = ~w23325 & ~w23326;
assign w23328 = (w23317 & w23326) | (w23317 & w27689) | (w23326 & w27689);
assign w23329 = w23317 & ~w23328;
assign w23330 = ~w23327 & ~w23328;
assign w23331 = ~w23329 & ~w23330;
assign w23332 = (~w23012 & w32467) | (~w23012 & w32468) | (w32467 & w32468);
assign w23333 = w23331 & w23332;
assign w23334 = ~w23331 & ~w23332;
assign w23335 = ~w23333 & ~w23334;
assign w23336 = b_48 & w10562;
assign w23337 = w10902 & w32469;
assign w23338 = b_47 & w10557;
assign w23339 = ~w23337 & ~w23338;
assign w23340 = ~w23336 & w23339;
assign w23341 = (w23340 & ~w7284) | (w23340 & w26478) | (~w7284 & w26478);
assign w23342 = (w7284 & w26725) | (w7284 & w26726) | (w26725 & w26726);
assign w23343 = (~w7284 & w27690) | (~w7284 & w27691) | (w27690 & w27691);
assign w23344 = ~w23341 & ~w23342;
assign w23345 = ~w23343 & ~w23344;
assign w23346 = w23335 & ~w23345;
assign w23347 = w23345 & w23335;
assign w23348 = ~w23335 & ~w23345;
assign w23349 = (~w23195 & w23184) | (~w23195 & w32470) | (w23184 & w32470);
assign w23350 = ~w23209 & ~w23349;
assign w23351 = (~w23350 & w23348) | (~w23350 & w27692) | (w23348 & w27692);
assign w23352 = ~w23348 & w27693;
assign w23353 = ~w23351 & ~w23352;
assign w23354 = ~w23308 & w23353;
assign w23355 = ~w23353 & ~w23308;
assign w23356 = w23353 & ~w23354;
assign w23357 = ~w23355 & ~w23356;
assign w23358 = (~w23298 & w23356) | (~w23298 & w32471) | (w23356 & w32471);
assign w23359 = ~w23298 & ~w23358;
assign w23360 = ~w23357 & ~w23358;
assign w23361 = ~w23359 & ~w23360;
assign w23362 = b_54 & w8526;
assign w23363 = w8886 & w32472;
assign w23364 = b_53 & w8521;
assign w23365 = ~w23363 & ~w23364;
assign w23366 = ~w23362 & w23365;
assign w23367 = (w23366 & ~w9134) | (w23366 & w32473) | (~w9134 & w32473);
assign w23368 = a_53 & ~w23367;
assign w23369 = w23367 & a_53;
assign w23370 = ~w23367 & ~w23368;
assign w23371 = ~w23369 & ~w23370;
assign w23372 = w23361 & w23371;
assign w23373 = ~w23361 & ~w23371;
assign w23374 = ~w23372 & ~w23373;
assign w23375 = ~w23297 & w23374;
assign w23376 = w23297 & ~w23374;
assign w23377 = ~w23375 & ~w23376;
assign w23378 = w23296 & ~w23377;
assign w23379 = ~w23296 & w23377;
assign w23380 = ~w23378 & ~w23379;
assign w23381 = ~w23286 & w23380;
assign w23382 = w23286 & ~w23380;
assign w23383 = ~w23381 & ~w23382;
assign w23384 = ~w23285 & w23383;
assign w23385 = w23383 & ~w23384;
assign w23386 = ~w23383 & ~w23285;
assign w23387 = ~w23385 & ~w23386;
assign w23388 = (~w23242 & ~w23244) | (~w23242 & w32474) | (~w23244 & w32474);
assign w23389 = w23387 & w23388;
assign w23390 = ~w23387 & ~w23388;
assign w23391 = ~w23389 & ~w23390;
assign w23392 = b_63 & w5962;
assign w23393 = w6246 & w32475;
assign w23394 = b_62 & w5957;
assign w23395 = ~w23393 & ~w23394;
assign w23396 = ~w23392 & w23395;
assign w23397 = (w23396 & ~w12646) | (w23396 & w32476) | (~w12646 & w32476);
assign w23398 = a_44 & ~w23397;
assign w23399 = w23397 & a_44;
assign w23400 = ~w23397 & ~w23398;
assign w23401 = ~w23399 & ~w23400;
assign w23402 = w23391 & ~w23401;
assign w23403 = w23391 & ~w23402;
assign w23404 = ~w23391 & ~w23401;
assign w23405 = ~w23403 & ~w23404;
assign w23406 = (~w23251 & ~w23252) | (~w23251 & w32477) | (~w23252 & w32477);
assign w23407 = w23405 & w23406;
assign w23408 = ~w23405 & ~w23406;
assign w23409 = ~w23407 & ~w23408;
assign w23410 = (~w23266 & w23140) | (~w23266 & w32478) | (w23140 & w32478);
assign w23411 = (w23409 & w23410) | (w23409 & w32479) | (w23410 & w32479);
assign w23412 = ~w23410 & w32480;
assign w23413 = ~w23411 & ~w23412;
assign w23414 = (~w13761 & w37768) | (~w13761 & w37769) | (w37768 & w37769);
assign w23415 = (w13761 & w37770) | (w13761 & w37771) | (w37770 & w37771);
assign w23416 = ~w23414 & ~w23415;
assign w23417 = (~w23384 & w23387) | (~w23384 & w32481) | (w23387 & w32481);
assign w23418 = w6246 & w32482;
assign w23419 = b_63 & w5957;
assign w23420 = ~w23418 & ~w23419;
assign w23421 = ~w12671 & w32483;
assign w23422 = (a_44 & w23421) | (a_44 & w32484) | (w23421 & w32484);
assign w23423 = ~w23421 & w32485;
assign w23424 = ~w23422 & ~w23423;
assign w23425 = ~w23417 & ~w23424;
assign w23426 = w23417 & w23424;
assign w23427 = ~w23425 & ~w23426;
assign w23428 = b_61 & w6761;
assign w23429 = w7075 & w32486;
assign w23430 = b_60 & w6756;
assign w23431 = ~w23429 & ~w23430;
assign w23432 = ~w23428 & w23431;
assign w23433 = (w23432 & ~w11901) | (w23432 & w32487) | (~w11901 & w32487);
assign w23434 = a_47 & ~w23433;
assign w23435 = w23433 & a_47;
assign w23436 = ~w23433 & ~w23434;
assign w23437 = ~w23435 & ~w23436;
assign w23438 = ~w23379 & ~w23381;
assign w23439 = (~w23373 & ~w23374) | (~w23373 & w32488) | (~w23374 & w32488);
assign w23440 = w12380 & w32490;
assign w23441 = b_43 & ~w12380;
assign w23442 = ~w23440 & ~w23441;
assign w23443 = ~a_41 & ~w22998;
assign w23444 = (~w23443 & w23311) | (~w23443 & w32491) | (w23311 & w32491);
assign w23445 = w23442 & ~w23444;
assign w23446 = w23444 & w23442;
assign w23447 = ~w23444 & ~w23445;
assign w23448 = ~w23446 & ~w23447;
assign w23449 = b_46 & w11620;
assign w23450 = w11969 & w32492;
assign w23451 = b_45 & w11615;
assign w23452 = ~w23450 & ~w23451;
assign w23453 = ~w23449 & w23452;
assign w23454 = w23452 & w32493;
assign w23455 = (~w23454 & w6974) | (~w23454 & w32494) | (w6974 & w32494);
assign w23456 = a_62 & ~w23455;
assign w23457 = (~w23448 & w23456) | (~w23448 & w32497) | (w23456 & w32497);
assign w23458 = ~w23456 & w32498;
assign w23459 = ~w23457 & ~w23458;
assign w23460 = (~w23331 & w32499) | (~w23331 & w32500) | (w32499 & w32500);
assign w23461 = (w23331 & w32501) | (w23331 & w32502) | (w32501 & w32502);
assign w23462 = ~w23460 & ~w23461;
assign w23463 = b_49 & w10562;
assign w23464 = w10902 & w32503;
assign w23465 = b_48 & w10557;
assign w23466 = ~w23464 & ~w23465;
assign w23467 = ~w23463 & w23466;
assign w23468 = (w23467 & ~w7859) | (w23467 & w27694) | (~w7859 & w27694);
assign w23469 = (w7859 & w32504) | (w7859 & w32505) | (w32504 & w32505);
assign w23470 = (~w7859 & w32506) | (~w7859 & w32507) | (w32506 & w32507);
assign w23471 = ~w23468 & ~w23469;
assign w23472 = ~w23470 & ~w23471;
assign w23473 = w23462 & ~w23472;
assign w23474 = w23462 & ~w23473;
assign w23475 = ~w23462 & ~w23472;
assign w23476 = ~w23474 & ~w23475;
assign w23477 = (~w27692 & w32508) | (~w27692 & w32509) | (w32508 & w32509);
assign w23478 = w23476 & w23477;
assign w23479 = ~w23476 & ~w23477;
assign w23480 = ~w23478 & ~w23479;
assign w23481 = b_52 & w9534;
assign w23482 = w9876 & w32510;
assign w23483 = b_51 & w9529;
assign w23484 = ~w23482 & ~w23483;
assign w23485 = ~w23481 & w23484;
assign w23486 = (w23485 & ~w8793) | (w23485 & w32511) | (~w8793 & w32511);
assign w23487 = a_56 & ~w23486;
assign w23488 = w23486 & a_56;
assign w23489 = ~w23486 & ~w23487;
assign w23490 = ~w23488 & ~w23489;
assign w23491 = w23480 & ~w23490;
assign w23492 = w23480 & ~w23491;
assign w23493 = ~w23480 & ~w23490;
assign w23494 = ~w23492 & ~w23493;
assign w23495 = ~w23354 & ~w23358;
assign w23496 = w23494 & w23495;
assign w23497 = ~w23494 & ~w23495;
assign w23498 = ~w23496 & ~w23497;
assign w23499 = b_55 & w8526;
assign w23500 = w8886 & w32512;
assign w23501 = b_54 & w8521;
assign w23502 = ~w23500 & ~w23501;
assign w23503 = ~w23499 & w23502;
assign w23504 = (w23503 & ~w9776) | (w23503 & w32513) | (~w9776 & w32513);
assign w23505 = a_53 & ~w23504;
assign w23506 = w23504 & a_53;
assign w23507 = ~w23504 & ~w23505;
assign w23508 = ~w23506 & ~w23507;
assign w23509 = w23498 & ~w23508;
assign w23510 = w23498 & ~w23509;
assign w23511 = ~w23498 & ~w23508;
assign w23512 = ~w23510 & ~w23511;
assign w23513 = ~w23439 & w23512;
assign w23514 = w23439 & ~w23512;
assign w23515 = ~w23513 & ~w23514;
assign w23516 = b_58 & w7613;
assign w23517 = w7941 & w32514;
assign w23518 = b_57 & w7608;
assign w23519 = ~w23517 & ~w23518;
assign w23520 = ~w23516 & w23519;
assign w23521 = (w23520 & ~w10476) | (w23520 & w32515) | (~w10476 & w32515);
assign w23522 = a_50 & ~w23521;
assign w23523 = w23521 & a_50;
assign w23524 = ~w23521 & ~w23522;
assign w23525 = ~w23523 & ~w23524;
assign w23526 = w23515 & w23525;
assign w23527 = ~w23515 & ~w23525;
assign w23528 = ~w23526 & ~w23527;
assign w23529 = ~w23438 & w23528;
assign w23530 = ~w23438 & ~w23529;
assign w23531 = w23528 & ~w23529;
assign w23532 = ~w23530 & ~w23531;
assign w23533 = ~w23437 & ~w23532;
assign w23534 = w23532 & ~w23437;
assign w23535 = ~w23532 & ~w23533;
assign w23536 = ~w23534 & ~w23535;
assign w23537 = w23427 & ~w23536;
assign w23538 = w23427 & ~w23537;
assign w23539 = ~w23536 & ~w23537;
assign w23540 = ~w23538 & ~w23539;
assign w23541 = (~w23402 & w23405) | (~w23402 & w32516) | (w23405 & w32516);
assign w23542 = w23540 & w23541;
assign w23543 = ~w23540 & ~w23541;
assign w23544 = ~w23542 & ~w23543;
assign w23545 = (~w13761 & w37772) | (~w13761 & w37773) | (w37772 & w37773);
assign w23546 = (w13761 & w37774) | (w13761 & w37775) | (w37774 & w37775);
assign w23547 = ~w23545 & ~w23546;
assign w23548 = ~w23425 & ~w23537;
assign w23549 = (~w23529 & w23532) | (~w23529 & w32517) | (w23532 & w32517);
assign w23550 = w6246 & w32518;
assign w23551 = (~w23550 & ~w12670) | (~w23550 & w32519) | (~w12670 & w32519);
assign w23552 = a_44 & ~w23551;
assign w23553 = w23551 & a_44;
assign w23554 = ~w23551 & ~w23552;
assign w23555 = ~w23553 & ~w23554;
assign w23556 = (~w23532 & w32520) | (~w23532 & w32521) | (w32520 & w32521);
assign w23557 = ~w23549 & ~w23556;
assign w23558 = ~w23555 & ~w23556;
assign w23559 = ~w23557 & ~w23558;
assign w23560 = b_59 & w7613;
assign w23561 = w7941 & w32522;
assign w23562 = b_58 & w7608;
assign w23563 = ~w23561 & ~w23562;
assign w23564 = ~w23560 & w23563;
assign w23565 = (w23564 & ~w11169) | (w23564 & w32523) | (~w11169 & w32523);
assign w23566 = a_50 & ~w23565;
assign w23567 = w23565 & a_50;
assign w23568 = ~w23565 & ~w23566;
assign w23569 = ~w23567 & ~w23568;
assign w23570 = (~w23497 & ~w23498) | (~w23497 & w32524) | (~w23498 & w32524);
assign w23571 = b_56 & w8526;
assign w23572 = w8886 & w32525;
assign w23573 = b_55 & w8521;
assign w23574 = ~w23572 & ~w23573;
assign w23575 = ~w23571 & w23574;
assign w23576 = (w23575 & ~w9798) | (w23575 & w32526) | (~w9798 & w32526);
assign w23577 = a_53 & ~w23576;
assign w23578 = w23576 & a_53;
assign w23579 = ~w23576 & ~w23577;
assign w23580 = ~w23578 & ~w23579;
assign w23581 = (~w23479 & ~w23480) | (~w23479 & w32527) | (~w23480 & w32527);
assign w23582 = b_53 & w9534;
assign w23583 = w9876 & w32528;
assign w23584 = b_52 & w9529;
assign w23585 = ~w23583 & ~w23584;
assign w23586 = ~w23582 & w23585;
assign w23587 = (w23586 & ~w9110) | (w23586 & w32529) | (~w9110 & w32529);
assign w23588 = a_56 & ~w23587;
assign w23589 = w23587 & a_56;
assign w23590 = ~w23587 & ~w23588;
assign w23591 = ~w23589 & ~w23590;
assign w23592 = (~w23460 & ~w23462) | (~w23460 & w32530) | (~w23462 & w32530);
assign w23593 = b_50 & w10562;
assign w23594 = w10902 & w32531;
assign w23595 = b_49 & w10557;
assign w23596 = ~w23594 & ~w23595;
assign w23597 = ~w23593 & w23596;
assign w23598 = (w23597 & ~w8162) | (w23597 & w27695) | (~w8162 & w27695);
assign w23599 = (w8162 & w32532) | (w8162 & w32533) | (w32532 & w32533);
assign w23600 = (~w8162 & w32534) | (~w8162 & w32535) | (w32534 & w32535);
assign w23601 = ~w23598 & ~w23599;
assign w23602 = ~w23600 & ~w23601;
assign w23603 = ~w23445 & ~w23457;
assign w23604 = w12380 & w32536;
assign w23605 = b_44 & ~w12380;
assign w23606 = ~w23604 & ~w23605;
assign w23607 = w23442 & ~w23606;
assign w23608 = ~w23442 & w23606;
assign w23609 = ~w23607 & ~w23608;
assign w23610 = b_47 & w11620;
assign w23611 = w11969 & w32537;
assign w23612 = b_46 & w11615;
assign w23613 = ~w23611 & ~w23612;
assign w23614 = ~w23610 & w23613;
assign w23615 = w23613 & w32538;
assign w23616 = (~w6998 & w26479) | (~w6998 & w26480) | (w26479 & w26480);
assign w23617 = (w6998 & w26481) | (w6998 & w26482) | (w26481 & w26482);
assign w23618 = ~w23616 & ~w23617;
assign w23619 = w23609 & ~w23618;
assign w23620 = ~w23609 & w23618;
assign w23621 = ~w23619 & ~w23620;
assign w23622 = ~w23603 & w23621;
assign w23623 = ~w23603 & ~w23622;
assign w23624 = w23621 & ~w23622;
assign w23625 = ~w23623 & ~w23624;
assign w23626 = ~w23602 & ~w23625;
assign w23627 = (w23602 & w23622) | (w23602 & w32539) | (w23622 & w32539);
assign w23628 = ~w23623 & w23627;
assign w23629 = ~w23626 & ~w23628;
assign w23630 = ~w23592 & w23629;
assign w23631 = ~w23629 & ~w23592;
assign w23632 = w23629 & ~w23630;
assign w23633 = (~w23591 & w23632) | (~w23591 & w32540) | (w23632 & w32540);
assign w23634 = ~w23632 & w32541;
assign w23635 = ~w23633 & ~w23634;
assign w23636 = ~w23581 & w23635;
assign w23637 = ~w23581 & ~w23636;
assign w23638 = w23635 & ~w23636;
assign w23639 = ~w23637 & ~w23638;
assign w23640 = ~w23580 & ~w23639;
assign w23641 = (w23580 & w23636) | (w23580 & w32542) | (w23636 & w32542);
assign w23642 = ~w23637 & w23641;
assign w23643 = ~w23640 & ~w23642;
assign w23644 = ~w23570 & w23643;
assign w23645 = w23570 & ~w23643;
assign w23646 = ~w23644 & ~w23645;
assign w23647 = ~w23569 & w23646;
assign w23648 = w23646 & ~w23647;
assign w23649 = ~w23646 & ~w23569;
assign w23650 = ~w23648 & ~w23649;
assign w23651 = ~w23439 & ~w23512;
assign w23652 = (~w23651 & w23515) | (~w23651 & w32543) | (w23515 & w32543);
assign w23653 = ~w23650 & ~w23652;
assign w23654 = ~w23650 & ~w23653;
assign w23655 = ~w23652 & ~w23653;
assign w23656 = ~w23654 & ~w23655;
assign w23657 = b_62 & w6761;
assign w23658 = w7075 & w32544;
assign w23659 = b_61 & w6756;
assign w23660 = ~w23658 & ~w23659;
assign w23661 = ~w23657 & w23660;
assign w23662 = (w23661 & ~w12273) | (w23661 & w32545) | (~w12273 & w32545);
assign w23663 = a_47 & ~w23662;
assign w23664 = w23662 & a_47;
assign w23665 = ~w23662 & ~w23663;
assign w23666 = ~w23664 & ~w23665;
assign w23667 = ~w23656 & ~w23666;
assign w23668 = ~w23656 & ~w23667;
assign w23669 = w23656 & ~w23666;
assign w23670 = ~w23668 & ~w23669;
assign w23671 = ~w23559 & w23670;
assign w23672 = w23559 & ~w23670;
assign w23673 = ~w23671 & ~w23672;
assign w23674 = ~w23548 & ~w23673;
assign w23675 = w23548 & w23673;
assign w23676 = ~w23674 & ~w23675;
assign w23677 = (~w13761 & w37776) | (~w13761 & w37777) | (w37776 & w37777);
assign w23678 = (w13761 & w37778) | (w13761 & w37779) | (w37778 & w37779);
assign w23679 = ~w23677 & ~w23678;
assign w23680 = b_63 & w6761;
assign w23681 = w7075 & w32546;
assign w23682 = b_62 & w6756;
assign w23683 = ~w23681 & ~w23682;
assign w23684 = ~w23680 & w23683;
assign w23685 = (w23684 & ~w12646) | (w23684 & w32547) | (~w12646 & w32547);
assign w23686 = a_47 & ~w23685;
assign w23687 = w23685 & a_47;
assign w23688 = ~w23685 & ~w23686;
assign w23689 = ~w23687 & ~w23688;
assign w23690 = (~w23644 & ~w23646) | (~w23644 & w32548) | (~w23646 & w32548);
assign w23691 = b_60 & w7613;
assign w23692 = w7941 & w32549;
assign w23693 = b_59 & w7608;
assign w23694 = ~w23692 & ~w23693;
assign w23695 = ~w23691 & w23694;
assign w23696 = (w23695 & ~w11196) | (w23695 & w32550) | (~w11196 & w32550);
assign w23697 = a_50 & ~w23696;
assign w23698 = w23696 & a_50;
assign w23699 = ~w23696 & ~w23697;
assign w23700 = ~w23698 & ~w23699;
assign w23701 = (~w23636 & w23639) | (~w23636 & w32551) | (w23639 & w32551);
assign w23702 = b_57 & w8526;
assign w23703 = w8886 & w32552;
assign w23704 = b_56 & w8521;
assign w23705 = ~w23703 & ~w23704;
assign w23706 = ~w23702 & w23705;
assign w23707 = (w23706 & ~w10452) | (w23706 & w32553) | (~w10452 & w32553);
assign w23708 = a_53 & ~w23707;
assign w23709 = w23707 & a_53;
assign w23710 = ~w23707 & ~w23708;
assign w23711 = ~w23709 & ~w23710;
assign w23712 = ~w23630 & ~w23633;
assign w23713 = b_54 & w9534;
assign w23714 = w9876 & w32554;
assign w23715 = b_53 & w9529;
assign w23716 = ~w23714 & ~w23715;
assign w23717 = ~w23713 & w23716;
assign w23718 = (w23717 & ~w9134) | (w23717 & w32555) | (~w9134 & w32555);
assign w23719 = a_56 & ~w23718;
assign w23720 = w23718 & a_56;
assign w23721 = ~w23718 & ~w23719;
assign w23722 = ~w23720 & ~w23721;
assign w23723 = (~w23622 & w23625) | (~w23622 & w32556) | (w23625 & w32556);
assign w23724 = (~w23607 & w23618) | (~w23607 & w26727) | (w23618 & w26727);
assign w23725 = w12380 & w32557;
assign w23726 = b_45 & ~w12380;
assign w23727 = ~w23725 & ~w23726;
assign w23728 = ~a_44 & ~w23727;
assign w23729 = a_44 & w23727;
assign w23730 = ~w23728 & ~w23729;
assign w23731 = ~w23442 & w23730;
assign w23732 = ~w23730 & ~w23442;
assign w23733 = w23730 & ~w23731;
assign w23734 = ~w23732 & ~w23733;
assign w23735 = (~w23618 & w27696) | (~w23618 & w27697) | (w27696 & w27697);
assign w23736 = ~w23724 & ~w23735;
assign w23737 = (w23618 & w32558) | (w23618 & w32559) | (w32558 & w32559);
assign w23738 = ~w23736 & ~w23737;
assign w23739 = b_48 & w11620;
assign w23740 = w11969 & w32560;
assign w23741 = b_47 & w11615;
assign w23742 = ~w23740 & ~w23741;
assign w23743 = ~w23739 & w23742;
assign w23744 = (w23743 & ~w7284) | (w23743 & w27698) | (~w7284 & w27698);
assign w23745 = (w7284 & w32561) | (w7284 & w32562) | (w32561 & w32562);
assign w23746 = (~w7284 & w32563) | (~w7284 & w32564) | (w32563 & w32564);
assign w23747 = ~w23744 & ~w23745;
assign w23748 = ~w23746 & ~w23747;
assign w23749 = (~w23748 & w23736) | (~w23748 & w32565) | (w23736 & w32565);
assign w23750 = ~w23738 & ~w23749;
assign w23751 = ~w23748 & ~w23749;
assign w23752 = ~w23750 & ~w23751;
assign w23753 = b_51 & w10562;
assign w23754 = w10902 & w32566;
assign w23755 = b_50 & w10557;
assign w23756 = ~w23754 & ~w23755;
assign w23757 = ~w23753 & w23756;
assign w23758 = (w23757 & ~w8186) | (w23757 & w27699) | (~w8186 & w27699);
assign w23759 = (w8186 & w32567) | (w8186 & w32568) | (w32567 & w32568);
assign w23760 = (~w8186 & w32569) | (~w8186 & w32570) | (w32569 & w32570);
assign w23761 = ~w23758 & ~w23759;
assign w23762 = ~w23760 & ~w23761;
assign w23763 = w23752 & w23762;
assign w23764 = ~w23752 & ~w23762;
assign w23765 = ~w23763 & ~w23764;
assign w23766 = ~w23723 & w23765;
assign w23767 = w23723 & ~w23765;
assign w23768 = ~w23766 & ~w23767;
assign w23769 = w23722 & ~w23768;
assign w23770 = ~w23722 & w23768;
assign w23771 = ~w23769 & ~w23770;
assign w23772 = ~w23712 & w23771;
assign w23773 = w23712 & ~w23771;
assign w23774 = ~w23772 & ~w23773;
assign w23775 = w23711 & ~w23774;
assign w23776 = ~w23711 & w23774;
assign w23777 = ~w23775 & ~w23776;
assign w23778 = ~w23701 & w23777;
assign w23779 = w23701 & ~w23777;
assign w23780 = ~w23778 & ~w23779;
assign w23781 = w23700 & ~w23780;
assign w23782 = ~w23700 & w23780;
assign w23783 = ~w23781 & ~w23782;
assign w23784 = ~w23690 & w23783;
assign w23785 = w23690 & ~w23783;
assign w23786 = ~w23784 & ~w23785;
assign w23787 = ~w23689 & w23786;
assign w23788 = w23786 & ~w23787;
assign w23789 = ~w23786 & ~w23689;
assign w23790 = ~w23788 & ~w23789;
assign w23791 = (~w23653 & w23656) | (~w23653 & w32571) | (w23656 & w32571);
assign w23792 = w23790 & w23791;
assign w23793 = ~w23790 & ~w23791;
assign w23794 = ~w23792 & ~w23793;
assign w23795 = (~w23556 & w23559) | (~w23556 & w32572) | (w23559 & w32572);
assign w23796 = w23794 & ~w23795;
assign w23797 = ~w23794 & w23795;
assign w23798 = ~w23796 & ~w23797;
assign w23799 = (~w13761 & w37780) | (~w13761 & w37781) | (w37780 & w37781);
assign w23800 = (w13761 & w37782) | (w13761 & w37783) | (w37782 & w37783);
assign w23801 = ~w23799 & ~w23800;
assign w23802 = w7075 & w32573;
assign w23803 = b_63 & w6756;
assign w23804 = ~w23802 & ~w23803;
assign w23805 = ~w12671 & w32574;
assign w23806 = (a_47 & w23805) | (a_47 & w32575) | (w23805 & w32575);
assign w23807 = ~w23805 & w32576;
assign w23808 = ~w23806 & ~w23807;
assign w23809 = (~w23808 & w23784) | (~w23808 & w32577) | (w23784 & w32577);
assign w23810 = ~w23784 & w32578;
assign w23811 = ~w23809 & ~w23810;
assign w23812 = b_61 & w7613;
assign w23813 = w7941 & w32579;
assign w23814 = b_60 & w7608;
assign w23815 = ~w23813 & ~w23814;
assign w23816 = ~w23812 & w23815;
assign w23817 = (w23816 & ~w11901) | (w23816 & w32580) | (~w11901 & w32580);
assign w23818 = a_50 & ~w23817;
assign w23819 = w23817 & a_50;
assign w23820 = ~w23817 & ~w23818;
assign w23821 = ~w23819 & ~w23820;
assign w23822 = ~w23776 & ~w23778;
assign w23823 = ~w23770 & ~w23772;
assign w23824 = b_55 & w9534;
assign w23825 = w9876 & w32581;
assign w23826 = b_54 & w9529;
assign w23827 = ~w23825 & ~w23826;
assign w23828 = ~w23824 & w23827;
assign w23829 = (w23828 & ~w9776) | (w23828 & w32582) | (~w9776 & w32582);
assign w23830 = a_56 & ~w23829;
assign w23831 = w23829 & a_56;
assign w23832 = ~w23829 & ~w23830;
assign w23833 = ~w23831 & ~w23832;
assign w23834 = (~w23764 & ~w23765) | (~w23764 & w32583) | (~w23765 & w32583);
assign w23835 = b_52 & w10562;
assign w23836 = w10902 & w32584;
assign w23837 = b_51 & w10557;
assign w23838 = ~w23836 & ~w23837;
assign w23839 = ~w23835 & w23838;
assign w23840 = (w23839 & ~w8793) | (w23839 & w26483) | (~w8793 & w26483);
assign w23841 = (w8793 & w32585) | (w8793 & w32586) | (w32585 & w32586);
assign w23842 = (~w8793 & w32587) | (~w8793 & w32588) | (w32587 & w32588);
assign w23843 = ~w23840 & ~w23841;
assign w23844 = ~w23842 & ~w23843;
assign w23845 = ~w23735 & ~w23749;
assign w23846 = w12380 & w32589;
assign w23847 = b_46 & ~w12380;
assign w23848 = ~w23846 & ~w23847;
assign w23849 = (~w23728 & ~w23730) | (~w23728 & w32590) | (~w23730 & w32590);
assign w23850 = ~w23848 & w23849;
assign w23851 = w23848 & ~w23849;
assign w23852 = ~w23850 & ~w23851;
assign w23853 = b_49 & w11620;
assign w23854 = w11969 & w32591;
assign w23855 = b_48 & w11615;
assign w23856 = ~w23854 & ~w23855;
assign w23857 = ~w23853 & w23856;
assign w23858 = (w23857 & ~w7859) | (w23857 & w25469) | (~w7859 & w25469);
assign w23859 = (w7859 & w25708) | (w7859 & w25709) | (w25708 & w25709);
assign w23860 = ~w23858 & ~w23859;
assign w23861 = ~w23860 & w32592;
assign w23862 = (w23852 & w23860) | (w23852 & w25470) | (w23860 & w25470);
assign w23863 = ~w23861 & ~w23862;
assign w23864 = (w23863 & w23749) | (w23863 & w32593) | (w23749 & w32593);
assign w23865 = ~w23845 & ~w23864;
assign w23866 = w23863 & ~w23864;
assign w23867 = ~w23865 & ~w23866;
assign w23868 = ~w23844 & ~w23867;
assign w23869 = (w23844 & w23864) | (w23844 & w32594) | (w23864 & w32594);
assign w23870 = ~w23865 & w23869;
assign w23871 = ~w23868 & ~w23870;
assign w23872 = ~w23834 & w23871;
assign w23873 = w23834 & ~w23871;
assign w23874 = ~w23872 & ~w23873;
assign w23875 = ~w23833 & w23874;
assign w23876 = w23874 & ~w23875;
assign w23877 = ~w23874 & ~w23833;
assign w23878 = ~w23876 & ~w23877;
assign w23879 = ~w23823 & w23878;
assign w23880 = w23823 & ~w23878;
assign w23881 = ~w23879 & ~w23880;
assign w23882 = b_58 & w8526;
assign w23883 = w8886 & w32595;
assign w23884 = b_57 & w8521;
assign w23885 = ~w23883 & ~w23884;
assign w23886 = ~w23882 & w23885;
assign w23887 = (w23886 & ~w10476) | (w23886 & w32596) | (~w10476 & w32596);
assign w23888 = a_53 & ~w23887;
assign w23889 = w23887 & a_53;
assign w23890 = ~w23887 & ~w23888;
assign w23891 = ~w23889 & ~w23890;
assign w23892 = w23881 & w23891;
assign w23893 = ~w23881 & ~w23891;
assign w23894 = ~w23892 & ~w23893;
assign w23895 = ~w23822 & w23894;
assign w23896 = ~w23822 & ~w23895;
assign w23897 = w23894 & ~w23895;
assign w23898 = ~w23896 & ~w23897;
assign w23899 = ~w23821 & ~w23898;
assign w23900 = w23898 & ~w23821;
assign w23901 = ~w23898 & ~w23899;
assign w23902 = ~w23900 & ~w23901;
assign w23903 = w23811 & ~w23902;
assign w23904 = w23902 & w23811;
assign w23905 = ~w23902 & ~w23903;
assign w23906 = ~w23904 & ~w23905;
assign w23907 = (~w23787 & w23791) | (~w23787 & w32597) | (w23791 & w32597);
assign w23908 = w23906 & w23907;
assign w23909 = ~w23906 & ~w23907;
assign w23910 = ~w23908 & ~w23909;
assign w23911 = (~w13761 & w37656) | (~w13761 & w37657) | (w37656 & w37657);
assign w23912 = (w13761 & w37784) | (w13761 & w37785) | (w37784 & w37785);
assign w23913 = ~w23911 & ~w23912;
assign w23914 = b_59 & w8526;
assign w23915 = w8886 & w32600;
assign w23916 = b_58 & w8521;
assign w23917 = ~w23915 & ~w23916;
assign w23918 = ~w23914 & w23917;
assign w23919 = (w23918 & ~w11169) | (w23918 & w32601) | (~w11169 & w32601);
assign w23920 = a_53 & ~w23919;
assign w23921 = w23919 & a_53;
assign w23922 = ~w23919 & ~w23920;
assign w23923 = ~w23921 & ~w23922;
assign w23924 = (~w23872 & ~w23874) | (~w23872 & w32602) | (~w23874 & w32602);
assign w23925 = b_56 & w9534;
assign w23926 = w9876 & w32603;
assign w23927 = b_55 & w9529;
assign w23928 = ~w23926 & ~w23927;
assign w23929 = ~w23925 & w23928;
assign w23930 = (w23929 & ~w9798) | (w23929 & w26486) | (~w9798 & w26486);
assign w23931 = (w9798 & w32604) | (w9798 & w32605) | (w32604 & w32605);
assign w23932 = (~w9798 & w32606) | (~w9798 & w32607) | (w32606 & w32607);
assign w23933 = ~w23930 & ~w23931;
assign w23934 = ~w23932 & ~w23933;
assign w23935 = (~w23864 & w23867) | (~w23864 & w32608) | (w23867 & w32608);
assign w23936 = b_53 & w10562;
assign w23937 = w10902 & w32609;
assign w23938 = b_52 & w10557;
assign w23939 = ~w23937 & ~w23938;
assign w23940 = ~w23936 & w23939;
assign w23941 = (w23940 & ~w9110) | (w23940 & w32610) | (~w9110 & w32610);
assign w23942 = a_59 & ~w23941;
assign w23943 = w23941 & a_59;
assign w23944 = ~w23941 & ~w23942;
assign w23945 = ~w23943 & ~w23944;
assign w23946 = ~w23851 & ~w23862;
assign w23947 = w12380 & w32611;
assign w23948 = b_47 & ~w12380;
assign w23949 = ~w23947 & ~w23948;
assign w23950 = w23848 & ~w23949;
assign w23951 = ~w23848 & w23949;
assign w23952 = (w23862 & w26487) | (w23862 & w26488) | (w26487 & w26488);
assign w23953 = ~w23946 & ~w23952;
assign w23954 = (~w23862 & w27700) | (~w23862 & w27701) | (w27700 & w27701);
assign w23955 = ~w23862 & w32612;
assign w23956 = b_50 & w11620;
assign w23957 = w11969 & w32613;
assign w23958 = b_49 & w11615;
assign w23959 = ~w23957 & ~w23958;
assign w23960 = ~w23956 & w23959;
assign w23961 = (w23960 & ~w8162) | (w23960 & w32614) | (~w8162 & w32614);
assign w23962 = a_62 & ~w23961;
assign w23963 = w23961 & a_62;
assign w23964 = ~w23961 & ~w23962;
assign w23965 = ~w23963 & ~w23964;
assign w23966 = (w23965 & w23953) | (w23965 & w32615) | (w23953 & w32615);
assign w23967 = ~w23953 & w32616;
assign w23968 = ~w23966 & ~w23967;
assign w23969 = ~w23945 & ~w23968;
assign w23970 = w23945 & w23968;
assign w23971 = ~w23969 & ~w23970;
assign w23972 = ~w23935 & w23971;
assign w23973 = ~w23935 & ~w23972;
assign w23974 = w23971 & ~w23972;
assign w23975 = ~w23973 & ~w23974;
assign w23976 = ~w23934 & ~w23975;
assign w23977 = (w23934 & w23972) | (w23934 & w32617) | (w23972 & w32617);
assign w23978 = ~w23973 & w23977;
assign w23979 = ~w23976 & ~w23978;
assign w23980 = ~w23924 & w23979;
assign w23981 = w23924 & ~w23979;
assign w23982 = ~w23980 & ~w23981;
assign w23983 = ~w23923 & w23982;
assign w23984 = w23982 & ~w23983;
assign w23985 = ~w23982 & ~w23923;
assign w23986 = ~w23984 & ~w23985;
assign w23987 = ~w23823 & ~w23878;
assign w23988 = (~w23987 & w23881) | (~w23987 & w32618) | (w23881 & w32618);
assign w23989 = ~w23986 & ~w23988;
assign w23990 = ~w23986 & ~w23989;
assign w23991 = w23986 & ~w23988;
assign w23992 = ~w23990 & ~w23991;
assign w23993 = b_62 & w7613;
assign w23994 = w7941 & w32619;
assign w23995 = b_61 & w7608;
assign w23996 = ~w23994 & ~w23995;
assign w23997 = ~w23993 & w23996;
assign w23998 = (w23997 & ~w12273) | (w23997 & w32620) | (~w12273 & w32620);
assign w23999 = a_50 & ~w23998;
assign w24000 = w23998 & a_50;
assign w24001 = ~w23998 & ~w23999;
assign w24002 = ~w24000 & ~w24001;
assign w24003 = (~w24002 & w23990) | (~w24002 & w32621) | (w23990 & w32621);
assign w24004 = ~w23992 & ~w24003;
assign w24005 = ~w24002 & ~w24003;
assign w24006 = ~w24004 & ~w24005;
assign w24007 = w7075 & w32622;
assign w24008 = (w9770 & w32623) | (w9770 & w32624) | (w32623 & w32624);
assign w24009 = (a_47 & w24008) | (a_47 & w32625) | (w24008 & w32625);
assign w24010 = ~w24008 & w32626;
assign w24011 = ~w24009 & ~w24010;
assign w24012 = (~w23898 & w32627) | (~w23898 & w32628) | (w32627 & w32628);
assign w24013 = (w23898 & w32629) | (w23898 & w32630) | (w32629 & w32630);
assign w24014 = ~w24012 & ~w24013;
assign w24015 = ~w24006 & w24014;
assign w24016 = ~w24006 & ~w24015;
assign w24017 = w24014 & ~w24015;
assign w24018 = ~w24016 & ~w24017;
assign w24019 = (~w23809 & w23902) | (~w23809 & w32631) | (w23902 & w32631);
assign w24020 = w24018 & w24019;
assign w24021 = ~w24018 & ~w24019;
assign w24022 = ~w24020 & ~w24021;
assign w24023 = (~w13761 & w37786) | (~w13761 & w37787) | (w37786 & w37787);
assign w24024 = (w13761 & w37788) | (w13761 & w37789) | (w37788 & w37789);
assign w24025 = ~w24023 & ~w24024;
assign w24026 = b_63 & w7613;
assign w24027 = w7941 & w32632;
assign w24028 = b_62 & w7608;
assign w24029 = ~w24027 & ~w24028;
assign w24030 = ~w24026 & w24029;
assign w24031 = (w24030 & ~w12646) | (w24030 & w32633) | (~w12646 & w32633);
assign w24032 = a_50 & ~w24031;
assign w24033 = w24031 & a_50;
assign w24034 = ~w24031 & ~w24032;
assign w24035 = ~w24033 & ~w24034;
assign w24036 = (~w23980 & ~w23982) | (~w23980 & w32634) | (~w23982 & w32634);
assign w24037 = b_60 & w8526;
assign w24038 = w8886 & w32635;
assign w24039 = b_59 & w8521;
assign w24040 = ~w24038 & ~w24039;
assign w24041 = ~w24037 & w24040;
assign w24042 = (w24041 & ~w11196) | (w24041 & w32636) | (~w11196 & w32636);
assign w24043 = a_53 & ~w24042;
assign w24044 = w24042 & a_53;
assign w24045 = ~w24042 & ~w24043;
assign w24046 = ~w24044 & ~w24045;
assign w24047 = (~w23972 & w23975) | (~w23972 & w32637) | (w23975 & w32637);
assign w24048 = b_57 & w9534;
assign w24049 = w9876 & w32638;
assign w24050 = b_56 & w9529;
assign w24051 = ~w24049 & ~w24050;
assign w24052 = ~w24048 & w24051;
assign w24053 = (w24052 & ~w10452) | (w24052 & w32639) | (~w10452 & w32639);
assign w24054 = a_56 & ~w24053;
assign w24055 = w24053 & a_56;
assign w24056 = ~w24053 & ~w24054;
assign w24057 = ~w24055 & ~w24056;
assign w24058 = (~w23965 & w23953) | (~w23965 & w32640) | (w23953 & w32640);
assign w24059 = ~w23969 & ~w24058;
assign w24060 = b_51 & w11620;
assign w24061 = w11969 & w32641;
assign w24062 = b_50 & w11615;
assign w24063 = ~w24061 & ~w24062;
assign w24064 = ~w24060 & w24063;
assign w24065 = (w24064 & ~w8186) | (w24064 & w26489) | (~w8186 & w26489);
assign w24066 = (w8186 & w27702) | (w8186 & w27703) | (w27702 & w27703);
assign w24067 = (~w8186 & w32642) | (~w8186 & w32643) | (w32642 & w32643);
assign w24068 = ~w24065 & ~w24066;
assign w24069 = ~w24067 & ~w24068;
assign w24070 = w12380 & w32644;
assign w24071 = b_48 & ~w12380;
assign w24072 = ~w24070 & ~w24071;
assign w24073 = a_47 & ~w23949;
assign w24074 = ~a_47 & w23949;
assign w24075 = ~w24073 & ~w24074;
assign w24076 = ~w24072 & ~w24075;
assign w24077 = w24072 & w24075;
assign w24078 = ~w24076 & ~w24077;
assign w24079 = (w24078 & w24068) | (w24078 & w32645) | (w24068 & w32645);
assign w24080 = ~w24069 & ~w24079;
assign w24081 = w24078 & ~w24079;
assign w24082 = ~w24080 & ~w24081;
assign w24083 = ~w23954 & ~w24082;
assign w24084 = w24082 & ~w23954;
assign w24085 = ~w24082 & ~w24083;
assign w24086 = b_54 & w10562;
assign w24087 = w10902 & w32646;
assign w24088 = b_53 & w10557;
assign w24089 = ~w24087 & ~w24088;
assign w24090 = ~w24086 & w24089;
assign w24091 = (w24090 & ~w9134) | (w24090 & w32647) | (~w9134 & w32647);
assign w24092 = a_59 & ~w24091;
assign w24093 = w24091 & a_59;
assign w24094 = ~w24091 & ~w24092;
assign w24095 = ~w24093 & ~w24094;
assign w24096 = ~w24085 & w32648;
assign w24097 = (~w24095 & w24085) | (~w24095 & w32649) | (w24085 & w32649);
assign w24098 = ~w24096 & ~w24097;
assign w24099 = ~w24059 & w24098;
assign w24100 = w24059 & ~w24098;
assign w24101 = ~w24099 & ~w24100;
assign w24102 = w24057 & ~w24101;
assign w24103 = ~w24057 & w24101;
assign w24104 = ~w24102 & ~w24103;
assign w24105 = ~w24047 & w24104;
assign w24106 = w24047 & ~w24104;
assign w24107 = ~w24105 & ~w24106;
assign w24108 = w24046 & ~w24107;
assign w24109 = ~w24046 & w24107;
assign w24110 = ~w24108 & ~w24109;
assign w24111 = ~w24036 & w24110;
assign w24112 = w24036 & ~w24110;
assign w24113 = ~w24111 & ~w24112;
assign w24114 = ~w24035 & w24113;
assign w24115 = w24113 & ~w24114;
assign w24116 = ~w24113 & ~w24035;
assign w24117 = ~w24115 & ~w24116;
assign w24118 = ~w23989 & ~w24003;
assign w24119 = w24117 & w24118;
assign w24120 = ~w24117 & ~w24118;
assign w24121 = ~w24119 & ~w24120;
assign w24122 = ~w24012 & ~w24015;
assign w24123 = ~w24121 & w24122;
assign w24124 = w24121 & ~w24122;
assign w24125 = ~w24123 & ~w24124;
assign w24126 = (~w13761 & w37790) | (~w13761 & w37791) | (w37790 & w37791);
assign w24127 = (w13761 & w37792) | (w13761 & w37793) | (w37792 & w37793);
assign w24128 = ~w24126 & ~w24127;
assign w24129 = w7941 & w32650;
assign w24130 = b_63 & w7608;
assign w24131 = ~w24129 & ~w24130;
assign w24132 = (w7616 & w12671) | (w7616 & w32651) | (w12671 & w32651);
assign w24133 = w24131 & ~w24132;
assign w24134 = (a_50 & w24132) | (a_50 & w32652) | (w24132 & w32652);
assign w24135 = ~w24132 & w32653;
assign w24136 = ~w24133 & ~w24134;
assign w24137 = ~w24135 & ~w24136;
assign w24138 = ~w24109 & ~w24111;
assign w24139 = b_61 & w8526;
assign w24140 = w8886 & w32654;
assign w24141 = b_60 & w8521;
assign w24142 = ~w24140 & ~w24141;
assign w24143 = ~w24139 & w24142;
assign w24144 = (w24143 & ~w11901) | (w24143 & w32655) | (~w11901 & w32655);
assign w24145 = a_53 & ~w24144;
assign w24146 = w24144 & a_53;
assign w24147 = ~w24144 & ~w24145;
assign w24148 = ~w24146 & ~w24147;
assign w24149 = ~w24103 & ~w24105;
assign w24150 = b_58 & w9534;
assign w24151 = w9876 & w32656;
assign w24152 = b_57 & w9529;
assign w24153 = ~w24151 & ~w24152;
assign w24154 = ~w24150 & w24153;
assign w24155 = (w24154 & ~w10476) | (w24154 & w32657) | (~w10476 & w32657);
assign w24156 = a_56 & ~w24155;
assign w24157 = w24155 & a_56;
assign w24158 = ~w24155 & ~w24156;
assign w24159 = ~w24157 & ~w24158;
assign w24160 = ~w24097 & ~w24099;
assign w24161 = b_55 & w10562;
assign w24162 = w10902 & w32658;
assign w24163 = b_54 & w10557;
assign w24164 = ~w24162 & ~w24163;
assign w24165 = ~w24161 & w24164;
assign w24166 = (w24165 & ~w9776) | (w24165 & w32659) | (~w9776 & w32659);
assign w24167 = a_59 & ~w24166;
assign w24168 = w24166 & a_59;
assign w24169 = ~w24166 & ~w24167;
assign w24170 = ~w24168 & ~w24169;
assign w24171 = (~w24079 & w24082) | (~w24079 & w32660) | (w24082 & w32660);
assign w24172 = w12380 & w32661;
assign w24173 = b_49 & ~w12380;
assign w24174 = ~w24172 & ~w24173;
assign w24175 = ~a_47 & ~w23949;
assign w24176 = (~w24175 & w24075) | (~w24175 & w32662) | (w24075 & w32662);
assign w24177 = w24174 & ~w24176;
assign w24178 = ~w24174 & w24176;
assign w24179 = ~w24177 & ~w24178;
assign w24180 = b_52 & w11620;
assign w24181 = w11969 & w32663;
assign w24182 = b_51 & w11615;
assign w24183 = ~w24181 & ~w24182;
assign w24184 = ~w24180 & w24183;
assign w24185 = w24183 & w32664;
assign w24186 = (~w24185 & w8793) | (~w24185 & w32665) | (w8793 & w32665);
assign w24187 = a_62 & ~w24186;
assign w24188 = (w24179 & w24187) | (w24179 & w32668) | (w24187 & w32668);
assign w24189 = ~w24187 & w32669;
assign w24190 = ~w24188 & ~w24189;
assign w24191 = ~w24171 & w24190;
assign w24192 = ~w24171 & ~w24191;
assign w24193 = w24171 & w24190;
assign w24194 = (~w24170 & w24192) | (~w24170 & w32670) | (w24192 & w32670);
assign w24195 = w24170 & ~w24193;
assign w24196 = ~w24192 & w24195;
assign w24197 = ~w24194 & ~w24196;
assign w24198 = ~w24160 & w24197;
assign w24199 = w24160 & ~w24197;
assign w24200 = ~w24198 & ~w24199;
assign w24201 = ~w24159 & w24200;
assign w24202 = w24159 & ~w24200;
assign w24203 = ~w24201 & ~w24202;
assign w24204 = ~w24149 & w24203;
assign w24205 = ~w24149 & ~w24204;
assign w24206 = w24203 & ~w24204;
assign w24207 = ~w24205 & ~w24206;
assign w24208 = ~w24148 & ~w24207;
assign w24209 = (w24148 & w24204) | (w24148 & w32671) | (w24204 & w32671);
assign w24210 = ~w24205 & w24209;
assign w24211 = ~w24208 & ~w24210;
assign w24212 = ~w24138 & w24211;
assign w24213 = w24138 & ~w24211;
assign w24214 = ~w24212 & ~w24213;
assign w24215 = ~w24137 & w24214;
assign w24216 = w24214 & ~w24215;
assign w24217 = ~w24214 & ~w24137;
assign w24218 = ~w24216 & ~w24217;
assign w24219 = (~w24114 & w24118) | (~w24114 & w32672) | (w24118 & w32672);
assign w24220 = w24218 & w24219;
assign w24221 = ~w24218 & ~w24219;
assign w24222 = ~w24220 & ~w24221;
assign w24223 = (~w13761 & w37794) | (~w13761 & w37795) | (w37794 & w37795);
assign w24224 = (w13761 & w37796) | (w13761 & w37797) | (w37796 & w37797);
assign w24225 = ~w24223 & ~w24224;
assign w24226 = b_59 & w9534;
assign w24227 = w9876 & w32673;
assign w24228 = b_58 & w9529;
assign w24229 = ~w24227 & ~w24228;
assign w24230 = ~w24226 & w24229;
assign w24231 = (w24230 & ~w11169) | (w24230 & w32674) | (~w11169 & w32674);
assign w24232 = a_56 & ~w24231;
assign w24233 = w24231 & a_56;
assign w24234 = ~w24231 & ~w24232;
assign w24235 = ~w24233 & ~w24234;
assign w24236 = ~w24191 & ~w24194;
assign w24237 = b_53 & w11620;
assign w24238 = w11969 & w32675;
assign w24239 = b_52 & w11615;
assign w24240 = ~w24238 & ~w24239;
assign w24241 = ~w24237 & w24240;
assign w24242 = (w24241 & ~w9110) | (w24241 & w26072) | (~w9110 & w26072);
assign w24243 = (w9110 & w26490) | (w9110 & w26491) | (w26490 & w26491);
assign w24244 = (~w9110 & w27704) | (~w9110 & w27705) | (w27704 & w27705);
assign w24245 = ~w24242 & ~w24243;
assign w24246 = ~w24244 & ~w24245;
assign w24247 = w12380 & w32676;
assign w24248 = b_50 & ~w12380;
assign w24249 = ~w24247 & ~w24248;
assign w24250 = w24174 & ~w24249;
assign w24251 = w24174 & ~w24250;
assign w24252 = ~w24249 & ~w24250;
assign w24253 = ~w24251 & ~w24252;
assign w24254 = (~w24253 & w24245) | (~w24253 & w27706) | (w24245 & w27706);
assign w24255 = ~w24246 & ~w24254;
assign w24256 = ~w24253 & ~w24254;
assign w24257 = ~w24255 & ~w24256;
assign w24258 = ~w24177 & ~w24188;
assign w24259 = w24257 & w24258;
assign w24260 = ~w24257 & ~w24258;
assign w24261 = ~w24259 & ~w24260;
assign w24262 = b_56 & w10562;
assign w24263 = w10902 & w32677;
assign w24264 = b_55 & w10557;
assign w24265 = ~w24263 & ~w24264;
assign w24266 = ~w24262 & w24265;
assign w24267 = (w24266 & ~w9798) | (w24266 & w32678) | (~w9798 & w32678);
assign w24268 = a_59 & ~w24267;
assign w24269 = w24267 & a_59;
assign w24270 = ~w24267 & ~w24268;
assign w24271 = ~w24269 & ~w24270;
assign w24272 = ~w24261 & w24271;
assign w24273 = w24261 & ~w24271;
assign w24274 = ~w24272 & ~w24273;
assign w24275 = ~w24236 & w24274;
assign w24276 = w24236 & ~w24274;
assign w24277 = ~w24275 & ~w24276;
assign w24278 = ~w24235 & w24277;
assign w24279 = w24277 & ~w24278;
assign w24280 = ~w24277 & ~w24235;
assign w24281 = ~w24279 & ~w24280;
assign w24282 = (~w24198 & ~w24200) | (~w24198 & w32679) | (~w24200 & w32679);
assign w24283 = w24281 & w24282;
assign w24284 = ~w24281 & ~w24282;
assign w24285 = ~w24283 & ~w24284;
assign w24286 = b_62 & w8526;
assign w24287 = w8886 & w32680;
assign w24288 = b_61 & w8521;
assign w24289 = ~w24287 & ~w24288;
assign w24290 = ~w24286 & w24289;
assign w24291 = (w24290 & ~w12273) | (w24290 & w32681) | (~w12273 & w32681);
assign w24292 = a_53 & ~w24291;
assign w24293 = w24291 & a_53;
assign w24294 = ~w24291 & ~w24292;
assign w24295 = ~w24293 & ~w24294;
assign w24296 = w24285 & ~w24295;
assign w24297 = w24285 & ~w24296;
assign w24298 = ~w24285 & ~w24295;
assign w24299 = ~w24297 & ~w24298;
assign w24300 = w7941 & w32682;
assign w24301 = (w9770 & w32683) | (w9770 & w32684) | (w32683 & w32684);
assign w24302 = (a_50 & w24301) | (a_50 & w32685) | (w24301 & w32685);
assign w24303 = ~w24301 & w32686;
assign w24304 = ~w24302 & ~w24303;
assign w24305 = (~w24207 & w32687) | (~w24207 & w32688) | (w32687 & w32688);
assign w24306 = (w24207 & w32689) | (w24207 & w32690) | (w32689 & w32690);
assign w24307 = ~w24305 & ~w24306;
assign w24308 = ~w24299 & w24307;
assign w24309 = ~w24299 & ~w24308;
assign w24310 = w24307 & ~w24308;
assign w24311 = ~w24309 & ~w24310;
assign w24312 = (~w24212 & ~w24214) | (~w24212 & w32691) | (~w24214 & w32691);
assign w24313 = w24311 & w24312;
assign w24314 = ~w24311 & ~w24312;
assign w24315 = ~w24313 & ~w24314;
assign w24316 = (~w13761 & w37798) | (~w13761 & w37799) | (w37798 & w37799);
assign w24317 = (w13761 & w37800) | (w13761 & w37801) | (w37800 & w37801);
assign w24318 = ~w24316 & ~w24317;
assign w24319 = (~w24275 & ~w24277) | (~w24275 & w32692) | (~w24277 & w32692);
assign w24320 = b_60 & w9534;
assign w24321 = w9876 & w32693;
assign w24322 = b_59 & w9529;
assign w24323 = ~w24321 & ~w24322;
assign w24324 = ~w24320 & w24323;
assign w24325 = (w24324 & ~w11196) | (w24324 & w32694) | (~w11196 & w32694);
assign w24326 = a_56 & ~w24325;
assign w24327 = w24325 & a_56;
assign w24328 = ~w24325 & ~w24326;
assign w24329 = ~w24327 & ~w24328;
assign w24330 = (~w24260 & ~w24261) | (~w24260 & w32695) | (~w24261 & w32695);
assign w24331 = b_57 & w10562;
assign w24332 = w10902 & w32696;
assign w24333 = b_56 & w10557;
assign w24334 = ~w24332 & ~w24333;
assign w24335 = ~w24331 & w24334;
assign w24336 = (w24335 & ~w10452) | (w24335 & w27707) | (~w10452 & w27707);
assign w24337 = (w10452 & w32697) | (w10452 & w32698) | (w32697 & w32698);
assign w24338 = (~w10452 & w32699) | (~w10452 & w32700) | (w32699 & w32700);
assign w24339 = ~w24336 & ~w24337;
assign w24340 = ~w24338 & ~w24339;
assign w24341 = b_54 & w11620;
assign w24342 = w11969 & w32701;
assign w24343 = b_53 & w11615;
assign w24344 = ~w24342 & ~w24343;
assign w24345 = ~w24341 & w24344;
assign w24346 = (w24345 & ~w9134) | (w24345 & w27708) | (~w9134 & w27708);
assign w24347 = (w9134 & w32702) | (w9134 & w32703) | (w32702 & w32703);
assign w24348 = (~w9134 & w32704) | (~w9134 & w32705) | (w32704 & w32705);
assign w24349 = ~w24346 & ~w24347;
assign w24350 = ~w24348 & ~w24349;
assign w24351 = ~w24250 & ~w24254;
assign w24352 = w12380 & w32706;
assign w24353 = b_51 & ~w12380;
assign w24354 = ~w24352 & ~w24353;
assign w24355 = ~a_50 & ~w24354;
assign w24356 = a_50 & w24354;
assign w24357 = ~w24355 & ~w24356;
assign w24358 = ~w24174 & w24357;
assign w24359 = w24174 & ~w24357;
assign w24360 = ~w24358 & ~w24359;
assign w24361 = (w24360 & w24254) | (w24360 & w32707) | (w24254 & w32707);
assign w24362 = ~w24351 & ~w24361;
assign w24363 = ~w24254 & w32708;
assign w24364 = (~w24350 & w24362) | (~w24350 & w32709) | (w24362 & w32709);
assign w24365 = w24350 & ~w24363;
assign w24366 = ~w24362 & w24365;
assign w24367 = ~w24364 & ~w24366;
assign w24368 = ~w24340 & w24367;
assign w24369 = ~w24367 & ~w24340;
assign w24370 = w24367 & ~w24368;
assign w24371 = (~w24330 & w24370) | (~w24330 & w32710) | (w24370 & w32710);
assign w24372 = ~w24370 & w32711;
assign w24373 = ~w24371 & ~w24372;
assign w24374 = ~w24329 & w24373;
assign w24375 = w24329 & ~w24373;
assign w24376 = ~w24374 & ~w24375;
assign w24377 = ~w24319 & w24376;
assign w24378 = w24319 & ~w24376;
assign w24379 = ~w24377 & ~w24378;
assign w24380 = b_63 & w8526;
assign w24381 = w8886 & w32712;
assign w24382 = b_62 & w8521;
assign w24383 = ~w24381 & ~w24382;
assign w24384 = ~w24380 & w24383;
assign w24385 = (w24384 & ~w12646) | (w24384 & w32713) | (~w12646 & w32713);
assign w24386 = a_53 & ~w24385;
assign w24387 = w24385 & a_53;
assign w24388 = ~w24385 & ~w24386;
assign w24389 = ~w24387 & ~w24388;
assign w24390 = w24379 & ~w24389;
assign w24391 = w24379 & ~w24390;
assign w24392 = ~w24379 & ~w24389;
assign w24393 = ~w24391 & ~w24392;
assign w24394 = (~w24284 & ~w24285) | (~w24284 & w32714) | (~w24285 & w32714);
assign w24395 = w24393 & w24394;
assign w24396 = ~w24393 & ~w24394;
assign w24397 = ~w24395 & ~w24396;
assign w24398 = ~w24308 & w32715;
assign w24399 = (w24397 & w24308) | (w24397 & w32716) | (w24308 & w32716);
assign w24400 = ~w24398 & ~w24399;
assign w24401 = (~w13761 & w37802) | (~w13761 & w37803) | (w37802 & w37803);
assign w24402 = (w13761 & w37804) | (w13761 & w37805) | (w37804 & w37805);
assign w24403 = ~w24401 & ~w24402;
assign w24404 = w8886 & w32717;
assign w24405 = b_63 & w8521;
assign w24406 = ~w24404 & ~w24405;
assign w24407 = (w8529 & w12671) | (w8529 & w32718) | (w12671 & w32718);
assign w24408 = w24406 & ~w24407;
assign w24409 = (a_53 & w24407) | (a_53 & w32719) | (w24407 & w32719);
assign w24410 = ~w24407 & w32720;
assign w24411 = ~w24408 & ~w24409;
assign w24412 = ~w24410 & ~w24411;
assign w24413 = ~w24374 & ~w24377;
assign w24414 = b_61 & w9534;
assign w24415 = w9876 & w32721;
assign w24416 = b_60 & w9529;
assign w24417 = ~w24415 & ~w24416;
assign w24418 = ~w24414 & w24417;
assign w24419 = (w24418 & ~w11901) | (w24418 & w32722) | (~w11901 & w32722);
assign w24420 = a_56 & ~w24419;
assign w24421 = w24419 & a_56;
assign w24422 = ~w24419 & ~w24420;
assign w24423 = ~w24421 & ~w24422;
assign w24424 = ~w24368 & ~w24371;
assign w24425 = b_58 & w10562;
assign w24426 = w10902 & w32723;
assign w24427 = b_57 & w10557;
assign w24428 = ~w24426 & ~w24427;
assign w24429 = ~w24425 & w24428;
assign w24430 = (w24429 & ~w10476) | (w24429 & w32724) | (~w10476 & w32724);
assign w24431 = a_59 & ~w24430;
assign w24432 = w24430 & a_59;
assign w24433 = ~w24430 & ~w24431;
assign w24434 = ~w24432 & ~w24433;
assign w24435 = w12380 & w32725;
assign w24436 = b_52 & ~w12380;
assign w24437 = ~w24435 & ~w24436;
assign w24438 = (~w24355 & ~w24357) | (~w24355 & w32726) | (~w24357 & w32726);
assign w24439 = ~w24437 & w24438;
assign w24440 = w24437 & ~w24438;
assign w24441 = ~w24439 & ~w24440;
assign w24442 = b_55 & w11620;
assign w24443 = w11969 & w32727;
assign w24444 = b_54 & w11615;
assign w24445 = ~w24443 & ~w24444;
assign w24446 = ~w24442 & w24445;
assign w24447 = (w24446 & ~w9776) | (w24446 & w25471) | (~w9776 & w25471);
assign w24448 = (w9776 & w26073) | (w9776 & w26074) | (w26073 & w26074);
assign w24449 = ~w24447 & ~w24448;
assign w24450 = ~w24449 & w32728;
assign w24451 = (w24441 & w24449) | (w24441 & w26494) | (w24449 & w26494);
assign w24452 = ~w24450 & ~w24451;
assign w24453 = (w24452 & w24364) | (w24452 & w32729) | (w24364 & w32729);
assign w24454 = ~w24364 & w32730;
assign w24455 = ~w24453 & ~w24454;
assign w24456 = ~w24434 & w24455;
assign w24457 = w24434 & ~w24455;
assign w24458 = ~w24456 & ~w24457;
assign w24459 = ~w24424 & w24458;
assign w24460 = ~w24424 & ~w24459;
assign w24461 = w24424 & w24458;
assign w24462 = (~w24423 & w24460) | (~w24423 & w32731) | (w24460 & w32731);
assign w24463 = w24423 & ~w24461;
assign w24464 = ~w24460 & w24463;
assign w24465 = ~w24462 & ~w24464;
assign w24466 = ~w24413 & w24465;
assign w24467 = w24413 & ~w24465;
assign w24468 = ~w24466 & ~w24467;
assign w24469 = ~w24412 & w24468;
assign w24470 = w24468 & ~w24469;
assign w24471 = ~w24468 & ~w24412;
assign w24472 = ~w24470 & ~w24471;
assign w24473 = ~w24390 & ~w24396;
assign w24474 = w24472 & w24473;
assign w24475 = ~w24472 & ~w24473;
assign w24476 = ~w24474 & ~w24475;
assign w24477 = (~w13761 & w37806) | (~w13761 & w37807) | (w37806 & w37807);
assign w24478 = (w13761 & w37808) | (w13761 & w37809) | (w37808 & w37809);
assign w24479 = ~w24477 & ~w24478;
assign w24480 = (~w24453 & ~w24455) | (~w24453 & w32732) | (~w24455 & w32732);
assign w24481 = ~w24440 & ~w24451;
assign w24482 = w12380 & w32733;
assign w24483 = b_53 & ~w12380;
assign w24484 = ~w24482 & ~w24483;
assign w24485 = w24437 & ~w24484;
assign w24486 = ~w24437 & w24484;
assign w24487 = (w24451 & w32734) | (w24451 & w32735) | (w32734 & w32735);
assign w24488 = ~w24481 & ~w24487;
assign w24489 = (~w24451 & w32736) | (~w24451 & w32737) | (w32736 & w32737);
assign w24490 = ~w24451 & w32738;
assign w24491 = b_56 & w11620;
assign w24492 = w11969 & w32739;
assign w24493 = b_55 & w11615;
assign w24494 = ~w24492 & ~w24493;
assign w24495 = ~w24491 & w24494;
assign w24496 = (w24495 & ~w9798) | (w24495 & w32740) | (~w9798 & w32740);
assign w24497 = a_62 & ~w24496;
assign w24498 = w24496 & a_62;
assign w24499 = ~w24496 & ~w24497;
assign w24500 = ~w24498 & ~w24499;
assign w24501 = (w24500 & w24488) | (w24500 & w32741) | (w24488 & w32741);
assign w24502 = ~w24488 & w32742;
assign w24503 = ~w24501 & ~w24502;
assign w24504 = b_59 & w10562;
assign w24505 = w10902 & w32743;
assign w24506 = b_58 & w10557;
assign w24507 = ~w24505 & ~w24506;
assign w24508 = ~w24504 & w24507;
assign w24509 = (w24508 & ~w11169) | (w24508 & w32744) | (~w11169 & w32744);
assign w24510 = a_59 & ~w24509;
assign w24511 = w24509 & a_59;
assign w24512 = ~w24509 & ~w24510;
assign w24513 = ~w24511 & ~w24512;
assign w24514 = ~w24503 & ~w24513;
assign w24515 = w24503 & w24513;
assign w24516 = ~w24514 & ~w24515;
assign w24517 = w24480 & ~w24516;
assign w24518 = ~w24480 & w24516;
assign w24519 = ~w24517 & ~w24518;
assign w24520 = b_62 & w9534;
assign w24521 = w9876 & w32745;
assign w24522 = b_61 & w9529;
assign w24523 = ~w24521 & ~w24522;
assign w24524 = ~w24520 & w24523;
assign w24525 = (w24524 & ~w12273) | (w24524 & w32746) | (~w12273 & w32746);
assign w24526 = a_56 & ~w24525;
assign w24527 = w24525 & a_56;
assign w24528 = ~w24525 & ~w24526;
assign w24529 = ~w24527 & ~w24528;
assign w24530 = w24519 & ~w24529;
assign w24531 = w24519 & ~w24530;
assign w24532 = ~w24519 & ~w24529;
assign w24533 = ~w24531 & ~w24532;
assign w24534 = w8886 & w32747;
assign w24535 = (w9770 & w32748) | (w9770 & w32749) | (w32748 & w32749);
assign w24536 = (a_53 & w24535) | (a_53 & w32750) | (w24535 & w32750);
assign w24537 = ~w24535 & w32751;
assign w24538 = ~w24536 & ~w24537;
assign w24539 = (~w24538 & w24462) | (~w24538 & w32752) | (w24462 & w32752);
assign w24540 = ~w24462 & w32753;
assign w24541 = ~w24539 & ~w24540;
assign w24542 = ~w24533 & w24541;
assign w24543 = ~w24541 & ~w24533;
assign w24544 = w24541 & ~w24542;
assign w24545 = ~w24543 & ~w24544;
assign w24546 = (~w24466 & ~w24468) | (~w24466 & w32754) | (~w24468 & w32754);
assign w24547 = w24545 & w24546;
assign w24548 = ~w24545 & ~w24546;
assign w24549 = ~w24547 & ~w24548;
assign w24550 = (~w13761 & w37810) | (~w13761 & w37811) | (w37810 & w37811);
assign w24551 = (w13761 & w37812) | (w13761 & w37813) | (w37812 & w37813);
assign w24552 = ~w24550 & ~w24551;
assign w24553 = (~w24539 & ~w24541) | (~w24539 & w32755) | (~w24541 & w32755);
assign w24554 = (~w24518 & ~w24519) | (~w24518 & w26963) | (~w24519 & w26963);
assign w24555 = b_63 & w9534;
assign w24556 = w9876 & w32756;
assign w24557 = b_62 & w9529;
assign w24558 = ~w24556 & ~w24557;
assign w24559 = ~w24555 & w24558;
assign w24560 = (w24559 & ~w12646) | (w24559 & w32757) | (~w12646 & w32757);
assign w24561 = a_56 & ~w24560;
assign w24562 = w24560 & a_56;
assign w24563 = ~w24560 & ~w24561;
assign w24564 = ~w24562 & ~w24563;
assign w24565 = ~w24554 & ~w24564;
assign w24566 = ~w24554 & ~w24565;
assign w24567 = w24554 & ~w24564;
assign w24568 = (~w24500 & w24488) | (~w24500 & w32758) | (w24488 & w32758);
assign w24569 = ~w24514 & ~w24568;
assign w24570 = b_60 & w10562;
assign w24571 = w10902 & w32759;
assign w24572 = b_59 & w10557;
assign w24573 = ~w24571 & ~w24572;
assign w24574 = ~w24570 & w24573;
assign w24575 = (w24574 & ~w11196) | (w24574 & w32760) | (~w11196 & w32760);
assign w24576 = a_59 & ~w24575;
assign w24577 = w24575 & a_59;
assign w24578 = ~w24575 & ~w24576;
assign w24579 = ~w24577 & ~w24578;
assign w24580 = a_53 & ~w24484;
assign w24581 = ~a_53 & w24484;
assign w24582 = ~w24580 & ~w24581;
assign w24583 = w12380 & w32761;
assign w24584 = b_54 & ~w12380;
assign w24585 = ~w24583 & ~w24584;
assign w24586 = w24582 & w24585;
assign w24587 = ~w24582 & ~w24585;
assign w24588 = ~w24586 & ~w24587;
assign w24589 = b_57 & w11620;
assign w24590 = w11969 & w32762;
assign w24591 = b_56 & w11615;
assign w24592 = ~w24590 & ~w24591;
assign w24593 = ~w24589 & w24592;
assign w24594 = (w24593 & ~w10452) | (w24593 & w26964) | (~w10452 & w26964);
assign w24595 = (w10452 & w27709) | (w10452 & w27710) | (w27709 & w27710);
assign w24596 = (~w10452 & w32763) | (~w10452 & w32764) | (w32763 & w32764);
assign w24597 = ~w24594 & ~w24595;
assign w24598 = ~w24596 & ~w24597;
assign w24599 = (w24588 & w24597) | (w24588 & w32765) | (w24597 & w32765);
assign w24600 = w24588 & ~w24599;
assign w24601 = ~w24598 & ~w24599;
assign w24602 = ~w24600 & ~w24601;
assign w24603 = ~w24489 & ~w24602;
assign w24604 = w24489 & w24602;
assign w24605 = ~w24603 & ~w24604;
assign w24606 = ~w24579 & w24605;
assign w24607 = ~w24605 & ~w24579;
assign w24608 = w24605 & ~w24606;
assign w24609 = ~w24607 & ~w24608;
assign w24610 = ~w24569 & ~w24609;
assign w24611 = w24609 & ~w24569;
assign w24612 = ~w24609 & ~w24610;
assign w24613 = ~w24611 & ~w24612;
assign w24614 = (w24613 & w24566) | (w24613 & w32766) | (w24566 & w32766);
assign w24615 = ~w24566 & w32767;
assign w24616 = ~w24614 & ~w24615;
assign w24617 = ~w24553 & ~w24616;
assign w24618 = w24553 & w24616;
assign w24619 = ~w24617 & ~w24618;
assign w24620 = (~w13761 & w37814) | (~w13761 & w37815) | (w37814 & w37815);
assign w24621 = (w13761 & w37816) | (w13761 & w37817) | (w37816 & w37817);
assign w24622 = ~w24620 & ~w24621;
assign w24623 = w9876 & w32768;
assign w24624 = b_63 & w9529;
assign w24625 = ~w24623 & ~w24624;
assign w24626 = (w9537 & w12671) | (w9537 & w32769) | (w12671 & w32769);
assign w24627 = w24625 & ~w24626;
assign w24628 = (a_56 & w24626) | (a_56 & w32770) | (w24626 & w32770);
assign w24629 = ~w24626 & w32771;
assign w24630 = ~w24627 & ~w24628;
assign w24631 = ~w24629 & ~w24630;
assign w24632 = (~w24606 & w24609) | (~w24606 & w32772) | (w24609 & w32772);
assign w24633 = b_61 & w10562;
assign w24634 = w10902 & w32773;
assign w24635 = b_60 & w10557;
assign w24636 = ~w24634 & ~w24635;
assign w24637 = ~w24633 & w24636;
assign w24638 = (w24637 & ~w11901) | (w24637 & w32774) | (~w11901 & w32774);
assign w24639 = a_59 & ~w24638;
assign w24640 = w24638 & a_59;
assign w24641 = ~w24638 & ~w24639;
assign w24642 = ~w24640 & ~w24641;
assign w24643 = (~w24599 & w24602) | (~w24599 & w32775) | (w24602 & w32775);
assign w24644 = w12380 & w32776;
assign w24645 = b_55 & ~w12380;
assign w24646 = ~w24644 & ~w24645;
assign w24647 = ~a_53 & ~w24484;
assign w24648 = (~w24647 & w24582) | (~w24647 & w32777) | (w24582 & w32777);
assign w24649 = w24646 & ~w24648;
assign w24650 = ~w24646 & w24648;
assign w24651 = ~w24649 & ~w24650;
assign w24652 = b_58 & w11620;
assign w24653 = w11969 & w32778;
assign w24654 = b_57 & w11615;
assign w24655 = ~w24653 & ~w24654;
assign w24656 = ~w24652 & w24655;
assign w24657 = w24655 & w32779;
assign w24658 = (~w24657 & w10476) | (~w24657 & w32780) | (w10476 & w32780);
assign w24659 = a_62 & ~w24658;
assign w24660 = (w24651 & w24659) | (w24651 & w32783) | (w24659 & w32783);
assign w24661 = ~w24659 & w32784;
assign w24662 = ~w24660 & ~w24661;
assign w24663 = ~w24643 & w24662;
assign w24664 = ~w24643 & ~w24663;
assign w24665 = w24643 & w24662;
assign w24666 = (~w24642 & w24664) | (~w24642 & w32785) | (w24664 & w32785);
assign w24667 = w24642 & ~w24665;
assign w24668 = ~w24664 & w24667;
assign w24669 = ~w24666 & ~w24668;
assign w24670 = ~w24632 & w24669;
assign w24671 = w24632 & ~w24669;
assign w24672 = ~w24670 & ~w24671;
assign w24673 = ~w24631 & w24672;
assign w24674 = w24672 & ~w24673;
assign w24675 = ~w24672 & ~w24631;
assign w24676 = ~w24674 & ~w24675;
assign w24677 = (~w24613 & w24566) | (~w24613 & w32786) | (w24566 & w32786);
assign w24678 = ~w24565 & ~w24677;
assign w24679 = ~w24676 & ~w24678;
assign w24680 = ~w24676 & ~w24679;
assign w24681 = ~w24678 & ~w24679;
assign w24682 = ~w24680 & ~w24681;
assign w24683 = (~w13761 & w37818) | (~w13761 & w37819) | (w37818 & w37819);
assign w24684 = (w13761 & w37820) | (w13761 & w37821) | (w37820 & w37821);
assign w24685 = ~w24683 & ~w24684;
assign w24686 = b_59 & w11620;
assign w24687 = w11969 & w32787;
assign w24688 = b_58 & w11615;
assign w24689 = ~w24687 & ~w24688;
assign w24690 = ~w24686 & w24689;
assign w24691 = (w24690 & ~w26965) | (w24690 & w32788) | (~w26965 & w32788);
assign w24692 = (w26965 & w32789) | (w26965 & w32790) | (w32789 & w32790);
assign w24693 = a_62 & ~w24692;
assign w24694 = ~w24691 & ~w24692;
assign w24695 = ~w24693 & ~w24694;
assign w24696 = w12380 & w32791;
assign w24697 = b_56 & ~w12380;
assign w24698 = ~w24696 & ~w24697;
assign w24699 = w24646 & ~w24698;
assign w24700 = w24646 & ~w24699;
assign w24701 = ~w24698 & ~w24699;
assign w24702 = ~w24700 & ~w24701;
assign w24703 = ~w24695 & ~w24702;
assign w24704 = ~w24695 & ~w24703;
assign w24705 = w24695 & ~w24702;
assign w24706 = ~w24649 & ~w24660;
assign w24707 = ~w24704 & w32792;
assign w24708 = (~w24706 & w24704) | (~w24706 & w32793) | (w24704 & w32793);
assign w24709 = ~w24707 & ~w24708;
assign w24710 = b_62 & w10562;
assign w24711 = w10902 & w32794;
assign w24712 = b_61 & w10557;
assign w24713 = ~w24711 & ~w24712;
assign w24714 = ~w24710 & w24713;
assign w24715 = (w24714 & ~w12273) | (w24714 & w32795) | (~w12273 & w32795);
assign w24716 = a_59 & ~w24715;
assign w24717 = w24715 & a_59;
assign w24718 = ~w24715 & ~w24716;
assign w24719 = ~w24717 & ~w24718;
assign w24720 = w24709 & ~w24719;
assign w24721 = w24709 & ~w24720;
assign w24722 = ~w24709 & ~w24719;
assign w24723 = ~w24721 & ~w24722;
assign w24724 = w9876 & w32796;
assign w24725 = (w9770 & w32797) | (w9770 & w32798) | (w32797 & w32798);
assign w24726 = (a_56 & w24725) | (a_56 & w32799) | (w24725 & w32799);
assign w24727 = ~w24725 & w32800;
assign w24728 = ~w24726 & ~w24727;
assign w24729 = (~w24728 & w24666) | (~w24728 & w32801) | (w24666 & w32801);
assign w24730 = ~w24666 & w32802;
assign w24731 = ~w24729 & ~w24730;
assign w24732 = ~w24723 & w24731;
assign w24733 = ~w24731 & ~w24723;
assign w24734 = w24731 & ~w24732;
assign w24735 = ~w24733 & ~w24734;
assign w24736 = (~w24670 & ~w24672) | (~w24670 & w32803) | (~w24672 & w32803);
assign w24737 = w24735 & w24736;
assign w24738 = ~w24735 & ~w24736;
assign w24739 = ~w24737 & ~w24738;
assign w24740 = (~w13761 & w37822) | (~w13761 & w37823) | (w37822 & w37823);
assign w24741 = (w13761 & w37824) | (w13761 & w37825) | (w37824 & w37825);
assign w24742 = ~w24740 & ~w24741;
assign w24743 = (~w24708 & ~w24709) | (~w24708 & w32804) | (~w24709 & w32804);
assign w24744 = b_63 & w10562;
assign w24745 = w10902 & w32805;
assign w24746 = b_62 & w10557;
assign w24747 = ~w24745 & ~w24746;
assign w24748 = ~w24744 & w24747;
assign w24749 = (w24748 & ~w12646) | (w24748 & w32806) | (~w12646 & w32806);
assign w24750 = a_59 & ~w24749;
assign w24751 = w24749 & a_59;
assign w24752 = ~w24749 & ~w24750;
assign w24753 = ~w24751 & ~w24752;
assign w24754 = ~w24743 & ~w24753;
assign w24755 = ~w24743 & ~w24754;
assign w24756 = w24743 & ~w24753;
assign w24757 = ~w24755 & ~w24756;
assign w24758 = w12380 & w32807;
assign w24759 = b_57 & ~w12380;
assign w24760 = ~w24758 & ~w24759;
assign w24761 = ~a_56 & ~w24760;
assign w24762 = w24760 & ~a_56;
assign w24763 = ~w24760 & ~w24761;
assign w24764 = ~w24762 & ~w24763;
assign w24765 = (~w24646 & w24763) | (~w24646 & w32808) | (w24763 & w32808);
assign w24766 = ~w24646 & ~w24765;
assign w24767 = ~w24764 & ~w24765;
assign w24768 = ~w24766 & ~w24767;
assign w24769 = (w24695 & w32810) | (w24695 & w32811) | (w32810 & w32811);
assign w24770 = (~w24695 & w32812) | (~w24695 & w32813) | (w32812 & w32813);
assign w24771 = ~w24769 & ~w24770;
assign w24772 = b_60 & w11620;
assign w24773 = w11969 & w32814;
assign w24774 = b_59 & w11615;
assign w24775 = ~w24773 & ~w24774;
assign w24776 = ~w24772 & w24775;
assign w24777 = (w24776 & ~w11196) | (w24776 & w32815) | (~w11196 & w32815);
assign w24778 = a_62 & ~w24777;
assign w24779 = w24777 & a_62;
assign w24780 = ~w24777 & ~w24778;
assign w24781 = ~w24779 & ~w24780;
assign w24782 = w24771 & ~w24781;
assign w24783 = ~w24771 & w24781;
assign w24784 = (~w24783 & w24755) | (~w24783 & w32816) | (w24755 & w32816);
assign w24785 = ~w24782 & w24784;
assign w24786 = ~w24757 & ~w24785;
assign w24787 = (~w24784 & w32818) | (~w24784 & w32819) | (w32818 & w32819);
assign w24788 = (~w24729 & ~w24731) | (~w24729 & w32820) | (~w24731 & w32820);
assign w24789 = ~w24786 & w32821;
assign w24790 = (~w24788 & w24786) | (~w24788 & w32822) | (w24786 & w32822);
assign w24791 = ~w24789 & ~w24790;
assign w24792 = (~w13761 & w37826) | (~w13761 & w37827) | (w37826 & w37827);
assign w24793 = (w13761 & w37828) | (w13761 & w37829) | (w37828 & w37829);
assign w24794 = ~w24792 & ~w24793;
assign w24795 = (~w24770 & ~w24771) | (~w24770 & w32823) | (~w24771 & w32823);
assign w24796 = w12380 & w32824;
assign w24797 = b_58 & ~w12380;
assign w24798 = ~w24796 & ~w24797;
assign w24799 = ~w24765 & w32825;
assign w24800 = (w24798 & w24765) | (w24798 & w32826) | (w24765 & w32826);
assign w24801 = ~w24799 & ~w24800;
assign w24802 = b_61 & w11620;
assign w24803 = w11969 & w32827;
assign w24804 = b_60 & w11615;
assign w24805 = ~w24803 & ~w24804;
assign w24806 = ~w24802 & w24805;
assign w24807 = w24805 & w32828;
assign w24808 = (~w24807 & w11901) | (~w24807 & w32829) | (w11901 & w32829);
assign w24809 = a_62 & ~w24808;
assign w24810 = (w24801 & w24809) | (w24801 & w32832) | (w24809 & w32832);
assign w24811 = ~w24809 & w32833;
assign w24812 = ~w24810 & ~w24811;
assign w24813 = ~w24795 & w24812;
assign w24814 = w24795 & ~w24812;
assign w24815 = ~w24813 & ~w24814;
assign w24816 = w10902 & w32834;
assign w24817 = b_63 & w10557;
assign w24818 = ~w24816 & ~w24817;
assign w24819 = (w10565 & w12671) | (w10565 & w32835) | (w12671 & w32835);
assign w24820 = w24818 & ~w24819;
assign w24821 = (a_59 & w24819) | (a_59 & w32836) | (w24819 & w32836);
assign w24822 = ~w24819 & w32837;
assign w24823 = ~w24820 & ~w24821;
assign w24824 = ~w24822 & ~w24823;
assign w24825 = w24815 & ~w24824;
assign w24826 = w24815 & ~w24825;
assign w24827 = ~w24815 & ~w24824;
assign w24828 = ~w24826 & ~w24827;
assign w24829 = (~w24754 & ~w24784) | (~w24754 & w32838) | (~w24784 & w32838);
assign w24830 = w24828 & w24829;
assign w24831 = ~w24828 & ~w24829;
assign w24832 = ~w24830 & ~w24831;
assign w24833 = (~w13761 & w37830) | (~w13761 & w37831) | (w37830 & w37831);
assign w24834 = (w13761 & w37832) | (w13761 & w37833) | (w37832 & w37833);
assign w24835 = ~w24833 & ~w24834;
assign w24836 = (~w24813 & ~w24815) | (~w24813 & w32839) | (~w24815 & w32839);
assign w24837 = ~w24800 & ~w24810;
assign w24838 = w12380 & w32840;
assign w24839 = b_59 & ~w12380;
assign w24840 = ~w24838 & ~w24839;
assign w24841 = w24798 & ~w24840;
assign w24842 = ~w24798 & w24840;
assign w24843 = (w24810 & w32842) | (w24810 & w32843) | (w32842 & w32843);
assign w24844 = ~w24837 & ~w24843;
assign w24845 = (~w24810 & w32844) | (~w24810 & w32845) | (w32844 & w32845);
assign w24846 = ~w24810 & w32846;
assign w24847 = ~w24844 & ~w24846;
assign w24848 = b_62 & w11620;
assign w24849 = w11969 & w32847;
assign w24850 = b_61 & w11615;
assign w24851 = ~w24849 & ~w24850;
assign w24852 = ~w24848 & w24851;
assign w24853 = (w24852 & ~w12273) | (w24852 & w32848) | (~w12273 & w32848);
assign w24854 = a_62 & ~w24853;
assign w24855 = w24853 & a_62;
assign w24856 = ~w24853 & ~w24854;
assign w24857 = ~w24855 & ~w24856;
assign w24858 = w10902 & w32849;
assign w24859 = (~w24858 & ~w12670) | (~w24858 & w32850) | (~w12670 & w32850);
assign w24860 = a_59 & ~w24859;
assign w24861 = w24859 & a_59;
assign w24862 = ~w24859 & ~w24860;
assign w24863 = ~w24861 & ~w24862;
assign w24864 = ~w24857 & ~w24863;
assign w24865 = ~w24857 & ~w24864;
assign w24866 = w24857 & ~w24863;
assign w24867 = ~w24865 & ~w24866;
assign w24868 = ~w24847 & w24867;
assign w24869 = w24847 & ~w24867;
assign w24870 = ~w24868 & ~w24869;
assign w24871 = ~w24836 & ~w24870;
assign w24872 = ~w24836 & ~w24871;
assign w24873 = ~w24870 & ~w24871;
assign w24874 = ~w24872 & ~w24873;
assign w24875 = (~w13761 & w37834) | (~w13761 & w37835) | (w37834 & w37835);
assign w24876 = (w13761 & w37836) | (w13761 & w37837) | (w37836 & w37837);
assign w24877 = ~w24875 & ~w24876;
assign w24878 = (~w24864 & w24867) | (~w24864 & w32851) | (w24867 & w32851);
assign w24879 = a_59 & ~w24840;
assign w24880 = ~a_59 & w24840;
assign w24881 = ~w24879 & ~w24880;
assign w24882 = w12380 & w32852;
assign w24883 = b_60 & ~w12380;
assign w24884 = ~w24882 & ~w24883;
assign w24885 = w24881 & w24884;
assign w24886 = ~w24881 & ~w24884;
assign w24887 = ~w24885 & ~w24886;
assign w24888 = b_63 & w11620;
assign w24889 = w11969 & w32853;
assign w24890 = b_62 & w11615;
assign w24891 = ~w24889 & ~w24890;
assign w24892 = ~w24888 & w24891;
assign w24893 = (w24892 & ~w12646) | (w24892 & w32854) | (~w12646 & w32854);
assign w24894 = a_62 & ~w24893;
assign w24895 = w24893 & a_62;
assign w24896 = ~w24893 & ~w24894;
assign w24897 = ~w24895 & ~w24896;
assign w24898 = (w24887 & w24896) | (w24887 & w32855) | (w24896 & w32855);
assign w24899 = w24887 & ~w24898;
assign w24900 = ~w24897 & ~w24898;
assign w24901 = ~w24899 & ~w24900;
assign w24902 = ~w24845 & ~w24901;
assign w24903 = w24845 & w24901;
assign w24904 = ~w24902 & ~w24903;
assign w24905 = ~w24878 & w24904;
assign w24906 = ~w24878 & ~w24905;
assign w24907 = w24904 & ~w24905;
assign w24908 = ~w24906 & ~w24907;
assign w24909 = (~w13761 & w37838) | (~w13761 & w37839) | (w37838 & w37839);
assign w24910 = (w13761 & w37840) | (w13761 & w37841) | (w37840 & w37841);
assign w24911 = ~w24909 & ~w24910;
assign w24912 = (~w24898 & w24901) | (~w24898 & w32856) | (w24901 & w32856);
assign w24913 = w12380 & w32857;
assign w24914 = b_61 & ~w12380;
assign w24915 = ~w24913 & ~w24914;
assign w24916 = ~a_59 & ~w24840;
assign w24917 = (~w24916 & w24881) | (~w24916 & w32858) | (w24881 & w32858);
assign w24918 = w24915 & ~w24917;
assign w24919 = ~w24915 & w24917;
assign w24920 = ~w24918 & ~w24919;
assign w24921 = w11969 & w32859;
assign w24922 = b_63 & w11615;
assign w24923 = ~w24921 & ~w24922;
assign w24924 = ~w11623 & w24923;
assign w24925 = ~w12671 & w32860;
assign w24926 = (a_62 & w24925) | (a_62 & w32861) | (w24925 & w32861);
assign w24927 = ~w24925 & w32862;
assign w24928 = ~w24926 & ~w24927;
assign w24929 = w24920 & ~w24928;
assign w24930 = ~w24920 & w24928;
assign w24931 = ~w24929 & ~w24930;
assign w24932 = (~w24901 & w32863) | (~w24901 & w32864) | (w32863 & w32864);
assign w24933 = ~w24912 & ~w24932;
assign w24934 = w24931 & ~w24932;
assign w24935 = ~w24933 & ~w24934;
assign w24936 = (~w13761 & w37842) | (~w13761 & w37843) | (w37842 & w37843);
assign w24937 = (w13761 & w37856) | (w13761 & w37857) | (w37856 & w37857);
assign w24938 = ~w24936 & ~w24937;
assign w24939 = (~w24918 & w24928) | (~w24918 & w32865) | (w24928 & w32865);
assign w24940 = w12380 & w32866;
assign w24941 = b_62 & ~w12380;
assign w24942 = ~w24940 & ~w24941;
assign w24943 = w24915 & ~w24942;
assign w24944 = ~w24915 & w24942;
assign w24945 = ~w24943 & ~w24944;
assign w24946 = w11969 & w32867;
assign w24947 = (w9770 & w32868) | (w9770 & w32869) | (w32868 & w32869);
assign w24948 = (a_62 & w24947) | (a_62 & w32870) | (w24947 & w32870);
assign w24949 = ~w24947 & w32871;
assign w24950 = ~w24948 & ~w24949;
assign w24951 = w24945 & ~w24950;
assign w24952 = ~w24945 & w24950;
assign w24953 = ~w24951 & ~w24952;
assign w24954 = ~w24939 & w24953;
assign w24955 = ~w24939 & ~w24954;
assign w24956 = w24939 & w24953;
assign w24957 = ~w24955 & ~w24956;
assign w24958 = (~w13761 & w37844) | (~w13761 & w37845) | (w37844 & w37845);
assign w24959 = (w13761 & w37846) | (w13761 & w37847) | (w37846 & w37847);
assign w24960 = ~w24958 & ~w24959;
assign w24961 = w12380 & w32875;
assign w24962 = b_63 & ~w12380;
assign w24963 = ~w24961 & ~w24962;
assign w24964 = ~a_62 & ~w24963;
assign w24965 = a_62 & w24963;
assign w24966 = ~w24964 & ~w24965;
assign w24967 = ~w24915 & w24966;
assign w24968 = w24915 & ~w24966;
assign w24969 = ~w24967 & ~w24968;
assign w24970 = (~w24950 & w32876) | (~w24950 & w32877) | (w32876 & w32877);
assign w24971 = (w24950 & w32878) | (w24950 & w32879) | (w32878 & w32879);
assign w24972 = ~w24970 & ~w24971;
assign w24973 = (~w13761 & w37848) | (~w13761 & w37849) | (w37848 & w37849);
assign w24974 = (w13761 & w37850) | (w13761 & w37851) | (w37850 & w37851);
assign w24975 = ~w24973 & ~w24974;
assign w24976 = (~w24964 & ~w24966) | (~w24964 & w32882) | (~w24966 & w32882);
assign w24977 = w12380 & w32883;
assign w24978 = ~w24976 & w24977;
assign w24979 = w24976 & ~w24977;
assign w24980 = ~w24978 & ~w24979;
assign w24981 = (w13761 & w37852) | (w13761 & w37853) | (w37852 & w37853);
assign w24982 = (~w13761 & w37854) | (~w13761 & w37855) | (w37854 & w37855);
assign w24983 = ~w24981 & ~w24982;
assign w24984 = w412 & b_0;
assign w24985 = w651 & b_0;
assign w24986 = w980 & b_0;
assign w24987 = w1289 & b_0;
assign w24988 = w1688 & b_0;
assign w24989 = w2152 & b_0;
assign w24990 = w35 & w25334;
assign w24991 = (w2291 & ~w2318) | (w2291 & w25335) | (~w2318 & w25335);
assign w24992 = w2192 & w2344;
assign w24993 = w2217 & w2367;
assign w24994 = ~w2303 & w25475;
assign w24995 = (~w2474 & w2303) | (~w2474 & w25476) | (w2303 & w25476);
assign w24996 = ~w2349 & w27257;
assign w24997 = w2532 & w32888;
assign w24998 = (a_26 & ~w2622) | (a_26 & w25336) | (~w2622 & w25336);
assign w24999 = ~w2511 & ~w2509;
assign w25000 = w2684 & w32889;
assign w25001 = ~w2517 & ~w2516;
assign w25002 = w2703 & w32890;
assign w25003 = w2721 & w32891;
assign w25004 = ~w2540 & w32892;
assign w25005 = ~w2659 & ~w2657;
assign w25006 = w2653 & ~w2817;
assign w25007 = w2633 & b_0;
assign w25008 = w2886 & w32893;
assign w25009 = ~w2711 & w26864;
assign w25010 = w3062 & w32894;
assign w25011 = w3222 & w32895;
assign w25012 = w3265 & w32896;
assign w25013 = w3283 & w32897;
assign w25014 = ~w3291 & w27373;
assign w25015 = w3209 & ~w3385;
assign w25016 = ~w3450 & ~w3449;
assign w25017 = ~w3490 & ~w3489;
assign w25018 = w3497 & w32898;
assign w25019 = w3327 & ~w3529;
assign w25020 = ~w3506 & ~w3505;
assign w25021 = w3435 & ~w3431;
assign w25022 = w3640 & w32899;
assign w25023 = w3696 & w32900;
assign w25024 = ~w3649 & ~w3648;
assign w25025 = w3873 & w32901;
assign w25026 = ~w3672 & ~w3670;
assign w25027 = w3891 & w32902;
assign w25028 = ~w3491 & w26865;
assign w25029 = w3909 & w32903;
assign w25030 = ~w3917 & ~w3916;
assign w25031 = w3926 & w32904;
assign w25032 = (w3727 & w3939) | (w3727 & w32905) | (w3939 & w32905);
assign w25033 = ~w3741 & ~w3740;
assign w25034 = w3984 & w32906;
assign w25035 = ~w4118 & ~w4117;
assign w25036 = ~w3934 & w27493;
assign w25037 = w4899 & w32907;
assign w25038 = ~w4854 & ~w4853;
assign w25039 = w4865 & w5104;
assign w25040 = w5382 & w32908;
assign w25041 = w5393 & w32909;
assign w25042 = w5346 & w5596;
assign w25043 = w5369 & w5617;
assign w25044 = w5637 & w32910;
assign w25045 = w5833 & w32911;
assign w25046 = ~w5842 & ~w5841;
assign w25047 = w6376 & w32912;
assign w25048 = w6639 & w32913;
assign w25049 = ~w6392 & w32914;
assign w25050 = w6420 & w6690;
assign w25051 = ~w6562 & ~w6560;
assign w25052 = ~w6941 & ~w6940;
assign w25053 = ~w6857 & w27258;
assign w25054 = ~w6821 & w27259;
assign w25055 = ~w7172 & ~w7171;
assign w25056 = w6882 & w7196;
assign w25057 = w7217 & w32915;
assign w25058 = ~w7243 & ~w7242;
assign w25059 = w6956 & w7261;
assign w25060 = ~w6995 & ~w6994;
assign w25061 = ~w7202 & ~w7201;
assign w25062 = ~w7190 & ~w7189;
assign w25063 = ~w7206 & ~w7498;
assign w25064 = w7206 & w7498;
assign w25065 = w7505 & w32916;
assign w25066 = w7523 & w32917;
assign w25067 = w7798 & w32918;
assign w25068 = ~w7513 & w26966;
assign w25069 = w7816 & w32919;
assign w25070 = w8102 & w32920;
assign w25071 = ~w8128 & ~w8127;
assign w25072 = w7844 & ~w7841;
assign w25073 = ~w8069 & ~w8068;
assign w25074 = w7904 & ~w8056;
assign w25075 = ~w8073 & ~w8409;
assign w25076 = w8073 & w8409;
assign w25077 = w8416 & w32921;
assign w25078 = w8434 & w32922;
assign w25079 = ~w8443 & ~w8442;
assign w25080 = w8717 & w32923;
assign w25081 = ~w8424 & w25477;
assign w25082 = w9035 & w32924;
assign w25083 = ~w9061 & ~w9060;
assign w25084 = (w8776 & w9084) | (w8776 & w32925) | (w9084 & w32925);
assign w25085 = w9118 & ~w9122;
assign w25086 = ~w8974 & w27121;
assign w25087 = w9384 & w32926;
assign w25088 = ~w9393 & ~w9392;
assign w25089 = ~w9301 & w26967;
assign w25090 = ~w9314 & ~w9312;
assign w25091 = w9724 & w32927;
assign w25092 = ~w9732 & ~w9731;
assign w25093 = w9415 & w9754;
assign w25094 = ~w9131 & ~w9130;
assign w25095 = w9439 & w9784;
assign w25096 = ~w9759 & w32928;
assign w25097 = ~w9748 & ~w9747;
assign w25098 = ~w9642 & w27122;
assign w25099 = (w9623 & w9977) | (w9623 & w25337) | (w9977 & w25337);
assign w25100 = w9659 & w10013;
assign w25101 = ~w9659 & ~w10013;
assign w25102 = w10064 & w32929;
assign w25103 = ~w10072 & ~w10071;
assign w25104 = w10081 & w32930;
assign w25105 = ~w10113 & ~w10112;
assign w25106 = ~w10097 & w32931;
assign w25107 = ~w10018 & w27197;
assign w25108 = ~w10118 & w26081;
assign w25109 = ~w10391 & w26741;
assign w25110 = (w10408 & ~w10778) | (w10408 & w25338) | (~w10778 & w25338);
assign w25111 = w10427 & w10810;
assign w25112 = ~w10821 & w26508;
assign w25113 = w10625 & ~w10621;
assign w25114 = (w10692 & w11022) | (w10692 & w25339) | (w11022 & w25339);
assign w25115 = (w10761 & w11080) | (w10761 & w27440) | (w11080 & w27440);
assign w25116 = ~w10473 & ~w10472;
assign w25117 = w11166 & w10472;
assign w25118 = w11166 & ~w25116;
assign w25119 = (w27242 & w27441) | (w27242 & w27442) | (w27441 & w27442);
assign w25120 = ~w10966 & w27443;
assign w25121 = ~w11001 & ~w10999;
assign w25122 = w11178 & w11535;
assign w25123 = ~w11445 & w27494;
assign w25124 = ~w11420 & w27260;
assign w25125 = ~w11462 & ~w11460;
assign w25126 = ~w11820 & w26082;
assign w25127 = w11770 & ~w11767;
assign w25128 = ~w12118 & ~w12117;
assign w25129 = ~w12171 & ~w12170;
assign w25130 = w11853 & w12206;
assign w25131 = w11911 & w12284;
assign w25132 = ~w12211 & w25478;
assign w25133 = ~w12229 & ~w12227;
assign w25134 = ~w12270 & ~w12269;
assign w25135 = w12654 & ~w12656;
assign w25136 = w12660 & ~w12657;
assign w25137 = ~w12542 & ~w12540;
assign w25138 = ~w12558 & ~w12557;
assign w25139 = ~w13033 & ~w13031;
assign w25140 = (~w13366 & w37658) | (~w13366 & w37659) | (w37658 & w37659);
assign w25141 = ~w13756 & ~w13755;
assign w25142 = ~w14122 & w32932;
assign w25143 = ~w14481 & w38070;
assign w25144 = w14834 & w14480;
assign w25145 = (w14834 & ~w14483) | (w14834 & w25144) | (~w14483 & w25144);
assign w25146 = w14832 & ~w15168;
assign w25147 = w15165 & ~w15506;
assign w25148 = ~w15503 & w15506;
assign w25149 = (~w15503 & ~w15165) | (~w15503 & w25148) | (~w15165 & w25148);
assign w25150 = ~w15844 & ~w25148;
assign w25151 = ~w15844 & ~w25149;
assign w25152 = w15841 & ~w16174;
assign w25153 = ~w16172 & w25719;
assign w25154 = (~w16171 & w16174) | (~w16171 & w25340) | (w16174 & w25340);
assign w25155 = ~w16489 & ~w25153;
assign w25156 = (~w16174 & w25720) | (~w16174 & w25721) | (w25720 & w25721);
assign w25157 = w16486 & ~w16803;
assign w25158 = ~w16801 & w32933;
assign w25159 = (~w16800 & w16803) | (~w16800 & w25341) | (w16803 & w25341);
assign w25160 = ~w17121 & ~w25158;
assign w25161 = (~w25341 & w32934) | (~w25341 & w32935) | (w32934 & w32935);
assign w25162 = (~w17118 & w25158) | (~w17118 & w25479) | (w25158 & w25479);
assign w25163 = (w25341 & w32936) | (w25341 & w32937) | (w32936 & w32937);
assign w25164 = ~w17417 & ~w17415;
assign w25165 = w17711 & w17415;
assign w25166 = w17711 & ~w25164;
assign w25167 = (w25490 & w32938) | (w25490 & w32939) | (w32938 & w32939);
assign w25168 = (~w17710 & ~w17711) | (~w17710 & w25342) | (~w17711 & w25342);
assign w25169 = ~w17990 & ~w17989;
assign w25170 = ~w18274 & w17989;
assign w25171 = (~w18274 & w17990) | (~w18274 & w25170) | (w17990 & w25170);
assign w25172 = (~w18271 & ~w17989) | (~w18271 & w32940) | (~w17989 & w32940);
assign w25173 = ~w18271 & ~w25171;
assign w25174 = ~w18548 & ~w25172;
assign w25175 = (~w18548 & w25171) | (~w18548 & w25480) | (w25171 & w25480);
assign w25176 = (~w18545 & w25172) | (~w18545 & w32941) | (w25172 & w32941);
assign w25177 = (~w25171 & w32941) | (~w25171 & w32942) | (w32941 & w32942);
assign w25178 = ~w18814 & w32943;
assign w25179 = w19079 & w18813;
assign w25180 = (w19079 & ~w18816) | (w19079 & w25179) | (~w18816 & w25179);
assign w25181 = (~w19077 & ~w19079) | (~w19077 & w26968) | (~w19079 & w26968);
assign w25182 = (w18816 & w32944) | (w18816 & w32945) | (w32944 & w32945);
assign w25183 = (~w26968 & w32946) | (~w26968 & w32947) | (w32946 & w32947);
assign w25184 = w19338 & ~w25182;
assign w25185 = (~w19337 & w25181) | (~w19337 & w32948) | (w25181 & w32948);
assign w25186 = (~w19337 & w25182) | (~w19337 & w32948) | (w25182 & w32948);
assign w25187 = (~w25181 & w25481) | (~w25181 & w32949) | (w25481 & w32949);
assign w25188 = (~w25182 & w32950) | (~w25182 & w32951) | (w32950 & w32951);
assign w25189 = (w25181 & w32952) | (w25181 & w32953) | (w32952 & w32953);
assign w25190 = (w25182 & w32954) | (w25182 & w32955) | (w32954 & w32955);
assign w25191 = w19831 & ~w19828;
assign w25192 = (w19828 & w20072) | (w19828 & w32956) | (w20072 & w32956);
assign w25193 = ~w20074 & ~w25191;
assign w25194 = (~w20071 & w20074) | (~w20071 & w25482) | (w20074 & w25482);
assign w25195 = (~w20071 & w25191) | (~w20071 & w25343) | (w25191 & w25343);
assign w25196 = (~w20074 & w32957) | (~w20074 & w32958) | (w32957 & w32958);
assign w25197 = ~w20308 & ~w25195;
assign w25198 = ~w20305 & ~w25196;
assign w25199 = (~w20305 & w25195) | (~w20305 & w25483) | (w25195 & w25483);
assign w25200 = (w20535 & w25196) | (w20535 & w26866) | (w25196 & w26866);
assign w25201 = (~w25195 & w26866) | (~w25195 & w32959) | (w26866 & w32959);
assign w25202 = (~w25196 & w26867) | (~w25196 & w26971) | (w26867 & w26971);
assign w25203 = (w25195 & w32960) | (w25195 & w32961) | (w32960 & w32961);
assign w25204 = (w25196 & w26973) | (w25196 & w32962) | (w26973 & w32962);
assign w25205 = (~w25195 & w32963) | (~w25195 & w32964) | (w32963 & w32964);
assign w25206 = w20753 & w20970;
assign w25207 = ~w20969 & ~w20970;
assign w25208 = (~w20969 & ~w20970) | (~w20969 & w25344) | (~w20970 & w25344);
assign w25209 = (~w21183 & w20970) | (~w21183 & w25484) | (w20970 & w25484);
assign w25210 = (~w25344 & w25484) | (~w25344 & w32965) | (w25484 & w32965);
assign w25211 = ~w21180 & ~w25209;
assign w25212 = (w25344 & w32966) | (w25344 & w32967) | (w32966 & w32967);
assign w25213 = (w21389 & w25209) | (w21389 & w26742) | (w25209 & w26742);
assign w25214 = (~w25208 & w26742) | (~w25208 & w26743) | (w26742 & w26743);
assign w25215 = (~w25209 & w26868) | (~w25209 & w26869) | (w26868 & w26869);
assign w25216 = (w25208 & w26869) | (w25208 & w32968) | (w26869 & w32968);
assign w25217 = (w25209 & w32969) | (w25209 & w32970) | (w32969 & w32970);
assign w25218 = ~w21584 & ~w25216;
assign w25219 = (~w25209 & w32971) | (~w25209 & w32972) | (w32971 & w32972);
assign w25220 = (~w21581 & w25216) | (~w21581 & w26870) | (w25216 & w26870);
assign w25221 = (w25209 & w32973) | (w25209 & w32974) | (w32973 & w32974);
assign w25222 = (~w25216 & w26974) | (~w25216 & w32975) | (w26974 & w32975);
assign w25223 = ~w21777 & ~w25221;
assign w25224 = (w25216 & w32976) | (w25216 & w32977) | (w32976 & w32977);
assign w25225 = ~w21962 & ~w21960;
assign w25226 = ~w22143 & w21960;
assign w25227 = ~w22143 & ~w25225;
assign w25228 = (~w22140 & w25225) | (~w22140 & w32978) | (w25225 & w32978);
assign w25229 = (~w22140 & w22143) | (~w22140 & w25346) | (w22143 & w25346);
assign w25230 = (~w22143 & w25486) | (~w22143 & w25487) | (w25486 & w25487);
assign w25231 = (~w25345 & w32979) | (~w25345 & w32980) | (w32979 & w32980);
assign w25232 = (w25345 & w32981) | (w25345 & w32982) | (w32981 & w32982);
assign w25233 = (~w25487 & w32983) | (~w25487 & w32984) | (w32983 & w32984);
assign w25234 = (w25487 & w32985) | (w25487 & w32986) | (w32985 & w32986);
assign w25235 = (~w25345 & w32987) | (~w25345 & w32988) | (w32987 & w32988);
assign w25236 = (w25345 & w32989) | (w25345 & w32990) | (w32989 & w32990);
assign w25237 = (~w25487 & w32991) | (~w25487 & w32992) | (w32991 & w32992);
assign w25238 = w22662 & ~w25237;
assign w25239 = w22662 & ~w25236;
assign w25240 = (~w22661 & w25236) | (~w22661 & w26871) | (w25236 & w26871);
assign w25241 = (~w22661 & w25237) | (~w22661 & w26871) | (w25237 & w26871);
assign w25242 = (~w25237 & w26976) | (~w25237 & w26977) | (w26976 & w26977);
assign w25243 = (~w25236 & w26976) | (~w25236 & w26977) | (w26976 & w26977);
assign w25244 = (w25236 & w32993) | (w25236 & w32994) | (w32993 & w32994);
assign w25245 = (w25237 & w32993) | (w25237 & w32994) | (w32993 & w32994);
assign w25246 = ~w22980 & ~w22978;
assign w25247 = w23127 & w22978;
assign w25248 = (w23127 & w22980) | (w23127 & w25247) | (w22980 & w25247);
assign w25249 = ~w23126 & ~w25248;
assign w25250 = (~w23126 & ~w22978) | (~w23126 & w32995) | (~w22978 & w32995);
assign w25251 = w23272 & ~w25250;
assign w25252 = (w23272 & w25248) | (w23272 & w25347) | (w25248 & w25347);
assign w25253 = (~w25248 & w25488) | (~w25248 & w32996) | (w25488 & w32996);
assign w25254 = (~w23270 & w25250) | (~w23270 & w25488) | (w25250 & w25488);
assign w25255 = (~w25250 & w25489) | (~w25250 & w32997) | (w25489 & w32997);
assign w25256 = (w25248 & w32998) | (w25248 & w32999) | (w32998 & w32999);
assign w25257 = (~w25248 & w33000) | (~w25248 & w33001) | (w33000 & w33001);
assign w25258 = (w25250 & w33002) | (w25250 & w33003) | (w33002 & w33003);
assign w25259 = (~w25250 & w33004) | (~w25250 & w33005) | (w33004 & w33005);
assign w25260 = (w25248 & w33006) | (w25248 & w33007) | (w33006 & w33007);
assign w25261 = (~w25248 & w33008) | (~w25248 & w33009) | (w33008 & w33009);
assign w25262 = (w25250 & w33010) | (w25250 & w33011) | (w33010 & w33011);
assign w25263 = (~w25250 & w33012) | (~w25250 & w33013) | (w33012 & w33013);
assign w25264 = (w25248 & w33014) | (w25248 & w33015) | (w33014 & w33015);
assign w25265 = (~w25248 & w33016) | (~w25248 & w33017) | (w33016 & w33017);
assign w25266 = ~w23674 & ~w25263;
assign w25267 = (w23798 & w25263) | (w23798 & w26872) | (w25263 & w26872);
assign w25268 = (w25248 & w33018) | (w25248 & w33019) | (w33018 & w33019);
assign w25269 = ~w23796 & ~w25268;
assign w25270 = (~w25263 & w26978) | (~w25263 & w26979) | (w26978 & w26979);
assign w25271 = (w25263 & w33020) | (w25263 & w33021) | (w33020 & w33021);
assign w25272 = (w23910 & w25268) | (w23910 & w26980) | (w25268 & w26980);
assign w25273 = w23909 & w24022;
assign w25274 = ~w24021 & ~w24022;
assign w25275 = (~w24021 & ~w24022) | (~w24021 & w25348) | (~w24022 & w25348);
assign w25276 = (w24125 & w24022) | (w24125 & w25722) | (w24022 & w25722);
assign w25277 = (~w25348 & w25722) | (~w25348 & w33022) | (w25722 & w33022);
assign w25278 = ~w24124 & ~w25276;
assign w25279 = (w25348 & w33023) | (w25348 & w33024) | (w33023 & w33024);
assign w25280 = (w24222 & w25276) | (w24222 & w26085) | (w25276 & w26085);
assign w25281 = (~w25275 & w26085) | (~w25275 & w26086) | (w26085 & w26086);
assign w25282 = (~w25276 & w33025) | (~w25276 & w33026) | (w33025 & w33026);
assign w25283 = (w25275 & w33026) | (w25275 & w33027) | (w33026 & w33027);
assign w25284 = (w25276 & w33028) | (w25276 & w33029) | (w33028 & w33029);
assign w25285 = (~w25275 & w33029) | (~w25275 & w33030) | (w33029 & w33030);
assign w25286 = (~w25276 & w33031) | (~w25276 & w33032) | (w33031 & w33032);
assign w25287 = (w25275 & w33032) | (w25275 & w33033) | (w33032 & w33033);
assign w25288 = (w25276 & w33034) | (w25276 & w33035) | (w33034 & w33035);
assign w25289 = w24400 & ~w25287;
assign w25290 = (~w25276 & w33036) | (~w25276 & w33037) | (w33036 & w33037);
assign w25291 = (~w24399 & w25287) | (~w24399 & w26874) | (w25287 & w26874);
assign w25292 = (w25276 & w33038) | (w25276 & w33039) | (w33038 & w33039);
assign w25293 = (~w25287 & w26981) | (~w25287 & w26982) | (w26981 & w26982);
assign w25294 = ~w24475 & ~w25292;
assign w25295 = (w25287 & w33040) | (w25287 & w33041) | (w33040 & w33041);
assign w25296 = (w24549 & w25292) | (w24549 & w33042) | (w25292 & w33042);
assign w25297 = (~w25287 & w33043) | (~w25287 & w33044) | (w33043 & w33044);
assign w25298 = w24548 & w24619;
assign w25299 = ~w24617 & ~w24619;
assign w25300 = (~w24617 & ~w24548) | (~w24617 & w25299) | (~w24548 & w25299);
assign w25301 = ~w24682 & ~w25299;
assign w25302 = ~w24682 & ~w25300;
assign w25303 = ~w24679 & ~w25301;
assign w25304 = (~w24679 & w25300) | (~w24679 & w33045) | (w25300 & w33045);
assign w25305 = (w24739 & w25301) | (w24739 & w25724) | (w25301 & w25724);
assign w25306 = (~w25300 & w33046) | (~w25300 & w33047) | (w33046 & w33047);
assign w25307 = (~w25301 & w26087) | (~w25301 & w26088) | (w26087 & w26088);
assign w25308 = (w25300 & w33048) | (w25300 & w33049) | (w33048 & w33049);
assign w25309 = (w25301 & w33050) | (w25301 & w33051) | (w33050 & w33051);
assign w25310 = w24791 & ~w25308;
assign w25311 = (~w25301 & w33052) | (~w25301 & w33053) | (w33052 & w33053);
assign w25312 = (~w24790 & w25308) | (~w24790 & w26513) | (w25308 & w26513);
assign w25313 = w24832 & ~w25311;
assign w25314 = (~w25308 & w33054) | (~w25308 & w33055) | (w33054 & w33055);
assign w25315 = (~w24831 & w25311) | (~w24831 & w26751) | (w25311 & w26751);
assign w25316 = (w25308 & w26983) | (w25308 & w26984) | (w26983 & w26984);
assign w25317 = (~w25311 & w33056) | (~w25311 & w33057) | (w33056 & w33057);
assign w25318 = (~w25308 & w33058) | (~w25308 & w33059) | (w33058 & w33059);
assign w25319 = (w25311 & w33060) | (w25311 & w33061) | (w33060 & w33061);
assign w25320 = (w25308 & w33062) | (w25308 & w33063) | (w33062 & w33063);
assign w25321 = (~w25311 & w33064) | (~w25311 & w33065) | (w33064 & w33065);
assign w25322 = (~w25308 & w33066) | (~w25308 & w33067) | (w33066 & w33067);
assign w25323 = (w25311 & w33068) | (w25311 & w33069) | (w33068 & w33069);
assign w25324 = (w25308 & w33070) | (w25308 & w33071) | (w33070 & w33071);
assign w25325 = (~w25311 & w33072) | (~w25311 & w33073) | (w33072 & w33073);
assign w25326 = ~w24935 & ~w25324;
assign w25327 = w24932 & ~w24957;
assign w25328 = ~w24955 & w33074;
assign w25329 = ~w24954 & ~w25327;
assign w25330 = w24972 & ~w25328;
assign w25331 = (w24972 & w25327) | (w24972 & w33075) | (w25327 & w33075);
assign w25332 = (~w24970 & w25328) | (~w24970 & w33076) | (w25328 & w33076);
assign w25333 = (~w25327 & w33076) | (~w25327 & w33077) | (w33076 & w33077);
assign w25334 = w2161 & a_26;
assign w25335 = w2307 & w2291;
assign w25336 = w2158 & w33078;
assign w25337 = w9612 & w27261;
assign w25338 = w10768 & w10408;
assign w25339 = w10681 & w27262;
assign w25340 = ~w15841 & ~w16171;
assign w25341 = ~w16486 & ~w16800;
assign w25342 = (~w17415 & w17707) | (~w17415 & w25491) | (w17707 & w25491);
assign w25343 = ~w20072 & w33079;
assign w25344 = ~w20753 & ~w20969;
assign w25345 = ~w21962 & w25346;
assign w25346 = ~w21960 & ~w22140;
assign w25347 = w23126 & w23272;
assign w25348 = ~w23909 & ~w24021;
assign w25349 = ~w54 & ~w53;
assign w25350 = w93 & b_0;
assign w25351 = w233 & b_0;
assign w25352 = w421 & w25725;
assign w25353 = w35 & w25726;
assign w25354 = w660 & w25492;
assign w25355 = w35 & w25493;
assign w25356 = w989 & w25494;
assign w25357 = w35 & w25495;
assign w25358 = w1298 & w25496;
assign w25359 = w35 & w25497;
assign w25360 = w1697 & w25498;
assign w25361 = w35 & w25499;
assign w25362 = w2161 & w25500;
assign w25363 = ~w24990 & a_26;
assign w25364 = w2488 & ~w2617;
assign w25365 = w2642 & w25501;
assign w25366 = w35 & w25502;
assign w25367 = w3189 & b_0;
assign w25368 = w3797 & b_0;
assign w25369 = w4493 & b_0;
assign w25370 = w5190 & b_0;
assign w25371 = w5956 & b_0;
assign w25372 = w7607 & b_0;
assign w25373 = w35 & w25503;
assign w25374 = (w7626 & w7967) | (w7626 & w26985) | (w7967 & w26985);
assign w25375 = ~w7967 & w26986;
assign w25376 = w7649 & w7991;
assign w25377 = (w7708 & w8027) | (w7708 & w26875) | (w8027 & w26875);
assign w25378 = w7751 & w8069;
assign w25379 = ~w7751 & ~w8069;
assign w25380 = w8084 & w33080;
assign w25381 = (a_11 & ~w8102) | (a_11 & w33081) | (~w8102 & w33081);
assign w25382 = a_11 & ~w25070;
assign w25383 = w8120 & w33082;
assign w25384 = w8137 & w33083;
assign w25385 = ~w7856 & ~w7855;
assign w25386 = (~w7855 & ~w7856) | (~w7855 & w33084) | (~w7856 & w33084);
assign w25387 = ~w7867 & ~w7866;
assign w25388 = (~w7866 & ~w7867) | (~w7866 & w25727) | (~w7867 & w25727);
assign w25389 = w8196 & w33085;
assign w25390 = w8207 & w33086;
assign w25391 = ~w8063 & ~w8062;
assign w25392 = ~w8004 & w26987;
assign w25393 = ~w7975 & w33087;
assign w25394 = ~w7950 & w25728;
assign w25395 = (~w8272 & w7950) | (~w8272 & w25729) | (w7950 & w25729);
assign w25396 = w8400 & w33088;
assign w25397 = (a_14 & ~w8416) | (a_14 & w33089) | (~w8416 & w33089);
assign w25398 = a_14 & ~w25077;
assign w25399 = (a_11 & ~w8434) | (a_11 & w33090) | (~w8434 & w33090);
assign w25400 = a_11 & ~w25078;
assign w25401 = ~w8391 & w27263;
assign w25402 = w8699 & w33091;
assign w25403 = (a_14 & ~w8717) | (a_14 & w33092) | (~w8717 & w33092);
assign w25404 = a_14 & ~w25080;
assign w25405 = w8735 & w33093;
assign w25406 = ~w8743 & ~w8742;
assign w25407 = w8751 & w33094;
assign w25408 = w8520 & b_0;
assign w25409 = w9017 & w33095;
assign w25410 = ~w8707 & w26876;
assign w25411 = (a_14 & ~w9035) | (a_14 & w33096) | (~w9035 & w33096);
assign w25412 = a_14 & ~w25082;
assign w25413 = w9053 & w33097;
assign w25414 = w9070 & w33098;
assign w25415 = w9143 & w33099;
assign w25416 = ~w9044 & w26752;
assign w25417 = w9366 & w33100;
assign w25418 = (a_14 & ~w9384) | (a_14 & w33101) | (~w9384 & w33101);
assign w25419 = a_14 & ~w25087;
assign w25420 = w9459 & w33102;
assign w25421 = w9706 & w33103;
assign w25422 = (a_14 & ~w9724) | (a_14 & w33104) | (~w9724 & w33104);
assign w25423 = a_14 & ~w25091;
assign w25424 = w9739 & w33105;
assign w25425 = w10046 & w33106;
assign w25426 = (a_14 & ~w10064) | (a_14 & w33107) | (~w10064 & w33107);
assign w25427 = a_14 & ~w25102;
assign w25428 = (a_11 & ~w10081) | (a_11 & w33108) | (~w10081 & w33108);
assign w25429 = a_11 & ~w25104;
assign w25430 = w10151 & w33109;
assign w25431 = w10161 & w33110;
assign w25432 = w10382 & w33111;
assign w25433 = w10754 & w33112;
assign w25434 = w11084 & w33113;
assign w25435 = w11118 & w33114;
assign w25436 = w11811 & w33115;
assign w25437 = w12197 & w33116;
assign w25438 = (w9770 & w33117) | (w9770 & w33118) | (w33117 & w33118);
assign w25439 = ~w12258 & w12259;
assign w25440 = w12258 & ~w12259;
assign w25441 = ~w11898 & ~w11897;
assign w25442 = (~w11897 & ~w11898) | (~w11897 & w33119) | (~w11898 & w33119);
assign w25443 = ~w1298 & w12316;
assign w25444 = w12156 & ~w12152;
assign w25445 = w12138 & ~w12134;
assign w25446 = (~w12187 & w12569) | (~w12187 & w25504) | (w12569 & w25504);
assign w25447 = ~w12282 & ~w12284;
assign w25448 = (~w12282 & ~w12284) | (~w12282 & w25730) | (~w12284 & w25730);
assign w25449 = ~w12570 & w26089;
assign w25450 = ~w12518 & ~w12517;
assign w25451 = w12944 & w33120;
assign w25452 = ~w13399 & ~w13398;
assign w25453 = (w9770 & w33121) | (w9770 & w33122) | (w33121 & w33122);
assign w25454 = ~w660 & w14159;
assign w25455 = ~w14428 & ~w14429;
assign w25456 = w14906 & w33123;
assign w25457 = ~w15424 & ~w15425;
assign w25458 = w15895 & w33124;
assign w25459 = ~w17180 & ~w17181;
assign w25460 = w21701 & w33125;
assign w25461 = w21859 & w33126;
assign w25462 = w21875 & w33127;
assign w25463 = w22365 & w33128;
assign w25464 = w22384 & w33129;
assign w25465 = w22402 & w33130;
assign w25466 = w22557 & w33131;
assign w25467 = w22574 & w33132;
assign w25468 = w22869 & w33133;
assign w25469 = w23856 & w33134;
assign w25470 = (~w7859 & w33135) | (~w7859 & w33136) | (w33135 & w33136);
assign w25471 = w24445 & w33137;
assign w25472 = (w25311 & w33138) | (w25311 & w33139) | (w33138 & w33139);
assign w25473 = (w25311 & w33142) | (w25311 & w33143) | (w33142 & w33143);
assign w25474 = (w25311 & w33145) | (w25311 & w33146) | (w33145 & w33146);
assign w25475 = ~w2302 & w2474;
assign w25476 = w2302 & ~w2474;
assign w25477 = ~w8425 & ~w8423;
assign w25478 = ~w12212 & ~w12210;
assign w25479 = w17121 & ~w17118;
assign w25480 = w18271 & ~w18548;
assign w25481 = w19337 & w19582;
assign w25482 = ~w19828 & ~w20071;
assign w25483 = ~w20306 & w33147;
assign w25484 = w20969 & ~w21183;
assign w25485 = ~w21181 & w33148;
assign w25486 = w22321 & w22140;
assign w25487 = (w22321 & w21960) | (w22321 & w25486) | (w21960 & w25486);
assign w25488 = ~w23272 & ~w23270;
assign w25489 = w23270 & w23413;
assign w25490 = ~w17417 & w25491;
assign w25491 = w17708 & ~w17415;
assign w25492 = ~w15 & a_14;
assign w25493 = w660 & a_14;
assign w25494 = ~w15 & a_17;
assign w25495 = w989 & a_17;
assign w25496 = ~w15 & a_20;
assign w25497 = w1298 & a_20;
assign w25498 = ~w15 & a_23;
assign w25499 = w1697 & a_23;
assign w25500 = ~w15 & a_26;
assign w25501 = ~w15 & a_29;
assign w25502 = w2642 & a_29;
assign w25503 = w7616 & a_50;
assign w25504 = ~w12568 & ~w12187;
assign w25505 = w421 & ~w25117;
assign w25506 = w421 & ~w25118;
assign w25507 = ~w81 & ~w80;
assign w25508 = ~w25354 & a_14;
assign w25509 = w664 & w648;
assign w25510 = ~w25355 & a_14;
assign w25511 = ~w666 & w868;
assign w25512 = w666 & ~w868;
assign w25513 = ~w25356 & a_17;
assign w25514 = w993 & w977;
assign w25515 = ~w25357 & a_17;
assign w25516 = ~w995 & w1175;
assign w25517 = w995 & ~w1175;
assign w25518 = ~w25358 & a_20;
assign w25519 = w1302 & w1286;
assign w25520 = ~w25359 & a_20;
assign w25521 = ~w1304 & w1553;
assign w25522 = w1304 & ~w1553;
assign w25523 = ~w25360 & a_23;
assign w25524 = w1701 & w1685;
assign w25525 = ~w25361 & a_23;
assign w25526 = ~w1703 & w1994;
assign w25527 = w1703 & ~w1994;
assign w25528 = ~w25362 & a_26;
assign w25529 = w2165 & w2149;
assign w25530 = w2152 & b_1;
assign w25531 = w2167 & w2474;
assign w25532 = w2152 & b_2;
assign w25533 = w2622 & w33149;
assign w25534 = ~w25365 & a_29;
assign w25535 = w2646 & w2630;
assign w25536 = ~w2646 & ~w2630;
assign w25537 = ~w25366 & a_29;
assign w25538 = ~w2846 & ~w2845;
assign w25539 = ~w2648 & w3004;
assign w25540 = w2648 & ~w3004;
assign w25541 = w2633 & b_2;
assign w25542 = (a_29 & ~w3178) | (a_29 & w25731) | (~w3178 & w25731);
assign w25543 = w3198 & w25732;
assign w25544 = w35 & w25733;
assign w25545 = w3806 & w25734;
assign w25546 = w35 & w25735;
assign w25547 = w4502 & w25736;
assign w25548 = w35 & w25737;
assign w25549 = w5199 & w25738;
assign w25550 = w35 & w25739;
assign w25551 = w5965 & w25740;
assign w25552 = w35 & w25741;
assign w25553 = w6755 & b_0;
assign w25554 = w7616 & w25742;
assign w25555 = ~w25373 & a_50;
assign w25556 = w8286 & ~w8504;
assign w25557 = w8529 & w25743;
assign w25558 = w35 & w25744;
assign w25559 = w8539 & ~w8912;
assign w25560 = (w8619 & w8974) | (w8619 & w27495) | (w8974 & w27495);
assign w25561 = (a_17 & ~w9017) | (a_17 & w33150) | (~w9017 & w33150);
assign w25562 = a_17 & ~w25409;
assign w25563 = w9035 & w33151;
assign w25564 = a_14 & w25082;
assign w25565 = (~w9096 & w25084) | (~w9096 & ~w8779) | (w25084 & ~w8779);
assign w25566 = ~w8790 & ~w8789;
assign w25567 = (~w8789 & ~w8790) | (~w8789 & w33152) | (~w8790 & w33152);
assign w25568 = a_11 & ~w9144;
assign w25569 = a_11 & ~w25415;
assign w25570 = ~w9002 & ~w9001;
assign w25571 = ~w8996 & ~w8995;
assign w25572 = ~w8990 & ~w8989;
assign w25573 = ~w8949 & w26988;
assign w25574 = w9200 & w33153;
assign w25575 = ~w8941 & w27264;
assign w25576 = ~w8930 & ~w8929;
assign w25577 = w9333 & w33154;
assign w25578 = (a_17 & ~w9366) | (a_17 & w33155) | (~w9366 & w33155);
assign w25579 = a_17 & ~w25417;
assign w25580 = a_14 & ~w25418;
assign w25581 = w25087 & a_14;
assign w25582 = w9441 & w9122;
assign w25583 = w9441 & ~w25085;
assign w25584 = w9267 & ~w9512;
assign w25585 = (~w9312 & ~w9314) | (~w9312 & w25745) | (~w9314 & w25745);
assign w25586 = (~w9312 & w25090) | (~w9312 & w25086) | (w25090 & w25086);
assign w25587 = w9688 & w33156;
assign w25588 = ~w9359 & ~w9357;
assign w25589 = (a_17 & ~w9706) | (a_17 & w33157) | (~w9706 & w33157);
assign w25590 = a_17 & ~w25421;
assign w25591 = a_14 & ~w25422;
assign w25592 = w25091 & a_14;
assign w25593 = (a_11 & ~w9739) | (a_11 & w33158) | (~w9739 & w33158);
assign w25594 = a_11 & ~w25424;
assign w25595 = w9820 & w33159;
assign w25596 = w9830 & w33160;
assign w25597 = w9528 & b_0;
assign w25598 = w10028 & w33161;
assign w25599 = (a_17 & ~w10046) | (a_17 & w33162) | (~w10046 & w33162);
assign w25600 = a_17 & ~w25425;
assign w25601 = ~w9715 & w26753;
assign w25602 = a_14 & ~w25426;
assign w25603 = w25102 & a_14;
assign w25604 = a_11 & ~w25428;
assign w25605 = w25104 & a_11;
assign w25606 = (w25097 & w27496) | (w25097 & w27497) | (w27496 & w27497);
assign w25607 = (a_11 & ~w10151) | (a_11 & w33163) | (~w10151 & w33163);
assign w25608 = a_11 & ~w25430;
assign w25609 = (a_14 & ~w10161) | (a_14 & w33164) | (~w10161 & w33164);
assign w25610 = a_14 & ~w25431;
assign w25611 = w10349 & w33165;
assign w25612 = (a_20 & ~w10382) | (a_20 & w33166) | (~w10382 & w33166);
assign w25613 = a_20 & ~w25432;
assign w25614 = w10400 & w33167;
assign w25615 = w10506 & w33168;
assign w25616 = w10736 & w33169;
assign w25617 = (a_20 & ~w10754) | (a_20 & w33170) | (~w10754 & w33170);
assign w25618 = a_20 & ~w25433;
assign w25619 = w10772 & w33171;
assign w25620 = w10789 & w33172;
assign w25621 = w11066 & w33173;
assign w25622 = (a_20 & ~w11084) | (a_20 & w33174) | (~w11084 & w33174);
assign w25623 = a_20 & ~w25434;
assign w25624 = w11101 & w33175;
assign w25625 = (a_14 & ~w11118) | (a_14 & w33176) | (~w11118 & w33176);
assign w25626 = a_14 & ~w25435;
assign w25627 = w11238 & w33177;
assign w25628 = w11249 & w33178;
assign w25629 = w11261 & w33179;
assign w25630 = w11469 & w33180;
assign w25631 = w11487 & w33181;
assign w25632 = w11760 & w33182;
assign w25633 = w11793 & w33183;
assign w25634 = (a_23 & ~w11811) | (a_23 & w33184) | (~w11811 & w33184);
assign w25635 = a_23 & ~w25436;
assign w25636 = w12163 & w33185;
assign w25637 = w12180 & w33186;
assign w25638 = (a_17 & ~w12197) | (a_17 & w33187) | (~w12197 & w33187);
assign w25639 = a_17 & ~w25437;
assign w25640 = w12303 & w33188;
assign w25641 = (a_20 & ~w12315) | (a_20 & w33189) | (~w12315 & w33189);
assign w25642 = (a_20 & ~w12316) | (a_20 & w25497) | (~w12316 & w25497);
assign w25643 = w12325 & w33190;
assign w25644 = w12337 & w33191;
assign w25645 = w12549 & w33192;
assign w25646 = w12706 & w33193;
assign w25647 = w12717 & w33194;
assign w25648 = w12926 & w33195;
assign w25649 = (a_26 & ~w12944) | (a_26 & w33196) | (~w12944 & w33196);
assign w25650 = a_26 & ~w25451;
assign w25651 = w13052 & w33197;
assign w25652 = w14051 & w33198;
assign w25653 = w15230 & w33199;
assign w25654 = a_29 & w15425;
assign w25655 = a_29 & ~w25457;
assign w25656 = ~a_29 & ~w15425;
assign w25657 = ~a_29 & w25457;
assign w25658 = (a_26 & ~w15895) | (a_26 & w33200) | (~w15895 & w33200);
assign w25659 = a_26 & ~w25458;
assign w25660 = a_26 & ~w25658;
assign w25661 = w25458 & a_26;
assign w25662 = w15801 & ~w15593;
assign w25663 = ~w16110 & ~w16111;
assign w25664 = w15905 & ~w16121;
assign w25665 = w15826 & ~w15564;
assign w25666 = (~w15525 & w33201) | (~w15525 & w33202) | (w33201 & w33202);
assign w25667 = (w16125 & w15888) | (w16125 & w33203) | (w15888 & w33203);
assign w25668 = ~w16234 & ~w16235;
assign w25669 = w16245 & w33204;
assign w25670 = ~w16460 & ~w16461;
assign w25671 = a_32 & w17181;
assign w25672 = a_32 & ~w25459;
assign w25673 = ~a_32 & ~w17181;
assign w25674 = ~a_32 & w25459;
assign w25675 = w17769 & w33205;
assign w25676 = w20482 & w33206;
assign w25677 = w20680 & w33207;
assign w25678 = w21120 & w33208;
assign w25679 = w21301 & w33209;
assign w25680 = (a_50 & ~w21701) | (a_50 & w33210) | (~w21701 & w33210);
assign w25681 = a_50 & ~w25460;
assign w25682 = w21800 & w33211;
assign w25683 = (a_53 & ~w21859) | (a_53 & w33212) | (~w21859 & w33212);
assign w25684 = a_53 & ~w25461;
assign w25685 = (a_50 & ~w21875) | (a_50 & w33213) | (~w21875 & w33213);
assign w25686 = a_50 & ~w25462;
assign w25687 = w21892 & w33214;
assign w25688 = w22020 & w33215;
assign w25689 = (a_59 & ~w22365) | (a_59 & w33216) | (~w22365 & w33216);
assign w25690 = a_59 & ~w25463;
assign w25691 = (a_56 & ~w22384) | (a_56 & w33217) | (~w22384 & w33217);
assign w25692 = a_56 & ~w25464;
assign w25693 = (a_53 & ~w22402) | (a_53 & w33218) | (~w22402 & w33218);
assign w25694 = a_53 & ~w25465;
assign w25695 = w22512 & w33219;
assign w25696 = w22539 & w33220;
assign w25697 = (a_56 & ~w22557) | (a_56 & w33221) | (~w22557 & w33221);
assign w25698 = a_56 & ~w25466;
assign w25699 = (a_53 & ~w22574) | (a_53 & w33222) | (~w22574 & w33222);
assign w25700 = a_53 & ~w25467;
assign w25701 = w22592 & w33223;
assign w25702 = w22747 & w33224;
assign w25703 = (a_59 & ~w22869) | (a_59 & w33225) | (~w22869 & w33225);
assign w25704 = a_59 & ~w25468;
assign w25705 = w22888 & w33226;
assign w25706 = w23021 & w33227;
assign w25707 = w23038 & w33228;
assign w25708 = (a_62 & ~w23856) | (a_62 & w33229) | (~w23856 & w33229);
assign w25709 = a_62 & ~w25469;
assign w25710 = w23856 & w33230;
assign w25711 = a_62 & w25469;
assign w25712 = (w25287 & w33231) | (w25287 & w33232) | (w33231 & w33232);
assign w25713 = (w25287 & w33235) | (w25287 & w33236) | (w33235 & w33236);
assign w25714 = (w25287 & w33239) | (w25287 & w33240) | (w33239 & w33240);
assign w25715 = (~w25324 & w33243) | (~w25324 & w33244) | (w33243 & w33244);
assign w25716 = (~w25311 & w33245) | (~w25311 & w33246) | (w33245 & w33246);
assign w25717 = (~w25324 & w33247) | (~w25324 & w33248) | (w33247 & w33248);
assign w25718 = (~w25311 & w33249) | (~w25311 & w33250) | (w33249 & w33250);
assign w25719 = ~w16173 & ~w16171;
assign w25720 = ~w16489 & w16171;
assign w25721 = (~w16489 & w15841) | (~w16489 & w25720) | (w15841 & w25720);
assign w25722 = w24021 & w24125;
assign w25723 = ~w24125 & ~w24124;
assign w25724 = w24679 & w24739;
assign w25725 = ~w15 & a_11;
assign w25726 = w421 & a_11;
assign w25727 = (~w7552 & ~w7848) | (~w7552 & w33251) | (~w7848 & w33251);
assign w25728 = ~w7949 & w8272;
assign w25729 = w7949 & ~w8272;
assign w25730 = ~w11911 & ~w12282;
assign w25731 = w2639 & w33252;
assign w25732 = ~w15 & a_32;
assign w25733 = w3198 & a_32;
assign w25734 = ~w15 & a_35;
assign w25735 = w3806 & a_35;
assign w25736 = ~w15 & a_38;
assign w25737 = w4502 & a_38;
assign w25738 = ~w15 & a_41;
assign w25739 = w5199 & a_41;
assign w25740 = ~w15 & a_44;
assign w25741 = w5965 & a_44;
assign w25742 = ~w15 & a_50;
assign w25743 = ~w15 & a_53;
assign w25744 = w8529 & a_53;
assign w25745 = ~w9312 & ~w8972;
assign w25746 = w102 & w26090;
assign w25747 = w126 & w80;
assign w25748 = w126 & ~w25507;
assign w25749 = ~w126 & ~w80;
assign w25750 = ~w126 & w25507;
assign w25751 = ~w135 & ~w102;
assign w25752 = ~w135 & ~w35;
assign w25753 = w242 & w26091;
assign w25754 = w35 & w26092;
assign w25755 = ~w25352 & a_11;
assign w25756 = w425 & w409;
assign w25757 = ~w25353 & a_11;
assign w25758 = ~w427 & w571;
assign w25759 = w427 & ~w571;
assign w25760 = w651 & b_1;
assign w25761 = w651 & b_2;
assign w25762 = (a_14 & ~w969) | (a_14 & w26093) | (~w969 & w26093);
assign w25763 = ~w1000 & ~w999;
assign w25764 = w980 & b_1;
assign w25765 = w980 & b_2;
assign w25766 = (a_17 & ~w1278) | (a_17 & w26094) | (~w1278 & w26094);
assign w25767 = w1309 & ~w1419;
assign w25768 = w1289 & b_1;
assign w25769 = w1289 & b_2;
assign w25770 = (a_20 & ~w1677) | (a_20 & w26095) | (~w1677 & w26095);
assign w25771 = w1708 & ~w1831;
assign w25772 = w1688 & b_1;
assign w25773 = w1688 & b_2;
assign w25774 = (a_23 & ~w2141) | (a_23 & w26096) | (~w2141 & w26096);
assign w25775 = ~w2319 & ~w2320;
assign w25776 = ~w2319 & w24991;
assign w25777 = ~w25538 & ~w2845;
assign w25778 = w2633 & b_1;
assign w25779 = w3178 & w33253;
assign w25780 = ~w25543 & a_32;
assign w25781 = w3202 & w3186;
assign w25782 = ~w3202 & ~w3186;
assign w25783 = ~w25544 & a_32;
assign w25784 = ~w3414 & ~w3413;
assign w25785 = ~w3204 & w3596;
assign w25786 = w3204 & ~w3596;
assign w25787 = ~w25545 & a_35;
assign w25788 = w3810 & w3794;
assign w25789 = ~w25546 & a_35;
assign w25790 = ~w3812 & w4242;
assign w25791 = w3812 & ~w4242;
assign w25792 = ~w25547 & a_38;
assign w25793 = w4506 & w4490;
assign w25794 = ~w25548 & a_38;
assign w25795 = ~w4508 & w4943;
assign w25796 = w4508 & ~w4943;
assign w25797 = ~w25549 & a_41;
assign w25798 = w5203 & w5187;
assign w25799 = ~w25550 & a_41;
assign w25800 = ~w5205 & w5693;
assign w25801 = w5205 & ~w5693;
assign w25802 = ~w25551 & a_44;
assign w25803 = w5969 & w5953;
assign w25804 = ~w25552 & a_44;
assign w25805 = ~w5971 & w6483;
assign w25806 = w5971 & ~w6483;
assign w25807 = w6764 & w26097;
assign w25808 = w35 & w26098;
assign w25809 = ~w25554 & a_50;
assign w25810 = w7620 & w7604;
assign w25811 = w7607 & b_1;
assign w25812 = w7622 & w8272;
assign w25813 = w7607 & b_2;
assign w25814 = (a_50 & ~w8509) | (a_50 & w26099) | (~w8509 & w26099);
assign w25815 = ~w25557 & a_53;
assign w25816 = w8533 & w8517;
assign w25817 = ~w25558 & a_53;
assign w25818 = ~w8535 & w9253;
assign w25819 = w8535 & ~w9253;
assign w25820 = w8520 & b_1;
assign w25821 = w8535 & w9253;
assign w25822 = w8520 & b_2;
assign w25823 = (a_53 & ~w9517) | (a_53 & w26100) | (~w9517 & w26100);
assign w25824 = w9537 & w26101;
assign w25825 = w35 & w26102;
assign w25826 = w9547 & ~w9902;
assign w25827 = w9605 & w9974;
assign w25828 = w9981 & w33254;
assign w25829 = ~w9988 & w25099;
assign w25830 = ~w9988 & ~w9989;
assign w25831 = (a_20 & ~w10028) | (a_20 & w33255) | (~w10028 & w33255);
assign w25832 = a_20 & ~w25598;
assign w25833 = a_17 & ~w25599;
assign w25834 = w25425 & a_17;
assign w25835 = (w10110 & ~w9805) | (w10110 & w27265) | (~w9805 & w27265);
assign w25836 = w9805 & w27266;
assign w25837 = a_11 & ~w25607;
assign w25838 = w25430 & a_11;
assign w25839 = a_14 & ~w25609;
assign w25840 = w25431 & a_14;
assign w25841 = w10197 & w33256;
assign w25842 = ~w9931 & w27267;
assign w25843 = ~w9926 & ~w9925;
assign w25844 = (a_26 & ~w10349) | (a_26 & w33257) | (~w10349 & w33257);
assign w25845 = a_26 & ~w25611;
assign w25846 = w10366 & w33258;
assign w25847 = a_20 & ~w25612;
assign w25848 = w25432 & a_20;
assign w25849 = (a_17 & ~w10400) | (a_17 & w33259) | (~w10400 & w33259);
assign w25850 = a_17 & ~w25614;
assign w25851 = ~w9795 & ~w9794;
assign w25852 = (~w9794 & ~w9795) | (~w9794 & w33260) | (~w9795 & w33260);
assign w25853 = w10125 & w26989;
assign w25854 = ~w10436 & w33261;
assign w25855 = w10495 & w33262;
assign w25856 = (a_11 & ~w10506) | (a_11 & w33263) | (~w10506 & w33263);
assign w25857 = a_11 & ~w25615;
assign w25858 = ~w10073 & w26877;
assign w25859 = ~w10295 & w27268;
assign w25860 = w10254 & ~w10540;
assign w25861 = w10685 & w33264;
assign w25862 = w10718 & w33265;
assign w25863 = ~w10357 & w27269;
assign w25864 = (a_23 & ~w10736) | (a_23 & w33266) | (~w10736 & w33266);
assign w25865 = a_23 & ~w25616;
assign w25866 = ~w10375 & ~w10373;
assign w25867 = a_20 & ~w25617;
assign w25868 = w25433 & a_20;
assign w25869 = (a_17 & ~w10772) | (a_17 & w33267) | (~w10772 & w33267);
assign w25870 = a_17 & ~w25619;
assign w25871 = ~w10779 & w25110;
assign w25872 = ~w10779 & ~w10780;
assign w25873 = (a_14 & ~w10789) | (a_14 & w33268) | (~w10789 & w33268);
assign w25874 = a_14 & ~w25620;
assign w25875 = ~w10804 & ~w10803;
assign w25876 = w10845 & w33269;
assign w25877 = w10856 & w33270;
assign w25878 = w10871 & w33271;
assign w25879 = w11026 & w33272;
assign w25880 = (a_23 & ~w11066) | (a_23 & w33273) | (~w11066 & w33273);
assign w25881 = a_23 & ~w25621;
assign w25882 = a_20 & ~w25622;
assign w25883 = w25434 & a_20;
assign w25884 = (a_17 & ~w11101) | (a_17 & w33274) | (~w11101 & w33274);
assign w25885 = a_17 & ~w25624;
assign w25886 = a_14 & ~w25625;
assign w25887 = w25435 & a_14;
assign w25888 = w11227 & w33275;
assign w25889 = (a_14 & ~w11238) | (a_14 & w33276) | (~w11238 & w33276);
assign w25890 = a_14 & ~w25627;
assign w25891 = (a_17 & ~w11249) | (a_17 & w33277) | (~w11249 & w33277);
assign w25892 = a_17 & ~w25628;
assign w25893 = (a_29 & ~w11261) | (a_29 & w33278) | (~w11261 & w33278);
assign w25894 = a_29 & ~w25629;
assign w25895 = w11283 & w33279;
assign w25896 = w11412 & w33280;
assign w25897 = w11453 & w33281;
assign w25898 = (a_23 & ~w11469) | (a_23 & w33282) | (~w11469 & w33282);
assign w25899 = a_23 & ~w25630;
assign w25900 = (a_20 & ~w11487) | (a_20 & w33283) | (~w11487 & w33283);
assign w25901 = a_20 & ~w25631;
assign w25902 = w11564 & w33284;
assign w25903 = w11742 & w33285;
assign w25904 = (a_32 & ~w11760) | (a_32 & w33286) | (~w11760 & w33286);
assign w25905 = a_32 & ~w25632;
assign w25906 = (a_26 & ~w11793) | (a_26 & w33287) | (~w11793 & w33287);
assign w25907 = a_26 & ~w25633;
assign w25908 = a_23 & ~w25634;
assign w25909 = w25436 & a_23;
assign w25910 = w11829 & w33288;
assign w25911 = w11845 & w33289;
assign w25912 = w11924 & w33290;
assign w25913 = w12092 & w33291;
assign w25914 = w12110 & w33292;
assign w25915 = w12145 & w33293;
assign w25916 = (a_23 & ~w12163) | (a_23 & w33294) | (~w12163 & w33294);
assign w25917 = a_23 & ~w25636;
assign w25918 = ~w25129 & ~w12170;
assign w25919 = (a_20 & ~w12180) | (a_20 & w33295) | (~w12180 & w33295);
assign w25920 = a_20 & ~w25637;
assign w25921 = w12197 & w33296;
assign w25922 = a_17 & w25437;
assign w25923 = ~w12204 & ~w12206;
assign w25924 = ~w12204 & ~w11855;
assign w25925 = (a_17 & ~w12303) | (a_17 & w33297) | (~w12303 & w33297);
assign w25926 = a_17 & ~w25640;
assign w25927 = a_20 & ~w25641;
assign w25928 = w12316 & w33298;
assign w25929 = (a_23 & ~w12325) | (a_23 & w33299) | (~w12325 & w33299);
assign w25930 = a_23 & ~w25643;
assign w25931 = (a_32 & ~w12337) | (a_32 & w33300) | (~w12337 & w33300);
assign w25932 = a_32 & ~w25644;
assign w25933 = w12509 & w33301;
assign w25934 = w12533 & w33302;
assign w25935 = (a_26 & ~w12549) | (a_26 & w33303) | (~w12549 & w33303);
assign w25936 = a_26 & ~w25645;
assign w25937 = (a_17 & ~w12706) | (a_17 & w33304) | (~w12706 & w33304);
assign w25938 = a_17 & ~w25646;
assign w25939 = (a_20 & ~w12717) | (a_20 & w33305) | (~w12717 & w33305);
assign w25940 = a_20 & ~w25647;
assign w25941 = w12728 & w33306;
assign w25942 = w12901 & w33307;
assign w25943 = (a_29 & ~w12926) | (a_29 & w33308) | (~w12926 & w33308);
assign w25944 = a_29 & ~w25648;
assign w25945 = a_26 & ~w25649;
assign w25946 = w25451 & a_26;
assign w25947 = (a_20 & ~w13052) | (a_20 & w33309) | (~w13052 & w33309);
assign w25948 = a_20 & ~w25651;
assign w25949 = w12955 & ~w12951;
assign w25950 = w13279 & w33310;
assign w25951 = w13296 & w33311;
assign w25952 = w13780 & w33312;
assign w25953 = (a_17 & ~w14051) | (a_17 & w33313) | (~w14051 & w33313);
assign w25954 = a_17 & ~w25652;
assign w25955 = (a_14 & ~w14158) | (a_14 & w33314) | (~w14158 & w33314);
assign w25956 = (a_14 & ~w14159) | (a_14 & w25493) | (~w14159 & w25493);
assign w25957 = a_14 & ~w25955;
assign w25958 = w14159 & w33315;
assign w25959 = w14043 & ~w13788;
assign w25960 = ~w14173 & ~w14174;
assign w25961 = w14184 & w33316;
assign w25962 = (~w27488 & w33317) | (~w27488 & w33318) | (w33317 & w33318);
assign w25963 = w14199 & w33319;
assign w25964 = a_26 & w14429;
assign w25965 = a_26 & ~w25455;
assign w25966 = ~a_26 & ~w14429;
assign w25967 = ~a_26 & w25455;
assign w25968 = w14069 & ~w14080;
assign w25969 = w14454 & ~w14153;
assign w25970 = w14167 & ~w14451;
assign w25971 = (a_23 & ~w14906) | (a_23 & w33320) | (~w14906 & w33320);
assign w25972 = a_23 & ~w25456;
assign w25973 = w15186 & w33321;
assign w25974 = w15214 & w33322;
assign w25975 = (a_32 & ~w15230) | (a_32 & w33323) | (~w15230 & w33323);
assign w25976 = a_32 & ~w25653;
assign w25977 = w15418 & ~w15429;
assign w25978 = w15586 & w33324;
assign w25979 = w15899 & ~w15902;
assign w25980 = a_29 & w16111;
assign w25981 = a_29 & ~w25663;
assign w25982 = ~a_29 & ~w16111;
assign w25983 = ~a_29 & w25663;
assign w25984 = w16218 & w33325;
assign w25985 = a_26 & w16235;
assign w25986 = a_26 & ~w25668;
assign w25987 = ~a_26 & ~w16235;
assign w25988 = ~a_26 & w25668;
assign w25989 = (a_29 & ~w16245) | (a_29 & w33326) | (~w16245 & w33326);
assign w25990 = a_29 & ~w25669;
assign w25991 = ~w15903 & w16121;
assign w25992 = ~w15903 & ~w15904;
assign w25993 = a_23 & w16461;
assign w25994 = a_23 & ~w25670;
assign w25995 = ~a_23 & ~w16461;
assign w25996 = ~a_23 & w25670;
assign w25997 = w17362 & ~w17185;
assign w25998 = w17681 & w33327;
assign w25999 = (a_29 & ~w17769) | (a_29 & w33328) | (~w17769 & w33328);
assign w26000 = a_29 & ~w25675;
assign w26001 = w17782 & w33329;
assign w26002 = w18050 & w33330;
assign w26003 = w18863 & w33331;
assign w26004 = (a_44 & ~w20482) | (a_44 & w33332) | (~w20482 & w33332);
assign w26005 = a_44 & ~w25676;
assign w26006 = w20664 & w33333;
assign w26007 = (a_44 & ~w20680) | (a_44 & w33334) | (~w20680 & w33334);
assign w26008 = a_44 & ~w25677;
assign w26009 = w20696 & w33335;
assign w26010 = (a_47 & ~w21120) | (a_47 & w33336) | (~w21120 & w33336);
assign w26011 = a_47 & ~w25678;
assign w26012 = w21285 & w33337;
assign w26013 = (a_47 & ~w21301) | (a_47 & w33338) | (~w21301 & w33338);
assign w26014 = a_47 & ~w25679;
assign w26015 = w21318 & w33339;
assign w26016 = w21494 & w33340;
assign w26017 = w21511 & w33341;
assign w26018 = w21626 & w33342;
assign w26019 = a_50 & ~w25680;
assign w26020 = w25460 & a_50;
assign w26021 = w21708 & ~w21710;
assign w26022 = w21717 & w33343;
assign w26023 = (a_56 & ~w21800) | (a_56 & w33344) | (~w21800 & w33344);
assign w26024 = a_56 & ~w25682;
assign w26025 = a_53 & ~w25683;
assign w26026 = w25461 & a_53;
assign w26027 = w21867 & ~w21869;
assign w26028 = a_50 & ~w25685;
assign w26029 = w25462 & a_50;
assign w26030 = w21883 & ~w21885;
assign w26031 = (a_47 & ~w21892) | (a_47 & w33345) | (~w21892 & w33345);
assign w26032 = a_47 & ~w25687;
assign w26033 = (a_62 & ~w22020) | (a_62 & w33346) | (~w22020 & w33346);
assign w26034 = a_62 & ~w25688;
assign w26035 = w22243 & w33347;
assign w26036 = a_59 & ~w25689;
assign w26037 = w25463 & a_59;
assign w26038 = a_56 & ~w25691;
assign w26039 = w25464 & a_56;
assign w26040 = a_53 & ~w25693;
assign w26041 = w25465 & a_53;
assign w26042 = w22419 & w33348;
assign w26043 = (a_62 & ~w22512) | (a_62 & w33349) | (~w22512 & w33349);
assign w26044 = a_62 & ~w25695;
assign w26045 = (a_59 & ~w22539) | (a_59 & w33350) | (~w22539 & w33350);
assign w26046 = a_59 & ~w25696;
assign w26047 = a_56 & ~w25697;
assign w26048 = w25466 & a_56;
assign w26049 = w22395 & ~w22391;
assign w26050 = a_53 & ~w25699;
assign w26051 = w25467 & a_53;
assign w26052 = w22413 & ~w22409;
assign w26053 = (a_50 & ~w22592) | (a_50 & w33351) | (~w22592 & w33351);
assign w26054 = a_50 & ~w25701;
assign w26055 = w22606 & ~w22617;
assign w26056 = (a_56 & ~w22747) | (a_56 & w33352) | (~w22747 & w33352);
assign w26057 = a_56 & ~w25702;
assign w26058 = w22833 & w33353;
assign w26059 = a_59 & ~w25703;
assign w26060 = w25468 & a_59;
assign w26061 = (a_56 & ~w22888) | (a_56 & w33354) | (~w22888 & w33354);
assign w26062 = a_56 & ~w25705;
assign w26063 = ~w22897 & w22898;
assign w26064 = w22897 & ~w22898;
assign w26065 = w22905 & w33355;
assign w26066 = (a_59 & ~w23021) | (a_59 & w33356) | (~w23021 & w33356);
assign w26067 = a_59 & ~w25706;
assign w26068 = (a_56 & ~w23038) | (a_56 & w33357) | (~w23038 & w33357);
assign w26069 = a_56 & ~w25707;
assign w26070 = w23056 & w33358;
assign w26071 = ~w23614 & ~w23615;
assign w26072 = w24240 & w33360;
assign w26073 = (a_62 & ~w24445) | (a_62 & w33361) | (~w24445 & w33361);
assign w26074 = a_62 & ~w25471;
assign w26075 = (w25268 & w33362) | (w25268 & w33363) | (w33362 & w33363);
assign w26076 = (w25263 & w33364) | (w25263 & w33365) | (w33364 & w33365);
assign w26077 = (~w25292 & w33366) | (~w25292 & w33367) | (w33366 & w33367);
assign w26078 = (~w25292 & w33368) | (~w25292 & w33369) | (w33368 & w33369);
assign w26079 = (~w25292 & w33370) | (~w25292 & w33371) | (w33370 & w33371);
assign w26080 = w24935 & w25714;
assign w26081 = ~w10119 & ~w10117;
assign w26082 = ~w11819 & ~w11818;
assign w26083 = ~w23413 & ~w23411;
assign w26084 = w23411 & w23544;
assign w26085 = w24124 & w24222;
assign w26086 = (w24222 & w24125) | (w24222 & w26085) | (w24125 & w26085);
assign w26087 = ~w24738 & ~w24739;
assign w26088 = (~w24738 & ~w24679) | (~w24738 & w26087) | (~w24679 & w26087);
assign w26089 = ~w12571 & ~w12569;
assign w26090 = ~w15 & a_5;
assign w26091 = ~w15 & a_8;
assign w26092 = w242 & a_8;
assign w26093 = w657 & w33372;
assign w26094 = w986 & w33373;
assign w26095 = w1295 & w33374;
assign w26096 = w1694 & w33375;
assign w26097 = ~w15 & a_47;
assign w26098 = w6764 & a_47;
assign w26099 = w7613 & w33376;
assign w26100 = w8526 & w33377;
assign w26101 = ~w15 & a_56;
assign w26102 = w9537 & a_56;
assign w26103 = ~w25746 & a_5;
assign w26104 = w106 & w90;
assign w26105 = w108 & w161;
assign w26106 = w125 & w187;
assign w26107 = ~w125 & ~w187;
assign w26108 = ~w25753 & a_8;
assign w26109 = w246 & w230;
assign w26110 = ~w25754 & a_8;
assign w26111 = ~w248 & w335;
assign w26112 = w248 & ~w335;
assign w26113 = w412 & b_1;
assign w26114 = w412 & b_2;
assign w26115 = (a_11 & ~w640) | (a_11 & w26514) | (~w640 & w26514);
assign w26116 = ~w671 & ~w670;
assign w26117 = w969 & w33378;
assign w26118 = ~w993 & ~w977;
assign w26119 = ~w1095 & ~w1094;
assign w26120 = w1278 & w33379;
assign w26121 = ~w1302 & ~w1286;
assign w26122 = ~w1448 & ~w1447;
assign w26123 = w1677 & w33380;
assign w26124 = ~w1701 & ~w1685;
assign w26125 = ~w1860 & ~w1859;
assign w26126 = w2141 & w33381;
assign w26127 = ~w2165 & ~w2149;
assign w26128 = w2152 & b_3;
assign w26129 = (a_26 & ~w2837) | (a_26 & w33382) | (~w2837 & w33382);
assign w26130 = w2849 & ~w3022;
assign w26131 = ~w3041 & ~w3039;
assign w26132 = ~w25784 & ~w3413;
assign w26133 = w3189 & b_1;
assign w26134 = w3189 & b_2;
assign w26135 = (a_32 & ~w3786) | (a_32 & w26515) | (~w3786 & w26515);
assign w26136 = ~w3817 & ~w3816;
assign w26137 = w3797 & b_1;
assign w26138 = w3797 & b_2;
assign w26139 = (a_35 & ~w4482) | (a_35 & w26516) | (~w4482 & w26516);
assign w26140 = ~w4513 & ~w4512;
assign w26141 = w4493 & b_1;
assign w26142 = w4493 & b_2;
assign w26143 = (a_38 & ~w5179) | (a_38 & w26517) | (~w5179 & w26517);
assign w26144 = ~w5210 & ~w5209;
assign w26145 = w5190 & b_1;
assign w26146 = w5190 & b_2;
assign w26147 = (a_41 & ~w5945) | (a_41 & w26518) | (~w5945 & w26518);
assign w26148 = ~w5976 & ~w5975;
assign w26149 = w5956 & b_1;
assign w26150 = w5956 & b_2;
assign w26151 = (a_44 & ~w6744) | (a_44 & w26990) | (~w6744 & w26990);
assign w26152 = ~w25807 & a_47;
assign w26153 = w6768 & w6752;
assign w26154 = ~w6775 & ~w6774;
assign w26155 = ~w25808 & a_47;
assign w26156 = ~w6770 & w7349;
assign w26157 = w6770 & ~w7349;
assign w26158 = w6755 & b_3;
assign w26159 = (a_47 & ~w7958) | (a_47 & w33383) | (~w7958 & w33383);
assign w26160 = ~w7967 & w26991;
assign w26161 = (~w7966 & w7592) | (~w7966 & w26992) | (w7592 & w26992);
assign w26162 = w8310 & w7973;
assign w26163 = w8310 & ~w7928;
assign w26164 = w8509 & w33384;
assign w26165 = ~w8533 & ~w8517;
assign w26166 = w7607 & b_3;
assign w26167 = (a_50 & ~w8903) | (a_50 & w33385) | (~w8903 & w33385);
assign w26168 = w8916 & ~w9271;
assign w26169 = w9517 & w33386;
assign w26170 = ~w25824 & a_56;
assign w26171 = w9541 & w9525;
assign w26172 = ~w9541 & ~w9525;
assign w26173 = ~w25825 & a_56;
assign w26174 = w8520 & b_3;
assign w26175 = (a_53 & ~w9893) | (a_53 & w33387) | (~w9893 & w33387);
assign w26176 = ~w9543 & w10240;
assign w26177 = w9543 & ~w10240;
assign w26178 = w9528 & b_1;
assign w26179 = w9543 & w10240;
assign w26180 = w9528 & b_2;
assign w26181 = (a_56 & ~w10545) | (a_56 & w27270) | (~w10545 & w27270);
assign w26182 = w10565 & w27271;
assign w26183 = w10258 & w10582;
assign w26184 = ~w10258 & ~w10582;
assign w26185 = ~w10277 & ~w10275;
assign w26186 = ~w10605 & ~w10604;
assign w26187 = ~w10289 & ~w10287;
assign w26188 = ~w10640 & ~w10639;
assign w26189 = w10667 & w33388;
assign w26190 = (a_32 & ~w10685) | (a_32 & w33389) | (~w10685 & w33389);
assign w26191 = a_32 & ~w25861;
assign w26192 = w10702 & w33390;
assign w26193 = (a_26 & ~w10718) | (a_26 & w33391) | (~w10718 & w33391);
assign w26194 = a_26 & ~w25862;
assign w26195 = a_17 & ~w25869;
assign w26196 = w25619 & a_17;
assign w26197 = a_14 & ~w25873;
assign w26198 = w25620 & a_14;
assign w26199 = (a_11 & ~w10845) | (a_11 & w33392) | (~w10845 & w33392);
assign w26200 = a_11 & ~w25876;
assign w26201 = (a_26 & ~w10856) | (a_26 & w33393) | (~w10856 & w33393);
assign w26202 = a_26 & ~w25877;
assign w26203 = ~w10711 & ~w10709;
assign w26204 = (a_44 & ~w10871) | (a_44 & w33394) | (~w10871 & w33394);
assign w26205 = a_44 & ~w25878;
assign w26206 = w10881 & w33395;
assign w26207 = w10556 & b_0;
assign w26208 = ~w10928 & ~w10927;
assign w26209 = w11008 & w33396;
assign w26210 = ~w10675 & w27272;
assign w26211 = (a_32 & ~w11026) | (a_32 & w33397) | (~w11026 & w33397);
assign w26212 = a_32 & ~w25879;
assign w26213 = ~w11033 & ~w11034;
assign w26214 = ~w11033 & w25114;
assign w26215 = w11042 & w33398;
assign w26216 = ~w11091 & w25115;
assign w26217 = ~w11091 & ~w11092;
assign w26218 = a_17 & ~w25884;
assign w26219 = w25624 & a_17;
assign w26220 = w10830 & w27273;
assign w26221 = ~w10473 & ~w10472;
assign w26222 = (~w10472 & ~w10473) | (~w10472 & w33399) | (~w10473 & w33399);
assign w26223 = w25118 | w25117;
assign w26224 = (w25117 & w25118) | (w25117 & w10448) | (w25118 & w10448);
assign w26225 = ~w11140 & w26754;
assign w26226 = (a_11 & ~w11227) | (a_11 & w33400) | (~w11227 & w33400);
assign w26227 = a_11 & ~w25888;
assign w26228 = a_14 & ~w25889;
assign w26229 = w25627 & a_14;
assign w26230 = a_17 & ~w25891;
assign w26231 = w25628 & a_17;
assign w26232 = a_29 & ~w25893;
assign w26233 = w25629 & a_29;
assign w26234 = (a_44 & ~w11283) | (a_44 & w33401) | (~w11283 & w33401);
assign w26235 = a_44 & ~w25895;
assign w26236 = w11394 & w33402;
assign w26237 = (a_35 & ~w11412) | (a_35 & w33403) | (~w11412 & w33403);
assign w26238 = a_35 & ~w25896;
assign w26239 = w11430 & w33404;
assign w26240 = (a_26 & ~w11453) | (a_26 & w33405) | (~w11453 & w33405);
assign w26241 = a_26 & ~w25897;
assign w26242 = a_20 & ~w25900;
assign w26243 = w25631 & a_20;
assign w26244 = w11253 & w11499;
assign w26245 = w25122 & w11535;
assign w26246 = (w11535 & w25122) | (w11535 & ~w11181) | (w25122 & ~w11181);
assign w26247 = w11553 & w33406;
assign w26248 = (a_14 & ~w11564) | (a_14 & w33407) | (~w11564 & w33407);
assign w26249 = a_14 & ~w25902;
assign w26250 = w11724 & w33408;
assign w26251 = (a_35 & ~w11742) | (a_35 & w33409) | (~w11742 & w33409);
assign w26252 = a_35 & ~w25903;
assign w26253 = a_32 & ~w25904;
assign w26254 = w25632 & a_32;
assign w26255 = w11777 & w33410;
assign w26256 = a_26 & ~w25906;
assign w26257 = w25633 & a_26;
assign w26258 = (a_20 & ~w11829) | (a_20 & w33411) | (~w11829 & w33411);
assign w26259 = a_20 & ~w25910;
assign w26260 = ~w11837 & ~w11836;
assign w26261 = (a_17 & ~w11845) | (a_17 & w33412) | (~w11845 & w33412);
assign w26262 = a_17 & ~w25911;
assign w26263 = ~w11866 & ~w11865;
assign w26264 = ~w11860 & ~w11859;
assign w26265 = (a_14 & ~w11924) | (a_14 & w33413) | (~w11924 & w33413);
assign w26266 = a_14 & ~w25912;
assign w26267 = w12074 & w33414;
assign w26268 = (a_35 & ~w12092) | (a_35 & w33415) | (~w12092 & w33415);
assign w26269 = a_35 & ~w25913;
assign w26270 = (a_32 & ~w12110) | (a_32 & w33416) | (~w12110 & w33416);
assign w26271 = a_32 & ~w25914;
assign w26272 = ~w25128 & ~w12117;
assign w26273 = w12127 & w33417;
assign w26274 = ~w11786 & ~w11784;
assign w26275 = (a_26 & ~w12145) | (a_26 & w33418) | (~w12145 & w33418);
assign w26276 = a_26 & ~w25915;
assign w26277 = (w25125 & w27498) | (w25125 & w27499) | (w27498 & w27499);
assign w26278 = a_23 & ~w25916;
assign w26279 = w25636 & a_23;
assign w26280 = ~w12171 & w11931;
assign w26281 = a_20 & ~w25919;
assign w26282 = w25637 & a_20;
assign w26283 = (~w11853 & w11571) | (~w11853 & w27500) | (w11571 & w27500);
assign w26284 = (~w11930 & ~w26283) | (~w11930 & w27759) | (~w26283 & w27759);
assign w26285 = w12292 & w33419;
assign w26286 = a_17 & ~w25925;
assign w26287 = w25640 & a_17;
assign w26288 = w11840 & ~w12187;
assign w26289 = w12491 & w33420;
assign w26290 = (a_35 & ~w12509) | (a_35 & w33421) | (~w12509 & w33421);
assign w26291 = a_35 & ~w25933;
assign w26292 = a_26 & ~w25935;
assign w26293 = w25645 & a_26;
assign w26294 = w12592 & w33422;
assign w26295 = ~w12606 & w27501;
assign w26296 = (~w12628 & w12606) | (~w12628 & w27502) | (w12606 & w27502);
assign w26297 = w12603 & ~w12599;
assign w26298 = w12695 & w33423;
assign w26299 = a_17 & ~w25937;
assign w26300 = w25646 & a_17;
assign w26301 = a_20 & ~w25939;
assign w26302 = w25647 & a_20;
assign w26303 = w12883 & w33424;
assign w26304 = (a_35 & ~w12901) | (a_35 & w33425) | (~w12901 & w33425);
assign w26305 = a_35 & ~w25942;
assign w26306 = w12961 & w33426;
assign w26307 = w12713 & ~w12974;
assign w26308 = a_20 & ~w25947;
assign w26309 = w25651 & a_20;
assign w26310 = w13227 & w33427;
assign w26311 = w13262 & w33428;
assign w26312 = (a_26 & ~w13279) | (a_26 & w33429) | (~w13279 & w33429);
assign w26313 = a_26 & ~w25950;
assign w26314 = ~w13287 & ~w13286;
assign w26315 = (a_23 & ~w13296) | (a_23 & w33430) | (~w13296 & w33430);
assign w26316 = a_23 & ~w25951;
assign w26317 = (w13367 & w13354) | (w13367 & w33431) | (w13354 & w33431);
assign w26318 = ~w13354 & w33432;
assign w26319 = ~w12991 & w27817;
assign w26320 = w13436 & w33433;
assign w26321 = (w13364 & ~w13341) | (w13364 & w33434) | (~w13341 & w33434);
assign w26322 = w13743 & ~w13730;
assign w26323 = ~w13752 & w13753;
assign w26324 = w13752 & ~w13753;
assign w26325 = w13766 & w33435;
assign w26326 = (a_20 & ~w13780) | (a_20 & w33436) | (~w13780 & w33436);
assign w26327 = a_20 & ~w25952;
assign w26328 = w14029 & w33437;
assign w26329 = a_17 & ~w25953;
assign w26330 = w25652 & a_17;
assign w26331 = ~w14075 & ~w14076;
assign w26332 = w14082 & ~w14069;
assign w26333 = ~w14093 & ~w14094;
assign w26334 = w14087 & ~w14098;
assign w26335 = a_17 & w14174;
assign w26336 = a_17 & ~w25960;
assign w26337 = ~a_17 & ~w14174;
assign w26338 = ~a_17 & w25960;
assign w26339 = (a_20 & ~w14184) | (a_20 & w33438) | (~w14184 & w33438);
assign w26340 = a_20 & ~w25961;
assign w26341 = (a_23 & ~w14199) | (a_23 & w33439) | (~w14199 & w33439);
assign w26342 = a_23 & ~w25963;
assign w26343 = w14167 & w14451;
assign w26344 = ~w14167 & ~w14451;
assign w26345 = w14522 & w33440;
assign w26346 = w14423 & ~w14433;
assign w26347 = w14551 & w33441;
assign w26348 = w14165 & ~w14816;
assign w26349 = ~w14165 & w14816;
assign w26350 = w14892 & w33442;
assign w26351 = a_23 & ~w25971;
assign w26352 = w25456 & a_23;
assign w26353 = (a_17 & ~w15186) | (a_17 & w33443) | (~w15186 & w33443);
assign w26354 = a_17 & ~w25973;
assign w26355 = w15200 & w33444;
assign w26356 = (a_26 & ~w15214) | (a_26 & w33445) | (~w15214 & w33445);
assign w26357 = a_26 & ~w25974;
assign w26358 = a_32 & ~w25975;
assign w26359 = w25653 & a_32;
assign w26360 = w15234 & ~w15236;
assign w26361 = w14916 & ~w15144;
assign w26362 = ~w15449 & ~w15450;
assign w26363 = (a_29 & ~w15586) | (a_29 & w33446) | (~w15586 & w33446);
assign w26364 = a_29 & ~w25978;
assign w26365 = (a_20 & ~w16218) | (a_20 & w33447) | (~w16218 & w33447);
assign w26366 = a_20 & ~w25984;
assign w26367 = a_29 & ~w25989;
assign w26368 = w25669 & a_29;
assign w26369 = (w16249 & w16102) | (w16249 & w33450) | (w16102 & w33450);
assign w26370 = ~w16450 & ~w16449;
assign w26371 = w16454 & ~w16465;
assign w26372 = w16539 & w33451;
assign w26373 = w16842 & w33452;
assign w26374 = ~w17042 & ~w17043;
assign w26375 = w17152 & w33453;
assign w26376 = ~w17372 & ~w17373;
assign w26377 = (a_32 & ~w17681) | (a_32 & w33454) | (~w17681 & w33454);
assign w26378 = a_32 & ~w25998;
assign w26379 = w17677 & w33455;
assign w26380 = a_29 & ~w25999;
assign w26381 = w25675 & a_29;
assign w26382 = (a_32 & ~w17782) | (a_32 & w33456) | (~w17782 & w33456);
assign w26383 = a_32 & ~w26001;
assign w26384 = (w17690 & w33457) | (w17690 & w33458) | (w33457 & w33458);
assign w26385 = w18037 & w33459;
assign w26386 = (a_29 & ~w18050) | (a_29 & w33460) | (~w18050 & w33460);
assign w26387 = a_29 & ~w26002;
assign w26388 = w18065 & w33461;
assign w26389 = w18598 & w33462;
assign w26390 = (a_29 & ~w18863) | (a_29 & w33463) | (~w18863 & w33463);
assign w26391 = a_29 & ~w26003;
assign w26392 = w18878 & w33464;
assign w26393 = w19630 & w33465;
assign w26394 = w20015 & w33466;
assign w26395 = w20220 & w33467;
assign w26396 = w20238 & w33468;
assign w26397 = w20376 & w33469;
assign w26398 = a_44 & ~w26004;
assign w26399 = w25676 & a_44;
assign w26400 = (w20489 & w20227) | (w20489 & w33470) | (w20227 & w33470);
assign w26401 = w20498 & w33471;
assign w26402 = w20647 & w33472;
assign w26403 = (a_47 & ~w20664) | (a_47 & w33473) | (~w20664 & w33473);
assign w26404 = a_47 & ~w26006;
assign w26405 = a_44 & ~w26007;
assign w26406 = w25677 & a_44;
assign w26407 = w20688 & ~w20690;
assign w26408 = (a_41 & ~w20696) | (a_41 & w33474) | (~w20696 & w33474);
assign w26409 = a_41 & ~w26009;
assign w26410 = w21028 & w33475;
assign w26411 = a_47 & ~w26010;
assign w26412 = w25678 & a_47;
assign w26413 = w21136 & w33476;
assign w26414 = (~w26705 & w33477) | (~w26705 & w33478) | (w33477 & w33478);
assign w26415 = w21268 & w33479;
assign w26416 = (a_50 & ~w21285) | (a_50 & w33480) | (~w21285 & w33480);
assign w26417 = a_50 & ~w26012;
assign w26418 = a_47 & ~w26013;
assign w26419 = w25679 & a_47;
assign w26420 = ~w21309 & w21311;
assign w26421 = w21309 & ~w21311;
assign w26422 = (a_44 & ~w21318) | (a_44 & w33481) | (~w21318 & w33481);
assign w26423 = a_44 & ~w26015;
assign w26424 = w21417 & w33482;
assign w26425 = w21457 & w33483;
assign w26426 = (a_50 & ~w21494) | (a_50 & w33484) | (~w21494 & w33484);
assign w26427 = a_50 & ~w26016;
assign w26428 = (a_47 & ~w21511) | (a_47 & w33485) | (~w21511 & w33485);
assign w26429 = a_47 & ~w26017;
assign w26430 = w21528 & w33486;
assign w26431 = w21603 & w33487;
assign w26432 = w21614 & w33488;
assign w26433 = (a_53 & ~w21626) | (a_53 & w33489) | (~w21626 & w33489);
assign w26434 = a_53 & ~w26018;
assign w26435 = w21705 & w21697;
assign w26436 = (a_47 & ~w21717) | (a_47 & w33490) | (~w21717 & w33490);
assign w26437 = a_47 & ~w26022;
assign w26438 = (~w26021 & w33491) | (~w26021 & w33492) | (w33491 & w33492);
assign w26439 = a_56 & ~w26023;
assign w26440 = w25682 & a_56;
assign w26441 = w21835 & w33493;
assign w26442 = a_47 & ~w26031;
assign w26443 = w25687 & a_47;
assign w26444 = w21908 & w33494;
assign w26445 = (a_53 & ~w22243) | (a_53 & w33495) | (~w22243 & w33495);
assign w26446 = a_53 & ~w26035;
assign w26447 = (a_50 & ~w22419) | (a_50 & w33496) | (~w22419 & w33496);
assign w26448 = a_50 & ~w26042;
assign w26449 = w22601 & ~w22603;
assign w26450 = w22611 & w33497;
assign w26451 = ~w22605 & ~w22617;
assign w26452 = w22652 & ~w22641;
assign w26453 = w22730 & w33498;
assign w26454 = a_56 & ~w26056;
assign w26455 = w25702 & a_56;
assign w26456 = ~w22754 & w22756;
assign w26457 = w22754 & ~w22756;
assign w26458 = w22763 & w33499;
assign w26459 = (a_50 & ~w22833) | (a_50 & w33500) | (~w22833 & w33500);
assign w26460 = a_50 & ~w26058;
assign w26461 = w22877 & ~w22880;
assign w26462 = a_56 & ~w26061;
assign w26463 = w25705 & a_56;
assign w26464 = (a_53 & ~w22905) | (a_53 & w33501) | (~w22905 & w33501);
assign w26465 = a_53 & ~w26065;
assign w26466 = w22927 & w33502;
assign w26467 = w22953 & ~w22955;
assign w26468 = a_59 & ~w26066;
assign w26469 = w25706 & a_59;
assign w26470 = a_56 & ~w26068;
assign w26471 = w25707 & a_56;
assign w26472 = ~w22895 & w22898;
assign w26473 = ~w22895 & ~w22896;
assign w26474 = (a_53 & ~w23056) | (a_53 & w33503) | (~w23056 & w33503);
assign w26475 = a_53 & ~w26070;
assign w26476 = w26721 & w33504;
assign w26477 = w23321 & w33505;
assign w26478 = w23339 & w33506;
assign w26479 = a_62 & w23615;
assign w26480 = a_62 & ~w26071;
assign w26481 = ~a_62 & ~w23615;
assign w26482 = ~a_62 & w26071;
assign w26483 = w23838 & w33507;
assign w26484 = (~w25237 & w33508) | (~w25237 & w33509) | (w33508 & w33509);
assign w26485 = (~w25236 & w33508) | (~w25236 & w33509) | (w33508 & w33509);
assign w26486 = w23928 & w33510;
assign w26487 = ~w23950 & ~w23951;
assign w26488 = ~w23849 & w33511;
assign w26489 = ~w11623 & w24064;
assign w26490 = (a_62 & ~w24240) | (a_62 & w33512) | (~w24240 & w33512);
assign w26491 = a_62 & ~w26072;
assign w26492 = a_62 & ~w26073;
assign w26493 = w25471 & a_62;
assign w26494 = (~w9776 & w33513) | (~w9776 & w33514) | (w33513 & w33514);
assign w26495 = (~w25263 & w33515) | (~w25263 & w33516) | (w33515 & w33516);
assign w26496 = (~w25263 & w33519) | (~w25263 & w33520) | (w33519 & w33520);
assign w26497 = (~w25263 & w33523) | (~w25263 & w33524) | (w33523 & w33524);
assign w26498 = (~w25263 & w33527) | (~w25263 & w33528) | (w33527 & w33528);
assign w26499 = (~w25263 & w33531) | (~w25263 & w33532) | (w33531 & w33532);
assign w26500 = w24957 & w25472;
assign w26501 = (w25324 & w33535) | (w25324 & w33536) | (w33535 & w33536);
assign w26502 = ~w24972 & w25473;
assign w26503 = (w25324 & w33537) | (w25324 & w33538) | (w33537 & w33538);
assign w26504 = w24980 & w25474;
assign w26505 = (w25324 & w33539) | (w25324 & w33540) | (w33539 & w33540);
assign w26506 = ~w24980 & ~w25474;
assign w26507 = (~w25324 & w33541) | (~w25324 & w33542) | (w33541 & w33542);
assign w26508 = ~w10822 & ~w10820;
assign w26509 = w22319 & w22494;
assign w26510 = ~w23543 & ~w23544;
assign w26511 = (~w23543 & ~w23411) | (~w23543 & w26510) | (~w23411 & w26510);
assign w26512 = w24221 & w24315;
assign w26513 = ~w24791 & ~w24790;
assign w26514 = w418 & w33543;
assign w26515 = w3195 & w33544;
assign w26516 = w3803 & w33545;
assign w26517 = w4499 & w33546;
assign w26518 = w5196 & w33547;
assign w26519 = ~w186 & ~w187;
assign w26520 = (~w186 & ~w187) | (~w186 & w26878) | (~w187 & w26878);
assign w26521 = w93 & b_2;
assign w26522 = (a_5 & ~w222) | (a_5 & w26993) | (~w222 & w26993);
assign w26523 = w176 & ~w162;
assign w26524 = w233 & b_1;
assign w26525 = w233 & b_2;
assign w26526 = (a_8 & ~w401) | (a_8 & w26994) | (~w401 & w26994);
assign w26527 = ~w432 & ~w431;
assign w26528 = w640 & w33548;
assign w26529 = ~w664 & ~w648;
assign w26530 = ~w780 & ~w779;
assign w26531 = ~w26119 & ~w1094;
assign w26532 = w1098 & ~w1193;
assign w26533 = ~w26122 & ~w1447;
assign w26534 = w1451 & ~w1571;
assign w26535 = ~w26125 & ~w1859;
assign w26536 = w1863 & ~w2012;
assign w26537 = w2492 & w2659;
assign w26538 = ~w2492 & ~w2659;
assign w26539 = w2633 & b_3;
assign w26540 = (a_29 & ~w3405) | (a_29 & w33549) | (~w3405 & w33549);
assign w26541 = w3786 & w33550;
assign w26542 = ~w3810 & ~w3794;
assign w26543 = ~w3846 & ~w3845;
assign w26544 = ~w4053 & ~w4052;
assign w26545 = w4482 & w33551;
assign w26546 = ~w4506 & ~w4490;
assign w26547 = w3797 & b_3;
assign w26548 = (a_35 & ~w4740) | (a_35 & w33552) | (~w4740 & w33552);
assign w26549 = w5179 & w33553;
assign w26550 = ~w5203 & ~w5187;
assign w26551 = w4493 & b_3;
assign w26552 = (a_38 & ~w5476) | (a_38 & w33554) | (~w5476 & w33554);
assign w26553 = ~w5493 & w26995;
assign w26554 = w5945 & w33555;
assign w26555 = ~w5969 & ~w5953;
assign w26556 = w5190 & b_3;
assign w26557 = (a_41 & ~w6263) | (a_41 & w33556) | (~w6263 & w33556);
assign w26558 = ~w6280 & w26996;
assign w26559 = ~w7109 & w26997;
assign w26560 = w6755 & b_1;
assign w26561 = (w7124 & w7393) | (w7124 & w26998) | (w7393 & w26998);
assign w26562 = w7195 & w7475;
assign w26563 = ~w7195 & ~w7475;
assign w26564 = w7489 & w33557;
assign w26565 = (a_11 & ~w7505) | (a_11 & w33558) | (~w7505 & w33558);
assign w26566 = a_11 & ~w25065;
assign w26567 = w7260 & w7549;
assign w26568 = w7265 & w7553;
assign w26569 = ~w7457 & w27712;
assign w26570 = ~w7387 & ~w7386;
assign w26571 = w6755 & b_2;
assign w26572 = (a_47 & ~w7596) | (a_47 & w27374) | (~w7596 & w27374);
assign w26573 = ~w7400 & ~w7398;
assign w26574 = ~w7433 & w27274;
assign w26575 = ~w7452 & ~w7451;
assign w26576 = w7780 & w33559;
assign w26577 = (a_11 & ~w7798) | (a_11 & w33560) | (~w7798 & w33560);
assign w26578 = a_11 & ~w25067;
assign w26579 = ~w7531 & w33561;
assign w26580 = ~w7281 & ~w7280;
assign w26581 = ~w7770 & w27275;
assign w26582 = w25385 | w25386;
assign w26583 = (w25386 & w25385) | (w25386 & ~w7281) | (w25385 & ~w7281);
assign w26584 = (a_8 & ~w8196) | (a_8 & w33562) | (~w8196 & w33562);
assign w26585 = a_8 & ~w25389;
assign w26586 = (a_20 & ~w8207) | (a_20 & w33563) | (~w8207 & w33563);
assign w26587 = a_20 & ~w25390;
assign w26588 = ~w7990 & ~w7651;
assign w26589 = ~w7990 & ~w7991;
assign w26590 = ~w8092 & w26999;
assign w26591 = (w8309 & w8551) | (w8309 & w27000) | (w8551 & w27000);
assign w26592 = w8663 & w33564;
assign w26593 = w8681 & w33565;
assign w26594 = (a_17 & ~w8699) | (a_17 & w33566) | (~w8699 & w33566);
assign w26595 = a_17 & ~w25402;
assign w26596 = (a_11 & ~w8735) | (a_11 & w33567) | (~w8735 & w33567);
assign w26597 = a_11 & ~w25405;
assign w26598 = ~w25406 & ~w8742;
assign w26599 = (a_8 & ~w8751) | (a_8 & w33568) | (~w8751 & w33568);
assign w26600 = a_8 & ~w25407;
assign w26601 = w8810 & w33569;
assign w26602 = w8821 & w33570;
assign w26603 = ~w8545 & w27276;
assign w26604 = ~w8911 & ~w8912;
assign w26605 = (w8927 & w8913) | (w8927 & w33571) | (w8913 & w33571);
assign w26606 = ~w8913 & w33572;
assign w26607 = a_11 & ~w9054;
assign w26608 = a_11 & ~w25413;
assign w26609 = (a_8 & ~w9070) | (a_8 & w33573) | (~w9070 & w33573);
assign w26610 = a_8 & ~w25414;
assign w26611 = w9144 & a_11;
assign w26612 = w25415 & a_11;
assign w26613 = (a_23 & ~w9333) | (a_23 & w33574) | (~w9333 & w33574);
assign w26614 = a_23 & ~w25577;
assign w26615 = w9350 & w33575;
assign w26616 = w9408 & w33576;
assign w26617 = w9229 & ~w9278;
assign w26618 = w9634 & w33577;
assign w26619 = w9652 & w33578;
assign w26620 = w9670 & w33579;
assign w26621 = (a_20 & ~w9688) | (a_20 & w33580) | (~w9688 & w33580);
assign w26622 = a_20 & ~w25587;
assign w26623 = a_17 & ~w25589;
assign w26624 = w25421 & a_17;
assign w26625 = a_11 & ~w25593;
assign w26626 = w25424 & a_11;
assign w26627 = (a_23 & ~w9820) | (a_23 & w33581) | (~w9820 & w33581);
assign w26628 = a_23 & ~w25595;
assign w26629 = (a_26 & ~w9830) | (a_26 & w33582) | (~w9830 & w33582);
assign w26630 = a_26 & ~w25596;
assign w26631 = ~w9554 & ~w9553;
assign w26632 = ~w9901 & ~w9902;
assign w26633 = (w9917 & w9903) | (w9917 & w33583) | (w9903 & w33583);
assign w26634 = ~w9903 & w33584;
assign w26635 = a_17 & ~w25849;
assign w26636 = w25614 & a_17;
assign w26637 = w10420 & w10804;
assign w26638 = ~w10420 & ~w10804;
assign w26639 = ~w10809 & ~w10810;
assign w26640 = (~w10809 & ~w10810) | (~w10809 & w27713) | (~w10810 & w27713);
assign w26641 = w35 & w27277;
assign w26642 = ~w26208 & ~w10927;
assign w26643 = ~w11091 & ~w25115;
assign w26644 = ~w11091 & w11092;
assign w26645 = ~w10953 & ~w10952;
assign w26646 = a_20 & ~w26258;
assign w26647 = w25910 & a_20;
assign w26648 = (w27437 & w33585) | (w27437 & w33586) | (w33585 & w33586);
assign w26649 = a_17 & ~w26261;
assign w26650 = w25911 & a_17;
assign w26651 = w11507 & w11860;
assign w26652 = ~w11507 & ~w11860;
assign w26653 = w11514 & w11866;
assign w26654 = ~w11514 & ~w11866;
assign w26655 = ~w11523 & ~w11521;
assign w26656 = w11533 & w11912;
assign w26657 = w26283 & w27760;
assign w26658 = w12188 & ~w11840;
assign w26659 = ~w12999 & w27503;
assign w26660 = (~w13021 & w12999) | (~w13021 & w27504) | (w12999 & w27504);
assign w26661 = (w13327 & ~w13315) | (w13327 & w27761) | (~w13315 & w27761);
assign w26662 = w13315 & w27762;
assign w26663 = ~w12999 & w27818;
assign w26664 = ~w13395 & w13396;
assign w26665 = w13395 & ~w13396;
assign w26666 = w13463 & w33587;
assign w26667 = ~w13330 & ~w13329;
assign w26668 = w13417 & ~w13749;
assign w26669 = ~w13417 & ~w13749;
assign w26670 = ~w13392 & ~w13390;
assign w26671 = (a_23 & ~w14029) | (a_23 & w33588) | (~w14029 & w33588);
assign w26672 = a_23 & ~w26328;
assign w26673 = (w13726 & w13429) | (w13726 & w33589) | (w13429 & w33589);
assign w26674 = w14116 & ~w14105;
assign w26675 = a_23 & ~w26341;
assign w26676 = w25963 & a_23;
assign w26677 = w14203 & ~w14205;
assign w26678 = ~w14923 & ~w14924;
assign w26679 = a_26 & ~w26356;
assign w26680 = w25974 & a_26;
assign w26681 = ~w15222 & w33590;
assign w26682 = w15910 & w33591;
assign w26683 = ~w16259 & ~w16260;
assign w26684 = w16448 & ~w16253;
assign w26685 = w16568 & w33592;
assign w26686 = w16548 & ~w16785;
assign w26687 = a_32 & w17043;
assign w26688 = a_32 & ~w26374;
assign w26689 = ~a_32 & ~w17043;
assign w26690 = ~a_32 & w26374;
assign w26691 = w17662 & w33593;
assign w26692 = w18466 & w33594;
assign w26693 = w18484 & w33595;
assign w26694 = w19779 & w33596;
assign w26695 = w19982 & w33597;
assign w26696 = w19999 & w33598;
assign w26697 = (a_41 & ~w20015) | (a_41 & w33599) | (~w20015 & w33599);
assign w26698 = a_41 & ~w26394;
assign w26699 = w20110 & w33600;
assign w26700 = (a_44 & ~w20220) | (a_44 & w33601) | (~w20220 & w33601);
assign w26701 = a_44 & ~w26395;
assign w26702 = w20504 & ~w20493;
assign w26703 = w20837 & w33602;
assign w26704 = w20893 & w33603;
assign w26705 = (w21127 & w20900) | (w21127 & w33604) | (w20900 & w33604);
assign w26706 = w21206 & w33605;
assign w26707 = (a_53 & ~w21268) | (a_53 & w33606) | (~w21268 & w33606);
assign w26708 = a_53 & ~w26415;
assign w26709 = (a_53 & ~w21417) | (a_53 & w33607) | (~w21417 & w33607);
assign w26710 = a_53 & ~w26424;
assign w26711 = w21428 & w33608;
assign w26712 = a_50 & ~w26426;
assign w26713 = w26016 & a_50;
assign w26714 = w21537 & w21329;
assign w26715 = (w21713 & w33609) | (w21713 & w33610) | (w33609 & w33610);
assign w26716 = w22049 & w33611;
assign w26717 = ~w22601 & ~w22603;
assign w26718 = (w25216 & w33612) | (w25216 & w33613) | (w33612 & w33613);
assign w26719 = (~w25221 & w33614) | (~w25221 & w33615) | (w33614 & w33615);
assign w26720 = w23065 & ~w23067;
assign w26721 = ~w23065 & ~w23067;
assign w26722 = w23202 & w33616;
assign w26723 = (a_62 & ~w23321) | (a_62 & w33617) | (~w23321 & w33617);
assign w26724 = a_62 & ~w26477;
assign w26725 = (a_59 & ~w23339) | (a_59 & w33618) | (~w23339 & w33618);
assign w26726 = a_59 & ~w26478;
assign w26727 = ~w23609 & ~w23607;
assign w26728 = (w25236 & w33619) | (w25236 & w33620) | (w33619 & w33620);
assign w26729 = (w25236 & w33621) | (w25236 & w33622) | (w33621 & w33622);
assign w26730 = (w25236 & w33623) | (w25236 & w33624) | (w33623 & w33624);
assign w26731 = (w25236 & w33625) | (w25236 & w33626) | (w33625 & w33626);
assign w26732 = (w25236 & w33627) | (w25236 & w33628) | (w33627 & w33628);
assign w26733 = (w25236 & w33629) | (w25236 & w33630) | (w33629 & w33630);
assign w26734 = (w25236 & w33631) | (w25236 & w33632) | (w33631 & w33632);
assign w26735 = w25712 & w24874;
assign w26736 = ~w24872 & w26077;
assign w26737 = w25713 & w24908;
assign w26738 = ~w24906 & w26078;
assign w26739 = (w25263 & w33633) | (w25263 & w33634) | (w33633 & w33634);
assign w26740 = (w25268 & w33635) | (w25268 & w33636) | (w33635 & w33636);
assign w26741 = ~w10390 & ~w10389;
assign w26742 = w21180 & w21389;
assign w26743 = w21389 & ~w25485;
assign w26744 = ~w22492 & ~w22494;
assign w26745 = ~w22492 & ~w26509;
assign w26746 = w23676 & w23543;
assign w26747 = (w23676 & w23544) | (w23676 & w26746) | (w23544 & w26746);
assign w26748 = ~w23676 & ~w23674;
assign w26749 = ~w24314 & ~w24315;
assign w26750 = (~w24314 & ~w24221) | (~w24314 & w26749) | (~w24221 & w26749);
assign w26751 = ~w24832 & ~w24831;
assign w26752 = ~w9043 & ~w9042;
assign w26753 = ~w9714 & ~w9713;
assign w26754 = ~w11139 & ~w11138;
assign w26755 = w210 & ~w26519;
assign w26756 = w210 & ~w26520;
assign w26757 = ~w246 & ~w230;
assign w26758 = w196 & w261;
assign w26759 = w209 & w306;
assign w26760 = ~w292 & w27278;
assign w26761 = ~w425 & ~w409;
assign w26762 = w233 & b_3;
assign w26763 = (a_8 & ~w498) | (a_8 & w33637) | (~w498 & w33637);
assign w26764 = ~w26530 & ~w779;
assign w26765 = ~w799 & ~w798;
assign w26766 = w783 & ~w886;
assign w26767 = w651 & b_3;
assign w26768 = (a_14 & ~w1086) | (a_14 & w33638) | (~w1086 & w33638);
assign w26769 = w980 & b_3;
assign w26770 = (a_17 & ~w1439) | (a_17 & w33639) | (~w1439 & w33639);
assign w26771 = ~w1590 & ~w1588;
assign w26772 = w1289 & b_3;
assign w26773 = (a_20 & ~w1851) | (a_20 & w33640) | (~w1851 & w33640);
assign w26774 = ~w2031 & ~w2029;
assign w26775 = w2172 & ~w2291;
assign w26776 = ~w2343 & ~w2344;
assign w26777 = ~w2343 & ~w2198;
assign w26778 = ~w2871 & ~w2870;
assign w26779 = ~w2894 & w27123;
assign w26780 = w3417 & ~w3614;
assign w26781 = ~w3633 & ~w3631;
assign w26782 = ~w26543 & ~w3845;
assign w26783 = ~w26544 & ~w4052;
assign w26784 = w4056 & ~w4260;
assign w26785 = ~w5731 & ~w5730;
assign w26786 = ~w6521 & ~w6520;
assign w26787 = ~w6768 & ~w6752;
assign w26788 = w5956 & b_3;
assign w26789 = (a_44 & ~w7092) | (a_44 & w33641) | (~w7092 & w33641);
assign w26790 = ~w7393 & w27001;
assign w26791 = (~w7391 & w6801) | (~w7391 & w33642) | (w6801 & w33642);
assign w26792 = ~w7650 & ~w7649;
assign w26793 = (~w7927 & w7991) | (~w7927 & w27002) | (w7991 & w27002);
assign w26794 = ~w8310 & ~w7973;
assign w26795 = ~w8310 & w7928;
assign w26796 = ~w8316 & w27003;
assign w26797 = ~w8563 & ~w8562;
assign w26798 = ~w8567 & w8577;
assign w26799 = w8567 & ~w8577;
assign w26800 = (w8327 & w8591) | (w8327 & w27004) | (w8591 & w27004);
assign w26801 = ~w8344 & w27505;
assign w26802 = ~w8386 & ~w8384;
assign w26803 = w25406 & w8442;
assign w26804 = w25406 & ~w25079;
assign w26805 = w8471 & w8801;
assign w26806 = (w26802 & w27375) | (w26802 & w27376) | (w27375 & w27376);
assign w26807 = ~w8656 & ~w8654;
assign w26808 = ~w8638 & w27506;
assign w26809 = ~w8585 & w27005;
assign w26810 = ~w8580 & ~w8579;
assign w26811 = ~w25083 & ~w9060;
assign w26812 = ~w9095 & w25565;
assign w26813 = w25084 & w27006;
assign w26814 = w25566 | w25567;
assign w26815 = (w25567 & w25566) | (w25567 & ~w8183) | (w25566 & ~w8183);
assign w26816 = ~w9007 & w27507;
assign w26817 = ~w8936 & ~w8935;
assign w26818 = (w9299 & w9577) | (w9299 & w27279) | (w9577 & w27279);
assign w26819 = ~w9589 & ~w9196;
assign w26820 = ~w9374 & w27007;
assign w26821 = ~w9560 & ~w9559;
assign w26822 = w10165 & w10412;
assign w26823 = w9528 & b_3;
assign w26824 = (a_56 & ~w10919) | (a_56 & w33643) | (~w10919 & w33643);
assign w26825 = ~w10606 & w27280;
assign w26826 = ~w11346 & ~w10931;
assign w26827 = w11346 & w10931;
assign w26828 = a_14 & ~w26248;
assign w26829 = w25902 & a_14;
assign w26830 = ~w11380 & w27444;
assign w26831 = w11346 & ~w10931;
assign w26832 = w11340 & ~w11598;
assign w26833 = ~w11663 & ~w11662;
assign w26834 = (w11909 & w11890) | (w11909 & w33644) | (w11890 & w33644);
assign w26835 = ~w11890 & w33645;
assign w26836 = (~w25440 & w27714) | (~w25440 & w27715) | (w27714 & w27715);
assign w26837 = w12999 & w33646;
assign w26838 = (~w13389 & ~w12999) | (~w13389 & w33647) | (~w12999 & w33647);
assign w26839 = w13383 & w13392;
assign w26840 = (w12677 & w13024) | (w12677 & w27839) | (w13024 & w27839);
assign w26841 = (~w25196 & w33650) | (~w25196 & w33651) | (w33650 & w33651);
assign w26842 = (~w25196 & w33653) | (~w25196 & w33654) | (w33653 & w33654);
assign w26843 = (w25195 & w33655) | (w25195 & w33656) | (w33655 & w33656);
assign w26844 = (~w25196 & w33657) | (~w25196 & w33658) | (w33657 & w33658);
assign w26845 = (~w25221 & w33659) | (~w25221 & w33660) | (w33659 & w33660);
assign w26846 = (~w25221 & w33662) | (~w25221 & w33663) | (w33662 & w33663);
assign w26847 = (~w25221 & w33665) | (~w25221 & w33666) | (w33665 & w33666);
assign w26848 = (~w25221 & w33668) | (~w25221 & w33669) | (w33668 & w33669);
assign w26849 = (~w25221 & w33671) | (~w25221 & w33672) | (w33671 & w33672);
assign w26850 = (~w25221 & w33674) | (~w25221 & w33675) | (w33674 & w33675);
assign w26851 = (~w25221 & w33677) | (~w25221 & w33678) | (w33677 & w33678);
assign w26852 = (w25221 & w33680) | (w25221 & w33681) | (w33680 & w33681);
assign w26853 = (~w25216 & w33682) | (~w25216 & w33683) | (w33682 & w33683);
assign w26854 = (~w25268 & w33684) | (~w25268 & w33685) | (w33684 & w33685);
assign w26855 = ~w24619 & w26495;
assign w26856 = (~w25268 & w33686) | (~w25268 & w33687) | (w33686 & w33687);
assign w26857 = w24682 & w26496;
assign w26858 = (~w25268 & w33688) | (~w25268 & w33689) | (w33688 & w33689);
assign w26859 = ~w24739 & w26497;
assign w26860 = (~w25268 & w33690) | (~w25268 & w33691) | (w33690 & w33691);
assign w26861 = ~w24791 & w26498;
assign w26862 = (~w25268 & w33692) | (~w25268 & w33693) | (w33692 & w33693);
assign w26863 = ~w24832 & w26499;
assign w26864 = ~w2712 & ~w2710;
assign w26865 = (~w3489 & ~w3675) | (~w3489 & w27124) | (~w3675 & w27124);
assign w26866 = w20305 & w20535;
assign w26867 = ~w20535 & ~w20533;
assign w26868 = ~w21387 & ~w21389;
assign w26869 = ~w21387 & ~w26742;
assign w26870 = w21584 & ~w21581;
assign w26871 = ~w22662 & ~w22661;
assign w26872 = w23674 & w23798;
assign w26873 = (w23798 & w23676) | (w23798 & w26872) | (w23676 & w26872);
assign w26874 = ~w24400 & ~w24399;
assign w26875 = w7697 & w27281;
assign w26876 = ~w8708 & ~w8706;
assign w26877 = (~w26822 & w27008) | (~w26822 & w27009) | (w27008 & w27009);
assign w26878 = ~w125 & ~w186;
assign w26879 = (w306 & w26759) | (w306 & w26756) | (w26759 & w26756);
assign w26880 = (w306 & w26759) | (w306 & w26755) | (w26759 & w26755);
assign w26881 = ~w259 & ~w261;
assign w26882 = (~w259 & ~w261) | (~w259 & w27282) | (~w261 & w27282);
assign w26883 = w305 & w368;
assign w26884 = ~w515 & w27283;
assign w26885 = w412 & b_3;
assign w26886 = (a_11 & ~w771) | (a_11 & w33694) | (~w771 & w33694);
assign w26887 = w893 & w1012;
assign w26888 = ~w1212 & ~w1210;
assign w26889 = ~w3052 & w27125;
assign w26890 = ~w3249 & ~w3248;
assign w26891 = w3383 & ~w3466;
assign w26892 = (w26891 & w33695) | (w26891 & w33696) | (w33695 & w33696);
assign w26893 = w3884 & ~w3880;
assign w26894 = w3189 & b_3;
assign w26895 = (a_32 & ~w4044) | (a_32 & w33697) | (~w4044 & w33697);
assign w26896 = (w4092 & ~w4080) | (w4092 & w27284) | (~w4080 & w27284);
assign w26897 = w4080 & w27285;
assign w26898 = w3866 & ~w3862;
assign w26899 = w4024 & ~w4070;
assign w26900 = ~w3833 & w33698;
assign w26901 = ~w4768 & ~w4766;
assign w26902 = w4984 & ~w4980;
assign w26903 = ~w5999 & ~w5998;
assign w26904 = (w6293 & ~w6232) | (w6293 & w27286) | (~w6232 & w27286);
assign w26905 = w6232 & w27287;
assign w26906 = ~w6798 & ~w6797;
assign w26907 = (w7122 & ~w7061) | (w7122 & w27288) | (~w7061 & w27288);
assign w26908 = w7061 & w27289;
assign w26909 = ~w7668 & ~w7667;
assign w26910 = (w26909 & w27126) | (w26909 & w27127) | (w27126 & w27127);
assign w26911 = w8329 & w8002;
assign w26912 = w8329 & ~w7906;
assign w26913 = w8953 & ~w8964;
assign w26914 = w9218 & ~w9286;
assign w26915 = ~w9295 & ~w9293;
assign w26916 = ~w10586 & w10589;
assign w26917 = w10556 & b_1;
assign w26918 = w10556 & b_2;
assign w26919 = (a_59 & ~w11603) | (a_59 & w33699) | (~w11603 & w33699);
assign w26920 = w11623 & w27445;
assign w26921 = ~w11362 & ~w11360;
assign w26922 = ~w11698 & ~w11697;
assign w26923 = ~w11634 & ~w11633;
assign w26924 = w11614 & b_0;
assign w26925 = w35 & w27446;
assign w26926 = ~w11995 & ~w11994;
assign w26927 = w12051 & ~w11700;
assign w26928 = ~w12910 & ~w12909;
assign w26929 = (w25182 & w33700) | (w25182 & w33701) | (w33700 & w33701);
assign w26930 = (w25182 & w33702) | (w25182 & w33703) | (w33702 & w33703);
assign w26931 = (~w25182 & w33704) | (~w25182 & w33705) | (w33704 & w33705);
assign w26932 = (w25205 & w25204) | (w25205 & ~w25189) | (w25204 & ~w25189);
assign w26933 = ~w21182 & w26841;
assign w26934 = (w25195 & w33706) | (w25195 & w33707) | (w33706 & w33707);
assign w26935 = ~w21779 & w26842;
assign w26936 = (w25195 & w33708) | (w25195 & w33709) | (w33708 & w33709);
assign w26937 = (~w21960 & w25225) | (~w21960 & w26844) | (w25225 & w26844);
assign w26938 = (w25195 & w33710) | (w25195 & w33711) | (w33710 & w33711);
assign w26939 = (w25229 & w25228) | (w25229 & w26844) | (w25228 & w26844);
assign w26940 = (w25195 & w33712) | (w25195 & w33713) | (w33712 & w33713);
assign w26941 = (w25233 & w25232) | (w25233 & w26844) | (w25232 & w26844);
assign w26942 = (w25195 & w33714) | (w25195 & w33715) | (w33714 & w33715);
assign w26943 = (w25237 & w25236) | (w25237 & w26844) | (w25236 & w26844);
assign w26944 = (w25195 & w33716) | (w25195 & w33717) | (w33716 & w33717);
assign w26945 = (w25241 & w25240) | (w25241 & w26844) | (w25240 & w26844);
assign w26946 = (w25195 & w33718) | (w25195 & w33719) | (w33718 & w33719);
assign w26947 = (w26485 & w26484) | (w26485 & ~w26844) | (w26484 & ~w26844);
assign w26948 = (~w25195 & w33720) | (~w25195 & w33721) | (w33720 & w33721);
assign w26949 = (w25237 & w33722) | (w25237 & w33723) | (w33722 & w33723);
assign w26950 = ~w24022 & w26728;
assign w26951 = (w25237 & w33724) | (w25237 & w33725) | (w33724 & w33725);
assign w26952 = ~w24125 & w26729;
assign w26953 = (w25237 & w33726) | (w25237 & w33727) | (w33726 & w33727);
assign w26954 = ~w24222 & w26730;
assign w26955 = (w25237 & w33728) | (w25237 & w33729) | (w33728 & w33729);
assign w26956 = ~w24315 & w26731;
assign w26957 = (w25237 & w33730) | (w25237 & w33731) | (w33730 & w33731);
assign w26958 = ~w24400 & w26732;
assign w26959 = (w25237 & w33732) | (w25237 & w33733) | (w33732 & w33733);
assign w26960 = ~w24476 & w26733;
assign w26961 = (w25237 & w33734) | (w25237 & w33735) | (w33734 & w33735);
assign w26962 = ~w24549 & w26734;
assign w26963 = (w24529 & ~w24516) | (w24529 & w33736) | (~w24516 & w33736);
assign w26964 = w24592 & w33737;
assign w26965 = (w9770 & w33738) | (w9770 & w33739) | (w33738 & w33739);
assign w26966 = ~w7514 & ~w7512;
assign w26967 = ~w9300 & ~w9299;
assign w26968 = ~w18813 & ~w19077;
assign w26969 = ~w19582 & ~w19581;
assign w26970 = (~w19581 & ~w19337) | (~w19581 & w26969) | (~w19337 & w26969);
assign w26971 = ~w20533 & ~w26866;
assign w26972 = w20754 & w20533;
assign w26973 = (w20754 & w20535) | (w20754 & w26972) | (w20535 & w26972);
assign w26974 = w21581 & ~w21780;
assign w26975 = ~w21779 & w33740;
assign w26976 = w22825 & w22661;
assign w26977 = (w22825 & w22662) | (w22825 & w26976) | (w22662 & w26976);
assign w26978 = ~w23796 & ~w23798;
assign w26979 = ~w23796 & ~w26872;
assign w26980 = ~w23795 & w33741;
assign w26981 = w24476 & w24399;
assign w26982 = (w24476 & w24400) | (w24476 & w26981) | (w24400 & w26981);
assign w26983 = (~w24831 & w26751) | (~w24831 & ~w24790) | (w26751 & ~w24790);
assign w26984 = (~w24831 & w26751) | (~w24831 & w26513) | (w26751 & w26513);
assign w26985 = w7968 & w7626;
assign w26986 = ~w7968 & ~w7626;
assign w26987 = ~w8003 & ~w8002;
assign w26988 = ~w8948 & ~w8947;
assign w26989 = (~w10457 & w10436) | (~w10457 & w33742) | (w10436 & w33742);
assign w26990 = w5962 & w33743;
assign w26991 = ~w7968 & ~w7966;
assign w26992 = ~w7627 & ~w7966;
assign w26993 = w99 & w33744;
assign w26994 = w239 & w33745;
assign w26995 = ~w5492 & ~w5491;
assign w26996 = ~w6279 & ~w6278;
assign w26997 = ~w7108 & ~w7107;
assign w26998 = w7392 & w7124;
assign w26999 = ~w8093 & ~w8091;
assign w27000 = w8297 & w27377;
assign w27001 = ~w7392 & ~w7391;
assign w27002 = (~w7927 & w7651) | (~w7927 & w27290) | (w7651 & w27290);
assign w27003 = ~w8315 & ~w8314;
assign w27004 = w8326 & w27291;
assign w27005 = ~w8586 & ~w8584;
assign w27006 = ~w9096 & ~w9095;
assign w27007 = ~w9375 & ~w9373;
assign w27008 = ~w10071 & ~w10412;
assign w27009 = (~w10166 & ~w10060) | (~w10166 & w27819) | (~w10060 & w27819);
assign w27010 = ~a_0 & ~a_1;
assign w27011 = w93 & b_1;
assign w27012 = w222 & w33746;
assign w27013 = w93 & b_3;
assign w27014 = (a_5 & ~w283) | (a_5 & w33747) | (~w283 & w33747);
assign w27015 = w401 & w33748;
assign w27016 = ~w367 & ~w368;
assign w27017 = (~w367 & ~w368) | (~w367 & w27292) | (~w368 & w27292);
assign w27018 = ~w609 & ~w608;
assign w27019 = ~w1120 & ~w1119;
assign w27020 = ~w1473 & ~w1472;
assign w27021 = ~w1885 & ~w1884;
assign w27022 = (w2728 & w2900) | (w2728 & w33749) | (w2900 & w33749);
assign w27023 = ~w3273 & w27293;
assign w27024 = w3902 & ~w3898;
assign w27025 = ~w25035 & ~w4117;
assign w27026 = w3849 & ~w4094;
assign w27027 = ~w4295 & ~w4294;
assign w27028 = ~w4279 & ~w4277;
assign w27029 = (w27026 & w33750) | (w27026 & w33751) | (w33750 & w33751);
assign w27030 = ~w4319 & ~w4317;
assign w27031 = ~w5233 & ~w5232;
assign w27032 = (w5506 & ~w5445) | (w5506 & w27294) | (~w5445 & w27294);
assign w27033 = w5445 & w27295;
assign w27034 = w6744 & w33752;
assign w27035 = ~w6816 & ~w6815;
assign w27036 = (w7988 & ~w7928) | (w7988 & w27296) | (~w7928 & w27296);
assign w27037 = w7928 & w27297;
assign w27038 = w8294 & ~w8290;
assign w27039 = ~w8562 & w26591;
assign w27040 = ~w8562 & w8563;
assign w27041 = ~w8562 & ~w26591;
assign w27042 = ~w8602 & w26800;
assign w27043 = ~w8602 & ~w8603;
assign w27044 = (~w8964 & w8951) | (~w8964 & w27378) | (w8951 & w27378);
assign w27045 = ~w8625 & ~w8975;
assign w27046 = (w8987 & ~w27045) | (w8987 & w27508) | (~w27045 & w27508);
assign w27047 = w27045 & w27509;
assign w27048 = ~w8604 & w27298;
assign w27049 = w9095 & w9435;
assign w27050 = w9418 & ~w9415;
assign w27051 = w9588 & ~w9468;
assign w27052 = ~w9589 & ~w9588;
assign w27053 = ~w9308 & ~w9306;
assign w27054 = ~w9320 & ~w9318;
assign w27055 = ~w9326 & ~w9324;
assign w27056 = ~w25092 & ~w9731;
assign w27057 = ~w9566 & ~w9565;
assign w27058 = w9840 & w27299;
assign w27059 = ~w9988 & ~w25830;
assign w27060 = ~w25099 & ~w9988;
assign w27061 = ~w9678 & w27300;
assign w27062 = ~w9782 & ~w9784;
assign w27063 = (~w9782 & ~w9784) | (~w9782 & w27301) | (~w9784 & w27301);
assign w27064 = ~w9939 & w27302;
assign w27065 = w10289 & w9930;
assign w27066 = w10289 & ~w9851;
assign w27067 = ~w10289 & ~w9930;
assign w27068 = ~w10289 & w9851;
assign w27069 = ~w10036 & w27716;
assign w27070 = w11683 & ~w11679;
assign w27071 = w11648 & ~w11644;
assign w27072 = ~w12049 & w11700;
assign w27073 = ~w12049 & ~w12050;
assign w27074 = w12384 & ~w12396;
assign w27075 = (~w25171 & w33753) | (~w25171 & w33754) | (w33753 & w33754);
assign w27076 = (w25172 & w33755) | (w25172 & w33753) | (w33755 & w33753);
assign w27077 = (w25189 & w33756) | (w25189 & w33757) | (w33756 & w33757);
assign w27078 = ~w20073 & w26929;
assign w27079 = (w25189 & w33758) | (w25189 & w33759) | (w33758 & w33759);
assign w27080 = ~w20307 & w26930;
assign w27081 = (w25189 & w33760) | (w25189 & w33761) | (w33760 & w33761);
assign w27082 = (w25182 & w33762) | (w25182 & w33763) | (w33762 & w33763);
assign w27083 = (w25189 & w33764) | (w25189 & w33765) | (w33764 & w33765);
assign w27084 = (w25182 & w33766) | (w25182 & w33767) | (w33766 & w33767);
assign w27085 = (w25189 & w33768) | (w25189 & w33769) | (w33768 & w33769);
assign w27086 = (w25182 & w33770) | (w25182 & w33771) | (w33770 & w33771);
assign w27087 = (w25189 & w33772) | (w25189 & w33773) | (w33772 & w33773);
assign w27088 = (w25182 & w33774) | (w25182 & w33775) | (w33774 & w33775);
assign w27089 = (w25216 & w33776) | (w25216 & w33777) | (w33776 & w33777);
assign w27090 = ~w23127 & w26845;
assign w27091 = (w25216 & w33778) | (w25216 & w33779) | (w33778 & w33779);
assign w27092 = ~w23272 & w26846;
assign w27093 = (w25216 & w33780) | (w25216 & w33781) | (w33780 & w33781);
assign w27094 = ~w23413 & w26847;
assign w27095 = (w25216 & w33782) | (w25216 & w33783) | (w33782 & w33783);
assign w27096 = ~w23544 & w26848;
assign w27097 = (w25216 & w33784) | (w25216 & w33785) | (w33784 & w33785);
assign w27098 = ~w23676 & w26849;
assign w27099 = (w25216 & w33786) | (w25216 & w33787) | (w33786 & w33787);
assign w27100 = ~w23798 & w26850;
assign w27101 = (w25216 & w33788) | (w25216 & w33789) | (w33788 & w33789);
assign w27102 = ~w23910 & w26851;
assign w27103 = (~w25216 & w33790) | (~w25216 & w33791) | (w33790 & w33791);
assign w27104 = (w25221 & w33792) | (w25221 & w33793) | (w33792 & w33793);
assign w27105 = (~w25216 & w33794) | (~w25216 & w33795) | (w33794 & w33795);
assign w27106 = (w25221 & w33796) | (w25221 & w33797) | (w33796 & w33797);
assign w27107 = (~w25216 & w33798) | (~w25216 & w33799) | (w33798 & w33799);
assign w27108 = (w25221 & w33800) | (w25221 & w33801) | (w33800 & w33801);
assign w27109 = (~w25216 & w33802) | (~w25216 & w33803) | (w33802 & w33803);
assign w27110 = (w25221 & w33804) | (w25221 & w33805) | (w33804 & w33805);
assign w27111 = (~w25216 & w33806) | (~w25216 & w33807) | (w33806 & w33807);
assign w27112 = (w25221 & w33808) | (w25221 & w33809) | (w33808 & w33809);
assign w27113 = (~w25216 & w33810) | (~w25216 & w33811) | (w33810 & w33811);
assign w27114 = (w25221 & w33812) | (w25221 & w33813) | (w33812 & w33813);
assign w27115 = (~w25216 & w33814) | (~w25216 & w33815) | (w33814 & w33815);
assign w27116 = (w25221 & w33816) | (w25221 & w33817) | (w33816 & w33817);
assign w27117 = (~w25216 & w33818) | (~w25216 & w33819) | (w33818 & w33819);
assign w27118 = (w25221 & w33820) | (w25221 & w33821) | (w33820 & w33821);
assign w27119 = (~w25216 & w33822) | (~w25216 & w33823) | (w33822 & w33823);
assign w27120 = (w25221 & w33824) | (w25221 & w33825) | (w33824 & w33825);
assign w27121 = ~w8973 & ~w8972;
assign w27122 = ~w9643 & ~w9641;
assign w27123 = ~w2895 & ~w2893;
assign w27124 = (w3685 & ~w3478) | (w3685 & w33826) | (~w3478 & w33826);
assign w27125 = ~w3053 & ~w3051;
assign w27126 = ~w7995 & ~w7667;
assign w27127 = ~w7995 & w7579;
assign w27128 = w451 & ~w27016;
assign w27129 = w451 & ~w27017;
assign w27130 = (w26779 & w33827) | (w26779 & w33828) | (w33827 & w33828);
assign w27131 = ~w4352 & ~w4351;
assign w27132 = w4121 & ~w4333;
assign w27133 = ~w4531 & ~w4530;
assign w27134 = ~w4525 & ~w4524;
assign w27135 = (w4787 & ~w4775) | (w4787 & w27303) | (~w4775 & w27303);
assign w27136 = w4775 & w27304;
assign w27137 = ~w4795 & w27379;
assign w27138 = w4709 & ~w4772;
assign w27139 = ~w5039 & w27305;
assign w27140 = w5667 & ~w5753;
assign w27141 = ~w6017 & ~w6016;
assign w27142 = w6457 & ~w6543;
assign w27143 = ~w7139 & w33829;
assign w27144 = ~w7138 & w27306;
assign w27145 = (w7549 & w26567) | (w7549 & w7261) | (w26567 & w7261);
assign w27146 = (w7549 & w26567) | (w7549 & w25059) | (w26567 & w25059);
assign w27147 = ~w7620 & ~w7604;
assign w27148 = ~w7737 & w33830;
assign w27149 = ~w7481 & w27307;
assign w27150 = (w7530 & w7824) | (w7530 & w33831) | (w7824 & w33831);
assign w27151 = (~w26579 & w7824) | (~w26579 & w33832) | (w7824 & w33832);
assign w27152 = w7754 & ~w7751;
assign w27153 = ~w7736 & w27308;
assign w27154 = ~w7691 & w27717;
assign w27155 = ~w8038 & w25377;
assign w27156 = ~w8038 & ~w8039;
assign w27157 = ~w7788 & w27309;
assign w27158 = (w25388 & w25387) | (w25388 & ~w7553) | (w25387 & ~w7553);
assign w27159 = (w25388 & w25387) | (w25388 & ~w26568) | (w25387 & ~w26568);
assign w27160 = w8024 & ~w8020;
assign w27161 = ~w8110 & w27310;
assign w27162 = ~w8368 & w27311;
assign w27163 = ~w8407 & ~w8409;
assign w27164 = (~w8407 & ~w8409) | (~w8407 & w27312) | (~w8409 & w27312);
assign w27165 = (w8967 & w8604) | (w8967 & w27380) | (w8604 & w27380);
assign w27166 = w9002 & w8670;
assign w27167 = w9002 & ~w8673;
assign w27168 = ~w9002 & ~w8670;
assign w27169 = ~w9002 & w8673;
assign w27170 = w9308 & w8965;
assign w27171 = w9308 & ~w27048;
assign w27172 = ~w9308 & ~w8965;
assign w27173 = ~w9308 & w27048;
assign w27174 = ~w9341 & w27313;
assign w27175 = ~w10006 & w9837;
assign w27176 = w9592 & ~w9955;
assign w27177 = ~w9972 & ~w9974;
assign w27178 = ~w9972 & ~w9611;
assign w27179 = w10513 & ~w10797;
assign w27180 = (w27179 & w27510) | (w27179 & w27511) | (w27510 & w27511);
assign w27181 = w10643 & ~w10982;
assign w27182 = (w27180 & w27314) | (w27180 & w27315) | (w27314 & w27315);
assign w27183 = ~w11374 & ~w11372;
assign w27184 = ~w11681 & w11683;
assign w27185 = w11681 & ~w11683;
assign w27186 = w26922 & w27447;
assign w27187 = ~w11640 & ~w11639;
assign w27188 = ~w26926 & ~w11994;
assign w27189 = ~w12051 & ~w11700;
assign w27190 = w12051 & w11700;
assign w27191 = w11614 & b_1;
assign w27192 = w11998 & ~w12412;
assign w27193 = ~w12460 & ~w12459;
assign w27194 = ~w12466 & ~w12464;
assign w27195 = w12484 & ~w12480;
assign w27196 = ~w13235 & ~w13234;
assign w27197 = ~w10019 & ~w10017;
assign w27198 = (~w450 & w27016) | (~w450 & w27381) | (w27016 & w27381);
assign w27199 = (~w450 & w27017) | (~w450 & w27381) | (w27017 & w27381);
assign w27200 = ~w527 & ~w526;
assign w27201 = w538 & ~w618;
assign w27202 = ~w694 & ~w693;
assign w27203 = ~w1349 & ~w1348;
assign w27204 = w1481 & ~w1477;
assign w27205 = ~w2911 & ~w2912;
assign w27206 = ~w2911 & w27022;
assign w27207 = w27316 | w27317;
assign w27208 = w27318 & w27319;
assign w27209 = ~w4590 & ~w4589;
assign w27210 = (w4571 & w4819) | (w4571 & w27320) | (w4819 & w27320);
assign w27211 = ~w5024 & ~w5022;
assign w27212 = w5277 & ~w5273;
assign w27213 = (w5291 & w5532) | (w5291 & w27321) | (w5532 & w27321);
assign w27214 = ~w5521 & ~w5520;
assign w27215 = ~w5515 & ~w5514;
assign w27216 = ~w5755 & ~w5667;
assign w27217 = w5755 & w5667;
assign w27218 = w5529 & ~w5525;
assign w27219 = ~w5782 & w33833;
assign w27220 = w6021 & w6308;
assign w27221 = ~w6021 & ~w6308;
assign w27222 = ~w5773 & w33834;
assign w27223 = ~w6302 & ~w6301;
assign w27224 = ~w6545 & ~w6457;
assign w27225 = w6545 & w6457;
assign w27226 = (w25051 & w33835) | (w25051 & w33836) | (w33835 & w33836);
assign w27227 = ~w25055 & ~w7171;
assign w27228 = w7157 & ~w7153;
assign w27229 = (w26575 & w27382) | (w26575 & w27383) | (w27382 & w27383);
assign w27230 = w26797 & w8563;
assign w27231 = w26797 & ~w26591;
assign w27232 = ~w8970 & ~w8850;
assign w27233 = (w25410 & w27512) | (w25410 & w27513) | (w27512 & w27513);
assign w27234 = w9609 & ~w9605;
assign w27235 = (~w9987 & ~w9839) | (~w9987 & w27514) | (~w9839 & w27514);
assign w27236 = w9839 & w27515;
assign w27237 = ~w9989 & ~w9629;
assign w27238 = ~w10342 & ~w10340;
assign w27239 = ~w10336 & ~w10335;
assign w27240 = ~w10302 & ~w10300;
assign w27241 = ~w10779 & ~w25872;
assign w27242 = (~w10779 & w10168) | (~w10779 & w27718) | (w10168 & w27718);
assign w27243 = w10660 & ~w10656;
assign w27244 = ~w10726 & w27322;
assign w27245 = (w25866 & w27323) | (w25866 & w27324) | (w27323 & w27324);
assign w27246 = ~w11016 & w27764;
assign w27247 = ~w11387 & ~w11385;
assign w27248 = (w11268 & w27448) | (w11268 & w27449) | (w27448 & w27449);
assign w27249 = (w25127 & w27719) | (w25127 & w27720) | (w27719 & w27720);
assign w27250 = w11614 & b_2;
assign w27251 = (a_62 & ~w12772) | (a_62 & w33837) | (~w12772 & w33837);
assign w27252 = ~w13110 & ~w13109;
assign w27253 = ~w12891 & w27450;
assign w27254 = ~w27196 & ~w13234;
assign w27255 = w12937 & ~w12933;
assign w27256 = ~w13383 & w13392;
assign w27257 = ~w2350 & ~w2348;
assign w27258 = ~w6858 & ~w6856;
assign w27259 = ~w6822 & ~w6820;
assign w27260 = ~w11421 & ~w11419;
assign w27261 = ~w9622 & ~w9987;
assign w27262 = ~w10691 & ~w11032;
assign w27263 = ~w8392 & ~w8390;
assign w27264 = ~w8942 & ~w8940;
assign w27265 = ~w10097 & w33838;
assign w27266 = (~w10110 & w10097) | (~w10110 & w33839) | (w10097 & w33839);
assign w27267 = ~w9932 & ~w9930;
assign w27268 = ~w10294 & ~w10293;
assign w27269 = ~w10358 & ~w10356;
assign w27270 = w9534 & w33840;
assign w27271 = ~w15 & a_59;
assign w27272 = ~w10676 & ~w10674;
assign w27273 = (~w11155 & w11140) | (~w11155 & w33841) | (w11140 & w33841);
assign w27274 = ~w7434 & ~w7432;
assign w27275 = ~w7771 & ~w7769;
assign w27276 = ~w8546 & ~w8544;
assign w27277 = w10565 & a_59;
assign w27278 = ~w293 & ~w291;
assign w27279 = w9298 & w33842;
assign w27280 = ~w10604 & ~w10957;
assign w27281 = ~w7707 & ~w8037;
assign w27282 = ~w196 & ~w259;
assign w27283 = ~w514 & ~w513;
assign w27284 = ~w3833 & w33843;
assign w27285 = (~w4092 & w3833) | (~w4092 & w33844) | (w3833 & w33844);
assign w27286 = ~w6280 & w33845;
assign w27287 = (~w6293 & w6280) | (~w6293 & w33846) | (w6280 & w33846);
assign w27288 = ~w7109 & w33847;
assign w27289 = (~w7122 & w7109) | (~w7122 & w33848) | (w7109 & w33848);
assign w27290 = w7638 & w33849;
assign w27291 = ~w8236 & ~w8601;
assign w27292 = ~w305 & ~w367;
assign w27293 = ~w3274 & ~w3272;
assign w27294 = ~w5493 & w33850;
assign w27295 = (~w5506 & w5493) | (~w5506 & w33851) | (w5493 & w33851);
assign w27296 = ~w7975 & w33852;
assign w27297 = (~w7988 & w7975) | (~w7988 & w33853) | (w7975 & w33853);
assign w27298 = ~w8602 & ~w8965;
assign w27299 = (~w9954 & w9939) | (~w9954 & w27384) | (w9939 & w27384);
assign w27300 = ~w9679 & ~w9677;
assign w27301 = ~w9439 & ~w9782;
assign w27302 = ~w9938 & ~w9937;
assign w27303 = w4709 & w4787;
assign w27304 = ~w4709 & ~w4787;
assign w27305 = ~w5040 & ~w5038;
assign w27306 = ~w7137 & ~w7136;
assign w27307 = ~w7480 & ~w7479;
assign w27308 = ~w7735 & ~w7734;
assign w27309 = ~w7789 & ~w7787;
assign w27310 = ~w8111 & ~w8109;
assign w27311 = ~w8369 & ~w8367;
assign w27312 = (~w8073 & w8396) | (~w8073 & w27820) | (w8396 & w27820);
assign w27313 = ~w9342 & ~w9340;
assign w27314 = (~w11125 & ~w11506) | (~w11125 & w33854) | (~w11506 & w33854);
assign w27315 = ~w11507 & ~w11127;
assign w27316 = w3503 & ~w25017;
assign w27317 = w3503 & ~w3372;
assign w27318 = ~w3503 & w25017;
assign w27319 = ~w3503 & w3372;
assign w27320 = w4560 & w27385;
assign w27321 = w5280 & w27386;
assign w27322 = ~w10727 & ~w10725;
assign w27323 = ~w10743 & ~w10373;
assign w27324 = ~w10743 & w10169;
assign w27325 = w27010 & b_1;
assign w27326 = (a_2 & ~w48) | (a_2 & w33855) | (~w48 & w33855);
assign w27327 = w318 & ~w314;
assign w27328 = w519 & w535;
assign w27329 = ~w519 & ~w535;
assign w27330 = (~w526 & w27200) | (~w526 & w27199) | (w27200 & w27199);
assign w27331 = ~w1018 & ~w1017;
assign w27332 = ~w1602 & ~w1600;
assign w27333 = ~w1748 & ~w1747;
assign w27334 = w1798 & ~w1897;
assign w27335 = w1893 & ~w1889;
assign w27336 = ~w4142 & ~w4141;
assign w27337 = (w27336 & w33856) | (w27336 & w33857) | (w33856 & w33857);
assign w27338 = ~w27209 & ~w4589;
assign w27339 = ~w4830 & w27210;
assign w27340 = ~w4830 & ~w4831;
assign w27341 = ~w5543 & w27213;
assign w27342 = ~w5543 & ~w5544;
assign w27343 = ~w6331 & ~w6330;
assign w27344 = (w27144 & w33858) | (w27144 & w33859) | (w33858 & w33859);
assign w27345 = ~w27002 & w33860;
assign w27346 = ~w8363 & ~w8362;
assign w27347 = w9287 & ~w9218;
assign w27348 = w9218 & ~w9287;
assign w27349 = ~w9588 & w25089;
assign w27350 = ~w9588 & ~w26818;
assign w27351 = ~w9607 & w9609;
assign w27352 = w9607 & ~w9609;
assign w27353 = w9574 & ~w9570;
assign w27354 = w10545 & w33861;
assign w27355 = ~w26182 & a_59;
assign w27356 = w10569 & w10553;
assign w27357 = ~w10569 & ~w10553;
assign w27358 = ~w10623 & w10625;
assign w27359 = w10623 & ~w10625;
assign w27360 = ~w26641 & a_59;
assign w27361 = ~w10984 & ~w10643;
assign w27362 = w10984 & w10643;
assign w27363 = (w25121 & w27516) | (w25121 & w27517) | (w27516 & w27517);
assign w27364 = ~w11837 & ~w26260;
assign w27365 = ~w12020 & ~w12019;
assign w27366 = w12367 & ~w12417;
assign w27367 = w12366 & ~w12435;
assign w27368 = ~w12498 & w12502;
assign w27369 = ~w12830 & w33862;
assign w27370 = ~w12782 & w33863;
assign w27371 = ~w27252 & ~w13109;
assign w27372 = ~w13235 & w13060;
assign w27373 = ~w3292 & ~w3290;
assign w27374 = w6761 & w33864;
assign w27375 = ~w8670 & ~w8384;
assign w27376 = ~w8670 & w8214;
assign w27377 = ~w8307 & ~w8561;
assign w27378 = w8851 & ~w8964;
assign w27379 = ~w4796 & ~w4794;
assign w27380 = w8602 & w8967;
assign w27381 = ~w451 & ~w450;
assign w27382 = (~w7451 & ~w7715) | (~w7451 & w33865) | (~w7715 & w33865);
assign w27383 = ~w7726 & w7175;
assign w27384 = ~w9936 & w33866;
assign w27385 = ~w4570 & ~w4829;
assign w27386 = ~w5290 & ~w5542;
assign w27387 = w8 & w33867;
assign w27388 = a_0 & b_1;
assign w27389 = w27010 & b_0;
assign w27390 = a_0 & b_3;
assign w27391 = w76 & w33868;
assign w27392 = ~w106 & ~w90;
assign w27393 = ~w42 & ~w67;
assign w27394 = w115 & ~w111;
assign w27395 = ~w462 & ~w461;
assign w27396 = (~w27198 & w27451) | (~w27198 & w27452) | (w27451 & w27452);
assign w27397 = (~w27199 & w27451) | (~w27199 & w27452) | (w27451 & w27452);
assign w27398 = w519 & ~w535;
assign w27399 = w719 & ~w723;
assign w27400 = ~w893 & ~w1012;
assign w27401 = ~w1126 & ~w1125;
assign w27402 = ~w2061 & ~w2060;
assign w27403 = ~w2212 & ~w2211;
assign w27404 = w2239 & ~w2235;
assign w27405 = w2385 & ~w2381;
assign w27406 = w2732 & ~w2728;
assign w27407 = w2932 & ~w2928;
assign w27408 = ~w3511 & w33869;
assign w27409 = ~w4147 & w27721;
assign w27410 = ~w5081 & ~w5079;
assign w27411 = w5139 & ~w5335;
assign w27412 = ~w5567 & ~w5566;
assign w27413 = ~w5561 & ~w5560;
assign w27414 = w27722 | w27723;
assign w27415 = w27724 & w27725;
assign w27416 = w5907 & ~w6083;
assign w27417 = w6079 & ~w6075;
assign w27418 = ~w27343 & ~w6330;
assign w27419 = w7596 & w33870;
assign w27420 = (w8203 & w27821) | (w8203 & w27822) | (w27821 & w27822);
assign w27421 = (w25081 & w27823) | (w25081 & w27824) | (w27823 & w27824);
assign w27422 = w9314 & w8972;
assign w27423 = w9314 & ~w25086;
assign w27424 = ~w9314 & ~w8972;
assign w27425 = ~w9314 & w25086;
assign w27426 = ~w27058 & ~w9954;
assign w27427 = ~w10167 & ~w10166;
assign w27428 = ~w10167 & ~w10412;
assign w27429 = ~w10421 & w27518;
assign w27430 = w10516 & ~w10692;
assign w27431 = ~w26214 & w26213;
assign w27432 = ~w11038 & w11048;
assign w27433 = w11038 & ~w11048;
assign w27434 = ~w11055 & w11059;
assign w27435 = w11077 & ~w11073;
assign w27436 = ~w11254 & w11499;
assign w27437 = ~w11495 & ~w11496;
assign w27438 = (w25151 & w25150) | (w25151 & ~w15168) | (w25150 & ~w15168);
assign w27439 = (w25151 & w25150) | (w25151 & w25146) | (w25150 & w25146);
assign w27440 = w10750 & w27825;
assign w27441 = ~w11108 & ~w25871;
assign w27442 = ~w11108 & w27241;
assign w27443 = ~w10965 & ~w10964;
assign w27444 = ~w11379 & ~w11378;
assign w27445 = ~w15 & a_62;
assign w27446 = w11623 & a_62;
assign w27447 = w11575 & ~w11712;
assign w27448 = ~w11713 & ~w11385;
assign w27449 = ~w11713 & w27247;
assign w27450 = ~w12892 & ~w12890;
assign w27451 = w549 & w526;
assign w27452 = w549 & ~w27200;
assign w27453 = ~w548 & ~w27397;
assign w27454 = ~w548 & ~w27396;
assign w27455 = ~w10571 & w11326;
assign w27456 = w10571 & ~w11326;
assign w27457 = w11387 & w10982;
assign w27458 = w11387 & ~w27181;
assign w27459 = ~w11387 & ~w10982;
assign w27460 = ~w11387 & w27181;
assign w27461 = ~w11344 & w10931;
assign w27462 = ~w11344 & ~w11345;
assign w27463 = ~w26920 & a_62;
assign w27464 = w11627 & w11611;
assign w27465 = ~w26833 & ~w11662;
assign w27466 = w11576 & w33871;
assign w27467 = (~w11678 & ~w11576) | (~w11678 & w33872) | (~w11576 & w33872);
assign w27468 = ~w26925 & a_62;
assign w27469 = w12034 & w27765;
assign w27470 = (~w12048 & ~w12034) | (~w12048 & w27777) | (~w12034 & w27777);
assign w27471 = w11753 & ~w11749;
assign w27472 = w11934 & ~w12031;
assign w27473 = w11629 & w12381;
assign w27474 = ~w11629 & w12381;
assign w27475 = w11666 & ~w12024;
assign w27476 = ~w12065 & w11933;
assign w27477 = w12103 & ~w12099;
assign w27478 = ~w13271 & w13272;
assign w27479 = w13271 & ~w13272;
assign w27480 = (a_23 & ~w13463) | (a_23 & w33873) | (~w13463 & w33873);
assign w27481 = a_23 & ~w26666;
assign w27482 = (w13317 & w37858) | (w13317 & w37859) | (w37858 & w37859);
assign w27483 = (~w13718 & w13330) | (~w13718 & w27482) | (w13330 & w27482);
assign w27484 = a_20 & ~w26326;
assign w27485 = w25952 & a_20;
assign w27486 = a_23 & ~w26671;
assign w27487 = w26328 & a_23;
assign w27488 = w14033 & ~w14036;
assign w27489 = a_20 & ~w26339;
assign w27490 = w25961 & a_20;
assign w27491 = (w14444 & w14191) | (w14444 & w33874) | (w14191 & w33874);
assign w27492 = w14802 & ~w14529;
assign w27493 = ~w3935 & ~w3933;
assign w27494 = ~w11444 & ~w11443;
assign w27495 = w8973 & w8619;
assign w27496 = (~w9747 & w10077) | (~w9747 & w27840) | (w10077 & w27840);
assign w27497 = ~w10088 & w9466;
assign w27498 = ~w11800 & ~w11460;
assign w27499 = ~w11800 & w11256;
assign w27500 = ~w11854 & ~w11853;
assign w27501 = ~w12616 & w12628;
assign w27502 = w12616 & ~w12628;
assign w27503 = ~w13009 & w13021;
assign w27504 = w13009 & ~w13021;
assign w27505 = ~w8345 & ~w8343;
assign w27506 = ~w8639 & ~w8637;
assign w27507 = ~w9008 & ~w9006;
assign w27508 = w25560 & w8987;
assign w27509 = ~w25560 & ~w8987;
assign w27510 = ~w11125 & ~w10797;
assign w27511 = ~w11125 & ~w10798;
assign w27512 = (~w8706 & ~w9013) | (~w8706 & w27826) | (~w9013 & w27826);
assign w27513 = ~w9024 & w8710;
assign w27514 = w9974 & ~w9987;
assign w27515 = ~w9974 & w9987;
assign w27516 = ~w11401 & ~w10999;
assign w27517 = ~w11401 & w10866;
assign w27518 = ~w10422 & ~w10420;
assign w27519 = w811 & ~w815;
assign w27520 = w816 & ~w907;
assign w27521 = ~w1224 & ~w1222;
assign w27522 = w1358 & ~w1354;
assign w27523 = w1386 & ~w1485;
assign w27524 = w1902 & ~w1914;
assign w27525 = ~w4375 & ~w4374;
assign w27526 = ~w5819 & ~w5817;
assign w27527 = ~w5796 & ~w5795;
assign w27528 = w6077 & ~w6079;
assign w27529 = ~w6077 & w6079;
assign w27530 = w5906 & ~w6100;
assign w27531 = ~w6366 & w33875;
assign w27532 = ~w6355 & ~w6354;
assign w27533 = ~w6591 & w33876;
assign w27534 = (w6897 & ~w6885) | (w6897 & w33877) | (~w6885 & w33877);
assign w27535 = w6885 & w33878;
assign w27536 = w6706 & ~w6882;
assign w27537 = ~w6587 & w33879;
assign w27538 = ~w7473 & ~w7475;
assign w27539 = ~w7473 & ~w7197;
assign w27540 = w8478 & ~w8746;
assign w27541 = w10342 & w10006;
assign w27542 = w10342 & w10007;
assign w27543 = ~w10342 & ~w10006;
assign w27544 = ~w10342 & ~w10007;
assign w27545 = ~w11033 & ~w26214;
assign w27546 = ~w11033 & ~w26213;
assign w27547 = w10841 & ~w11131;
assign w27548 = ~w11051 & ~w11050;
assign w27549 = ~w11697 & w11575;
assign w27550 = w11735 & ~w11731;
assign w27551 = ~w12136 & w12138;
assign w27552 = w12136 & ~w12138;
assign w27553 = w25446 & ~w12570;
assign w27554 = w12622 & w33880;
assign w27555 = w12121 & ~w12523;
assign w27556 = w13015 & w33881;
assign w27557 = w13321 & w33882;
assign w27558 = (a_17 & ~w13436) | (a_17 & w33883) | (~w13436 & w33883);
assign w27559 = a_17 & ~w26320;
assign w27560 = w13048 & ~w13312;
assign w27561 = w13449 & w33884;
assign w27562 = ~w13714 & ~w13715;
assign w27563 = ~w12985 & w27778;
assign w27564 = ~w13329 & ~w13718;
assign w27565 = w13793 & w33885;
assign w27566 = ~w13719 & w13708;
assign w27567 = w14212 & w33886;
assign w27568 = w14536 & w33887;
assign w27569 = (~w26677 & w33888) | (~w26677 & w33889) | (w33888 & w33889);
assign w27570 = (a_26 & ~w14551) | (a_26 & w33890) | (~w14551 & w33890);
assign w27571 = a_26 & ~w26347;
assign w27572 = w14788 & w33891;
assign w27573 = ~w14867 & ~w14868;
assign w27574 = w14878 & w33892;
assign w27575 = w14784 & ~w14796;
assign w27576 = w14560 & w14777;
assign w27577 = a_26 & w14924;
assign w27578 = a_26 & ~w26678;
assign w27579 = ~a_26 & ~w14924;
assign w27580 = ~a_26 & w26678;
assign w27581 = ~w15153 & ~w15152;
assign w27582 = (a_23 & ~w15200) | (a_23 & w33893) | (~w15200 & w33893);
assign w27583 = a_23 & ~w26355;
assign w27584 = w15456 & w15443;
assign w27585 = (w9770 & w33894) | (w9770 & w33895) | (w33894 & w33895);
assign w27586 = (w15804 & w15578) | (w15804 & w33896) | (w15578 & w33896);
assign w27587 = a_32 & w16260;
assign w27588 = a_32 & ~w26683;
assign w27589 = ~a_32 & ~w16260;
assign w27590 = ~a_32 & w26683;
assign w27591 = ~w16464 & w25664;
assign w27592 = (~w16464 & w15903) | (~w16464 & w33897) | (w15903 & w33897);
assign w27593 = (a_29 & ~w16568) | (a_29 & w33898) | (~w16568 & w33898);
assign w27594 = a_29 & ~w26685;
assign w27595 = w16769 & w33899;
assign w27596 = ~w16779 & ~w16778;
assign w27597 = (a_29 & ~w16842) | (a_29 & w33900) | (~w16842 & w33900);
assign w27598 = a_29 & ~w26373;
assign w27599 = (w17048 & w17035) | (w17048 & w33901) | (w17035 & w33901);
assign w27600 = a_29 & w17373;
assign w27601 = a_29 & ~w26376;
assign w27602 = ~a_29 & ~w17373;
assign w27603 = ~a_29 & w26376;
assign w27604 = w17480 & w33902;
assign w27605 = (a_35 & ~w17662) | (a_35 & w33903) | (~w17662 & w33903);
assign w27606 = a_35 & ~w26691;
assign w27607 = a_32 & ~w26382;
assign w27608 = w26001 & a_32;
assign w27609 = ~w17969 & ~w17970;
assign w27610 = ~w17690 & w33904;
assign w27611 = w17968 & ~w17791;
assign w27612 = (a_32 & ~w18065) | (a_32 & w33905) | (~w18065 & w33905);
assign w27613 = a_32 & ~w26388;
assign w27614 = w18241 & w33906;
assign w27615 = (a_38 & ~w18466) | (a_38 & w33907) | (~w18466 & w33907);
assign w27616 = a_38 & ~w26692;
assign w27617 = (a_35 & ~w18484) | (a_35 & w33908) | (~w18484 & w33908);
assign w27618 = a_35 & ~w26693;
assign w27619 = w18757 & w33909;
assign w27620 = w19033 & w33910;
assign w27621 = w19274 & w33911;
assign w27622 = w19292 & w33912;
assign w27623 = w19520 & w33913;
assign w27624 = (a_41 & ~w19779) | (a_41 & w33914) | (~w19779 & w33914);
assign w27625 = a_41 & ~w26694;
assign w27626 = w19964 & w33915;
assign w27627 = (a_47 & ~w19982) | (a_47 & w33916) | (~w19982 & w33916);
assign w27628 = a_47 & ~w26695;
assign w27629 = (a_44 & ~w19999) | (a_44 & w33917) | (~w19999 & w33917);
assign w27630 = a_44 & ~w26696;
assign w27631 = a_41 & ~w26697;
assign w27632 = w26394 & a_41;
assign w27633 = w20023 & ~w20026;
assign w27634 = (a_47 & ~w20110) | (a_47 & w33918) | (~w20110 & w33918);
assign w27635 = a_47 & ~w26699;
assign w27636 = w20121 & w33919;
assign w27637 = a_44 & ~w26700;
assign w27638 = w26395 & a_44;
assign w27639 = (a_41 & ~w20238) | (a_41 & w33920) | (~w20238 & w33920);
assign w27640 = a_41 & ~w26396;
assign w27641 = w20278 & ~w20345;
assign w27642 = w20703 & ~w20564;
assign w27643 = ~w20703 & ~w20704;
assign w27644 = w20798 & w33921;
assign w27645 = (a_47 & ~w20893) | (a_47 & w33922) | (~w20893 & w33922);
assign w27646 = a_47 & ~w26704;
assign w27647 = w20910 & w33923;
assign w27648 = w21325 & ~w21199;
assign w27649 = ~w21325 & ~w21326;
assign w27650 = (w21573 & w21559) | (w21573 & w33924) | (w21559 & w33924);
assign w27651 = w21534 & ~w21523;
assign w27652 = (w21517 & w21503) | (w21517 & w33925) | (w21503 & w33925);
assign w27653 = a_53 & ~w26433;
assign w27654 = w26018 & a_53;
assign w27655 = w21637 & w33926;
assign w27656 = a_47 & ~w26436;
assign w27657 = w26022 & a_47;
assign w27658 = w21728 & ~w21620;
assign w27659 = w21620 & ~w21728;
assign w27660 = (w21923 & w21920) | (w21923 & w33927) | (w21920 & w33927);
assign w27661 = ~w21920 & w33928;
assign w27662 = w21769 & ~w21758;
assign w27663 = w21990 & w33929;
assign w27664 = (a_53 & ~w22049) | (a_53 & w33930) | (~w22049 & w33930);
assign w27665 = a_53 & ~w26716;
assign w27666 = w22066 & w33931;
assign w27667 = w22186 & w33932;
assign w27668 = a_53 & ~w26445;
assign w27669 = w26035 & a_53;
assign w27670 = w22250 & ~w22252;
assign w27671 = ~w22450 & w22451;
assign w27672 = w22450 & ~w22451;
assign w27673 = ~w22638 & w22639;
assign w27674 = w22638 & ~w22639;
assign w27675 = (a_59 & ~w22730) | (a_59 & w33933) | (~w22730 & w33933);
assign w27676 = a_59 & ~w26453;
assign w27677 = w22751 & w22743;
assign w27678 = ~w22877 & ~w22880;
assign w27679 = ~w22936 & w22937;
assign w27680 = w22936 & ~w22937;
assign w27681 = w22840 & ~w22913;
assign w27682 = ~w23102 & w23103;
assign w27683 = w23102 & ~w23103;
assign w27684 = (a_59 & ~w23202) | (a_59 & w33934) | (~w23202 & w33934);
assign w27685 = a_59 & ~w26722;
assign w27686 = w23302 & w33935;
assign w27687 = a_62 & ~w26723;
assign w27688 = w26477 & a_62;
assign w27689 = (~w6682 & w33936) | (~w6682 & w33937) | (w33936 & w33937);
assign w27690 = a_59 & ~w26725;
assign w27691 = w26478 & a_59;
assign w27692 = w23347 & ~w23350;
assign w27693 = ~w23347 & w23350;
assign w27694 = w23466 & w33938;
assign w27695 = w23596 & w33939;
assign w27696 = (w23607 & w23733) | (w23607 & w33940) | (w23733 & w33940);
assign w27697 = (~w26727 & w23733) | (~w26727 & w33941) | (w23733 & w33941);
assign w27698 = w23742 & w33942;
assign w27699 = w23756 & w33943;
assign w27700 = ~w23951 & ~w26487;
assign w27701 = ~w23951 & ~w26488;
assign w27702 = (a_62 & ~w24063) | (a_62 & w33944) | (~w24063 & w33944);
assign w27703 = (a_62 & ~w24064) | (a_62 & w27446) | (~w24064 & w27446);
assign w27704 = a_62 & ~w26490;
assign w27705 = w26072 & a_62;
assign w27706 = (~w9110 & w33945) | (~w9110 & w33946) | (w33945 & w33946);
assign w27707 = w24334 & w33947;
assign w27708 = w24344 & w33948;
assign w27709 = (a_62 & ~w24592) | (a_62 & w33950) | (~w24592 & w33950);
assign w27710 = a_62 & ~w26964;
assign w27711 = (a_62 & ~w24689) | (a_62 & w33951) | (~w24689 & w33951);
assign w27712 = ~w7458 & ~w7456;
assign w27713 = ~w10427 & ~w10809;
assign w27714 = w12278 & w12259;
assign w27715 = (w12278 & w12256) | (w12278 & w33952) | (w12256 & w33952);
assign w27716 = ~w10037 & ~w10035;
assign w27717 = ~w7692 & ~w7690;
assign w27718 = ~w10409 & ~w10779;
assign w27719 = ~w12118 & ~w11767;
assign w27720 = ~w12118 & w11574;
assign w27721 = ~w4148 & ~w4146;
assign w27722 = w6098 & w5907;
assign w27723 = (w6098 & w6085) | (w6098 & w33953) | (w6085 & w33953);
assign w27724 = ~w6098 & ~w5907;
assign w27725 = ~w6085 & w33954;
assign w27726 = ~w708 & ~w707;
assign w27727 = w900 & w1018;
assign w27728 = ~w900 & ~w1018;
assign w27729 = w1024 & ~w1134;
assign w27730 = w1135 & ~w1130;
assign w27731 = w1488 & w33955;
assign w27732 = ~w1769 & w33956;
assign w27733 = (w1772 & w33957) | (w1772 & w33958) | (w33957 & w33958);
assign w27734 = ~w4614 & ~w4613;
assign w27735 = ~w6106 & w33959;
assign w27736 = ~w6632 & ~w6630;
assign w27737 = (w27736 & w33960) | (w27736 & w33961) | (w33960 & w33961);
assign w27738 = w7228 & ~w7224;
assign w27739 = ~w8022 & w8024;
assign w27740 = w8022 & ~w8024;
assign w27741 = w7809 & ~w7805;
assign w27742 = w7823 & w25071;
assign w27743 = ~w25071 & ~w8127;
assign w27744 = (~w8127 & ~w25071) | (~w8127 & w33962) | (~w25071 & w33962);
assign w27745 = ~w8757 & w8746;
assign w27746 = ~w8757 & ~w8744;
assign w27747 = (w26598 & w33963) | (w26598 & w33964) | (w33963 & w33964);
assign w27748 = w9403 & ~w9414;
assign w27749 = ~w9397 & w9400;
assign w27750 = w9699 & ~w9695;
assign w27751 = ~w10053 & w10056;
assign w27752 = w11097 & ~w11107;
assign w27753 = ~w11255 & ~w11254;
assign w27754 = ~w11255 & ~w11499;
assign w27755 = w12122 & ~w12133;
assign w27756 = ~w12122 & ~w12133;
assign w27757 = (w25146 & w33965) | (w25146 & w33966) | (w33965 & w33966);
assign w27758 = (w25155 & w25156) | (w25155 & w27438) | (w25156 & w27438);
assign w27759 = ~w11930 & w12206;
assign w27760 = ~w11930 & ~w12206;
assign w27761 = (w26307 & w33967) | (w26307 & w33968) | (w33967 & w33968);
assign w27762 = (~w26307 & w33969) | (~w26307 & w33970) | (w33969 & w33970);
assign w27763 = (~w15436 & w15221) | (~w15436 & w33971) | (w15221 & w33971);
assign w27764 = ~w11017 & ~w11015;
assign w27765 = ~w11934 & ~w12048;
assign w27766 = w732 & w707;
assign w27767 = w732 & ~w27726;
assign w27768 = w12954 & w33972;
assign w27769 = (~w12967 & ~w12954) | (~w12967 & w33973) | (~w12954 & w33973);
assign w27770 = ~w26314 & w33974;
assign w27771 = (w13442 & ~w13311) | (w13442 & w33975) | (~w13311 & w33975);
assign w27772 = w13442 & w13315;
assign w27773 = w13311 & w33976;
assign w27774 = ~w13442 & ~w13315;
assign w27775 = (w25163 & w25162) | (w25163 & ~w27757) | (w25162 & ~w27757);
assign w27776 = w17078 & ~w17089;
assign w27777 = w11934 & ~w12048;
assign w27778 = (~w13718 & ~w12980) | (~w13718 & w33978) | (~w12980 & w33978);
assign w27779 = (~w731 & ~w732) | (~w731 & w33979) | (~w732 & w33979);
assign w27780 = (~w731 & w27726) | (~w731 & w33980) | (w27726 & w33980);
assign w27781 = w12299 & ~w12576;
assign w27782 = (~w13302 & w26314) | (~w13302 & w33981) | (w26314 & w33981);
assign w27783 = w12970 & ~w13307;
assign w27784 = ~w13704 & ~w13703;
assign w27785 = (~w13398 & ~w13399) | (~w13398 & w27827) | (~w13399 & w27827);
assign w27786 = (~w13398 & w25452) | (~w13398 & w25139) | (w25452 & w25139);
assign w27787 = ~w13415 & w13749;
assign w27788 = ~w13415 & ~w13416;
assign w27789 = ~w27784 & ~w13444;
assign w27790 = (w13696 & w13290) | (w13696 & w33982) | (w13290 & w33982);
assign w27791 = w13695 & ~w13485;
assign w27792 = ~w13456 & w33983;
assign w27793 = w14100 & ~w14087;
assign w27794 = ~w13742 & w13730;
assign w27795 = ~w13742 & ~w13744;
assign w27796 = ~w14088 & w33984;
assign w27797 = (~w14136 & w14098) | (~w14136 & w33985) | (w14098 & w33985);
assign w27798 = ~w307 & w11623;
assign w27799 = ~w14070 & w33986;
assign w27800 = (~w14468 & w14080) | (~w14468 & w33987) | (w14080 & w33987);
assign w27801 = (a_23 & ~w14536) | (a_23 & w33988) | (~w14536 & w33988);
assign w27802 = a_23 & ~w27568;
assign w27803 = (a_20 & ~w14892) | (a_20 & w33989) | (~w14892 & w33989);
assign w27804 = a_20 & ~w26350;
assign w27805 = (w14780 & w14543) | (w14780 & w33990) | (w14543 & w33990);
assign w27806 = a_17 & ~w26353;
assign w27807 = w25973 & a_17;
assign w27808 = a_23 & ~w27582;
assign w27809 = w26355 & a_23;
assign w27810 = (w15461 & w15193) | (w15461 & w33991) | (w15193 & w33991);
assign w27811 = (~w15221 & w33992) | (~w15221 & w33993) | (w33992 & w33993);
assign w27812 = w15812 & w33994;
assign w27813 = w15566 & ~w15826;
assign w27814 = w15868 & w33995;
assign w27815 = ~w16127 & ~w16126;
assign w27816 = w16131 & ~w16142;
assign w27817 = (~w12988 & ~w13333) | (~w12988 & w33996) | (~w13333 & w33996);
assign w27818 = ~w13009 & ~w13021;
assign w27819 = w10070 & ~w10166;
assign w27820 = (w8406 & ~w8072) | (w8406 & w33997) | (~w8072 & w33997);
assign w27821 = (~w8390 & ~w8677) | (~w8390 & w33998) | (~w8677 & w33998);
assign w27822 = ~w8688 & w25401;
assign w27823 = (~w8423 & ~w8713) | (~w8423 & w33999) | (~w8713 & w33999);
assign w27824 = ~w8724 & w8427;
assign w27825 = ~w10760 & ~w11090;
assign w27826 = (w9023 & ~w8695) | (w9023 & w34000) | (~w8695 & w34000);
assign w27827 = ~w13398 & ~w13031;
assign w27828 = (w9745 & ~w9467) | (w9745 & w34001) | (~w9467 & w34001);
assign w27829 = w9467 & w34002;
assign w27830 = ~w10409 & ~w10408;
assign w27831 = w11097 & w11107;
assign w27832 = ~w11097 & ~w11107;
assign w27833 = w11127 & w10797;
assign w27834 = w11127 & w10798;
assign w27835 = ~w11127 & ~w10797;
assign w27836 = ~w11127 & ~w10798;
assign w27837 = ~w12606 & w34003;
assign w27838 = ~w12583 & w12288;
assign w27839 = ~w12678 & w34004;
assign w27840 = (~w9734 & w34005) | (~w9734 & w34006) | (w34005 & w34006);
assign w27841 = w34007 & w17;
assign w27842 = (~w17 & ~a_2) | (~w17 & ~w1) | (~a_2 & ~w1);
assign w27843 = a_0 & b_2;
assign w27844 = a_0 & b_4;
assign w27845 = w27010 & b_2;
assign w27846 = w76 & w34008;
assign w27847 = (a_2 & ~w76) | (a_2 & w34009) | (~w76 & w34009);
assign w27848 = (a_2 & ~w76) | (a_2 & w34010) | (~w76 & w34010);
assign w27849 = ~b_0 & a_5;
assign w27850 = a_0 & b_5;
assign w27851 = w27010 & b_3;
assign w27852 = w122 & w34011;
assign w27853 = a_0 & b_6;
assign w27854 = w27010 & b_4;
assign w27855 = w183 & w34012;
assign w27856 = a_0 & b_7;
assign w27857 = w27010 & b_5;
assign w27858 = ~w210 & w26520;
assign w27859 = ~w210 & w26519;
assign w27860 = w206 & w34013;
assign w27861 = ~b_0 & a_8;
assign w27862 = a_0 & b_8;
assign w27863 = w27010 & b_6;
assign w27864 = (~w209 & w26520) | (~w209 & w34014) | (w26520 & w34014);
assign w27865 = (~w209 & w26519) | (~w209 & w34014) | (w26519 & w34014);
assign w27866 = ~w307 & w12;
assign w27867 = (a_2 & ~w302) | (a_2 & w34015) | (~w302 & w34015);
assign w27868 = ~w27867 & a_2;
assign w27869 = w93 & b_4;
assign w27870 = w325 & w34016;
assign w27871 = a_0 & b_9;
assign w27872 = w27010 & b_7;
assign w27873 = ~w305 & ~w368;
assign w27874 = w364 & w34017;
assign w27875 = w93 & b_5;
assign w27876 = w389 & w34018;
assign w27877 = w248 & w335;
assign w27878 = w349 & ~w396;
assign w27879 = ~b_0 & a_11;
assign w27880 = a_0 & b_10;
assign w27881 = w27010 & b_8;
assign w27882 = ~w451 & w27017;
assign w27883 = ~w451 & w27016;
assign w27884 = w447 & w34019;
assign w27885 = ~w437 & w34020;
assign w27886 = w93 & b_6;
assign w27887 = ~w307 & w102;
assign w27888 = (a_5 & ~w471) | (a_5 & w34021) | (~w471 & w34021);
assign w27889 = ~w27888 & a_5;
assign w27890 = a_0 & b_11;
assign w27891 = w27010 & b_9;
assign w27892 = w527 & ~w27199;
assign w27893 = w527 & ~w27198;
assign w27894 = ~w527 & w27199;
assign w27895 = ~w527 & w27198;
assign w27896 = w523 & w34022;
assign w27897 = a_0 & b_12;
assign w27898 = w27010 & b_10;
assign w27899 = (w27198 & w34023) | (w27198 & w34024) | (w34023 & w34024);
assign w27900 = ~w549 & w27330;
assign w27901 = w545 & w34025;
assign w27902 = w233 & b_4;
assign w27903 = w561 & w34026;
assign w27904 = w93 & b_7;
assign w27905 = w600 & w34027;
assign w27906 = w233 & b_5;
assign w27907 = w628 & w34028;
assign w27908 = w427 & w571;
assign w27909 = w585 & ~w635;
assign w27910 = ~b_0 & a_14;
assign w27911 = w93 & b_8;
assign w27912 = w686 & w34029;
assign w27913 = a_0 & b_13;
assign w27914 = w27010 & b_11;
assign w27915 = w703 & w34030;
assign w27916 = a_0 & b_14;
assign w27917 = w27010 & b_12;
assign w27918 = ~w732 & ~w707;
assign w27919 = ~w732 & w27726;
assign w27920 = w728 & w34031;
assign w27921 = w93 & b_9;
assign w27922 = w744 & w34032;
assign w27923 = ~w676 & w34033;
assign w27924 = w233 & b_6;
assign w27925 = ~w307 & w242;
assign w27926 = (a_8 & ~w789) | (a_8 & w34034) | (~w789 & w34034);
assign w27927 = ~w27926 & a_8;
assign w27928 = a_0 & b_15;
assign w27929 = w27010 & b_13;
assign w27930 = w824 & ~w27779;
assign w27931 = w824 & ~w27780;
assign w27932 = ~w824 & w27779;
assign w27933 = ~w824 & w27780;
assign w27934 = w820 & w34035;
assign w27935 = ~w805 & ~w804;
assign w27936 = w93 & b_10;
assign w27937 = w837 & w34036;
assign w27938 = w233 & b_7;
assign w27939 = w848 & w34037;
assign w27940 = w412 & b_4;
assign w27941 = w858 & w34038;
assign w27942 = a_0 & b_16;
assign w27943 = w27010 & b_14;
assign w27944 = (~w823 & w27779) | (~w823 & w34039) | (w27779 & w34039);
assign w27945 = (~w823 & w27780) | (~w823 & w34039) | (w27780 & w34039);
assign w27946 = w919 & w34040;
assign w27947 = w833 & ~w900;
assign w27948 = w93 & b_11;
assign w27949 = w936 & w34041;
assign w27950 = w233 & b_8;
assign w27951 = w946 & w34042;
assign w27952 = w412 & b_5;
assign w27953 = w957 & w34043;
assign w27954 = w666 & w868;
assign w27955 = w882 & ~w964;
assign w27956 = ~b_0 & a_17;
assign w27957 = a_0 & b_17;
assign w27958 = w27010 & b_15;
assign w27959 = ~w923 & ~w922;
assign w27960 = w1035 & w922;
assign w27961 = w1035 & ~w27959;
assign w27962 = ~w1035 & ~w922;
assign w27963 = ~w1035 & w27959;
assign w27964 = w1031 & w34044;
assign w27965 = w93 & b_12;
assign w27966 = w1048 & w34045;
assign w27967 = w233 & b_9;
assign w27968 = w1059 & w34046;
assign w27969 = ~w1006 & ~w1005;
assign w27970 = w412 & b_6;
assign w27971 = ~w307 & w421;
assign w27972 = (a_11 & ~w1104) | (a_11 & w34047) | (~w1104 & w34047);
assign w27973 = ~w27972 & a_11;
assign w27974 = w93 & b_13;
assign w27975 = w1143 & w34048;
assign w27976 = w233 & b_10;
assign w27977 = w1154 & w34049;
assign w27978 = w1066 & ~w1113;
assign w27979 = w651 & b_4;
assign w27980 = w1165 & w34050;
assign w27981 = w412 & b_7;
assign w27982 = w1203 & w34051;
assign w27983 = a_0 & b_18;
assign w27984 = w27010 & b_16;
assign w27985 = (~w1034 & ~w1035) | (~w1034 & w34052) | (~w1035 & w34052);
assign w27986 = (~w1034 & w27959) | (~w1034 & w34053) | (w27959 & w34053);
assign w27987 = w1235 & ~w27985;
assign w27988 = w1235 & ~w27986;
assign w27989 = ~w1235 & w27985;
assign w27990 = ~w1235 & w27986;
assign w27991 = w1231 & w34054;
assign w27992 = w93 & b_14;
assign w27993 = w1255 & w34055;
assign w27994 = w651 & b_5;
assign w27995 = w1266 & w34056;
assign w27996 = w995 & w1175;
assign w27997 = w1189 & ~w1273;
assign w27998 = ~b_0 & a_20;
assign w27999 = w412 & b_8;
assign w28000 = w1322 & w34057;
assign w28001 = w233 & b_11;
assign w28002 = w1340 & w34058;
assign w28003 = ~w1218 & ~w1217;
assign w28004 = a_0 & b_19;
assign w28005 = w27010 & b_17;
assign w28006 = (~w1234 & w27985) | (~w1234 & w34059) | (w27985 & w34059);
assign w28007 = w1369 & ~w28006;
assign w28008 = (~w27986 & w34060) | (~w27986 & w34061) | (w34060 & w34061);
assign w28009 = ~w1369 & w28006;
assign w28010 = (w27986 & w34062) | (w27986 & w34063) | (w34062 & w34063);
assign w28011 = ~w12 & w1366;
assign w28012 = w93 & b_15;
assign w28013 = w1390 & w34064;
assign w28014 = w233 & b_12;
assign w28015 = w1400 & w34065;
assign w28016 = w412 & b_9;
assign w28017 = w1411 & w34066;
assign w28018 = ~w1315 & ~w1313;
assign w28019 = w651 & b_6;
assign w28020 = ~w307 & w660;
assign w28021 = (a_14 & ~w1457) | (a_14 & w34067) | (~w1457 & w34067);
assign w28022 = ~w28021 & a_14;
assign w28023 = a_0 & b_20;
assign w28024 = w27010 & b_18;
assign w28025 = w1368 & w1500;
assign w28026 = ~w1368 & ~w1500;
assign w28027 = w1496 & w34068;
assign w28028 = ~w1379 & w34069;
assign w28029 = w233 & b_13;
assign w28030 = w1521 & w34070;
assign w28031 = w412 & b_10;
assign w28032 = w1532 & w34071;
assign w28033 = w1418 & ~w1466;
assign w28034 = w980 & b_4;
assign w28035 = w1543 & w34072;
assign w28036 = w651 & b_7;
assign w28037 = w1581 & w34073;
assign w28038 = w93 & b_16;
assign w28039 = w1609 & w34074;
assign w28040 = a_0 & b_21;
assign w28041 = w27010 & b_19;
assign w28042 = ~w1499 & ~w1500;
assign w28043 = (~w1499 & ~w1500) | (~w1499 & w34075) | (~w1500 & w34075);
assign w28044 = w1631 & ~w28042;
assign w28045 = w1631 & ~w28043;
assign w28046 = ~w1631 & w28042;
assign w28047 = ~w1631 & w28043;
assign w28048 = w1627 & w34076;
assign w28049 = w1513 & ~w1509;
assign w28050 = w233 & b_14;
assign w28051 = w1653 & w34077;
assign w28052 = ~w1596 & ~w1595;
assign w28053 = w980 & b_5;
assign w28054 = w1665 & w34078;
assign w28055 = w1304 & w1553;
assign w28056 = w1567 & ~w1672;
assign w28057 = ~b_0 & a_23;
assign w28058 = w651 & b_8;
assign w28059 = w1721 & w34079;
assign w28060 = w412 & b_11;
assign w28061 = w1739 & w34080;
assign w28062 = w93 & b_17;
assign w28063 = w1761 & w34081;
assign w28064 = a_0 & b_22;
assign w28065 = w27010 & b_20;
assign w28066 = (~w1630 & w28042) | (~w1630 & w34082) | (w28042 & w34082);
assign w28067 = (~w1630 & w28043) | (~w1630 & w34082) | (w28043 & w34082);
assign w28068 = w1783 & ~w28066;
assign w28069 = w1783 & ~w28067;
assign w28070 = ~w1783 & w28066;
assign w28071 = ~w1783 & w28067;
assign w28072 = w1779 & w34083;
assign w28073 = ~w1754 & ~w1752;
assign w28074 = w233 & b_15;
assign w28075 = w1802 & w34084;
assign w28076 = w412 & b_12;
assign w28077 = w1812 & w34085;
assign w28078 = w651 & b_9;
assign w28079 = w1823 & w34086;
assign w28080 = ~w1714 & ~w1712;
assign w28081 = w980 & b_6;
assign w28082 = ~w307 & w989;
assign w28083 = (a_17 & ~w1869) | (a_17 & w34087) | (~w1869 & w34087);
assign w28084 = ~w28083 & a_17;
assign w28085 = w1898 & ~w1798;
assign w28086 = ~w1898 & ~w1798;
assign w28087 = w93 & b_18;
assign w28088 = w1908 & w34088;
assign w28089 = a_0 & b_23;
assign w28090 = w27010 & b_21;
assign w28091 = (~w1782 & w28067) | (~w1782 & w34089) | (w28067 & w34089);
assign w28092 = (~w28066 & w34090) | (~w28066 & w34091) | (w34090 & w34091);
assign w28093 = (~w28067 & w34090) | (~w28067 & w34091) | (w34090 & w34091);
assign w28094 = (w28066 & w34092) | (w28066 & w34093) | (w34092 & w34093);
assign w28095 = ~w1930 & w28091;
assign w28096 = w1926 & w34094;
assign w28097 = ~w1794 & ~w1793;
assign w28098 = w93 & b_19;
assign w28099 = w1951 & w34095;
assign w28100 = w412 & b_13;
assign w28101 = w1962 & w34096;
assign w28102 = w651 & b_10;
assign w28103 = w1973 & w34097;
assign w28104 = w1830 & ~w1878;
assign w28105 = w1289 & b_4;
assign w28106 = w1984 & w34098;
assign w28107 = w980 & b_7;
assign w28108 = w2022 & w34099;
assign w28109 = w233 & b_16;
assign w28110 = w2052 & w34100;
assign w28111 = a_0 & b_24;
assign w28112 = w27010 & b_22;
assign w28113 = w1929 & w2080;
assign w28114 = ~w1929 & ~w2080;
assign w28115 = w2076 & w34101;
assign w28116 = w2093 & ~w2089;
assign w28117 = a_0 & b_25;
assign w28118 = w27010 & b_23;
assign w28119 = ~w2079 & ~w2080;
assign w28120 = (~w2079 & ~w2080) | (~w2079 & w34102) | (~w2080 & w34102);
assign w28121 = w2105 & ~w28119;
assign w28122 = w2105 & ~w28120;
assign w28123 = ~w2105 & w28119;
assign w28124 = ~w2105 & w28120;
assign w28125 = w2101 & w34103;
assign w28126 = w412 & b_14;
assign w28127 = w2118 & w34104;
assign w28128 = w1289 & b_5;
assign w28129 = w2129 & w34105;
assign w28130 = w1703 & w1994;
assign w28131 = w2008 & ~w2136;
assign w28132 = ~b_0 & a_26;
assign w28133 = w980 & b_8;
assign w28134 = w2185 & w34106;
assign w28135 = w651 & b_11;
assign w28136 = w2203 & w34107;
assign w28137 = ~w2037 & ~w2036;
assign w28138 = w233 & b_17;
assign w28139 = w2228 & w34108;
assign w28140 = w93 & b_20;
assign w28141 = w2246 & w34109;
assign w28142 = w2242 & w2252;
assign w28143 = ~w2242 & ~w2252;
assign w28144 = ~w2261 & ~w2259;
assign w28145 = w2242 & ~w2252;
assign w28146 = ~w2218 & w34110;
assign w28147 = w651 & b_12;
assign w28148 = w2273 & w34111;
assign w28149 = w980 & b_9;
assign w28150 = w2283 & w34112;
assign w28151 = ~w2178 & ~w2176;
assign w28152 = w1688 & b_3;
assign w28153 = (a_23 & ~w2311) | (a_23 & w34113) | (~w2311 & w34113);
assign w28154 = ~w2319 & ~w2173;
assign w28155 = ~w2319 & ~w25775;
assign w28156 = ~w2173 & w25775;
assign w28157 = w1289 & b_6;
assign w28158 = ~w307 & w1298;
assign w28159 = (a_20 & ~w2328) | (a_20 & w34114) | (~w2328 & w34114);
assign w28160 = ~w28159 & a_20;
assign w28161 = ~w2324 & w2335;
assign w28162 = w2324 & ~w2335;
assign w28163 = ~w2192 & ~w2344;
assign w28164 = w412 & b_15;
assign w28165 = w2358 & w34115;
assign w28166 = w233 & b_18;
assign w28167 = w2374 & w34116;
assign w28168 = w93 & b_21;
assign w28169 = w2392 & w34117;
assign w28170 = a_0 & b_26;
assign w28171 = w27010 & b_24;
assign w28172 = (~w2104 & w28119) | (~w2104 & w34118) | (w28119 & w34118);
assign w28173 = (~w2104 & w28120) | (~w2104 & w34118) | (w28120 & w34118);
assign w28174 = w2413 & ~w28172;
assign w28175 = w2413 & ~w28173;
assign w28176 = ~w2413 & w28172;
assign w28177 = ~w2413 & w28173;
assign w28178 = w2409 & w34119;
assign w28179 = w93 & b_22;
assign w28180 = w2432 & w34120;
assign w28181 = w651 & b_13;
assign w28182 = w2442 & w34121;
assign w28183 = w980 & b_10;
assign w28184 = w2453 & w34122;
assign w28185 = w1688 & b_4;
assign w28186 = w2464 & w34123;
assign w28187 = w1289 & b_7;
assign w28188 = w2502 & w34124;
assign w28189 = w412 & b_16;
assign w28190 = (a_11 & ~w2532) | (a_11 & w34125) | (~w2532 & w34125);
assign w28191 = a_11 & ~w24997;
assign w28192 = a_11 & ~w28190;
assign w28193 = w24997 & a_11;
assign w28194 = w233 & b_19;
assign w28195 = w2550 & w34126;
assign w28196 = ~w2400 & w34127;
assign w28197 = a_0 & b_27;
assign w28198 = w27010 & b_25;
assign w28199 = (~w2412 & w28173) | (~w2412 & w34128) | (w28173 & w34128);
assign w28200 = (~w28172 & w34129) | (~w28172 & w34130) | (w34129 & w34130);
assign w28201 = (~w28173 & w34129) | (~w28173 & w34130) | (w34129 & w34130);
assign w28202 = (w28172 & w34131) | (w28172 & w34132) | (w34131 & w34132);
assign w28203 = ~w2579 & w28199;
assign w28204 = w2575 & w34133;
assign w28205 = ~w2590 & ~w2589;
assign w28206 = w93 & b_23;
assign w28207 = w2598 & w34134;
assign w28208 = w2323 & ~w2492;
assign w28209 = w1688 & b_5;
assign w28210 = w2610 & w34135;
assign w28211 = ~b_0 & a_29;
assign w28212 = w1289 & b_8;
assign w28213 = w2666 & w34136;
assign w28214 = w980 & b_11;
assign w28215 = (a_17 & ~w2684) | (a_17 & w34137) | (~w2684 & w34137);
assign w28216 = a_17 & ~w25000;
assign w28217 = a_17 & ~w28215;
assign w28218 = w25000 & a_17;
assign w28219 = w651 & b_14;
assign w28220 = (a_14 & ~w2703) | (a_14 & w34138) | (~w2703 & w34138);
assign w28221 = a_14 & ~w25002;
assign w28222 = a_14 & ~w28220;
assign w28223 = w25002 & a_14;
assign w28224 = w2698 & ~w2709;
assign w28225 = ~w2698 & ~w2709;
assign w28226 = ~w2521 & w2525;
assign w28227 = w412 & b_17;
assign w28228 = (a_11 & ~w2721) | (a_11 & w34139) | (~w2721 & w34139);
assign w28229 = a_11 & ~w25003;
assign w28230 = a_11 & ~w28228;
assign w28231 = w25003 & a_11;
assign w28232 = w233 & b_20;
assign w28233 = w2739 & w34140;
assign w28234 = ~w2559 & ~w2558;
assign w28235 = a_0 & b_28;
assign w28236 = w27010 & b_26;
assign w28237 = ~w2578 & ~w28200;
assign w28238 = ~w2578 & ~w28201;
assign w28239 = w2764 & w34141;
assign w28240 = ~w2754 & w34142;
assign w28241 = w93 & b_24;
assign w28242 = w2787 & w34143;
assign w28243 = w980 & b_12;
assign w28244 = w2798 & w34144;
assign w28245 = w1289 & b_9;
assign w28246 = w2809 & w34145;
assign w28247 = w1688 & b_6;
assign w28248 = ~w307 & w1697;
assign w28249 = (a_23 & ~w2855) | (a_23 & w34146) | (~w2855 & w34146);
assign w28250 = ~w28249 & a_23;
assign w28251 = w2695 & ~w2691;
assign w28252 = w651 & b_15;
assign w28253 = (a_14 & ~w2886) | (a_14 & w34147) | (~w2886 & w34147);
assign w28254 = a_14 & ~w25008;
assign w28255 = a_14 & ~w28253;
assign w28256 = w25008 & a_14;
assign w28257 = w412 & b_18;
assign w28258 = w2904 & w34148;
assign w28259 = ~w2911 & ~w2734;
assign w28260 = ~w2911 & ~w27205;
assign w28261 = ~w2734 & w27205;
assign w28262 = w233 & b_21;
assign w28263 = w2921 & w34149;
assign w28264 = w28261 & w34150;
assign w28265 = (~w2927 & ~w28261) | (~w2927 & w34151) | (~w28261 & w34151);
assign w28266 = a_0 & b_29;
assign w28267 = w27010 & b_27;
assign w28268 = ~w2768 & ~w2767;
assign w28269 = w2951 & w2767;
assign w28270 = w2951 & ~w28268;
assign w28271 = ~w2951 & ~w2767;
assign w28272 = ~w2951 & w28268;
assign w28273 = w2947 & w34152;
assign w28274 = w34153 & w34154;
assign w28275 = w980 & b_13;
assign w28276 = w2972 & w34155;
assign w28277 = w1289 & b_10;
assign w28278 = w2983 & w34156;
assign w28279 = w2816 & ~w2864;
assign w28280 = w2152 & b_4;
assign w28281 = w2994 & w34157;
assign w28282 = w1688 & b_7;
assign w28283 = w3032 & w34158;
assign w28284 = w2879 & ~w2875;
assign w28285 = w651 & b_16;
assign w28286 = (a_14 & ~w3062) | (a_14 & w34159) | (~w3062 & w34159);
assign w28287 = a_14 & ~w25010;
assign w28288 = a_14 & ~w28286;
assign w28289 = w25010 & a_14;
assign w28290 = w412 & b_19;
assign w28291 = w3080 & w34160;
assign w28292 = w233 & b_22;
assign w28293 = w3097 & w34161;
assign w28294 = w93 & b_25;
assign w28295 = w3113 & w34162;
assign w28296 = (w2757 & w34163) | (w2757 & w34164) | (w34163 & w34164);
assign w28297 = a_0 & b_30;
assign w28298 = w27010 & b_28;
assign w28299 = (~w2950 & ~w2951) | (~w2950 & w34165) | (~w2951 & w34165);
assign w28300 = (~w2950 & w28268) | (~w2950 & w34166) | (w28268 & w34166);
assign w28301 = w3135 & ~w28299;
assign w28302 = w3135 & ~w28300;
assign w28303 = ~w3135 & w28299;
assign w28304 = ~w3135 & w28300;
assign w28305 = w3131 & w34167;
assign w28306 = ~w2780 & w34168;
assign w28307 = w980 & b_14;
assign w28308 = w3155 & w34169;
assign w28309 = w2152 & b_5;
assign w28310 = w3166 & w34170;
assign w28311 = w2648 & w3004;
assign w28312 = w3018 & ~w3173;
assign w28313 = ~b_0 & a_32;
assign w28314 = w1688 & b_8;
assign w28315 = (a_23 & ~w3222) | (a_23 & w34171) | (~w3222 & w34171);
assign w28316 = a_23 & ~w25011;
assign w28317 = w1289 & b_11;
assign w28318 = w3240 & w34172;
assign w28319 = ~w3047 & ~w3046;
assign w28320 = w651 & b_17;
assign w28321 = (a_14 & ~w3265) | (a_14 & w34173) | (~w3265 & w34173);
assign w28322 = a_14 & ~w25012;
assign w28323 = w3265 & w34174;
assign w28324 = a_14 & w25012;
assign w28325 = w412 & b_20;
assign w28326 = (a_11 & ~w3283) | (a_11 & w34175) | (~w3283 & w34175);
assign w28327 = a_11 & ~w25013;
assign w28328 = a_11 & ~w28326;
assign w28329 = w25013 & a_11;
assign w28330 = w233 & b_23;
assign w28331 = w3302 & w34176;
assign w28332 = ~w3106 & ~w3104;
assign w28333 = w93 & b_26;
assign w28334 = w3320 & w34177;
assign w28335 = a_0 & b_31;
assign w28336 = w27010 & b_29;
assign w28337 = (~w3134 & w28299) | (~w3134 & w34178) | (w28299 & w34178);
assign w28338 = w3342 & ~w28337;
assign w28339 = (~w28300 & w34179) | (~w28300 & w34180) | (w34179 & w34180);
assign w28340 = ~w3342 & w28337;
assign w28341 = (w28300 & w34181) | (w28300 & w34182) | (w34181 & w34182);
assign w28342 = ~w12 & w3339;
assign w28343 = w233 & b_24;
assign w28344 = w3364 & w34183;
assign w28345 = w980 & b_15;
assign w28346 = w3376 & w34184;
assign w28347 = w2152 & b_6;
assign w28348 = ~w307 & w2161;
assign w28349 = (a_26 & ~w3423) | (a_26 & w34185) | (~w3423 & w34185);
assign w28350 = ~w28349 & a_26;
assign w28351 = ~w3215 & ~w3213;
assign w28352 = ~w3433 & w3435;
assign w28353 = w3433 & ~w3435;
assign w28354 = w1688 & b_9;
assign w28355 = w3442 & w34186;
assign w28356 = ~w25016 & ~w3449;
assign w28357 = w1289 & b_12;
assign w28358 = w3458 & w34187;
assign w28359 = ~w3454 & w3464;
assign w28360 = w3454 & ~w3464;
assign w28361 = w651 & b_18;
assign w28362 = w3482 & w34188;
assign w28363 = ~w25017 & ~w3489;
assign w28364 = w412 & b_21;
assign w28365 = (a_11 & ~w3497) | (a_11 & w34189) | (~w3497 & w34189);
assign w28366 = a_11 & ~w25018;
assign w28367 = a_11 & ~w28365;
assign w28368 = w25018 & a_11;
assign w28369 = ~w3309 & w3313;
assign w28370 = w93 & b_27;
assign w28371 = w3521 & w34190;
assign w28372 = ~w3528 & ~w3529;
assign w28373 = ~w3528 & w25019;
assign w28374 = a_0 & b_32;
assign w28375 = w27010 & b_30;
assign w28376 = ~w3341 & ~w28339;
assign w28377 = (~w28337 & w34192) | (~w28337 & w34193) | (w34192 & w34193);
assign w28378 = (w3542 & w28339) | (w3542 & w34192) | (w28339 & w34192);
assign w28379 = (w28337 & w34194) | (w28337 & w34195) | (w34194 & w34195);
assign w28380 = ~w3542 & w28376;
assign w28381 = w3538 & w34196;
assign w28382 = w3553 & ~w3557;
assign w28383 = w233 & b_25;
assign w28384 = w3562 & w34197;
assign w28385 = w1289 & b_13;
assign w28386 = w3575 & w34198;
assign w28387 = w2633 & b_4;
assign w28388 = w3586 & w34199;
assign w28389 = w2152 & b_7;
assign w28390 = w3624 & w34200;
assign w28391 = w1688 & b_10;
assign w28392 = (a_23 & ~w3640) | (a_23 & w34201) | (~w3640 & w34201);
assign w28393 = a_23 & ~w25022;
assign w28394 = w980 & b_16;
assign w28395 = w3663 & w34202;
assign w28396 = w651 & b_19;
assign w28397 = w3679 & w34203;
assign w28398 = w412 & b_22;
assign w28399 = (a_11 & ~w3696) | (a_11 & w34204) | (~w3696 & w34204);
assign w28400 = a_11 & ~w25023;
assign w28401 = a_11 & ~w28399;
assign w28402 = w25023 & a_11;
assign w28403 = w93 & b_28;
assign w28404 = w3720 & w34205;
assign w28405 = a_0 & b_33;
assign w28406 = w27010 & b_31;
assign w28407 = ~w3541 & ~w28377;
assign w28408 = (~w28339 & w34206) | (~w28339 & w34207) | (w34206 & w34207);
assign w28409 = w3737 & w34208;
assign w28410 = ~w3752 & ~w3750;
assign w28411 = w2152 & b_8;
assign w28412 = w3763 & w34209;
assign w28413 = w2633 & b_5;
assign w28414 = w3774 & w34210;
assign w28415 = w3204 & w3596;
assign w28416 = w3610 & ~w3781;
assign w28417 = ~b_0 & a_35;
assign w28418 = w1688 & b_11;
assign w28419 = w3838 & w34211;
assign w28420 = w1289 & b_14;
assign w28421 = w3855 & w34212;
assign w28422 = w980 & b_17;
assign w28423 = (a_17 & ~w3873) | (a_17 & w34213) | (~w3873 & w34213);
assign w28424 = a_17 & ~w25025;
assign w28425 = a_17 & ~w28423;
assign w28426 = w25025 & a_17;
assign w28427 = ~w3882 & w3884;
assign w28428 = w3882 & ~w3884;
assign w28429 = w651 & b_20;
assign w28430 = (a_14 & ~w3891) | (a_14 & w34214) | (~w3891 & w34214);
assign w28431 = a_14 & ~w25027;
assign w28432 = a_14 & ~w28430;
assign w28433 = w25027 & a_14;
assign w28434 = w412 & b_23;
assign w28435 = (a_11 & ~w3909) | (a_11 & w34215) | (~w3909 & w34215);
assign w28436 = a_11 & ~w25029;
assign w28437 = a_11 & ~w28435;
assign w28438 = w25029 & a_11;
assign w28439 = w233 & b_26;
assign w28440 = (a_8 & ~w3926) | (a_8 & w34216) | (~w3926 & w34216);
assign w28441 = a_8 & ~w25031;
assign w28442 = a_8 & ~w28440;
assign w28443 = w25031 & a_8;
assign w28444 = ~w3710 & w34217;
assign w28445 = w93 & b_29;
assign w28446 = w3943 & w34218;
assign w28447 = ~w3951 & ~w3950;
assign w28448 = a_0 & b_34;
assign w28449 = w27010 & b_32;
assign w28450 = w3964 & w3740;
assign w28451 = w3964 & ~w25033;
assign w28452 = ~w3964 & ~w3740;
assign w28453 = ~w3964 & w25033;
assign w28454 = w3960 & w34219;
assign w28455 = w3956 & w3972;
assign w28456 = ~w3956 & ~w3972;
assign w28457 = w3956 & ~w3972;
assign w28458 = w233 & b_27;
assign w28459 = (a_8 & ~w3984) | (a_8 & w34220) | (~w3984 & w34220);
assign w28460 = a_8 & ~w25034;
assign w28461 = a_8 & ~w28459;
assign w28462 = w25034 & a_8;
assign w28463 = w412 & b_24;
assign w28464 = w3994 & w34221;
assign w28465 = w1289 & b_15;
assign w28466 = w4006 & w34222;
assign w28467 = w2152 & b_9;
assign w28468 = w4017 & w34223;
assign w28469 = ~w3823 & ~w3822;
assign w28470 = w2633 & b_6;
assign w28471 = ~w307 & w2642;
assign w28472 = (a_29 & ~w4062) | (a_29 & w34224) | (~w4062 & w34224);
assign w28473 = ~w28472 & a_29;
assign w28474 = w4072 & ~w4024;
assign w28475 = ~w4072 & w4024;
assign w28476 = w1688 & b_12;
assign w28477 = w4086 & w34225;
assign w28478 = w980 & b_18;
assign w28479 = w4110 & w34226;
assign w28480 = w651 & b_21;
assign w28481 = w4127 & w34227;
assign w28482 = w93 & b_30;
assign w28483 = w4157 & w34228;
assign w28484 = ~w4165 & w3950;
assign w28485 = ~w4165 & ~w4164;
assign w28486 = a_0 & b_35;
assign w28487 = w27010 & b_33;
assign w28488 = (~w3963 & ~w3964) | (~w3963 & w34229) | (~w3964 & w34229);
assign w28489 = (~w3963 & w25033) | (~w3963 & w34230) | (w25033 & w34230);
assign w28490 = w4178 & ~w28488;
assign w28491 = w4178 & ~w28489;
assign w28492 = ~w4178 & w28488;
assign w28493 = ~w4178 & w28489;
assign w28494 = w4174 & w34231;
assign w28495 = w4170 & w4186;
assign w28496 = ~w4170 & ~w4186;
assign w28497 = w93 & b_31;
assign w28498 = w4196 & w34232;
assign w28499 = w412 & b_25;
assign w28500 = w4208 & w34233;
assign w28501 = w4001 & ~w4135;
assign w28502 = ~w4100 & w34234;
assign w28503 = w1688 & b_13;
assign w28504 = w4221 & w34235;
assign w28505 = w3189 & b_4;
assign w28506 = w4232 & w34236;
assign w28507 = w2633 & b_7;
assign w28508 = w4270 & w34237;
assign w28509 = w2152 & b_10;
assign w28510 = w4286 & w34238;
assign w28511 = w1289 & b_16;
assign w28512 = w4310 & w34239;
assign w28513 = w980 & b_19;
assign w28514 = w4326 & w34240;
assign w28515 = w651 & b_22;
assign w28516 = w4343 & w34241;
assign w28517 = w233 & b_28;
assign w28518 = w4366 & w34242;
assign w28519 = a_0 & b_36;
assign w28520 = w27010 & b_34;
assign w28521 = (~w4177 & w28488) | (~w4177 & w34243) | (w28488 & w34243);
assign w28522 = w4392 & ~w28521;
assign w28523 = (~w28489 & w34244) | (~w28489 & w34245) | (w34244 & w34245);
assign w28524 = ~w4392 & w28521;
assign w28525 = (w28489 & w34246) | (w28489 & w34247) | (w34246 & w34247);
assign w28526 = ~w12 & w4389;
assign w28527 = w4170 & ~w4186;
assign w28528 = ~w4402 & w34248;
assign w28529 = w93 & b_32;
assign w28530 = w4414 & w34249;
assign w28531 = w233 & b_29;
assign w28532 = w4425 & w34250;
assign w28533 = w1688 & b_14;
assign w28534 = w4437 & w34251;
assign w28535 = w2152 & b_11;
assign w28536 = w4448 & w34252;
assign w28537 = w2633 & b_8;
assign w28538 = w4459 & w34253;
assign w28539 = w3189 & b_5;
assign w28540 = w4470 & w34254;
assign w28541 = w3812 & w4242;
assign w28542 = w4256 & ~w4477;
assign w28543 = ~b_0 & a_38;
assign w28544 = w1289 & b_17;
assign w28545 = w4546 & w34255;
assign w28546 = w980 & b_20;
assign w28547 = w4564 & w34256;
assign w28548 = w651 & b_23;
assign w28549 = w4582 & w34257;
assign w28550 = ~w4590 & w4433;
assign w28551 = w412 & b_26;
assign w28552 = w4599 & w34258;
assign w28553 = ~w4381 & ~w4379;
assign w28554 = a_0 & b_37;
assign w28555 = w27010 & b_35;
assign w28556 = ~w4391 & ~w28523;
assign w28557 = (~w28521 & w34260) | (~w28521 & w34261) | (w34260 & w34261);
assign w28558 = (w4633 & w28523) | (w4633 & w34260) | (w28523 & w34260);
assign w28559 = (w28521 & w34262) | (w28521 & w34263) | (w34262 & w34263);
assign w28560 = ~w4633 & w28556;
assign w28561 = w4629 & w34264;
assign w28562 = a_0 & b_38;
assign w28563 = w27010 & b_36;
assign w28564 = (~w28523 & w34265) | (~w28523 & w34266) | (w34265 & w34266);
assign w28565 = (w4655 & w28557) | (w4655 & w34267) | (w28557 & w34267);
assign w28566 = (w28523 & w34268) | (w28523 & w34269) | (w34268 & w34269);
assign w28567 = ~w28557 & w34270;
assign w28568 = ~w4655 & w28564;
assign w28569 = w4651 & w34271;
assign w28570 = w4622 & ~w4618;
assign w28571 = w93 & b_33;
assign w28572 = w4668 & w34272;
assign w28573 = w233 & b_30;
assign w28574 = w4679 & w34273;
assign w28575 = ~w4608 & ~w4607;
assign w28576 = w412 & b_27;
assign w28577 = w4690 & w34274;
assign w28578 = w1688 & b_15;
assign w28579 = w4701 & w34275;
assign w28580 = w2633 & b_9;
assign w28581 = w4713 & w34276;
assign w28582 = ~w4519 & ~w4518;
assign w28583 = w3189 & b_6;
assign w28584 = ~w307 & w3198;
assign w28585 = (a_32 & ~w4758) | (a_32 & w34277) | (~w4758 & w34277);
assign w28586 = ~w28585 & a_32;
assign w28587 = w2152 & b_12;
assign w28588 = w4781 & w34278;
assign w28589 = w1289 & b_18;
assign w28590 = w4805 & w34279;
assign w28591 = w980 & b_21;
assign w28592 = w4823 & w34280;
assign w28593 = w651 & b_24;
assign w28594 = w4839 & w34281;
assign w28595 = ~w4644 & ~w4643;
assign w28596 = a_0 & b_39;
assign w28597 = w27010 & b_37;
assign w28598 = w4654 & w4885;
assign w28599 = ~w4654 & ~w4885;
assign w28600 = w4881 & w34282;
assign w28601 = ~w4860 & ~w4859;
assign w28602 = w233 & b_31;
assign w28603 = (a_8 & ~w4899) | (a_8 & w34283) | (~w4899 & w34283);
assign w28604 = a_8 & ~w25037;
assign w28605 = w4899 & w34284;
assign w28606 = a_8 & w25037;
assign w28607 = w651 & b_25;
assign w28608 = w4911 & w34285;
assign w28609 = ~w4790 & ~w4789;
assign w28610 = w2152 & b_13;
assign w28611 = w4923 & w34286;
assign w28612 = w3797 & b_4;
assign w28613 = w4933 & w34287;
assign w28614 = w3189 & b_7;
assign w28615 = w4973 & w34288;
assign w28616 = w2633 & b_10;
assign w28617 = w4991 & w34289;
assign w28618 = w1688 & b_16;
assign w28619 = w5015 & w34290;
assign w28620 = w1289 & b_19;
assign w28621 = w5031 & w34291;
assign w28622 = w980 & b_22;
assign w28623 = w5049 & w34292;
assign w28624 = w412 & b_28;
assign w28625 = w5072 & w34293;
assign w28626 = w93 & b_34;
assign w28627 = w5095 & w34294;
assign w28628 = ~w5103 & ~w5104;
assign w28629 = ~w5103 & ~w4867;
assign w28630 = w93 & b_35;
assign w28631 = w5121 & w34295;
assign w28632 = w5088 & ~w5085;
assign w28633 = w233 & b_32;
assign w28634 = w5132 & w34296;
assign w28635 = w651 & b_26;
assign w28636 = w5145 & w34297;
assign w28637 = w2152 & b_14;
assign w28638 = w5155 & w34298;
assign w28639 = w3797 & b_5;
assign w28640 = w5167 & w34299;
assign w28641 = w4508 & w4943;
assign w28642 = w4957 & ~w5174;
assign w28643 = ~b_0 & a_41;
assign w28644 = w3189 & b_8;
assign w28645 = w5225 & w34300;
assign w28646 = w2633 & b_11;
assign w28647 = w5242 & w34301;
assign w28648 = w4919 & ~w5005;
assign w28649 = w1688 & b_17;
assign w28650 = w5266 & w34302;
assign w28651 = w1289 & b_20;
assign w28652 = w5284 & w34303;
assign w28653 = w980 & b_23;
assign w28654 = w5302 & w34304;
assign w28655 = w412 & b_29;
assign w28656 = w5327 & w34305;
assign w28657 = a_0 & b_40;
assign w28658 = w27010 & b_38;
assign w28659 = ~w4884 & ~w4885;
assign w28660 = (~w4884 & ~w4885) | (~w4884 & w34306) | (~w4885 & w34306);
assign w28661 = w5360 & ~w28659;
assign w28662 = w5360 & ~w28660;
assign w28663 = ~w5360 & w28659;
assign w28664 = ~w5360 & w28660;
assign w28665 = w5356 & w34307;
assign w28666 = ~w5371 & ~w5369;
assign w28667 = w5117 & ~w5346;
assign w28668 = ~w5341 & w5128;
assign w28669 = w233 & b_33;
assign w28670 = (a_8 & ~w5382) | (a_8 & w34308) | (~w5382 & w34308);
assign w28671 = a_8 & ~w25040;
assign w28672 = w5382 & w34309;
assign w28673 = a_8 & w25040;
assign w28674 = w412 & b_30;
assign w28675 = (a_11 & ~w5393) | (a_11 & w34310) | (~w5393 & w34310);
assign w28676 = a_11 & ~w25041;
assign w28677 = a_11 & ~w28675;
assign w28678 = w25041 & a_11;
assign w28679 = w651 & b_27;
assign w28680 = w5404 & w34311;
assign w28681 = w1688 & b_18;
assign w28682 = w5416 & w34312;
assign w28683 = w5259 & ~w5255;
assign w28684 = w2152 & b_15;
assign w28685 = w5427 & w34313;
assign w28686 = w2633 & b_12;
assign w28687 = w5438 & w34314;
assign w28688 = ~w5215 & w34315;
assign w28689 = w3797 & b_6;
assign w28690 = ~w307 & w3806;
assign w28691 = (a_35 & ~w5449) | (a_35 & w34316) | (~w5449 & w34316);
assign w28692 = ~w28691 & a_35;
assign w28693 = w3189 & b_9;
assign w28694 = w5500 & w34317;
assign w28695 = w1289 & b_21;
assign w28696 = w5536 & w34318;
assign w28697 = ~w5543 & ~w27342;
assign w28698 = ~w5543 & ~w27341;
assign w28699 = ~w27341 & w27342;
assign w28700 = w980 & b_24;
assign w28701 = w5552 & w34319;
assign w28702 = ~w5548 & w5558;
assign w28703 = w5548 & ~w5558;
assign w28704 = w5309 & w5561;
assign w28705 = ~w5309 & ~w5561;
assign w28706 = w5317 & w5567;
assign w28707 = ~w5317 & ~w5567;
assign w28708 = w93 & b_36;
assign w28709 = w5587 & w34320;
assign w28710 = a_0 & b_41;
assign w28711 = w27010 & b_39;
assign w28712 = (~w5359 & w28659) | (~w5359 & w34321) | (w28659 & w34321);
assign w28713 = (~w5359 & w28660) | (~w5359 & w34321) | (w28660 & w34321);
assign w28714 = w5606 & ~w28712;
assign w28715 = w5606 & ~w28713;
assign w28716 = ~w5606 & w28712;
assign w28717 = ~w5606 & w28713;
assign w28718 = w5602 & w34322;
assign w28719 = w5597 & w5614;
assign w28720 = ~w5597 & ~w5614;
assign w28721 = ~w5594 & ~w5596;
assign w28722 = ~w5594 & ~w5376;
assign w28723 = w93 & b_37;
assign w28724 = w5625 & w34323;
assign w28725 = w5378 & ~w5577;
assign w28726 = w412 & b_31;
assign w28727 = (a_11 & ~w5637) | (a_11 & w34324) | (~w5637 & w34324);
assign w28728 = a_11 & ~w25044;
assign w28729 = a_11 & ~w28727;
assign w28730 = w25044 & a_11;
assign w28731 = w980 & b_25;
assign w28732 = w5649 & w34325;
assign w28733 = w1688 & b_19;
assign w28734 = w5659 & w34326;
assign w28735 = ~w5509 & ~w5508;
assign w28736 = w3189 & b_10;
assign w28737 = w5672 & w34327;
assign w28738 = w4493 & b_4;
assign w28739 = w5683 & w34328;
assign w28740 = w3797 & b_7;
assign w28741 = w5722 & w34329;
assign w28742 = w2633 & b_13;
assign w28743 = w5746 & w34330;
assign w28744 = w2152 & b_16;
assign w28745 = w5763 & w34331;
assign w28746 = w1289 & b_22;
assign w28747 = w5787 & w34332;
assign w28748 = w651 & b_28;
assign w28749 = w5810 & w34333;
assign w28750 = w233 & b_34;
assign w28751 = (a_8 & ~w5833) | (a_8 & w34334) | (~w5833 & w34334);
assign w28752 = a_8 & ~w25045;
assign w28753 = a_8 & ~w28751;
assign w28754 = w25045 & a_8;
assign w28755 = a_0 & b_42;
assign w28756 = w27010 & b_40;
assign w28757 = (~w5605 & w28713) | (~w5605 & w34335) | (w28713 & w34335);
assign w28758 = (~w28712 & w34336) | (~w28712 & w34337) | (w34336 & w34337);
assign w28759 = (~w28713 & w34336) | (~w28713 & w34337) | (w34336 & w34337);
assign w28760 = (w28712 & w34338) | (w28712 & w34339) | (w34338 & w34339);
assign w28761 = ~w5861 & w28757;
assign w28762 = w5857 & w34340;
assign w28763 = a_0 & b_43;
assign w28764 = w27010 & b_41;
assign w28765 = ~w5860 & ~w28759;
assign w28766 = (w5885 & w28758) | (w5885 & w34341) | (w28758 & w34341);
assign w28767 = (w5885 & w28759) | (w5885 & w34341) | (w28759 & w34341);
assign w28768 = ~w28758 & w34342;
assign w28769 = ~w5885 & w28765;
assign w28770 = w5881 & w34343;
assign w28771 = w412 & b_32;
assign w28772 = w5899 & w34344;
assign w28773 = ~w5801 & w34345;
assign w28774 = w980 & b_26;
assign w28775 = w5911 & w34346;
assign w28776 = w2633 & b_14;
assign w28777 = w5921 & w34347;
assign w28778 = w4493 & b_5;
assign w28779 = w5933 & w34348;
assign w28780 = w5205 & w5693;
assign w28781 = w5707 & ~w5940;
assign w28782 = ~b_0 & a_44;
assign w28783 = w3797 & b_8;
assign w28784 = w5991 & w34349;
assign w28785 = w3189 & b_11;
assign w28786 = w6008 & w34350;
assign w28787 = w2152 & b_17;
assign w28788 = w6032 & w34351;
assign w28789 = w1688 & b_20;
assign w28790 = w6050 & w34352;
assign w28791 = w1289 & b_23;
assign w28792 = w6068 & w34353;
assign w28793 = w651 & b_29;
assign w28794 = w6092 & w34354;
assign w28795 = w233 & b_35;
assign w28796 = w6117 & w34355;
assign w28797 = ~w6125 & ~w6124;
assign w28798 = w93 & b_38;
assign w28799 = w6134 & w34356;
assign w28800 = w5874 & ~w5870;
assign w28801 = w93 & b_39;
assign w28802 = w6160 & w34357;
assign w28803 = w412 & b_33;
assign w28804 = w6170 & w34358;
assign w28805 = w651 & b_30;
assign w28806 = w6181 & w34359;
assign w28807 = w980 & b_27;
assign w28808 = w6192 & w34360;
assign w28809 = w2152 & b_18;
assign w28810 = w6204 & w34361;
assign w28811 = w2633 & b_15;
assign w28812 = w6214 & w34362;
assign w28813 = w3189 & b_12;
assign w28814 = w6225 & w34363;
assign w28815 = ~w5981 & w34364;
assign w28816 = w4493 & b_6;
assign w28817 = ~w307 & w4502;
assign w28818 = (a_38 & ~w6236) | (a_38 & w34365) | (~w6236 & w34365);
assign w28819 = ~w28818 & a_38;
assign w28820 = w3797 & b_9;
assign w28821 = w6287 & w34366;
assign w28822 = w1688 & b_21;
assign w28823 = w6323 & w34367;
assign w28824 = w1289 & b_24;
assign w28825 = w6340 & w34368;
assign w28826 = w233 & b_36;
assign w28827 = (a_8 & ~w6376) | (a_8 & w34369) | (~w6376 & w34369);
assign w28828 = a_8 & ~w25047;
assign w28829 = a_8 & ~w28827;
assign w28830 = w25047 & a_8;
assign w28831 = a_0 & b_44;
assign w28832 = w27010 & b_42;
assign w28833 = (~w28759 & w34370) | (~w28759 & w34371) | (w34370 & w34371);
assign w28834 = (w28758 & w34372) | (w28758 & w34373) | (w34372 & w34373);
assign w28835 = (w28759 & w34372) | (w28759 & w34373) | (w34372 & w34373);
assign w28836 = (~w28758 & w34374) | (~w28758 & w34375) | (w34374 & w34375);
assign w28837 = ~w6405 & w28833;
assign w28838 = w6401 & w34376;
assign w28839 = ~w6361 & ~w6360;
assign w28840 = w651 & b_31;
assign w28841 = w6427 & w34377;
assign w28842 = w6199 & ~w6348;
assign w28843 = w1289 & b_25;
assign w28844 = w6439 & w34378;
assign w28845 = w2152 & b_19;
assign w28846 = w6449 & w34379;
assign w28847 = ~w6307 & ~w6308;
assign w28848 = ~w6307 & ~w6027;
assign w28849 = ~w6296 & ~w6295;
assign w28850 = w3797 & b_10;
assign w28851 = w6462 & w34380;
assign w28852 = w5190 & b_4;
assign w28853 = w6473 & w34381;
assign w28854 = w4493 & b_7;
assign w28855 = w6512 & w34382;
assign w28856 = w3189 & b_13;
assign w28857 = w6536 & w34383;
assign w28858 = w2633 & b_16;
assign w28859 = w6553 & w34384;
assign w28860 = w1688 & b_22;
assign w28861 = w6577 & w34385;
assign w28862 = w980 & b_28;
assign w28863 = w6600 & w34386;
assign w28864 = w412 & b_34;
assign w28865 = w6623 & w34387;
assign w28866 = w233 & b_37;
assign w28867 = (a_8 & ~w6639) | (a_8 & w34388) | (~w6639 & w34388);
assign w28868 = a_8 & ~w25048;
assign w28869 = w6639 & w34389;
assign w28870 = a_8 & w25048;
assign w28871 = w93 & b_40;
assign w28872 = w6657 & w34390;
assign w28873 = a_0 & b_45;
assign w28874 = w27010 & b_43;
assign w28875 = w6404 & w6679;
assign w28876 = ~w6404 & ~w6679;
assign w28877 = w6675 & w34391;
assign w28878 = w651 & b_32;
assign w28879 = w6698 & w34392;
assign w28880 = ~w6609 & ~w6607;
assign w28881 = w1289 & b_26;
assign w28882 = w6710 & w34393;
assign w28883 = w3189 & b_14;
assign w28884 = w6720 & w34394;
assign w28885 = w5190 & b_5;
assign w28886 = w6732 & w34395;
assign w28887 = w5971 & w6483;
assign w28888 = w6497 & ~w6739;
assign w28889 = ~b_0 & a_47;
assign w28890 = w4493 & b_8;
assign w28891 = w6790 & w34396;
assign w28892 = w3797 & b_11;
assign w28893 = w6807 & w34397;
assign w28894 = w2633 & b_17;
assign w28895 = w6831 & w34398;
assign w28896 = w2152 & b_20;
assign w28897 = w6849 & w34399;
assign w28898 = ~w6567 & w34400;
assign w28899 = w1688 & b_23;
assign w28900 = w6867 & w34401;
assign w28901 = w980 & b_29;
assign w28902 = w6891 & w34402;
assign w28903 = w6423 & ~w6613;
assign w28904 = w412 & b_35;
assign w28905 = w6915 & w34403;
assign w28906 = w233 & b_38;
assign w28907 = w6933 & w34404;
assign w28908 = w6646 & w25052;
assign w28909 = w93 & b_41;
assign w28910 = w6949 & w34405;
assign w28911 = a_0 & b_46;
assign w28912 = w27010 & b_44;
assign w28913 = ~w6678 & ~w6679;
assign w28914 = (~w6678 & ~w6679) | (~w6678 & w34406) | (~w6679 & w34406);
assign w28915 = w6971 & ~w28913;
assign w28916 = w6971 & ~w28914;
assign w28917 = ~w6971 & w28913;
assign w28918 = ~w6971 & w28914;
assign w28919 = w6967 & w34407;
assign w28920 = ~w6689 & ~w6690;
assign w28921 = ~w6689 & ~w6417;
assign w28922 = a_0 & b_47;
assign w28923 = w27010 & b_45;
assign w28924 = (~w6970 & w28913) | (~w6970 & w34408) | (w28913 & w34408);
assign w28925 = (~w6970 & w28914) | (~w6970 & w34408) | (w28914 & w34408);
assign w28926 = w6995 & ~w28924;
assign w28927 = w6995 & ~w28925;
assign w28928 = ~w6995 & w28924;
assign w28929 = ~w6995 & w28925;
assign w28930 = w6991 & w34409;
assign w28931 = w651 & b_33;
assign w28932 = w7008 & w34410;
assign w28933 = w980 & b_30;
assign w28934 = w7019 & w34411;
assign w28935 = w1289 & b_27;
assign w28936 = w7030 & w34412;
assign w28937 = w3189 & b_15;
assign w28938 = w7043 & w34413;
assign w28939 = w3797 & b_12;
assign w28940 = w7054 & w34414;
assign w28941 = ~w6780 & w34415;
assign w28942 = w5190 & b_6;
assign w28943 = ~w307 & w5199;
assign w28944 = (a_41 & ~w7065) | (a_41 & w34416) | (~w7065 & w34416);
assign w28945 = ~w28944 & a_41;
assign w28946 = w4493 & b_9;
assign w28947 = w7116 & w34417;
assign w28948 = w2633 & b_18;
assign w28949 = w7146 & w34418;
assign w28950 = ~w7140 & ~w7152;
assign w28951 = w2152 & b_21;
assign w28952 = w7164 & w34419;
assign w28953 = ~w7172 & w7038;
assign w28954 = w1688 & b_24;
assign w28955 = w7181 & w34420;
assign w28956 = w412 & b_36;
assign w28957 = (a_11 & ~w7217) | (a_11 & w34421) | (~w7217 & w34421);
assign w28958 = a_11 & ~w25057;
assign w28959 = a_11 & ~w28957;
assign w28960 = w25057 & a_11;
assign w28961 = w233 & b_39;
assign w28962 = w7235 & w34422;
assign w28963 = ~w25058 & ~w7242;
assign w28964 = w93 & b_42;
assign w28965 = w7252 & w34423;
assign w28966 = ~w6980 & w6984;
assign w28967 = w7269 & ~w7265;
assign w28968 = a_0 & b_48;
assign w28969 = w27010 & b_46;
assign w28970 = (~w6994 & w25060) | (~w6994 & w28924) | (w25060 & w28924);
assign w28971 = (~w6994 & w25060) | (~w6994 & w28925) | (w25060 & w28925);
assign w28972 = (~w28924 & w34424) | (~w28924 & w34425) | (w34424 & w34425);
assign w28973 = (~w28925 & w34424) | (~w28925 & w34425) | (w34424 & w34425);
assign w28974 = (w28924 & w34426) | (w28924 & w34427) | (w34426 & w34427);
assign w28975 = (w28925 & w34426) | (w28925 & w34427) | (w34426 & w34427);
assign w28976 = w7277 & w34428;
assign w28977 = ~w7260 & ~w7261;
assign w28978 = ~w7260 & ~w6962;
assign w28979 = w980 & b_31;
assign w28980 = w7295 & w34429;
assign w28981 = w1688 & b_25;
assign w28982 = w7306 & w34430;
assign w28983 = w3797 & b_13;
assign w28984 = w7317 & w34431;
assign w28985 = ~w7125 & ~w7124;
assign w28986 = w4493 & b_10;
assign w28987 = w7328 & w34432;
assign w28988 = w5956 & b_4;
assign w28989 = w7339 & w34433;
assign w28990 = w5190 & b_7;
assign w28991 = w7378 & w34434;
assign w28992 = w7129 & w7400;
assign w28993 = ~w7129 & ~w7400;
assign w28994 = w3189 & b_16;
assign w28995 = w7407 & w34435;
assign w28996 = w2633 & b_19;
assign w28997 = w7425 & w34436;
assign w28998 = w2152 & b_22;
assign w28999 = w7443 & w34437;
assign w29000 = w1289 & b_28;
assign w29001 = w7466 & w34438;
assign w29002 = w651 & b_34;
assign w29003 = (a_14 & ~w7489) | (a_14 & w34439) | (~w7489 & w34439);
assign w29004 = a_14 & ~w26564;
assign w29005 = a_14 & ~w29003;
assign w29006 = w26564 & a_14;
assign w29007 = w412 & b_37;
assign w29008 = a_11 & ~w26565;
assign w29009 = w25065 & a_11;
assign w29010 = w233 & b_40;
assign w29011 = (a_8 & ~w7523) | (a_8 & w34440) | (~w7523 & w34440);
assign w29012 = a_8 & ~w25066;
assign w29013 = a_8 & ~w29011;
assign w29014 = w25066 & a_8;
assign w29015 = w93 & b_43;
assign w29016 = w7540 & w34441;
assign w29017 = w7290 & w34442;
assign w29018 = (~w7289 & ~w7290) | (~w7289 & w34443) | (~w7290 & w34443);
assign w29019 = w1688 & b_26;
assign w29020 = w7562 & w34444;
assign w29021 = w3797 & b_14;
assign w29022 = w7572 & w34445;
assign w29023 = w5956 & b_5;
assign w29024 = w7584 & w34446;
assign w29025 = w6770 & w7349;
assign w29026 = w7363 & ~w7591;
assign w29027 = ~b_0 & a_50;
assign w29028 = w5190 & b_8;
assign w29029 = w7642 & w34447;
assign w29030 = w4493 & b_11;
assign w29031 = w7659 & w34448;
assign w29032 = w3189 & b_17;
assign w29033 = w7683 & w34449;
assign w29034 = w2633 & b_20;
assign w29035 = w7701 & w34450;
assign w29036 = w2152 & b_23;
assign w29037 = w7719 & w34451;
assign w29038 = w1289 & b_29;
assign w29039 = w7744 & w34452;
assign w29040 = ~w7738 & ~w7750;
assign w29041 = w980 & b_32;
assign w29042 = w7762 & w34453;
assign w29043 = w651 & b_35;
assign w29044 = (a_14 & ~w7780) | (a_14 & w34454) | (~w7780 & w34454);
assign w29045 = a_14 & ~w26576;
assign w29046 = a_14 & ~w29044;
assign w29047 = w26576 & a_14;
assign w29048 = ~w7496 & ~w7498;
assign w29049 = ~w7496 & ~w7212;
assign w29050 = w412 & b_38;
assign w29051 = a_11 & ~w26577;
assign w29052 = w25067 & a_11;
assign w29053 = w233 & b_41;
assign w29054 = (a_8 & ~w7816) | (a_8 & w34455) | (~w7816 & w34455);
assign w29055 = a_8 & ~w25069;
assign w29056 = a_8 & ~w29054;
assign w29057 = w25069 & a_8;
assign w29058 = ~w7530 & w7246;
assign w29059 = w93 & b_44;
assign w29060 = w7834 & w34456;
assign w29061 = ~w7828 & ~w7840;
assign w29062 = a_0 & b_49;
assign w29063 = w27010 & b_47;
assign w29064 = (w28924 & w34457) | (w28924 & w34458) | (w34457 & w34458);
assign w29065 = (w28925 & w34457) | (w28925 & w34458) | (w34457 & w34458);
assign w29066 = w7856 & ~w29064;
assign w29067 = w7856 & ~w29065;
assign w29068 = ~w7856 & w29064;
assign w29069 = ~w7856 & w29065;
assign w29070 = w7852 & w34459;
assign w29071 = w980 & b_33;
assign w29072 = w7875 & w34460;
assign w29073 = w1289 & b_30;
assign w29074 = w7886 & w34461;
assign w29075 = w1688 & b_27;
assign w29076 = w7897 & w34462;
assign w29077 = w3797 & b_15;
assign w29078 = w7910 & w34463;
assign w29079 = w4493 & b_12;
assign w29080 = w7921 & w34464;
assign w29081 = ~w7632 & w34465;
assign w29082 = w5956 & b_6;
assign w29083 = ~w307 & w5965;
assign w29084 = (a_44 & ~w7932) | (a_44 & w34466) | (~w7932 & w34466);
assign w29085 = ~w29084 & a_44;
assign w29086 = w5190 & b_9;
assign w29087 = w7982 & w34467;
assign w29088 = w3189 & b_18;
assign w29089 = w8013 & w34468;
assign w29090 = w2633 & b_21;
assign w29091 = w8031 & w34469;
assign w29092 = w2152 & b_24;
assign w29093 = w8048 & w34470;
assign w29094 = w651 & b_36;
assign w29095 = (a_14 & ~w8084) | (a_14 & w34471) | (~w8084 & w34471);
assign w29096 = a_14 & ~w25380;
assign w29097 = a_14 & ~w29095;
assign w29098 = w25380 & a_14;
assign w29099 = w412 & b_39;
assign w29100 = w8102 & w34472;
assign w29101 = a_11 & w25070;
assign w29102 = w233 & b_42;
assign w29103 = (a_8 & ~w8120) | (a_8 & w34473) | (~w8120 & w34473);
assign w29104 = a_8 & ~w25383;
assign w29105 = a_8 & ~w29103;
assign w29106 = w25383 & a_8;
assign w29107 = w93 & b_45;
assign w29108 = (a_5 & ~w8137) | (a_5 & w34474) | (~w8137 & w34474);
assign w29109 = a_5 & ~w25384;
assign w29110 = a_5 & ~w29108;
assign w29111 = w25384 & a_5;
assign w29112 = a_0 & b_50;
assign w29113 = w27010 & b_48;
assign w29114 = (w26583 & w26582) | (w26583 & w28971) | (w26582 & w28971);
assign w29115 = (~w28970 & w34475) | (~w28970 & w34476) | (w34475 & w34476);
assign w29116 = (~w28971 & w34475) | (~w28971 & w34476) | (w34475 & w34476);
assign w29117 = (w28970 & w34477) | (w28970 & w34478) | (w34477 & w34478);
assign w29118 = ~w8159 & w29114;
assign w29119 = w8155 & w34479;
assign w29120 = a_0 & b_51;
assign w29121 = w27010 & b_49;
assign w29122 = ~w8158 & ~w29116;
assign w29123 = (w8183 & w29115) | (w8183 & w34480) | (w29115 & w34480);
assign w29124 = (w8183 & w29116) | (w8183 & w34480) | (w29116 & w34480);
assign w29125 = ~w29115 & w34481;
assign w29126 = ~w29116 & w34481;
assign w29127 = w8179 & w34482;
assign w29128 = ~w8144 & w8148;
assign w29129 = w233 & b_43;
assign w29130 = a_8 & ~w26584;
assign w29131 = w25389 & a_8;
assign w29132 = w1289 & b_31;
assign w29133 = a_20 & ~w26586;
assign w29134 = w25390 & a_20;
assign w29135 = w2152 & b_25;
assign w29136 = w8219 & w34483;
assign w29137 = w3797 & b_16;
assign w29138 = w8230 & w34484;
assign w29139 = w4493 & b_13;
assign w29140 = w8241 & w34485;
assign w29141 = w5190 & b_10;
assign w29142 = w8252 & w34486;
assign w29143 = w6755 & b_4;
assign w29144 = w8262 & w34487;
assign w29145 = w5956 & b_7;
assign w29146 = w8301 & w34488;
assign w29147 = w3189 & b_19;
assign w29148 = w8336 & w34489;
assign w29149 = w2633 & b_22;
assign w29150 = w8354 & w34490;
assign w29151 = w1688 & b_28;
assign w29152 = w8377 & w34491;
assign w29153 = w980 & b_34;
assign w29154 = (a_17 & ~w8400) | (a_17 & w34492) | (~w8400 & w34492);
assign w29155 = a_17 & ~w25396;
assign w29156 = a_17 & ~w29154;
assign w29157 = w25396 & a_17;
assign w29158 = w651 & b_37;
assign w29159 = a_14 & ~w25397;
assign w29160 = w25077 & a_14;
assign w29161 = w412 & b_40;
assign w29162 = a_11 & ~w25399;
assign w29163 = w25078 & a_11;
assign w29164 = w93 & b_46;
assign w29165 = w8458 & w34493;
assign w29166 = w8168 & w8473;
assign w29167 = ~w8168 & ~w8473;
assign w29168 = ~w8467 & ~w8466;
assign w29169 = w4493 & b_14;
assign w29170 = w8485 & w34494;
assign w29171 = w6755 & b_5;
assign w29172 = w8497 & w34495;
assign w29173 = ~b_0 & a_53;
assign w29174 = w5956 & b_8;
assign w29175 = w8555 & w34496;
assign w29176 = w5190 & b_11;
assign w29177 = w8571 & w34497;
assign w29178 = w3797 & b_17;
assign w29179 = w8595 & w34498;
assign w29180 = w3189 & b_20;
assign w29181 = w8612 & w34499;
assign w29182 = w2633 & b_23;
assign w29183 = w8630 & w34500;
assign w29184 = w2152 & b_26;
assign w29185 = w8647 & w34501;
assign w29186 = w1688 & b_29;
assign w29187 = (a_23 & ~w8663) | (a_23 & w34502) | (~w8663 & w34502);
assign w29188 = a_23 & ~w26592;
assign w29189 = a_23 & ~w29187;
assign w29190 = w26592 & a_23;
assign w29191 = w1289 & b_32;
assign w29192 = (a_20 & ~w8681) | (a_20 & w34503) | (~w8681 & w34503);
assign w29193 = a_20 & ~w26593;
assign w29194 = a_20 & ~w29192;
assign w29195 = w26593 & a_20;
assign w29196 = w980 & b_35;
assign w29197 = a_17 & ~w26594;
assign w29198 = w25402 & a_17;
assign w29199 = w651 & b_38;
assign w29200 = a_14 & ~w25403;
assign w29201 = w25080 & a_14;
assign w29202 = w412 & b_41;
assign w29203 = a_11 & ~w26596;
assign w29204 = w25405 & a_11;
assign w29205 = w233 & b_44;
assign w29206 = a_8 & ~w26599;
assign w29207 = w25407 & a_8;
assign w29208 = ~w8449 & w34504;
assign w29209 = w93 & b_47;
assign w29210 = w8769 & w34505;
assign w29211 = a_0 & b_52;
assign w29212 = w27010 & b_50;
assign w29213 = (~w29116 & w34506) | (~w29116 & w34507) | (w34506 & w34507);
assign w29214 = (w29115 & w34508) | (w29115 & w34509) | (w34508 & w34509);
assign w29215 = (w29116 & w34508) | (w29116 & w34509) | (w34508 & w34509);
assign w29216 = (~w29115 & w34510) | (~w29115 & w34511) | (w34510 & w34511);
assign w29217 = ~w8790 & w29213;
assign w29218 = w8786 & w34512;
assign w29219 = ~w8471 & ~w8801;
assign w29220 = ~w8777 & w34513;
assign w29221 = w1289 & b_33;
assign w29222 = (a_20 & ~w8810) | (a_20 & w34514) | (~w8810 & w34514);
assign w29223 = a_20 & ~w26601;
assign w29224 = a_20 & ~w29222;
assign w29225 = w26601 & a_20;
assign w29226 = w1688 & b_30;
assign w29227 = (a_23 & ~w8821) | (a_23 & w34515) | (~w8821 & w34515);
assign w29228 = a_23 & ~w26602;
assign w29229 = a_23 & ~w29227;
assign w29230 = w26602 & a_23;
assign w29231 = w2152 & b_27;
assign w29232 = w8832 & w34516;
assign w29233 = w3189 & b_21;
assign w29234 = w8844 & w34517;
assign w29235 = w4493 & b_15;
assign w29236 = w8855 & w34518;
assign w29237 = w5190 & b_12;
assign w29238 = w8866 & w34519;
assign w29239 = w5956 & b_9;
assign w29240 = w8876 & w34520;
assign w29241 = w6755 & b_6;
assign w29242 = ~w307 & w6764;
assign w29243 = (a_47 & ~w8920) | (a_47 & w34521) | (~w8920 & w34521);
assign w29244 = ~w29243 & a_47;
assign w29245 = w3797 & b_18;
assign w29246 = w8958 & w34522;
assign w29247 = w2633 & b_24;
assign w29248 = w8981 & w34523;
assign w29249 = w980 & b_36;
assign w29250 = a_17 & ~w25561;
assign w29251 = w25409 & a_17;
assign w29252 = w651 & b_39;
assign w29253 = w412 & b_42;
assign w29254 = w9054 & a_11;
assign w29255 = w25413 & a_11;
assign w29256 = w233 & b_45;
assign w29257 = a_8 & ~w26609;
assign w29258 = w25414 & a_8;
assign w29259 = w93 & b_48;
assign w29260 = w9088 & w34524;
assign w29261 = ~w8806 & ~w26813;
assign w29262 = ~w9095 & w8477;
assign w29263 = (~w9095 & ~w27006) | (~w9095 & w34525) | (~w27006 & w34525);
assign w29264 = a_0 & b_53;
assign w29265 = w27010 & b_51;
assign w29266 = (w26815 & w26814) | (w26815 & w29122) | (w26814 & w29122);
assign w29267 = (w29115 & w34528) | (w29115 & w34529) | (w34528 & w34529);
assign w29268 = (~w29122 & w34530) | (~w29122 & w34531) | (w34530 & w34531);
assign w29269 = (~w29115 & w34532) | (~w29115 & w34533) | (w34532 & w34533);
assign w29270 = ~w9107 & w29266;
assign w29271 = w9103 & w34534;
assign w29272 = (w29261 & w34535) | (w29261 & w34536) | (w34535 & w34536);
assign w29273 = (~w29261 & w34537) | (~w29261 & w34538) | (w34537 & w34538);
assign w29274 = (w29261 & w34539) | (w29261 & w34540) | (w34539 & w34540);
assign w29275 = a_0 & b_54;
assign w29276 = w27010 & b_52;
assign w29277 = (w29122 & w34541) | (w29122 & w34542) | (w34541 & w34542);
assign w29278 = (w9131 & w29267) | (w9131 & w34543) | (w29267 & w34543);
assign w29279 = (~w29122 & w34544) | (~w29122 & w34545) | (w34544 & w34545);
assign w29280 = ~w29267 & w34546;
assign w29281 = (w29122 & w34547) | (w29122 & w34548) | (w34547 & w34548);
assign w29282 = w9127 & w34549;
assign w29283 = w412 & b_43;
assign w29284 = w2152 & b_28;
assign w29285 = w9157 & w34550;
assign w29286 = w2633 & b_25;
assign w29287 = w9168 & w34551;
assign w29288 = w3189 & b_22;
assign w29289 = w9178 & w34552;
assign w29290 = w3797 & b_19;
assign w29291 = w9189 & w34553;
assign w29292 = w4493 & b_16;
assign w29293 = (a_38 & ~w9200) | (a_38 & w34554) | (~w9200 & w34554);
assign w29294 = a_38 & ~w25574;
assign w29295 = a_38 & ~w29293;
assign w29296 = w25574 & a_38;
assign w29297 = w5190 & b_13;
assign w29298 = w9211 & w34555;
assign w29299 = w5956 & b_10;
assign w29300 = w9222 & w34556;
assign w29301 = w6755 & b_7;
assign w29302 = w9233 & w34557;
assign w29303 = w7607 & b_4;
assign w29304 = w9243 & w34558;
assign w29305 = w1688 & b_31;
assign w29306 = a_23 & ~w26613;
assign w29307 = w25577 & a_23;
assign w29308 = w1289 & b_34;
assign w29309 = (a_20 & ~w9350) | (a_20 & w34559) | (~w9350 & w34559);
assign w29310 = a_20 & ~w26615;
assign w29311 = a_20 & ~w29309;
assign w29312 = w26615 & a_20;
assign w29313 = w980 & b_37;
assign w29314 = a_17 & ~w25578;
assign w29315 = w25417 & a_17;
assign w29316 = w651 & b_40;
assign w29317 = w233 & b_46;
assign w29318 = (a_8 & ~w9408) | (a_8 & w34560) | (~w9408 & w34560);
assign w29319 = a_8 & ~w26616;
assign w29320 = a_8 & ~w29318;
assign w29321 = w26616 & a_8;
assign w29322 = ~w9077 & w9418;
assign w29323 = w9077 & ~w9418;
assign w29324 = w93 & b_49;
assign w29325 = w9426 & w34561;
assign w29326 = ~w9434 & ~w9435;
assign w29327 = (~w9434 & ~w9435) | (~w9434 & w34562) | (~w9435 & w34562);
assign w29328 = w93 & b_50;
assign w29329 = w9449 & w34563;
assign w29330 = w233 & b_47;
assign w29331 = (a_8 & ~w9459) | (a_8 & w34564) | (~w9459 & w34564);
assign w29332 = a_8 & ~w25420;
assign w29333 = a_8 & ~w29331;
assign w29334 = w25420 & a_8;
assign w29335 = w5190 & b_14;
assign w29336 = w9472 & w34565;
assign w29337 = w5956 & b_11;
assign w29338 = w9483 & w34566;
assign w29339 = w6755 & b_8;
assign w29340 = w9494 & w34567;
assign w29341 = w7607 & b_5;
assign w29342 = w9505 & w34568;
assign w29343 = ~b_0 & a_56;
assign w29344 = w4493 & b_17;
assign w29345 = w9581 & w34569;
assign w29346 = w3797 & b_20;
assign w29347 = w9598 & w34570;
assign w29348 = w3189 & b_23;
assign w29349 = w9616 & w34571;
assign w29350 = w2633 & b_26;
assign w29351 = (a_29 & ~w9634) | (a_29 & w34572) | (~w9634 & w34572);
assign w29352 = a_29 & ~w26618;
assign w29353 = a_29 & ~w29351;
assign w29354 = w26618 & a_29;
assign w29355 = w2152 & b_29;
assign w29356 = (a_26 & ~w9652) | (a_26 & w34573) | (~w9652 & w34573);
assign w29357 = a_26 & ~w26619;
assign w29358 = a_26 & ~w29356;
assign w29359 = w26619 & a_26;
assign w29360 = w1688 & b_32;
assign w29361 = (a_23 & ~w9670) | (a_23 & w34574) | (~w9670 & w34574);
assign w29362 = a_23 & ~w26620;
assign w29363 = a_23 & ~w29361;
assign w29364 = w26620 & a_23;
assign w29365 = w1289 & b_35;
assign w29366 = a_20 & ~w26621;
assign w29367 = w25587 & a_20;
assign w29368 = w980 & b_38;
assign w29369 = w651 & b_41;
assign w29370 = w412 & b_44;
assign w29371 = ~w9754 & ~w9415;
assign w29372 = ~w9754 & w27050;
assign w29373 = a_0 & b_55;
assign w29374 = w27010 & b_53;
assign w29375 = (~w29267 & w34575) | (~w29267 & w34576) | (w34575 & w34576);
assign w29376 = (~w9130 & w25094) | (~w9130 & w29277) | (w25094 & w29277);
assign w29377 = w9768 & w34577;
assign w29378 = ~w9439 & ~w9784;
assign w29379 = a_0 & b_56;
assign w29380 = w27010 & b_54;
assign w29381 = ~w9773 & ~w9772;
assign w29382 = w9795 & w9772;
assign w29383 = w9795 & ~w29381;
assign w29384 = ~w9795 & ~w9772;
assign w29385 = ~w9795 & w29381;
assign w29386 = w9791 & w34578;
assign w29387 = w233 & b_48;
assign w29388 = w9809 & w34579;
assign w29389 = w1688 & b_33;
assign w29390 = a_23 & ~w26627;
assign w29391 = w25595 & a_23;
assign w29392 = w2152 & b_30;
assign w29393 = a_26 & ~w26629;
assign w29394 = w25596 & a_26;
assign w29395 = w5190 & b_15;
assign w29396 = w9844 & w34580;
assign w29397 = w5956 & b_12;
assign w29398 = w9855 & w34581;
assign w29399 = w6755 & b_9;
assign w29400 = w9866 & w34582;
assign w29401 = w7607 & b_6;
assign w29402 = ~w307 & w7616;
assign w29403 = (a_50 & ~w9910) | (a_50 & w34583) | (~w9910 & w34583);
assign w29404 = ~w29403 & a_50;
assign w29405 = w4493 & b_18;
assign w29406 = w9948 & w34584;
assign w29407 = w3797 & b_21;
assign w29408 = w9965 & w34585;
assign w29409 = w3189 & b_24;
assign w29410 = (a_32 & ~w9981) | (a_32 & w34586) | (~w9981 & w34586);
assign w29411 = a_32 & ~w25828;
assign w29412 = a_32 & ~w29410;
assign w29413 = w25828 & a_32;
assign w29414 = w2633 & b_27;
assign w29415 = w9998 & w34587;
assign w29416 = w1289 & b_36;
assign w29417 = a_20 & ~w25831;
assign w29418 = w25598 & a_20;
assign w29419 = w980 & b_39;
assign w29420 = w651 & b_42;
assign w29421 = w412 & b_45;
assign w29422 = w93 & b_51;
assign w29423 = w10104 & w34588;
assign w29424 = w93 & b_52;
assign w29425 = w10129 & w34589;
assign w29426 = w233 & b_49;
assign w29427 = w10140 & w34590;
assign w29428 = w412 & b_46;
assign w29429 = w651 & b_43;
assign w29430 = w2633 & b_28;
assign w29431 = w10175 & w34591;
assign w29432 = w4493 & b_19;
assign w29433 = w10186 & w34592;
assign w29434 = w5190 & b_16;
assign w29435 = (a_41 & ~w10197) | (a_41 & w34593) | (~w10197 & w34593);
assign w29436 = a_41 & ~w25841;
assign w29437 = a_41 & ~w29435;
assign w29438 = w25841 & a_41;
assign w29439 = w5956 & b_13;
assign w29440 = w10208 & w34594;
assign w29441 = w6755 & b_10;
assign w29442 = w10219 & w34595;
assign w29443 = w8520 & b_4;
assign w29444 = w10230 & w34596;
assign w29445 = w7607 & b_7;
assign w29446 = w10268 & w34597;
assign w29447 = w3797 & b_22;
assign w29448 = w10309 & w34598;
assign w29449 = w3189 & b_25;
assign w29450 = w10327 & w34599;
assign w29451 = w2152 & b_31;
assign w29452 = a_26 & ~w25844;
assign w29453 = w25611 & a_26;
assign w29454 = w1688 & b_34;
assign w29455 = (a_23 & ~w10366) | (a_23 & w34600) | (~w10366 & w34600);
assign w29456 = a_23 & ~w25846;
assign w29457 = a_23 & ~w29455;
assign w29458 = w25846 & a_23;
assign w29459 = w1289 & b_37;
assign w29460 = w980 & b_40;
assign w29461 = a_0 & b_57;
assign w29462 = w27010 & b_55;
assign w29463 = w25851 | w25852;
assign w29464 = (w25852 & w25851) | (w25852 & ~w9773) | (w25851 & ~w9773);
assign w29465 = w10449 & ~w29464;
assign w29466 = w10449 & ~w29463;
assign w29467 = ~w10449 & w29464;
assign w29468 = ~w10449 & w29463;
assign w29469 = w10445 & w34601;
assign w29470 = a_0 & b_58;
assign w29471 = w27010 & b_56;
assign w29472 = (~w10448 & w29463) | (~w10448 & w34602) | (w29463 & w34602);
assign w29473 = (~w10448 & w29464) | (~w10448 & w34602) | (w29464 & w34602);
assign w29474 = (~w29464 & w34603) | (~w29464 & w34604) | (w34603 & w34604);
assign w29475 = (~w29463 & w34603) | (~w29463 & w34604) | (w34603 & w34604);
assign w29476 = (w29464 & w34605) | (w29464 & w34606) | (w34605 & w34606);
assign w29477 = (w29463 & w34605) | (w29463 & w34606) | (w34605 & w34606);
assign w29478 = w10469 & w34607;
assign w29479 = w93 & b_53;
assign w29480 = w10485 & w34608;
assign w29481 = w233 & b_50;
assign w29482 = (a_8 & ~w10495) | (a_8 & w34609) | (~w10495 & w34609);
assign w29483 = a_8 & ~w25855;
assign w29484 = a_8 & ~w29482;
assign w29485 = w25855 & a_8;
assign w29486 = w412 & b_47;
assign w29487 = a_11 & ~w25856;
assign w29488 = w25615 & a_11;
assign w29489 = w7607 & b_8;
assign w29490 = w10522 & w34610;
assign w29491 = w8520 & b_5;
assign w29492 = w10533 & w34611;
assign w29493 = ~b_0 & a_59;
assign w29494 = w6755 & b_11;
assign w29495 = w10597 & w34612;
assign w29496 = w5956 & b_14;
assign w29497 = w10614 & w34613;
assign w29498 = w5190 & b_17;
assign w29499 = w10632 & w34614;
assign w29500 = w4493 & b_20;
assign w29501 = w10649 & w34615;
assign w29502 = w3797 & b_23;
assign w29503 = (a_35 & ~w10667) | (a_35 & w34616) | (~w10667 & w34616);
assign w29504 = a_35 & ~w26189;
assign w29505 = a_35 & ~w29503;
assign w29506 = w26189 & a_35;
assign w29507 = w3189 & b_26;
assign w29508 = a_32 & ~w26190;
assign w29509 = w25861 & a_32;
assign w29510 = w2633 & b_29;
assign w29511 = (a_29 & ~w10702) | (a_29 & w34617) | (~w10702 & w34617);
assign w29512 = a_29 & ~w26192;
assign w29513 = a_29 & ~w29511;
assign w29514 = w26192 & a_29;
assign w29515 = w2152 & b_32;
assign w29516 = a_26 & ~w26193;
assign w29517 = w25862 & a_26;
assign w29518 = w1688 & b_35;
assign w29519 = a_23 & ~w25864;
assign w29520 = w25616 & a_23;
assign w29521 = w1289 & b_38;
assign w29522 = w980 & b_41;
assign w29523 = w651 & b_44;
assign w29524 = ~w10427 & ~w10810;
assign w29525 = w10816 & w10434;
assign w29526 = w10816 & ~w10125;
assign w29527 = ~w10816 & ~w10434;
assign w29528 = ~w10816 & w10125;
assign w29529 = w233 & b_51;
assign w29530 = w10834 & w34618;
assign w29531 = w412 & b_48;
assign w29532 = a_11 & ~w26199;
assign w29533 = w25876 & a_11;
assign w29534 = w2152 & b_33;
assign w29535 = a_26 & ~w26201;
assign w29536 = w25877 & a_26;
assign w29537 = w5956 & b_15;
assign w29538 = a_44 & ~w26204;
assign w29539 = w25878 & a_44;
assign w29540 = w6755 & b_12;
assign w29541 = (a_47 & ~w10881) | (a_47 & w34619) | (~w10881 & w34619);
assign w29542 = a_47 & ~w26206;
assign w29543 = a_47 & ~w29541;
assign w29544 = w26206 & a_47;
assign w29545 = w7607 & b_9;
assign w29546 = w10892 & w34620;
assign w29547 = w8520 & b_6;
assign w29548 = ~w307 & w8529;
assign w29549 = (a_53 & ~w10937) | (a_53 & w34621) | (~w10937 & w34621);
assign w29550 = ~w29549 & a_53;
assign w29551 = w5190 & b_18;
assign w29552 = w10975 & w34622;
assign w29553 = w4493 & b_21;
assign w29554 = w10992 & w34623;
assign w29555 = w3797 & b_24;
assign w29556 = (a_35 & ~w11008) | (a_35 & w34624) | (~w11008 & w34624);
assign w29557 = a_35 & ~w26209;
assign w29558 = a_35 & ~w29556;
assign w29559 = w26209 & a_35;
assign w29560 = w3189 & b_27;
assign w29561 = a_32 & ~w26211;
assign w29562 = w25879 & a_32;
assign w29563 = w2633 & b_30;
assign w29564 = (a_29 & ~w11042) | (a_29 & w34625) | (~w11042 & w34625);
assign w29565 = a_29 & ~w26215;
assign w29566 = a_29 & ~w29564;
assign w29567 = w26215 & a_29;
assign w29568 = w1688 & b_36;
assign w29569 = a_23 & ~w25880;
assign w29570 = w25621 & a_23;
assign w29571 = w1289 & b_39;
assign w29572 = w980 & b_42;
assign w29573 = w651 & b_45;
assign w29574 = w93 & b_54;
assign w29575 = w11149 & w34626;
assign w29576 = a_0 & b_59;
assign w29577 = w27010 & b_57;
assign w29578 = (w29463 & w34627) | (w29463 & w34628) | (w34627 & w34628);
assign w29579 = (w29464 & w34627) | (w29464 & w34628) | (w34627 & w34628);
assign w29580 = (w26224 & w26223) | (w26224 & w29466) | (w26223 & w29466);
assign w29581 = (w26224 & w26223) | (w26224 & w29465) | (w26223 & w29465);
assign w29582 = ~w11166 & w29579;
assign w29583 = ~w11166 & w29578;
assign w29584 = w11162 & w34629;
assign w29585 = (~w10820 & w11178) | (~w10820 & w34630) | (w11178 & w34630);
assign w29586 = ~w11180 & w25112;
assign w29587 = ~w11180 & w34631;
assign w29588 = (~w11143 & w34632) | (~w11143 & w34633) | (w34632 & w34633);
assign w29589 = w27010 & b_58;
assign w29590 = ~w11165 & ~w29581;
assign w29591 = (w11193 & w29580) | (w11193 & w34634) | (w29580 & w34634);
assign w29592 = (w11193 & w29581) | (w11193 & w34634) | (w29581 & w34634);
assign w29593 = ~w29580 & w34635;
assign w29594 = ~w11193 & w29590;
assign w29595 = ~w12 & w11190;
assign w29596 = w93 & b_55;
assign w29597 = w11205 & w34636;
assign w29598 = w233 & b_52;
assign w29599 = w11216 & w34637;
assign w29600 = w412 & b_49;
assign w29601 = a_11 & ~w26226;
assign w29602 = w25888 & a_11;
assign w29603 = w651 & b_46;
assign w29604 = w980 & b_43;
assign w29605 = w2633 & b_31;
assign w29606 = w5190 & b_19;
assign w29607 = w11272 & w34638;
assign w29608 = w5956 & b_16;
assign w29609 = a_44 & ~w26234;
assign w29610 = w25895 & a_44;
assign w29611 = w6755 & b_13;
assign w29612 = w11294 & w34639;
assign w29613 = w7607 & b_10;
assign w29614 = w11305 & w34640;
assign w29615 = w9528 & b_4;
assign w29616 = w11316 & w34641;
assign w29617 = w8520 & b_7;
assign w29618 = w11353 & w34642;
assign w29619 = w4493 & b_22;
assign w29620 = (a_38 & ~w11394) | (a_38 & w34643) | (~w11394 & w34643);
assign w29621 = a_38 & ~w26236;
assign w29622 = a_38 & ~w29620;
assign w29623 = w26236 & a_38;
assign w29624 = w3797 & b_25;
assign w29625 = a_35 & ~w26237;
assign w29626 = w25896 & a_35;
assign w29627 = w3189 & b_28;
assign w29628 = (a_32 & ~w11430) | (a_32 & w34644) | (~w11430 & w34644);
assign w29629 = a_32 & ~w26239;
assign w29630 = a_32 & ~w29628;
assign w29631 = w26239 & a_32;
assign w29632 = w2152 & b_34;
assign w29633 = a_26 & ~w26240;
assign w29634 = w25897 & a_26;
assign w29635 = w1688 & b_37;
assign w29636 = a_23 & ~w25898;
assign w29637 = w25630 & a_23;
assign w29638 = w1289 & b_40;
assign w29639 = w233 & b_53;
assign w29640 = w11542 & w34645;
assign w29641 = w412 & b_50;
assign w29642 = (a_11 & ~w11553) | (a_11 & w34646) | (~w11553 & w34646);
assign w29643 = a_11 & ~w26247;
assign w29644 = a_11 & ~w29642;
assign w29645 = w26247 & a_11;
assign w29646 = w651 & b_47;
assign w29647 = w8520 & b_8;
assign w29648 = w11580 & w34647;
assign w29649 = w9528 & b_5;
assign w29650 = w11591 & w34648;
assign w29651 = w10571 & w11326;
assign w29652 = ~b_0 & a_62;
assign w29653 = ~w11627 & ~w11611;
assign w29654 = w7607 & b_11;
assign w29655 = w11655 & w34649;
assign w29656 = w6755 & b_14;
assign w29657 = w11672 & w34650;
assign w29658 = w5956 & b_17;
assign w29659 = w11690 & w34651;
assign w29660 = w5190 & b_20;
assign w29661 = w11706 & w34652;
assign w29662 = w4493 & b_23;
assign w29663 = (a_38 & ~w11724) | (a_38 & w34653) | (~w11724 & w34653);
assign w29664 = a_38 & ~w26250;
assign w29665 = a_38 & ~w29663;
assign w29666 = w26250 & a_38;
assign w29667 = w3797 & b_26;
assign w29668 = a_35 & ~w26251;
assign w29669 = w25903 & a_35;
assign w29670 = w3189 & b_29;
assign w29671 = w2633 & b_32;
assign w29672 = (a_29 & ~w11777) | (a_29 & w34654) | (~w11777 & w34654);
assign w29673 = a_29 & ~w26255;
assign w29674 = a_29 & ~w29672;
assign w29675 = w26255 & a_29;
assign w29676 = w2152 & b_35;
assign w29677 = w1688 & b_38;
assign w29678 = ~w11476 & w11821;
assign w29679 = w11476 & ~w11821;
assign w29680 = w1289 & b_41;
assign w29681 = ~w11836 & ~w26260;
assign w29682 = w980 & b_44;
assign w29683 = w93 & b_56;
assign w29684 = w11881 & w34655;
assign w29685 = a_0 & b_61;
assign w29686 = w27010 & b_59;
assign w29687 = (~w29581 & w34656) | (~w29581 & w34657) | (w34656 & w34657);
assign w29688 = (w29580 & w34658) | (w29580 & w34659) | (w34658 & w34659);
assign w29689 = (w29581 & w34658) | (w29581 & w34659) | (w34658 & w34659);
assign w29690 = (~w29580 & w34660) | (~w29580 & w34661) | (w34660 & w34661);
assign w29691 = ~w11898 & w29687;
assign w29692 = w11894 & w34662;
assign w29693 = (w11201 & ~w11526) | (w11201 & w34663) | (~w11526 & w34663);
assign w29694 = ~w11911 & ~w11912;
assign w29695 = ~w11911 & ~w11536;
assign w29696 = (w11906 & ~w11877) | (w11906 & w34664) | (~w11877 & w34664);
assign w29697 = w651 & b_48;
assign w29698 = a_14 & ~w26265;
assign w29699 = w25912 & a_14;
assign w29700 = w6755 & b_15;
assign w29701 = w11938 & w34665;
assign w29702 = w7607 & b_12;
assign w29703 = w11948 & w34666;
assign w29704 = w8520 & b_9;
assign w29705 = w11959 & w34667;
assign w29706 = w10556 & b_3;
assign w29707 = (a_59 & ~w11986) | (a_59 & w34668) | (~w11986 & w34668);
assign w29708 = w9528 & b_6;
assign w29709 = ~w307 & w9537;
assign w29710 = (a_56 & ~w12004) | (a_56 & w34669) | (~w12004 & w34669);
assign w29711 = ~w29710 & a_56;
assign w29712 = w5956 & b_18;
assign w29713 = w12042 & w34670;
assign w29714 = w5190 & b_21;
assign w29715 = w12058 & w34671;
assign w29716 = w4493 & b_24;
assign w29717 = (a_38 & ~w12074) | (a_38 & w34672) | (~w12074 & w34672);
assign w29718 = a_38 & ~w26267;
assign w29719 = a_38 & ~w29717;
assign w29720 = w26267 & a_38;
assign w29721 = w3797 & b_27;
assign w29722 = a_35 & ~w26268;
assign w29723 = w25913 & a_35;
assign w29724 = w3189 & b_30;
assign w29725 = a_32 & ~w26270;
assign w29726 = w25914 & a_32;
assign w29727 = w2633 & b_33;
assign w29728 = (a_29 & ~w12127) | (a_29 & w34673) | (~w12127 & w34673);
assign w29729 = a_29 & ~w26273;
assign w29730 = a_29 & ~w29728;
assign w29731 = w26273 & a_29;
assign w29732 = w2152 & b_36;
assign w29733 = a_26 & ~w26275;
assign w29734 = w25915 & a_26;
assign w29735 = w1688 & b_39;
assign w29736 = w1289 & b_42;
assign w29737 = w980 & b_45;
assign w29738 = w412 & b_51;
assign w29739 = w12220 & w34674;
assign w29740 = w233 & b_54;
assign w29741 = w12236 & w34675;
assign w29742 = w93 & b_57;
assign w29743 = (w9770 & w34676) | (w9770 & w34677) | (w34676 & w34677);
assign w29744 = w11874 & ~w11870;
assign w29745 = a_0 & b_62;
assign w29746 = w27010 & b_60;
assign w29747 = (~w29581 & w34678) | (~w29581 & w34679) | (w34678 & w34679);
assign w29748 = (w29580 & w34680) | (w29580 & w34681) | (w34680 & w34681);
assign w29749 = (w29581 & w34680) | (w29581 & w34681) | (w34680 & w34681);
assign w29750 = (~w29580 & w34682) | (~w29580 & w34683) | (w34682 & w34683);
assign w29751 = (~w29581 & w34682) | (~w29581 & w34683) | (w34682 & w34683);
assign w29752 = w12266 & w34684;
assign w29753 = w651 & b_49;
assign w29754 = (a_14 & ~w12292) | (a_14 & w34685) | (~w12292 & w34685);
assign w29755 = a_14 & ~w26285;
assign w29756 = a_14 & ~w29754;
assign w29757 = w26285 & a_14;
assign w29758 = w980 & b_46;
assign w29759 = w1289 & b_43;
assign w29760 = w1688 & b_40;
assign w29761 = a_23 & ~w25929;
assign w29762 = w25643 & a_23;
assign w29763 = w3189 & b_31;
assign w29764 = a_32 & ~w25931;
assign w29765 = w25644 & a_32;
assign w29766 = w5956 & b_19;
assign w29767 = w12348 & w34686;
assign w29768 = w7607 & b_13;
assign w29769 = w12359 & w34687;
assign w29770 = w11966 & ~w12013;
assign w29771 = w9528 & b_7;
assign w29772 = w12371 & w34688;
assign w29773 = w10556 & b_4;
assign w29774 = w12404 & w34689;
assign w29775 = w8520 & b_10;
assign w29776 = w12427 & w34690;
assign w29777 = w6755 & b_16;
assign w29778 = w12451 & w34691;
assign w29779 = w5190 & b_22;
assign w29780 = w12473 & w34692;
assign w29781 = w4493 & b_25;
assign w29782 = (a_38 & ~w12491) | (a_38 & w34693) | (~w12491 & w34693);
assign w29783 = a_38 & ~w26289;
assign w29784 = a_38 & ~w29782;
assign w29785 = w26289 & a_38;
assign w29786 = w3797 & b_28;
assign w29787 = a_35 & ~w26290;
assign w29788 = w25933 & a_35;
assign w29789 = w2633 & b_34;
assign w29790 = (a_29 & ~w12533) | (a_29 & w34694) | (~w12533 & w34694);
assign w29791 = a_29 & ~w25934;
assign w29792 = a_29 & ~w29790;
assign w29793 = w25934 & a_29;
assign w29794 = w2152 & b_37;
assign w29795 = ~w12573 & ~w12309;
assign w29796 = w12573 & ~w12309;
assign w29797 = w412 & b_52;
assign w29798 = (a_11 & ~w12592) | (a_11 & w34695) | (~w12592 & w34695);
assign w29799 = a_11 & ~w26294;
assign w29800 = a_11 & ~w29798;
assign w29801 = w26294 & a_11;
assign w29802 = w233 & b_55;
assign w29803 = w12610 & w34696;
assign w29804 = w93 & b_58;
assign w29805 = (a_5 & ~w12622) | (a_5 & w34697) | (~w12622 & w34697);
assign w29806 = a_5 & ~w27554;
assign w29807 = a_5 & ~w29805;
assign w29808 = w27554 & a_5;
assign w29809 = (w12255 & ~w12232) | (w12255 & w34698) | (~w12232 & w34698);
assign w29810 = a_0 & b_63;
assign w29811 = w27010 & b_61;
assign w29812 = (~w29580 & w34699) | (~w29580 & w34700) | (w34699 & w34700);
assign w29813 = (~w29747 & w34701) | (~w29747 & w34702) | (w34701 & w34702);
assign w29814 = (w29580 & w34703) | (w29580 & w34704) | (w34703 & w34704);
assign w29815 = (w29747 & w34705) | (w29747 & w34706) | (w34705 & w34706);
assign w29816 = (~w29580 & w34707) | (~w29580 & w34708) | (w34707 & w34708);
assign w29817 = w12639 & w34709;
assign w29818 = (w12651 & w12631) | (w12651 & w34710) | (w12631 & w34710);
assign w29819 = w27010 & b_62;
assign w29820 = ~b_62 & ~w29814;
assign w29821 = (~w29747 & w34713) | (~w29747 & w34714) | (w34713 & w34714);
assign w29822 = b_63 & ~w29820;
assign w29823 = (~w29747 & w34715) | (~w29747 & w34716) | (w34715 & w34716);
assign w29824 = (~w9770 & w34717) | (~w9770 & w34718) | (w34717 & w34718);
assign w29825 = (a_2 & w12667) | (a_2 & w34719) | (w12667 & w34719);
assign w29826 = ~w29825 & a_2;
assign w29827 = w412 & b_53;
assign w29828 = w12684 & w34720;
assign w29829 = w651 & b_50;
assign w29830 = (a_14 & ~w12695) | (a_14 & w34721) | (~w12695 & w34721);
assign w29831 = a_14 & ~w26298;
assign w29832 = a_14 & ~w29830;
assign w29833 = w26298 & a_14;
assign w29834 = w980 & b_47;
assign w29835 = w1289 & b_44;
assign w29836 = w3189 & b_32;
assign w29837 = (a_32 & ~w12728) | (a_32 & w34722) | (~w12728 & w34722);
assign w29838 = a_32 & ~w25941;
assign w29839 = a_32 & ~w29837;
assign w29840 = w25941 & a_32;
assign w29841 = w5956 & b_20;
assign w29842 = w12738 & w34723;
assign w29843 = w7607 & b_14;
assign w29844 = w12748 & w34724;
assign w29845 = w9528 & b_8;
assign w29846 = w12758 & w34725;
assign w29847 = a_63 & b_0;
assign w29848 = w10556 & b_5;
assign w29849 = w12791 & w34726;
assign w29850 = w8520 & b_11;
assign w29851 = w12815 & w34727;
assign w29852 = w6755 & b_17;
assign w29853 = w12840 & w34728;
assign w29854 = w5190 & b_23;
assign w29855 = w12865 & w34729;
assign w29856 = w4493 & b_26;
assign w29857 = (a_38 & ~w12883) | (a_38 & w34730) | (~w12883 & w34730);
assign w29858 = a_38 & ~w26303;
assign w29859 = a_38 & ~w29857;
assign w29860 = w26303 & a_38;
assign w29861 = w3797 & b_29;
assign w29862 = a_35 & ~w26304;
assign w29863 = w25942 & a_35;
assign w29864 = w2633 & b_35;
assign w29865 = a_29 & ~w25943;
assign w29866 = w25648 & a_29;
assign w29867 = w2152 & b_38;
assign w29868 = w1688 & b_41;
assign w29869 = (a_23 & ~w12961) | (a_23 & w34731) | (~w12961 & w34731);
assign w29870 = a_23 & ~w26306;
assign w29871 = a_23 & ~w29869;
assign w29872 = w26306 & a_23;
assign w29873 = w233 & b_56;
assign w29874 = w13003 & w34732;
assign w29875 = w93 & b_59;
assign w29876 = (a_5 & ~w13015) | (a_5 & w34733) | (~w13015 & w34733);
assign w29877 = a_5 & ~w27556;
assign w29878 = a_5 & ~w29876;
assign w29879 = w27556 & a_5;
assign w29880 = w651 & b_51;
assign w29881 = w13040 & w34734;
assign w29882 = w1289 & b_45;
assign w29883 = ~w12824 & ~w12823;
assign w29884 = w8520 & b_12;
assign w29885 = w13068 & w34735;
assign w29886 = a_63 & b_1;
assign w29887 = w11614 & b_3;
assign w29888 = (a_62 & ~w13083) | (a_62 & w34736) | (~w13083 & w34736);
assign w29889 = ~w13093 & w34737;
assign w29890 = (w12780 & w13093) | (w12780 & w34738) | (w13093 & w34738);
assign w29891 = w10556 & b_6;
assign w29892 = ~w307 & w10565;
assign w29893 = (a_59 & ~w13101) | (a_59 & w34739) | (~w13101 & w34739);
assign w29894 = ~w29893 & a_59;
assign w29895 = w9528 & b_9;
assign w29896 = w13119 & w34740;
assign w29897 = w7607 & b_15;
assign w29898 = w13142 & w34741;
assign w29899 = w6755 & b_18;
assign w29900 = w13158 & w34742;
assign w29901 = w5956 & b_21;
assign w29902 = w13175 & w34743;
assign w29903 = w5190 & b_24;
assign w29904 = w13191 & w34744;
assign w29905 = w4493 & b_27;
assign w29906 = w13209 & w34745;
assign w29907 = w3797 & b_30;
assign w29908 = (a_35 & ~w13227) | (a_35 & w34746) | (~w13227 & w34746);
assign w29909 = a_35 & ~w26310;
assign w29910 = a_35 & ~w29908;
assign w29911 = w26310 & a_35;
assign w29912 = w3189 & b_33;
assign w29913 = w13244 & w34747;
assign w29914 = ~w12915 & w12919;
assign w29915 = w2633 & b_36;
assign w29916 = (a_29 & ~w13262) | (a_29 & w34748) | (~w13262 & w34748);
assign w29917 = a_29 & ~w26311;
assign w29918 = a_29 & ~w29916;
assign w29919 = w26311 & a_29;
assign w29920 = w2152 & b_39;
assign w29921 = a_26 & ~w26312;
assign w29922 = w25950 & a_26;
assign w29923 = w13059 & ~w13286;
assign w29924 = w1688 & b_42;
assign w29925 = a_23 & ~w26315;
assign w29926 = w25951 & a_23;
assign w29927 = w12954 & w34749;
assign w29928 = w980 & b_48;
assign w29929 = (a_17 & ~w13321) | (a_17 & w34750) | (~w13321 & w34750);
assign w29930 = a_17 & ~w27557;
assign w29931 = a_17 & ~w29929;
assign w29932 = w27557 & a_17;
assign w29933 = w412 & b_54;
assign w29934 = w13345 & w34751;
assign w29935 = w233 & b_57;
assign w29936 = w13358 & w34752;
assign w29937 = ~w12996 & ~w12994;
assign w29938 = w93 & b_60;
assign w29939 = w13374 & w34753;
assign w29940 = ~w29820 & w34754;
assign w29941 = (~w29747 & w34755) | (~w29747 & w34756) | (w34755 & w34756);
assign w29942 = w27010 & b_63;
assign w29943 = w13387 & a_2;
assign w29944 = w93 & b_61;
assign w29945 = w13408 & w34757;
assign w29946 = w412 & b_55;
assign w29947 = w13422 & w34758;
assign w29948 = w980 & b_49;
assign w29949 = a_17 & ~w27558;
assign w29950 = w26320 & a_17;
assign w29951 = w1289 & b_46;
assign w29952 = (a_20 & ~w13449) | (a_20 & w34759) | (~w13449 & w34759);
assign w29953 = a_20 & ~w27561;
assign w29954 = a_20 & ~w29952;
assign w29955 = w27561 & a_20;
assign w29956 = w13308 & ~w13303;
assign w29957 = w1688 & b_43;
assign w29958 = a_23 & ~w27480;
assign w29959 = w26666 & a_23;
assign w29960 = w2152 & b_40;
assign w29961 = w13476 & w34760;
assign w29962 = ~w13269 & w13272;
assign w29963 = ~w13269 & ~w13270;
assign w29964 = w13255 & ~w13251;
assign w29965 = w2633 & b_37;
assign w29966 = ~w13488 & ~w2642;
assign w29967 = ~w13492 & ~w13493;
assign w29968 = ~a_29 & ~w13493;
assign w29969 = ~a_29 & w29967;
assign w29970 = w3797 & b_31;
assign w29971 = w13503 & w34761;
assign w29972 = w5956 & b_22;
assign w29973 = w13513 & w34762;
assign w29974 = w8520 & b_13;
assign w29975 = w13523 & w34763;
assign w29976 = a_63 & b_2;
assign w29977 = w11614 & b_4;
assign w29978 = ~w13536 & ~w11623;
assign w29979 = ~w13540 & ~w13541;
assign w29980 = w13091 & w13548;
assign w29981 = ~w13091 & ~w13548;
assign w29982 = w10556 & b_7;
assign w29983 = w13555 & w34764;
assign w29984 = w9528 & b_10;
assign w29985 = w13572 & w34765;
assign w29986 = w13127 & w13581;
assign w29987 = ~w13127 & ~w13581;
assign w29988 = w13064 & ~w13132;
assign w29989 = w7607 & b_16;
assign w29990 = w13596 & w34766;
assign w29991 = ~w13151 & ~w13149;
assign w29992 = w6755 & b_19;
assign w29993 = w13614 & w34767;
assign w29994 = ~w12851 & w34768;
assign w29995 = w5190 & b_25;
assign w29996 = w13639 & w34769;
assign w29997 = w4493 & b_28;
assign w29998 = w13657 & w34770;
assign w29999 = w13220 & ~w13216;
assign w30000 = w3189 & b_34;
assign w30001 = ~w13675 & ~w3198;
assign w30002 = ~w13679 & ~w13680;
assign w30003 = ~a_32 & ~w13680;
assign w30004 = ~a_32 & w30002;
assign w30005 = w13223 & w34771;
assign w30006 = ~w13683 & ~w13060;
assign w30007 = ~w13697 & ~w13696;
assign w30008 = w651 & b_52;
assign w30009 = ~w13710 & ~w660;
assign w30010 = a_14 & w13715;
assign w30011 = a_14 & ~w27562;
assign w30012 = ~a_14 & ~w13715;
assign w30013 = ~a_14 & w27562;
assign w30014 = w13721 & ~w13708;
assign w30015 = w233 & b_58;
assign w30016 = w13734 & w34772;
assign w30017 = w13756 & ~w12665;
assign w30018 = w13756 & ~w27785;
assign w30019 = ~w13756 & w12665;
assign w30020 = ~w13756 & w27785;
assign w30021 = w651 & b_53;
assign w30022 = (a_14 & ~w13766) | (a_14 & w34773) | (~w13766 & w34773);
assign w30023 = a_14 & ~w26325;
assign w30024 = a_14 & ~w30022;
assign w30025 = w26325 & a_14;
assign w30026 = w1289 & b_47;
assign w30027 = (w13786 & w13290) | (w13786 & w34774) | (w13290 & w34774);
assign w30028 = w13786 & w27790;
assign w30029 = ~w13290 & w34775;
assign w30030 = ~w13786 & ~w27790;
assign w30031 = w2152 & b_41;
assign w30032 = (a_26 & ~w13793) | (a_26 & w34776) | (~w13793 & w34776);
assign w30033 = a_26 & ~w27565;
assign w30034 = a_26 & ~w30032;
assign w30035 = w27565 & a_26;
assign w30036 = w13691 & ~w13497;
assign w30037 = w13509 & ~w13668;
assign w30038 = w3189 & b_35;
assign w30039 = ~w13805 & ~w3198;
assign w30040 = ~w13809 & ~w13810;
assign w30041 = ~a_32 & ~w13810;
assign w30042 = ~a_32 & w30040;
assign w30043 = w3797 & b_32;
assign w30044 = w13820 & w34777;
assign w30045 = w13663 & ~w13652;
assign w30046 = w8520 & b_14;
assign w30047 = w13831 & w34778;
assign w30048 = w11614 & b_5;
assign w30049 = w13841 & w34779;
assign w30050 = a_63 & b_3;
assign w30051 = w34780 & w13843;
assign w30052 = ~w13535 & ~w13533;
assign w30053 = w10556 & b_8;
assign w30054 = w13866 & w34781;
assign w30055 = (~w13096 & w34782) | (~w13096 & w34783) | (w34782 & w34783);
assign w30056 = w9528 & b_11;
assign w30057 = w13884 & w34784;
assign w30058 = w13578 & ~w13894;
assign w30059 = w13529 & ~w13582;
assign w30060 = w7607 & b_17;
assign w30061 = w13910 & w34785;
assign w30062 = w13602 & ~w13591;
assign w30063 = w6755 & b_20;
assign w30064 = w13928 & w34786;
assign w30065 = w13620 & ~w13609;
assign w30066 = w5956 & b_23;
assign w30067 = w13947 & w34787;
assign w30068 = w13519 & ~w13625;
assign w30069 = w5190 & b_26;
assign w30070 = w13965 & w34788;
assign w30071 = (w13645 & w13632) | (w13645 & w34789) | (w13632 & w34789);
assign w30072 = w4493 & b_29;
assign w30073 = w13983 & w34790;
assign w30074 = w13674 & ~w13684;
assign w30075 = w2633 & b_38;
assign w30076 = ~w14005 & ~w2642;
assign w30077 = ~w14009 & ~w14010;
assign w30078 = ~a_29 & ~w14010;
assign w30079 = ~a_29 & w30077;
assign w30080 = ~w14013 & w13684;
assign w30081 = ~w14013 & ~w30074;
assign w30082 = w1688 & b_44;
assign w30083 = ~w14035 & ~w14034;
assign w30084 = ~w14035 & w14036;
assign w30085 = ~w14034 & ~w14036;
assign w30086 = w980 & b_50;
assign w30087 = w13702 & ~w13458;
assign w30088 = (~w14057 & w13456) | (~w14057 & w34791) | (w13456 & w34791);
assign w30089 = ~w14060 & ~w14047;
assign w30090 = w14060 & w14047;
assign w30091 = w412 & b_56;
assign w30092 = ~w14071 & ~w421;
assign w30093 = a_11 & w14076;
assign w30094 = a_11 & ~w26331;
assign w30095 = ~a_11 & ~w14076;
assign w30096 = ~a_11 & w26331;
assign w30097 = w233 & b_59;
assign w30098 = ~w14089 & ~w242;
assign w30099 = a_8 & w14094;
assign w30100 = a_8 & ~w26333;
assign w30101 = ~a_8 & ~w14094;
assign w30102 = ~a_8 & w26333;
assign w30103 = w93 & b_62;
assign w30104 = (w9770 & w34792) | (w9770 & w34793) | (w34792 & w34793);
assign w30105 = w14109 & w34794;
assign w30106 = (~a_5 & ~w14109) | (~a_5 & w34795) | (~w14109 & w34795);
assign w30107 = ~w14113 & w26322;
assign w30108 = ~w14113 & ~w27794;
assign w30109 = ~w14113 & ~w26322;
assign w30110 = ~w14113 & w27794;
assign w30111 = (w13755 & w14122) | (w13755 & w34796) | (w14122 & w34796);
assign w30112 = ~w14124 & ~w25141;
assign w30113 = ~w14123 & ~w13755;
assign w30114 = ~w13756 & w30113;
assign w30115 = w93 & b_63;
assign w30116 = ~w102 & ~w14131;
assign w30117 = w412 & b_57;
assign w30118 = (w9770 & w34797) | (w9770 & w34798) | (w34797 & w34798);
assign w30119 = w14065 & ~w13775;
assign w30120 = w651 & b_54;
assign w30121 = (w13703 & w34799) | (w13703 & w34800) | (w34799 & w34800);
assign w30122 = (~w14164 & w14059) | (~w14164 & w34801) | (w14059 & w34801);
assign w30123 = (w13703 & w34802) | (w13703 & w34803) | (w34802 & w34803);
assign w30124 = (w14164 & w14059) | (w14164 & w34804) | (w14059 & w34804);
assign w30125 = w980 & b_51;
assign w30126 = ~w14169 & ~w989;
assign w30127 = w1289 & b_48;
assign w30128 = w1688 & b_45;
assign w30129 = w14021 & ~w13802;
assign w30130 = ~w14203 & ~w14204;
assign w30131 = w2633 & b_39;
assign w30132 = (a_29 & ~w14212) | (a_29 & w34805) | (~w14212 & w34805);
assign w30133 = a_29 & ~w27567;
assign w30134 = a_29 & ~w30132;
assign w30135 = w27567 & a_29;
assign w30136 = (w14218 & w13804) | (w14218 & w34806) | (w13804 & w34806);
assign w30137 = ~w13804 & w34807;
assign w30138 = w3797 & b_33;
assign w30139 = w14225 & w34808;
assign w30140 = w6755 & b_21;
assign w30141 = w14235 & w34809;
assign w30142 = w9528 & b_12;
assign w30143 = w14245 & w34810;
assign w30144 = w11614 & b_6;
assign w30145 = (a_62 & ~w14255) | (a_62 & w34811) | (~w14255 & w34811);
assign w30146 = ~w30145 & a_62;
assign w30147 = a_63 & b_4;
assign w30148 = ~w14257 & w34812;
assign w30149 = w10556 & b_9;
assign w30150 = w14281 & w34813;
assign w30151 = (w13872 & w13858) | (w13872 & w34814) | (w13858 & w34814);
assign w30152 = w13890 & ~w13879;
assign w30153 = w8520 & b_15;
assign w30154 = w14307 & w34815;
assign w30155 = w14302 & ~w14313;
assign w30156 = (w13837 & w13895) | (w13837 & w34816) | (w13895 & w34816);
assign w30157 = w7607 & b_18;
assign w30158 = w14325 & w34817;
assign w30159 = w13916 & ~w13905;
assign w30160 = w13934 & ~w13923;
assign w30161 = w5956 & b_24;
assign w30162 = w14350 & w34818;
assign w30163 = w13953 & ~w13940;
assign w30164 = w5190 & b_27;
assign w30165 = w14368 & w34819;
assign w30166 = (w13971 & w13957) | (w13971 & w34820) | (w13957 & w34820);
assign w30167 = w4493 & b_30;
assign w30168 = w14386 & w34821;
assign w30169 = (w13989 & w13975) | (w13989 & w34822) | (w13975 & w34822);
assign w30170 = w3189 & b_36;
assign w30171 = ~w14404 & ~w3198;
assign w30172 = ~w14408 & ~w14409;
assign w30173 = ~a_32 & ~w14409;
assign w30174 = ~a_32 & w30172;
assign w30175 = ~w14412 & w13993;
assign w30176 = (~w14412 & w13993) | (~w14412 & w34823) | (w13993 & w34823);
assign w30177 = w14412 & ~w13993;
assign w30178 = ~w13993 & w34824;
assign w30179 = w2152 & b_42;
assign w30180 = ~w14424 & ~w2161;
assign w30181 = ~w14432 & w14014;
assign w30182 = (~w14432 & w14014) | (~w14432 & w34825) | (w14014 & w34825);
assign w30183 = w14432 & w14014;
assign w30184 = (w14432 & w14014) | (w14432 & w34826) | (w14014 & w34826);
assign w30185 = w14434 & ~w14423;
assign w30186 = (~w14440 & ~w14205) | (~w14440 & w34827) | (~w14205 & w34827);
assign w30187 = w14205 & w34828;
assign w30188 = w233 & b_60;
assign w30189 = ~w14460 & ~w242;
assign w30190 = ~w14464 & ~w14465;
assign w30191 = ~a_8 & ~w14465;
assign w30192 = ~a_8 & w30190;
assign w30193 = ~w14456 & w34829;
assign w30194 = ~w14483 & w14121;
assign w30195 = ~w14483 & ~w25142;
assign w30196 = ~w14482 & ~w14121;
assign w30197 = ~w14482 & w25142;
assign w30198 = (~w14480 & w14483) | (~w14480 & w34830) | (w14483 & w34830);
assign w30199 = (~w14480 & w25143) | (~w14480 & w25142) | (w25143 & w25142);
assign w30200 = ~w14476 & ~w14137;
assign w30201 = w14458 & ~w14469;
assign w30202 = w233 & b_61;
assign w30203 = w14493 & w34831;
assign w30204 = (~w14083 & w34832) | (~w14083 & w34833) | (w34832 & w34833);
assign w30205 = (~w14499 & w14469) | (~w14499 & w34834) | (w14469 & w34834);
assign w30206 = w412 & b_58;
assign w30207 = w14507 & w34835;
assign w30208 = w14447 & ~w14178;
assign w30209 = w980 & b_52;
assign w30210 = (a_17 & ~w14522) | (a_17 & w34836) | (~w14522 & w34836);
assign w30211 = a_17 & ~w26345;
assign w30212 = a_17 & ~w30210;
assign w30213 = w26345 & a_17;
assign w30214 = w1688 & b_46;
assign w30215 = a_23 & ~w27801;
assign w30216 = w27568 & a_23;
assign w30217 = w2152 & b_43;
assign w30218 = a_26 & ~w27570;
assign w30219 = w26347 & a_26;
assign w30220 = (~w14017 & w34837) | (~w14017 & w34838) | (w34837 & w34838);
assign w30221 = ~w14557 & ~w26346;
assign w30222 = (w14017 & w34839) | (w14017 & w34840) | (w34839 & w34840);
assign w30223 = ~w14557 & w26346;
assign w30224 = w2633 & b_40;
assign w30225 = w14564 & w34841;
assign w30226 = w14419 & ~w14220;
assign w30227 = (w14231 & w14396) | (w14231 & w34842) | (w14396 & w34842);
assign w30228 = w14392 & ~w14381;
assign w30229 = (w14374 & w14361) | (w14374 & w34843) | (w14361 & w34843);
assign w30230 = w14241 & ~w14336;
assign w30231 = (w14331 & w14317) | (w14331 & w34844) | (w14317 & w34844);
assign w30232 = (w14287 & w14273) | (w14287 & w34845) | (w14273 & w34845);
assign w30233 = w10556 & b_10;
assign w30234 = w14583 & w34846;
assign w30235 = a_63 & b_5;
assign w30236 = ~w14266 & ~w14598;
assign w30237 = w14266 & w14598;
assign w30238 = w11614 & b_7;
assign w30239 = w14605 & w34847;
assign w30240 = w14616 & ~w14579;
assign w30241 = w9528 & b_13;
assign w30242 = w14626 & w34848;
assign w30243 = (w14251 & ~w14290) | (w14251 & w34849) | (~w14290 & w34849);
assign w30244 = ~w14635 & w14636;
assign w30245 = w14635 & ~w14636;
assign w30246 = w8520 & b_16;
assign w30247 = w14643 & w34850;
assign w30248 = w7607 & b_19;
assign w30249 = w14661 & w34851;
assign w30250 = ~w14670 & ~w14578;
assign w30251 = w14670 & w14578;
assign w30252 = w6755 & b_22;
assign w30253 = w14677 & w34852;
assign w30254 = w5956 & b_25;
assign w30255 = w14693 & w34853;
assign w30256 = w14356 & ~w14345;
assign w30257 = w5190 & b_28;
assign w30258 = w14711 & w34854;
assign w30259 = ~w14719 & ~w14718;
assign w30260 = ~w30259 & ~w14718;
assign w30261 = w4493 & b_31;
assign w30262 = w14728 & w34855;
assign w30263 = w3797 & b_34;
assign w30264 = w14745 & w34856;
assign w30265 = w3189 & b_37;
assign w30266 = w14761 & w34857;
assign w30267 = w14403 & ~w14413;
assign w30268 = w14560 & ~w14777;
assign w30269 = ~w14560 & w14777;
assign w30270 = w1289 & b_49;
assign w30271 = (a_20 & ~w14788) | (a_20 & w34858) | (~w14788 & w34858);
assign w30272 = a_20 & ~w27572;
assign w30273 = a_20 & ~w30271;
assign w30274 = w27572 & a_20;
assign w30275 = w651 & b_55;
assign w30276 = w14810 & w34859;
assign w30277 = (w25144 & ~w14483) | (w25144 & w34860) | (~w14483 & w34860);
assign w30278 = (w25144 & w25145) | (w25144 & ~w25142) | (w25145 & ~w25142);
assign w30279 = w14824 & ~w14516;
assign w30280 = w233 & b_62;
assign w30281 = (w9770 & w34861) | (w9770 & w34862) | (w34861 & w34862);
assign w30282 = w14841 & w34863;
assign w30283 = (~a_8 & ~w14841) | (~a_8 & w34864) | (~w14841 & w34864);
assign w30284 = w412 & b_59;
assign w30285 = w14852 & w34865;
assign w30286 = w14806 & ~w14818;
assign w30287 = w651 & b_56;
assign w30288 = ~w14863 & ~w660;
assign w30289 = a_14 & w14868;
assign w30290 = a_14 & ~w27573;
assign w30291 = ~a_14 & ~w14868;
assign w30292 = ~a_14 & w27573;
assign w30293 = w980 & b_53;
assign w30294 = (a_17 & ~w14878) | (a_17 & w34866) | (~w14878 & w34866);
assign w30295 = a_17 & ~w27574;
assign w30296 = a_17 & ~w30294;
assign w30297 = w27574 & a_17;
assign w30298 = w1289 & b_50;
assign w30299 = a_20 & ~w27803;
assign w30300 = w26350 & a_20;
assign w30301 = w1688 & b_47;
assign w30302 = w14558 & ~w14912;
assign w30303 = ~w14558 & ~w14912;
assign w30304 = w14558 & w14912;
assign w30305 = ~w14774 & ~w14572;
assign w30306 = w2152 & b_44;
assign w30307 = ~w14919 & ~w2161;
assign w30308 = w2633 & b_41;
assign w30309 = w14934 & w34867;
assign w30310 = (~w14757 & w14768) | (~w14757 & w34868) | (w14768 & w34868);
assign w30311 = w3189 & b_38;
assign w30312 = w14947 & w34869;
assign w30313 = (w14953 & w14741) | (w14953 & w34870) | (w14741 & w34870);
assign w30314 = ~w14741 & w34871;
assign w30315 = w3797 & b_35;
assign w30316 = w14960 & w34872;
assign w30317 = w14575 & ~w14735;
assign w30318 = w4493 & b_32;
assign w30319 = w14971 & w34873;
assign w30320 = w14611 & ~w14600;
assign w30321 = w14595 & ~w14979;
assign w30322 = a_63 & b_6;
assign w30323 = w11614 & b_8;
assign w30324 = ~w14987 & ~w11623;
assign w30325 = ~w14991 & ~w14992;
assign w30326 = ~a_62 & ~w14992;
assign w30327 = ~a_62 & w30325;
assign w30328 = w14994 & w14986;
assign w30329 = ~w14994 & ~w14986;
assign w30330 = w10556 & b_11;
assign w30331 = w15004 & w34874;
assign w30332 = w9528 & b_14;
assign w30333 = w15022 & w34875;
assign w30334 = w8520 & b_17;
assign w30335 = w15040 & w34876;
assign w30336 = w14654 & ~w14650;
assign w30337 = w7607 & b_20;
assign w30338 = w15058 & w34877;
assign w30339 = w14670 & ~w14578;
assign w30340 = w6755 & b_23;
assign w30341 = w15077 & w34878;
assign w30342 = w14577 & ~w14684;
assign w30343 = ~w15086 & w15087;
assign w30344 = w15086 & ~w15087;
assign w30345 = w5956 & b_26;
assign w30346 = w15094 & w34879;
assign w30347 = w14704 & ~w14700;
assign w30348 = ~w15103 & w15104;
assign w30349 = w15103 & ~w15104;
assign w30350 = w5190 & b_29;
assign w30351 = w15111 & w34880;
assign w30352 = w34881 & w14941;
assign w30353 = (~w14941 & w34882) | (~w14941 & w34883) | (w34882 & w34883);
assign w30354 = ~w15159 & ~w15158;
assign w30355 = w14828 & ~w14500;
assign w30356 = ~w14832 & w15168;
assign w30357 = ~w15167 & w34884;
assign w30358 = ~w30354 & ~w14846;
assign w30359 = w15157 & ~w14861;
assign w30360 = w233 & b_63;
assign w30361 = ~w242 & ~w15174;
assign w30362 = w980 & b_54;
assign w30363 = (w15147 & w14899) | (w15147 & w34885) | (w14899 & w34885);
assign w30364 = w1688 & b_48;
assign w30365 = w15140 & ~w14928;
assign w30366 = w2152 & b_45;
assign w30367 = w34886 & w14941;
assign w30368 = w14942 & ~w15220;
assign w30369 = ~w14942 & ~w15220;
assign w30370 = ~w14941 & w34887;
assign w30371 = w3189 & b_39;
assign w30372 = (w14966 & w14967) | (w14966 & w34888) | (w14967 & w34888);
assign w30373 = ~w15234 & ~w15235;
assign w30374 = w4493 & b_33;
assign w30375 = w15243 & w34889;
assign w30376 = w6755 & b_24;
assign w30377 = w15253 & w34890;
assign w30378 = (w15064 & w15050) | (w15064 & w34891) | (w15050 & w34891);
assign w30379 = w7607 & b_21;
assign w30380 = w15264 & w34892;
assign w30381 = w15046 & ~w15035;
assign w30382 = (w15010 & w14978) | (w15010 & w34893) | (w14978 & w34893);
assign w30383 = a_63 & b_7;
assign w30384 = ~w15277 & ~w15278;
assign w30385 = w14984 & w30384;
assign w30386 = ~w15278 & ~w30384;
assign w30387 = ~w15278 & ~w30385;
assign w30388 = ~w30385 & w30384;
assign w30389 = w11614 & b_9;
assign w30390 = w15285 & w34894;
assign w30391 = w15281 & w15291;
assign w30392 = ~w15281 & ~w15291;
assign w30393 = w10556 & b_12;
assign w30394 = w15298 & w34895;
assign w30395 = w9528 & b_15;
assign w30396 = w15314 & w34896;
assign w30397 = w15028 & ~w15017;
assign w30398 = w8520 & b_18;
assign w30399 = w15332 & w34897;
assign w30400 = w15344 & ~w15270;
assign w30401 = (w15083 & w15068) | (w15083 & w34898) | (w15068 & w34898);
assign w30402 = w5956 & b_27;
assign w30403 = w15363 & w34899;
assign w30404 = w15100 & ~w15089;
assign w30405 = w5190 & b_30;
assign w30406 = w15381 & w34900;
assign w30407 = w15117 & ~w15106;
assign w30408 = w14977 & ~w15121;
assign w30409 = ~w15397 & w15398;
assign w30410 = w15397 & ~w15398;
assign w30411 = w3797 & b_36;
assign w30412 = w15405 & w34901;
assign w30413 = (~w15413 & ~w15236) | (~w15413 & w34902) | (~w15236 & w34902);
assign w30414 = w15412 & ~w15413;
assign w30415 = ~w15412 & ~w15413;
assign w30416 = ~w15412 & w30414;
assign w30417 = w15133 & ~w14955;
assign w30418 = w2633 & b_42;
assign w30419 = ~w15420 & ~w2642;
assign w30420 = ~w15221 & w34903;
assign w30421 = (~w15221 & w33590) | (~w15221 & w34904) | (w33590 & w34904);
assign w30422 = (~w15436 & w15221) | (~w15436 & w34905) | (w15221 & w34905);
assign w30423 = ~w14914 & w15144;
assign w30424 = ~w14914 & ~w14915;
assign w30425 = w1289 & b_51;
assign w30426 = ~w15445 & ~w1298;
assign w30427 = a_20 & w15450;
assign w30428 = a_20 & ~w26362;
assign w30429 = ~a_20 & ~w15450;
assign w30430 = ~a_20 & w26362;
assign w30431 = w651 & b_57;
assign w30432 = (w9770 & w34906) | (w9770 & w34907) | (w34906 & w34907);
assign w30433 = w15151 & ~w14887;
assign w30434 = ~w15478 & ~w15465;
assign w30435 = w15478 & w15465;
assign w30436 = ~w27581 & ~w14872;
assign w30437 = w412 & b_60;
assign w30438 = ~w15484 & ~w421;
assign w30439 = ~w15488 & ~w15489;
assign w30440 = ~a_11 & ~w15489;
assign w30441 = ~a_11 & w30439;
assign w30442 = w15495 & ~w15482;
assign w30443 = w15182 & w15499;
assign w30444 = ~w15182 & ~w15499;
assign w30445 = (~w15506 & w25147) | (~w15506 & ~w15168) | (w25147 & ~w15168);
assign w30446 = (~w15506 & w25147) | (~w15506 & w25146) | (w25147 & w25146);
assign w30447 = ~w15505 & w30357;
assign w30448 = ~w25146 & w34908;
assign w30449 = (w25148 & w25149) | (w25148 & ~w25146) | (w25149 & ~w25146);
assign w30450 = w412 & b_61;
assign w30451 = w15515 & w34909;
assign w30452 = ~w15483 & w34910;
assign w30453 = (~w15521 & w15483) | (~w15521 & w34911) | (w15483 & w34911);
assign w30454 = w15478 & ~w15465;
assign w30455 = w651 & b_58;
assign w30456 = w15529 & w34912;
assign w30457 = ~w15476 & w34913;
assign w30458 = (~w15535 & w15476) | (~w15535 & w34914) | (w15476 & w34914);
assign w30459 = w980 & b_55;
assign w30460 = w15542 & w34915;
assign w30461 = w1289 & b_52;
assign w30462 = w15557 & w34916;
assign w30463 = ~w15444 & w34917;
assign w30464 = (~w15563 & w15444) | (~w15563 & w34918) | (w15444 & w34918);
assign w30465 = w2152 & b_46;
assign w30466 = w15571 & w34919;
assign w30467 = w27811 & ~w15224;
assign w30468 = (~w15224 & w27811) | (~w15224 & ~w15223) | (w27811 & ~w15223);
assign w30469 = w2633 & b_43;
assign w30470 = a_29 & ~w26363;
assign w30471 = w25978 & a_29;
assign w30472 = ~w15419 & w34920;
assign w30473 = ~w15592 & ~w15432;
assign w30474 = (~w15592 & w15419) | (~w15592 & w34921) | (w15419 & w34921);
assign w30475 = ~w15592 & w15432;
assign w30476 = (~w26360 & w34922) | (~w26360 & w34923) | (w34922 & w34923);
assign w30477 = w3189 & b_40;
assign w30478 = w15601 & w34924;
assign w30479 = (w15249 & ~w15390) | (w15249 & w34925) | (~w15390 & w34925);
assign w30480 = (w15387 & w15373) | (w15387 & w34926) | (w15373 & w34926);
assign w30481 = w15369 & ~w15358;
assign w30482 = w7607 & b_22;
assign w30483 = w15619 & w34927;
assign w30484 = w9528 & b_16;
assign w30485 = w15629 & w34928;
assign w30486 = w15281 & ~w15291;
assign w30487 = w11614 & b_10;
assign w30488 = w15641 & w34929;
assign w30489 = a_63 & b_8;
assign w30490 = w15656 & ~w30386;
assign w30491 = w15656 & ~w30387;
assign w30492 = ~w15656 & w30386;
assign w30493 = ~w15656 & w30387;
assign w30494 = w10556 & b_13;
assign w30495 = w15666 & w34930;
assign w30496 = w15320 & ~w15309;
assign w30497 = ~w15681 & w15682;
assign w30498 = w15681 & ~w15682;
assign w30499 = w8520 & b_19;
assign w30500 = w15689 & w34931;
assign w30501 = w15338 & ~w15327;
assign w30502 = w6755 & b_25;
assign w30503 = w15715 & w34932;
assign w30504 = (w15259 & w15260) | (w15259 & w34933) | (w15260 & w34933);
assign w30505 = ~w15724 & w15725;
assign w30506 = w15724 & ~w15725;
assign w30507 = w5956 & b_28;
assign w30508 = w15732 & w34934;
assign w30509 = ~w15740 & ~w15739;
assign w30510 = w5190 & b_31;
assign w30511 = w15749 & w34935;
assign w30512 = w4493 & b_34;
assign w30513 = w15766 & w34936;
assign w30514 = w3797 & b_37;
assign w30515 = w15782 & w34937;
assign w30516 = w15411 & ~w15400;
assign w30517 = w15791 & ~w15793;
assign w30518 = w34938 & w15597;
assign w30519 = w1688 & b_49;
assign w30520 = (a_23 & ~w15812) | (a_23 & w34939) | (~w15812 & w34939);
assign w30521 = a_23 & ~w27812;
assign w30522 = a_23 & ~w30520;
assign w30523 = w27812 & a_23;
assign w30524 = ~w15209 & w15440;
assign w30525 = ~w15832 & ~w15831;
assign w30526 = w15524 & w15837;
assign w30527 = ~w15524 & ~w15837;
assign w30528 = (w15168 & w34940) | (w15168 & w34941) | (w34940 & w34941);
assign w30529 = ~w15843 & w30449;
assign w30530 = (~w25146 & w34942) | (~w25146 & w34943) | (w34942 & w34943);
assign w30531 = w15524 & ~w15837;
assign w30532 = w651 & b_59;
assign w30533 = w15853 & w34944;
assign w30534 = (w15830 & w15549) | (w15830 & w34945) | (w15549 & w34945);
assign w30535 = w1289 & b_53;
assign w30536 = (a_20 & ~w15868) | (a_20 & w34946) | (~w15868 & w34946);
assign w30537 = a_20 & ~w27814;
assign w30538 = a_20 & ~w30536;
assign w30539 = w27814 & a_20;
assign w30540 = (w15874 & w15819) | (w15874 & w34947) | (w15819 & w34947);
assign w30541 = ~w15806 & w34948;
assign w30542 = ~w15819 & w34949;
assign w30543 = (~w15874 & w15806) | (~w15874 & w34950) | (w15806 & w34950);
assign w30544 = w1688 & b_50;
assign w30545 = w15881 & w34951;
assign w30546 = w2152 & b_47;
assign w30547 = ~w15901 & ~w15900;
assign w30548 = ~w15901 & w15902;
assign w30549 = w3189 & b_41;
assign w30550 = (a_32 & ~w15910) | (a_32 & w34952) | (~w15910 & w34952);
assign w30551 = a_32 & ~w26682;
assign w30552 = a_32 & ~w30550;
assign w30553 = w26682 & a_32;
assign w30554 = (w15916 & ~w15778) | (w15916 & w34953) | (~w15778 & w34953);
assign w30555 = w15778 & w34954;
assign w30556 = w3797 & b_38;
assign w30557 = w15923 & w34955;
assign w30558 = w15612 & ~w15773;
assign w30559 = w4493 & b_35;
assign w30560 = w15934 & w34956;
assign w30561 = w15613 & ~w15756;
assign w30562 = w5190 & b_32;
assign w30563 = w15945 & w34957;
assign w30564 = w11614 & b_11;
assign w30565 = w15955 & w34958;
assign w30566 = a_63 & b_9;
assign w30567 = w15650 & ~w15965;
assign w30568 = w15959 & ~w15970;
assign w30569 = w15647 & ~w15657;
assign w30570 = w10556 & b_14;
assign w30571 = w15983 & w34959;
assign w30572 = w15978 & ~w15989;
assign w30573 = w9528 & b_17;
assign w30574 = w16001 & w34960;
assign w30575 = ~w16010 & w16011;
assign w30576 = w16010 & ~w16011;
assign w30577 = w8520 & b_20;
assign w30578 = w16018 & w34961;
assign w30579 = w15700 & ~w15696;
assign w30580 = ~w16027 & w16028;
assign w30581 = w16027 & ~w16028;
assign w30582 = w7607 & b_23;
assign w30583 = w16035 & w34962;
assign w30584 = w6755 & b_26;
assign w30585 = w16053 & w34963;
assign w30586 = w5956 & b_29;
assign w30587 = w16071 & w34964;
assign w30588 = w16089 & ~w15940;
assign w30589 = w2633 & b_44;
assign w30590 = ~w16106 & ~w2642;
assign w30591 = ~w15597 & w34965;
assign w30592 = (~w15597 & w34966) | (~w15597 & w34967) | (w34966 & w34967);
assign w30593 = ~w15597 & w34968;
assign w30594 = (~w15597 & w34969) | (~w15597 & w34970) | (w34969 & w34970);
assign w30595 = w16115 & ~w16105;
assign w30596 = ~w27815 & ~w16127;
assign w30597 = w980 & b_56;
assign w30598 = ~w16133 & ~w989;
assign w30599 = ~w16137 & ~w16138;
assign w30600 = ~a_17 & ~w16138;
assign w30601 = ~a_17 & w30599;
assign w30602 = (w15458 & w34971) | (w15458 & w34972) | (w34971 & w34972);
assign w30603 = ~w16141 & ~w25665;
assign w30604 = (~w15458 & w34973) | (~w15458 & w34974) | (w34973 & w34974);
assign w30605 = ~w16141 & w25665;
assign w30606 = w16144 & ~w16131;
assign w30607 = w34975 & w15860;
assign w30608 = ~w15476 & w34976;
assign w30609 = w412 & b_62;
assign w30610 = (w9770 & w34977) | (w9770 & w34978) | (w34977 & w34978);
assign w30611 = w16158 & w34979;
assign w30612 = (~a_11 & ~w16158) | (~a_11 & w34980) | (~w16158 & w34980);
assign w30613 = ~w16162 & w16154;
assign w30614 = (w15525 & w34981) | (w15525 & w34982) | (w34981 & w34982);
assign w30615 = w16162 & w16153;
assign w30616 = (w25146 & w34983) | (w25146 & w34984) | (w34983 & w34984);
assign w30617 = (~w16174 & w25152) | (~w16174 & w27438) | (w25152 & w27438);
assign w30618 = ~w27438 & w34985;
assign w30619 = ~w16173 & w30530;
assign w30620 = (~w25146 & w34986) | (~w25146 & w34987) | (w34986 & w34987);
assign w30621 = w16153 & ~w16163;
assign w30622 = w412 & b_63;
assign w30623 = ~w421 & ~w16180;
assign w30624 = ~w15860 & w34988;
assign w30625 = (~w16185 & w15860) | (~w16185 & w34989) | (w15860 & w34989);
assign w30626 = w651 & b_60;
assign w30627 = ~w16189 & ~w660;
assign w30628 = ~w16193 & ~w16194;
assign w30629 = ~a_14 & ~w16194;
assign w30630 = ~a_14 & w30628;
assign w30631 = ~w16197 & w16142;
assign w30632 = ~w16197 & ~w27816;
assign w30633 = w16197 & ~w16142;
assign w30634 = w16197 & w27816;
assign w30635 = w980 & b_57;
assign w30636 = w16204 & w34990;
assign w30637 = ~w27815 & ~w15876;
assign w30638 = w1289 & b_54;
assign w30639 = a_20 & ~w26365;
assign w30640 = w25984 & a_20;
assign w30641 = w2152 & b_48;
assign w30642 = ~w16230 & ~w2161;
assign w30643 = (~w15611 & w34991) | (~w15611 & w34992) | (w34991 & w34992);
assign w30644 = (~w15611 & w34993) | (~w15611 & w34994) | (w34993 & w34994);
assign w30645 = (w15611 & w34995) | (w15611 & w34996) | (w34995 & w34996);
assign w30646 = (w15611 & w34997) | (w15611 & w34998) | (w34997 & w34998);
assign w30647 = w2633 & b_45;
assign w30648 = ~w16249 & ~w16250;
assign w30649 = w3189 & b_42;
assign w30650 = ~w16255 & ~w3198;
assign w30651 = ~w16263 & w16094;
assign w30652 = (~w16263 & w16094) | (~w16263 & w34999) | (w16094 & w34999);
assign w30653 = w16263 & ~w16094;
assign w30654 = ~w16094 & w35000;
assign w30655 = w3797 & b_39;
assign w30656 = w16270 & w35001;
assign w30657 = w5190 & b_33;
assign w30658 = w16281 & w35002;
assign w30659 = w16041 & ~w16030;
assign w30660 = w7607 & b_24;
assign w30661 = w16292 & w35003;
assign w30662 = w16024 & ~w16013;
assign w30663 = w8520 & b_21;
assign w30664 = w16303 & w35004;
assign w30665 = (w16007 & w15993) | (w16007 & w35005) | (w15993 & w35005);
assign w30666 = a_63 & b_10;
assign w30667 = w15967 & ~w16318;
assign w30668 = ~w15967 & ~w16318;
assign w30669 = w11614 & b_12;
assign w30670 = w16326 & w35006;
assign w30671 = w16321 & ~w16332;
assign w30672 = w10556 & b_15;
assign w30673 = w16340 & w35007;
assign w30674 = ~w16349 & w16350;
assign w30675 = w16349 & ~w16350;
assign w30676 = w9528 & b_18;
assign w30677 = w16357 & w35008;
assign w30678 = w16368 & ~w16309;
assign w30679 = w16309 & ~w16368;
assign w30680 = w6755 & b_27;
assign w30681 = w16385 & w35009;
assign w30682 = w16059 & ~w16048;
assign w30683 = w5956 & b_30;
assign w30684 = w16403 & w35010;
assign w30685 = w16077 & ~w16066;
assign w30686 = w15951 & ~w16081;
assign w30687 = w4493 & b_36;
assign w30688 = w16428 & w35011;
assign w30689 = ~w16252 & ~w16448;
assign w30690 = w16252 & w16448;
assign w30691 = w1688 & b_51;
assign w30692 = ~w16456 & ~w1697;
assign w30693 = w16467 & ~w16454;
assign w30694 = w16227 & ~w16472;
assign w30695 = ~w16478 & ~w16477;
assign w30696 = w16188 & w16482;
assign w30697 = (~w16482 & w16150) | (~w16482 & w35012) | (w16150 & w35012);
assign w30698 = ~w16485 & w16163;
assign w30699 = ~w16485 & ~w30621;
assign w30700 = (~w27438 & w35013) | (~w27438 & w35014) | (w35013 & w35014);
assign w30701 = ~w16488 & w30620;
assign w30702 = (~w27438 & w35015) | (~w27438 & w35016) | (w35015 & w35016);
assign w30703 = ~w16150 & w35017;
assign w30704 = ~w30695 & ~w16198;
assign w30705 = w651 & b_61;
assign w30706 = w16499 & w35018;
assign w30707 = w980 & b_58;
assign w30708 = w16512 & w35019;
assign w30709 = ~w16211 & w35020;
assign w30710 = (~w16518 & w16211) | (~w16518 & w35021) | (w16211 & w35021);
assign w30711 = w1289 & b_55;
assign w30712 = w16525 & w35022;
assign w30713 = (w16531 & w16225) | (w16531 & w35023) | (w16225 & w35023);
assign w30714 = ~w16225 & w35024;
assign w30715 = w1688 & b_52;
assign w30716 = (a_23 & ~w16539) | (a_23 & w35025) | (~w16539 & w35025);
assign w30717 = a_23 & ~w26372;
assign w30718 = a_23 & ~w30716;
assign w30719 = w26372 & a_23;
assign w30720 = ~w16545 & w16465;
assign w30721 = ~w16545 & ~w26371;
assign w30722 = ~w16545 & ~w16465;
assign w30723 = ~w16545 & w26371;
assign w30724 = w2152 & b_49;
assign w30725 = w16553 & w35026;
assign w30726 = (w16117 & w35027) | (w16117 & w35028) | (w35027 & w35028);
assign w30727 = w2633 & b_46;
assign w30728 = a_29 & ~w27593;
assign w30729 = w26685 & a_29;
assign w30730 = (w16276 & w16277) | (w16276 & w35029) | (w16277 & w35029);
assign w30731 = (w16434 & w16420) | (w16434 & w35030) | (w16420 & w35030);
assign w30732 = w16287 & ~w16414;
assign w30733 = (w16409 & w16395) | (w16409 & w35031) | (w16395 & w35031);
assign w30734 = (w16391 & ~w16378) | (w16391 & w35032) | (~w16378 & w35032);
assign w30735 = w8520 & b_22;
assign w30736 = w16587 & w35033;
assign w30737 = ~w16315 & w16318;
assign w30738 = (~w16315 & ~w15967) | (~w16315 & w30737) | (~w15967 & w30737);
assign w30739 = w11614 & b_13;
assign w30740 = w16598 & w35034;
assign w30741 = a_63 & b_11;
assign w30742 = w35035 & w16600;
assign w30743 = w10556 & b_16;
assign w30744 = w16625 & w35036;
assign w30745 = w16619 & ~w16631;
assign w30746 = w16346 & ~w16333;
assign w30747 = w9528 & b_19;
assign w30748 = w16643 & w35037;
assign w30749 = w16363 & ~w16352;
assign w30750 = w16652 & ~w16653;
assign w30751 = ~w16652 & w16653;
assign w30752 = w7607 & b_25;
assign w30753 = w16668 & w35038;
assign w30754 = w16662 & ~w16674;
assign w30755 = (w16298 & ~w16372) | (w16298 & w35039) | (~w16372 & w35039);
assign w30756 = w6755 & b_28;
assign w30757 = w16686 & w35040;
assign w30758 = (w16381 & w35041) | (w16381 & w35042) | (w35041 & w35042);
assign w30759 = ~w16693 & ~w16694;
assign w30760 = w5956 & b_31;
assign w30761 = w16704 & w35043;
assign w30762 = ~w16713 & ~w16581;
assign w30763 = w16713 & w16581;
assign w30764 = w5190 & b_34;
assign w30765 = w16720 & w35044;
assign w30766 = w4493 & b_37;
assign w30767 = w16736 & w35045;
assign w30768 = ~w16745 & ~w16579;
assign w30769 = w16745 & w16579;
assign w30770 = w3797 & b_40;
assign w30771 = w16752 & w35046;
assign w30772 = w3189 & b_43;
assign w30773 = (a_32 & ~w16769) | (a_32 & w35047) | (~w16769 & w35047);
assign w30774 = a_32 & ~w27595;
assign w30775 = a_32 & ~w30773;
assign w30776 = w27595 & a_32;
assign w30777 = (~w16097 & w35048) | (~w16097 & w35049) | (w35048 & w35049);
assign w30778 = ~w30777 & ~w16775;
assign w30779 = ~w16445 & w35050;
assign w30780 = (~w16764 & w16445) | (~w16764 & w35051) | (w16445 & w35051);
assign w30781 = w16784 & ~w16785;
assign w30782 = ~w16784 & ~w16785;
assign w30783 = ~w16784 & w30781;
assign w30784 = ~w16792 & ~w16791;
assign w30785 = ~w30784 & ~w16792;
assign w30786 = w16508 & w16796;
assign w30787 = ~w16508 & ~w16796;
assign w30788 = w16186 & ~w16799;
assign w30789 = ~w16186 & ~w16799;
assign w30790 = (w27438 & w35052) | (w27438 & w35053) | (w35052 & w35053);
assign w30791 = (~w16803 & w25157) | (~w16803 & w27757) | (w25157 & w27757);
assign w30792 = ~w27757 & w35054;
assign w30793 = ~w16802 & w30702;
assign w30794 = (~w27438 & w35055) | (~w27438 & w35056) | (w35055 & w35056);
assign w30795 = w16508 & ~w16796;
assign w30796 = w980 & b_59;
assign w30797 = w16812 & w35057;
assign w30798 = w16790 & ~w16533;
assign w30799 = w1688 & b_53;
assign w30800 = w16827 & w35058;
assign w30801 = (w16783 & w16560) | (w16783 & w35059) | (w16560 & w35059);
assign w30802 = w2633 & b_47;
assign w30803 = a_29 & ~w27597;
assign w30804 = w26373 & a_29;
assign w30805 = (w16445 & w35060) | (w16445 & w35061) | (w35060 & w35061);
assign w30806 = (~w16445 & w35062) | (~w16445 & w35063) | (w35062 & w35063);
assign w30807 = w3797 & b_41;
assign w30808 = w16857 & w35064;
assign w30809 = w16745 & ~w16579;
assign w30810 = w4493 & b_38;
assign w30811 = w16869 & w35065;
assign w30812 = w16580 & ~w16727;
assign w30813 = w5190 & b_35;
assign w30814 = w16880 & w35066;
assign w30815 = w16713 & ~w16581;
assign w30816 = w5956 & b_32;
assign w30817 = w16892 & w35067;
assign w30818 = w6755 & b_29;
assign w30819 = w16902 & w35068;
assign w30820 = w16679 & ~w16675;
assign w30821 = a_63 & b_12;
assign w30822 = w16607 & ~w16913;
assign w30823 = w11614 & b_14;
assign w30824 = w16922 & w35069;
assign w30825 = (~w16924 & w35070) | (~w16924 & w35071) | (w35070 & w35071);
assign w30826 = w35072 & w16924;
assign w30827 = w16594 & ~w16614;
assign w30828 = w10556 & b_17;
assign w30829 = w16937 & w35073;
assign w30830 = w16636 & ~w16632;
assign w30831 = w9528 & b_20;
assign w30832 = w16955 & w35074;
assign w30833 = w8520 & b_23;
assign w30834 = w16973 & w35075;
assign w30835 = w16583 & ~w16657;
assign w30836 = w7607 & b_26;
assign w30837 = w16991 & w35076;
assign w30838 = ~w17000 & w16908;
assign w30839 = ~w17014 & w16886;
assign w30840 = ~w17021 & ~w16876;
assign w30841 = w3189 & b_44;
assign w30842 = ~w17038 & ~w3198;
assign w30843 = ~w16748 & w35077;
assign w30844 = ~w16748 & w35078;
assign w30845 = ~w17049 & ~w17037;
assign w30846 = ~w17050 & ~w17049;
assign w30847 = ~w17050 & w17037;
assign w30848 = w16851 & ~w17053;
assign w30849 = (~w27596 & w16564) | (~w27596 & w35079) | (w16564 & w35079);
assign w30850 = w2152 & b_50;
assign w30851 = ~w17059 & ~w2161;
assign w30852 = ~w17063 & ~w17064;
assign w30853 = ~a_26 & ~w17064;
assign w30854 = ~a_26 & w30852;
assign w30855 = w35080 & w16834;
assign w30856 = w16784 & ~w16546;
assign w30857 = w1289 & b_56;
assign w30858 = ~w17080 & ~w1298;
assign w30859 = ~w17084 & ~w17085;
assign w30860 = ~a_20 & ~w17085;
assign w30861 = ~a_20 & w30859;
assign w30862 = ~w17088 & w16546;
assign w30863 = (~w17088 & w16546) | (~w17088 & w35081) | (w16546 & w35081);
assign w30864 = w16821 & ~w17096;
assign w30865 = ~w16211 & w35082;
assign w30866 = w651 & b_62;
assign w30867 = (w9770 & w35083) | (w9770 & w35084) | (w35083 & w35084);
assign w30868 = w17105 & w35085;
assign w30869 = (~a_14 & ~w17105) | (~a_14 & w35086) | (~w17105 & w35086);
assign w30870 = w17101 & ~w17109;
assign w30871 = ~w17101 & ~w17109;
assign w30872 = (w27438 & w35087) | (w27438 & w35088) | (w35087 & w35088);
assign w30873 = (w25160 & w25161) | (w25160 & w27757) | (w25161 & w27757);
assign w30874 = (~w27757 & w35089) | (~w27757 & w35090) | (w35089 & w35090);
assign w30875 = ~w17120 & w30794;
assign w30876 = w17100 & ~w17110;
assign w30877 = w651 & b_63;
assign w30878 = ~w660 & ~w17127;
assign w30879 = ~w16819 & w35091;
assign w30880 = (~w17132 & w16819) | (~w17132 & w35092) | (w16819 & w35092);
assign w30881 = w1289 & b_57;
assign w30882 = w17139 & w35093;
assign w30883 = (w17145 & w16834) | (w17145 & w35094) | (w16834 & w35094);
assign w30884 = ~w16834 & w35095;
assign w30885 = w1688 & b_54;
assign w30886 = (a_23 & ~w17152) | (a_23 & w35096) | (~w17152 & w35096);
assign w30887 = a_23 & ~w26375;
assign w30888 = a_23 & ~w30886;
assign w30889 = w26375 & a_23;
assign w30890 = w17057 & ~w17068;
assign w30891 = w2152 & b_51;
assign w30892 = w17166 & w35097;
assign w30893 = (~w16778 & w35098) | (~w16778 & w35099) | (w35098 & w35099);
assign w30894 = (w16778 & w35100) | (w16778 & w35101) | (w35100 & w35101);
assign w30895 = (w16863 & ~w17030) | (w16863 & w35102) | (~w17030 & w35102);
assign w30896 = w3189 & b_45;
assign w30897 = ~w17176 & ~w3198;
assign w30898 = w3797 & b_42;
assign w30899 = w17191 & w35103;
assign w30900 = w16875 & ~w17023;
assign w30901 = w4493 & b_39;
assign w30902 = w17202 & w35104;
assign w30903 = w16886 & ~w17015;
assign w30904 = w16908 & ~w17001;
assign w30905 = w16979 & ~w16968;
assign w30906 = w8520 & b_24;
assign w30907 = w17215 & w35105;
assign w30908 = w16961 & ~w16950;
assign w30909 = w35106 & w16924;
assign w30910 = a_63 & b_13;
assign w30911 = w11614 & b_15;
assign w30912 = ~w17231 & ~w11623;
assign w30913 = ~w17235 & ~w17236;
assign w30914 = ~a_62 & ~w17236;
assign w30915 = (w1038 & w35107) | (w1038 & w35108) | (w35107 & w35108);
assign w30916 = (~w1038 & w35109) | (~w1038 & w35110) | (w35109 & w35110);
assign w30917 = w10556 & b_18;
assign w30918 = w17247 & w35111;
assign w30919 = (w16943 & w16930) | (w16943 & w35112) | (w16930 & w35112);
assign w30920 = w9528 & b_21;
assign w30921 = w17265 & w35113;
assign w30922 = w7607 & b_27;
assign w30923 = w17287 & w35114;
assign w30924 = (w16997 & w16983) | (w16997 & w35115) | (w16983 & w35115);
assign w30925 = w6755 & b_30;
assign w30926 = w17306 & w35116;
assign w30927 = w5956 & b_33;
assign w30928 = w17322 & w35117;
assign w30929 = (w16898 & ~w17008) | (w16898 & w35118) | (~w17008 & w35118);
assign w30930 = w5190 & b_36;
assign w30931 = w17340 & w35119;
assign w30932 = ~w17047 & ~w17049;
assign w30933 = ~w17035 & w35120;
assign w30934 = w2633 & b_48;
assign w30935 = ~w17368 & ~w2642;
assign w30936 = ~w17389 & ~w17388;
assign w30937 = w980 & b_60;
assign w30938 = ~w17395 & ~w989;
assign w30939 = ~w17399 & ~w17400;
assign w30940 = ~a_17 & ~w17400;
assign w30941 = ~a_17 & w30939;
assign w30942 = (w16786 & w35121) | (w16786 & w35122) | (w35121 & w35122);
assign w30943 = ~w17403 & ~w27776;
assign w30944 = ~w17391 & w35123;
assign w30945 = w17135 & w17411;
assign w30946 = ~w17135 & ~w17411;
assign w30947 = (w27757 & w35124) | (w27757 & w35125) | (w35124 & w35125);
assign w30948 = (w27438 & w35126) | (w27438 & w35127) | (w35126 & w35127);
assign w30949 = (~w27757 & w35128) | (~w27757 & w35129) | (w35128 & w35129);
assign w30950 = (~w27438 & w35130) | (~w27438 & w35131) | (w35130 & w35131);
assign w30951 = w17393 & ~w17404;
assign w30952 = w980 & b_61;
assign w30953 = w17425 & w35132;
assign w30954 = ~w17431 & w17404;
assign w30955 = ~w17431 & ~w30951;
assign w30956 = w1289 & b_58;
assign w30957 = w17439 & w35133;
assign w30958 = (~w17075 & w35134) | (~w17075 & w35135) | (w35134 & w35135);
assign w30959 = w17387 & ~w17161;
assign w30960 = w1688 & b_55;
assign w30961 = w17454 & w35136;
assign w30962 = w2152 & b_52;
assign w30963 = w17467 & w35137;
assign w30964 = (~w17054 & w35138) | (~w17054 & w35139) | (w35138 & w35139);
assign w30965 = (w17054 & w35140) | (w17054 & w35141) | (w35140 & w35141);
assign w30966 = w2633 & b_49;
assign w30967 = (a_29 & ~w17480) | (a_29 & w35142) | (~w17480 & w35142);
assign w30968 = a_29 & ~w27604;
assign w30969 = a_29 & ~w30967;
assign w30970 = w27604 & a_29;
assign w30971 = ~w17377 & w17366;
assign w30972 = w17208 & ~w17350;
assign w30973 = (w17346 & w17332) | (w17346 & w35143) | (w17332 & w35143);
assign w30974 = w17328 & ~w17317;
assign w30975 = w17312 & ~w17299;
assign w30976 = a_63 & b_14;
assign w30977 = w17500 & ~w16912;
assign w30978 = w11614 & b_16;
assign w30979 = w17510 & w35144;
assign w30980 = w35145 & w17512;
assign w30981 = w10556 & b_19;
assign w30982 = w17528 & w35146;
assign w30983 = w17253 & ~w17241;
assign w30984 = ~w17537 & w17538;
assign w30985 = w17537 & ~w17538;
assign w30986 = w9528 & b_22;
assign w30987 = w17545 & w35147;
assign w30988 = ~w17553 & ~w17552;
assign w30989 = w8520 & b_25;
assign w30990 = w17562 & w35148;
assign w30991 = w17221 & ~w17275;
assign w30992 = ~w17571 & w17572;
assign w30993 = w17571 & ~w17572;
assign w30994 = w7607 & b_28;
assign w30995 = w17579 & w35149;
assign w30996 = (w17293 & w17211) | (w17293 & w35150) | (w17211 & w35150);
assign w30997 = ~w17588 & w17589;
assign w30998 = w17588 & ~w17589;
assign w30999 = w6755 & b_31;
assign w31000 = w17596 & w35151;
assign w31001 = w5956 & b_34;
assign w31002 = w17613 & w35152;
assign w31003 = w5190 & b_37;
assign w31004 = w17629 & w35153;
assign w31005 = w4493 & b_40;
assign w31006 = w17646 & w35154;
assign w31007 = w3797 & b_43;
assign w31008 = a_35 & ~w27605;
assign w31009 = w26691 & a_35;
assign w31010 = w17197 & ~w17356;
assign w31011 = w3189 & b_46;
assign w31012 = a_32 & ~w26377;
assign w31013 = w25998 & a_32;
assign w31014 = (~w17676 & ~w17677) | (~w17676 & w35155) | (~w17677 & w35155);
assign w31015 = ~w17691 & ~w17690;
assign w31016 = ~w17697 & ~w17696;
assign w31017 = ~w17703 & ~w17702;
assign w31018 = (~w17415 & w25164) | (~w17415 & w27775) | (w25164 & w27775);
assign w31019 = (w27757 & w35157) | (w27757 & w35158) | (w35157 & w35158);
assign w31020 = (w27438 & w35159) | (w27438 & w35160) | (w35159 & w35160);
assign w31021 = (~w27438 & w35161) | (~w27438 & w35162) | (w35161 & w35162);
assign w31022 = ~w17711 & w31018;
assign w31023 = (w17701 & w17446) | (w17701 & w35163) | (w17446 & w35163);
assign w31024 = w980 & b_62;
assign w31025 = (w9770 & w35164) | (w9770 & w35165) | (w35164 & w35165);
assign w31026 = w17718 & w35166;
assign w31027 = (~a_17 & ~w17718) | (~a_17 & w35167) | (~w17718 & w35167);
assign w31028 = w1289 & b_59;
assign w31029 = w17729 & w35168;
assign w31030 = (~w31016 & w17450) | (~w31016 & w35169) | (w17450 & w35169);
assign w31031 = w1688 & b_56;
assign w31032 = ~w17740 & ~w1697;
assign w31033 = ~w17744 & ~w17745;
assign w31034 = ~a_23 & ~w17745;
assign w31035 = ~a_23 & w31033;
assign w31036 = (w17384 & w35170) | (w17384 & w35171) | (w35170 & w35171);
assign w31037 = (~w17384 & w35172) | (~w17384 & w35173) | (w35172 & w35173);
assign w31038 = w2152 & b_53;
assign w31039 = w17755 & w35174;
assign w31040 = ~w31015 & ~w17489;
assign w31041 = w2633 & b_50;
assign w31042 = (~w17775 & w17677) | (~w17775 & w35176) | (w17677 & w35176);
assign w31043 = ~w17677 & w35177;
assign w31044 = w3189 & b_47;
assign w31045 = w17673 & ~w17669;
assign w31046 = w4493 & b_41;
assign w31047 = w17796 & w35178;
assign w31048 = w5190 & b_38;
assign w31049 = w17808 & w35179;
assign w31050 = w5956 & b_35;
assign w31051 = w17819 & w35180;
assign w31052 = w7607 & b_29;
assign w31053 = w17831 & w35181;
assign w31054 = w17521 & ~w17517;
assign w31055 = a_63 & b_15;
assign w31056 = ~w17499 & ~w17840;
assign w31057 = w17499 & w17840;
assign w31058 = w11614 & b_17;
assign w31059 = ~w17844 & ~w11623;
assign w31060 = ~w17848 & ~w17849;
assign w31061 = ~a_62 & ~w17849;
assign w31062 = ~a_62 & w31060;
assign w31063 = (w1372 & w35182) | (w1372 & w35183) | (w35182 & w35183);
assign w31064 = (~w1372 & w35184) | (~w1372 & w35185) | (w35184 & w35185);
assign w31065 = w17853 & w17517;
assign w31066 = w17853 & ~w31054;
assign w31067 = ~w17853 & ~w17517;
assign w31068 = ~w17853 & w31054;
assign w31069 = w10556 & b_20;
assign w31070 = w17860 & w35186;
assign w31071 = w9528 & b_23;
assign w31072 = w17878 & w35187;
assign w31073 = w8520 & b_26;
assign w31074 = w17895 & w35188;
assign w31075 = w6755 & b_32;
assign w31076 = w17920 & w35189;
assign w31077 = ~w17929 & w17825;
assign w31078 = w17939 & ~w17814;
assign w31079 = w17814 & ~w17939;
assign w31080 = w3797 & b_44;
assign w31081 = w17958 & w35190;
assign w31082 = ~w17976 & ~w17975;
assign w31083 = ~w31082 & ~w17976;
assign w31084 = ~w17983 & ~w17982;
assign w31085 = ~w31017 & ~w17432;
assign w31086 = (~w27757 & w35191) | (~w27757 & w35192) | (w35191 & w35192);
assign w31087 = (~w27438 & w35193) | (~w27438 & w35194) | (w35193 & w35194);
assign w31088 = ~w17990 & w31087;
assign w31089 = (~w27757 & w35195) | (~w27757 & w35196) | (w35195 & w35196);
assign w31090 = (~w27438 & w35197) | (~w27438 & w35198) | (w35197 & w35198);
assign w31091 = (~w31084 & w17715) | (~w31084 & w35200) | (w17715 & w35200);
assign w31092 = w17981 & ~w17738;
assign w31093 = w980 & b_63;
assign w31094 = ~w989 & ~w17996;
assign w31095 = w1289 & b_60;
assign w31096 = w18008 & w35201;
assign w31097 = ~w31082 & ~w17749;
assign w31098 = w1688 & b_57;
assign w31099 = w18022 & w35202;
assign w31100 = w17974 & ~w17764;
assign w31101 = w2152 & b_54;
assign w31102 = (a_26 & ~w18037) | (a_26 & w35203) | (~w18037 & w35203);
assign w31103 = a_26 & ~w26385;
assign w31104 = a_26 & ~w31102;
assign w31105 = w26385 & a_26;
assign w31106 = (~w17690 & w35204) | (~w17690 & w35205) | (w35204 & w35205);
assign w31107 = (w17690 & w35206) | (w17690 & w35207) | (w35206 & w35207);
assign w31108 = w2633 & b_51;
assign w31109 = a_29 & ~w26386;
assign w31110 = w26002 & a_29;
assign w31111 = ~w17789 & w35208;
assign w31112 = ~w18056 & w17792;
assign w31113 = w3189 & b_48;
assign w31114 = a_32 & ~w27612;
assign w31115 = w26388 & a_32;
assign w31116 = (w17964 & w17950) | (w17964 & w35209) | (w17950 & w35209);
assign w31117 = w17802 & ~w17944;
assign w31118 = w4493 & b_42;
assign w31119 = w18079 & w35210;
assign w31120 = w5190 & b_39;
assign w31121 = w18090 & w35211;
assign w31122 = w17825 & ~w17930;
assign w31123 = (w17884 & w17871) | (w17884 & w35212) | (w17871 & w35212);
assign w31124 = w9528 & b_24;
assign w31125 = w18102 & w35213;
assign w31126 = w17866 & ~w17854;
assign w31127 = w11614 & b_18;
assign w31128 = w18113 & w35214;
assign w31129 = a_63 & b_16;
assign w31130 = w35215 & w18115;
assign w31131 = w18123 & ~w18124;
assign w31132 = ~w18123 & ~w18124;
assign w31133 = ~w18123 & w31131;
assign w31134 = (w18125 & w35216) | (w18125 & w35217) | (w35216 & w35217);
assign w31135 = (~w18125 & w35218) | (~w18125 & w35219) | (w35218 & w35219);
assign w31136 = w10556 & b_21;
assign w31137 = w18136 & w35220;
assign w31138 = w8520 & b_27;
assign w31139 = w18158 & w35221;
assign w31140 = (w17901 & w17888) | (w17901 & w35222) | (w17888 & w35222);
assign w31141 = w7607 & b_30;
assign w31142 = w18178 & w35223;
assign w31143 = w17837 & ~w17906;
assign w31144 = w6755 & b_33;
assign w31145 = w18195 & w35224;
assign w31146 = (w17926 & w17912) | (w17926 & w35225) | (w17912 & w35225);
assign w31147 = w5956 & b_36;
assign w31148 = w18213 & w35226;
assign w31149 = w18209 & w18219;
assign w31150 = ~w18209 & ~w18219;
assign w31151 = w3797 & b_45;
assign w31152 = (a_35 & ~w18241) | (a_35 & w35227) | (~w18241 & w35227);
assign w31153 = a_35 & ~w27614;
assign w31154 = a_35 & ~w31152;
assign w31155 = w27614 & a_35;
assign w31156 = ~w18253 & ~w18252;
assign w31157 = w18031 & ~w18259;
assign w31158 = w18258 & ~w18259;
assign w31159 = ~w18258 & ~w18259;
assign w31160 = ~w18258 & w31158;
assign w31161 = w18004 & w18267;
assign w31162 = ~w18004 & ~w18267;
assign w31163 = (w27438 & w35228) | (w27438 & w35229) | (w35228 & w35229);
assign w31164 = (w27757 & w35230) | (w27757 & w35231) | (w35230 & w35231);
assign w31165 = (~w27757 & w35232) | (~w27757 & w35233) | (w35232 & w35233);
assign w31166 = ~w18273 & w31090;
assign w31167 = (~w27438 & w35234) | (~w27438 & w35235) | (w35234 & w35235);
assign w31168 = ~w18018 & ~w18017;
assign w31169 = w1289 & b_61;
assign w31170 = w18283 & w35237;
assign w31171 = w1688 & b_58;
assign w31172 = w18296 & w35238;
assign w31173 = (w18302 & w18029) | (w18302 & w35239) | (w18029 & w35239);
assign w31174 = (w18029 & w35240) | (w18029 & w35241) | (w35240 & w35241);
assign w31175 = ~w18029 & w35242;
assign w31176 = (~w18029 & w35243) | (~w18029 & w35244) | (w35243 & w35244);
assign w31177 = w2633 & b_52;
assign w31178 = w18309 & w35245;
assign w31179 = ~w31156 & ~w18058;
assign w31180 = w18315 & ~w18058;
assign w31181 = w18315 & w31179;
assign w31182 = ~w18315 & w18058;
assign w31183 = ~w18315 & ~w31179;
assign w31184 = w18096 & ~w18223;
assign w31185 = w18209 & ~w18219;
assign w31186 = (w18201 & w18187) | (w18201 & w35246) | (w18187 & w35246);
assign w31187 = w9528 & b_25;
assign w31188 = w18326 & w35247;
assign w31189 = (~w18127 & w35248) | (~w18127 & w35249) | (w35248 & w35249);
assign w31190 = w11614 & b_19;
assign w31191 = w18337 & w35250;
assign w31192 = a_63 & b_17;
assign w31193 = w35251 & w18339;
assign w31194 = w10556 & b_22;
assign w31195 = w18363 & w35252;
assign w31196 = ~w18358 & w18369;
assign w31197 = w18358 & ~w18369;
assign w31198 = (w18108 & ~w18145) | (w18108 & w35253) | (~w18145 & w35253);
assign w31199 = ~w18378 & w18379;
assign w31200 = w18378 & ~w18379;
assign w31201 = w8520 & b_28;
assign w31202 = w18386 & w35254;
assign w31203 = w18164 & ~w18152;
assign w31204 = ~w18395 & w18396;
assign w31205 = w18395 & ~w18396;
assign w31206 = w7607 & b_31;
assign w31207 = w18403 & w35255;
assign w31208 = w18184 & ~w18171;
assign w31209 = w18409 & ~w18171;
assign w31210 = ~w18171 & w35256;
assign w31211 = (~w18174 & w35257) | (~w18174 & w35258) | (w35257 & w35258);
assign w31212 = (w18174 & w35259) | (w18174 & w35260) | (w35259 & w35260);
assign w31213 = w6755 & b_34;
assign w31214 = w18417 & w35261;
assign w31215 = w5956 & b_37;
assign w31216 = w18433 & w35262;
assign w31217 = w5190 & b_40;
assign w31218 = w18450 & w35263;
assign w31219 = w4493 & b_43;
assign w31220 = a_38 & ~w27615;
assign w31221 = w26692 & a_38;
assign w31222 = (w18085 & w18086) | (w18085 & w35264) | (w18086 & w35264);
assign w31223 = w3797 & b_46;
assign w31224 = a_35 & ~w27617;
assign w31225 = w26693 & a_35;
assign w31226 = (w18247 & ~w18234) | (w18247 & w35265) | (~w18234 & w35265);
assign w31227 = ~w18493 & w18494;
assign w31228 = w18493 & ~w18494;
assign w31229 = w3189 & b_49;
assign w31230 = w18501 & w35266;
assign w31231 = w18251 & ~w18073;
assign w31232 = w2152 & b_55;
assign w31233 = w18523 & w35267;
assign w31234 = w18292 & w18541;
assign w31235 = ~w18292 & ~w18541;
assign w31236 = w18002 & ~w18544;
assign w31237 = (w27438 & w35268) | (w27438 & w35269) | (w35268 & w35269);
assign w31238 = (w27757 & w35270) | (w27757 & w35271) | (w35270 & w35271);
assign w31239 = (~w27757 & w35272) | (~w27757 & w35273) | (w35272 & w35273);
assign w31240 = ~w18547 & w31167;
assign w31241 = (~w25146 & w37860) | (~w25146 & w37861) | (w37860 & w37861);
assign w31242 = w18292 & ~w18541;
assign w31243 = w1688 & b_59;
assign w31244 = w18557 & w35277;
assign w31245 = w18519 & ~w18531;
assign w31246 = w2152 & b_56;
assign w31247 = w18571 & w35278;
assign w31248 = ~w18317 & w18577;
assign w31249 = w18317 & ~w18577;
assign w31250 = w2633 & b_53;
assign w31251 = w18584 & w35279;
assign w31252 = (~w18497 & w18508) | (~w18497 & w35280) | (w18508 & w35280);
assign w31253 = w3189 & b_50;
assign w31254 = (a_32 & ~w18598) | (a_32 & w35281) | (~w18598 & w35281);
assign w31255 = a_32 & ~w26389;
assign w31256 = a_32 & ~w31254;
assign w31257 = w26389 & a_32;
assign w31258 = (w18604 & ~w18480) | (w18604 & w35282) | (~w18480 & w35282);
assign w31259 = w18480 & w35283;
assign w31260 = w5190 & b_41;
assign w31261 = w18611 & w35284;
assign w31262 = w5956 & b_38;
assign w31263 = w18623 & w35285;
assign w31264 = w18322 & ~w18424;
assign w31265 = w8520 & b_29;
assign w31266 = w18634 & w35286;
assign w31267 = w18333 & ~w18371;
assign w31268 = w10556 & b_23;
assign w31269 = w18645 & w35287;
assign w31270 = a_63 & b_18;
assign w31271 = w18122 & ~w18347;
assign w31272 = w11614 & b_20;
assign w31273 = w18662 & w35288;
assign w31274 = (~w18664 & w35289) | (~w18664 & ~w18658) | (w35289 & ~w18658);
assign w31275 = w35290 & w18664;
assign w31276 = w18128 & ~w18353;
assign w31277 = w9528 & b_26;
assign w31278 = w18684 & w35291;
assign w31279 = w7607 & b_32;
assign w31280 = w18709 & w35292;
assign w31281 = (~w18174 & w35293) | (~w18174 & w35294) | (w35293 & w35294);
assign w31282 = w6755 & b_35;
assign w31283 = w18728 & w35295;
assign w31284 = w18739 & ~w18629;
assign w31285 = w18629 & ~w18739;
assign w31286 = w18319 & ~w18457;
assign w31287 = ~w18749 & w18750;
assign w31288 = w18749 & ~w18750;
assign w31289 = w4493 & b_44;
assign w31290 = (a_38 & ~w18757) | (a_38 & w35296) | (~w18757 & w35296);
assign w31291 = a_38 & ~w27619;
assign w31292 = a_38 & ~w31290;
assign w31293 = w27619 & a_38;
assign w31294 = w18477 & ~w18473;
assign w31295 = w3797 & b_47;
assign w31296 = w18775 & w35297;
assign w31297 = ~w18787 & ~w18786;
assign w31298 = ~w18793 & ~w18792;
assign w31299 = w18537 & ~w18304;
assign w31300 = w1289 & b_62;
assign w31301 = (w9770 & w35298) | (w9770 & w35299) | (w35298 & w35299);
assign w31302 = w18801 & w35300;
assign w31303 = (~a_20 & ~w18801) | (~a_20 & w35301) | (~w18801 & w35301);
assign w31304 = w18808 & ~w18797;
assign w31305 = (w27757 & w35302) | (w27757 & w35303) | (w35302 & w35303);
assign w31306 = (w27438 & w35304) | (w27438 & w35305) | (w35304 & w35305);
assign w31307 = (~w27757 & w35306) | (~w27757 & w35307) | (w35306 & w35307);
assign w31308 = (~w27438 & w35308) | (~w27438 & w35309) | (w35308 & w35309);
assign w31309 = (~w27757 & w35310) | (~w27757 & w35311) | (w35310 & w35311);
assign w31310 = (~w27438 & w35312) | (~w27438 & w35313) | (w35312 & w35313);
assign w31311 = (~w31298 & w18564) | (~w31298 & w35314) | (w18564 & w35314);
assign w31312 = w1289 & b_63;
assign w31313 = ~w1298 & ~w18822;
assign w31314 = w1688 & b_60;
assign w31315 = w18834 & w35315;
assign w31316 = (w18516 & w35316) | (w18516 & w35317) | (w35316 & w35317);
assign w31317 = ~w31316 & ~w18840;
assign w31318 = w2152 & b_57;
assign w31319 = w18849 & w35318;
assign w31320 = (~w31297 & w18591) | (~w31297 & w35319) | (w18591 & w35319);
assign w31321 = w2633 & b_54;
assign w31322 = a_29 & ~w26390;
assign w31323 = w26003 & a_29;
assign w31324 = (w18496 & w35320) | (w18496 & w35321) | (w35320 & w35321);
assign w31325 = (~w18496 & w35322) | (~w18496 & w35323) | (w35322 & w35323);
assign w31326 = w3189 & b_51;
assign w31327 = (a_32 & ~w18878) | (a_32 & w35324) | (~w18878 & w35324);
assign w31328 = a_32 & ~w26392;
assign w31329 = a_32 & ~w31327;
assign w31330 = w26392 & a_32;
assign w31331 = (w18781 & w18767) | (w18781 & w35325) | (w18767 & w35325);
assign w31332 = (w18617 & w18619) | (w18617 & w35326) | (w18619 & w35326);
assign w31333 = w5190 & b_42;
assign w31334 = w18892 & w35327;
assign w31335 = w5956 & b_39;
assign w31336 = w18903 & w35328;
assign w31337 = w18734 & ~w18723;
assign w31338 = w6755 & b_36;
assign w31339 = w18914 & w35329;
assign w31340 = (w18715 & w18701) | (w18715 & w35330) | (w18701 & w35330);
assign w31341 = w7607 & b_33;
assign w31342 = w18925 & w35331;
assign w31343 = w18640 & ~w18695;
assign w31344 = (w18651 & w18670) | (w18651 & w35332) | (w18670 & w35332);
assign w31345 = w10556 & b_24;
assign w31346 = w18937 & w35333;
assign w31347 = a_63 & b_19;
assign w31348 = w11614 & b_21;
assign w31349 = ~w18951 & ~w11623;
assign w31350 = ~w18955 & ~w18956;
assign w31351 = ~a_62 & ~w18956;
assign w31352 = (w1933 & w35334) | (w1933 & w35335) | (w35334 & w35335);
assign w31353 = (~w1933 & w35336) | (~w1933 & w35337) | (w35336 & w35337);
assign w31354 = w9528 & b_27;
assign w31355 = w18973 & w35338;
assign w31356 = (w18690 & w18677) | (w18690 & w35339) | (w18677 & w35339);
assign w31357 = w8520 & b_30;
assign w31358 = w18993 & w35340;
assign w31359 = w4493 & b_45;
assign w31360 = (a_38 & ~w19033) | (a_38 & w35341) | (~w19033 & w35341);
assign w31361 = a_38 & ~w27620;
assign w31362 = a_38 & ~w31360;
assign w31363 = w27620 & a_38;
assign w31364 = w18763 & ~w18752;
assign w31365 = w3797 & b_48;
assign w31366 = w19051 & w35342;
assign w31367 = ~w19059 & ~w19058;
assign w31368 = w18830 & ~w19073;
assign w31369 = ~w18830 & w19073;
assign w31370 = (w27757 & w35343) | (w27757 & w35344) | (w35343 & w35344);
assign w31371 = (w27438 & w35345) | (w27438 & w35346) | (w35345 & w35346);
assign w31372 = w19070 & ~w18842;
assign w31373 = w1688 & b_61;
assign w31374 = w19087 & w35347;
assign w31375 = w2152 & b_58;
assign w31376 = w19101 & w35348;
assign w31377 = w19066 & ~w18858;
assign w31378 = w19063 & ~w18871;
assign w31379 = w2633 & b_55;
assign w31380 = w19116 & w35349;
assign w31381 = w3189 & b_52;
assign w31382 = w19129 & w35350;
assign w31383 = ~w31367 & ~w18886;
assign w31384 = (w19057 & w19043) | (w19057 & w35351) | (w19043 & w35351);
assign w31385 = (w18931 & w19002) | (w18931 & w35352) | (w19002 & w35352);
assign w31386 = a_63 & b_20;
assign w31387 = w11614 & b_22;
assign w31388 = w19154 & w35353;
assign w31389 = w35354 & w19156;
assign w31390 = w10556 & b_25;
assign w31391 = w19173 & w35355;
assign w31392 = w35356 & w19164;
assign w31393 = w18943 & ~w18961;
assign w31394 = w9528 & b_28;
assign w31395 = w19191 & w35357;
assign w31396 = (w18979 & w18933) | (w18979 & w35358) | (w18933 & w35358);
assign w31397 = (w19187 & w35359) | (w19187 & w35360) | (w35359 & w35360);
assign w31398 = w35361 & ~w19187;
assign w31399 = w8520 & b_31;
assign w31400 = w19207 & w35362;
assign w31401 = w18999 & ~w18986;
assign w31402 = w19213 & ~w18986;
assign w31403 = ~w18986 & w35363;
assign w31404 = ~w19216 & ~w19203;
assign w31405 = w19216 & w19203;
assign w31406 = w7607 & b_34;
assign w31407 = w19223 & w35364;
assign w31408 = w6755 & b_37;
assign w31409 = w19239 & w35365;
assign w31410 = w18920 & ~w19009;
assign w31411 = ~w19248 & w19249;
assign w31412 = w19248 & ~w19249;
assign w31413 = w5956 & b_40;
assign w31414 = w19256 & w35366;
assign w31415 = (w18909 & w18910) | (w18909 & w35367) | (w18910 & w35367);
assign w31416 = w5190 & b_43;
assign w31417 = (a_41 & ~w19274) | (a_41 & w35368) | (~w19274 & w35368);
assign w31418 = a_41 & ~w27621;
assign w31419 = a_41 & ~w31417;
assign w31420 = w27621 & a_41;
assign w31421 = (w18898 & w18899) | (w18898 & w35369) | (w18899 & w35369);
assign w31422 = w4493 & b_46;
assign w31423 = (a_38 & ~w19292) | (a_38 & w35370) | (~w19292 & w35370);
assign w31424 = a_38 & ~w27622;
assign w31425 = a_38 & ~w31423;
assign w31426 = w27622 & a_38;
assign w31427 = w19039 & ~w19027;
assign w31428 = ~w19301 & w19302;
assign w31429 = w19301 & ~w19302;
assign w31430 = w3797 & b_49;
assign w31431 = w19309 & w35371;
assign w31432 = ~w19317 & ~w19316;
assign w31433 = ~w19323 & ~w19322;
assign w31434 = w19096 & ~w19329;
assign w31435 = w19328 & ~w19329;
assign w31436 = ~w19328 & ~w19329;
assign w31437 = ~w19328 & w31435;
assign w31438 = (~w27757 & w35372) | (~w27757 & w35373) | (w35372 & w35373);
assign w31439 = (~w27438 & w35374) | (~w27438 & w35375) | (w35374 & w35375);
assign w31440 = (w27757 & w35376) | (w27757 & w35377) | (w35376 & w35377);
assign w31441 = (w27438 & w35378) | (w27438 & w35379) | (w35378 & w35379);
assign w31442 = w19327 & ~w19110;
assign w31443 = w1688 & b_62;
assign w31444 = (w9770 & w35380) | (w9770 & w35381) | (w35380 & w35381);
assign w31445 = w19345 & w35382;
assign w31446 = (~a_23 & ~w19345) | (~a_23 & w35383) | (~w19345 & w35383);
assign w31447 = w2152 & b_59;
assign w31448 = w19356 & w35384;
assign w31449 = ~w31433 & ~w19363;
assign w31450 = (w19321 & w19136) | (w19321 & w35385) | (w19136 & w35385);
assign w31451 = w2633 & b_56;
assign w31452 = ~w19369 & ~w2642;
assign w31453 = ~w19373 & ~w19374;
assign w31454 = ~a_29 & ~w19374;
assign w31455 = ~a_29 & w31453;
assign w31456 = w3189 & b_53;
assign w31457 = w19384 & w35386;
assign w31458 = w19305 & w35387;
assign w31459 = (~w19390 & ~w19305) | (~w19390 & w35388) | (~w19305 & w35388);
assign w31460 = w5956 & b_41;
assign w31461 = w19397 & w35389;
assign w31462 = w6755 & b_38;
assign w31463 = w19408 & w35390;
assign w31464 = w19141 & ~w19230;
assign w31465 = (~w19167 & w35391) | (~w19167 & w35392) | (w35391 & w35392);
assign w31466 = w10556 & b_26;
assign w31467 = w19419 & w35393;
assign w31468 = w19165 & ~w19161;
assign w31469 = a_63 & b_21;
assign w31470 = w18947 & ~w19145;
assign w31471 = w11614 & b_23;
assign w31472 = ~w19433 & ~w11623;
assign w31473 = ~w19437 & ~w19438;
assign w31474 = ~a_62 & ~w19438;
assign w31475 = ~a_62 & w31473;
assign w31476 = (w2108 & w35394) | (w2108 & w35395) | (w35394 & w35395);
assign w31477 = (~w2108 & w35396) | (~w2108 & w35397) | (w35396 & w35397);
assign w31478 = w19442 & w19161;
assign w31479 = w19442 & ~w31468;
assign w31480 = ~w19442 & ~w19161;
assign w31481 = ~w19442 & w31468;
assign w31482 = w19448 & w19180;
assign w31483 = w19448 & ~w31465;
assign w31484 = ~w19448 & ~w19180;
assign w31485 = ~w19448 & w31465;
assign w31486 = w9528 & b_29;
assign w31487 = w19455 & w35398;
assign w31488 = w8520 & b_32;
assign w31489 = w19473 & w35399;
assign w31490 = ~w19216 & w19203;
assign w31491 = w7607 & b_35;
assign w31492 = w19492 & w35400;
assign w31493 = w35401 & ~w19501;
assign w31494 = (w19501 & w35402) | (w19501 & w19414) | (w35402 & w19414);
assign w31495 = w19267 & ~w19263;
assign w31496 = ~w19512 & w19513;
assign w31497 = w19512 & ~w19513;
assign w31498 = w5190 & b_44;
assign w31499 = (a_41 & ~w19520) | (a_41 & w35403) | (~w19520 & w35403);
assign w31500 = a_41 & ~w27623;
assign w31501 = a_41 & ~w31499;
assign w31502 = w27623 & a_41;
assign w31503 = w19285 & ~w19281;
assign w31504 = w4493 & b_47;
assign w31505 = w19538 & w35404;
assign w31506 = w3797 & b_50;
assign w31507 = w19556 & w35405;
assign w31508 = ~w19568 & ~w19567;
assign w31509 = ~w19574 & ~w19573;
assign w31510 = w19328 & ~w19094;
assign w31511 = (~w27757 & w35406) | (~w27757 & w35407) | (w35406 & w35407);
assign w31512 = (~w27438 & w35408) | (~w27438 & w35409) | (w35408 & w35409);
assign w31513 = (w27757 & w35410) | (w27757 & w35411) | (w35410 & w35411);
assign w31514 = (w27438 & w35412) | (w27438 & w35413) | (w35412 & w35413);
assign w31515 = (~w27757 & w35415) | (~w27757 & w35416) | (w35415 & w35416);
assign w31516 = ~w31509 & ~w19350;
assign w31517 = w19572 & ~w19366;
assign w31518 = w1688 & b_63;
assign w31519 = ~w1697 & ~w19588;
assign w31520 = w2152 & b_60;
assign w31521 = w19600 & w35417;
assign w31522 = (~w31508 & w19368) | (~w31508 & w35418) | (w19368 & w35418);
assign w31523 = w2633 & b_57;
assign w31524 = w19614 & w35419;
assign w31525 = w19305 & w35420;
assign w31526 = (w19318 & w35421) | (w19318 & w35422) | (w35421 & w35422);
assign w31527 = (~w19318 & w35423) | (~w19318 & w35424) | (w35423 & w35424);
assign w31528 = w3189 & b_54;
assign w31529 = (a_32 & ~w19630) | (a_32 & w35425) | (~w19630 & w35425);
assign w31530 = a_32 & ~w26393;
assign w31531 = a_32 & ~w31529;
assign w31532 = w26393 & a_32;
assign w31533 = (w19562 & w19548) | (w19562 & w35426) | (w19548 & w35426);
assign w31534 = w3797 & b_51;
assign w31535 = w19643 & w35427;
assign w31536 = (w19544 & w19530) | (w19544 & w35428) | (w19530 & w35428);
assign w31537 = (w19403 & ~w19506) | (w19403 & w35429) | (~w19506 & w35429);
assign w31538 = w5956 & b_42;
assign w31539 = w19655 & w35430;
assign w31540 = (w19479 & w19466) | (w19479 & w35431) | (w19466 & w35431);
assign w31541 = w8520 & b_33;
assign w31542 = w19667 & w35432;
assign w31543 = w19461 & ~w19449;
assign w31544 = a_63 & b_22;
assign w31545 = w11614 & b_24;
assign w31546 = ~w19682 & ~w11623;
assign w31547 = ~w19686 & ~w19687;
assign w31548 = ~a_62 & ~w19687;
assign w31549 = (w2416 & w35433) | (w2416 & w35434) | (w35433 & w35434);
assign w31550 = (~w2416 & w35435) | (~w2416 & w35436) | (w35435 & w35436);
assign w31551 = w10556 & b_27;
assign w31552 = w19698 & w35437;
assign w31553 = w19425 & ~w19443;
assign w31554 = w9528 & b_30;
assign w31555 = w19716 & w35438;
assign w31556 = w7607 & b_36;
assign w31557 = w19738 & w35439;
assign w31558 = (w19498 & w19483) | (w19498 & w35440) | (w19483 & w35440);
assign w31559 = w6755 & b_39;
assign w31560 = w19757 & w35441;
assign w31561 = w5190 & b_45;
assign w31562 = a_41 & ~w27624;
assign w31563 = w26694 & a_41;
assign w31564 = w19526 & ~w19515;
assign w31565 = ~w19788 & w19789;
assign w31566 = w19788 & ~w19789;
assign w31567 = w4493 & b_48;
assign w31568 = w19796 & w35442;
assign w31569 = w19596 & w19824;
assign w31570 = ~w19596 & ~w19824;
assign w31571 = (w27757 & w35443) | (w27757 & w35444) | (w35443 & w35444);
assign w31572 = (w27438 & w35445) | (w27438 & w35446) | (w35445 & w35446);
assign w31573 = (~w27757 & w35447) | (~w27757 & w35448) | (w35447 & w35448);
assign w31574 = (~w27438 & w35449) | (~w27438 & w35450) | (w35449 & w35450);
assign w31575 = w19596 & ~w19824;
assign w31576 = w19820 & ~w19609;
assign w31577 = w2152 & b_61;
assign w31578 = w19841 & w35451;
assign w31579 = w19817 & ~w19623;
assign w31580 = w2633 & b_58;
assign w31581 = w19855 & w35452;
assign w31582 = w3189 & b_55;
assign w31583 = w19868 & w35453;
assign w31584 = w19813 & ~w19638;
assign w31585 = w19649 & ~w19806;
assign w31586 = w19802 & ~w19791;
assign w31587 = w19661 & ~w19767;
assign w31588 = w19763 & ~w19750;
assign w31589 = w8520 & b_34;
assign w31590 = w19886 & w35454;
assign w31591 = w19704 & ~w19692;
assign w31592 = a_63 & b_23;
assign w31593 = w11614 & b_25;
assign w31594 = w19907 & w35455;
assign w31595 = w35456 & w19909;
assign w31596 = w10556 & b_28;
assign w31597 = w19924 & w35457;
assign w31598 = w9528 & b_31;
assign w31599 = w19940 & w35458;
assign w31600 = w19722 & ~w19711;
assign w31601 = (w19673 & w19674) | (w19673 & w35459) | (w19674 & w35459);
assign w31602 = ~w19956 & w19957;
assign w31603 = w19956 & ~w19957;
assign w31604 = w7607 & b_37;
assign w31605 = (a_50 & ~w19964) | (a_50 & w35460) | (~w19964 & w35460);
assign w31606 = a_50 & ~w27626;
assign w31607 = a_50 & ~w31605;
assign w31608 = w27626 & a_50;
assign w31609 = (w19744 & w19663) | (w19744 & w35461) | (w19663 & w35461);
assign w31610 = w6755 & b_40;
assign w31611 = a_47 & ~w27627;
assign w31612 = w26695 & a_47;
assign w31613 = w5956 & b_43;
assign w31614 = a_44 & ~w27629;
assign w31615 = w26696 & a_44;
assign w31616 = w5190 & b_46;
assign w31617 = (w19785 & ~w19772) | (w19785 & w35462) | (~w19772 & w35462);
assign w31618 = w4493 & b_49;
assign w31619 = w20032 & w35463;
assign w31620 = ~w20027 & ~w20038;
assign w31621 = w20027 & w20038;
assign w31622 = ~w20040 & ~w20039;
assign w31623 = w3797 & b_52;
assign w31624 = w20049 & w35464;
assign w31625 = ~w20063 & ~w20062;
assign w31626 = w19850 & w20067;
assign w31627 = ~w19850 & ~w20067;
assign w31628 = (w27757 & w35465) | (w27757 & w35466) | (w35465 & w35466);
assign w31629 = (w27438 & w35467) | (w27438 & w35468) | (w35467 & w35468);
assign w31630 = (~w27757 & w35469) | (~w27757 & w35470) | (w35469 & w35470);
assign w31631 = (~w27438 & w35471) | (~w27438 & w35472) | (w35471 & w35472);
assign w31632 = w19850 & ~w20067;
assign w31633 = w2633 & b_59;
assign w31634 = w20083 & w35473;
assign w31635 = (~w20061 & w19875) | (~w20061 & w35474) | (w19875 & w35474);
assign w31636 = w3189 & b_56;
assign w31637 = ~w20095 & ~w3198;
assign w31638 = ~w20099 & ~w20100;
assign w31639 = ~a_32 & ~w20100;
assign w31640 = ~a_32 & w31638;
assign w31641 = ~w20045 & w35475;
assign w31642 = (w20103 & w20045) | (w20103 & w35476) | (w20045 & w35476);
assign w31643 = w6755 & b_41;
assign w31644 = a_47 & ~w27634;
assign w31645 = w26699 & a_47;
assign w31646 = w7607 & b_38;
assign w31647 = (a_50 & ~w20121) | (a_50 & w35477) | (~w20121 & w35477);
assign w31648 = a_50 & ~w27636;
assign w31649 = a_50 & ~w31647;
assign w31650 = w27636 & a_50;
assign w31651 = w19894 & ~w19914;
assign w31652 = w19678 & ~w19898;
assign w31653 = w11614 & b_26;
assign w31654 = ~w20136 & ~w11623;
assign w31655 = ~w20140 & ~w20141;
assign w31656 = ~a_62 & ~w20141;
assign w31657 = ~a_62 & w31655;
assign w31658 = (w2771 & w35478) | (w2771 & w35479) | (w35478 & w35479);
assign w31659 = (~w2771 & w35480) | (~w2771 & w35481) | (w35480 & w35481);
assign w31660 = w20145 & w19914;
assign w31661 = w20145 & ~w31651;
assign w31662 = ~w20145 & ~w19914;
assign w31663 = ~w20145 & w31651;
assign w31664 = w10556 & b_29;
assign w31665 = w20152 & w35482;
assign w31666 = (w19893 & w19920) | (w19893 & w35483) | (w19920 & w35483);
assign w31667 = w9528 & b_32;
assign w31668 = w20170 & w35484;
assign w31669 = ~w19936 & ~w19948;
assign w31670 = w8520 & b_35;
assign w31671 = w20188 & w35485;
assign w31672 = ~w20197 & w20127;
assign w31673 = ~w19990 & w35486;
assign w31674 = w5956 & b_44;
assign w31675 = w5190 & b_47;
assign w31676 = a_41 & ~w27639;
assign w31677 = w26396 & a_41;
assign w31678 = ~w20022 & ~w20024;
assign w31679 = ~w20022 & w20026;
assign w31680 = w4493 & b_50;
assign w31681 = w20256 & w35487;
assign w31682 = ~w20265 & ~w20043;
assign w31683 = w20265 & w20043;
assign w31684 = w3797 & b_53;
assign w31685 = w20272 & w35488;
assign w31686 = w35489 & w20090;
assign w31687 = ~w31625 & ~w20289;
assign w31688 = w2152 & b_62;
assign w31689 = (w9770 & w35490) | (w9770 & w35491) | (w35490 & w35491);
assign w31690 = w20293 & w35492;
assign w31691 = (~a_26 & ~w20293) | (~a_26 & w35493) | (~w20293 & w35493);
assign w31692 = w20300 & ~w20288;
assign w31693 = (w27757 & w35494) | (w27757 & w35495) | (w35494 & w35495);
assign w31694 = (w27438 & w35496) | (w27438 & w35497) | (w35496 & w35497);
assign w31695 = (~w27757 & w35498) | (~w27757 & w35499) | (w35498 & w35499);
assign w31696 = (~w27438 & w35500) | (~w27438 & w35501) | (w35500 & w35501);
assign w31697 = (~w27757 & w35502) | (~w27757 & w35503) | (w35502 & w35503);
assign w31698 = (~w27438 & w35504) | (~w27438 & w35505) | (w35504 & w35505);
assign w31699 = w2152 & b_63;
assign w31700 = ~w2161 & ~w20313;
assign w31701 = ~w20090 & w35506;
assign w31702 = (~w20318 & w20090) | (~w20318 & w35507) | (w20090 & w35507);
assign w31703 = w2633 & b_60;
assign w31704 = w20324 & w35508;
assign w31705 = ~w20281 & ~w20104;
assign w31706 = w3189 & b_57;
assign w31707 = w20338 & w35509;
assign w31708 = w20265 & ~w20043;
assign w31709 = w3797 & b_54;
assign w31710 = w20353 & w35510;
assign w31711 = (w20262 & w20248) | (w20262 & w35511) | (w20248 & w35511);
assign w31712 = w4493 & b_51;
assign w31713 = w20364 & w35512;
assign w31714 = (w20244 & w20231) | (w20244 & w35513) | (w20231 & w35513);
assign w31715 = w20116 & ~w20206;
assign w31716 = w6755 & b_42;
assign w31717 = (a_47 & ~w20376) | (a_47 & w35514) | (~w20376 & w35514);
assign w31718 = a_47 & ~w26397;
assign w31719 = a_47 & ~w31717;
assign w31720 = w26397 & a_47;
assign w31721 = w20127 & ~w20198;
assign w31722 = w20176 & ~w20165;
assign w31723 = w9528 & b_33;
assign w31724 = w20388 & w35515;
assign w31725 = w20158 & ~w20146;
assign w31726 = w10556 & b_30;
assign w31727 = w20399 & w35516;
assign w31728 = a_63 & b_25;
assign w31729 = w11614 & b_27;
assign w31730 = ~w20413 & ~w11623;
assign w31731 = ~w20417 & ~w20418;
assign w31732 = ~a_62 & ~w20418;
assign w31733 = ~a_62 & w31731;
assign w31734 = (w2954 & w35517) | (w2954 & w35518) | (w35517 & w35518);
assign w31735 = (~w2954 & w35519) | (~w2954 & w35520) | (w35519 & w35520);
assign w31736 = w8520 & b_36;
assign w31737 = w20441 & w35521;
assign w31738 = (w20194 & w20180) | (w20194 & w35522) | (w20180 & w35522);
assign w31739 = w7607 & b_39;
assign w31740 = w20460 & w35523;
assign w31741 = w5956 & b_45;
assign w31742 = ~w20489 & ~w20490;
assign w31743 = w5190 & b_48;
assign w31744 = (a_41 & ~w20498) | (a_41 & w35524) | (~w20498 & w35524);
assign w31745 = a_41 & ~w26401;
assign w31746 = a_41 & ~w31744;
assign w31747 = w26401 & a_41;
assign w31748 = w20491 & w35525;
assign w31749 = (~w20504 & ~w20491) | (~w20504 & w35526) | (~w20491 & w35526);
assign w31750 = ~w20507 & w20370;
assign w31751 = ~w20285 & w35527;
assign w31752 = (~w20529 & w20285) | (~w20529 & w35528) | (w20285 & w35528);
assign w31753 = (w25200 & w25201) | (w25200 & ~w31515) | (w25201 & ~w31515);
assign w31754 = (w27438 & w35529) | (w27438 & w35530) | (w35529 & w35530);
assign w31755 = w2633 & b_61;
assign w31756 = w20543 & w35531;
assign w31757 = ~w20331 & w35532;
assign w31758 = (~w20549 & w20331) | (~w20549 & w35533) | (w20331 & w35533);
assign w31759 = w3797 & b_55;
assign w31760 = w20556 & w35534;
assign w31761 = (w20370 & w20371) | (w20370 & w31750) | (w20371 & w31750);
assign w31762 = w20382 & ~w20470;
assign w31763 = w20466 & ~w20453;
assign w31764 = w10556 & b_31;
assign w31765 = w20570 & w35535;
assign w31766 = w20405 & ~w20423;
assign w31767 = a_63 & b_26;
assign w31768 = w20410 & w20589;
assign w31769 = ~w20410 & ~w20589;
assign w31770 = w11614 & b_28;
assign w31771 = w20596 & w35536;
assign w31772 = w9528 & b_34;
assign w31773 = w20613 & w35537;
assign w31774 = w20394 & ~w20429;
assign w31775 = ~w20622 & w20623;
assign w31776 = w20622 & ~w20623;
assign w31777 = w8520 & b_37;
assign w31778 = w20630 & w35538;
assign w31779 = (w20447 & w20384) | (w20447 & w35539) | (w20384 & w35539);
assign w31780 = ~w20639 & w20640;
assign w31781 = w20639 & ~w20640;
assign w31782 = w7607 & b_40;
assign w31783 = (a_50 & ~w20647) | (a_50 & w35540) | (~w20647 & w35540);
assign w31784 = a_50 & ~w26402;
assign w31785 = a_50 & ~w31783;
assign w31786 = w26402 & a_50;
assign w31787 = w6755 & b_43;
assign w31788 = a_47 & ~w26403;
assign w31789 = w26006 & a_47;
assign w31790 = w5956 & b_46;
assign w31791 = ~w20476 & w20488;
assign w31792 = ~w20688 & ~w20689;
assign w31793 = w5190 & b_49;
assign w31794 = a_41 & ~w26408;
assign w31795 = w26009 & a_41;
assign w31796 = ~w20691 & ~w20702;
assign w31797 = w20691 & w20702;
assign w31798 = w20704 & ~w20703;
assign w31799 = w4493 & b_52;
assign w31800 = w20711 & w35541;
assign w31801 = (~w20564 & w35542) | (~w20564 & w35543) | (w35542 & w35543);
assign w31802 = (w20564 & w35544) | (w20564 & w35545) | (w35544 & w35545);
assign w31803 = w20359 & ~w20516;
assign w31804 = w3189 & b_58;
assign w31805 = w20735 & w35546;
assign w31806 = w20522 & ~w20348;
assign w31807 = w20552 & ~w20748;
assign w31808 = ~w20552 & w20748;
assign w31809 = ~w20319 & ~w20751;
assign w31810 = w20319 & w20751;
assign w31811 = (~w27757 & w35547) | (~w27757 & w35548) | (w35547 & w35548);
assign w31812 = (~w27438 & w35549) | (~w27438 & w35550) | (w35549 & w35550);
assign w31813 = (w27757 & w35551) | (w27757 & w35552) | (w35551 & w35552);
assign w31814 = (w27438 & w35553) | (w27438 & w35554) | (w35553 & w35554);
assign w31815 = (~w20731 & w20742) | (~w20731 & w35555) | (w20742 & w35555);
assign w31816 = ~w20760 & ~w2642;
assign w31817 = (w9770 & w35556) | (w9770 & w35557) | (w35556 & w35557);
assign w31818 = w20762 & a_29;
assign w31819 = ~w20762 & ~a_29;
assign w31820 = w3189 & b_59;
assign w31821 = w20773 & w35558;
assign w31822 = w20728 & ~w20724;
assign w31823 = w3797 & b_56;
assign w31824 = w20787 & w35559;
assign w31825 = w7607 & b_41;
assign w31826 = (a_50 & ~w20798) | (a_50 & w35560) | (~w20798 & w35560);
assign w31827 = a_50 & ~w27644;
assign w31828 = a_50 & ~w31826;
assign w31829 = w27644 & a_50;
assign w31830 = w8520 & b_38;
assign w31831 = w20809 & w35561;
assign w31832 = w10556 & b_32;
assign w31833 = w20820 & w35562;
assign w31834 = a_63 & b_27;
assign w31835 = w20409 & ~w20584;
assign w31836 = w11614 & b_29;
assign w31837 = (a_62 & ~w20837) | (a_62 & w35563) | (~w20837 & w35563);
assign w31838 = a_62 & ~w26703;
assign w31839 = a_62 & ~w31837;
assign w31840 = w26703 & a_62;
assign w31841 = (w3345 & w35564) | (w3345 & w35565) | (w35564 & w35565);
assign w31842 = (~w3345 & w35566) | (~w3345 & w35567) | (w35566 & w35567);
assign w31843 = w20602 & ~w20590;
assign w31844 = w20606 & ~w20579;
assign w31845 = w9528 & b_35;
assign w31846 = w20860 & w35568;
assign w31847 = w20856 & w20866;
assign w31848 = ~w20856 & ~w20866;
assign w31849 = w20869 & w20815;
assign w31850 = w6755 & b_44;
assign w31851 = a_47 & ~w27645;
assign w31852 = w26704 & a_47;
assign w31853 = ~w20902 & w20903;
assign w31854 = w20902 & ~w20903;
assign w31855 = w5956 & b_47;
assign w31856 = (a_44 & ~w20910) | (a_44 & w35569) | (~w20910 & w35569);
assign w31857 = a_44 & ~w27647;
assign w31858 = a_44 & ~w31856;
assign w31859 = w27647 & a_44;
assign w31860 = ~w20687 & ~w20689;
assign w31861 = ~w20687 & w20690;
assign w31862 = ~w20919 & w20920;
assign w31863 = w20919 & ~w20920;
assign w31864 = w5190 & b_50;
assign w31865 = w20927 & w35570;
assign w31866 = w4493 & b_53;
assign w31867 = w20944 & w35571;
assign w31868 = ~w20962 & ~w20961;
assign w31869 = (w27081 & w27082) | (w27081 & w31241) | (w27082 & w31241);
assign w31870 = (~w27438 & w35572) | (~w27438 & w35573) | (w35572 & w35573);
assign w31871 = (~w31868 & w20758) | (~w31868 & w35574) | (w20758 & w35574);
assign w31872 = w20960 & ~w20782;
assign w31873 = w2633 & b_63;
assign w31874 = ~w29820 & w35575;
assign w31875 = (~w29747 & w35576) | (~w29747 & w35577) | (w35576 & w35577);
assign w31876 = w20976 & a_29;
assign w31877 = ~w20976 & a_29;
assign w31878 = w3189 & b_60;
assign w31879 = w20989 & w35578;
assign w31880 = (w20793 & w20794) | (w20793 & w35579) | (w20794 & w35579);
assign w31881 = (w20950 & w20937) | (w20950 & w35580) | (w20937 & w35580);
assign w31882 = w4493 & b_54;
assign w31883 = w21005 & w35581;
assign w31884 = w20933 & ~w20922;
assign w31885 = w5190 & b_51;
assign w31886 = w21016 & w35582;
assign w31887 = w20916 & ~w20905;
assign w31888 = (w20804 & ~w20877) | (w20804 & w35583) | (~w20877 & w35583);
assign w31889 = w7607 & b_42;
assign w31890 = (a_50 & ~w21028) | (a_50 & w35584) | (~w21028 & w35584);
assign w31891 = a_50 & ~w26410;
assign w31892 = a_50 & ~w31890;
assign w31893 = w26410 & a_50;
assign w31894 = w20815 & ~w20870;
assign w31895 = (w20826 & w20845) | (w20826 & w35585) | (w20845 & w35585);
assign w31896 = w10556 & b_33;
assign w31897 = w21040 & w35586;
assign w31898 = a_63 & b_28;
assign w31899 = ~w21051 & ~w21052;
assign w31900 = ~w20830 & w35588;
assign w31901 = ~w21052 & ~w31899;
assign w31902 = ~w21052 & ~w31900;
assign w31903 = ~w31900 & w31899;
assign w31904 = w11614 & b_30;
assign w31905 = w21060 & w35589;
assign w31906 = w21056 & w21066;
assign w31907 = ~w21056 & ~w21066;
assign w31908 = w9528 & b_36;
assign w31909 = w21079 & w35590;
assign w31910 = w20856 & ~w20866;
assign w31911 = w8520 & b_39;
assign w31912 = w21098 & w35591;
assign w31913 = w21093 & w21104;
assign w31914 = ~w21093 & ~w21104;
assign w31915 = w6755 & b_45;
assign w31916 = ~w21127 & ~w21128;
assign w31917 = w5956 & b_48;
assign w31918 = (a_44 & ~w21136) | (a_44 & w35592) | (~w21136 & w35592);
assign w31919 = a_44 & ~w26413;
assign w31920 = a_44 & ~w31918;
assign w31921 = w26413 & a_44;
assign w31922 = w21129 & w35593;
assign w31923 = (~w21142 & ~w21129) | (~w21142 & w35594) | (~w21129 & w35594);
assign w31924 = w35595 & w35596;
assign w31925 = w35597 | w35598;
assign w31926 = w3797 & b_57;
assign w31927 = w21163 & w35599;
assign w31928 = w20985 & w21176;
assign w31929 = ~w20985 & ~w21176;
assign w31930 = (~w27757 & w35600) | (~w27757 & w35601) | (w35600 & w35601);
assign w31931 = (~w27438 & w35602) | (~w27438 & w35603) | (w35602 & w35603);
assign w31932 = (~w27757 & w35604) | (~w27757 & w35605) | (w35604 & w35605);
assign w31933 = (~w27438 & w35606) | (~w27438 & w35607) | (w35606 & w35607);
assign w31934 = w4493 & b_55;
assign w31935 = w21191 & w35608;
assign w31936 = w21034 & ~w21108;
assign w31937 = w21093 & ~w21104;
assign w31938 = w9528 & b_37;
assign w31939 = (a_56 & ~w21206) | (a_56 & w35609) | (~w21206 & w35609);
assign w31940 = a_56 & ~w26706;
assign w31941 = a_56 & ~w31939;
assign w31942 = w26706 & a_56;
assign w31943 = w21056 & ~w21066;
assign w31944 = a_63 & b_29;
assign w31945 = (~w31901 & w21223) | (~w31901 & w35610) | (w21223 & w35610);
assign w31946 = ~w21224 & ~w31902;
assign w31947 = ~w21224 & ~w31945;
assign w31948 = ~w21224 & ~w31946;
assign w31949 = w11614 & b_31;
assign w31950 = w21232 & w35611;
assign w31951 = w10556 & b_34;
assign w31952 = w21245 & w35612;
assign w31953 = w21085 & ~w21073;
assign w31954 = ~w21260 & w21261;
assign w31955 = w21260 & ~w21261;
assign w31956 = w8520 & b_40;
assign w31957 = a_53 & ~w26707;
assign w31958 = w26415 & a_53;
assign w31959 = w7607 & b_43;
assign w31960 = a_50 & ~w26416;
assign w31961 = w26012 & a_50;
assign w31962 = w6755 & b_46;
assign w31963 = ~w21114 & w21126;
assign w31964 = w5956 & b_49;
assign w31965 = a_44 & ~w26422;
assign w31966 = w26015 & a_44;
assign w31967 = w21326 & ~w21325;
assign w31968 = w21326 & w27649;
assign w31969 = w5190 & b_52;
assign w31970 = w21334 & w35613;
assign w31971 = ~w21330 & w21340;
assign w31972 = w21330 & ~w21340;
assign w31973 = w21011 & ~w21151;
assign w31974 = ~w21349 & w21350;
assign w31975 = w21349 & ~w21350;
assign w31976 = w3797 & b_58;
assign w31977 = w21357 & w35614;
assign w31978 = (w21169 & w21001) | (w21169 & w35615) | (w21001 & w35615);
assign w31979 = ~w21366 & w21367;
assign w31980 = w21366 & ~w21367;
assign w31981 = w21173 & ~w20998;
assign w31982 = w3189 & b_61;
assign w31983 = w21375 & w35616;
assign w31984 = (~w21371 & w35617) | (~w21371 & ~w21370) | (w35617 & ~w21370);
assign w31985 = w35618 & w21371;
assign w31986 = w3189 & b_62;
assign w31987 = (w9770 & w35619) | (w9770 & w35620) | (w35619 & w35620);
assign w31988 = w21395 & w35621;
assign w31989 = (~a_32 & ~w21395) | (~a_32 & w35622) | (~w21395 & w35622);
assign w31990 = w21364 & ~w21399;
assign w31991 = (w21399 & ~w21353) | (w21399 & w35623) | (~w21353 & w35623);
assign w31992 = w4493 & b_56;
assign w31993 = w21406 & w35624;
assign w31994 = w8520 & b_41;
assign w31995 = a_53 & ~w26709;
assign w31996 = w26424 & a_53;
assign w31997 = w9528 & b_38;
assign w31998 = (a_56 & ~w21428) | (a_56 & w35625) | (~w21428 & w35625);
assign w31999 = a_56 & ~w26711;
assign w32000 = a_56 & ~w31998;
assign w32001 = w26711 & a_56;
assign w32002 = w21214 & ~w21252;
assign w32003 = w10556 & b_35;
assign w32004 = w21439 & w35626;
assign w32005 = w21238 & ~w21225;
assign w32006 = w21050 & ~w21218;
assign w32007 = w11614 & b_32;
assign w32008 = (a_62 & ~w21457) | (a_62 & w35627) | (~w21457 & w35627);
assign w32009 = a_62 & ~w26425;
assign w32010 = a_62 & ~w32008;
assign w32011 = w26425 & a_62;
assign w32012 = (w3967 & w35628) | (w3967 & w35629) | (w35628 & w35629);
assign w32013 = (~w3967 & w35630) | (~w3967 & w35631) | (w35630 & w35631);
assign w32014 = w35632 & w21446;
assign w32015 = ~w21471 & w21434;
assign w32016 = w7607 & b_44;
assign w32017 = w21200 & ~w21292;
assign w32018 = w6755 & b_47;
assign w32019 = a_47 & ~w26428;
assign w32020 = w26017 & a_47;
assign w32021 = ~w21308 & w21311;
assign w32022 = ~w21308 & ~w21310;
assign w32023 = ~w21520 & w21521;
assign w32024 = w21520 & ~w21521;
assign w32025 = w5956 & b_50;
assign w32026 = (a_44 & ~w21528) | (a_44 & w35633) | (~w21528 & w35633);
assign w32027 = a_44 & ~w26430;
assign w32028 = a_44 & ~w32026;
assign w32029 = w26430 & a_44;
assign w32030 = w5190 & b_53;
assign w32031 = w21543 & w35634;
assign w32032 = w21538 & w35635;
assign w32033 = (w21549 & ~w21538) | (w21549 & w35636) | (~w21538 & w35636);
assign w32034 = w3797 & b_59;
assign w32035 = w21567 & w35637;
assign w32036 = ~w21575 & ~w21574;
assign w32037 = w21382 & ~w21579;
assign w32038 = (~w27757 & w35638) | (~w27757 & w35639) | (w35638 & w35639);
assign w32039 = (~w27438 & w35640) | (~w27438 & w35641) | (w35640 & w35641);
assign w32040 = w3189 & b_63;
assign w32041 = ~w3198 & ~w21590;
assign w32042 = w5190 & b_54;
assign w32043 = (a_41 & ~w21603) | (a_41 & w35642) | (~w21603 & w35642);
assign w32044 = a_41 & ~w26431;
assign w32045 = a_41 & ~w32043;
assign w32046 = w26431 & a_41;
assign w32047 = w5956 & b_51;
assign w32048 = (a_44 & ~w21614) | (a_44 & w35643) | (~w21614 & w35643);
assign w32049 = a_44 & ~w26432;
assign w32050 = a_44 & ~w32048;
assign w32051 = w26432 & a_44;
assign w32052 = w21423 & ~w21480;
assign w32053 = w8520 & b_42;
assign w32054 = w21434 & ~w21472;
assign w32055 = w9528 & b_39;
assign w32056 = (a_56 & ~w21637) | (a_56 & w35644) | (~w21637 & w35644);
assign w32057 = a_56 & ~w27655;
assign w32058 = a_56 & ~w32056;
assign w32059 = w27655 & a_56;
assign w32060 = a_63 & b_31;
assign w32061 = ~w21450 & w35645;
assign w32062 = ~w21649 & ~w21650;
assign w32063 = ~w21649 & w32061;
assign w32064 = ~w21649 & ~w32062;
assign w32065 = ~w32061 & ~w21649;
assign w32066 = w32062 & ~w32061;
assign w32067 = w11614 & b_33;
assign w32068 = w21659 & w35646;
assign w32069 = w21654 & ~w21665;
assign w32070 = w10556 & b_36;
assign w32071 = w21673 & w35647;
assign w32072 = w7607 & b_45;
assign w32073 = ~w21707 & ~w21706;
assign w32074 = ~w21707 & ~w21697;
assign w32075 = ~w21489 & w21500;
assign w32076 = ~w21708 & ~w21709;
assign w32077 = w6755 & b_48;
assign w32078 = w21711 & w21723;
assign w32079 = ~w21711 & ~w21723;
assign w32080 = w21599 & w21738;
assign w32081 = ~w21599 & ~w21738;
assign w32082 = w4493 & b_57;
assign w32083 = w21745 & w35648;
assign w32084 = (w21412 & w21413) | (w21412 & w35649) | (w21413 & w35649);
assign w32085 = w3797 & b_60;
assign w32086 = w21763 & w35650;
assign w32087 = w21598 & w21773;
assign w32088 = ~w21598 & ~w21773;
assign w32089 = (~w27757 & w35651) | (~w27757 & w35652) | (w35651 & w35652);
assign w32090 = (~w27438 & w35653) | (~w27438 & w35654) | (w35653 & w35654);
assign w32091 = (~w27757 & w35655) | (~w27757 & w35656) | (w35655 & w35656);
assign w32092 = (~w27438 & w35657) | (~w27438 & w35658) | (w35657 & w35658);
assign w32093 = w21598 & ~w21773;
assign w32094 = w5190 & b_55;
assign w32095 = w21788 & w35659;
assign w32096 = w9528 & b_40;
assign w32097 = w21679 & ~w21666;
assign w32098 = ~w12380 & w35660;
assign w32099 = (a_32 & w12380) | (a_32 & w35661) | (w12380 & w35661);
assign w32100 = ~w21815 & ~w32064;
assign w32101 = ~w21815 & ~w32065;
assign w32102 = ~w21815 & ~w32100;
assign w32103 = ~w21815 & ~w32101;
assign w32104 = w11614 & b_34;
assign w32105 = w21822 & w35662;
assign w32106 = w21818 & w21828;
assign w32107 = ~w21818 & ~w21828;
assign w32108 = w10556 & b_37;
assign w32109 = (a_59 & ~w21835) | (a_59 & w35663) | (~w21835 & w35663);
assign w32110 = a_59 & ~w26441;
assign w32111 = a_59 & ~w32109;
assign w32112 = w26441 & a_59;
assign w32113 = w21643 & ~w21683;
assign w32114 = w8520 & b_43;
assign w32115 = w21632 & ~w21689;
assign w32116 = ~w21867 & ~w21868;
assign w32117 = w7607 & b_46;
assign w32118 = ~w21870 & ~w21881;
assign w32119 = ~w21870 & w21881;
assign w32120 = ~w21695 & ~w21706;
assign w32121 = ~w21695 & ~w21697;
assign w32122 = w6755 & b_49;
assign w32123 = ~w21899 & w21888;
assign w32124 = ~w21899 & ~w21796;
assign w32125 = ~w21899 & ~w21888;
assign w32126 = ~w21899 & w21796;
assign w32127 = w5956 & b_52;
assign w32128 = (a_44 & ~w21908) | (a_44 & w35664) | (~w21908 & w35664);
assign w32129 = a_44 & ~w26444;
assign w32130 = a_44 & ~w32128;
assign w32131 = w26444 & a_44;
assign w32132 = w21609 & ~w21733;
assign w32133 = w4493 & b_58;
assign w32134 = w21930 & w35665;
assign w32135 = (~w32080 & w35666) | (~w32080 & w35667) | (w35666 & w35667);
assign w32136 = ~w21939 & w21940;
assign w32137 = w21939 & ~w21940;
assign w32138 = w3797 & b_61;
assign w32139 = w21948 & w35668;
assign w32140 = (~w21944 & w35669) | (~w21944 & ~w21943) | (w35669 & ~w21943);
assign w32141 = w35670 & w21944;
assign w32142 = w21596 & w21959;
assign w32143 = ~w21596 & ~w21959;
assign w32144 = w3797 & b_62;
assign w32145 = (w9770 & w35671) | (w9770 & w35672) | (w35671 & w35672);
assign w32146 = w21968 & w35673;
assign w32147 = (~a_35 & ~w21968) | (~a_35 & w35674) | (~w21968 & w35674);
assign w32148 = w21937 & ~w21972;
assign w32149 = (w21972 & ~w21926) | (w21972 & w35675) | (~w21926 & w35675);
assign w32150 = w5190 & b_56;
assign w32151 = w21979 & w35676;
assign w32152 = w21795 & ~w21916;
assign w32153 = w9528 & b_41;
assign w32154 = (a_56 & ~w21990) | (a_56 & w35677) | (~w21990 & w35677);
assign w32155 = a_56 & ~w27663;
assign w32156 = a_56 & ~w32154;
assign w32157 = w27663 & a_56;
assign w32158 = w10556 & b_38;
assign w32159 = w22001 & w35678;
assign w32160 = w21818 & ~w21828;
assign w32161 = a_63 & b_33;
assign w32162 = w21648 & ~w21809;
assign w32163 = w11614 & b_35;
assign w32164 = a_62 & ~w26033;
assign w32165 = w25688 & a_62;
assign w32166 = (w4636 & w35679) | (w4636 & w35680) | (w35679 & w35680);
assign w32167 = (~w4636 & w35681) | (~w4636 & w35682) | (w35681 & w35682);
assign w32168 = w21816 & w22027;
assign w32169 = ~w32168 & w22027;
assign w32170 = w22030 & ~w22007;
assign w32171 = w8520 & b_44;
assign w32172 = a_53 & ~w27664;
assign w32173 = w26716 & a_53;
assign w32174 = ~w21866 & ~w21868;
assign w32175 = ~w21866 & w21869;
assign w32176 = ~w22058 & w22059;
assign w32177 = w22058 & ~w22059;
assign w32178 = w7607 & b_47;
assign w32179 = (a_50 & ~w22066) | (a_50 & w35683) | (~w22066 & w35683);
assign w32180 = a_50 & ~w27666;
assign w32181 = a_50 & ~w32179;
assign w32182 = w27666 & a_50;
assign w32183 = ~w21882 & ~w21884;
assign w32184 = ~w21882 & w21885;
assign w32185 = w6755 & b_50;
assign w32186 = w22084 & w35684;
assign w32187 = w5956 & b_53;
assign w32188 = w22101 & w35685;
assign w32189 = w4493 & b_59;
assign w32190 = w22125 & w35686;
assign w32191 = ~w22133 & ~w22132;
assign w32192 = ~w32191 & ~w22133;
assign w32193 = (~w27757 & w35687) | (~w27757 & w35688) | (w35687 & w35688);
assign w32194 = (~w27438 & w35689) | (~w27438 & w35690) | (w35689 & w35690);
assign w32195 = (~w27757 & w35691) | (~w27757 & w35692) | (w35691 & w35692);
assign w32196 = (~w27438 & w35693) | (~w27438 & w35694) | (w35693 & w35694);
assign w32197 = ~w32191 & ~w21973;
assign w32198 = w22131 & ~w22120;
assign w32199 = w3797 & b_63;
assign w32200 = ~w3806 & ~w22149;
assign w32201 = (w22107 & w22094) | (w22107 & w35695) | (w22094 & w35695);
assign w32202 = w5956 & b_54;
assign w32203 = w22163 & w35696;
assign w32204 = (w22090 & w22076) | (w22090 & w35697) | (w22076 & w35697);
assign w32205 = w6755 & b_51;
assign w32206 = w22174 & w35698;
assign w32207 = w22072 & ~w22061;
assign w32208 = (w21996 & w21997) | (w21996 & w35699) | (w21997 & w35699);
assign w32209 = w9528 & b_42;
assign w32210 = (a_56 & ~w22186) | (a_56 & w35700) | (~w22186 & w35700);
assign w32211 = a_56 & ~w27667;
assign w32212 = a_56 & ~w32210;
assign w32213 = w27667 & a_56;
assign w32214 = a_63 & b_34;
assign w32215 = ~w22198 & ~w22199;
assign w32216 = ~w22013 & w35702;
assign w32217 = ~w22198 & ~w32215;
assign w32218 = ~w22198 & ~w32216;
assign w32219 = ~w32216 & w32215;
assign w32220 = w11614 & b_36;
assign w32221 = w22207 & w35703;
assign w32222 = w22202 & ~w22213;
assign w32223 = w10556 & b_39;
assign w32224 = w22221 & w35704;
assign w32225 = w8520 & b_45;
assign w32226 = (w22055 & w22041) | (w22055 & w35705) | (w22041 & w35705);
assign w32227 = ~w22250 & ~w22251;
assign w32228 = w7607 & b_48;
assign w32229 = w22257 & w35706;
assign w32230 = w22252 & w35707;
assign w32231 = (~w22263 & ~w22252) | (~w22263 & w35708) | (~w22252 & w35708);
assign w32232 = ~w22266 & w22180;
assign w32233 = w5190 & b_57;
assign w32234 = w22287 & w35709;
assign w32235 = w21985 & ~w22111;
assign w32236 = w4493 & b_60;
assign w32237 = w22305 & w35710;
assign w32238 = w22157 & w22315;
assign w32239 = ~w22157 & ~w22315;
assign w32240 = (~w27757 & w35711) | (~w27757 & w35712) | (w35711 & w35712);
assign w32241 = (~w27438 & w35713) | (~w27438 & w35714) | (w35713 & w35714);
assign w32242 = w22180 & ~w22267;
assign w32243 = w6755 & b_52;
assign w32244 = w22329 & w35715;
assign w32245 = a_63 & b_35;
assign w32246 = w22345 & ~w32217;
assign w32247 = w22345 & ~w32218;
assign w32248 = ~w22345 & w32217;
assign w32249 = ~w22345 & w32218;
assign w32250 = w11614 & b_37;
assign w32251 = w22352 & w35716;
assign w32252 = w10556 & b_40;
assign w32253 = w22227 & ~w22214;
assign w32254 = w9528 & b_43;
assign w32255 = w22379 & ~w22390;
assign w32256 = w22192 & ~w22231;
assign w32257 = w8520 & b_46;
assign w32258 = w22249 & ~w22237;
assign w32259 = w22411 & ~w22413;
assign w32260 = w7607 & b_49;
assign w32261 = a_50 & ~w26447;
assign w32262 = w26042 & a_50;
assign w32263 = w22415 & w22425;
assign w32264 = ~w22415 & ~w22425;
assign w32265 = w5956 & b_55;
assign w32266 = w22441 & w35717;
assign w32267 = w22169 & ~w22275;
assign w32268 = w5190 & b_58;
assign w32269 = w22458 & w35718;
assign w32270 = (w22293 & w22159) | (w22293 & w35719) | (w22159 & w35719);
assign w32271 = w4493 & b_61;
assign w32272 = w22476 & w35720;
assign w32273 = (w22311 & w22297) | (w22311 & w35721) | (w22297 & w35721);
assign w32274 = w22157 & ~w22315;
assign w32275 = w22155 & w22490;
assign w32276 = ~w22155 & ~w22490;
assign w32277 = w22469 & ~w22465;
assign w32278 = w4493 & b_62;
assign w32279 = (w9770 & w35722) | (w9770 & w35723) | (w35722 & w35723);
assign w32280 = w22501 & w35724;
assign w32281 = (~a_38 & ~w22501) | (~a_38 & w35725) | (~w22501 & w35725);
assign w32282 = w11614 & b_38;
assign w32283 = a_62 & ~w26043;
assign w32284 = w25695 & a_62;
assign w32285 = a_63 & b_36;
assign w32286 = w22339 & ~w22522;
assign w32287 = (~w5363 & w35726) | (~w5363 & w35727) | (w35726 & w35727);
assign w32288 = w10556 & b_41;
assign w32289 = a_59 & ~w26045;
assign w32290 = w25696 & a_59;
assign w32291 = w9528 & b_44;
assign w32292 = w8520 & b_47;
assign w32293 = w7607 & b_50;
assign w32294 = a_50 & ~w26053;
assign w32295 = w25701 & a_50;
assign w32296 = ~w22427 & ~w22428;
assign w32297 = w6755 & b_53;
assign w32298 = (a_47 & ~w22611) | (a_47 & w35728) | (~w22611 & w35728);
assign w32299 = a_47 & ~w26450;
assign w32300 = a_47 & ~w32298;
assign w32301 = w26450 & a_47;
assign w32302 = w5956 & b_56;
assign w32303 = w22629 & w35729;
assign w32304 = ~w22448 & w22451;
assign w32305 = ~w22448 & ~w22449;
assign w32306 = w5190 & b_59;
assign w32307 = w22646 & w35730;
assign w32308 = ~w22654 & ~w22653;
assign w32309 = w22487 & ~w22483;
assign w32310 = (~w27757 & w35731) | (~w27757 & w35732) | (w35731 & w35732);
assign w32311 = (~w27438 & w35733) | (~w27438 & w35734) | (w35733 & w35734);
assign w32312 = (~w27757 & w35735) | (~w27757 & w35736) | (w35735 & w35736);
assign w32313 = (~w27438 & w35737) | (~w27438 & w35738) | (w35737 & w35738);
assign w32314 = ~w32308 & ~w22506;
assign w32315 = w4493 & b_63;
assign w32316 = ~w4502 & ~w22668;
assign w32317 = w6755 & b_54;
assign w32318 = w22682 & w35739;
assign w32319 = (w22598 & w22584) | (w22598 & w35740) | (w22584 & w35740);
assign w32320 = w7607 & b_51;
assign w32321 = w22693 & w35741;
assign w32322 = (w22580 & w22566) | (w22580 & w35742) | (w22566 & w35742);
assign w32323 = a_63 & b_37;
assign w32324 = w22524 & ~w22708;
assign w32325 = ~w22524 & ~w22708;
assign w32326 = w11614 & b_39;
assign w32327 = w22716 & w35743;
assign w32328 = w22711 & ~w22722;
assign w32329 = w10556 & b_42;
assign w32330 = a_59 & ~w27675;
assign w32331 = w26453 & a_59;
assign w32332 = (w22545 & w22532) | (w22545 & w35744) | (w22532 & w35744);
assign w32333 = w9528 & b_45;
assign w32334 = ~w22753 & ~w22752;
assign w32335 = ~w22753 & ~w22743;
assign w32336 = (w22563 & w22549) | (w22563 & w35745) | (w22549 & w35745);
assign w32337 = w8520 & b_48;
assign w32338 = (a_53 & ~w22763) | (a_53 & w35746) | (~w22763 & w35746);
assign w32339 = a_53 & ~w26458;
assign w32340 = a_53 & ~w32338;
assign w32341 = w26458 & a_53;
assign w32342 = w22774 & ~w22699;
assign w32343 = w22699 & ~w22774;
assign w32344 = w5956 & b_57;
assign w32345 = w22791 & w35747;
assign w32346 = (w22635 & w22621) | (w22635 & w35748) | (w22621 & w35748);
assign w32347 = w5190 & b_60;
assign w32348 = w22809 & w35749;
assign w32349 = (~w27757 & w35750) | (~w27757 & w35751) | (w35750 & w35751);
assign w32350 = (~w27438 & w35752) | (~w27438 & w35753) | (w35752 & w35753);
assign w32351 = w7607 & b_52;
assign w32352 = a_50 & ~w26459;
assign w32353 = w26058 & a_50;
assign w32354 = (~w26457 & w35754) | (~w26457 & w35755) | (w35754 & w35755);
assign w32355 = ~w22705 & w22708;
assign w32356 = (~w22705 & ~w22524) | (~w22705 & w32355) | (~w22524 & w32355);
assign w32357 = a_63 & b_38;
assign w32358 = w22849 & ~w32355;
assign w32359 = w22849 & ~w32356;
assign w32360 = ~w22849 & w32355;
assign w32361 = ~w22849 & w32356;
assign w32362 = w11614 & b_40;
assign w32363 = w22856 & w35756;
assign w32364 = w10556 & b_43;
assign w32365 = w22865 & ~w22875;
assign w32366 = w22865 & w22875;
assign w32367 = w22736 & ~w22723;
assign w32368 = w9528 & b_46;
assign w32369 = w27678 & w35757;
assign w32370 = (~w22894 & ~w27678) | (~w22894 & w35758) | (~w27678 & w35758);
assign w32371 = (~w22752 & w22739) | (~w22752 & w35759) | (w22739 & w35759);
assign w32372 = ~w22742 & ~w22743;
assign w32373 = w8520 & b_49;
assign w32374 = a_53 & ~w26464;
assign w32375 = w26065 & a_53;
assign w32376 = w6755 & b_55;
assign w32377 = (a_47 & ~w22927) | (a_47 & w35760) | (~w22927 & w35760);
assign w32378 = a_47 & ~w26466;
assign w32379 = a_47 & ~w32377;
assign w32380 = w26466 & a_47;
assign w32381 = w22688 & ~w22779;
assign w32382 = w5956 & b_58;
assign w32383 = w22944 & w35761;
assign w32384 = (w22797 & w22678) | (w22797 & w35762) | (w22678 & w35762);
assign w32385 = w5190 & b_61;
assign w32386 = w22962 & w35763;
assign w32387 = (w22815 & w22801) | (w22815 & w35764) | (w22801 & w35764);
assign w32388 = w22819 & ~w22674;
assign w32389 = ~w22951 & w22955;
assign w32390 = ~w22951 & ~w22952;
assign w32391 = w5190 & b_62;
assign w32392 = (w9770 & w35765) | (w9770 & w35766) | (w35765 & w35766);
assign w32393 = w22987 & w35767;
assign w32394 = (~a_41 & ~w22987) | (~a_41 & w35768) | (~w22987 & w35768);
assign w32395 = w22862 & ~w22850;
assign w32396 = a_63 & b_39;
assign w32397 = w22843 & ~w22999;
assign w32398 = w11614 & b_41;
assign w32399 = ~w23004 & ~w11623;
assign w32400 = ~w23008 & ~w23009;
assign w32401 = ~a_62 & ~w23009;
assign w32402 = ~a_62 & w32400;
assign w32403 = (w5888 & w35769) | (w5888 & w35770) | (w35769 & w35770);
assign w32404 = (~w5888 & w35771) | (~w5888 & w35772) | (w35771 & w35772);
assign w32405 = w10556 & b_44;
assign w32406 = ~w22876 & w22880;
assign w32407 = ~w22876 & ~w22878;
assign w32408 = w9528 & b_47;
assign w32409 = w8520 & b_50;
assign w32410 = a_53 & ~w26474;
assign w32411 = w26070 & a_53;
assign w32412 = w7607 & b_53;
assign w32413 = w23075 & w35773;
assign w32414 = w6755 & b_56;
assign w32415 = w23093 & w35774;
assign w32416 = w5956 & b_59;
assign w32417 = w23110 & w35775;
assign w32418 = ~w23118 & ~w23117;
assign w32419 = ~w32418 & ~w23118;
assign w32420 = w22973 & ~w22969;
assign w32421 = ~w32418 & ~w22992;
assign w32422 = w23116 & ~w23105;
assign w32423 = w5190 & b_63;
assign w32424 = ~w5199 & ~w23133;
assign w32425 = w6755 & b_57;
assign w32426 = w23145 & w35776;
assign w32427 = w7607 & b_54;
assign w32428 = w23155 & w35777;
assign w32429 = w23062 & ~w23051;
assign w32430 = w8520 & b_51;
assign w32431 = w23166 & w35778;
assign w32432 = (w23044 & w23031) | (w23044 & w35779) | (w23031 & w35779);
assign w32433 = (w23027 & w22995) | (w23027 & w35780) | (w22995 & w35780);
assign w32434 = a_63 & b_40;
assign w32435 = w23001 & ~w23182;
assign w32436 = ~w23001 & ~w23182;
assign w32437 = w11614 & b_42;
assign w32438 = w23189 & w35781;
assign w32439 = w23185 & w23195;
assign w32440 = ~w23185 & ~w23195;
assign w32441 = w10556 & b_45;
assign w32442 = a_59 & ~w27684;
assign w32443 = w26722 & a_59;
assign w32444 = w9528 & b_48;
assign w32445 = w23218 & w35782;
assign w32446 = w23230 & ~w23172;
assign w32447 = w23237 & ~w23161;
assign w32448 = w23068 & w23241;
assign w32449 = ~w23068 & ~w23241;
assign w32450 = (w23099 & w23085) | (w23099 & w35783) | (w23085 & w35783);
assign w32451 = w5956 & b_60;
assign w32452 = w23256 & w35784;
assign w32453 = w23141 & w23266;
assign w32454 = ~w23141 & ~w23266;
assign w32455 = w6755 & b_58;
assign w32456 = w23279 & w35785;
assign w32457 = w7607 & b_55;
assign w32458 = w23290 & w35786;
assign w32459 = w23224 & ~w23213;
assign w32460 = w9528 & b_49;
assign w32461 = (a_56 & ~w23302) | (a_56 & w35787) | (~w23302 & w35787);
assign w32462 = a_56 & ~w27686;
assign w32463 = a_56 & ~w32461;
assign w32464 = w27686 & a_56;
assign w32465 = a_63 & b_41;
assign w32466 = w11614 & b_43;
assign w32467 = ~w23179 & w23182;
assign w32468 = (~w23179 & ~w23001) | (~w23179 & w32467) | (~w23001 & w32467);
assign w32469 = w10556 & b_46;
assign w32470 = w23185 & ~w23195;
assign w32471 = w23355 & ~w23298;
assign w32472 = w8520 & b_52;
assign w32473 = w23365 & w35788;
assign w32474 = w23151 & ~w23242;
assign w32475 = w5956 & b_61;
assign w32476 = w23395 & w35789;
assign w32477 = w23262 & ~w23251;
assign w32478 = w23141 & ~w23266;
assign w32479 = w23139 & w23409;
assign w32480 = ~w23139 & ~w23409;
assign w32481 = w23388 & ~w23384;
assign w32482 = w5956 & b_62;
assign w32483 = (w9770 & w35790) | (w9770 & w35791) | (w35790 & w35791);
assign w32484 = w23420 & w35792;
assign w32485 = (~a_44 & ~w23420) | (~a_44 & w35793) | (~w23420 & w35793);
assign w32486 = w6755 & b_59;
assign w32487 = w23431 & w35794;
assign w32488 = w23297 & ~w23373;
assign w32489 = w23332 & ~w23328;
assign w32490 = a_63 & b_42;
assign w32491 = w23314 & ~w23443;
assign w32492 = w11614 & b_44;
assign w32493 = ~w23449 & ~w11623;
assign w32494 = ~w23453 & ~w23454;
assign w32495 = ~a_62 & ~w23454;
assign w32496 = ~a_62 & w32494;
assign w32497 = (w6974 & w35795) | (w6974 & w35796) | (w35795 & w35796);
assign w32498 = (~w6974 & w35797) | (~w6974 & w35798) | (w35797 & w35798);
assign w32499 = w23459 & w23328;
assign w32500 = w23459 & ~w32489;
assign w32501 = ~w23459 & ~w23328;
assign w32502 = ~w23459 & w32489;
assign w32503 = w10556 & b_47;
assign w32504 = (a_59 & ~w23466) | (a_59 & w35799) | (~w23466 & w35799);
assign w32505 = a_59 & ~w27694;
assign w32506 = a_59 & ~w32504;
assign w32507 = w27694 & a_59;
assign w32508 = ~w23346 & w23350;
assign w32509 = ~w23346 & ~w23348;
assign w32510 = w9528 & b_50;
assign w32511 = w23484 & w35800;
assign w32512 = w8520 & b_53;
assign w32513 = w23502 & w35801;
assign w32514 = w7607 & b_56;
assign w32515 = w23519 & w35802;
assign w32516 = w23406 & ~w23402;
assign w32517 = w23437 & ~w23529;
assign w32518 = w5956 & b_63;
assign w32519 = ~w5965 & ~w23550;
assign w32520 = ~w23555 & w23529;
assign w32521 = (~w23555 & w23529) | (~w23555 & w35803) | (w23529 & w35803);
assign w32522 = w7607 & b_57;
assign w32523 = w23563 & w35804;
assign w32524 = w23508 & ~w23497;
assign w32525 = w8520 & b_54;
assign w32526 = w23574 & w35805;
assign w32527 = w23490 & ~w23479;
assign w32528 = w9528 & b_51;
assign w32529 = w23585 & w35806;
assign w32530 = w23472 & ~w23460;
assign w32531 = w10556 & b_48;
assign w32532 = (a_59 & ~w23596) | (a_59 & w35807) | (~w23596 & w35807);
assign w32533 = a_59 & ~w27695;
assign w32534 = a_59 & ~w32532;
assign w32535 = w27695 & a_59;
assign w32536 = a_63 & b_43;
assign w32537 = w11614 & b_45;
assign w32538 = ~w23610 & ~w11623;
assign w32539 = ~w23621 & w23602;
assign w32540 = w23631 & ~w23591;
assign w32541 = w23591 & ~w23631;
assign w32542 = ~w23635 & w23580;
assign w32543 = (w23525 & w23512) | (w23525 & w35808) | (w23512 & w35808);
assign w32544 = w6755 & b_60;
assign w32545 = w23660 & w35809;
assign w32546 = w6755 & b_61;
assign w32547 = w23683 & w35810;
assign w32548 = w23569 & ~w23644;
assign w32549 = w7607 & b_58;
assign w32550 = w23694 & w35811;
assign w32551 = w23580 & ~w23636;
assign w32552 = w8520 & b_55;
assign w32553 = w23705 & w35812;
assign w32554 = w9528 & b_52;
assign w32555 = w23716 & w35813;
assign w32556 = w23602 & ~w23622;
assign w32557 = a_63 & b_44;
assign w32558 = ~w23734 & ~w27697;
assign w32559 = ~w23734 & ~w27696;
assign w32560 = w11614 & b_46;
assign w32561 = (a_62 & ~w23742) | (a_62 & w35814) | (~w23742 & w35814);
assign w32562 = a_62 & ~w27698;
assign w32563 = a_62 & ~w32561;
assign w32564 = w27698 & a_62;
assign w32565 = w23737 & ~w23748;
assign w32566 = w10556 & b_49;
assign w32567 = (a_59 & ~w23756) | (a_59 & w35815) | (~w23756 & w35815);
assign w32568 = a_59 & ~w27699;
assign w32569 = a_59 & ~w32567;
assign w32570 = w27699 & a_59;
assign w32571 = w23666 & ~w23653;
assign w32572 = w23670 & ~w23556;
assign w32573 = w6755 & b_62;
assign w32574 = (w9770 & w35816) | (w9770 & w35817) | (w35816 & w35817);
assign w32575 = w23804 & w35818;
assign w32576 = (~a_47 & ~w23804) | (~a_47 & w35819) | (~w23804 & w35819);
assign w32577 = w23782 & ~w23808;
assign w32578 = (w23808 & ~w23780) | (w23808 & w35820) | (~w23780 & w35820);
assign w32579 = w7607 & b_59;
assign w32580 = w23815 & w35821;
assign w32581 = w9528 & b_53;
assign w32582 = w23827 & w35822;
assign w32583 = w23723 & ~w23764;
assign w32584 = w10556 & b_50;
assign w32585 = (a_59 & ~w23838) | (a_59 & w35823) | (~w23838 & w35823);
assign w32586 = a_59 & ~w26483;
assign w32587 = a_59 & ~w32585;
assign w32588 = w26483 & a_59;
assign w32589 = a_63 & b_45;
assign w32590 = w23442 & ~w23728;
assign w32591 = w11614 & b_47;
assign w32592 = (w7859 & w35824) | (w7859 & w35825) | (w35824 & w35825);
assign w32593 = w23735 & w23863;
assign w32594 = ~w23863 & w23844;
assign w32595 = w8520 & b_56;
assign w32596 = w23885 & w35826;
assign w32597 = ~w23788 & w35827;
assign w32598 = (w27757 & w35828) | (w27757 & w35829) | (w35828 & w35829);
assign w32599 = (w27438 & w35830) | (w27438 & w35831) | (w35830 & w35831);
assign w32600 = w8520 & b_57;
assign w32601 = w23917 & w35832;
assign w32602 = w23833 & ~w23872;
assign w32603 = w9528 & b_54;
assign w32604 = (a_56 & ~w23928) | (a_56 & w35833) | (~w23928 & w35833);
assign w32605 = a_56 & ~w26486;
assign w32606 = a_56 & ~w32604;
assign w32607 = w26486 & a_56;
assign w32608 = w23844 & ~w23864;
assign w32609 = w10556 & b_51;
assign w32610 = w23939 & w35834;
assign w32611 = a_63 & b_46;
assign w32612 = ~w26488 & w26487;
assign w32613 = w11614 & b_48;
assign w32614 = w23959 & w35835;
assign w32615 = w23955 & w23965;
assign w32616 = ~w23955 & ~w23965;
assign w32617 = ~w23971 & w23934;
assign w32618 = w23891 & ~w23987;
assign w32619 = w7607 & b_60;
assign w32620 = w23996 & w35836;
assign w32621 = w23991 & ~w24002;
assign w32622 = w6755 & b_63;
assign w32623 = (~w24007 & w29820) | (~w24007 & w35837) | (w29820 & w35837);
assign w32624 = (w29747 & w35838) | (w29747 & w35839) | (w35838 & w35839);
assign w32625 = ~w24007 & w35818;
assign w32626 = (~a_47 & w24007) | (~a_47 & w35819) | (w24007 & w35819);
assign w32627 = ~w24011 & w23895;
assign w32628 = (~w24011 & w23895) | (~w24011 & w35840) | (w23895 & w35840);
assign w32629 = w24011 & ~w23895;
assign w32630 = ~w23895 & w35841;
assign w32631 = ~w23811 & ~w23809;
assign w32632 = w7607 & b_61;
assign w32633 = w24029 & w35842;
assign w32634 = (w23923 & ~w23979) | (w23923 & w35843) | (~w23979 & w35843);
assign w32635 = w8520 & b_58;
assign w32636 = w24040 & w35844;
assign w32637 = w23934 & ~w23972;
assign w32638 = w9528 & b_55;
assign w32639 = w24051 & w35845;
assign w32640 = w23955 & ~w23965;
assign w32641 = w11614 & b_49;
assign w32642 = a_62 & ~w27702;
assign w32643 = w24064 & w35846;
assign w32644 = a_63 & b_47;
assign w32645 = (~w8186 & w35847) | (~w8186 & w35848) | (w35847 & w35848);
assign w32646 = w10556 & b_52;
assign w32647 = w24089 & w35849;
assign w32648 = ~w24084 & w24095;
assign w32649 = w24084 & ~w24095;
assign w32650 = w7607 & b_62;
assign w32651 = (~w9770 & w35850) | (~w9770 & w35851) | (w35850 & w35851);
assign w32652 = ~w24131 & a_50;
assign w32653 = w24131 & a_50;
assign w32654 = w8520 & b_59;
assign w32655 = w24142 & w35852;
assign w32656 = w9528 & b_56;
assign w32657 = w24153 & w35853;
assign w32658 = w10556 & b_53;
assign w32659 = w24164 & w35854;
assign w32660 = w23954 & ~w24079;
assign w32661 = a_63 & b_48;
assign w32662 = w24072 & ~w24175;
assign w32663 = w11614 & b_50;
assign w32664 = ~w24180 & ~w11623;
assign w32665 = ~w24184 & ~w24185;
assign w32666 = ~a_62 & ~w24185;
assign w32667 = ~a_62 & w32665;
assign w32668 = (w8793 & w35855) | (w8793 & w35856) | (w35855 & w35856);
assign w32669 = (~w8793 & w35857) | (~w8793 & w35858) | (w35857 & w35858);
assign w32670 = w35859 & w24171;
assign w32671 = ~w24203 & w24148;
assign w32672 = ~w24115 & w35860;
assign w32673 = w9528 & b_57;
assign w32674 = w24229 & w35861;
assign w32675 = w11614 & b_51;
assign w32676 = a_63 & b_49;
assign w32677 = w10556 & b_54;
assign w32678 = w24265 & w35862;
assign w32679 = (w24159 & w24160) | (w24159 & w35863) | (w24160 & w35863);
assign w32680 = w8520 & b_60;
assign w32681 = w24289 & w35864;
assign w32682 = w7607 & b_63;
assign w32683 = (~w24300 & w29820) | (~w24300 & w35865) | (w29820 & w35865);
assign w32684 = (w29747 & w35866) | (w29747 & w35867) | (w35866 & w35867);
assign w32685 = ~w24300 & w35868;
assign w32686 = (~a_50 & w24300) | (~a_50 & w35869) | (w24300 & w35869);
assign w32687 = ~w24304 & w24204;
assign w32688 = (~w24304 & w24204) | (~w24304 & w35870) | (w24204 & w35870);
assign w32689 = w24304 & ~w24204;
assign w32690 = ~w24204 & w35871;
assign w32691 = w24137 & ~w24212;
assign w32692 = (w24235 & w24236) | (w24235 & w35872) | (w24236 & w35872);
assign w32693 = w9528 & b_58;
assign w32694 = w24323 & w35873;
assign w32695 = w24271 & ~w24260;
assign w32696 = w10556 & b_55;
assign w32697 = (a_59 & ~w24334) | (a_59 & w35874) | (~w24334 & w35874);
assign w32698 = a_59 & ~w27707;
assign w32699 = a_59 & ~w32697;
assign w32700 = w27707 & a_59;
assign w32701 = w11614 & b_52;
assign w32702 = (a_62 & ~w24344) | (a_62 & w35875) | (~w24344 & w35875);
assign w32703 = a_62 & ~w27708;
assign w32704 = a_62 & ~w32702;
assign w32705 = w27708 & a_62;
assign w32706 = a_63 & b_50;
assign w32707 = w24250 & w24360;
assign w32708 = ~w32707 & w24360;
assign w32709 = w24363 & ~w24350;
assign w32710 = w24369 & ~w24330;
assign w32711 = w24330 & ~w24369;
assign w32712 = w8520 & b_61;
assign w32713 = w24383 & w35876;
assign w32714 = (w24295 & w24281) | (w24295 & w35877) | (w24281 & w35877);
assign w32715 = ~w24305 & ~w24397;
assign w32716 = w24305 & w24397;
assign w32717 = w8520 & b_62;
assign w32718 = (~w9770 & w35878) | (~w9770 & w35879) | (w35878 & w35879);
assign w32719 = ~w24406 & a_53;
assign w32720 = w24406 & a_53;
assign w32721 = w9528 & b_59;
assign w32722 = w24417 & w35880;
assign w32723 = w10556 & b_56;
assign w32724 = w24428 & w35881;
assign w32725 = a_63 & b_51;
assign w32726 = w24174 & ~w24355;
assign w32727 = w11614 & b_53;
assign w32728 = (w9776 & w35882) | (w9776 & w35883) | (w35882 & w35883);
assign w32729 = w24361 & w24452;
assign w32730 = ~w24361 & ~w24452;
assign w32731 = w24461 & ~w24423;
assign w32732 = w24434 & ~w24453;
assign w32733 = a_63 & b_52;
assign w32734 = ~w24485 & ~w24486;
assign w32735 = ~w24438 & w35884;
assign w32736 = ~w24486 & ~w32734;
assign w32737 = ~w24486 & ~w32735;
assign w32738 = ~w32735 & w32734;
assign w32739 = w11614 & b_54;
assign w32740 = w24494 & w35885;
assign w32741 = w24490 & w24500;
assign w32742 = ~w24490 & ~w24500;
assign w32743 = w10556 & b_57;
assign w32744 = w24507 & w35886;
assign w32745 = w9528 & b_60;
assign w32746 = w24523 & w35887;
assign w32747 = w8520 & b_63;
assign w32748 = (~w24534 & w29820) | (~w24534 & w35888) | (w29820 & w35888);
assign w32749 = (w29747 & w35889) | (w29747 & w35890) | (w35889 & w35890);
assign w32750 = ~w24534 & w35891;
assign w32751 = (~a_53 & w24534) | (~a_53 & w35892) | (w24534 & w35892);
assign w32752 = w24459 & ~w24538;
assign w32753 = (w24538 & w24424) | (w24538 & w35893) | (w24424 & w35893);
assign w32754 = w24412 & ~w24466;
assign w32755 = w24533 & ~w24539;
assign w32756 = w9528 & b_61;
assign w32757 = w24558 & w35894;
assign w32758 = w24490 & ~w24500;
assign w32759 = w10556 & b_58;
assign w32760 = w24573 & w35895;
assign w32761 = a_63 & b_53;
assign w32762 = w11614 & b_55;
assign w32763 = a_62 & ~w27709;
assign w32764 = w26964 & a_62;
assign w32765 = (~w10452 & w35896) | (~w10452 & w35897) | (w35896 & w35897);
assign w32766 = w24567 & w24613;
assign w32767 = ~w24567 & ~w24613;
assign w32768 = w9528 & b_62;
assign w32769 = (~w9770 & w35898) | (~w9770 & w35899) | (w35898 & w35899);
assign w32770 = ~w24625 & a_56;
assign w32771 = w24625 & a_56;
assign w32772 = w24569 & ~w24606;
assign w32773 = w10556 & b_59;
assign w32774 = w24636 & w35900;
assign w32775 = w24489 & ~w24599;
assign w32776 = a_63 & b_54;
assign w32777 = w24585 & ~w24647;
assign w32778 = w11614 & b_56;
assign w32779 = ~w24652 & ~w11623;
assign w32780 = ~w24656 & ~w24657;
assign w32781 = ~a_62 & ~w24657;
assign w32782 = ~a_62 & w32780;
assign w32783 = (w10476 & w35901) | (w10476 & w35902) | (w35901 & w35902);
assign w32784 = (~w10476 & w35903) | (~w10476 & w35904) | (w35903 & w35904);
assign w32785 = w35905 & w24643;
assign w32786 = w24567 & ~w24613;
assign w32787 = w11614 & b_57;
assign w32788 = (w9770 & w35906) | (w9770 & w35907) | (w35906 & w35907);
assign w32789 = w27711 & a_62;
assign w32790 = (~w9770 & w35908) | (~w9770 & w35909) | (w35908 & w35909);
assign w32791 = a_63 & b_55;
assign w32792 = ~w24705 & w24706;
assign w32793 = w24705 & ~w24706;
assign w32794 = w10556 & b_60;
assign w32795 = w24713 & w35910;
assign w32796 = w9528 & b_63;
assign w32797 = (~w24724 & w29820) | (~w24724 & w35911) | (w29820 & w35911);
assign w32798 = (w29747 & w35912) | (w29747 & w35913) | (w35912 & w35913);
assign w32799 = ~w24724 & w35914;
assign w32800 = (~a_56 & w24724) | (~a_56 & w35915) | (w24724 & w35915);
assign w32801 = w24663 & ~w24728;
assign w32802 = (w24728 & w24643) | (w24728 & w35916) | (w24643 & w35916);
assign w32803 = (w24631 & w24632) | (w24631 & w35917) | (w24632 & w35917);
assign w32804 = (~w32793 & w35918) | (~w32793 & w35919) | (w35918 & w35919);
assign w32805 = w10556 & b_61;
assign w32806 = w24747 & w35920;
assign w32807 = a_63 & b_56;
assign w32808 = w24762 & ~w24646;
assign w32809 = w24702 & ~w24699;
assign w32810 = w24768 & ~w24699;
assign w32811 = w24768 & w32809;
assign w32812 = ~w24768 & w24699;
assign w32813 = ~w24768 & ~w32809;
assign w32814 = w11614 & b_58;
assign w32815 = w24775 & w35921;
assign w32816 = w35922 & w24743;
assign w32817 = w24782 & ~w24783;
assign w32818 = ~w24782 & ~w24783;
assign w32819 = ~w24782 & w32817;
assign w32820 = w24723 & ~w24729;
assign w32821 = ~w24787 & w24788;
assign w32822 = w24787 & ~w24788;
assign w32823 = w24781 & ~w24770;
assign w32824 = a_63 & b_57;
assign w32825 = ~w24761 & ~w24798;
assign w32826 = w24761 & w24798;
assign w32827 = w11614 & b_59;
assign w32828 = ~w24802 & ~w11623;
assign w32829 = ~w24806 & ~w24807;
assign w32830 = ~a_62 & ~w24807;
assign w32831 = ~a_62 & w32829;
assign w32832 = (w11901 & w35923) | (w11901 & w35924) | (w35923 & w35924);
assign w32833 = (~w11901 & w35925) | (~w11901 & w35926) | (w35925 & w35926);
assign w32834 = w10556 & b_62;
assign w32835 = (~w9770 & w35927) | (~w9770 & w35928) | (w35927 & w35928);
assign w32836 = ~w24818 & a_59;
assign w32837 = w24818 & a_59;
assign w32838 = (w24782 & w24743) | (w24782 & w35929) | (w24743 & w35929);
assign w32839 = (w24824 & w24795) | (w24824 & w35930) | (w24795 & w35930);
assign w32840 = a_63 & b_58;
assign w32841 = (w24765 & w35931) | (w24765 & w35932) | (w35931 & w35932);
assign w32842 = ~w24841 & ~w24842;
assign w32843 = ~w24841 & w32841;
assign w32844 = ~w24842 & ~w32842;
assign w32845 = (~w24842 & ~w32841) | (~w24842 & w35933) | (~w32841 & w35933);
assign w32846 = (~w32841 & w32842) | (~w32841 & w35934) | (w32842 & w35934);
assign w32847 = w11614 & b_60;
assign w32848 = w24851 & w35935;
assign w32849 = w10556 & b_63;
assign w32850 = ~w10565 & ~w24858;
assign w32851 = w24847 & ~w24864;
assign w32852 = a_63 & b_59;
assign w32853 = w11614 & b_61;
assign w32854 = w24891 & w35936;
assign w32855 = w35937 & w24893;
assign w32856 = w24845 & ~w24898;
assign w32857 = a_63 & b_60;
assign w32858 = w24884 & ~w24916;
assign w32859 = w11614 & b_62;
assign w32860 = (w9770 & w35938) | (w9770 & w35939) | (w35938 & w35939);
assign w32861 = w24924 & a_62;
assign w32862 = (~a_62 & ~w24923) | (~a_62 & w35940) | (~w24923 & w35940);
assign w32863 = w24931 & w24898;
assign w32864 = w24931 & ~w32856;
assign w32865 = ~w24920 & ~w24918;
assign w32866 = a_63 & b_61;
assign w32867 = w11614 & b_63;
assign w32868 = (~w24946 & w29820) | (~w24946 & w35941) | (w29820 & w35941);
assign w32869 = (w29747 & w35942) | (w29747 & w35943) | (w35942 & w35943);
assign w32870 = ~w24946 & w35944;
assign w32871 = (~a_62 & w24946) | (~a_62 & w35940) | (w24946 & w35940);
assign w32872 = (~w25221 & w35945) | (~w25221 & w35946) | (w35945 & w35946);
assign w32873 = (w25216 & w35947) | (w25216 & w35948) | (w35947 & w35948);
assign w32874 = ~w24945 & ~w24943;
assign w32875 = a_63 & b_62;
assign w32876 = w24969 & w24943;
assign w32877 = w24969 & ~w32874;
assign w32878 = ~w24969 & ~w24943;
assign w32879 = ~w24969 & w32874;
assign w32880 = (~w25221 & w35949) | (~w25221 & w35950) | (w35949 & w35950);
assign w32881 = (w25216 & w35951) | (w25216 & w35952) | (w35951 & w35952);
assign w32882 = w24915 & ~w24964;
assign w32883 = a_63 & b_63;
assign w32884 = (~w25221 & w35953) | (~w25221 & w35954) | (w35953 & w35954);
assign w32885 = (w25216 & w35955) | (w25216 & w35956) | (w35955 & w35956);
assign w32886 = (w25221 & w35957) | (w25221 & w35958) | (w35957 & w35958);
assign w32887 = (~w25216 & w35959) | (~w25216 & w35960) | (w35959 & w35960);
assign w32888 = ~w2529 & ~w421;
assign w32889 = ~w2681 & ~w989;
assign w32890 = ~w2700 & ~w660;
assign w32891 = ~w2718 & ~w421;
assign w32892 = ~w2541 & ~w2539;
assign w32893 = ~w2883 & ~w660;
assign w32894 = ~w3059 & ~w660;
assign w32895 = ~w3219 & ~w1697;
assign w32896 = ~w3262 & ~w660;
assign w32897 = ~w3280 & ~w421;
assign w32898 = ~w3494 & ~w421;
assign w32899 = ~w3637 & ~w1697;
assign w32900 = ~w3693 & ~w421;
assign w32901 = ~w3870 & ~w989;
assign w32902 = ~w3888 & ~w660;
assign w32903 = ~w3906 & ~w421;
assign w32904 = ~w3923 & ~w242;
assign w32905 = w3716 & w35961;
assign w32906 = ~w3981 & ~w242;
assign w32907 = ~w4896 & ~w242;
assign w32908 = ~w5379 & ~w242;
assign w32909 = ~w5390 & ~w421;
assign w32910 = ~w5634 & ~w421;
assign w32911 = ~w5830 & ~w242;
assign w32912 = ~w6373 & ~w242;
assign w32913 = ~w6636 & ~w242;
assign w32914 = ~w6391 & ~w6390;
assign w32915 = ~w7214 & ~w421;
assign w32916 = ~w7502 & ~w421;
assign w32917 = ~w7520 & ~w242;
assign w32918 = ~w7795 & ~w421;
assign w32919 = ~w7813 & ~w242;
assign w32920 = ~w8099 & ~w421;
assign w32921 = ~w8413 & ~w660;
assign w32922 = ~w8431 & ~w421;
assign w32923 = ~w8714 & ~w660;
assign w32924 = ~w9032 & ~w660;
assign w32925 = w8765 & w35962;
assign w32926 = ~w9381 & ~w660;
assign w32927 = ~w9721 & ~w660;
assign w32928 = ~w9760 & ~w9758;
assign w32929 = ~w10061 & ~w660;
assign w32930 = ~w10078 & ~w421;
assign w32931 = ~w10096 & ~w10095;
assign w32932 = ~w14123 & ~w14121;
assign w32933 = ~w16802 & ~w16800;
assign w32934 = ~w17121 & w16800;
assign w32935 = (~w17121 & w16801) | (~w17121 & w35963) | (w16801 & w35963);
assign w32936 = (~w17118 & w25479) | (~w17118 & ~w16800) | (w25479 & ~w16800);
assign w32937 = (~w16801 & w35964) | (~w16801 & w35965) | (w35964 & w35965);
assign w32938 = (~w17710 & ~w17711) | (~w17710 & w17707) | (~w17711 & w17707);
assign w32939 = (~w17417 & w35966) | (~w17417 & w35967) | (w35966 & w35967);
assign w32940 = ~w18272 & w35968;
assign w32941 = w18548 & ~w18545;
assign w32942 = ~w18545 & ~w25480;
assign w32943 = ~w18815 & ~w18813;
assign w32944 = ~w19077 & ~w19079;
assign w32945 = ~w19077 & ~w25179;
assign w32946 = w19338 & w19077;
assign w32947 = w19338 & w19079;
assign w32948 = ~w19337 & ~w19338;
assign w32949 = (w19582 & w19338) | (w19582 & w25481) | (w19338 & w25481);
assign w32950 = w19337 & w19582;
assign w32951 = (w19582 & w25481) | (w19582 & w19338) | (w25481 & w19338);
assign w32952 = (~w19581 & w26969) | (~w19581 & ~w19337) | (w26969 & ~w19337);
assign w32953 = (~w19338 & w35969) | (~w19338 & w26970) | (w35969 & w26970);
assign w32954 = w26970 | w26969;
assign w32955 = (w26969 & w26970) | (w26969 & ~w19338) | (w26970 & ~w19338);
assign w32956 = w20073 & w19828;
assign w32957 = ~w20308 & w20071;
assign w32958 = ~w20308 & ~w25482;
assign w32959 = w20535 & ~w25483;
assign w32960 = (~w20533 & w26867) | (~w20533 & ~w20305) | (w26867 & ~w20305);
assign w32961 = (~w20533 & w26867) | (~w20533 & w25483) | (w26867 & w25483);
assign w32962 = (w20754 & w26866) | (w20754 & w26972) | (w26866 & w26972);
assign w32963 = (w26972 & w26973) | (w26972 & w20305) | (w26973 & w20305);
assign w32964 = (w26972 & w26973) | (w26972 & ~w25483) | (w26973 & ~w25483);
assign w32965 = ~w21183 & w20970;
assign w32966 = (~w21180 & w25485) | (~w21180 & ~w20969) | (w25485 & ~w20969);
assign w32967 = (~w21180 & w25485) | (~w21180 & ~w20970) | (w25485 & ~w20970);
assign w32968 = (~w21387 & w25485) | (~w21387 & w26868) | (w25485 & w26868);
assign w32969 = (~w21584 & w21389) | (~w21584 & w35970) | (w21389 & w35970);
assign w32970 = (~w21584 & w26742) | (~w21584 & w35970) | (w26742 & w35970);
assign w32971 = ~w21581 & ~w32969;
assign w32972 = (~w26742 & w26870) | (~w26742 & w35971) | (w26870 & w35971);
assign w32973 = (~w21780 & w26974) | (~w21780 & w32969) | (w26974 & w32969);
assign w32974 = (w26742 & w35972) | (w26742 & w35973) | (w35972 & w35973);
assign w32975 = (~w21780 & ~w21584) | (~w21780 & w26974) | (~w21584 & w26974);
assign w32976 = (~w21777 & w26975) | (~w21777 & ~w21581) | (w26975 & ~w21581);
assign w32977 = (w21584 & w35974) | (w21584 & w32976) | (w35974 & w32976);
assign w32978 = ~w22142 & w35975;
assign w32979 = ~w22143 & w25486;
assign w32980 = (w25486 & ~w22143) | (w25486 & w22321) | (~w22143 & w22321);
assign w32981 = (w22143 & w35976) | (w22143 & w32983) | (w35976 & w32983);
assign w32982 = (~w22319 & w22143) | (~w22319 & w32983) | (w22143 & w32983);
assign w32983 = (~w22319 & ~w22140) | (~w22319 & w35976) | (~w22140 & w35976);
assign w32984 = ~w22142 & w35977;
assign w32985 = (w22140 & w35978) | (w22140 & w35979) | (w35978 & w35979);
assign w32986 = (w22142 & w35980) | (w22142 & w35981) | (w35980 & w35981);
assign w32987 = (~w22143 & w35979) | (~w22143 & w35982) | (w35979 & w35982);
assign w32988 = (~w22143 & w35978) | (~w22143 & w35982) | (w35978 & w35982);
assign w32989 = (w22143 & w35983) | (w22143 & w32991) | (w35983 & w32991);
assign w32990 = (w22143 & w35984) | (w22143 & w32991) | (w35984 & w32991);
assign w32991 = (w26744 & w26745) | (w26744 & ~w25486) | (w26745 & ~w25486);
assign w32992 = (~w22142 & w35985) | (~w22142 & w35986) | (w35985 & w35986);
assign w32993 = ~w22823 & ~w26976;
assign w32994 = ~w22823 & ~w26977;
assign w32995 = ~w23126 & ~w23127;
assign w32996 = ~w23270 & ~w25347;
assign w32997 = (w23413 & w23272) | (w23413 & w25489) | (w23272 & w25489);
assign w32998 = (w23413 & w25489) | (w23413 & w23272) | (w25489 & w23272);
assign w32999 = (w23413 & w25489) | (w23413 & w25347) | (w25489 & w25347);
assign w33000 = ~w23411 & ~w32998;
assign w33001 = (~w25347 & w26083) | (~w25347 & w35987) | (w26083 & w35987);
assign w33002 = (~w23411 & w26083) | (~w23411 & ~w23270) | (w26083 & ~w23270);
assign w33003 = (~w23411 & w26083) | (~w23411 & w25488) | (w26083 & w25488);
assign w33004 = (~w26083 & w26084) | (~w26083 & w35988) | (w26084 & w35988);
assign w33005 = (~w25488 & w26084) | (~w25488 & w35989) | (w26084 & w35989);
assign w33006 = (w23544 & w26084) | (w23544 & w32998) | (w26084 & w32998);
assign w33007 = (w25347 & w35990) | (w25347 & w35991) | (w35990 & w35991);
assign w33008 = (w26510 & w26511) | (w26510 & ~w32998) | (w26511 & ~w32998);
assign w33009 = (~w25347 & w35992) | (~w25347 & w35993) | (w35992 & w35993);
assign w33010 = (w26083 & w26511) | (w26083 & w35994) | (w26511 & w35994);
assign w33011 = (w25488 & w26511) | (w25488 & w35995) | (w26511 & w35995);
assign w33012 = (~w26083 & w35996) | (~w26083 & w35997) | (w35996 & w35997);
assign w33013 = (~w25488 & w35996) | (~w25488 & w35998) | (w35996 & w35998);
assign w33014 = (w32998 & w35999) | (w32998 & w36000) | (w35999 & w36000);
assign w33015 = w23676 & ~w33009;
assign w33016 = (~w32998 & w36001) | (~w32998 & w36002) | (w36001 & w36002);
assign w33017 = (~w23674 & w26748) | (~w23674 & w33009) | (w26748 & w33009);
assign w33018 = (w32998 & w36003) | (w32998 & w36004) | (w36003 & w36004);
assign w33019 = (w26872 & w26873) | (w26872 & ~w33009) | (w26873 & ~w33009);
assign w33020 = (w23910 & w23798) | (w23910 & w36005) | (w23798 & w36005);
assign w33021 = (w23910 & w26872) | (w23910 & w36005) | (w26872 & w36005);
assign w33022 = w24125 & w24022;
assign w33023 = (~w24124 & w25723) | (~w24124 & ~w24021) | (w25723 & ~w24021);
assign w33024 = (~w24124 & w25723) | (~w24124 & ~w24022) | (w25723 & ~w24022);
assign w33025 = ~w24221 & ~w24222;
assign w33026 = ~w24221 & ~w26085;
assign w33027 = ~w24221 & ~w26086;
assign w33028 = (w24315 & w26512) | (w24315 & w24222) | (w26512 & w24222);
assign w33029 = (w24315 & w26512) | (w24315 & w26085) | (w26512 & w26085);
assign w33030 = (w24315 & w26512) | (w24315 & w26086) | (w26512 & w26086);
assign w33031 = (w26749 & w26750) | (w26749 & ~w24222) | (w26750 & ~w24222);
assign w33032 = (w26749 & w26750) | (w26749 & ~w26085) | (w26750 & ~w26085);
assign w33033 = (w26749 & w26750) | (w26749 & ~w26086) | (w26750 & ~w26086);
assign w33034 = (w26085 & w36006) | (w26085 & w36007) | (w36006 & w36007);
assign w33035 = w24400 & ~w33031;
assign w33036 = (~w26085 & w36008) | (~w26085 & w36009) | (w36008 & w36009);
assign w33037 = (~w24399 & w26874) | (~w24399 & w33031) | (w26874 & w33031);
assign w33038 = (w26085 & w36010) | (w26085 & w36011) | (w36010 & w36011);
assign w33039 = (w26981 & w26982) | (w26981 & ~w33031) | (w26982 & ~w33031);
assign w33040 = ~w24475 & ~w26981;
assign w33041 = ~w24475 & ~w26982;
assign w33042 = w24475 & w24549;
assign w33043 = (w24549 & w26981) | (w24549 & w33042) | (w26981 & w33042);
assign w33044 = (w24549 & w26982) | (w24549 & w33042) | (w26982 & w33042);
assign w33045 = w24682 & ~w24679;
assign w33046 = w24679 & w24739;
assign w33047 = (w24739 & w25724) | (w24739 & ~w24682) | (w25724 & ~w24682);
assign w33048 = w26088 | w26087;
assign w33049 = (w26087 & w26088) | (w26087 & w24682) | (w26088 & w24682);
assign w33050 = (w24791 & w24739) | (w24791 & w36012) | (w24739 & w36012);
assign w33051 = w24791 & ~w26088;
assign w33052 = (~w24790 & w26513) | (~w24790 & w26087) | (w26513 & w26087);
assign w33053 = (~w24790 & w26513) | (~w24790 & w26088) | (w26513 & w26088);
assign w33054 = w24832 & w24790;
assign w33055 = (w24832 & w24791) | (w24832 & w33054) | (w24791 & w33054);
assign w33056 = ~w24874 & w24831;
assign w33057 = (~w24874 & w24832) | (~w24874 & w33056) | (w24832 & w33056);
assign w33058 = (~w26751 & w33056) | (~w26751 & w36013) | (w33056 & w36013);
assign w33059 = (~w26513 & w33056) | (~w26513 & w36014) | (w33056 & w36014);
assign w33060 = (~w24871 & ~w24831) | (~w24871 & w36015) | (~w24831 & w36015);
assign w33061 = ~w24871 & ~w33057;
assign w33062 = ~w24871 & ~w33058;
assign w33063 = ~w24871 & ~w33059;
assign w33064 = ~w24908 & ~w33060;
assign w33065 = (~w24908 & w33057) | (~w24908 & w36016) | (w33057 & w36016);
assign w33066 = (~w24908 & w33058) | (~w24908 & w36016) | (w33058 & w36016);
assign w33067 = (~w24908 & w33059) | (~w24908 & w36016) | (w33059 & w36016);
assign w33068 = (~w24905 & w33060) | (~w24905 & w36017) | (w33060 & w36017);
assign w33069 = (~w33057 & w36017) | (~w33057 & w36018) | (w36017 & w36018);
assign w33070 = (~w33058 & w36017) | (~w33058 & w36018) | (w36017 & w36018);
assign w33071 = (~w33059 & w36017) | (~w33059 & w36018) | (w36017 & w36018);
assign w33072 = (~w33060 & w36019) | (~w33060 & w36020) | (w36019 & w36020);
assign w33073 = (w33057 & w36020) | (w33057 & w36021) | (w36020 & w36021);
assign w33074 = ~w24956 & ~w24954;
assign w33075 = ~w24939 & w36022;
assign w33076 = ~w24972 & ~w24970;
assign w33077 = ~w24970 & ~w33075;
assign w33078 = b_4 & a_26;
assign w33079 = ~w20073 & ~w20071;
assign w33080 = ~w8081 & ~w660;
assign w33081 = w418 & w36023;
assign w33082 = ~w8117 & ~w242;
assign w33083 = ~w8134 & ~w102;
assign w33084 = ~w7855 & ~w7280;
assign w33085 = ~w8193 & ~w242;
assign w33086 = ~w8204 & ~w1298;
assign w33087 = ~w7974 & ~w7973;
assign w33088 = ~w8397 & ~w989;
assign w33089 = w657 & w36024;
assign w33090 = w418 & w36025;
assign w33091 = ~w8696 & ~w989;
assign w33092 = w657 & w36026;
assign w33093 = ~w8732 & ~w421;
assign w33094 = ~w8748 & ~w242;
assign w33095 = ~w9014 & ~w989;
assign w33096 = w657 & w36027;
assign w33097 = ~w9050 & ~w421;
assign w33098 = ~w9067 & ~w242;
assign w33099 = ~w9140 & ~w421;
assign w33100 = ~w9363 & ~w989;
assign w33101 = w657 & w36028;
assign w33102 = ~w9456 & ~w242;
assign w33103 = ~w9703 & ~w989;
assign w33104 = w657 & w36029;
assign w33105 = ~w9736 & ~w421;
assign w33106 = ~w10043 & ~w989;
assign w33107 = w657 & w36030;
assign w33108 = w418 & w36031;
assign w33109 = ~w10148 & ~w421;
assign w33110 = ~w10158 & ~w660;
assign w33111 = ~w10379 & ~w1298;
assign w33112 = ~w10751 & ~w1298;
assign w33113 = ~w11081 & ~w1298;
assign w33114 = ~w11115 & ~w660;
assign w33115 = ~w11808 & ~w1697;
assign w33116 = ~w12194 & ~w989;
assign w33117 = w102 & ~w29581;
assign w33118 = w102 & ~w29580;
assign w33119 = ~w11897 & ~w11192;
assign w33120 = ~w12941 & ~w2161;
assign w33121 = (w25505 & w25506) | (w25505 & w29473) | (w25506 & w29473);
assign w33122 = (w25505 & w25506) | (w25505 & w29472) | (w25506 & w29472);
assign w33123 = ~w14903 & ~w1697;
assign w33124 = ~w15892 & ~w2161;
assign w33125 = ~w21698 & ~w7616;
assign w33126 = ~w21856 & ~w8529;
assign w33127 = ~w21872 & ~w7616;
assign w33128 = ~w22362 & ~w10565;
assign w33129 = ~w22381 & ~w9537;
assign w33130 = ~w22399 & ~w8529;
assign w33131 = ~w22554 & ~w9537;
assign w33132 = ~w22571 & ~w8529;
assign w33133 = ~w22866 & ~w10565;
assign w33134 = ~w23853 & ~w11623;
assign w33135 = w23852 & w25711;
assign w33136 = w23852 & w25710;
assign w33137 = ~w24442 & ~w11623;
assign w33138 = (w33060 & w36032) | (w33060 & w36033) | (w36032 & w36033);
assign w33139 = (~w33057 & w36033) | (~w33057 & w36034) | (w36033 & w36034);
assign w33140 = (w25328 & ~w25327) | (w25328 & w36035) | (~w25327 & w36035);
assign w33141 = (w25328 & w25329) | (w25328 & w24935) | (w25329 & w24935);
assign w33142 = (w33060 & w36036) | (w33060 & w36037) | (w36036 & w36037);
assign w33143 = (~w33057 & w36037) | (~w33057 & w36038) | (w36037 & w36038);
assign w33144 = (w25332 & w25333) | (w25332 & w24935) | (w25333 & w24935);
assign w33145 = (w33060 & w36039) | (w33060 & w36040) | (w36039 & w36040);
assign w33146 = (~w33057 & w36040) | (~w33057 & w36041) | (w36040 & w36041);
assign w33147 = ~w20307 & ~w20305;
assign w33148 = ~w21182 & ~w21180;
assign w33149 = (a_26 & ~w2158) | (a_26 & w36042) | (~w2158 & w36042);
assign w33150 = w986 & w36043;
assign w33151 = (a_14 & ~w657) | (a_14 & w36044) | (~w657 & w36044);
assign w33152 = ~w8789 & ~w8182;
assign w33153 = ~w9197 & ~w4502;
assign w33154 = ~w9330 & ~w1697;
assign w33155 = w986 & w36045;
assign w33156 = ~w9685 & ~w1298;
assign w33157 = w986 & w36046;
assign w33158 = w418 & w36047;
assign w33159 = ~w9817 & ~w1697;
assign w33160 = ~w9827 & ~w2161;
assign w33161 = ~w10025 & ~w1298;
assign w33162 = w986 & w36048;
assign w33163 = w418 & w36049;
assign w33164 = w657 & w36050;
assign w33165 = ~w10346 & ~w2161;
assign w33166 = w1295 & w36051;
assign w33167 = ~w10397 & ~w989;
assign w33168 = ~w10503 & ~w421;
assign w33169 = ~w10733 & ~w1697;
assign w33170 = w1295 & w36052;
assign w33171 = ~w10769 & ~w989;
assign w33172 = ~w10786 & ~w660;
assign w33173 = ~w11063 & ~w1697;
assign w33174 = w1295 & w36053;
assign w33175 = ~w11098 & ~w989;
assign w33176 = w657 & w36054;
assign w33177 = ~w11235 & ~w660;
assign w33178 = ~w11246 & ~w989;
assign w33179 = ~w11258 & ~w2642;
assign w33180 = ~w11466 & ~w1697;
assign w33181 = ~w11484 & ~w1298;
assign w33182 = ~w11757 & ~w3198;
assign w33183 = ~w11790 & ~w2161;
assign w33184 = w1694 & w36055;
assign w33185 = ~w12160 & ~w1697;
assign w33186 = ~w12177 & ~w1298;
assign w33187 = w986 & w36056;
assign w33188 = ~w12300 & ~w989;
assign w33189 = w1295 & w36057;
assign w33190 = ~w12322 & ~w1697;
assign w33191 = ~w12334 & ~w3198;
assign w33192 = ~w12546 & ~w2161;
assign w33193 = ~w12703 & ~w989;
assign w33194 = ~w12714 & ~w1298;
assign w33195 = ~w12923 & ~w2642;
assign w33196 = w2158 & w36058;
assign w33197 = ~w13049 & ~w1298;
assign w33198 = ~w14048 & ~w989;
assign w33199 = ~w15227 & ~w3198;
assign w33200 = w2158 & w36059;
assign w33201 = w15552 & w36060;
assign w33202 = w15831 & ~w30608;
assign w33203 = w15887 & w16125;
assign w33204 = ~w16242 & ~w2642;
assign w33205 = ~w17766 & ~w2642;
assign w33206 = ~w20479 & ~w5965;
assign w33207 = ~w20677 & ~w5965;
assign w33208 = ~w21117 & ~w6764;
assign w33209 = ~w21298 & ~w6764;
assign w33210 = w7613 & w36061;
assign w33211 = ~w21797 & ~w9537;
assign w33212 = w8526 & w36062;
assign w33213 = w7613 & w36063;
assign w33214 = ~w21889 & ~w6764;
assign w33215 = ~w22017 & ~w11623;
assign w33216 = w10562 & w36064;
assign w33217 = w9534 & w36065;
assign w33218 = w8526 & w36066;
assign w33219 = ~w22509 & ~w11623;
assign w33220 = ~w22536 & ~w10565;
assign w33221 = w9534 & w36067;
assign w33222 = w8526 & w36068;
assign w33223 = ~w22589 & ~w7616;
assign w33224 = ~w22744 & ~w9537;
assign w33225 = w10562 & w36069;
assign w33226 = ~w22885 & ~w9537;
assign w33227 = ~w23018 & ~w10565;
assign w33228 = ~w23035 & ~w9537;
assign w33229 = w11620 & w36070;
assign w33230 = (a_62 & ~w11620) | (a_62 & w36071) | (~w11620 & w36071);
assign w33231 = (w25316 & w25315) | (w25316 & ~w33043) | (w25315 & ~w33043);
assign w33232 = (~w26982 & w33233) | (~w26982 & w33234) | (w33233 & w33234);
assign w33233 = (w25316 & w25315) | (w25316 & ~w24549) | (w25315 & ~w24549);
assign w33234 = (w25316 & w25315) | (w25316 & ~w33042) | (w25315 & ~w33042);
assign w33235 = (w25320 & w25319) | (w25320 & ~w33043) | (w25319 & ~w33043);
assign w33236 = (~w26982 & w33237) | (~w26982 & w33238) | (w33237 & w33238);
assign w33237 = (w25320 & w25319) | (w25320 & ~w24549) | (w25319 & ~w24549);
assign w33238 = (w25320 & w25319) | (w25320 & ~w33042) | (w25319 & ~w33042);
assign w33239 = (w25324 & w25323) | (w25324 & ~w33043) | (w25323 & ~w33043);
assign w33240 = (~w26982 & w33241) | (~w26982 & w33242) | (w33241 & w33242);
assign w33241 = (w25324 & w25323) | (w25324 & ~w24549) | (w25323 & ~w24549);
assign w33242 = (w25324 & w25323) | (w25324 & ~w33042) | (w25323 & ~w33042);
assign w33243 = w25327 & ~w24957;
assign w33244 = (~w24957 & w25327) | (~w24957 & ~w24935) | (w25327 & ~w24935);
assign w33245 = (~w33060 & w36072) | (~w33060 & w36073) | (w36072 & w36073);
assign w33246 = (w33057 & w36073) | (w33057 & w36074) | (w36073 & w36074);
assign w33247 = w25331 & w25330;
assign w33248 = (w25330 & w25331) | (w25330 & ~w24935) | (w25331 & ~w24935);
assign w33249 = (~w33060 & w36075) | (~w33060 & w36076) | (w36075 & w36076);
assign w33250 = (w33057 & w36076) | (w33057 & w36077) | (w36076 & w36077);
assign w33251 = w7864 & ~w7552;
assign w33252 = b_4 & a_29;
assign w33253 = (a_29 & ~w2639) | (a_29 & w36078) | (~w2639 & w36078);
assign w33254 = ~w9978 & ~w3198;
assign w33255 = w1295 & w36079;
assign w33256 = ~w10194 & ~w5199;
assign w33257 = w2158 & w36080;
assign w33258 = ~w10363 & ~w1697;
assign w33259 = w986 & w36081;
assign w33260 = ~w9794 & ~w9772;
assign w33261 = ~w10435 & ~w10434;
assign w33262 = ~w10492 & ~w242;
assign w33263 = w418 & w36082;
assign w33264 = ~w10682 & ~w3198;
assign w33265 = ~w10715 & ~w2161;
assign w33266 = w1694 & w36083;
assign w33267 = w986 & w36084;
assign w33268 = w657 & w36085;
assign w33269 = ~w10842 & ~w421;
assign w33270 = ~w10853 & ~w2161;
assign w33271 = ~w10868 & ~w5965;
assign w33272 = ~w11023 & ~w3198;
assign w33273 = w1694 & w36086;
assign w33274 = w986 & w36087;
assign w33275 = ~w11224 & ~w421;
assign w33276 = w657 & w36088;
assign w33277 = w986 & w36089;
assign w33278 = w2639 & w36090;
assign w33279 = ~w11280 & ~w5965;
assign w33280 = ~w11409 & ~w3806;
assign w33281 = ~w11450 & ~w2161;
assign w33282 = w1694 & w36091;
assign w33283 = w1295 & w36092;
assign w33284 = ~w11561 & ~w660;
assign w33285 = ~w11739 & ~w3806;
assign w33286 = w3195 & w36093;
assign w33287 = w2158 & w36094;
assign w33288 = ~w11826 & ~w1298;
assign w33289 = ~w11842 & ~w989;
assign w33290 = ~w11921 & ~w660;
assign w33291 = ~w12089 & ~w3806;
assign w33292 = ~w12107 & ~w3198;
assign w33293 = ~w12142 & ~w2161;
assign w33294 = w1694 & w36095;
assign w33295 = w1295 & w36096;
assign w33296 = (a_17 & ~w986) | (a_17 & w36097) | (~w986 & w36097);
assign w33297 = w986 & w36098;
assign w33298 = ~w1298 & a_20;
assign w33299 = w1694 & w36099;
assign w33300 = w3195 & w36100;
assign w33301 = ~w12506 & ~w3806;
assign w33302 = ~w12530 & ~w2642;
assign w33303 = w2158 & w36101;
assign w33304 = w986 & w36102;
assign w33305 = w1295 & w36103;
assign w33306 = ~w12725 & ~w3198;
assign w33307 = ~w12898 & ~w3806;
assign w33308 = w2639 & w36104;
assign w33309 = w1295 & w36105;
assign w33310 = ~w13276 & ~w2161;
assign w33311 = ~w13293 & ~w1697;
assign w33312 = ~w13777 & ~w1298;
assign w33313 = w986 & w36106;
assign w33314 = w657 & w36107;
assign w33315 = ~w660 & a_14;
assign w33316 = ~w14181 & ~w1298;
assign w33317 = ~w14023 & w36108;
assign w33318 = w14025 & w14036;
assign w33319 = ~w14196 & ~w1697;
assign w33320 = w1694 & w36109;
assign w33321 = ~w15183 & ~w989;
assign w33322 = ~w15211 & ~w2161;
assign w33323 = w3195 & w36110;
assign w33324 = ~w15583 & ~w2642;
assign w33325 = ~w16215 & ~w1298;
assign w33326 = w2639 & w36111;
assign w33327 = ~w17678 & ~w3198;
assign w33328 = w2639 & w36112;
assign w33329 = ~w17779 & ~w3198;
assign w33330 = ~w18047 & ~w2642;
assign w33331 = ~w18860 & ~w2642;
assign w33332 = w5962 & w36113;
assign w33333 = ~w20661 & ~w6764;
assign w33334 = w5962 & w36114;
assign w33335 = ~w20693 & ~w5199;
assign w33336 = w6761 & w36115;
assign w33337 = ~w21282 & ~w7616;
assign w33338 = w6761 & w36116;
assign w33339 = ~w21315 & ~w5965;
assign w33340 = ~w21491 & ~w7616;
assign w33341 = ~w21508 & ~w6764;
assign w33342 = ~w21623 & ~w8529;
assign w33343 = ~w21714 & ~w6764;
assign w33344 = w9534 & w36117;
assign w33345 = w6761 & w36118;
assign w33346 = w11620 & w36119;
assign w33347 = ~w22240 & ~w8529;
assign w33348 = ~w22416 & ~w7616;
assign w33349 = w11620 & w36120;
assign w33350 = w10562 & w36121;
assign w33351 = w7613 & w36122;
assign w33352 = w9534 & w36123;
assign w33353 = ~w22830 & ~w7616;
assign w33354 = w9534 & w36124;
assign w33355 = ~w22902 & ~w8529;
assign w33356 = w10562 & w36125;
assign w33357 = w9534 & w36126;
assign w33358 = ~w23053 & ~w8529;
assign w33359 = w23848 & ~w23951;
assign w33360 = ~w24237 & ~w11623;
assign w33361 = w11620 & w36127;
assign w33362 = (w25296 & w25297) | (w25296 & w23910) | (w25297 & w23910);
assign w33363 = (w25296 & w25297) | (w25296 & w26980) | (w25297 & w26980);
assign w33364 = (w25296 & w25297) | (w25296 & w33020) | (w25297 & w33020);
assign w33365 = (w26872 & w33362) | (w26872 & w36128) | (w33362 & w36128);
assign w33366 = ~w24873 & w33234;
assign w33367 = ~w24873 & w33233;
assign w33368 = ~w24907 & w33238;
assign w33369 = ~w24907 & w33237;
assign w33370 = w24935 & w33242;
assign w33371 = w24935 & w33241;
assign w33372 = b_4 & a_14;
assign w33373 = b_4 & a_17;
assign w33374 = b_4 & a_20;
assign w33375 = b_4 & a_23;
assign w33376 = b_4 & a_50;
assign w33377 = b_4 & a_53;
assign w33378 = (a_14 & ~w657) | (a_14 & w36129) | (~w657 & w36129);
assign w33379 = (a_17 & ~w986) | (a_17 & w36130) | (~w986 & w36130);
assign w33380 = (a_20 & ~w1295) | (a_20 & w36131) | (~w1295 & w36131);
assign w33381 = (a_23 & ~w1694) | (a_23 & w36132) | (~w1694 & w36132);
assign w33382 = w2158 & w36133;
assign w33383 = w6761 & w36134;
assign w33384 = (a_50 & ~w7613) | (a_50 & w36135) | (~w7613 & w36135);
assign w33385 = w7613 & w36136;
assign w33386 = (a_53 & ~w8526) | (a_53 & w36137) | (~w8526 & w36137);
assign w33387 = w8526 & w36138;
assign w33388 = ~w10664 & ~w3806;
assign w33389 = w3195 & w36139;
assign w33390 = ~w10699 & ~w2642;
assign w33391 = w2158 & w36140;
assign w33392 = w418 & w36141;
assign w33393 = w2158 & w36142;
assign w33394 = w5962 & w36143;
assign w33395 = ~w10878 & ~w6764;
assign w33396 = ~w11005 & ~w3806;
assign w33397 = w3195 & w36144;
assign w33398 = ~w11039 & ~w2642;
assign w33399 = ~w10472 & ~w10448;
assign w33400 = w418 & w36145;
assign w33401 = w5962 & w36146;
assign w33402 = ~w11391 & ~w4502;
assign w33403 = w3803 & w36147;
assign w33404 = ~w11427 & ~w3198;
assign w33405 = w2158 & w36148;
assign w33406 = ~w11550 & ~w421;
assign w33407 = w657 & w36149;
assign w33408 = ~w11721 & ~w4502;
assign w33409 = w3803 & w36150;
assign w33410 = ~w11774 & ~w2642;
assign w33411 = w1295 & w36151;
assign w33412 = w986 & w36152;
assign w33413 = w657 & w36153;
assign w33414 = ~w12071 & ~w4502;
assign w33415 = w3803 & w36154;
assign w33416 = w3195 & w36155;
assign w33417 = ~w12124 & ~w2642;
assign w33418 = w2158 & w36156;
assign w33419 = ~w12289 & ~w660;
assign w33420 = ~w12488 & ~w4502;
assign w33421 = w3803 & w36157;
assign w33422 = ~w12589 & ~w421;
assign w33423 = ~w12692 & ~w660;
assign w33424 = ~w12880 & ~w4502;
assign w33425 = w3803 & w36158;
assign w33426 = ~w12958 & ~w1697;
assign w33427 = ~w13224 & ~w3806;
assign w33428 = ~w13259 & ~w2642;
assign w33429 = w2158 & w36159;
assign w33430 = w1694 & w36160;
assign w33431 = w13364 & w13367;
assign w33432 = ~w13364 & ~w13367;
assign w33433 = ~w13433 & ~w989;
assign w33434 = w13351 & w13364;
assign w33435 = ~w13763 & ~w660;
assign w33436 = w1295 & w36161;
assign w33437 = ~w14026 & ~w1697;
assign w33438 = w1295 & w36162;
assign w33439 = w1694 & w36163;
assign w33440 = ~w14519 & ~w989;
assign w33441 = ~w14548 & ~w2161;
assign w33442 = ~w14889 & ~w1298;
assign w33443 = w986 & w36164;
assign w33444 = ~w15197 & ~w1697;
assign w33445 = w2158 & w36165;
assign w33446 = w2639 & w36166;
assign w33447 = w1295 & w36167;
assign w33448 = w16105 & ~w30592;
assign w33449 = w16105 & ~w30591;
assign w33450 = (w15794 & w36168) | (w15794 & w36169) | (w36168 & w36169);
assign w33451 = ~w16536 & ~w1697;
assign w33452 = ~w16839 & ~w2642;
assign w33453 = ~w17149 & ~w1697;
assign w33454 = w3195 & w36170;
assign w33455 = ~w17687 & w17676;
assign w33456 = w3195 & w36171;
assign w33457 = ~w17970 & w17775;
assign w33458 = ~w17970 & w31043;
assign w33459 = ~w18034 & ~w2161;
assign w33460 = w2639 & w36172;
assign w33461 = ~w18062 & ~w3198;
assign w33462 = ~w18595 & ~w3198;
assign w33463 = w2639 & w36173;
assign w33464 = ~w18875 & ~w3198;
assign w33465 = ~w19627 & ~w3198;
assign w33466 = ~w20012 & ~w5199;
assign w33467 = ~w20217 & ~w5965;
assign w33468 = ~w20235 & ~w5199;
assign w33469 = ~w20373 & ~w6764;
assign w33470 = w20215 & w20489;
assign w33471 = ~w20495 & ~w5199;
assign w33472 = ~w20644 & ~w7616;
assign w33473 = w6761 & w36174;
assign w33474 = w5196 & w36175;
assign w33475 = ~w21025 & ~w7616;
assign w33476 = ~w21133 & ~w5965;
assign w33477 = (w21116 & w36176) | (w21116 & w21142) | (w36176 & w21142);
assign w33478 = ~w20900 & w36177;
assign w33479 = ~w21265 & ~w8529;
assign w33480 = w7613 & w36178;
assign w33481 = w5962 & w36179;
assign w33482 = ~w21414 & ~w8529;
assign w33483 = ~w21454 & ~w11623;
assign w33484 = w7613 & w36180;
assign w33485 = w6761 & w36181;
assign w33486 = ~w21525 & ~w5965;
assign w33487 = ~w21600 & ~w5199;
assign w33488 = ~w21611 & ~w5965;
assign w33489 = w8526 & w36182;
assign w33490 = w6761 & w36183;
assign w33491 = w21723 & ~w21709;
assign w33492 = w21723 & w21710;
assign w33493 = ~w21832 & ~w10565;
assign w33494 = ~w21905 & ~w5965;
assign w33495 = w8526 & w36184;
assign w33496 = w7613 & w36185;
assign w33497 = ~w22608 & ~w6764;
assign w33498 = ~w22727 & ~w10565;
assign w33499 = ~w22760 & ~w8529;
assign w33500 = w7613 & w36186;
assign w33501 = w8526 & w36187;
assign w33502 = ~w22924 & ~w6764;
assign w33503 = w8526 & w36188;
assign w33504 = (~w23081 & w23063) | (~w23081 & w36189) | (w23063 & w36189);
assign w33505 = ~w23318 & ~w11623;
assign w33506 = ~w23336 & ~w10565;
assign w33507 = ~w23835 & ~w10565;
assign w33508 = (w25271 & w25272) | (w25271 & ~w32993) | (w25272 & ~w32993);
assign w33509 = (w25271 & w25272) | (w25271 & ~w32994) | (w25272 & ~w32994);
assign w33510 = ~w23925 & ~w9537;
assign w33511 = w33359 & ~w23950;
assign w33512 = w11620 & w36190;
assign w33513 = w24441 & w26493;
assign w33514 = w24441 & w26492;
assign w33515 = (~w33020 & w36191) | (~w33020 & w36192) | (w36191 & w36192);
assign w33516 = ~w24548 & ~w33365;
assign w33517 = (~w25297 & w36193) | (~w25297 & w36191) | (w36193 & w36191);
assign w33518 = (~w25297 & w36194) | (~w25297 & w36191) | (w36194 & w36191);
assign w33519 = (~w33020 & w36195) | (~w33020 & w36196) | (w36195 & w36196);
assign w33520 = (w25299 & w25300) | (w25299 & ~w33365) | (w25300 & ~w33365);
assign w33521 = (~w25297 & w36197) | (~w25297 & w36195) | (w36197 & w36195);
assign w33522 = (~w25297 & w36198) | (~w25297 & w36195) | (w36198 & w36195);
assign w33523 = (~w33020 & w36199) | (~w33020 & w36200) | (w36199 & w36200);
assign w33524 = (w25304 & w25303) | (w25304 & ~w33365) | (w25303 & ~w33365);
assign w33525 = (~w25297 & w36201) | (~w25297 & w36199) | (w36201 & w36199);
assign w33526 = (~w25297 & w36202) | (~w25297 & w36199) | (w36202 & w36199);
assign w33527 = (~w33020 & w36203) | (~w33020 & w36204) | (w36203 & w36204);
assign w33528 = (w25308 & w25307) | (w25308 & ~w33365) | (w25307 & ~w33365);
assign w33529 = (~w25297 & w36205) | (~w25297 & w36203) | (w36205 & w36203);
assign w33530 = (~w25297 & w36206) | (~w25297 & w36203) | (w36206 & w36203);
assign w33531 = (~w33020 & w36207) | (~w33020 & w36208) | (w36207 & w36208);
assign w33532 = (w25311 & w25312) | (w25311 & ~w33365) | (w25312 & ~w33365);
assign w33533 = (~w25297 & w36209) | (~w25297 & w36207) | (w36209 & w36207);
assign w33534 = (~w25297 & w36210) | (~w25297 & w36207) | (w36210 & w36207);
assign w33535 = w24957 & ~w24932;
assign w33536 = w24935 & w33535;
assign w33537 = ~w24972 & w33141;
assign w33538 = ~w24972 & w33140;
assign w33539 = w24980 & w33144;
assign w33540 = (w24980 & w25333) | (w24980 & w36211) | (w25333 & w36211);
assign w33541 = ~w24980 & ~w33144;
assign w33542 = ~w25333 & w36212;
assign w33543 = b_4 & a_11;
assign w33544 = b_4 & a_32;
assign w33545 = b_4 & a_35;
assign w33546 = b_4 & a_38;
assign w33547 = b_4 & a_41;
assign w33548 = (a_11 & ~w418) | (a_11 & w36213) | (~w418 & w36213);
assign w33549 = w2639 & w36214;
assign w33550 = (a_32 & ~w3195) | (a_32 & w36215) | (~w3195 & w36215);
assign w33551 = (a_35 & ~w3803) | (a_35 & w36216) | (~w3803 & w36216);
assign w33552 = w3803 & w36217;
assign w33553 = (a_38 & ~w4499) | (a_38 & w36218) | (~w4499 & w36218);
assign w33554 = w4499 & w36219;
assign w33555 = (a_41 & ~w5196) | (a_41 & w36220) | (~w5196 & w36220);
assign w33556 = w5196 & w36221;
assign w33557 = ~w7486 & ~w660;
assign w33558 = w418 & w36222;
assign w33559 = ~w7777 & ~w660;
assign w33560 = w418 & w36223;
assign w33561 = ~w7532 & ~w7530;
assign w33562 = w239 & w36224;
assign w33563 = w1295 & w36225;
assign w33564 = ~w8660 & ~w1697;
assign w33565 = ~w8678 & ~w1298;
assign w33566 = w986 & w36226;
assign w33567 = w418 & w36227;
assign w33568 = w239 & w36228;
assign w33569 = ~w8807 & ~w1298;
assign w33570 = ~w8818 & ~w1697;
assign w33571 = ~w26604 & w8927;
assign w33572 = w26604 & ~w8927;
assign w33573 = w239 & w36229;
assign w33574 = w1694 & w36230;
assign w33575 = ~w9347 & ~w1298;
assign w33576 = ~w9405 & ~w242;
assign w33577 = ~w9631 & ~w2642;
assign w33578 = ~w9649 & ~w2161;
assign w33579 = ~w9667 & ~w1697;
assign w33580 = w1295 & w36231;
assign w33581 = w1694 & w36232;
assign w33582 = w2158 & w36233;
assign w33583 = ~w26632 & w9917;
assign w33584 = w26632 & ~w9917;
assign w33585 = ~w11836 & ~w11495;
assign w33586 = ~w11836 & w11096;
assign w33587 = ~w13460 & ~w1697;
assign w33588 = w1694 & w36234;
assign w33589 = w13428 & w13726;
assign w33590 = ~w15436 & w15220;
assign w33591 = ~w15907 & ~w3198;
assign w33592 = ~w16565 & ~w2642;
assign w33593 = ~w17659 & ~w3806;
assign w33594 = ~w18463 & ~w4502;
assign w33595 = ~w18481 & ~w3806;
assign w33596 = ~w19776 & ~w5199;
assign w33597 = ~w19979 & ~w6764;
assign w33598 = ~w19996 & ~w5965;
assign w33599 = w5196 & w36235;
assign w33600 = ~w20107 & ~w6764;
assign w33601 = w5962 & w36236;
assign w33602 = ~w20834 & ~w11623;
assign w33603 = ~w20890 & ~w6764;
assign w33604 = w20888 & w21127;
assign w33605 = ~w21203 & ~w9537;
assign w33606 = w8526 & w36237;
assign w33607 = w8526 & w36238;
assign w33608 = ~w21425 & ~w9537;
assign w33609 = ~w21898 & ~w26438;
assign w33610 = (w26021 & w36239) | (w26021 & w36240) | (w36239 & w36240);
assign w33611 = ~w22046 & ~w8529;
assign w33612 = (w25245 & w25244) | (w25245 & w32976) | (w25244 & w32976);
assign w33613 = (w25245 & w25244) | (w25245 & w32977) | (w25244 & w32977);
assign w33614 = w25244 & w25245;
assign w33615 = (w25245 & w25244) | (w25245 & ~w21777) | (w25244 & ~w21777);
assign w33616 = ~w23199 & ~w10565;
assign w33617 = w11620 & w36241;
assign w33618 = w10562 & w36242;
assign w33619 = ~w23909 & ~w33508;
assign w33620 = (w32994 & w36243) | (w32994 & w36244) | (w36243 & w36244);
assign w33621 = (w25274 & w25275) | (w25274 & ~w33508) | (w25275 & ~w33508);
assign w33622 = (w32994 & w36245) | (w32994 & w36246) | (w36245 & w36246);
assign w33623 = (w25279 & w25278) | (w25279 & ~w33508) | (w25278 & ~w33508);
assign w33624 = (w32994 & w36247) | (w32994 & w36248) | (w36247 & w36248);
assign w33625 = (w25282 & w25283) | (w25282 & ~w33508) | (w25283 & ~w33508);
assign w33626 = (w32994 & w36249) | (w32994 & w36250) | (w36249 & w36250);
assign w33627 = (w25286 & w25287) | (w25286 & ~w33508) | (w25287 & ~w33508);
assign w33628 = (w32994 & w36251) | (w32994 & w36252) | (w36251 & w36252);
assign w33629 = (w25290 & w25291) | (w25290 & ~w33508) | (w25291 & ~w33508);
assign w33630 = (w32994 & w36253) | (w32994 & w36254) | (w36253 & w36254);
assign w33631 = (w25294 & w25295) | (w25294 & ~w33508) | (w25295 & ~w33508);
assign w33632 = (w32994 & w36255) | (w32994 & w36256) | (w36255 & w36256);
assign w33633 = (w33020 & w36257) | (w33020 & w36258) | (w36257 & w36258);
assign w33634 = (w25325 & w25326) | (w25325 & w33365) | (w25326 & w33365);
assign w33635 = (w25297 & w36259) | (w25297 & w36257) | (w36259 & w36257);
assign w33636 = (w25297 & w36260) | (w25297 & w36257) | (w36260 & w36257);
assign w33637 = w239 & w36261;
assign w33638 = w657 & w36262;
assign w33639 = w986 & w36263;
assign w33640 = w1295 & w36264;
assign w33641 = w5962 & w36265;
assign w33642 = ~w7125 & ~w7391;
assign w33643 = w9534 & w36266;
assign w33644 = (~w11529 & w36267) | (~w11529 & w36268) | (w36267 & w36268);
assign w33645 = (w11529 & w36269) | (w11529 & w36270) | (w36269 & w36270);
assign w33646 = (w13389 & w13008) | (w13389 & w36271) | (w13008 & w36271);
assign w33647 = ~w13008 & w36272;
assign w33648 = (w25483 & w36273) | (w25483 & w33650) | (w36273 & w33650);
assign w33649 = (~w26973 & w36274) | (~w26973 & w36273) | (w36274 & w36273);
assign w33650 = (w25207 & w25208) | (w25207 & ~w26973) | (w25208 & ~w26973);
assign w33651 = (~w26866 & w36275) | (~w26866 & w36273) | (w36275 & w36273);
assign w33652 = (w25483 & w36276) | (w25483 & w33653) | (w36276 & w33653);
assign w33653 = (w25219 & w25220) | (w25219 & ~w26973) | (w25220 & ~w26973);
assign w33654 = (w25219 & w25220) | (w25219 & ~w32962) | (w25220 & ~w32962);
assign w33655 = (w25483 & w36277) | (w25483 & w33657) | (w36277 & w33657);
assign w33656 = (w25223 & w25224) | (w25223 & ~w32963) | (w25224 & ~w32963);
assign w33657 = (w25223 & w25224) | (w25223 & ~w26973) | (w25224 & ~w26973);
assign w33658 = (w25223 & w25224) | (w25223 & ~w32962) | (w25224 & ~w32962);
assign w33659 = (w25244 & w36278) | (w25244 & w36279) | (w36278 & w36279);
assign w33660 = (w25244 & w36280) | (w25244 & w36279) | (w36280 & w36279);
assign w33661 = (w32977 & w36279) | (w32977 & w36281) | (w36279 & w36281);
assign w33662 = (w25244 & w36282) | (w25244 & w36283) | (w36282 & w36283);
assign w33663 = (w25244 & w36284) | (w25244 & w36283) | (w36284 & w36283);
assign w33664 = (w32977 & w36283) | (w32977 & w36285) | (w36283 & w36285);
assign w33665 = (w25244 & w36286) | (w25244 & w36287) | (w36286 & w36287);
assign w33666 = (w25244 & w36288) | (w25244 & w36287) | (w36288 & w36287);
assign w33667 = (w32977 & w36287) | (w32977 & w36289) | (w36287 & w36289);
assign w33668 = (w25244 & w36290) | (w25244 & w36291) | (w36290 & w36291);
assign w33669 = (w25244 & w36292) | (w25244 & w36291) | (w36292 & w36291);
assign w33670 = (w32977 & w36291) | (w32977 & w36293) | (w36291 & w36293);
assign w33671 = (w25244 & w36294) | (w25244 & w36295) | (w36294 & w36295);
assign w33672 = (w25244 & w36296) | (w25244 & w36295) | (w36296 & w36295);
assign w33673 = (w32977 & w36295) | (w32977 & w36297) | (w36295 & w36297);
assign w33674 = (w25244 & w36298) | (w25244 & w36299) | (w36298 & w36299);
assign w33675 = (w25244 & w36300) | (w25244 & w36299) | (w36300 & w36299);
assign w33676 = (w32977 & w36299) | (w32977 & w36301) | (w36299 & w36301);
assign w33677 = (w25244 & w36302) | (w25244 & w36303) | (w36302 & w36303);
assign w33678 = (w25244 & w36304) | (w25244 & w36303) | (w36304 & w36303);
assign w33679 = (w32977 & w36303) | (w32977 & w36305) | (w36303 & w36305);
assign w33680 = (~w25244 & w36306) | (~w25244 & w36307) | (w36306 & w36307);
assign w33681 = (~w25244 & w36308) | (~w25244 & w36307) | (w36308 & w36307);
assign w33682 = (w26076 & w26075) | (w26076 & ~w33612) | (w26075 & ~w33612);
assign w33683 = (~w32977 & w36307) | (~w32977 & w36309) | (w36307 & w36309);
assign w33684 = ~w24619 & w33518;
assign w33685 = ~w24619 & w33517;
assign w33686 = w24682 & w33522;
assign w33687 = w24682 & w33521;
assign w33688 = ~w24739 & w33526;
assign w33689 = ~w24739 & w33525;
assign w33690 = ~w24791 & w33530;
assign w33691 = ~w24791 & w33529;
assign w33692 = ~w24832 & w33534;
assign w33693 = ~w24832 & w33533;
assign w33694 = w418 & w36310;
assign w33695 = ~w3653 & ~w3466;
assign w33696 = ~w3653 & ~w3467;
assign w33697 = w3195 & w36311;
assign w33698 = (~w3827 & ~w4076) | (~w3827 & w36312) | (~w4076 & w36312);
assign w33699 = w10562 & w36313;
assign w33700 = (~w19828 & w25191) | (~w19828 & w32955) | (w25191 & w32955);
assign w33701 = (w26970 & ~w19828) | (w26970 & w36314) | (~w19828 & w36314);
assign w33702 = (w25194 & w25195) | (w25194 & w32955) | (w25195 & w32955);
assign w33703 = (w26970 & w36315) | (w26970 & w36316) | (w36315 & w36316);
assign w33704 = (w25204 & w25205) | (w25204 & ~w32955) | (w25205 & ~w32955);
assign w33705 = (w25204 & w25205) | (w25204 & ~w32954) | (w25205 & ~w32954);
assign w33706 = ~w21182 & w33649;
assign w33707 = ~w21182 & w33648;
assign w33708 = (~w32963 & w36317) | (~w32963 & w36318) | (w36317 & w36318);
assign w33709 = ~w21779 & w33652;
assign w33710 = (~w32963 & w36319) | (~w32963 & w36320) | (w36319 & w36320);
assign w33711 = (~w21960 & w25225) | (~w21960 & w33655) | (w25225 & w33655);
assign w33712 = (~w32963 & w36321) | (~w32963 & w36322) | (w36321 & w36322);
assign w33713 = (w25229 & w25228) | (w25229 & w33655) | (w25228 & w33655);
assign w33714 = (~w32963 & w36323) | (~w32963 & w36324) | (w36323 & w36324);
assign w33715 = (w25233 & w25232) | (w25233 & w33655) | (w25232 & w33655);
assign w33716 = (~w32963 & w36325) | (~w32963 & w36326) | (w36325 & w36326);
assign w33717 = (w25237 & w25236) | (w25237 & w33655) | (w25236 & w33655);
assign w33718 = (~w32963 & w36327) | (~w32963 & w36328) | (w36327 & w36328);
assign w33719 = (w25241 & w25240) | (w25241 & w33655) | (w25240 & w33655);
assign w33720 = (w32963 & w36329) | (w32963 & w36330) | (w36329 & w36330);
assign w33721 = (w26484 & w26485) | (w26484 & ~w33655) | (w26485 & ~w33655);
assign w33722 = ~w33508 & w36331;
assign w33723 = ~w24022 & w33620;
assign w33724 = (~w33508 & w36332) | (~w33508 & w36333) | (w36332 & w36333);
assign w33725 = ~w24125 & w33622;
assign w33726 = (~w33508 & w36334) | (~w33508 & w36335) | (w36334 & w36335);
assign w33727 = ~w24222 & w33624;
assign w33728 = (~w33508 & w36336) | (~w33508 & w36337) | (w36336 & w36337);
assign w33729 = ~w24315 & w33626;
assign w33730 = (~w33508 & w36338) | (~w33508 & w36339) | (w36338 & w36339);
assign w33731 = ~w24400 & w33628;
assign w33732 = (~w33508 & w36340) | (~w33508 & w36341) | (w36340 & w36341);
assign w33733 = ~w24476 & w33630;
assign w33734 = (~w33508 & w36342) | (~w33508 & w36343) | (w36342 & w36343);
assign w33735 = ~w24549 & w33632;
assign w33736 = w24480 & w24529;
assign w33737 = ~w24589 & ~w11623;
assign w33738 = w11623 & ~w29581;
assign w33739 = w11623 & ~w29580;
assign w33740 = ~w21778 & ~w21777;
assign w33741 = w23794 & w23910;
assign w33742 = w36344 & ~w10433;
assign w33743 = b_4 & a_44;
assign w33744 = b_4 & a_5;
assign w33745 = b_4 & a_8;
assign w33746 = (a_5 & ~w99) | (a_5 & w36345) | (~w99 & w36345);
assign w33747 = w99 & w36346;
assign w33748 = (a_8 & ~w239) | (a_8 & w36347) | (~w239 & w36347);
assign w33749 = w2717 & w36348;
assign w33750 = ~w4300 & ~w4094;
assign w33751 = ~w4300 & ~w4095;
assign w33752 = (a_44 & ~w5962) | (a_44 & w36349) | (~w5962 & w36349);
assign w33753 = (w25189 & w25190) | (w25189 & w32941) | (w25190 & w32941);
assign w33754 = (w25189 & w25190) | (w25189 & w32942) | (w25190 & w32942);
assign w33755 = (w25189 & w25190) | (w25189 & ~w18545) | (w25190 & ~w18545);
assign w33756 = ~w20073 & ~w19828;
assign w33757 = w19831 & w33756;
assign w33758 = (w20074 & w36350) | (w20074 & w36351) | (w36350 & w36351);
assign w33759 = (w25191 & w36350) | (w25191 & w36352) | (w36350 & w36352);
assign w33760 = (~w25196 & w36353) | (~w25196 & w36354) | (w36353 & w36354);
assign w33761 = (w25195 & w36355) | (w25195 & w36356) | (w36355 & w36356);
assign w33762 = (w32954 & w36357) | (w32954 & w36358) | (w36357 & w36358);
assign w33763 = (w32955 & w36357) | (w32955 & w36358) | (w36357 & w36358);
assign w33764 = (~w25196 & w36359) | (~w25196 & w36360) | (w36359 & w36360);
assign w33765 = (w25195 & w36361) | (w25195 & w36362) | (w36361 & w36362);
assign w33766 = (w32954 & w36363) | (w32954 & w36364) | (w36363 & w36364);
assign w33767 = (w32955 & w36363) | (w32955 & w36364) | (w36363 & w36364);
assign w33768 = (~w25196 & w36365) | (~w25196 & w36366) | (w36365 & w36366);
assign w33769 = (w25195 & w36367) | (w25195 & w36368) | (w36367 & w36368);
assign w33770 = (w32954 & w36369) | (w32954 & w36370) | (w36369 & w36370);
assign w33771 = (w32955 & w36369) | (w32955 & w36370) | (w36369 & w36370);
assign w33772 = (~w25196 & w36371) | (~w25196 & w36372) | (w36371 & w36372);
assign w33773 = (w25195 & w36373) | (w25195 & w36374) | (w36373 & w36374);
assign w33774 = (w32954 & w36375) | (w32954 & w36376) | (w36375 & w36376);
assign w33775 = (w32955 & w36375) | (w32955 & w36376) | (w36375 & w36376);
assign w33776 = (w33612 & w36377) | (w33612 & w36378) | (w36377 & w36378);
assign w33777 = ~w23127 & w33661;
assign w33778 = (w33612 & w36379) | (w33612 & w36380) | (w36379 & w36380);
assign w33779 = ~w23272 & w33664;
assign w33780 = (w33612 & w36381) | (w33612 & w36382) | (w36381 & w36382);
assign w33781 = ~w23413 & w33667;
assign w33782 = (w33612 & w36383) | (w33612 & w36384) | (w36383 & w36384);
assign w33783 = ~w23544 & w33670;
assign w33784 = (w33612 & w36385) | (w33612 & w36386) | (w36385 & w36386);
assign w33785 = ~w23676 & w33673;
assign w33786 = (w33612 & w36387) | (w33612 & w36388) | (w36387 & w36388);
assign w33787 = ~w23798 & w33676;
assign w33788 = (w33612 & w36389) | (w33612 & w36390) | (w36389 & w36390);
assign w33789 = ~w23910 & w33679;
assign w33790 = (~w33612 & w36391) | (~w33612 & w36392) | (w36391 & w36392);
assign w33791 = (w24619 & w25298) | (w24619 & w33683) | (w25298 & w33683);
assign w33792 = (w24619 & w25298) | (w24619 & w33681) | (w25298 & w33681);
assign w33793 = (w24619 & w25298) | (w24619 & w33680) | (w25298 & w33680);
assign w33794 = (~w33612 & w36393) | (~w33612 & w36394) | (w36393 & w36394);
assign w33795 = (w25301 & w25302) | (w25301 & w33683) | (w25302 & w33683);
assign w33796 = (w25301 & w25302) | (w25301 & w33681) | (w25302 & w33681);
assign w33797 = (w25301 & w25302) | (w25301 & w33680) | (w25302 & w33680);
assign w33798 = (~w33612 & w36395) | (~w33612 & w36396) | (w36395 & w36396);
assign w33799 = (w25305 & w25306) | (w25305 & w33683) | (w25306 & w33683);
assign w33800 = (w25305 & w25306) | (w25305 & w33681) | (w25306 & w33681);
assign w33801 = (w25305 & w25306) | (w25305 & w33680) | (w25306 & w33680);
assign w33802 = (~w33612 & w36397) | (~w33612 & w36398) | (w36397 & w36398);
assign w33803 = (w25309 & w25310) | (w25309 & w33683) | (w25310 & w33683);
assign w33804 = (w25309 & w25310) | (w25309 & w33681) | (w25310 & w33681);
assign w33805 = (w25309 & w25310) | (w25309 & w33680) | (w25310 & w33680);
assign w33806 = (~w33612 & w36399) | (~w33612 & w36400) | (w36399 & w36400);
assign w33807 = (w25313 & w25314) | (w25313 & w33683) | (w25314 & w33683);
assign w33808 = (w25313 & w25314) | (w25313 & w33681) | (w25314 & w33681);
assign w33809 = (w25313 & w25314) | (w25313 & w33680) | (w25314 & w33680);
assign w33810 = (~w33612 & w36401) | (~w33612 & w36402) | (w36401 & w36402);
assign w33811 = (w25318 & w25317) | (w25318 & w33683) | (w25317 & w33683);
assign w33812 = (w25318 & w25317) | (w25318 & w33681) | (w25317 & w33681);
assign w33813 = (w25318 & w25317) | (w25318 & w33680) | (w25317 & w33680);
assign w33814 = (~w33612 & w36403) | (~w33612 & w36404) | (w36403 & w36404);
assign w33815 = (w25322 & w25321) | (w25322 & w33683) | (w25321 & w33683);
assign w33816 = (w25322 & w25321) | (w25322 & w33681) | (w25321 & w33681);
assign w33817 = (w25322 & w25321) | (w25322 & w33680) | (w25321 & w33680);
assign w33818 = (~w33612 & w36405) | (~w33612 & w36406) | (w36405 & w36406);
assign w33819 = (w25716 & w25715) | (w25716 & w33683) | (w25715 & w33683);
assign w33820 = (w25716 & w25715) | (w25716 & w33681) | (w25715 & w33681);
assign w33821 = (w25716 & w25715) | (w25716 & w33680) | (w25715 & w33680);
assign w33822 = (~w33612 & w36407) | (~w33612 & w36408) | (w36407 & w36408);
assign w33823 = (w25718 & w25717) | (w25718 & w33683) | (w25717 & w33683);
assign w33824 = (w25718 & w25717) | (w25718 & w33681) | (w25717 & w33681);
assign w33825 = (w25718 & w25717) | (w25718 & w33680) | (w25717 & w33680);
assign w33826 = w3488 & w3685;
assign w33827 = ~w3069 & ~w2893;
assign w33828 = ~w3069 & w2897;
assign w33829 = w7039 & ~w7152;
assign w33830 = (w7302 & w36409) | (w7302 & w36410) | (w36409 & w36410);
assign w33831 = ~w7812 & w36411;
assign w33832 = w7825 & ~w26579;
assign w33833 = (~w5776 & ~w6046) | (~w5776 & w36412) | (~w6046 & w36412);
assign w33834 = ~w5770 & ~w6039;
assign w33835 = ~w6838 & ~w6560;
assign w33836 = ~w6838 & w6456;
assign w33837 = w11620 & w36413;
assign w33838 = (w10110 & w10094) | (w10110 & w36414) | (w10094 & w36414);
assign w33839 = ~w10094 & w36415;
assign w33840 = b_4 & a_56;
assign w33841 = ~w11137 & w36416;
assign w33842 = ~w9206 & ~w9587;
assign w33843 = (w4092 & ~w3826) | (w4092 & w36417) | (~w3826 & w36417);
assign w33844 = w3826 & w36418;
assign w33845 = (w6293 & w6277) | (w6293 & w36419) | (w6277 & w36419);
assign w33846 = ~w6277 & w36420;
assign w33847 = (w7122 & w7106) | (w7122 & w36421) | (w7106 & w36421);
assign w33848 = ~w7106 & w36422;
assign w33849 = ~w7648 & ~w7927;
assign w33850 = (w5506 & w5490) | (w5506 & w36423) | (w5490 & w36423);
assign w33851 = ~w5490 & w36424;
assign w33852 = (w7988 & w7972) | (w7988 & w36425) | (w7972 & w36425);
assign w33853 = ~w7972 & w36426;
assign w33854 = (w11244 & w11114) | (w11244 & w36427) | (w11114 & w36427);
assign w33855 = w8 & w36428;
assign w33856 = ~w4356 & ~w4141;
assign w33857 = ~w4356 & w3920;
assign w33858 = ~w7414 & ~w7136;
assign w33859 = ~w7414 & w7039;
assign w33860 = ~w7991 & ~w7927;
assign w33861 = (a_56 & ~w9534) | (a_56 & w36429) | (~w9534 & w36429);
assign w33862 = ~w12831 & ~w12829;
assign w33863 = ~w12781 & ~w12780;
assign w33864 = b_4 & a_47;
assign w33865 = (w7725 & ~w7439) | (w7725 & w36430) | (~w7439 & w36430);
assign w33866 = ~w9850 & ~w9954;
assign w33867 = w27844 & a_2;
assign w33868 = ~w27387 & a_2;
assign w33869 = ~w3512 & ~w3510;
assign w33870 = (a_47 & ~w6761) | (a_47 & w36431) | (~w6761 & w36431);
assign w33871 = w26833 & ~w11678;
assign w33872 = ~w26833 & ~w11678;
assign w33873 = w1694 & w36432;
assign w33874 = ~w14442 & w36433;
assign w33875 = ~w6367 & ~w6365;
assign w33876 = ~w6592 & ~w6590;
assign w33877 = w6706 & w6897;
assign w33878 = ~w6706 & ~w6897;
assign w33879 = ~w6585 & ~w6874;
assign w33880 = ~w12619 & ~w102;
assign w33881 = ~w13012 & ~w102;
assign w33882 = ~w13318 & ~w989;
assign w33883 = w986 & w36434;
assign w33884 = ~w13446 & ~w1298;
assign w33885 = ~w13790 & ~w2161;
assign w33886 = ~w14209 & ~w2642;
assign w33887 = ~w14533 & ~w1697;
assign w33888 = w14440 & ~w14204;
assign w33889 = w14440 & w14205;
assign w33890 = w2158 & w36435;
assign w33891 = ~w14785 & ~w1298;
assign w33892 = ~w14875 & ~w989;
assign w33893 = w1694 & w36436;
assign w33894 = w660 & ~w29581;
assign w33895 = w660 & ~w29580;
assign w33896 = w15577 & w15804;
assign w33897 = ~w16121 & ~w16464;
assign w33898 = w2639 & w36437;
assign w33899 = ~w16766 & ~w3198;
assign w33900 = w2639 & w36438;
assign w33901 = w17036 & w17048;
assign w33902 = ~w17477 & ~w2642;
assign w33903 = w3803 & w36439;
assign w33904 = w31042 & ~w17969;
assign w33905 = w3195 & w36440;
assign w33906 = ~w18238 & ~w3806;
assign w33907 = w4499 & w36441;
assign w33908 = w3803 & w36442;
assign w33909 = ~w18754 & ~w4502;
assign w33910 = ~w19030 & ~w4502;
assign w33911 = ~w19271 & ~w5199;
assign w33912 = ~w19289 & ~w4502;
assign w33913 = ~w19517 & ~w5199;
assign w33914 = w5196 & w36443;
assign w33915 = ~w19961 & ~w7616;
assign w33916 = w6761 & w36444;
assign w33917 = w5962 & w36445;
assign w33918 = w6761 & w36446;
assign w33919 = ~w20118 & ~w7616;
assign w33920 = w5196 & w36447;
assign w33921 = ~w20795 & ~w7616;
assign w33922 = w6761 & w36448;
assign w33923 = ~w20907 & ~w5965;
assign w33924 = ~w21352 & w36449;
assign w33925 = w21504 & w21517;
assign w33926 = ~w21634 & ~w9537;
assign w33927 = w21794 & w21923;
assign w33928 = ~w21794 & ~w21923;
assign w33929 = ~w21987 & ~w9537;
assign w33930 = w8526 & w36450;
assign w33931 = ~w22063 & ~w7616;
assign w33932 = ~w22183 & ~w9537;
assign w33933 = w10562 & w36451;
assign w33934 = w10562 & w36452;
assign w33935 = ~w23299 & ~w9537;
assign w33936 = w23317 & w27688;
assign w33937 = w23317 & w27687;
assign w33938 = ~w23463 & ~w10565;
assign w33939 = ~w23593 & ~w10565;
assign w33940 = w36453 & ~w23730;
assign w33941 = w23732 & ~w26727;
assign w33942 = ~w23739 & ~w11623;
assign w33943 = ~w23753 & ~w10565;
assign w33944 = w11620 & w36454;
assign w33945 = ~w24253 & w27705;
assign w33946 = ~w24253 & w27704;
assign w33947 = ~w24331 & ~w10565;
assign w33948 = ~w24341 & ~w11623;
assign w33949 = w24437 & ~w24486;
assign w33950 = w11620 & w36455;
assign w33951 = w11620 & w36456;
assign w33952 = ~w12245 & w12278;
assign w33953 = ~w6082 & w36457;
assign w33954 = (~w6098 & w6082) | (~w6098 & w36458) | (w6082 & w36458);
assign w33955 = (~w27522 & w36459) | (~w27522 & w36460) | (w36459 & w36460);
assign w33956 = ~w1770 & ~w1768;
assign w33957 = ~w1915 & ~w1768;
assign w33958 = ~w1915 & w27732;
assign w33959 = ~w6107 & ~w6105;
assign w33960 = ~w6922 & ~w6630;
assign w33961 = ~w6922 & w6422;
assign w33962 = (~w7823 & ~w8116) | (~w7823 & w36461) | (~w8116 & w36461);
assign w33963 = ~w9061 & ~w8742;
assign w33964 = ~w9061 & w8478;
assign w33965 = (~w25148 & w36462) | (~w25148 & w36463) | (w36462 & w36463);
assign w33966 = (~w25149 & w36462) | (~w25149 & w36463) | (w36462 & w36463);
assign w33967 = (w13327 & ~w12973) | (w13327 & w36464) | (~w12973 & w36464);
assign w33968 = w13327 & w12977;
assign w33969 = w12973 & w36465;
assign w33970 = ~w13327 & ~w12977;
assign w33971 = w14942 & ~w15436;
assign w33972 = ~w12955 & w12967;
assign w33973 = w12955 & ~w12967;
assign w33974 = ~w13059 & ~w13302;
assign w33975 = w13058 & w13442;
assign w33976 = ~w13058 & ~w13442;
assign w33977 = (w25153 & w36466) | (w25153 & w36467) | (w36466 & w36467);
assign w33978 = w12712 & ~w13718;
assign w33979 = ~w707 & ~w731;
assign w33980 = ~w732 & ~w731;
assign w33981 = w13059 & ~w13302;
assign w33982 = w13486 & w36468;
assign w33983 = ~w13455 & ~w14057;
assign w33984 = ~w14097 & ~w14136;
assign w33985 = ~w14087 & ~w14136;
assign w33986 = ~w14079 & ~w14468;
assign w33987 = (~w14468 & w14067) | (~w14468 & w36469) | (w14067 & w36469);
assign w33988 = w1694 & w36470;
assign w33989 = w1295 & w36471;
assign w33990 = w14542 & w14780;
assign w33991 = w15192 & w15461;
assign w33992 = w15436 & w15220;
assign w33993 = w15436 & ~w30368;
assign w33994 = ~w15809 & ~w1697;
assign w33995 = ~w15865 & ~w1298;
assign w33996 = (w13046 & ~w12987) | (w13046 & w36472) | (~w12987 & w36472);
assign w33997 = w7881 & w8406;
assign w33998 = (w8687 & ~w8389) | (w8687 & w36473) | (~w8389 & w36473);
assign w33999 = (w8723 & ~w8412) | (w8723 & w36474) | (~w8412 & w36474);
assign w34000 = w8705 & w9023;
assign w34001 = ~w25092 & w9745;
assign w34002 = w25092 & ~w9745;
assign w34003 = ~w12616 & ~w12628;
assign w34004 = (w12677 & ~w12606) | (w12677 & w36475) | (~w12606 & w36475);
assign w34005 = w10087 & w9745;
assign w34006 = w10087 & ~w27829;
assign w34007 = ~w0 & a_2;
assign w34008 = ~w73 & ~w12;
assign w34009 = w27387 & a_2;
assign w34010 = (a_2 & w27387) | (a_2 & w12) | (w27387 & w12);
assign w34011 = ~w119 & ~w12;
assign w34012 = ~w180 & ~w12;
assign w34013 = ~w203 & ~w12;
assign w34014 = ~w210 & ~w209;
assign w34015 = w8 & w36476;
assign w34016 = ~w322 & ~w102;
assign w34017 = ~w361 & ~w12;
assign w34018 = ~w386 & ~w102;
assign w34019 = ~w444 & ~w12;
assign w34020 = ~w438 & ~w436;
assign w34021 = w99 & w36477;
assign w34022 = ~w520 & ~w12;
assign w34023 = ~w549 & ~w526;
assign w34024 = ~w549 & w27200;
assign w34025 = ~w542 & ~w12;
assign w34026 = ~w558 & ~w242;
assign w34027 = ~w597 & ~w102;
assign w34028 = ~w625 & ~w242;
assign w34029 = ~w683 & ~w102;
assign w34030 = ~w700 & ~w12;
assign w34031 = ~w725 & ~w12;
assign w34032 = ~w741 & ~w102;
assign w34033 = ~w677 & ~w675;
assign w34034 = w239 & w36478;
assign w34035 = ~w817 & ~w12;
assign w34036 = ~w834 & ~w102;
assign w34037 = ~w845 & ~w242;
assign w34038 = ~w855 & ~w421;
assign w34039 = ~w824 & ~w823;
assign w34040 = ~w916 & ~w12;
assign w34041 = ~w933 & ~w102;
assign w34042 = ~w943 & ~w242;
assign w34043 = ~w954 & ~w421;
assign w34044 = ~w1028 & ~w12;
assign w34045 = ~w1045 & ~w102;
assign w34046 = ~w1056 & ~w242;
assign w34047 = w418 & w36479;
assign w34048 = ~w1140 & ~w102;
assign w34049 = ~w1151 & ~w242;
assign w34050 = ~w1162 & ~w660;
assign w34051 = ~w1200 & ~w421;
assign w34052 = ~w922 & ~w1034;
assign w34053 = ~w1035 & ~w1034;
assign w34054 = ~w1228 & ~w12;
assign w34055 = ~w1252 & ~w102;
assign w34056 = ~w1263 & ~w660;
assign w34057 = ~w1319 & ~w421;
assign w34058 = ~w1337 & ~w242;
assign w34059 = ~w1235 & ~w1234;
assign w34060 = w1369 & w1234;
assign w34061 = w1369 & ~w34059;
assign w34062 = ~w1369 & ~w1234;
assign w34063 = ~w1369 & w34059;
assign w34064 = ~w1387 & ~w102;
assign w34065 = ~w1397 & ~w242;
assign w34066 = ~w1408 & ~w421;
assign w34067 = w657 & w36480;
assign w34068 = ~w1493 & ~w12;
assign w34069 = ~w1380 & ~w1378;
assign w34070 = ~w1518 & ~w242;
assign w34071 = ~w1529 & ~w421;
assign w34072 = ~w1540 & ~w989;
assign w34073 = ~w1578 & ~w660;
assign w34074 = ~w1606 & ~w102;
assign w34075 = ~w1368 & ~w1499;
assign w34076 = ~w1624 & ~w12;
assign w34077 = ~w1650 & ~w242;
assign w34078 = ~w1662 & ~w989;
assign w34079 = ~w1718 & ~w660;
assign w34080 = ~w1736 & ~w421;
assign w34081 = ~w1758 & ~w102;
assign w34082 = ~w1631 & ~w1630;
assign w34083 = ~w1776 & ~w12;
assign w34084 = ~w1799 & ~w242;
assign w34085 = ~w1809 & ~w421;
assign w34086 = ~w1820 & ~w660;
assign w34087 = w986 & w36481;
assign w34088 = ~w1905 & ~w102;
assign w34089 = ~w1783 & ~w1782;
assign w34090 = w1930 & w1782;
assign w34091 = w1930 & ~w34089;
assign w34092 = ~w1930 & ~w1782;
assign w34093 = ~w1930 & w34089;
assign w34094 = ~w1923 & ~w12;
assign w34095 = ~w1948 & ~w102;
assign w34096 = ~w1959 & ~w421;
assign w34097 = ~w1970 & ~w660;
assign w34098 = ~w1981 & ~w1298;
assign w34099 = ~w2019 & ~w989;
assign w34100 = ~w2049 & ~w242;
assign w34101 = ~w2073 & ~w12;
assign w34102 = ~w1929 & ~w2079;
assign w34103 = ~w2098 & ~w12;
assign w34104 = ~w2115 & ~w421;
assign w34105 = ~w2126 & ~w1298;
assign w34106 = ~w2182 & ~w989;
assign w34107 = ~w2200 & ~w660;
assign w34108 = ~w2225 & ~w242;
assign w34109 = ~w2243 & ~w102;
assign w34110 = ~w2219 & ~w2217;
assign w34111 = ~w2270 & ~w660;
assign w34112 = ~w2280 & ~w989;
assign w34113 = w1694 & w36482;
assign w34114 = w1295 & w36483;
assign w34115 = ~w2355 & ~w421;
assign w34116 = ~w2371 & ~w242;
assign w34117 = ~w2389 & ~w102;
assign w34118 = ~w2105 & ~w2104;
assign w34119 = ~w2406 & ~w12;
assign w34120 = ~w2429 & ~w102;
assign w34121 = ~w2439 & ~w660;
assign w34122 = ~w2450 & ~w989;
assign w34123 = ~w2461 & ~w1697;
assign w34124 = ~w2499 & ~w1298;
assign w34125 = w418 & w36484;
assign w34126 = ~w2547 & ~w242;
assign w34127 = ~w2401 & ~w2399;
assign w34128 = ~w2413 & ~w2412;
assign w34129 = w2579 & w2412;
assign w34130 = w2579 & ~w34128;
assign w34131 = ~w2579 & ~w2412;
assign w34132 = ~w2579 & w34128;
assign w34133 = ~w2572 & ~w12;
assign w34134 = ~w2595 & ~w102;
assign w34135 = ~w2607 & ~w1697;
assign w34136 = ~w2663 & ~w1298;
assign w34137 = w986 & w36485;
assign w34138 = w657 & w36486;
assign w34139 = w418 & w36487;
assign w34140 = ~w2736 & ~w242;
assign w34141 = ~w2761 & ~w12;
assign w34142 = ~w2755 & ~w2753;
assign w34143 = ~w2784 & ~w102;
assign w34144 = ~w2795 & ~w989;
assign w34145 = ~w2806 & ~w1298;
assign w34146 = w1694 & w36488;
assign w34147 = w657 & w36489;
assign w34148 = ~w2901 & ~w421;
assign w34149 = ~w2918 & ~w242;
assign w34150 = ~w27206 & ~w2927;
assign w34151 = w27206 & ~w2927;
assign w34152 = ~w2944 & ~w12;
assign w34153 = (~w2757 & w36490) | (~w2757 & w36491) | (w36490 & w36491);
assign w34154 = ~w2938 & w36492;
assign w34155 = ~w2969 & ~w989;
assign w34156 = ~w2980 & ~w1298;
assign w34157 = ~w2991 & ~w2161;
assign w34158 = ~w3029 & ~w1697;
assign w34159 = w657 & w36493;
assign w34160 = ~w3077 & ~w421;
assign w34161 = ~w3094 & ~w242;
assign w34162 = ~w3110 & ~w102;
assign w34163 = (~w2753 & ~w2935) | (~w2753 & w36494) | (~w2935 & w36494);
assign w34164 = ~w2936 & w28240;
assign w34165 = ~w2767 & ~w2950;
assign w34166 = ~w2951 & ~w2950;
assign w34167 = ~w3128 & ~w12;
assign w34168 = ~w2778 & ~w2960;
assign w34169 = ~w3152 & ~w989;
assign w34170 = ~w3163 & ~w2161;
assign w34171 = w1694 & w36495;
assign w34172 = ~w3237 & ~w1298;
assign w34173 = w657 & w36496;
assign w34174 = (a_14 & ~w657) | (a_14 & w36497) | (~w657 & w36497);
assign w34175 = w418 & w36498;
assign w34176 = ~w3299 & ~w242;
assign w34177 = ~w3317 & ~w102;
assign w34178 = ~w3135 & ~w3134;
assign w34179 = w3342 & w3134;
assign w34180 = w3342 & ~w34178;
assign w34181 = ~w3342 & ~w3134;
assign w34182 = ~w3342 & w34178;
assign w34183 = ~w3361 & ~w242;
assign w34184 = ~w3373 & ~w989;
assign w34185 = w2158 & w36499;
assign w34186 = ~w3439 & ~w1697;
assign w34187 = ~w3455 & ~w1298;
assign w34188 = ~w3479 & ~w660;
assign w34189 = w418 & w36500;
assign w34190 = ~w3518 & ~w102;
assign w34191 = ~w3342 & ~w3341;
assign w34192 = w3542 & w3341;
assign w34193 = w3542 & ~w34191;
assign w34194 = ~w3542 & ~w3341;
assign w34195 = ~w3542 & w34191;
assign w34196 = ~w3535 & ~w12;
assign w34197 = ~w3559 & ~w242;
assign w34198 = ~w3572 & ~w1298;
assign w34199 = ~w3583 & ~w2642;
assign w34200 = ~w3621 & ~w2161;
assign w34201 = w1694 & w36501;
assign w34202 = ~w3660 & ~w989;
assign w34203 = ~w3676 & ~w660;
assign w34204 = w418 & w36502;
assign w34205 = ~w3717 & ~w102;
assign w34206 = ~w3541 & ~w3542;
assign w34207 = (~w3541 & ~w3542) | (~w3541 & w36503) | (~w3542 & w36503);
assign w34208 = ~w3734 & ~w12;
assign w34209 = ~w3760 & ~w2161;
assign w34210 = ~w3771 & ~w2642;
assign w34211 = ~w3835 & ~w1697;
assign w34212 = ~w3852 & ~w1298;
assign w34213 = w986 & w36504;
assign w34214 = w657 & w36505;
assign w34215 = w418 & w36506;
assign w34216 = w239 & w36507;
assign w34217 = ~w3711 & ~w3709;
assign w34218 = ~w3940 & ~w102;
assign w34219 = ~w3957 & ~w12;
assign w34220 = w239 & w36508;
assign w34221 = ~w3991 & ~w421;
assign w34222 = ~w4003 & ~w1298;
assign w34223 = ~w4014 & ~w2161;
assign w34224 = w2639 & w36509;
assign w34225 = ~w4083 & ~w1697;
assign w34226 = ~w4107 & ~w989;
assign w34227 = ~w4124 & ~w660;
assign w34228 = ~w4154 & ~w102;
assign w34229 = ~w3740 & ~w3963;
assign w34230 = ~w3964 & ~w3963;
assign w34231 = ~w4171 & ~w12;
assign w34232 = ~w4193 & ~w102;
assign w34233 = ~w4205 & ~w421;
assign w34234 = ~w4101 & ~w4099;
assign w34235 = ~w4218 & ~w1697;
assign w34236 = ~w4229 & ~w3198;
assign w34237 = ~w4267 & ~w2642;
assign w34238 = ~w4283 & ~w2161;
assign w34239 = ~w4307 & ~w1298;
assign w34240 = ~w4323 & ~w989;
assign w34241 = ~w4340 & ~w660;
assign w34242 = ~w4363 & ~w242;
assign w34243 = ~w4178 & ~w4177;
assign w34244 = w4392 & w4177;
assign w34245 = w4392 & ~w34243;
assign w34246 = ~w4392 & ~w4177;
assign w34247 = ~w4392 & w34243;
assign w34248 = ~w4403 & ~w4401;
assign w34249 = ~w4411 & ~w102;
assign w34250 = ~w4422 & ~w242;
assign w34251 = ~w4434 & ~w1697;
assign w34252 = ~w4445 & ~w2161;
assign w34253 = ~w4456 & ~w2642;
assign w34254 = ~w4467 & ~w3198;
assign w34255 = ~w4543 & ~w1298;
assign w34256 = ~w4561 & ~w989;
assign w34257 = ~w4579 & ~w660;
assign w34258 = ~w4596 & ~w421;
assign w34259 = ~w4392 & ~w4391;
assign w34260 = w4633 & w4391;
assign w34261 = w4633 & ~w34259;
assign w34262 = ~w4633 & ~w4391;
assign w34263 = ~w4633 & w34259;
assign w34264 = ~w4626 & ~w12;
assign w34265 = ~w4632 & ~w4633;
assign w34266 = (~w4632 & ~w4633) | (~w4632 & w36510) | (~w4633 & w36510);
assign w34267 = w4632 & w4655;
assign w34268 = w4655 & ~w34265;
assign w34269 = w4655 & ~w34266;
assign w34270 = ~w4632 & ~w4655;
assign w34271 = ~w4648 & ~w12;
assign w34272 = ~w4665 & ~w102;
assign w34273 = ~w4676 & ~w242;
assign w34274 = ~w4687 & ~w421;
assign w34275 = ~w4698 & ~w1697;
assign w34276 = ~w4710 & ~w2642;
assign w34277 = w3195 & w36511;
assign w34278 = ~w4778 & ~w2161;
assign w34279 = ~w4802 & ~w1298;
assign w34280 = ~w4820 & ~w989;
assign w34281 = ~w4836 & ~w660;
assign w34282 = ~w4878 & ~w12;
assign w34283 = w239 & w36512;
assign w34284 = (a_8 & ~w239) | (a_8 & w36513) | (~w239 & w36513);
assign w34285 = ~w4908 & ~w660;
assign w34286 = ~w4920 & ~w2161;
assign w34287 = ~w4930 & ~w3806;
assign w34288 = ~w4970 & ~w3198;
assign w34289 = ~w4988 & ~w2642;
assign w34290 = ~w5012 & ~w1697;
assign w34291 = ~w5028 & ~w1298;
assign w34292 = ~w5046 & ~w989;
assign w34293 = ~w5069 & ~w421;
assign w34294 = ~w5092 & ~w102;
assign w34295 = ~w5118 & ~w102;
assign w34296 = ~w5129 & ~w242;
assign w34297 = ~w5142 & ~w660;
assign w34298 = ~w5152 & ~w2161;
assign w34299 = ~w5164 & ~w3806;
assign w34300 = ~w5222 & ~w3198;
assign w34301 = ~w5239 & ~w2642;
assign w34302 = ~w5263 & ~w1697;
assign w34303 = ~w5281 & ~w1298;
assign w34304 = ~w5299 & ~w989;
assign w34305 = ~w5324 & ~w421;
assign w34306 = ~w4654 & ~w4884;
assign w34307 = ~w5353 & ~w12;
assign w34308 = w239 & w36514;
assign w34309 = (a_8 & ~w239) | (a_8 & w36515) | (~w239 & w36515);
assign w34310 = w418 & w36516;
assign w34311 = ~w5401 & ~w660;
assign w34312 = ~w5413 & ~w1697;
assign w34313 = ~w5424 & ~w2161;
assign w34314 = ~w5435 & ~w2642;
assign w34315 = ~w5216 & ~w5214;
assign w34316 = w3803 & w36517;
assign w34317 = ~w5497 & ~w3198;
assign w34318 = ~w5533 & ~w1298;
assign w34319 = ~w5549 & ~w989;
assign w34320 = ~w5584 & ~w102;
assign w34321 = ~w5360 & ~w5359;
assign w34322 = ~w5599 & ~w12;
assign w34323 = ~w5622 & ~w102;
assign w34324 = w418 & w36518;
assign w34325 = ~w5646 & ~w989;
assign w34326 = ~w5656 & ~w1697;
assign w34327 = ~w5669 & ~w3198;
assign w34328 = ~w5680 & ~w4502;
assign w34329 = ~w5719 & ~w3806;
assign w34330 = ~w5743 & ~w2642;
assign w34331 = ~w5760 & ~w2161;
assign w34332 = ~w5784 & ~w1298;
assign w34333 = ~w5807 & ~w660;
assign w34334 = w239 & w36519;
assign w34335 = ~w5606 & ~w5605;
assign w34336 = w5861 & w5605;
assign w34337 = w5861 & ~w34335;
assign w34338 = ~w5861 & ~w5605;
assign w34339 = ~w5861 & w34335;
assign w34340 = ~w5854 & ~w12;
assign w34341 = w5860 & w5885;
assign w34342 = ~w5860 & ~w5885;
assign w34343 = ~w5878 & ~w12;
assign w34344 = ~w5896 & ~w421;
assign w34345 = ~w5802 & ~w5800;
assign w34346 = ~w5908 & ~w989;
assign w34347 = ~w5918 & ~w2642;
assign w34348 = ~w5930 & ~w4502;
assign w34349 = ~w5988 & ~w3806;
assign w34350 = ~w6005 & ~w3198;
assign w34351 = ~w6029 & ~w2161;
assign w34352 = ~w6047 & ~w1697;
assign w34353 = ~w6065 & ~w1298;
assign w34354 = ~w6089 & ~w660;
assign w34355 = ~w6114 & ~w242;
assign w34356 = ~w6131 & ~w102;
assign w34357 = ~w6157 & ~w102;
assign w34358 = ~w6167 & ~w421;
assign w34359 = ~w6178 & ~w660;
assign w34360 = ~w6189 & ~w989;
assign w34361 = ~w6201 & ~w2161;
assign w34362 = ~w6211 & ~w2642;
assign w34363 = ~w6222 & ~w3198;
assign w34364 = ~w5982 & ~w5980;
assign w34365 = w4499 & w36520;
assign w34366 = ~w6284 & ~w3806;
assign w34367 = ~w6320 & ~w1697;
assign w34368 = ~w6337 & ~w1298;
assign w34369 = w239 & w36521;
assign w34370 = ~w5884 & ~w5885;
assign w34371 = (~w5884 & ~w5885) | (~w5884 & w36522) | (~w5885 & w36522);
assign w34372 = w6405 & ~w34370;
assign w34373 = w6405 & ~w34371;
assign w34374 = ~w6405 & w34370;
assign w34375 = ~w6405 & w34371;
assign w34376 = ~w6398 & ~w12;
assign w34377 = ~w6424 & ~w660;
assign w34378 = ~w6436 & ~w1298;
assign w34379 = ~w6446 & ~w2161;
assign w34380 = ~w6459 & ~w3806;
assign w34381 = ~w6470 & ~w5199;
assign w34382 = ~w6509 & ~w4502;
assign w34383 = ~w6533 & ~w3198;
assign w34384 = ~w6550 & ~w2642;
assign w34385 = ~w6574 & ~w1697;
assign w34386 = ~w6597 & ~w989;
assign w34387 = ~w6620 & ~w421;
assign w34388 = w239 & w36523;
assign w34389 = (a_8 & ~w239) | (a_8 & w36524) | (~w239 & w36524);
assign w34390 = ~w6654 & ~w102;
assign w34391 = ~w6672 & ~w12;
assign w34392 = ~w6695 & ~w660;
assign w34393 = ~w6707 & ~w1298;
assign w34394 = ~w6717 & ~w3198;
assign w34395 = ~w6729 & ~w5199;
assign w34396 = ~w6787 & ~w4502;
assign w34397 = ~w6804 & ~w3806;
assign w34398 = ~w6828 & ~w2642;
assign w34399 = ~w6846 & ~w2161;
assign w34400 = ~w6568 & ~w6566;
assign w34401 = ~w6864 & ~w1697;
assign w34402 = ~w6888 & ~w989;
assign w34403 = ~w6912 & ~w421;
assign w34404 = ~w6930 & ~w242;
assign w34405 = ~w6946 & ~w102;
assign w34406 = ~w6404 & ~w6678;
assign w34407 = ~w6964 & ~w12;
assign w34408 = ~w6971 & ~w6970;
assign w34409 = ~w6988 & ~w12;
assign w34410 = ~w7005 & ~w660;
assign w34411 = ~w7016 & ~w989;
assign w34412 = ~w7027 & ~w1298;
assign w34413 = ~w7040 & ~w3198;
assign w34414 = ~w7051 & ~w3806;
assign w34415 = ~w6781 & ~w6779;
assign w34416 = w5196 & w36525;
assign w34417 = ~w7113 & ~w4502;
assign w34418 = ~w7143 & ~w2642;
assign w34419 = ~w7161 & ~w2161;
assign w34420 = ~w7178 & ~w1697;
assign w34421 = w418 & w36526;
assign w34422 = ~w7232 & ~w242;
assign w34423 = ~w7249 & ~w102;
assign w34424 = w7281 & w6994;
assign w34425 = w7281 & ~w25060;
assign w34426 = ~w7281 & ~w6994;
assign w34427 = ~w7281 & w25060;
assign w34428 = ~w7274 & ~w12;
assign w34429 = ~w7292 & ~w989;
assign w34430 = ~w7303 & ~w1697;
assign w34431 = ~w7314 & ~w3806;
assign w34432 = ~w7325 & ~w4502;
assign w34433 = ~w7336 & ~w5965;
assign w34434 = ~w7375 & ~w5199;
assign w34435 = ~w7404 & ~w3198;
assign w34436 = ~w7422 & ~w2642;
assign w34437 = ~w7440 & ~w2161;
assign w34438 = ~w7463 & ~w1298;
assign w34439 = w657 & w36527;
assign w34440 = w239 & w36528;
assign w34441 = ~w7537 & ~w102;
assign w34442 = ~w7549 & w7289;
assign w34443 = w7549 & ~w7289;
assign w34444 = ~w7559 & ~w1697;
assign w34445 = ~w7569 & ~w3806;
assign w34446 = ~w7581 & ~w5965;
assign w34447 = ~w7639 & ~w5199;
assign w34448 = ~w7656 & ~w4502;
assign w34449 = ~w7680 & ~w3198;
assign w34450 = ~w7698 & ~w2642;
assign w34451 = ~w7716 & ~w2161;
assign w34452 = ~w7741 & ~w1298;
assign w34453 = ~w7759 & ~w989;
assign w34454 = w657 & w36529;
assign w34455 = w239 & w36530;
assign w34456 = ~w7831 & ~w102;
assign w34457 = (~w7280 & ~w7281) | (~w7280 & w36531) | (~w7281 & w36531);
assign w34458 = (~w7280 & w26580) | (~w7280 & w25060) | (w26580 & w25060);
assign w34459 = ~w7849 & ~w12;
assign w34460 = ~w7872 & ~w989;
assign w34461 = ~w7883 & ~w1298;
assign w34462 = ~w7894 & ~w1697;
assign w34463 = ~w7907 & ~w3806;
assign w34464 = ~w7918 & ~w4502;
assign w34465 = ~w7633 & ~w7631;
assign w34466 = w5962 & w36532;
assign w34467 = ~w7979 & ~w5199;
assign w34468 = ~w8010 & ~w3198;
assign w34469 = ~w8028 & ~w2642;
assign w34470 = ~w8045 & ~w2161;
assign w34471 = w657 & w36533;
assign w34472 = (a_11 & ~w418) | (a_11 & w36534) | (~w418 & w36534);
assign w34473 = w239 & w36535;
assign w34474 = w99 & w36536;
assign w34475 = w8159 & ~w26583;
assign w34476 = w8159 & ~w26582;
assign w34477 = ~w8159 & w26583;
assign w34478 = ~w8159 & w26582;
assign w34479 = ~w8152 & ~w12;
assign w34480 = w8158 & w8183;
assign w34481 = ~w8158 & ~w8183;
assign w34482 = ~w8176 & ~w12;
assign w34483 = ~w8216 & ~w2161;
assign w34484 = ~w8227 & ~w3806;
assign w34485 = ~w8238 & ~w4502;
assign w34486 = ~w8249 & ~w5199;
assign w34487 = ~w8259 & ~w6764;
assign w34488 = ~w8298 & ~w5965;
assign w34489 = ~w8333 & ~w3198;
assign w34490 = ~w8351 & ~w2642;
assign w34491 = ~w8374 & ~w1697;
assign w34492 = w986 & w36537;
assign w34493 = ~w8455 & ~w102;
assign w34494 = ~w8482 & ~w4502;
assign w34495 = ~w8494 & ~w6764;
assign w34496 = ~w8552 & ~w5965;
assign w34497 = ~w8568 & ~w5199;
assign w34498 = ~w8592 & ~w3806;
assign w34499 = ~w8609 & ~w3198;
assign w34500 = ~w8627 & ~w2642;
assign w34501 = ~w8644 & ~w2161;
assign w34502 = w1694 & w36538;
assign w34503 = w1295 & w36539;
assign w34504 = ~w8450 & ~w8448;
assign w34505 = ~w8766 & ~w102;
assign w34506 = ~w8183 & ~w8182;
assign w34507 = (~w8182 & ~w8183) | (~w8182 & w36540) | (~w8183 & w36540);
assign w34508 = w8790 & ~w34507;
assign w34509 = w8790 & ~w34506;
assign w34510 = ~w8790 & w34507;
assign w34511 = ~w8790 & w34506;
assign w34512 = ~w8783 & ~w12;
assign w34513 = ~w8778 & ~w8776;
assign w34514 = w1295 & w36541;
assign w34515 = w1694 & w36542;
assign w34516 = ~w8829 & ~w2161;
assign w34517 = ~w8841 & ~w3198;
assign w34518 = ~w8852 & ~w4502;
assign w34519 = ~w8863 & ~w5199;
assign w34520 = ~w8873 & ~w5965;
assign w34521 = w6761 & w36543;
assign w34522 = ~w8955 & ~w3806;
assign w34523 = ~w8978 & ~w2642;
assign w34524 = ~w9085 & ~w102;
assign w34525 = ~w25084 & ~w9095;
assign w34526 = w26814 & w26815;
assign w34527 = (w26815 & w26814) | (w26815 & ~w8158) | (w26814 & ~w8158);
assign w34528 = w9107 & ~w34527;
assign w34529 = w9107 & ~w34526;
assign w34530 = w9107 & ~w26815;
assign w34531 = w9107 & ~w26814;
assign w34532 = ~w9107 & w34527;
assign w34533 = ~w9107 & w34526;
assign w34534 = ~w9100 & ~w12;
assign w34535 = (w9115 & ~w25565) | (w9115 & w36544) | (~w25565 & w36544);
assign w34536 = ~w8806 & w36545;
assign w34537 = w25565 & w36546;
assign w34538 = (~w9115 & w8806) | (~w9115 & w36547) | (w8806 & w36547);
assign w34539 = (~w9115 & ~w25565) | (~w9115 & w36548) | (~w25565 & w36548);
assign w34540 = ~w8806 & w36549;
assign w34541 = ~w9106 & ~w34531;
assign w34542 = (~w9106 & w26815) | (~w9106 & w36550) | (w26815 & w36550);
assign w34543 = w9106 & w9131;
assign w34544 = (~w26815 & w34543) | (~w26815 & w36551) | (w34543 & w36551);
assign w34545 = (w9131 & w34531) | (w9131 & w34543) | (w34531 & w34543);
assign w34546 = ~w9106 & ~w9131;
assign w34547 = (w26815 & w34546) | (w26815 & w36552) | (w34546 & w36552);
assign w34548 = ~w34531 & w34546;
assign w34549 = ~w9124 & ~w12;
assign w34550 = ~w9154 & ~w2161;
assign w34551 = ~w9165 & ~w2642;
assign w34552 = ~w9175 & ~w3198;
assign w34553 = ~w9186 & ~w3806;
assign w34554 = w4499 & w36553;
assign w34555 = ~w9208 & ~w5199;
assign w34556 = ~w9219 & ~w5965;
assign w34557 = ~w9230 & ~w6764;
assign w34558 = ~w9240 & ~w7616;
assign w34559 = w1295 & w36554;
assign w34560 = w239 & w36555;
assign w34561 = ~w9423 & ~w102;
assign w34562 = ~w9095 & ~w9434;
assign w34563 = ~w9446 & ~w102;
assign w34564 = w239 & w36556;
assign w34565 = ~w9469 & ~w5199;
assign w34566 = ~w9480 & ~w5965;
assign w34567 = ~w9491 & ~w6764;
assign w34568 = ~w9502 & ~w7616;
assign w34569 = ~w9578 & ~w4502;
assign w34570 = ~w9595 & ~w3806;
assign w34571 = ~w9613 & ~w3198;
assign w34572 = w2639 & w36557;
assign w34573 = w2158 & w36558;
assign w34574 = w1694 & w36559;
assign w34575 = ~w9131 & ~w9130;
assign w34576 = (~w9130 & ~w9131) | (~w9130 & w36560) | (~w9131 & w36560);
assign w34577 = ~w9765 & ~w12;
assign w34578 = ~w9788 & ~w12;
assign w34579 = ~w9806 & ~w242;
assign w34580 = ~w9841 & ~w5199;
assign w34581 = ~w9852 & ~w5965;
assign w34582 = ~w9863 & ~w6764;
assign w34583 = w7613 & w36561;
assign w34584 = ~w9945 & ~w4502;
assign w34585 = ~w9962 & ~w3806;
assign w34586 = w3195 & w36562;
assign w34587 = ~w9995 & ~w2642;
assign w34588 = ~w10101 & ~w102;
assign w34589 = ~w10126 & ~w102;
assign w34590 = ~w10137 & ~w242;
assign w34591 = ~w10172 & ~w2642;
assign w34592 = ~w10183 & ~w4502;
assign w34593 = w5196 & w36563;
assign w34594 = ~w10205 & ~w5965;
assign w34595 = ~w10216 & ~w6764;
assign w34596 = ~w10227 & ~w8529;
assign w34597 = ~w10265 & ~w7616;
assign w34598 = ~w10306 & ~w3806;
assign w34599 = ~w10324 & ~w3198;
assign w34600 = w1694 & w36564;
assign w34601 = ~w10442 & ~w12;
assign w34602 = ~w10449 & ~w10448;
assign w34603 = w10473 & w10448;
assign w34604 = w10473 & ~w34602;
assign w34605 = ~w10473 & ~w10448;
assign w34606 = ~w10473 & w34602;
assign w34607 = ~w10466 & ~w12;
assign w34608 = ~w10482 & ~w102;
assign w34609 = w239 & w36565;
assign w34610 = ~w10519 & ~w7616;
assign w34611 = ~w10530 & ~w8529;
assign w34612 = ~w10594 & ~w6764;
assign w34613 = ~w10611 & ~w5965;
assign w34614 = ~w10629 & ~w5199;
assign w34615 = ~w10646 & ~w4502;
assign w34616 = w3803 & w36566;
assign w34617 = w2639 & w36567;
assign w34618 = ~w10831 & ~w242;
assign w34619 = w6761 & w36568;
assign w34620 = ~w10889 & ~w7616;
assign w34621 = w8526 & w36569;
assign w34622 = ~w10972 & ~w5199;
assign w34623 = ~w10989 & ~w4502;
assign w34624 = w3803 & w36570;
assign w34625 = w2639 & w36571;
assign w34626 = ~w11146 & ~w102;
assign w34627 = w26221 | w26222;
assign w34628 = (w26222 & w26221) | (w26222 & ~w10449) | (w26221 & ~w10449);
assign w34629 = ~w11159 & ~w12;
assign w34630 = w11177 & ~w10820;
assign w34631 = ~w11179 & ~w11178;
assign w34632 = w11174 & w11155;
assign w34633 = w11174 & ~w26220;
assign w34634 = w11165 & w11193;
assign w34635 = ~w11165 & ~w11193;
assign w34636 = ~w11202 & ~w102;
assign w34637 = ~w11213 & ~w242;
assign w34638 = ~w11269 & ~w5199;
assign w34639 = ~w11291 & ~w6764;
assign w34640 = ~w11302 & ~w7616;
assign w34641 = ~w11313 & ~w9537;
assign w34642 = ~w11350 & ~w8529;
assign w34643 = w4499 & w36572;
assign w34644 = w3195 & w36573;
assign w34645 = ~w11539 & ~w242;
assign w34646 = w418 & w36574;
assign w34647 = ~w11577 & ~w8529;
assign w34648 = ~w11588 & ~w9537;
assign w34649 = ~w11652 & ~w7616;
assign w34650 = ~w11669 & ~w6764;
assign w34651 = ~w11687 & ~w5965;
assign w34652 = ~w11703 & ~w5199;
assign w34653 = w4499 & w36575;
assign w34654 = w2639 & w36576;
assign w34655 = ~w11878 & ~w102;
assign w34656 = ~w11192 & ~w11193;
assign w34657 = (~w11192 & ~w11193) | (~w11192 & w36577) | (~w11193 & w36577);
assign w34658 = w11898 & ~w34656;
assign w34659 = w11898 & ~w34657;
assign w34660 = ~w11898 & w34656;
assign w34661 = ~w11898 & w34657;
assign w34662 = ~w11891 & ~w12;
assign w34663 = w11211 & w11201;
assign w34664 = w11887 & w11906;
assign w34665 = ~w11935 & ~w6764;
assign w34666 = ~w11945 & ~w7616;
assign w34667 = ~w11956 & ~w8529;
assign w34668 = w10562 & w36578;
assign w34669 = w9534 & w36579;
assign w34670 = ~w12039 & ~w5965;
assign w34671 = ~w12055 & ~w5199;
assign w34672 = w4499 & w36580;
assign w34673 = w2639 & w36581;
assign w34674 = ~w12217 & ~w421;
assign w34675 = ~w12233 & ~w242;
assign w34676 = w12250 & w29583;
assign w34677 = w12250 & w29582;
assign w34678 = (w25442 & w25441) | (w25442 & ~w11193) | (w25441 & ~w11193);
assign w34679 = (w25442 & w25441) | (w25442 & ~w34634) | (w25441 & ~w34634);
assign w34680 = w12270 & ~w34679;
assign w34681 = w12270 & ~w34678;
assign w34682 = ~w12270 & w34679;
assign w34683 = ~w12270 & w34678;
assign w34684 = ~w12263 & ~w12;
assign w34685 = w657 & w36582;
assign w34686 = ~w12345 & ~w5965;
assign w34687 = ~w12356 & ~w7616;
assign w34688 = ~w12368 & ~w9537;
assign w34689 = ~w12401 & ~w10565;
assign w34690 = ~w12424 & ~w8529;
assign w34691 = ~w12448 & ~w6764;
assign w34692 = ~w12470 & ~w5199;
assign w34693 = w4499 & w36583;
assign w34694 = w2639 & w36584;
assign w34695 = w418 & w36585;
assign w34696 = ~w12607 & ~w242;
assign w34697 = w99 & w36586;
assign w34698 = w12242 & w12255;
assign w34699 = (~w12269 & w25134) | (~w12269 & w34679) | (w25134 & w34679);
assign w34700 = (~w12269 & w25134) | (~w12269 & w34678) | (w25134 & w34678);
assign w34701 = ~w12643 & w12269;
assign w34702 = ~w12643 & ~w25134;
assign w34703 = (~w34678 & w34701) | (~w34678 & w34702) | (w34701 & w34702);
assign w34704 = (~w34679 & w34701) | (~w34679 & w34702) | (w34701 & w34702);
assign w34705 = w12643 & ~w12269;
assign w34706 = w12643 & w25134;
assign w34707 = (w34678 & w34705) | (w34678 & w34706) | (w34705 & w34706);
assign w34708 = (w34679 & w34705) | (w34679 & w34706) | (w34705 & w34706);
assign w34709 = ~w12636 & ~w12;
assign w34710 = (~w12245 & w36587) | (~w12245 & w36588) | (w36587 & w36588);
assign w34711 = (~b_62 & w12643) | (~b_62 & w36589) | (w12643 & w36589);
assign w34712 = (~b_62 & w25134) | (~b_62 & w36590) | (w25134 & w36590);
assign w34713 = b_63 & ~w34711;
assign w34714 = b_63 & ~w34712;
assign w34715 = w12641 & w12269;
assign w34716 = (w12641 & w12270) | (w12641 & w34715) | (w12270 & w34715);
assign w34717 = ~w29812 & w36591;
assign w34718 = (~w29747 & w36592) | (~w29747 & w36593) | (w36592 & w36593);
assign w34719 = w4 & w36594;
assign w34720 = ~w12681 & ~w421;
assign w34721 = w657 & w36595;
assign w34722 = w3195 & w36596;
assign w34723 = ~w12735 & ~w5965;
assign w34724 = ~w12745 & ~w7616;
assign w34725 = ~w12755 & ~w9537;
assign w34726 = ~w12788 & ~w10565;
assign w34727 = ~w12812 & ~w8529;
assign w34728 = ~w12837 & ~w6764;
assign w34729 = ~w12862 & ~w5199;
assign w34730 = w4499 & w36597;
assign w34731 = w1694 & w36598;
assign w34732 = ~w13000 & ~w242;
assign w34733 = w99 & w36599;
assign w34734 = ~w13037 & ~w660;
assign w34735 = ~w13065 & ~w8529;
assign w34736 = w11620 & w36600;
assign w34737 = ~w13092 & ~w12780;
assign w34738 = w13092 & w12780;
assign w34739 = w10562 & w36601;
assign w34740 = ~w13116 & ~w9537;
assign w34741 = ~w13139 & ~w7616;
assign w34742 = ~w13155 & ~w6764;
assign w34743 = ~w13172 & ~w5965;
assign w34744 = ~w13188 & ~w5199;
assign w34745 = ~w13206 & ~w4502;
assign w34746 = w3803 & w36602;
assign w34747 = ~w13241 & ~w3198;
assign w34748 = w2639 & w36603;
assign w34749 = ~w12955 & ~w12967;
assign w34750 = w986 & w36604;
assign w34751 = ~w13342 & ~w421;
assign w34752 = ~w13355 & ~w242;
assign w34753 = ~w13371 & ~w102;
assign w34754 = ~w8 & w29810;
assign w34755 = w12 & w34713;
assign w34756 = ~w34712 & w36605;
assign w34757 = ~w13405 & ~w102;
assign w34758 = ~w13419 & ~w421;
assign w34759 = w1295 & w36606;
assign w34760 = ~w13473 & ~w2161;
assign w34761 = ~w13500 & ~w3806;
assign w34762 = ~w13510 & ~w5965;
assign w34763 = ~w13520 & ~w8529;
assign w34764 = ~w13552 & ~w10565;
assign w34765 = ~w13569 & ~w9537;
assign w34766 = ~w13593 & ~w7616;
assign w34767 = ~w13611 & ~w6764;
assign w34768 = ~w12848 & ~w13165;
assign w34769 = ~w13636 & ~w5199;
assign w34770 = ~w13654 & ~w4502;
assign w34771 = ~w13233 & ~w13683;
assign w34772 = ~w13731 & ~w242;
assign w34773 = w657 & w36607;
assign w34774 = w13469 & w13786;
assign w34775 = ~w13469 & ~w13786;
assign w34776 = w2158 & w36608;
assign w34777 = ~w13817 & ~w3806;
assign w34778 = ~w13828 & ~w8529;
assign w34779 = ~w13838 & ~w11623;
assign w34780 = (a_62 & w13853) | (a_62 & w36609) | (w13853 & w36609);
assign w34781 = ~w13863 & ~w10565;
assign w34782 = w13561 & ~w13548;
assign w34783 = w13561 & ~w29980;
assign w34784 = ~w13881 & ~w9537;
assign w34785 = ~w13907 & ~w7616;
assign w34786 = ~w13925 & ~w6764;
assign w34787 = ~w13944 & ~w5965;
assign w34788 = ~w13962 & ~w5199;
assign w34789 = ~w13629 & w36610;
assign w34790 = ~w13980 & ~w4502;
assign w34791 = ~w33983 & ~w14057;
assign w34792 = (w14109 & w29812) | (w14109 & w36611) | (w29812 & w36611);
assign w34793 = (w29747 & w36612) | (w29747 & w36613) | (w36612 & w36613);
assign w34794 = ~w102 & a_5;
assign w34795 = w102 & ~a_5;
assign w34796 = w14123 & w13755;
assign w34797 = w14145 & w29583;
assign w34798 = w14145 & w29582;
assign w34799 = ~w14164 & ~w14057;
assign w34800 = ~w13456 & w36614;
assign w34801 = (~w14164 & w14045) | (~w14164 & w36615) | (w14045 & w36615);
assign w34802 = w14164 & ~w14057;
assign w34803 = ~w13456 & w36616;
assign w34804 = (w14164 & w14045) | (w14164 & w36617) | (w14045 & w36617);
assign w34805 = w2639 & w36618;
assign w34806 = w13813 & w14218;
assign w34807 = ~w13813 & ~w14218;
assign w34808 = ~w14222 & ~w3806;
assign w34809 = ~w14232 & ~w6764;
assign w34810 = ~w14242 & ~w9537;
assign w34811 = w11620 & w36619;
assign w34812 = w30146 & ~w14269;
assign w34813 = ~w14278 & ~w10565;
assign w34814 = w13859 & w13872;
assign w34815 = ~w14304 & ~w8529;
assign w34816 = ~w13893 & w13837;
assign w34817 = ~w14322 & ~w7616;
assign w34818 = ~w14347 & ~w5965;
assign w34819 = ~w14365 & ~w5199;
assign w34820 = w13958 & w13971;
assign w34821 = ~w14383 & ~w4502;
assign w34822 = (~w13635 & w36620) | (~w13635 & w36621) | (w36620 & w36621);
assign w34823 = ~w13826 & ~w14412;
assign w34824 = w13826 & w14412;
assign w34825 = w14003 & ~w14432;
assign w34826 = w14003 & w14432;
assign w34827 = ~w30130 & ~w14440;
assign w34828 = w30130 & ~w14440;
assign w34829 = (w14154 & w36622) | (w14154 & w14468) | (w36622 & w14468);
assign w34830 = ~w14480 & ~w14121;
assign w34831 = ~w14490 & ~w242;
assign w34832 = ~w14070 & w36623;
assign w34833 = (w14080 & w36624) | (w14080 & w36625) | (w36624 & w36625);
assign w34834 = (~w14499 & w14456) | (~w14499 & w36626) | (w14456 & w36626);
assign w34835 = ~w14504 & ~w421;
assign w34836 = w986 & w36627;
assign w34837 = ~w14557 & w30182;
assign w34838 = w14014 & w36628;
assign w34839 = ~w14557 & ~w30182;
assign w34840 = (~w14557 & ~w14014) | (~w14557 & w36629) | (~w14014 & w36629);
assign w34841 = ~w14561 & ~w2642;
assign w34842 = ~w14395 & w14231;
assign w34843 = ~w14358 & w36630;
assign w34844 = (~w13898 & w36631) | (~w13898 & w36632) | (w36631 & w36632);
assign w34845 = w14274 & w14287;
assign w34846 = ~w14580 & ~w10565;
assign w34847 = ~w14602 & ~w11623;
assign w34848 = ~w14623 & ~w9537;
assign w34849 = (~w13862 & w36633) | (~w13862 & w36634) | (w36633 & w36634);
assign w34850 = ~w14640 & ~w8529;
assign w34851 = ~w14658 & ~w7616;
assign w34852 = ~w14674 & ~w6764;
assign w34853 = ~w14690 & ~w5965;
assign w34854 = ~w14708 & ~w5199;
assign w34855 = ~w14725 & ~w4502;
assign w34856 = ~w14742 & ~w3806;
assign w34857 = ~w14758 & ~w3198;
assign w34858 = w1295 & w36635;
assign w34859 = ~w14807 & ~w660;
assign w34860 = (w14834 & w25144) | (w14834 & w14121) | (w25144 & w14121);
assign w34861 = (w14841 & w29812) | (w14841 & w36636) | (w29812 & w36636);
assign w34862 = (w29747 & w36637) | (w29747 & w36638) | (w36637 & w36638);
assign w34863 = ~w242 & a_8;
assign w34864 = w242 & ~a_8;
assign w34865 = ~w14849 & ~w421;
assign w34866 = w986 & w36639;
assign w34867 = ~w14931 & ~w2642;
assign w34868 = w14767 & ~w14757;
assign w34869 = ~w14944 & ~w3198;
assign w34870 = w14751 & w14953;
assign w34871 = ~w14751 & ~w14953;
assign w34872 = ~w14957 & ~w3806;
assign w34873 = ~w14968 & ~w4502;
assign w34874 = ~w15001 & ~w10565;
assign w34875 = ~w15019 & ~w9537;
assign w34876 = ~w15037 & ~w8529;
assign w34877 = ~w15055 & ~w7616;
assign w34878 = ~w15074 & ~w6764;
assign w34879 = ~w15091 & ~w5965;
assign w34880 = ~w15108 & ~w5199;
assign w34881 = ~w15135 & w36640;
assign w34882 = (w14940 & w15135) | (w14940 & w36641) | (w15135 & w36641);
assign w34883 = w15135 | w15136;
assign w34884 = ~w15166 & ~w15165;
assign w34885 = w14898 & w15147;
assign w34886 = (~w14940 & w15135) | (~w14940 & w36642) | (w15135 & w36642);
assign w34887 = ~w14940 & w15220;
assign w34888 = ~w15126 & w14966;
assign w34889 = ~w15240 & ~w4502;
assign w34890 = ~w15250 & ~w6764;
assign w34891 = w15051 & w15064;
assign w34892 = ~w15261 & ~w7616;
assign w34893 = ~w14997 & w15010;
assign w34894 = ~w15282 & ~w11623;
assign w34895 = ~w15295 & ~w10565;
assign w34896 = ~w15311 & ~w9537;
assign w34897 = ~w15329 & ~w8529;
assign w34898 = ~w15069 & w36643;
assign w34899 = ~w15360 & ~w5965;
assign w34900 = ~w15378 & ~w5199;
assign w34901 = ~w15402 & ~w3806;
assign w34902 = (~w30373 & w15401) | (~w30373 & w36644) | (w15401 & w36644);
assign w34903 = w30369 & ~w15436;
assign w34904 = (w15220 & ~w15436) | (w15220 & w30369) | (~w15436 & w30369);
assign w34905 = ~w30369 & ~w15436;
assign w34906 = w15470 & w29583;
assign w34907 = w15470 & w29582;
assign w34908 = (~w15505 & w15164) | (~w15505 & w36645) | (w15164 & w36645);
assign w34909 = ~w15512 & ~w421;
assign w34910 = ~w15492 & ~w15521;
assign w34911 = ~w34910 & ~w15521;
assign w34912 = ~w15526 & ~w660;
assign w34913 = ~w15475 & w15535;
assign w34914 = w15475 & ~w15535;
assign w34915 = ~w15539 & ~w989;
assign w34916 = ~w15554 & ~w1298;
assign w34917 = (~w15453 & w15562) | (~w15453 & w36646) | (w15562 & w36646);
assign w34918 = (w15453 & w15562) | (w15453 & w36647) | (w15562 & w36647);
assign w34919 = ~w15568 & ~w2161;
assign w34920 = (~w15428 & w15591) | (~w15428 & w36648) | (w15591 & w36648);
assign w34921 = (w15428 & w15591) | (w15428 & w36649) | (w15591 & w36649);
assign w34922 = w15401 & w36650;
assign w34923 = (~w15129 & w36651) | (~w15129 & w36652) | (w36651 & w36652);
assign w34924 = ~w15598 & ~w3198;
assign w34925 = w15391 & w15249;
assign w34926 = w15374 & w15387;
assign w34927 = ~w15616 & ~w7616;
assign w34928 = ~w15626 & ~w9537;
assign w34929 = ~w15638 & ~w11623;
assign w34930 = ~w15663 & ~w10565;
assign w34931 = ~w15686 & ~w8529;
assign w34932 = ~w15712 & ~w6764;
assign w34933 = ~w15348 & w15259;
assign w34934 = ~w15729 & ~w5965;
assign w34935 = ~w15746 & ~w5199;
assign w34936 = ~w15763 & ~w4502;
assign w34937 = ~w15779 & ~w3806;
assign w34938 = ~w15797 & ~w15607;
assign w34939 = w1694 & w36653;
assign w34940 = w15506 & w36654;
assign w34941 = ~w15843 & w25149;
assign w34942 = (~w15841 & w25148) | (~w15841 & w36655) | (w25148 & w36655);
assign w34943 = (~w15841 & w25149) | (~w15841 & w36655) | (w25149 & w36655);
assign w34944 = ~w15850 & ~w660;
assign w34945 = w15548 & w15830;
assign w34946 = w1295 & w36656;
assign w34947 = w15818 & w15874;
assign w34948 = (w15874 & w15581) | (w15874 & w36657) | (w15581 & w36657);
assign w34949 = ~w15818 & ~w15874;
assign w34950 = ~w15581 & w36658;
assign w34951 = ~w15878 & ~w1697;
assign w34952 = w3195 & w36659;
assign w34953 = w15788 & w15916;
assign w34954 = ~w15788 & ~w15916;
assign w34955 = ~w15920 & ~w3806;
assign w34956 = ~w15931 & ~w4502;
assign w34957 = ~w15942 & ~w5199;
assign w34958 = ~w15952 & ~w11623;
assign w34959 = ~w15980 & ~w10565;
assign w34960 = ~w15998 & ~w9537;
assign w34961 = ~w16015 & ~w8529;
assign w34962 = ~w16032 & ~w7616;
assign w34963 = ~w16050 & ~w6764;
assign w34964 = ~w16068 & ~w5965;
assign w34965 = ~w15607 & ~w16114;
assign w34966 = ~w16114 & ~w15797;
assign w34967 = (~w16114 & ~w15797) | (~w16114 & w34965) | (~w15797 & w34965);
assign w34968 = ~w15607 & w16114;
assign w34969 = w16114 & ~w15797;
assign w34970 = (w16114 & ~w15797) | (w16114 & w34968) | (~w15797 & w34968);
assign w34971 = ~w16141 & ~w15563;
assign w34972 = ~w15444 & w36660;
assign w34973 = ~w16141 & w15563;
assign w34974 = (~w16141 & w15444) | (~w16141 & w36661) | (w15444 & w36661);
assign w34975 = ~w16149 & ~w15859;
assign w34976 = ~w15475 & ~w15535;
assign w34977 = (w16158 & w29812) | (w16158 & w36662) | (w29812 & w36662);
assign w34978 = (w29747 & w36663) | (w29747 & w36664) | (w36663 & w36664);
assign w34979 = ~w421 & a_11;
assign w34980 = w421 & ~a_11;
assign w34981 = ~w16162 & ~w33202;
assign w34982 = (~w16162 & ~w15552) | (~w16162 & w36665) | (~w15552 & w36665);
assign w34983 = (~w25148 & w36666) | (~w25148 & w36667) | (w36666 & w36667);
assign w34984 = (~w25149 & w36666) | (~w25149 & w36667) | (w36666 & w36667);
assign w34985 = ~w15841 & ~w16173;
assign w34986 = (w25148 & w36668) | (w25148 & w36669) | (w36668 & w36669);
assign w34987 = (w25149 & w36668) | (w25149 & w36669) | (w36668 & w36669);
assign w34988 = ~w15859 & ~w16185;
assign w34989 = w15859 & ~w16185;
assign w34990 = ~w16201 & ~w989;
assign w34991 = (~w15597 & w36670) | (~w15597 & w36671) | (w36670 & w36671);
assign w34992 = ~w15597 & w36672;
assign w34993 = ~w16238 & ~w33449;
assign w34994 = ~w16238 & ~w33448;
assign w34995 = (w15597 & w36673) | (w15597 & w36674) | (w36673 & w36674);
assign w34996 = (w16238 & w15597) | (w16238 & w36675) | (w15597 & w36675);
assign w34997 = w16238 & w33449;
assign w34998 = w16238 & w33448;
assign w34999 = (~w16263 & w15928) | (~w16263 & w36676) | (w15928 & w36676);
assign w35000 = ~w15928 & w36677;
assign w35001 = ~w16267 & ~w3806;
assign w35002 = ~w16278 & ~w5199;
assign w35003 = ~w16289 & ~w7616;
assign w35004 = ~w16300 & ~w8529;
assign w35005 = ~w15676 & w36678;
assign w35006 = ~w16323 & ~w11623;
assign w35007 = ~w16337 & ~w10565;
assign w35008 = ~w16354 & ~w9537;
assign w35009 = ~w16382 & ~w6764;
assign w35010 = ~w16400 & ~w5965;
assign w35011 = ~w16425 & ~w4502;
assign w35012 = ~w30625 & ~w16482;
assign w35013 = ~w16488 & w25153;
assign w35014 = ~w16488 & w25154;
assign w35015 = (~w16486 & w25153) | (~w16486 & w36679) | (w25153 & w36679);
assign w35016 = ~w16486 & ~w25156;
assign w35017 = w30625 & ~w16482;
assign w35018 = ~w16496 & ~w660;
assign w35019 = ~w16509 & ~w989;
assign w35020 = ~w16210 & w16518;
assign w35021 = w16210 & ~w16518;
assign w35022 = ~w16522 & ~w1298;
assign w35023 = w16224 & w16531;
assign w35024 = ~w16224 & ~w16531;
assign w35025 = w1694 & w36680;
assign w35026 = ~w16550 & ~w2161;
assign w35027 = ~w26370 & ~w30644;
assign w35028 = ~w26370 & ~w30643;
assign w35029 = ~w16437 & w16276;
assign w35030 = w16421 & w16434;
assign w35031 = w16396 & w16409;
assign w35032 = w16288 & w16391;
assign w35033 = ~w16584 & ~w8529;
assign w35034 = ~w16595 & ~w11623;
assign w35035 = w16613 & a_62;
assign w35036 = ~w16622 & ~w10565;
assign w35037 = ~w16640 & ~w9537;
assign w35038 = ~w16665 & ~w7616;
assign w35039 = w16299 & w16298;
assign w35040 = ~w16683 & ~w6764;
assign w35041 = ~w16692 & ~w30734;
assign w35042 = w16378 & w36681;
assign w35043 = ~w16701 & ~w5965;
assign w35044 = ~w16717 & ~w5199;
assign w35045 = ~w16733 & ~w4502;
assign w35046 = ~w16749 & ~w3806;
assign w35047 = w3195 & w36682;
assign w35048 = (w16094 & w36683) | (w16094 & w36684) | (w36683 & w36684);
assign w35049 = w16094 & w36683;
assign w35050 = w30778 & w16764;
assign w35051 = ~w30778 & ~w16764;
assign w35052 = (~w25153 & w36685) | (~w25153 & w36686) | (w36685 & w36686);
assign w35053 = (~w16803 & w25157) | (~w16803 & w25156) | (w25157 & w25156);
assign w35054 = ~w16486 & ~w16802;
assign w35055 = (w25153 & w36687) | (w25153 & w36688) | (w36687 & w36688);
assign w35056 = (w25158 & w25159) | (w25158 & ~w25156) | (w25159 & ~w25156);
assign w35057 = ~w16809 & ~w989;
assign w35058 = ~w16824 & ~w1697;
assign w35059 = ~w16781 & w36689;
assign w35060 = ~w16848 & ~w16775;
assign w35061 = (~w16097 & w36690) | (~w16097 & w36691) | (w36690 & w36691);
assign w35062 = ~w16848 & ~w35060;
assign w35063 = ~w16848 & ~w35061;
assign w35064 = ~w16854 & ~w3806;
assign w35065 = ~w16866 & ~w4502;
assign w35066 = ~w16877 & ~w5199;
assign w35067 = ~w16889 & ~w5965;
assign w35068 = ~w16899 & ~w6764;
assign w35069 = ~w16919 & ~w11623;
assign w35070 = (~a_62 & w16917) | (~a_62 & w36692) | (w16917 & w36692);
assign w35071 = w16917 | w36693;
assign w35072 = ~w16917 & w36694;
assign w35073 = ~w16934 & ~w10565;
assign w35074 = ~w16952 & ~w9537;
assign w35075 = ~w16970 & ~w8529;
assign w35076 = ~w16988 & ~w7616;
assign w35077 = ~w16758 & ~w17046;
assign w35078 = ~w16758 & w17046;
assign w35079 = w16574 & ~w27596;
assign w35080 = (~w16833 & w17073) | (~w16833 & w36695) | (w17073 & w36695);
assign w35081 = (~w17088 & ~w16563) | (~w17088 & w36696) | (~w16563 & w36696);
assign w35082 = ~w16210 & ~w16518;
assign w35083 = (w17105 & w29812) | (w17105 & w36697) | (w29812 & w36697);
assign w35084 = (w29747 & w36698) | (w29747 & w36699) | (w36698 & w36699);
assign w35085 = ~w660 & a_14;
assign w35086 = w660 & ~a_14;
assign w35087 = (~w25153 & w36700) | (~w25153 & w36701) | (w36700 & w36701);
assign w35088 = (w25160 & w25161) | (w25160 & w25156) | (w25161 & w25156);
assign w35089 = ~w17120 & w25158;
assign w35090 = (w25341 & w36702) | (w25341 & w36703) | (w36702 & w36703);
assign w35091 = ~w16818 & ~w17132;
assign w35092 = w16818 & ~w17132;
assign w35093 = ~w17136 & ~w1298;
assign w35094 = w16833 & w17145;
assign w35095 = ~w16833 & ~w17145;
assign w35096 = w1694 & w36704;
assign w35097 = ~w17163 & ~w2161;
assign w35098 = w17172 & w16848;
assign w35099 = (~w16445 & w36705) | (~w16445 & w36706) | (w36705 & w36706);
assign w35100 = ~w17172 & ~w16848;
assign w35101 = (w16445 & w36707) | (w16445 & w36708) | (w36707 & w36708);
assign w35102 = ~w16864 & w36709;
assign w35103 = ~w17188 & ~w3806;
assign w35104 = ~w17199 & ~w4502;
assign w35105 = ~w17212 & ~w8529;
assign w35106 = (a_62 & w16917) | (a_62 & w36710) | (w16917 & w36710);
assign w35107 = w17230 & w30914;
assign w35108 = w30913 & w36711;
assign w35109 = ~w17230 & ~w30914;
assign w35110 = (~w17230 & ~w30913) | (~w17230 & w36712) | (~w30913 & w36712);
assign w35111 = ~w17244 & ~w10565;
assign w35112 = w16929 & w16943;
assign w35113 = ~w17262 & ~w9537;
assign w35114 = ~w17284 & ~w7616;
assign w35115 = w16984 & w16997;
assign w35116 = ~w17303 & ~w6764;
assign w35117 = ~w17319 & ~w5965;
assign w35118 = ~w16696 & w36713;
assign w35119 = ~w17337 & ~w5199;
assign w35120 = ~w17036 & ~w17047;
assign w35121 = (w16546 & w36714) | (w16546 & w36715) | (w36714 & w36715);
assign w35122 = w16546 & w36714;
assign w35123 = (w17148 & w36716) | (w17148 & w17403) | (w36716 & w17403);
assign w35124 = (~w25158 & w36717) | (~w25158 & w36718) | (w36717 & w36718);
assign w35125 = (~w25341 & w36719) | (~w25341 & w36720) | (w36719 & w36720);
assign w35126 = (w25156 & w36721) | (w25156 & w36722) | (w36721 & w36722);
assign w35127 = (~w25153 & w36723) | (~w25153 & w36724) | (w36723 & w36724);
assign w35128 = (w25158 & w36725) | (w25158 & w36726) | (w36725 & w36726);
assign w35129 = (w25341 & w36727) | (w25341 & w36728) | (w36727 & w36728);
assign w35130 = (~w25156 & w36729) | (~w25156 & w36730) | (w36729 & w36730);
assign w35131 = (w25153 & w36731) | (w25153 & w36732) | (w36731 & w36732);
assign w35132 = ~w17422 & ~w989;
assign w35133 = ~w17436 & ~w1298;
assign w35134 = ~w30936 & w17145;
assign w35135 = ~w30936 & ~w30884;
assign w35136 = ~w17451 & ~w1697;
assign w35137 = ~w17464 & ~w2161;
assign w35138 = w17473 & w17172;
assign w35139 = (~w16778 & w36733) | (~w16778 & w36734) | (w36733 & w36734);
assign w35140 = ~w17473 & ~w17172;
assign w35141 = (w16778 & w36735) | (w16778 & w36736) | (w36735 & w36736);
assign w35142 = w2639 & w36737;
assign w35143 = (~w17011 & w36738) | (~w17011 & w36739) | (w36738 & w36739);
assign w35144 = ~w17507 & ~w11623;
assign w35145 = ~w17506 & a_62;
assign w35146 = ~w17525 & ~w10565;
assign w35147 = ~w17542 & ~w9537;
assign w35148 = ~w17559 & ~w8529;
assign w35149 = ~w17576 & ~w7616;
assign w35150 = ~w17280 & w17293;
assign w35151 = ~w17593 & ~w6764;
assign w35152 = ~w17610 & ~w5965;
assign w35153 = ~w17626 & ~w5199;
assign w35154 = ~w17643 & ~w4502;
assign w35155 = w17687 & ~w17676;
assign w35156 = (w25153 & w36741) | (w25153 & w36742) | (w36741 & w36742);
assign w35157 = (~w25158 & w36743) | (~w25158 & w36744) | (w36743 & w36744);
assign w35158 = (~w25341 & w36745) | (~w25341 & w36746) | (w36745 & w36746);
assign w35159 = (w25156 & w36747) | (w25156 & w36748) | (w36747 & w36748);
assign w35160 = (~w25153 & w36749) | (~w25153 & w36750) | (w36749 & w36750);
assign w35161 = ~w17711 & w35156;
assign w35162 = (~w25156 & w36751) | (~w25156 & w36752) | (w36751 & w36752);
assign w35163 = w17445 & w17701;
assign w35164 = (w17718 & w29812) | (w17718 & w36753) | (w29812 & w36753);
assign w35165 = (w29747 & w36754) | (w29747 & w36755) | (w36754 & w36755);
assign w35166 = ~w989 & a_17;
assign w35167 = w989 & ~a_17;
assign w35168 = ~w17726 & ~w1298;
assign w35169 = w17460 & ~w31016;
assign w35170 = ~w17748 & ~w17473;
assign w35171 = (w17054 & w36756) | (w17054 & w36757) | (w36756 & w36757);
assign w35172 = w17748 & w17473;
assign w35173 = (~w17054 & w36758) | (~w17054 & w36759) | (w36758 & w36759);
assign w35174 = ~w17752 & ~w2161;
assign w35175 = ~w17687 & ~w17775;
assign w35176 = w17687 & ~w17775;
assign w35177 = ~w17687 & w17775;
assign w35178 = ~w17793 & ~w4502;
assign w35179 = ~w17805 & ~w5199;
assign w35180 = ~w17816 & ~w5965;
assign w35181 = ~w17828 & ~w7616;
assign w35182 = w17843 & w31061;
assign w35183 = w17843 & w31062;
assign w35184 = ~w17843 & ~w31061;
assign w35185 = ~w17843 & ~w31062;
assign w35186 = ~w17857 & ~w10565;
assign w35187 = ~w17875 & ~w9537;
assign w35188 = ~w17892 & ~w8529;
assign w35189 = ~w17917 & ~w6764;
assign w35190 = ~w17955 & ~w3806;
assign w35191 = (w25158 & w36760) | (w25158 & w36761) | (w36760 & w36761);
assign w35192 = (w25341 & w36762) | (w25341 & w36763) | (w36762 & w36763);
assign w35193 = (~w25156 & w36764) | (~w25156 & w36765) | (w36764 & w36765);
assign w35194 = (w25168 & w25167) | (w25168 & w33977) | (w25167 & w33977);
assign w35195 = (w25158 & w36766) | (w25158 & w36767) | (w36766 & w36767);
assign w35196 = ~w17990 & w35192;
assign w35197 = (w33977 & w36768) | (w33977 & w36769) | (w36768 & w36769);
assign w35198 = (~w25156 & w36770) | (~w25156 & w36771) | (w36770 & w36771);
assign w35199 = (w25158 & w36772) | (w25158 & w36773) | (w36772 & w36773);
assign w35200 = w17722 & ~w31084;
assign w35201 = ~w18005 & ~w1298;
assign w35202 = ~w18019 & ~w1697;
assign w35203 = w2158 & w36774;
assign w35204 = w18043 & w17775;
assign w35205 = (w18043 & w17677) | (w18043 & w36775) | (w17677 & w36775);
assign w35206 = ~w18043 & ~w17775;
assign w35207 = ~w17677 & w36776;
assign w35208 = ~w17788 & ~w18056;
assign w35209 = ~w17657 & w36777;
assign w35210 = ~w18076 & ~w4502;
assign w35211 = ~w18087 & ~w5199;
assign w35212 = ~w17868 & w36778;
assign w35213 = ~w18099 & ~w9537;
assign w35214 = ~w18110 & ~w11623;
assign w35215 = ~w18124 & a_62;
assign w35216 = ~w17851 & w36779;
assign w35217 = ~w17851 & w36780;
assign w35218 = (w31132 & w17851) | (w31132 & w36781) | (w17851 & w36781);
assign w35219 = (w31133 & w17851) | (w31133 & w36782) | (w17851 & w36782);
assign w35220 = ~w18133 & ~w10565;
assign w35221 = ~w18155 & ~w8529;
assign w35222 = ~w17554 & w36783;
assign w35223 = ~w18175 & ~w7616;
assign w35224 = ~w18192 & ~w6764;
assign w35225 = ~w17591 & w36784;
assign w35226 = ~w18210 & ~w5965;
assign w35227 = w3803 & w36785;
assign w35228 = (~w33977 & w36786) | (~w33977 & w36787) | (w36786 & w36787);
assign w35229 = (w25156 & w36788) | (w25156 & w36789) | (w36788 & w36789);
assign w35230 = (~w25158 & w36790) | (~w25158 & w36791) | (w36790 & w36791);
assign w35231 = (w25170 & w25171) | (w25170 & ~w35192) | (w25171 & ~w35192);
assign w35232 = ~w18273 & w35199;
assign w35233 = (w35192 & w36792) | (w35192 & w36793) | (w36792 & w36793);
assign w35234 = (w25172 & w25173) | (w25172 & w35194) | (w25173 & w35194);
assign w35235 = (~w25156 & w36794) | (~w25156 & w36795) | (w36794 & w36795);
assign w35236 = (w25158 & w36796) | (w25158 & w36797) | (w36796 & w36797);
assign w35237 = ~w18280 & ~w1298;
assign w35238 = ~w18293 & ~w1697;
assign w35239 = w18028 & w18302;
assign w35240 = w18302 & w18258;
assign w35241 = w18258 & w35239;
assign w35242 = ~w18028 & ~w18302;
assign w35243 = ~w18302 & ~w18258;
assign w35244 = (~w18302 & ~w18258) | (~w18302 & w35242) | (~w18258 & w35242);
assign w35245 = ~w18306 & ~w2642;
assign w35246 = w18188 & w18201;
assign w35247 = ~w18323 & ~w9537;
assign w35248 = w18142 & w18129;
assign w35249 = w18142 & ~w31135;
assign w35250 = ~w18334 & ~w11623;
assign w35251 = w18352 & a_62;
assign w35252 = ~w18360 & ~w10565;
assign w35253 = w18109 & w18108;
assign w35254 = ~w18383 & ~w8529;
assign w35255 = ~w18400 & ~w7616;
assign w35256 = w18184 & w18409;
assign w35257 = ~w18399 & ~w31210;
assign w35258 = ~w18399 & ~w31209;
assign w35259 = w18399 & w31210;
assign w35260 = w18399 & w31209;
assign w35261 = ~w18414 & ~w6764;
assign w35262 = ~w18430 & ~w5965;
assign w35263 = ~w18447 & ~w5199;
assign w35264 = ~w18228 & w18085;
assign w35265 = w18075 & w18247;
assign w35266 = ~w18498 & ~w3198;
assign w35267 = ~w18520 & ~w2161;
assign w35268 = (~w33977 & w36798) | (~w33977 & w36799) | (w36798 & w36799);
assign w35269 = (w25156 & w36800) | (w25156 & w36801) | (w36800 & w36801);
assign w35270 = (~w25158 & w36802) | (~w25158 & w36803) | (w36802 & w36803);
assign w35271 = (w25175 & w25174) | (w25175 & ~w35192) | (w25174 & ~w35192);
assign w35272 = ~w18547 & w35236;
assign w35273 = (w35192 & w36804) | (w35192 & w36805) | (w36804 & w36805);
assign w35274 = (w25177 & w25176) | (w25177 & w35194) | (w25176 & w35194);
assign w35275 = (w25158 & w36808) | (w25158 & w36809) | (w36808 & w36809);
assign w35276 = (w25177 & w25176) | (w25177 & w35192) | (w25176 & w35192);
assign w35277 = ~w18554 & ~w1697;
assign w35278 = ~w18568 & ~w2161;
assign w35279 = ~w18581 & ~w2642;
assign w35280 = w18507 & ~w18497;
assign w35281 = w3195 & w36810;
assign w35282 = w18490 & w18604;
assign w35283 = ~w18490 & ~w18604;
assign w35284 = ~w18608 & ~w5199;
assign w35285 = ~w18620 & ~w5965;
assign w35286 = ~w18631 & ~w8529;
assign w35287 = ~w18642 & ~w10565;
assign w35288 = ~w18659 & ~w11623;
assign w35289 = ~w18658 & ~a_62;
assign w35290 = w18658 & a_62;
assign w35291 = ~w18681 & ~w9537;
assign w35292 = ~w18706 & ~w7616;
assign w35293 = w18399 & ~w31210;
assign w35294 = w18399 & ~w31209;
assign w35295 = ~w18725 & ~w6764;
assign w35296 = w4499 & w36811;
assign w35297 = ~w18772 & ~w3806;
assign w35298 = (w18801 & w29812) | (w18801 & w36812) | (w29812 & w36812);
assign w35299 = (w29747 & w36813) | (w29747 & w36814) | (w36813 & w36814);
assign w35300 = ~w1298 & a_20;
assign w35301 = w1298 & ~a_20;
assign w35302 = ~w18816 & ~w35275;
assign w35303 = (~w35192 & w36815) | (~w35192 & w36816) | (w36815 & w36816);
assign w35304 = (w25156 & w36817) | (w25156 & w36818) | (w36817 & w36818);
assign w35305 = (~w35194 & w36815) | (~w35194 & w36816) | (w36815 & w36816);
assign w35306 = ~w18815 & w35275;
assign w35307 = (w35192 & w36819) | (w35192 & w36820) | (w36819 & w36820);
assign w35308 = (~w25156 & w36821) | (~w25156 & w36822) | (w36821 & w36822);
assign w35309 = (w35194 & w36819) | (w35194 & w36820) | (w36819 & w36820);
assign w35310 = (~w18813 & w25178) | (~w18813 & w35275) | (w25178 & w35275);
assign w35311 = (w35192 & w36823) | (w35192 & w36824) | (w36823 & w36824);
assign w35312 = (~w25156 & w36825) | (~w25156 & w36826) | (w36825 & w36826);
assign w35313 = (w35194 & w36823) | (w35194 & w36824) | (w36823 & w36824);
assign w35314 = w18563 & ~w31298;
assign w35315 = ~w18831 & ~w1697;
assign w35316 = ~w18840 & ~w18577;
assign w35317 = w18317 & w35316;
assign w35318 = ~w18846 & ~w2161;
assign w35319 = w18590 & ~w31297;
assign w35320 = ~w18869 & ~w18604;
assign w35321 = w18480 & w36827;
assign w35322 = ~w18869 & ~w35320;
assign w35323 = (~w18869 & ~w18480) | (~w18869 & w36828) | (~w18480 & w36828);
assign w35324 = w3195 & w36829;
assign w35325 = w18768 & w18781;
assign w35326 = ~w18743 & w18617;
assign w35327 = ~w18889 & ~w5199;
assign w35328 = ~w18900 & ~w5965;
assign w35329 = ~w18911 & ~w6764;
assign w35330 = ~w18398 & w36830;
assign w35331 = ~w18922 & ~w7616;
assign w35332 = ~w18669 & w18651;
assign w35333 = ~w18934 & ~w10565;
assign w35334 = w18950 & w31351;
assign w35335 = w31350 & w36831;
assign w35336 = ~w18950 & ~w31351;
assign w35337 = (~w18950 & ~w31350) | (~w18950 & w36832) | (~w31350 & w36832);
assign w35338 = ~w18970 & ~w9537;
assign w35339 = w18641 & w18690;
assign w35340 = ~w18990 & ~w8529;
assign w35341 = w4499 & w36833;
assign w35342 = ~w19048 & ~w3806;
assign w35343 = (w25179 & w25180) | (w25179 & ~w35275) | (w25180 & ~w35275);
assign w35344 = (~w35192 & w36834) | (~w35192 & w36835) | (w36834 & w36835);
assign w35345 = (w25156 & w36836) | (w25156 & w36837) | (w36836 & w36837);
assign w35346 = (~w35194 & w36834) | (~w35194 & w36835) | (w36834 & w36835);
assign w35347 = ~w19084 & ~w1697;
assign w35348 = ~w19098 & ~w2161;
assign w35349 = ~w19113 & ~w2642;
assign w35350 = ~w19126 & ~w3198;
assign w35351 = w19044 & w19057;
assign w35352 = w18932 & w18931;
assign w35353 = ~w19151 & ~w11623;
assign w35354 = w19150 & a_62;
assign w35355 = ~w19170 & ~w10565;
assign w35356 = ~w19179 & ~w19165;
assign w35357 = ~w19188 & ~w9537;
assign w35358 = ~w18966 & w18979;
assign w35359 = (~w18969 & w36838) | (~w18969 & w36839) | (w36838 & w36839);
assign w35360 = (~w18969 & w31396) | (~w18969 & w36840) | (w31396 & w36840);
assign w35361 = (w18969 & w36841) | (w18969 & w36842) | (w36841 & w36842);
assign w35362 = ~w19204 & ~w8529;
assign w35363 = w18999 & w19213;
assign w35364 = ~w19220 & ~w7616;
assign w35365 = ~w19236 & ~w6764;
assign w35366 = ~w19253 & ~w5965;
assign w35367 = ~w19014 & w18909;
assign w35368 = w5196 & w36843;
assign w35369 = ~w19020 & w18898;
assign w35370 = w4499 & w36844;
assign w35371 = ~w19306 & ~w3806;
assign w35372 = (w25181 & w25182) | (w25181 & w35275) | (w25182 & w35275);
assign w35373 = (w35192 & w36845) | (w35192 & w36846) | (w36845 & w36846);
assign w35374 = (~w25156 & w36847) | (~w25156 & w36848) | (w36847 & w36848);
assign w35375 = (w35194 & w36845) | (w35194 & w36846) | (w36845 & w36846);
assign w35376 = (w25183 & w25184) | (w25183 & ~w35275) | (w25184 & ~w35275);
assign w35377 = (~w35192 & w36849) | (~w35192 & w36850) | (w36849 & w36850);
assign w35378 = (w25156 & w36851) | (w25156 & w36852) | (w36851 & w36852);
assign w35379 = (~w35194 & w36849) | (~w35194 & w36850) | (w36849 & w36850);
assign w35380 = (w19345 & w29812) | (w19345 & w36853) | (w29812 & w36853);
assign w35381 = (w29747 & w36854) | (w29747 & w36855) | (w36854 & w36855);
assign w35382 = ~w1697 & a_23;
assign w35383 = w1697 & ~a_23;
assign w35384 = ~w19353 & ~w2161;
assign w35385 = w19135 & w19321;
assign w35386 = ~w19381 & ~w3198;
assign w35387 = ~w19315 & w19390;
assign w35388 = w19315 & ~w19390;
assign w35389 = ~w19394 & ~w5965;
assign w35390 = ~w19405 & ~w6764;
assign w35391 = w19184 & w19179;
assign w35392 = w19184 & ~w31392;
assign w35393 = ~w19416 & ~w10565;
assign w35394 = w19432 & w31474;
assign w35395 = w19432 & w31475;
assign w35396 = ~w19432 & ~w31474;
assign w35397 = ~w19432 & ~w31475;
assign w35398 = ~w19452 & ~w9537;
assign w35399 = ~w19470 & ~w8529;
assign w35400 = ~w19489 & ~w7616;
assign w35401 = ~w19414 & ~w19415;
assign w35402 = w19414 & w19415;
assign w35403 = w5196 & w36856;
assign w35404 = ~w19535 & ~w4502;
assign w35405 = ~w19553 & ~w3806;
assign w35406 = (w25185 & w25186) | (w25185 & w35275) | (w25186 & w35275);
assign w35407 = (w35192 & w36857) | (w35192 & w36858) | (w36857 & w36858);
assign w35408 = (~w25156 & w36859) | (~w25156 & w36860) | (w36859 & w36860);
assign w35409 = (w35194 & w36857) | (w35194 & w36858) | (w36857 & w36858);
assign w35410 = (w25187 & w25188) | (w25187 & ~w35275) | (w25188 & ~w35275);
assign w35411 = (~w35192 & w36861) | (~w35192 & w36862) | (w36861 & w36862);
assign w35412 = (w25156 & w36863) | (w25156 & w36864) | (w36863 & w36864);
assign w35413 = (~w35194 & w36861) | (~w35194 & w36862) | (w36861 & w36862);
assign w35414 = (w33977 & w36865) | (w33977 & w36866) | (w36865 & w36866);
assign w35415 = (w25158 & w36869) | (w25158 & w36870) | (w36869 & w36870);
assign w35416 = (w27076 & w27075) | (w27076 & w35192) | (w27075 & w35192);
assign w35417 = ~w19597 & ~w2161;
assign w35418 = w19377 & ~w31508;
assign w35419 = ~w19611 & ~w2642;
assign w35420 = ~w19315 & ~w19390;
assign w35421 = ~w19620 & ~w19390;
assign w35422 = w19305 & w36871;
assign w35423 = ~w19620 & ~w35421;
assign w35424 = (~w19620 & ~w19305) | (~w19620 & w36872) | (~w19305 & w36872);
assign w35425 = w3195 & w36873;
assign w35426 = ~w19304 & w36874;
assign w35427 = ~w19640 & ~w3806;
assign w35428 = w19531 & w19544;
assign w35429 = ~w19251 & w36875;
assign w35430 = ~w19652 & ~w5965;
assign w35431 = ~w19463 & w36876;
assign w35432 = ~w19664 & ~w8529;
assign w35433 = w19681 & w31548;
assign w35434 = w31547 & w36877;
assign w35435 = ~w19681 & ~w31548;
assign w35436 = (~w19681 & ~w31547) | (~w19681 & w36878) | (~w31547 & w36878);
assign w35437 = ~w19695 & ~w10565;
assign w35438 = ~w19713 & ~w9537;
assign w35439 = ~w19735 & ~w7616;
assign w35440 = ~w19484 & w36879;
assign w35441 = ~w19754 & ~w6764;
assign w35442 = ~w19793 & ~w4502;
assign w35443 = ~w19831 & ~w35415;
assign w35444 = (~w35192 & w36880) | (~w35192 & w36881) | (w36880 & w36881);
assign w35445 = (w25156 & w36882) | (w25156 & w36883) | (w36882 & w36883);
assign w35446 = (~w33977 & w36884) | (~w33977 & w36885) | (w36884 & w36885);
assign w35447 = ~w19830 & w35415;
assign w35448 = (w35192 & w36886) | (w35192 & w36887) | (w36886 & w36887);
assign w35449 = (~w25156 & w36888) | (~w25156 & w36889) | (w36888 & w36889);
assign w35450 = (w33977 & w36890) | (w33977 & w36891) | (w36890 & w36891);
assign w35451 = ~w19838 & ~w2161;
assign w35452 = ~w19852 & ~w2642;
assign w35453 = ~w19865 & ~w3198;
assign w35454 = ~w19883 & ~w8529;
assign w35455 = ~w19904 & ~w11623;
assign w35456 = w19903 & a_62;
assign w35457 = ~w19921 & ~w10565;
assign w35458 = ~w19937 & ~w9537;
assign w35459 = ~w19725 & w19673;
assign w35460 = w7613 & w36892;
assign w35461 = ~w19731 & w19744;
assign w35462 = (~w19509 & w36893) | (~w19509 & w36894) | (w36893 & w36894);
assign w35463 = ~w20029 & ~w4502;
assign w35464 = ~w20046 & ~w3806;
assign w35465 = (w25192 & w25193) | (w25192 & ~w35415) | (w25193 & ~w35415);
assign w35466 = (~w35192 & w36895) | (~w35192 & w36896) | (w36895 & w36896);
assign w35467 = (w25156 & w36897) | (w25156 & w36898) | (w36897 & w36898);
assign w35468 = (~w33977 & w36899) | (~w33977 & w36900) | (w36899 & w36900);
assign w35469 = (w27077 & w27078) | (w27077 & w35275) | (w27078 & w35275);
assign w35470 = (w35192 & w36901) | (w35192 & w36902) | (w36901 & w36902);
assign w35471 = (~w25156 & w36903) | (~w25156 & w36904) | (w36903 & w36904);
assign w35472 = (w35194 & w36901) | (w35194 & w36902) | (w36901 & w36902);
assign w35473 = ~w20080 & ~w2642;
assign w35474 = w19874 & ~w20061;
assign w35475 = ~w20055 & ~w20103;
assign w35476 = w20055 & w20103;
assign w35477 = w7613 & w36905;
assign w35478 = w20135 & w31656;
assign w35479 = w20135 & w31657;
assign w35480 = ~w20135 & ~w31656;
assign w35481 = ~w20135 & ~w31657;
assign w35482 = ~w20149 & ~w10565;
assign w35483 = w19930 & w19893;
assign w35484 = ~w20167 & ~w9537;
assign w35485 = ~w20185 & ~w8529;
assign w35486 = ~w19991 & ~w19989;
assign w35487 = ~w20253 & ~w4502;
assign w35488 = ~w20269 & ~w3806;
assign w35489 = w20284 & ~w20089;
assign w35490 = (w20293 & w29812) | (w20293 & w36906) | (w29812 & w36906);
assign w35491 = (w29747 & w36907) | (w29747 & w36908) | (w36907 & w36908);
assign w35492 = ~w2161 & a_26;
assign w35493 = w2161 & ~a_26;
assign w35494 = (w25196 & w25197) | (w25196 & ~w35415) | (w25197 & ~w35415);
assign w35495 = (~w35192 & w36909) | (~w35192 & w36910) | (w36909 & w36910);
assign w35496 = (w25156 & w36911) | (w25156 & w36912) | (w36911 & w36912);
assign w35497 = (~w33977 & w36913) | (~w33977 & w36914) | (w36913 & w36914);
assign w35498 = (w27079 & w27080) | (w27079 & w35275) | (w27080 & w35275);
assign w35499 = (w35192 & w36915) | (w35192 & w36916) | (w36915 & w36916);
assign w35500 = (~w25156 & w36917) | (~w25156 & w36918) | (w36917 & w36918);
assign w35501 = (w35194 & w36915) | (w35194 & w36916) | (w36915 & w36916);
assign w35502 = (w25198 & w25199) | (w25198 & w35415) | (w25199 & w35415);
assign w35503 = (w35192 & w36919) | (w35192 & w36920) | (w36919 & w36920);
assign w35504 = (~w25156 & w36921) | (~w25156 & w36922) | (w36921 & w36922);
assign w35505 = (w33977 & w36923) | (w33977 & w36924) | (w36923 & w36924);
assign w35506 = ~w20089 & ~w20318;
assign w35507 = w20089 & ~w20318;
assign w35508 = ~w20321 & ~w2642;
assign w35509 = ~w20335 & ~w3198;
assign w35510 = ~w20350 & ~w3806;
assign w35511 = w20249 & w20262;
assign w35512 = ~w20361 & ~w4502;
assign w35513 = w20230 & w20244;
assign w35514 = w6761 & w36925;
assign w35515 = ~w20385 & ~w9537;
assign w35516 = ~w20396 & ~w10565;
assign w35517 = w20412 & w31732;
assign w35518 = w20412 & w31733;
assign w35519 = ~w20412 & ~w31732;
assign w35520 = ~w20412 & ~w31733;
assign w35521 = ~w20438 & ~w8529;
assign w35522 = w20181 & w20194;
assign w35523 = ~w20457 & ~w7616;
assign w35524 = w5196 & w36926;
assign w35525 = w31742 & w20504;
assign w35526 = ~w31742 & ~w20504;
assign w35527 = w31702 & w20529;
assign w35528 = ~w31702 & ~w20529;
assign w35529 = (w25156 & w36927) | (w25156 & w36928) | (w36927 & w36928);
assign w35530 = (~w33977 & w36929) | (~w33977 & w36930) | (w36929 & w36930);
assign w35531 = ~w20540 & ~w2642;
assign w35532 = ~w20330 & ~w20549;
assign w35533 = ~w35532 & ~w20549;
assign w35534 = ~w20553 & ~w3806;
assign w35535 = ~w20567 & ~w10565;
assign w35536 = ~w20593 & ~w11623;
assign w35537 = ~w20610 & ~w9537;
assign w35538 = ~w20627 & ~w8529;
assign w35539 = ~w20434 & w20447;
assign w35540 = w7613 & w36931;
assign w35541 = ~w20708 & ~w4502;
assign w35542 = w20717 & ~w27643;
assign w35543 = (w20717 & ~w27643) | (w20717 & w36932) | (~w27643 & w36932);
assign w35544 = ~w20717 & w27643;
assign w35545 = w27643 & w36933;
assign w35546 = ~w20732 & ~w3198;
assign w35547 = (w25202 & w25203) | (w25202 & w35415) | (w25203 & w35415);
assign w35548 = (w35192 & w36934) | (w35192 & w36935) | (w36934 & w36935);
assign w35549 = (~w25156 & w36936) | (~w25156 & w36937) | (w36936 & w36937);
assign w35550 = (w33977 & w36938) | (w33977 & w36939) | (w36938 & w36939);
assign w35551 = (w26932 & w26931) | (w26932 & ~w35275) | (w26931 & ~w35275);
assign w35552 = (~w35192 & w36940) | (~w35192 & w36941) | (w36940 & w36941);
assign w35553 = (w25156 & w36942) | (w25156 & w36943) | (w36942 & w36943);
assign w35554 = (~w35194 & w36940) | (~w35194 & w36941) | (w36940 & w36941);
assign w35555 = w20741 & ~w20731;
assign w35556 = (w20761 & w29812) | (w20761 & w36944) | (w29812 & w36944);
assign w35557 = (w29747 & w36945) | (w29747 & w36946) | (w36945 & w36946);
assign w35558 = ~w20770 & ~w3198;
assign w35559 = ~w20784 & ~w3806;
assign w35560 = w7613 & w36947;
assign w35561 = ~w20806 & ~w8529;
assign w35562 = ~w20817 & ~w10565;
assign w35563 = w11620 & w36948;
assign w35564 = ~w20833 & ~w31840;
assign w35565 = ~w20833 & ~w31839;
assign w35566 = w20833 & w31840;
assign w35567 = w20833 & w31839;
assign w35568 = ~w20857 & ~w9537;
assign w35569 = w5962 & w36949;
assign w35570 = ~w20924 & ~w5199;
assign w35571 = ~w20941 & ~w4502;
assign w35572 = (~w25156 & w36950) | (~w25156 & w36951) | (w36950 & w36951);
assign w35573 = (w35194 & w36952) | (w35194 & w36953) | (w36952 & w36953);
assign w35574 = w20766 & ~w31868;
assign w35575 = b_63 & w2642;
assign w35576 = w2642 & w34713;
assign w35577 = ~w34712 & w35575;
assign w35578 = ~w20986 & ~w3198;
assign w35579 = ~w20953 & w20793;
assign w35580 = (w20564 & w36954) | (w20564 & w36955) | (w36954 & w36955);
assign w35581 = ~w21002 & ~w4502;
assign w35582 = ~w21013 & ~w5199;
assign w35583 = ~w20642 & w36956;
assign w35584 = w7613 & w36957;
assign w35585 = ~w20844 & w20826;
assign w35586 = ~w21037 & ~w10565;
assign w35587 = w20829 & ~w21052;
assign w35588 = w35587 & ~w21051;
assign w35589 = ~w21057 & ~w11623;
assign w35590 = ~w21076 & ~w9537;
assign w35591 = ~w21095 & ~w8529;
assign w35592 = w5962 & w36958;
assign w35593 = w31916 & w21142;
assign w35594 = ~w31916 & ~w21142;
assign w35595 = ~w21022 & ~w21023;
assign w35596 = ~w21022 & ~w21145;
assign w35597 = w21022 & w21023;
assign w35598 = w21022 & w21145;
assign w35599 = ~w21160 & ~w3806;
assign w35600 = (w26934 & w26933) | (w26934 & w35415) | (w26933 & w35415);
assign w35601 = (w35192 & w36959) | (w35192 & w36960) | (w36959 & w36960);
assign w35602 = (~w25156 & w36961) | (~w25156 & w36962) | (w36961 & w36962);
assign w35603 = (w33977 & w36963) | (w33977 & w36964) | (w36963 & w36964);
assign w35604 = (w27083 & w27084) | (w27083 & w35275) | (w27084 & w35275);
assign w35605 = (w35192 & w36965) | (w35192 & w36966) | (w36965 & w36966);
assign w35606 = (~w25156 & w36967) | (~w25156 & w36968) | (w36967 & w36968);
assign w35607 = (w35194 & w36965) | (w35194 & w36966) | (w36965 & w36966);
assign w35608 = ~w21188 & ~w4502;
assign w35609 = w9534 & w36969;
assign w35610 = w21222 & ~w31901;
assign w35611 = ~w21229 & ~w11623;
assign w35612 = ~w21242 & ~w10565;
assign w35613 = ~w21331 & ~w5199;
assign w35614 = ~w21354 & ~w3806;
assign w35615 = ~w21156 & w21169;
assign w35616 = ~w21372 & ~w3198;
assign w35617 = ~w21370 & w21381;
assign w35618 = w21370 & ~w21381;
assign w35619 = (w21395 & w29812) | (w21395 & w36970) | (w29812 & w36970);
assign w35620 = (w29747 & w36971) | (w29747 & w36972) | (w36971 & w36972);
assign w35621 = ~w3198 & a_32;
assign w35622 = w3198 & ~a_32;
assign w35623 = w21363 & w21399;
assign w35624 = ~w21403 & ~w4502;
assign w35625 = w9534 & w36973;
assign w35626 = ~w21436 & ~w10565;
assign w35627 = w11620 & w36974;
assign w35628 = ~w21453 & ~w32011;
assign w35629 = ~w21453 & ~w32010;
assign w35630 = w21453 & w32011;
assign w35631 = w21453 & w32010;
assign w35632 = ~w21445 & w21464;
assign w35633 = w5962 & w36975;
assign w35634 = ~w21540 & ~w5199;
assign w35635 = (~w21199 & w36976) | (~w21199 & w36977) | (w36976 & w36977);
assign w35636 = (w21199 & w36978) | (w21199 & w36979) | (w36978 & w36979);
assign w35637 = ~w21564 & ~w3806;
assign w35638 = (w27085 & w27086) | (w27085 & w35275) | (w27086 & w35275);
assign w35639 = (w35192 & w36980) | (w35192 & w36981) | (w36980 & w36981);
assign w35640 = (~w25156 & w36982) | (~w25156 & w36983) | (w36982 & w36983);
assign w35641 = (w35194 & w36980) | (w35194 & w36981) | (w36980 & w36981);
assign w35642 = w5196 & w36984;
assign w35643 = w5962 & w36985;
assign w35644 = w9534 & w36986;
assign w35645 = w21449 & ~w21650;
assign w35646 = ~w21656 & ~w11623;
assign w35647 = ~w21670 & ~w10565;
assign w35648 = ~w21742 & ~w4502;
assign w35649 = ~w21552 & w21412;
assign w35650 = ~w21760 & ~w3806;
assign w35651 = (w26936 & w26935) | (w26936 & w35415) | (w26935 & w35415);
assign w35652 = (w35192 & w36987) | (w35192 & w36988) | (w36987 & w36988);
assign w35653 = (~w25156 & w36989) | (~w25156 & w36990) | (w36989 & w36990);
assign w35654 = (w33977 & w36991) | (w33977 & w36992) | (w36991 & w36992);
assign w35655 = (w26844 & w26843) | (w26844 & w35415) | (w26843 & w35415);
assign w35656 = (w35192 & w36993) | (w35192 & w36994) | (w36993 & w36994);
assign w35657 = (~w25156 & w36995) | (~w25156 & w36996) | (w36995 & w36996);
assign w35658 = (w33977 & w36997) | (w33977 & w36998) | (w36997 & w36998);
assign w35659 = ~w21785 & ~w5199;
assign w35660 = b_33 & ~a_32;
assign w35661 = ~b_33 & a_32;
assign w35662 = ~w21819 & ~w11623;
assign w35663 = w10562 & w36999;
assign w35664 = w5962 & w37000;
assign w35665 = ~w21927 & ~w4502;
assign w35666 = w21751 & ~w21738;
assign w35667 = w21751 & ~w21550;
assign w35668 = ~w21945 & ~w3806;
assign w35669 = ~w21943 & w21954;
assign w35670 = w21943 & ~w21954;
assign w35671 = (w21968 & w29812) | (w21968 & w37001) | (w29812 & w37001);
assign w35672 = (w29747 & w37002) | (w29747 & w37003) | (w37002 & w37003);
assign w35673 = ~w3806 & a_35;
assign w35674 = w3806 & ~a_35;
assign w35675 = w21936 & w21972;
assign w35676 = ~w21976 & ~w5199;
assign w35677 = w9534 & w37004;
assign w35678 = ~w21998 & ~w10565;
assign w35679 = ~w22016 & ~w32165;
assign w35680 = ~w22016 & ~w32164;
assign w35681 = w22016 & w32165;
assign w35682 = w22016 & w32164;
assign w35683 = w7613 & w37005;
assign w35684 = ~w22081 & ~w6764;
assign w35685 = ~w22098 & ~w5965;
assign w35686 = ~w22122 & ~w4502;
assign w35687 = (w26938 & w26937) | (w26938 & w35415) | (w26937 & w35415);
assign w35688 = (w35192 & w37006) | (w35192 & w37007) | (w37006 & w37007);
assign w35689 = (~w25156 & w37008) | (~w25156 & w37009) | (w37008 & w37009);
assign w35690 = (w33977 & w37010) | (w33977 & w37011) | (w37010 & w37011);
assign w35691 = (w26940 & w26939) | (w26940 & w35415) | (w26939 & w35415);
assign w35692 = (w35192 & w37012) | (w35192 & w37013) | (w37012 & w37013);
assign w35693 = (~w25156 & w37014) | (~w25156 & w37015) | (w37014 & w37015);
assign w35694 = (w33977 & w37016) | (w33977 & w37017) | (w37016 & w37017);
assign w35695 = (w32126 & w37018) | (w32126 & w37019) | (w37018 & w37019);
assign w35696 = ~w22160 & ~w5965;
assign w35697 = w22077 & w22090;
assign w35698 = ~w22171 & ~w6764;
assign w35699 = ~w22034 & w21996;
assign w35700 = w9534 & w37020;
assign w35701 = w22012 & ~w22199;
assign w35702 = w35701 & ~w22198;
assign w35703 = ~w22204 & ~w11623;
assign w35704 = ~w22218 & ~w10565;
assign w35705 = ~w21854 & w37021;
assign w35706 = ~w22254 & ~w7616;
assign w35707 = w32227 & w22263;
assign w35708 = ~w32227 & ~w22263;
assign w35709 = ~w22284 & ~w5199;
assign w35710 = ~w22302 & ~w4502;
assign w35711 = (w26942 & w26941) | (w26942 & w35415) | (w26941 & w35415);
assign w35712 = (w35192 & w37022) | (w35192 & w37023) | (w37022 & w37023);
assign w35713 = (~w25156 & w37024) | (~w25156 & w37025) | (w37024 & w37025);
assign w35714 = (w33977 & w37026) | (w33977 & w37027) | (w37026 & w37027);
assign w35715 = ~w22326 & ~w6764;
assign w35716 = ~w22349 & ~w11623;
assign w35717 = ~w22438 & ~w5965;
assign w35718 = ~w22455 & ~w5199;
assign w35719 = ~w22280 & w22293;
assign w35720 = ~w22473 & ~w4502;
assign w35721 = w22298 & w22311;
assign w35722 = (w22501 & w29812) | (w22501 & w37028) | (w29812 & w37028);
assign w35723 = (w29747 & w37029) | (w29747 & w37030) | (w37029 & w37030);
assign w35724 = ~w4502 & a_38;
assign w35725 = w4502 & ~a_38;
assign w35726 = (w32284 & w22526) | (w32284 & w37031) | (w22526 & w37031);
assign w35727 = (w32283 & w22526) | (w32283 & w37032) | (w22526 & w37032);
assign w35728 = w6761 & w37033;
assign w35729 = ~w22626 & ~w5965;
assign w35730 = ~w22643 & ~w5199;
assign w35731 = (w26944 & w26943) | (w26944 & w35415) | (w26943 & w35415);
assign w35732 = (w35192 & w37034) | (w35192 & w37035) | (w37034 & w37035);
assign w35733 = (~w25156 & w37036) | (~w25156 & w37037) | (w37036 & w37037);
assign w35734 = (w33977 & w37038) | (w33977 & w37039) | (w37038 & w37039);
assign w35735 = (w26946 & w26945) | (w26946 & w35415) | (w26945 & w35415);
assign w35736 = (w35192 & w37040) | (w35192 & w37041) | (w37040 & w37041);
assign w35737 = (~w25156 & w37042) | (~w25156 & w37043) | (w37042 & w37043);
assign w35738 = (w33977 & w37044) | (w33977 & w37045) | (w37044 & w37045);
assign w35739 = ~w22679 & ~w6764;
assign w35740 = (w22412 & w37046) | (w22412 & w37047) | (w37046 & w37047);
assign w35741 = ~w22690 & ~w7616;
assign w35742 = w22567 & w22580;
assign w35743 = ~w22713 & ~w11623;
assign w35744 = w22531 & w22545;
assign w35745 = ~w22377 & w37048;
assign w35746 = w8526 & w37049;
assign w35747 = ~w22788 & ~w5965;
assign w35748 = ~w22435 & w37050;
assign w35749 = ~w22806 & ~w5199;
assign w35750 = (w27087 & w27088) | (w27087 & w35275) | (w27088 & w35275);
assign w35751 = (w35192 & w37051) | (w35192 & w37052) | (w37051 & w37052);
assign w35752 = (~w25156 & w37053) | (~w25156 & w37054) | (w37053 & w37054);
assign w35753 = (w27087 & w27088) | (w27087 & w35274) | (w27088 & w35274);
assign w35754 = (~w22553 & w37055) | (~w22553 & w37056) | (w37055 & w37056);
assign w35755 = w22769 & ~w22755;
assign w35756 = ~w22853 & ~w11623;
assign w35757 = (~w22894 & w22876) | (~w22894 & w37057) | (w22876 & w37057);
assign w35758 = ~w22876 & w37058;
assign w35759 = (~w22535 & w37059) | (~w22535 & w37060) | (w37059 & w37060);
assign w35760 = w6761 & w37061;
assign w35761 = ~w22941 & ~w5965;
assign w35762 = ~w22784 & w22797;
assign w35763 = ~w22959 & ~w5199;
assign w35764 = (~w22625 & w37062) | (~w22625 & w37063) | (w37062 & w37063);
assign w35765 = (w22987 & w29812) | (w22987 & w37064) | (w29812 & w37064);
assign w35766 = (w29747 & w37065) | (w29747 & w37066) | (w37065 & w37066);
assign w35767 = ~w5199 & a_41;
assign w35768 = w5199 & ~a_41;
assign w35769 = w23003 & w32401;
assign w35770 = w23003 & w32402;
assign w35771 = ~w23003 & ~w32401;
assign w35772 = ~w23003 & ~w32402;
assign w35773 = ~w23072 & ~w7616;
assign w35774 = ~w23090 & ~w6764;
assign w35775 = ~w23107 & ~w5965;
assign w35776 = ~w23142 & ~w6764;
assign w35777 = ~w23152 & ~w7616;
assign w35778 = ~w23163 & ~w8529;
assign w35779 = w23030 & w23044;
assign w35780 = ~w23014 & w23027;
assign w35781 = ~w23186 & ~w11623;
assign w35782 = ~w23215 & ~w9537;
assign w35783 = ~w22921 & w37067;
assign w35784 = ~w23253 & ~w5965;
assign w35785 = ~w23276 & ~w6764;
assign w35786 = ~w23287 & ~w7616;
assign w35787 = w9534 & w37068;
assign w35788 = ~w23362 & ~w8529;
assign w35789 = ~w23392 & ~w5965;
assign w35790 = (w23420 & w29812) | (w23420 & w37069) | (w29812 & w37069);
assign w35791 = (w29747 & w37070) | (w29747 & w37071) | (w37070 & w37071);
assign w35792 = ~w5965 & a_44;
assign w35793 = w5965 & ~a_44;
assign w35794 = ~w23428 & ~w6764;
assign w35795 = (w32495 & w23447) | (w32495 & w37072) | (w23447 & w37072);
assign w35796 = (w32496 & w23447) | (w32496 & w37073) | (w23447 & w37073);
assign w35797 = ~w23447 & w37074;
assign w35798 = ~w23447 & w37075;
assign w35799 = w10562 & w37076;
assign w35800 = ~w23481 & ~w9537;
assign w35801 = ~w23499 & ~w8529;
assign w35802 = ~w23516 & ~w7616;
assign w35803 = ~w23437 & ~w23555;
assign w35804 = ~w23560 & ~w7616;
assign w35805 = ~w23571 & ~w8529;
assign w35806 = ~w23582 & ~w9537;
assign w35807 = w10562 & w37077;
assign w35808 = w23439 & w23525;
assign w35809 = ~w23657 & ~w6764;
assign w35810 = ~w23680 & ~w6764;
assign w35811 = ~w23691 & ~w7616;
assign w35812 = ~w23702 & ~w8529;
assign w35813 = ~w23713 & ~w9537;
assign w35814 = w11620 & w37078;
assign w35815 = w10562 & w37079;
assign w35816 = (w23804 & w29812) | (w23804 & w37080) | (w29812 & w37080);
assign w35817 = (w29747 & w37081) | (w29747 & w37082) | (w37081 & w37082);
assign w35818 = ~w6764 & a_47;
assign w35819 = w6764 & ~a_47;
assign w35820 = w23700 & w23808;
assign w35821 = ~w23812 & ~w7616;
assign w35822 = ~w23824 & ~w9537;
assign w35823 = w10562 & w37083;
assign w35824 = ~w23852 & ~w25710;
assign w35825 = ~w23852 & ~w25711;
assign w35826 = ~w23882 & ~w8529;
assign w35827 = ~w23789 & ~w23787;
assign w35828 = (w26948 & w26947) | (w26948 & ~w35415) | (w26947 & ~w35415);
assign w35829 = (~w35192 & w37084) | (~w35192 & w37085) | (w37084 & w37085);
assign w35830 = (w25156 & w37086) | (w25156 & w37087) | (w37086 & w37087);
assign w35831 = (w26948 & w26947) | (w26948 & ~w35414) | (w26947 & ~w35414);
assign w35832 = ~w23914 & ~w8529;
assign w35833 = w9534 & w37088;
assign w35834 = ~w23936 & ~w10565;
assign w35835 = ~w23956 & ~w11623;
assign w35836 = ~w23993 & ~w7616;
assign w35837 = ~b_63 & ~w24007;
assign w35838 = ~w24007 & ~w34713;
assign w35839 = ~w24007 & ~w34714;
assign w35840 = (~w24011 & w23820) | (~w24011 & w37089) | (w23820 & w37089);
assign w35841 = ~w23820 & w37090;
assign w35842 = ~w24026 & ~w7616;
assign w35843 = w23924 & w23923;
assign w35844 = ~w24037 & ~w8529;
assign w35845 = ~w24048 & ~w9537;
assign w35846 = ~w11623 & a_62;
assign w35847 = w24078 & w32643;
assign w35848 = w24078 & w32642;
assign w35849 = ~w24086 & ~w10565;
assign w35850 = ~w29812 & w37091;
assign w35851 = (~w29747 & w37092) | (~w29747 & w37093) | (w37092 & w37093);
assign w35852 = ~w24139 & ~w8529;
assign w35853 = ~w24150 & ~w9537;
assign w35854 = ~w24161 & ~w10565;
assign w35855 = w24179 & w32666;
assign w35856 = w24179 & w32667;
assign w35857 = ~w24179 & ~w32666;
assign w35858 = ~w24179 & ~w32667;
assign w35859 = ~w24170 & w24190;
assign w35860 = ~w24116 & ~w24114;
assign w35861 = ~w24226 & ~w9537;
assign w35862 = ~w24262 & ~w10565;
assign w35863 = ~w24197 & w24159;
assign w35864 = ~w24286 & ~w8529;
assign w35865 = ~b_63 & ~w24300;
assign w35866 = ~w24300 & ~w34713;
assign w35867 = ~w24300 & ~w34714;
assign w35868 = ~w7616 & a_50;
assign w35869 = w7616 & ~a_50;
assign w35870 = (~w24304 & w24147) | (~w24304 & w37094) | (w24147 & w37094);
assign w35871 = ~w24147 & w37095;
assign w35872 = ~w24274 & w24235;
assign w35873 = ~w24320 & ~w9537;
assign w35874 = w10562 & w37096;
assign w35875 = w11620 & w37097;
assign w35876 = ~w24380 & ~w8529;
assign w35877 = (~w24200 & w37098) | (~w24200 & w37099) | (w37098 & w37099);
assign w35878 = ~w29812 & w37100;
assign w35879 = (~w29747 & w37101) | (~w29747 & w37102) | (w37101 & w37102);
assign w35880 = ~w24414 & ~w9537;
assign w35881 = ~w24425 & ~w10565;
assign w35882 = ~w24441 & ~w26493;
assign w35883 = ~w24441 & ~w26492;
assign w35884 = w33949 & ~w24485;
assign w35885 = ~w24491 & ~w11623;
assign w35886 = ~w24504 & ~w10565;
assign w35887 = ~w24520 & ~w9537;
assign w35888 = ~b_63 & ~w24534;
assign w35889 = ~w24534 & ~w34713;
assign w35890 = ~w24534 & ~w34714;
assign w35891 = ~w8529 & a_53;
assign w35892 = w8529 & ~a_53;
assign w35893 = ~w24458 & w24538;
assign w35894 = ~w24555 & ~w9537;
assign w35895 = ~w24570 & ~w10565;
assign w35896 = w24588 & w32764;
assign w35897 = w24588 & w32763;
assign w35898 = ~w29812 & w37103;
assign w35899 = (~w29747 & w37104) | (~w29747 & w37105) | (w37104 & w37105);
assign w35900 = ~w24633 & ~w10565;
assign w35901 = w24651 & w32781;
assign w35902 = w24651 & w32782;
assign w35903 = ~w24651 & ~w32781;
assign w35904 = ~w24651 & ~w32782;
assign w35905 = ~w24642 & w24662;
assign w35906 = w24690 & w29583;
assign w35907 = w24690 & w29582;
assign w35908 = (a_62 & w27711) | (a_62 & ~w29583) | (w27711 & ~w29583);
assign w35909 = (a_62 & w27711) | (a_62 & ~w29582) | (w27711 & ~w29582);
assign w35910 = ~w24710 & ~w10565;
assign w35911 = ~b_63 & ~w24724;
assign w35912 = ~w24724 & ~w34713;
assign w35913 = ~w24724 & ~w34714;
assign w35914 = ~w9537 & a_56;
assign w35915 = w9537 & ~a_56;
assign w35916 = ~w24662 & w24728;
assign w35917 = ~w24669 & w24631;
assign w35918 = w24719 & w24706;
assign w35919 = w24719 & ~w24704;
assign w35920 = ~w24744 & ~w10565;
assign w35921 = ~w24772 & ~w11623;
assign w35922 = ~w24783 & ~w24753;
assign w35923 = w24801 & w32830;
assign w35924 = w24801 & w32831;
assign w35925 = ~w24801 & ~w32830;
assign w35926 = ~w24801 & ~w32831;
assign w35927 = ~w29812 & w37106;
assign w35928 = (~w29747 & w37107) | (~w29747 & w37108) | (w37107 & w37108);
assign w35929 = w24753 & w24782;
assign w35930 = ~w24812 & w24824;
assign w35931 = ~w24842 & w24798;
assign w35932 = ~w24842 & w32826;
assign w35933 = w24841 & ~w24842;
assign w35934 = ~w24841 & w35933;
assign w35935 = ~w24848 & ~w11623;
assign w35936 = ~w24888 & ~w11623;
assign w35937 = w24887 & a_62;
assign w35938 = (w24923 & w29812) | (w24923 & w37109) | (w29812 & w37109);
assign w35939 = w24923 & ~w29823;
assign w35940 = w11623 & ~a_62;
assign w35941 = ~b_63 & ~w24946;
assign w35942 = ~w24946 & ~w34713;
assign w35943 = ~w24946 & ~w34714;
assign w35944 = ~w11623 & a_62;
assign w35945 = (w26500 & w26501) | (w26500 & ~w33681) | (w26501 & ~w33681);
assign w35946 = (w26500 & w26501) | (w26500 & ~w33680) | (w26501 & ~w33680);
assign w35947 = (w33612 & w37110) | (w33612 & w37111) | (w37110 & w37111);
assign w35948 = (w26500 & w26501) | (w26500 & ~w33683) | (w26501 & ~w33683);
assign w35949 = (w26502 & w26503) | (w26502 & ~w33681) | (w26503 & ~w33681);
assign w35950 = (w26502 & w26503) | (w26502 & ~w33680) | (w26503 & ~w33680);
assign w35951 = (w33612 & w37112) | (w33612 & w37113) | (w37112 & w37113);
assign w35952 = (w26502 & w26503) | (w26502 & ~w33683) | (w26503 & ~w33683);
assign w35953 = (w26504 & w26505) | (w26504 & ~w33681) | (w26505 & ~w33681);
assign w35954 = (w26504 & w26505) | (w26504 & ~w33680) | (w26505 & ~w33680);
assign w35955 = (w33612 & w37114) | (w33612 & w37115) | (w37114 & w37115);
assign w35956 = (w26504 & w26505) | (w26504 & ~w33683) | (w26505 & ~w33683);
assign w35957 = (w26506 & w26507) | (w26506 & w33681) | (w26507 & w33681);
assign w35958 = (w26506 & w26507) | (w26506 & w33680) | (w26507 & w33680);
assign w35959 = (~w33612 & w37116) | (~w33612 & w37117) | (w37116 & w37117);
assign w35960 = (w26506 & w26507) | (w26506 & w33683) | (w26507 & w33683);
assign w35961 = ~w3726 & ~w3949;
assign w35962 = ~w8775 & ~w9094;
assign w35963 = w16802 & ~w17121;
assign w35964 = w17121 & ~w17118;
assign w35965 = (~w17118 & w25479) | (~w17118 & ~w16802) | (w25479 & ~w16802);
assign w35966 = ~w17711 & ~w17710;
assign w35967 = (~w17710 & ~w17711) | (~w17710 & ~w17415) | (~w17711 & ~w17415);
assign w35968 = ~w18273 & ~w18271;
assign w35969 = ~w19582 & ~w19581;
assign w35970 = w21387 & ~w21584;
assign w35971 = ~w21581 & ~w35970;
assign w35972 = (~w21780 & w26974) | (~w21780 & ~w21584) | (w26974 & ~w21584);
assign w35973 = (~w21780 & w26974) | (~w21780 & w35970) | (w26974 & w35970);
assign w35974 = w33740 & w37118;
assign w35975 = ~w22141 & ~w22140;
assign w35976 = ~w22319 & ~w22321;
assign w35977 = ~w22141 & ~w22319;
assign w35978 = w26509 & w22494;
assign w35979 = (w22494 & w26509) | (w22494 & w22321) | (w26509 & w22321);
assign w35980 = w26509 | w22494;
assign w35981 = (w22494 & w26509) | (w22494 & w22141) | (w26509 & w22141);
assign w35982 = (w22140 & w35978) | (w22140 & w35979) | (w35978 & w35979);
assign w35983 = (w26744 & w26745) | (w26744 & ~w22321) | (w26745 & ~w22321);
assign w35984 = w26745 | w26744;
assign w35985 = w26745 & w26744;
assign w35986 = (w26744 & w26745) | (w26744 & ~w22141) | (w26745 & ~w22141);
assign w35987 = ~w23411 & ~w25489;
assign w35988 = ~w23269 & w37119;
assign w35989 = (w23544 & w23413) | (w23544 & w26084) | (w23413 & w26084);
assign w35990 = (w23544 & w26084) | (w23544 & w23413) | (w26084 & w23413);
assign w35991 = (w23544 & w26084) | (w23544 & w25489) | (w26084 & w25489);
assign w35992 = (w26510 & w26511) | (w26510 & ~w23413) | (w26511 & ~w23413);
assign w35993 = (w26510 & w26511) | (w26510 & ~w25489) | (w26511 & ~w25489);
assign w35994 = (~w23543 & w26510) | (~w23543 & ~w23270) | (w26510 & ~w23270);
assign w35995 = (~w23413 & w37120) | (~w23413 & w26511) | (w37120 & w26511);
assign w35996 = (w26746 & w26747) | (w26746 & w23411) | (w26747 & w23411);
assign w35997 = (w26746 & w26747) | (w26746 & w23270) | (w26747 & w23270);
assign w35998 = (w23413 & w37121) | (w23413 & w35996) | (w37121 & w35996);
assign w35999 = (w23676 & w23544) | (w23676 & w26746) | (w23544 & w26746);
assign w36000 = w23676 & ~w26511;
assign w36001 = (~w23674 & w26748) | (~w23674 & w26510) | (w26748 & w26510);
assign w36002 = (~w23674 & w26748) | (~w23674 & w26511) | (w26748 & w26511);
assign w36003 = (w26872 & w26873) | (w26872 & ~w26510) | (w26873 & ~w26510);
assign w36004 = (w26872 & w26873) | (w26872 & ~w26511) | (w26873 & ~w26511);
assign w36005 = ~w23795 & w33741;
assign w36006 = (w24400 & w24315) | (w24400 & w37122) | (w24315 & w37122);
assign w36007 = w24400 & ~w26750;
assign w36008 = (~w24315 & w37123) | (~w24315 & w37124) | (w37123 & w37124);
assign w36009 = (~w24399 & w26874) | (~w24399 & w26750) | (w26874 & w26750);
assign w36010 = (w24315 & w37125) | (w24315 & w37126) | (w37125 & w37126);
assign w36011 = (w26981 & w26982) | (w26981 & ~w26750) | (w26982 & ~w26750);
assign w36012 = w24738 & w24791;
assign w36013 = ~w24874 & w24790;
assign w36014 = (~w24874 & w24832) | (~w24874 & w33056) | (w24832 & w33056);
assign w36015 = w24874 & ~w24871;
assign w36016 = w24871 & ~w24908;
assign w36017 = w24908 & ~w24905;
assign w36018 = (~w24905 & w24908) | (~w24905 & w37127) | (w24908 & w37127);
assign w36019 = ~w24935 & w24905;
assign w36020 = (~w24935 & ~w24908) | (~w24935 & w36019) | (~w24908 & w36019);
assign w36021 = ~w24935 & ~w36018;
assign w36022 = w24953 & w24972;
assign w36023 = b_41 & a_11;
assign w36024 = b_39 & a_14;
assign w36025 = b_42 & a_11;
assign w36026 = b_40 & a_14;
assign w36027 = b_41 & a_14;
assign w36028 = b_42 & a_14;
assign w36029 = b_43 & a_14;
assign w36030 = b_44 & a_14;
assign w36031 = b_47 & a_11;
assign w36032 = ~w24932 & ~w36019;
assign w36033 = (w24908 & w37128) | (w24908 & w36032) | (w37128 & w36032);
assign w36034 = (~w24932 & w36018) | (~w24932 & w37128) | (w36018 & w37128);
assign w36035 = ~w24954 | w25328;
assign w36036 = (w25328 & w25329) | (w25328 & ~w36019) | (w25329 & ~w36019);
assign w36037 = (w24908 & w33141) | (w24908 & w36036) | (w33141 & w36036);
assign w36038 = (w36018 & w37129) | (w36018 & w33141) | (w37129 & w33141);
assign w36039 = (w25332 & w25333) | (w25332 & ~w36019) | (w25333 & ~w36019);
assign w36040 = (w24908 & w33144) | (w24908 & w36039) | (w33144 & w36039);
assign w36041 = (w36018 & w37130) | (w36018 & w33144) | (w37130 & w33144);
assign w36042 = ~w33078 & a_26;
assign w36043 = b_38 & a_17;
assign w36044 = ~b_41 & a_14;
assign w36045 = b_39 & a_17;
assign w36046 = b_40 & a_17;
assign w36047 = b_46 & a_11;
assign w36048 = b_41 & a_17;
assign w36049 = b_48 & a_11;
assign w36050 = b_45 & a_14;
assign w36051 = b_39 & a_20;
assign w36052 = b_40 & a_20;
assign w36053 = b_41 & a_20;
assign w36054 = b_47 & a_14;
assign w36055 = b_40 & a_23;
assign w36056 = b_47 & a_17;
assign w36057 = b_45 & a_20;
assign w36058 = b_40 & a_26;
assign w36059 = b_49 & a_26;
assign w36060 = ~w15830 & w15535;
assign w36061 = b_47 & a_50;
assign w36062 = b_45 & a_53;
assign w36063 = b_48 & a_50;
assign w36064 = b_42 & a_59;
assign w36065 = b_45 & a_56;
assign w36066 = b_48 & a_53;
assign w36067 = b_46 & a_56;
assign w36068 = b_49 & a_53;
assign w36069 = b_45 & a_59;
assign w36070 = b_49 & a_62;
assign w36071 = ~b_49 & a_62;
assign w36072 = (~w24957 & w25327) | (~w24957 & w36019) | (w25327 & w36019);
assign w36073 = (~w24908 & w33244) | (~w24908 & w36072) | (w33244 & w36072);
assign w36074 = (~w36018 & w33243) | (~w36018 & w33244) | (w33243 & w33244);
assign w36075 = (w25330 & w25331) | (w25330 & w36019) | (w25331 & w36019);
assign w36076 = (~w24908 & w33248) | (~w24908 & w36075) | (w33248 & w36075);
assign w36077 = (~w36018 & w33247) | (~w36018 & w33248) | (w33247 & w33248);
assign w36078 = ~w33252 & a_29;
assign w36079 = b_38 & a_20;
assign w36080 = b_33 & a_26;
assign w36081 = b_42 & a_17;
assign w36082 = b_49 & a_11;
assign w36083 = b_37 & a_23;
assign w36084 = b_43 & a_17;
assign w36085 = b_46 & a_14;
assign w36086 = b_38 & a_23;
assign w36087 = b_44 & a_17;
assign w36088 = b_48 & a_14;
assign w36089 = b_45 & a_17;
assign w36090 = b_33 & a_29;
assign w36091 = b_39 & a_23;
assign w36092 = b_42 & a_20;
assign w36093 = b_31 & a_32;
assign w36094 = b_37 & a_26;
assign w36095 = b_41 & a_23;
assign w36096 = b_44 & a_20;
assign w36097 = ~b_47 & a_17;
assign w36098 = b_48 & a_17;
assign w36099 = b_42 & a_23;
assign w36100 = b_33 & a_32;
assign w36101 = b_39 & a_26;
assign w36102 = b_49 & a_17;
assign w36103 = b_46 & a_20;
assign w36104 = b_37 & a_29;
assign w36105 = b_47 & a_20;
assign w36106 = b_52 & a_17;
assign w36107 = b_56 & a_14;
assign w36108 = (w13803 & w37131) | (w13803 & ~w14034) | (w37131 & ~w14034);
assign w36109 = b_49 & a_23;
assign w36110 = b_41 & a_32;
assign w36111 = b_47 & a_29;
assign w36112 = b_52 & a_29;
assign w36113 = b_47 & a_44;
assign w36114 = b_48 & a_44;
assign w36115 = b_47 & a_47;
assign w36116 = b_48 & a_47;
assign w36117 = b_42 & a_56;
assign w36118 = b_51 & a_47;
assign w36119 = b_37 & a_62;
assign w36120 = b_40 & a_62;
assign w36121 = b_43 & a_59;
assign w36122 = b_52 & a_50;
assign w36123 = b_47 & a_56;
assign w36124 = b_48 & a_56;
assign w36125 = b_46 & a_59;
assign w36126 = b_49 & a_56;
assign w36127 = b_55 & a_62;
assign w36128 = (w25296 & w25297) | (w25296 & w36005) | (w25297 & w36005);
assign w36129 = ~w33372 & a_14;
assign w36130 = ~w33373 & a_17;
assign w36131 = ~w33374 & a_20;
assign w36132 = ~w33375 & a_23;
assign w36133 = b_5 & a_26;
assign w36134 = b_5 & a_47;
assign w36135 = ~w33376 & a_50;
assign w36136 = b_5 & a_50;
assign w36137 = ~w33377 & a_53;
assign w36138 = b_5 & a_53;
assign w36139 = b_28 & a_32;
assign w36140 = b_34 & a_26;
assign w36141 = b_50 & a_11;
assign w36142 = b_35 & a_26;
assign w36143 = b_17 & a_44;
assign w36144 = b_29 & a_32;
assign w36145 = b_51 & a_11;
assign w36146 = b_18 & a_44;
assign w36147 = b_27 & a_35;
assign w36148 = b_36 & a_26;
assign w36149 = b_49 & a_14;
assign w36150 = b_28 & a_35;
assign w36151 = b_43 & a_20;
assign w36152 = b_46 & a_17;
assign w36153 = b_50 & a_14;
assign w36154 = b_29 & a_35;
assign w36155 = b_32 & a_32;
assign w36156 = b_38 & a_26;
assign w36157 = b_30 & a_35;
assign w36158 = b_31 & a_35;
assign w36159 = b_41 & a_26;
assign w36160 = b_44 & a_23;
assign w36161 = b_49 & a_20;
assign w36162 = b_50 & a_20;
assign w36163 = b_47 & a_23;
assign w36164 = b_56 & a_17;
assign w36165 = b_47 & a_26;
assign w36166 = b_45 & a_29;
assign w36167 = b_56 & a_20;
assign w36168 = w16249 & ~w15916;
assign w36169 = w15778 & w37132;
assign w36170 = b_48 & a_32;
assign w36171 = b_49 & a_32;
assign w36172 = b_53 & a_29;
assign w36173 = b_56 & a_29;
assign w36174 = b_45 & a_47;
assign w36175 = b_51 & a_41;
assign w36176 = w21142 & w21126;
assign w36177 = (w21142 & w20884) | (w21142 & w37133) | (w20884 & w37133);
assign w36178 = b_45 & a_50;
assign w36179 = b_51 & a_44;
assign w36180 = b_46 & a_50;
assign w36181 = b_49 & a_47;
assign w36182 = b_44 & a_53;
assign w36183 = b_50 & a_47;
assign w36184 = b_47 & a_53;
assign w36185 = b_51 & a_50;
assign w36186 = b_54 & a_50;
assign w36187 = b_51 & a_53;
assign w36188 = b_52 & a_53;
assign w36189 = ~w23052 & ~w23081;
assign w36190 = b_53 & a_62;
assign w36191 = (~w25292 & w37134) | (~w25292 & w37135) | (w37134 & w37135);
assign w36192 = (w25287 & w37136) | (w25287 & w37137) | (w37136 & w37137);
assign w36193 = ~w24548 & ~w26980;
assign w36194 = ~w24548 & ~w23910;
assign w36195 = (~w25292 & w37138) | (~w25292 & w37139) | (w37138 & w37139);
assign w36196 = (w25287 & w37140) | (w25287 & w37141) | (w37140 & w37141);
assign w36197 = (w25299 & w25300) | (w25299 & ~w26980) | (w25300 & ~w26980);
assign w36198 = (w25299 & w25300) | (w25299 & ~w23910) | (w25300 & ~w23910);
assign w36199 = (~w25292 & w37142) | (~w25292 & w37143) | (w37142 & w37143);
assign w36200 = (w25287 & w37144) | (w25287 & w37145) | (w37144 & w37145);
assign w36201 = (w25304 & w25303) | (w25304 & ~w26980) | (w25303 & ~w26980);
assign w36202 = (w25304 & w25303) | (w25304 & ~w23910) | (w25303 & ~w23910);
assign w36203 = (~w25292 & w37146) | (~w25292 & w37147) | (w37146 & w37147);
assign w36204 = (w25287 & w37148) | (w25287 & w37149) | (w37148 & w37149);
assign w36205 = (w25308 & w25307) | (w25308 & ~w26980) | (w25307 & ~w26980);
assign w36206 = (w25308 & w25307) | (w25308 & ~w23910) | (w25307 & ~w23910);
assign w36207 = (~w25292 & w37150) | (~w25292 & w37151) | (w37150 & w37151);
assign w36208 = (w25287 & w37152) | (w25287 & w37153) | (w37152 & w37153);
assign w36209 = (w25311 & w25312) | (w25311 & ~w26980) | (w25312 & ~w26980);
assign w36210 = (w25311 & w25312) | (w25311 & ~w23910) | (w25312 & ~w23910);
assign w36211 = (w25328 & w37154) | (w25328 & w37155) | (w37154 & w37155);
assign w36212 = (~w25328 & w37156) | (~w25328 & w37157) | (w37156 & w37157);
assign w36213 = ~w33543 & a_11;
assign w36214 = b_5 & a_29;
assign w36215 = ~w33544 & a_32;
assign w36216 = ~w33545 & a_35;
assign w36217 = b_5 & a_35;
assign w36218 = ~w33546 & a_38;
assign w36219 = b_5 & a_38;
assign w36220 = ~w33547 & a_41;
assign w36221 = b_5 & a_41;
assign w36222 = b_39 & a_11;
assign w36223 = b_40 & a_11;
assign w36224 = b_45 & a_8;
assign w36225 = b_33 & a_20;
assign w36226 = b_37 & a_17;
assign w36227 = b_43 & a_11;
assign w36228 = b_46 & a_8;
assign w36229 = b_47 & a_8;
assign w36230 = b_33 & a_23;
assign w36231 = b_37 & a_20;
assign w36232 = b_35 & a_23;
assign w36233 = b_32 & a_26;
assign w36234 = b_46 & a_23;
assign w36235 = b_48 & a_41;
assign w36236 = b_46 & a_44;
assign w36237 = b_42 & a_53;
assign w36238 = b_43 & a_53;
assign w36239 = ~w21898 & w21709;
assign w36240 = ~w21898 & ~w21710;
assign w36241 = b_45 & a_62;
assign w36242 = b_48 & a_59;
assign w36243 = (~w25263 & w37158) | (~w25263 & w37159) | (w37158 & w37159);
assign w36244 = (~w25268 & w37160) | (~w25268 & w37161) | (w37160 & w37161);
assign w36245 = (~w25263 & w37162) | (~w25263 & w37163) | (w37162 & w37163);
assign w36246 = (~w25268 & w37164) | (~w25268 & w37165) | (w37164 & w37165);
assign w36247 = (~w25263 & w37166) | (~w25263 & w37167) | (w37166 & w37167);
assign w36248 = (~w25268 & w37168) | (~w25268 & w37169) | (w37168 & w37169);
assign w36249 = (~w25263 & w37170) | (~w25263 & w37171) | (w37170 & w37171);
assign w36250 = (~w25268 & w37172) | (~w25268 & w37173) | (w37172 & w37173);
assign w36251 = (~w25263 & w37174) | (~w25263 & w37175) | (w37174 & w37175);
assign w36252 = (~w25268 & w37176) | (~w25268 & w37177) | (w37176 & w37177);
assign w36253 = (~w25263 & w37178) | (~w25263 & w37179) | (w37178 & w37179);
assign w36254 = (~w25268 & w37180) | (~w25268 & w37181) | (w37180 & w37181);
assign w36255 = (~w25263 & w37182) | (~w25263 & w37183) | (w37182 & w37183);
assign w36256 = (~w25268 & w37184) | (~w25268 & w37185) | (w37184 & w37185);
assign w36257 = (w25292 & w37186) | (w25292 & w37187) | (w37186 & w37187);
assign w36258 = (~w25287 & w37188) | (~w25287 & w37189) | (w37188 & w37189);
assign w36259 = (w25325 & w25326) | (w25325 & w26980) | (w25326 & w26980);
assign w36260 = (w25325 & w25326) | (w25325 & w23910) | (w25326 & w23910);
assign w36261 = b_5 & a_8;
assign w36262 = b_5 & a_14;
assign w36263 = b_5 & a_17;
assign w36264 = b_5 & a_20;
assign w36265 = b_5 & a_44;
assign w36266 = b_5 & a_56;
assign w36267 = (~w11526 & w37190) | (~w11526 & w37191) | (w37190 & w37191);
assign w36268 = (w11906 & ~w11526) | (w11906 & w37192) | (~w11526 & w37192);
assign w36269 = (w11526 & w37193) | (w11526 & w37194) | (w37193 & w37194);
assign w36270 = w11526 & w37195;
assign w36271 = w13007 & w13389;
assign w36272 = ~w13007 & ~w13389;
assign w36273 = (w25207 & w25208) | (w25207 & ~w26972) | (w25208 & ~w26972);
assign w36274 = (w25207 & w25208) | (w25207 & ~w20305) | (w25208 & ~w20305);
assign w36275 = (w25207 & w25208) | (w25207 & ~w20754) | (w25208 & ~w20754);
assign w36276 = (w25219 & w25220) | (w25219 & ~w26972) | (w25220 & ~w26972);
assign w36277 = (w25223 & w25224) | (w25223 & ~w26972) | (w25224 & ~w26972);
assign w36278 = (~w22978 & w25246) | (~w22978 & ~w21777) | (w25246 & ~w21777);
assign w36279 = (w25237 & w37196) | (w25237 & w37197) | (w37196 & w37197);
assign w36280 = ~w22980 & ~w22978;
assign w36281 = (w25236 & w37196) | (w25236 & w37197) | (w37196 & w37197);
assign w36282 = (w25250 & w25249) | (w25250 & ~w21777) | (w25249 & ~w21777);
assign w36283 = (w25237 & w37198) | (w25237 & w37199) | (w37198 & w37199);
assign w36284 = ~w25248 & w37200;
assign w36285 = (w25236 & w37198) | (w25236 & w37199) | (w37198 & w37199);
assign w36286 = (w25254 & w25253) | (w25254 & ~w21777) | (w25253 & ~w21777);
assign w36287 = (w25237 & w37201) | (w25237 & w37202) | (w37201 & w37202);
assign w36288 = w25253 & w25254;
assign w36289 = (w25236 & w37201) | (w25236 & w37202) | (w37201 & w37202);
assign w36290 = (w25258 & w25257) | (w25258 & ~w21777) | (w25257 & ~w21777);
assign w36291 = (w25237 & w37203) | (w25237 & w37204) | (w37203 & w37204);
assign w36292 = w25257 & w25258;
assign w36293 = (w25236 & w37203) | (w25236 & w37204) | (w37203 & w37204);
assign w36294 = (w25262 & w25261) | (w25262 & ~w21777) | (w25261 & ~w21777);
assign w36295 = (w25237 & w37205) | (w25237 & w37206) | (w37205 & w37206);
assign w36296 = w25261 & w25262;
assign w36297 = (w25236 & w37205) | (w25236 & w37206) | (w37205 & w37206);
assign w36298 = (w25266 & w25265) | (w25266 & ~w21777) | (w25265 & ~w21777);
assign w36299 = (w25237 & w37207) | (w25237 & w37208) | (w37207 & w37208);
assign w36300 = w25265 & w25266;
assign w36301 = (w25236 & w37207) | (w25236 & w37208) | (w37207 & w37208);
assign w36302 = (w25270 & w25269) | (w25270 & ~w21777) | (w25269 & ~w21777);
assign w36303 = (w25237 & w37209) | (w25237 & w37210) | (w37209 & w37210);
assign w36304 = w25269 & w25270;
assign w36305 = (w25236 & w37209) | (w25236 & w37210) | (w37209 & w37210);
assign w36306 = (w26076 & w26075) | (w26076 & w21777) | (w26075 & w21777);
assign w36307 = (~w25237 & w37211) | (~w25237 & w37212) | (w37211 & w37212);
assign w36308 = w26075 | w26076;
assign w36309 = (~w25236 & w37211) | (~w25236 & w37212) | (w37211 & w37212);
assign w36310 = b_5 & a_11;
assign w36311 = b_5 & a_32;
assign w36312 = (w4023 & ~w3826) | (w4023 & w37213) | (~w3826 & w37213);
assign w36313 = b_4 & a_59;
assign w36314 = (~w19828 & w25191) | (~w19828 & w26969) | (w25191 & w26969);
assign w36315 = w25195 | w25194;
assign w36316 = (w25194 & w25195) | (w25194 & w26969) | (w25195 & w26969);
assign w36317 = (~w25209 & w37214) | (~w25209 & w37215) | (w37214 & w37215);
assign w36318 = (w25216 & w37216) | (w25216 & w37217) | (w37216 & w37217);
assign w36319 = (~w25221 & w37218) | (~w25221 & w37219) | (w37218 & w37219);
assign w36320 = (w25216 & w37220) | (w25216 & w37221) | (w37220 & w37221);
assign w36321 = (~w25221 & w37222) | (~w25221 & w37223) | (w37222 & w37223);
assign w36322 = (w25216 & w37224) | (w25216 & w37225) | (w37224 & w37225);
assign w36323 = (~w25221 & w37226) | (~w25221 & w37227) | (w37226 & w37227);
assign w36324 = (w25216 & w37228) | (w25216 & w37229) | (w37228 & w37229);
assign w36325 = (~w25221 & w37230) | (~w25221 & w37231) | (w37230 & w37231);
assign w36326 = (w25216 & w37232) | (w25216 & w37233) | (w37232 & w37233);
assign w36327 = (~w25221 & w37234) | (~w25221 & w37235) | (w37234 & w37235);
assign w36328 = (w25216 & w37236) | (w25216 & w37237) | (w37236 & w37237);
assign w36329 = (w25221 & w37238) | (w25221 & w37239) | (w37238 & w37239);
assign w36330 = (~w25216 & w37240) | (~w25216 & w37241) | (w37240 & w37241);
assign w36331 = ~w23909 & ~w24022;
assign w36332 = ~w24022 & w37242;
assign w36333 = (w25348 & w37242) | (w25348 & w37243) | (w37242 & w37243);
assign w36334 = ~w24222 & w25279;
assign w36335 = ~w25276 & w37244;
assign w36336 = (~w25276 & w37245) | (~w25276 & w37246) | (w37245 & w37246);
assign w36337 = (w25275 & w37246) | (w25275 & w37247) | (w37246 & w37247);
assign w36338 = (~w25276 & w37248) | (~w25276 & w37249) | (w37248 & w37249);
assign w36339 = (w25275 & w37249) | (w25275 & w37250) | (w37249 & w37250);
assign w36340 = (~w25276 & w37251) | (~w25276 & w37252) | (w37251 & w37252);
assign w36341 = (w25287 & w37253) | (w25287 & w37254) | (w37253 & w37254);
assign w36342 = ~w25292 & w37255;
assign w36343 = (w25287 & w37256) | (w25287 & w37257) | (w37256 & w37257);
assign w36344 = ~w10457 & ~w10135;
assign w36345 = ~w33744 & a_5;
assign w36346 = b_5 & a_5;
assign w36347 = ~w33745 & a_8;
assign w36348 = (~w2727 & w2909) | (~w2727 & w37258) | (w2909 & w37258);
assign w36349 = ~w33743 & a_44;
assign w36350 = ~w20307 & ~w20071;
assign w36351 = ~w20307 & w25482;
assign w36352 = ~w20307 & w25343;
assign w36353 = ~w20753 & ~w26973;
assign w36354 = (~w26866 & w37259) | (~w26866 & w37260) | (w37259 & w37260);
assign w36355 = (~w26973 & w37261) | (~w26973 & w37260) | (w37261 & w37260);
assign w36356 = (w25483 & w37260) | (w25483 & w36353) | (w37260 & w36353);
assign w36357 = (~w25196 & w36353) | (~w25196 & w37262) | (w36353 & w37262);
assign w36358 = (w25195 & w37263) | (w25195 & w37264) | (w37263 & w37264);
assign w36359 = (w25212 & w25211) | (w25212 & ~w26973) | (w25211 & ~w26973);
assign w36360 = (~w26866 & w37265) | (~w26866 & w37266) | (w37265 & w37266);
assign w36361 = (~w26973 & w37267) | (~w26973 & w37266) | (w37267 & w37266);
assign w36362 = (w25483 & w37266) | (w25483 & w36359) | (w37266 & w36359);
assign w36363 = (~w25196 & w36359) | (~w25196 & w37268) | (w36359 & w37268);
assign w36364 = (w25195 & w37269) | (w25195 & w37270) | (w37269 & w37270);
assign w36365 = (w25215 & w25216) | (w25215 & ~w26973) | (w25216 & ~w26973);
assign w36366 = (~w26866 & w37271) | (~w26866 & w37272) | (w37271 & w37272);
assign w36367 = (~w26973 & w37273) | (~w26973 & w37272) | (w37273 & w37272);
assign w36368 = (w25483 & w37272) | (w25483 & w36365) | (w37272 & w36365);
assign w36369 = (~w25196 & w36365) | (~w25196 & w37274) | (w36365 & w37274);
assign w36370 = (w25195 & w37275) | (w25195 & w37276) | (w37275 & w37276);
assign w36371 = (w26719 & w26718) | (w26719 & ~w26973) | (w26718 & ~w26973);
assign w36372 = (w26719 & w26718) | (w26719 & ~w32962) | (w26718 & ~w32962);
assign w36373 = (w26719 & w26718) | (w26719 & ~w32963) | (w26718 & ~w32963);
assign w36374 = (w25483 & w37277) | (w25483 & w36371) | (w37277 & w36371);
assign w36375 = (~w25196 & w36371) | (~w25196 & w36372) | (w36371 & w36372);
assign w36376 = (w25195 & w36373) | (w25195 & w37278) | (w36373 & w37278);
assign w36377 = ~w23127 & ~w22978;
assign w36378 = ~w22980 & w36377;
assign w36379 = ~w23272 & w25250;
assign w36380 = ~w25248 & w37279;
assign w36381 = (w25250 & w37280) | (w25250 & w37281) | (w37280 & w37281);
assign w36382 = (~w25248 & w37281) | (~w25248 & w37282) | (w37281 & w37282);
assign w36383 = (w25250 & w37283) | (w25250 & w37284) | (w37283 & w37284);
assign w36384 = (~w25248 & w37285) | (~w25248 & w37286) | (w37285 & w37286);
assign w36385 = (w25250 & w37287) | (w25250 & w37288) | (w37287 & w37288);
assign w36386 = (~w25248 & w37289) | (~w25248 & w37290) | (w37289 & w37290);
assign w36387 = ~w25263 & w37291;
assign w36388 = (~w25248 & w37292) | (~w25248 & w37293) | (w37292 & w37293);
assign w36389 = (~w25263 & w37294) | (~w25263 & w37295) | (w37294 & w37295);
assign w36390 = ~w25268 & w37296;
assign w36391 = (w25263 & w37297) | (w25263 & w37298) | (w37297 & w37298);
assign w36392 = (w25268 & w37299) | (w25268 & w37300) | (w37299 & w37300);
assign w36393 = (w25263 & w37301) | (w25263 & w37302) | (w37301 & w37302);
assign w36394 = (w25268 & w37303) | (w25268 & w37304) | (w37303 & w37304);
assign w36395 = (w25263 & w37305) | (w25263 & w37306) | (w37305 & w37306);
assign w36396 = (w25268 & w37307) | (w25268 & w37308) | (w37307 & w37308);
assign w36397 = (w25263 & w37309) | (w25263 & w37310) | (w37309 & w37310);
assign w36398 = (w25268 & w37311) | (w25268 & w37312) | (w37311 & w37312);
assign w36399 = (w25263 & w37313) | (w25263 & w37314) | (w37313 & w37314);
assign w36400 = (w25268 & w37315) | (w25268 & w37316) | (w37315 & w37316);
assign w36401 = (w25263 & w37317) | (w25263 & w37318) | (w37317 & w37318);
assign w36402 = (w25268 & w37319) | (w25268 & w37320) | (w37319 & w37320);
assign w36403 = (w25263 & w37321) | (w25263 & w37322) | (w37321 & w37322);
assign w36404 = (w25268 & w37323) | (w25268 & w37324) | (w37323 & w37324);
assign w36405 = (w25263 & w37325) | (w25263 & w37326) | (w37325 & w37326);
assign w36406 = (w25268 & w37327) | (w25268 & w37328) | (w37327 & w37328);
assign w36407 = (w25263 & w37329) | (w25263 & w37330) | (w37329 & w37330);
assign w36408 = (w25268 & w37331) | (w25268 & w37332) | (w37331 & w37332);
assign w36409 = (~w7750 & ~w7455) | (~w7750 & w37333) | (~w7455 & w37333);
assign w36410 = ~w7750 & w26569;
assign w36411 = w7519 & w37334;
assign w36412 = (w6056 & ~w5775) | (w6056 & w37335) | (~w5775 & w37335);
assign w36413 = b_4 & a_62;
assign w36414 = w9815 & w10110;
assign w36415 = ~w9815 & ~w10110;
assign w36416 = ~w10840 & ~w11155;
assign w36417 = w3769 & w4092;
assign w36418 = ~w3769 & ~w4092;
assign w36419 = w6243 & w6293;
assign w36420 = ~w6243 & ~w6293;
assign w36421 = w7072 & w7122;
assign w36422 = ~w7072 & ~w7122;
assign w36423 = w5456 & w5506;
assign w36424 = ~w5456 & ~w5506;
assign w36425 = w7939 & w7988;
assign w36426 = ~w7939 & ~w7988;
assign w36427 = w11124 & w11244;
assign w36428 = w27390 & a_2;
assign w36429 = ~w33840 & a_56;
assign w36430 = w7449 & w7725;
assign w36431 = ~w33864 & a_47;
assign w36432 = b_45 & a_23;
assign w36433 = (~w14207 & w37336) | (~w14207 & w37337) | (w37336 & w37337);
assign w36434 = b_51 & a_17;
assign w36435 = b_45 & a_26;
assign w36436 = b_50 & a_23;
assign w36437 = b_48 & a_29;
assign w36438 = b_49 & a_29;
assign w36439 = b_45 & a_35;
assign w36440 = b_50 & a_32;
assign w36441 = b_45 & a_38;
assign w36442 = b_48 & a_35;
assign w36443 = b_47 & a_41;
assign w36444 = b_42 & a_47;
assign w36445 = b_45 & a_44;
assign w36446 = b_43 & a_47;
assign w36447 = b_49 & a_41;
assign w36448 = b_46 & a_47;
assign w36449 = (w21573 & ~w21346) | (w21573 & w37338) | (~w21346 & w37338);
assign w36450 = b_46 & a_53;
assign w36451 = b_44 & a_59;
assign w36452 = b_47 & a_59;
assign w36453 = w23607 & ~w23442;
assign w36454 = b_51 & a_62;
assign w36455 = b_57 & a_62;
assign w36456 = b_59 & a_62;
assign w36457 = ~w5917 & w6098;
assign w36458 = w5917 & ~w6098;
assign w36459 = w1353 & w37339;
assign w36460 = (~w1508 & w1355) | (~w1508 & w37340) | (w1355 & w37340);
assign w36461 = (w8126 & ~w7812) | (w8126 & w37341) | (~w7812 & w37341);
assign w36462 = w25156 & w25155;
assign w36463 = (w25155 & w25156) | (w25155 & ~w15844) | (w25156 & ~w15844);
assign w36464 = w12723 & w13327;
assign w36465 = ~w12723 & ~w13327;
assign w36466 = w25163 | w25162;
assign w36467 = (w25162 & w25163) | (w25162 & w16489) | (w25163 & w16489);
assign w36468 = (w13469 & w13693) | (w13469 & w37342) | (w13693 & w37342);
assign w36469 = w37343 & ~w13776;
assign w36470 = b_48 & a_23;
assign w36471 = b_52 & a_20;
assign w36472 = w12701 & w13046;
assign w36473 = w8213 & w8687;
assign w36474 = w8422 & w8723;
assign w36475 = w12616 & w12677;
assign w36476 = w27862 & a_2;
assign w36477 = b_8 & a_5;
assign w36478 = b_8 & a_8;
assign w36479 = b_8 & a_11;
assign w36480 = b_8 & a_14;
assign w36481 = b_8 & a_17;
assign w36482 = b_5 & a_23;
assign w36483 = b_8 & a_20;
assign w36484 = b_18 & a_11;
assign w36485 = b_13 & a_17;
assign w36486 = b_16 & a_14;
assign w36487 = b_19 & a_11;
assign w36488 = b_8 & a_23;
assign w36489 = b_17 & a_14;
assign w36490 = w2752 & w37344;
assign w36491 = ~w2959 & ~w28240;
assign w36492 = (w2935 & w37345) | (w2935 & ~w2959) | (w37345 & ~w2959);
assign w36493 = b_18 & a_14;
assign w36494 = (w2793 & ~w2752) | (w2793 & w37346) | (~w2752 & w37346);
assign w36495 = b_10 & a_23;
assign w36496 = b_19 & a_14;
assign w36497 = ~b_19 & a_14;
assign w36498 = b_22 & a_11;
assign w36499 = b_8 & a_26;
assign w36500 = b_23 & a_11;
assign w36501 = b_12 & a_23;
assign w36502 = b_24 & a_11;
assign w36503 = ~w3341 & ~w3541;
assign w36504 = b_19 & a_17;
assign w36505 = b_22 & a_14;
assign w36506 = b_25 & a_11;
assign w36507 = b_28 & a_8;
assign w36508 = b_29 & a_8;
assign w36509 = b_8 & a_29;
assign w36510 = ~w4391 & ~w4632;
assign w36511 = b_8 & a_32;
assign w36512 = b_33 & a_8;
assign w36513 = ~b_33 & a_8;
assign w36514 = b_35 & a_8;
assign w36515 = ~b_35 & a_8;
assign w36516 = b_32 & a_11;
assign w36517 = b_8 & a_35;
assign w36518 = b_33 & a_11;
assign w36519 = b_36 & a_8;
assign w36520 = b_8 & a_38;
assign w36521 = b_38 & a_8;
assign w36522 = ~w5860 & ~w5884;
assign w36523 = b_39 & a_8;
assign w36524 = ~b_39 & a_8;
assign w36525 = b_8 & a_41;
assign w36526 = b_38 & a_11;
assign w36527 = b_36 & a_14;
assign w36528 = b_42 & a_8;
assign w36529 = b_37 & a_14;
assign w36530 = b_43 & a_8;
assign w36531 = ~w7280 & ~w6994;
assign w36532 = b_8 & a_44;
assign w36533 = b_38 & a_14;
assign w36534 = ~b_41 & a_11;
assign w36535 = b_44 & a_8;
assign w36536 = b_47 & a_5;
assign w36537 = b_36 & a_17;
assign w36538 = b_31 & a_23;
assign w36539 = b_34 & a_20;
assign w36540 = ~w8182 & ~w8158;
assign w36541 = b_35 & a_20;
assign w36542 = b_32 & a_23;
assign w36543 = b_8 & a_47;
assign w36544 = w9084 & w37347;
assign w36545 = (w8192 & w37348) | (w8192 & w37349) | (w37348 & w37349);
assign w36546 = (~w9115 & ~w9084) | (~w9115 & w37350) | (~w9084 & w37350);
assign w36547 = (~w8192 & w37351) | (~w8192 & w37352) | (w37351 & w37352);
assign w36548 = w9084 & w37353;
assign w36549 = (w8192 & w37354) | (w8192 & w37355) | (w37354 & w37355);
assign w36550 = ~w9107 & ~w9106;
assign w36551 = w9131 & ~w36550;
assign w36552 = ~w9131 & w36550;
assign w36553 = b_18 & a_38;
assign w36554 = b_36 & a_20;
assign w36555 = b_48 & a_8;
assign w36556 = b_49 & a_8;
assign w36557 = b_28 & a_29;
assign w36558 = b_31 & a_26;
assign w36559 = b_34 & a_23;
assign w36560 = ~w9130 & ~w9106;
assign w36561 = b_8 & a_50;
assign w36562 = b_26 & a_32;
assign w36563 = b_18 & a_41;
assign w36564 = b_36 & a_23;
assign w36565 = b_52 & a_8;
assign w36566 = b_25 & a_35;
assign w36567 = b_31 & a_29;
assign w36568 = b_14 & a_47;
assign w36569 = b_8 & a_53;
assign w36570 = b_26 & a_35;
assign w36571 = b_32 & a_29;
assign w36572 = b_24 & a_38;
assign w36573 = b_30 & a_32;
assign w36574 = b_52 & a_11;
assign w36575 = b_25 & a_38;
assign w36576 = b_34 & a_29;
assign w36577 = ~w11165 & ~w11192;
assign w36578 = b_5 & a_59;
assign w36579 = b_8 & a_56;
assign w36580 = b_26 & a_38;
assign w36581 = b_35 & a_29;
assign w36582 = b_51 & a_14;
assign w36583 = b_27 & a_38;
assign w36584 = b_36 & a_29;
assign w36585 = b_54 & a_11;
assign w36586 = b_60 & a_5;
assign w36587 = (~w12232 & w37356) | (~w12232 & w37357) | (w37356 & w37357);
assign w36588 = (w12651 & ~w12232) | (w12651 & w37358) | (~w12232 & w37358);
assign w36589 = ~w12269 & ~b_62;
assign w36590 = w12643 & ~b_62;
assign w36591 = ~w8 & w37359;
assign w36592 = w12 & w34715;
assign w36593 = w12 & w34716;
assign w36594 = b_63 & a_2;
assign w36595 = b_52 & a_14;
assign w36596 = b_34 & a_32;
assign w36597 = b_28 & a_38;
assign w36598 = b_43 & a_23;
assign w36599 = b_61 & a_5;
assign w36600 = b_5 & a_62;
assign w36601 = b_8 & a_59;
assign w36602 = b_32 & a_35;
assign w36603 = b_38 & a_29;
assign w36604 = b_50 & a_17;
assign w36605 = ~w8 & w29810;
assign w36606 = b_48 & a_20;
assign w36607 = b_55 & a_14;
assign w36608 = b_43 & a_26;
assign w36609 = w37360 & w13850;
assign w36610 = (w13627 & w37361) | (w13627 & w13645) | (w37361 & w13645);
assign w36611 = ~w12641 & w14109;
assign w36612 = w14109 & ~w34715;
assign w36613 = w14109 & ~w34716;
assign w36614 = w33983 & ~w14164;
assign w36615 = w14046 & ~w14164;
assign w36616 = w33983 & w14164;
assign w36617 = w14046 & w14164;
assign w36618 = b_41 & a_29;
assign w36619 = b_8 & a_62;
assign w36620 = (w13632 & w37362) | (w13632 & w37363) | (w37362 & w37363);
assign w36621 = (w13989 & w13632) | (w13989 & w37364) | (w13632 & w37364);
assign w36622 = w14468 & w14454;
assign w36623 = w33986 & ~w14499;
assign w36624 = ~w14499 & ~w14468;
assign w36625 = (w14067 & w36624) | (w14067 & w37365) | (w36624 & w37365);
assign w36626 = w37366 & ~w14154;
assign w36627 = b_54 & a_17;
assign w36628 = (~w14432 & w14556) | (~w14432 & w37367) | (w14556 & w37367);
assign w36629 = (w14432 & w14556) | (w14432 & w37368) | (w14556 & w37368);
assign w36630 = (w14346 & w37369) | (w14346 & w14374) | (w37369 & w14374);
assign w36631 = w14331 & w30156;
assign w36632 = (w14331 & w13895) | (w14331 & w37370) | (w13895 & w37370);
assign w36633 = w14251 & w30151;
assign w36634 = w14251 & ~w13861;
assign w36635 = b_51 & a_20;
assign w36636 = ~w12641 & w14841;
assign w36637 = w14841 & ~w34715;
assign w36638 = w14841 & ~w34716;
assign w36639 = b_55 & a_17;
assign w36640 = ~w15136 & ~w14940;
assign w36641 = w15136 & w14940;
assign w36642 = w15136 & ~w14940;
assign w36643 = (w15083 & ~w14657) | (w15083 & w37371) | (~w14657 & w37371);
assign w36644 = ~w15411 & ~w30373;
assign w36645 = w15163 & ~w15505;
assign w36646 = w15561 & ~w15453;
assign w36647 = w15561 & w15453;
assign w36648 = w15590 & ~w15428;
assign w36649 = w15590 & w15428;
assign w36650 = ~w15411 & ~w15235;
assign w36651 = w15412 & w30372;
assign w36652 = w15412 & ~w15127;
assign w36653 = b_51 & a_23;
assign w36654 = ~w15503 & ~w15843;
assign w36655 = ~w15842 & w37372;
assign w36656 = b_55 & a_20;
assign w36657 = w15804 & w15874;
assign w36658 = ~w15804 & ~w15874;
assign w36659 = b_43 & a_32;
assign w36660 = w34917 & ~w16141;
assign w36661 = ~w34917 & ~w16141;
assign w36662 = ~w12641 & w16158;
assign w36663 = w16158 & ~w34715;
assign w36664 = w16158 & ~w34716;
assign w36665 = (~w16162 & w15830) | (~w16162 & w37373) | (w15830 & w37373);
assign w36666 = w25152 & ~w16174;
assign w36667 = (~w16174 & w25152) | (~w16174 & ~w15844) | (w25152 & ~w15844);
assign w36668 = w25154 | w25153;
assign w36669 = (w25153 & w25154) | (w25153 & w15844) | (w25154 & w15844);
assign w36670 = (~w15797 & w37374) | (~w15797 & w36672) | (w37374 & w36672);
assign w36671 = ~w15797 & w37374;
assign w36672 = ~w15607 & w37374;
assign w36673 = (w15797 & w37375) | (w15797 & w36675) | (w37375 & w36675);
assign w36674 = (w16238 & w15797) | (w16238 & w37375) | (w15797 & w37375);
assign w36675 = (w16238 & w15607) | (w16238 & w37375) | (w15607 & w37375);
assign w36676 = w15927 & ~w16263;
assign w36677 = ~w15927 & w16263;
assign w36678 = (w16007 & w15662) | (w16007 & w37376) | (w15662 & w37376);
assign w36679 = w16489 & ~w16486;
assign w36680 = b_54 & a_23;
assign w36681 = ~w16288 & ~w16692;
assign w36682 = b_45 & a_32;
assign w36683 = (~w16263 & w16774) | (~w16263 & w37377) | (w16774 & w37377);
assign w36684 = ~w16775 & w34999;
assign w36685 = w25157 & ~w16803;
assign w36686 = (~w16803 & w25157) | (~w16803 & ~w16489) | (w25157 & ~w16489);
assign w36687 = (w25341 & w37378) | (w25341 & w37379) | (w37378 & w37379);
assign w36688 = (w25158 & w25159) | (w25158 & w16489) | (w25159 & w16489);
assign w36689 = (~w16577 & w37380) | (~w16577 & w16559) | (w37380 & w16559);
assign w36690 = w16094 & w37381;
assign w36691 = (w16094 & w37381) | (w16094 & w37382) | (w37381 & w37382);
assign w36692 = w37383 & w16914;
assign w36693 = w16912 & w16914;
assign w36694 = (~w16914 & w37384) | (~w16914 & a_62) | (w37384 & a_62);
assign w36695 = w37385 & ~w17070;
assign w36696 = ~w16781 & w37386;
assign w36697 = ~w12641 & w17105;
assign w36698 = w17105 & ~w34715;
assign w36699 = w17105 & ~w34716;
assign w36700 = w25161 & w25160;
assign w36701 = (w25160 & w25161) | (w25160 & ~w16489) | (w25161 & ~w16489);
assign w36702 = (~w16493 & w37387) | (~w16493 & w37388) | (w37387 & w37388);
assign w36703 = ~w16801 & w37389;
assign w36704 = b_56 & a_23;
assign w36705 = w17172 & ~w35060;
assign w36706 = (w16097 & w37390) | (w16097 & w37391) | (w37390 & w37391);
assign w36707 = ~w17172 & w35060;
assign w36708 = (~w16097 & w37392) | (~w16097 & w37393) | (w37392 & w37393);
assign w36709 = (w16863 & ~w16732) | (w16863 & w37394) | (~w16732 & w37394);
assign w36710 = w37395 & w16914;
assign w36711 = ~a_62 & w17230;
assign w36712 = a_62 & ~w17230;
assign w36713 = (w16898 & ~w16682) | (w16898 & w37396) | (~w16682 & w37396);
assign w36714 = ~w17403 & ~w17088;
assign w36715 = (~w16563 & w36714) | (~w16563 & w37397) | (w36714 & w37397);
assign w36716 = w17403 & ~w30936;
assign w36717 = w17417 & w17118;
assign w36718 = (w17417 & ~w17121) | (w17417 & w36717) | (~w17121 & w36717);
assign w36719 = w17417 & ~w32936;
assign w36720 = w17417 & ~w32937;
assign w36721 = (~w25158 & w36717) | (~w25158 & w37398) | (w36717 & w37398);
assign w36722 = (~w25341 & w36719) | (~w25341 & w36720) | (w36719 & w36720);
assign w36723 = w17417 & ~w36467;
assign w36724 = ~w25163 & w37399;
assign w36725 = ~w17417 & ~w17118;
assign w36726 = w17121 & w36725;
assign w36727 = ~w17417 & w32936;
assign w36728 = ~w17417 & w32937;
assign w36729 = (w25158 & w36725) | (w25158 & w37400) | (w36725 & w37400);
assign w36730 = (w25341 & w36727) | (w25341 & w36728) | (w36727 & w36728);
assign w36731 = ~w17417 & w36467;
assign w36732 = (~w17417 & w25163) | (~w17417 & w37401) | (w25163 & w37401);
assign w36733 = w17473 & ~w35100;
assign w36734 = (~w16445 & w37402) | (~w16445 & w37403) | (w37402 & w37403);
assign w36735 = ~w17473 & w35100;
assign w36736 = (w16445 & w37404) | (w16445 & w37405) | (w37404 & w37405);
assign w36737 = b_51 & a_29;
assign w36738 = (~w17008 & w37406) | (~w17008 & w37407) | (w37406 & w37407);
assign w36739 = (w17346 & ~w17008) | (w17346 & w37408) | (~w17008 & w37408);
assign w36740 = (w25341 & w37411) | (w25341 & w37412) | (w37411 & w37412);
assign w36741 = (~w17415 & w25164) | (~w17415 & w36467) | (w25164 & w36467);
assign w36742 = (w25163 & w37413) | (w25163 & w37414) | (w37413 & w37414);
assign w36743 = (~w25164 & w37415) | (~w25164 & w37416) | (w37415 & w37416);
assign w36744 = (w25165 & w25166) | (w25165 & ~w25479) | (w25166 & ~w25479);
assign w36745 = (w25165 & w25166) | (w25165 & ~w32936) | (w25166 & ~w32936);
assign w36746 = (w25165 & w25166) | (w25165 & ~w32937) | (w25166 & ~w32937);
assign w36747 = (~w25158 & w37417) | (~w25158 & w36744) | (w37417 & w36744);
assign w36748 = (~w25341 & w36745) | (~w25341 & w36746) | (w36745 & w36746);
assign w36749 = (w25165 & w25166) | (w25165 & ~w36467) | (w25166 & ~w36467);
assign w36750 = (~w25163 & w37418) | (~w25163 & w37419) | (w37418 & w37419);
assign w36751 = (w25158 & w37420) | (w25158 & w37421) | (w37420 & w37421);
assign w36752 = ~w17711 & w36740;
assign w36753 = ~w12641 & w17718;
assign w36754 = w17718 & ~w34715;
assign w36755 = w17718 & ~w34716;
assign w36756 = ~w17748 & w35140;
assign w36757 = (w16778 & w37422) | (w16778 & w37423) | (w37422 & w37423);
assign w36758 = w17748 & ~w35140;
assign w36759 = (~w16778 & w37424) | (~w16778 & w37425) | (w37424 & w37425);
assign w36760 = (w25168 & w25167) | (w25168 & ~w17118) | (w25167 & ~w17118);
assign w36761 = (w25168 & w25167) | (w25168 & w25479) | (w25167 & w25479);
assign w36762 = (w25168 & w25167) | (w25168 & w32936) | (w25167 & w32936);
assign w36763 = (w25168 & w25167) | (w25168 & w32937) | (w25167 & w32937);
assign w36764 = (w25158 & w36760) | (w25158 & w36761) | (w36760 & w36761);
assign w36765 = (w25341 & w36762) | (w25341 & w36763) | (w36762 & w36763);
assign w36766 = ~w17990 & w36760;
assign w36767 = (w25479 & w37426) | (w25479 & w37427) | (w37426 & w37427);
assign w36768 = (w25342 & w37428) | (w25342 & w37429) | (w37428 & w37429);
assign w36769 = (~w17989 & w25169) | (~w17989 & w25167) | (w25169 & w25167);
assign w36770 = (w25158 & w36772) | (w25158 & w36773) | (w36772 & w36773);
assign w36771 = (~w17989 & w25169) | (~w17989 & w36765) | (w25169 & w36765);
assign w36772 = (~w17989 & w25169) | (~w17989 & w36760) | (w25169 & w36760);
assign w36773 = (w25479 & w37430) | (w25479 & w36769) | (w37430 & w36769);
assign w36774 = b_56 & a_26;
assign w36775 = ~w35175 & w18043;
assign w36776 = w35175 & ~w18043;
assign w36777 = (w17964 & w17642) | (w17964 & w37431) | (w17642 & w37431);
assign w36778 = (w17856 & w37432) | (w17856 & w17884) | (w37432 & w17884);
assign w36779 = (~w17503 & w37433) | (~w17503 & w37434) | (w37433 & w37434);
assign w36780 = ~w17842 & ~w31133;
assign w36781 = (w17503 & w37435) | (w17503 & w37436) | (w37435 & w37436);
assign w36782 = w17842 & w31133;
assign w36783 = (w17901 & ~w17541) | (w17901 & w37437) | (~w17541 & w37437);
assign w36784 = (w17926 & ~w17575) | (w17926 & w37438) | (~w17575 & w37438);
assign w36785 = b_47 & a_35;
assign w36786 = (~w25342 & w37439) | (~w25342 & w37440) | (w37439 & w37440);
assign w36787 = (w25170 & w25171) | (w25170 & ~w25167) | (w25171 & ~w25167);
assign w36788 = (~w25158 & w36790) | (~w25158 & w36791) | (w36790 & w36791);
assign w36789 = (w25170 & w25171) | (w25170 & ~w36765) | (w25171 & ~w36765);
assign w36790 = (w25170 & w25171) | (w25170 & ~w36760) | (w25171 & ~w36760);
assign w36791 = (~w25479 & w37441) | (~w25479 & w36787) | (w37441 & w36787);
assign w36792 = ~w18273 & ~w17989;
assign w36793 = ~w17990 & w36792;
assign w36794 = (w25158 & w36796) | (w25158 & w36797) | (w36796 & w36797);
assign w36795 = (w25172 & w25173) | (w25172 & w36765) | (w25173 & w36765);
assign w36796 = (w25172 & w25173) | (w25172 & w36760) | (w25173 & w36760);
assign w36797 = (w25479 & w37442) | (w25479 & w37443) | (w37442 & w37443);
assign w36798 = (~w25342 & w37444) | (~w25342 & w37445) | (w37444 & w37445);
assign w36799 = (w25174 & w25175) | (w25174 & ~w25167) | (w25175 & ~w25167);
assign w36800 = (~w25158 & w36802) | (~w25158 & w36803) | (w36802 & w36803);
assign w36801 = (w25174 & w25175) | (w25174 & ~w36765) | (w25175 & ~w36765);
assign w36802 = (w25174 & w25175) | (w25174 & ~w36760) | (w25175 & ~w36760);
assign w36803 = (~w25479 & w37446) | (~w25479 & w36799) | (w37446 & w36799);
assign w36804 = ~w18547 & w25172;
assign w36805 = ~w25171 & w37447;
assign w36806 = (w25158 & w36808) | (w25158 & w36809) | (w36808 & w36809);
assign w36807 = (w25176 & w25177) | (w25176 & w36765) | (w25177 & w36765);
assign w36808 = (w25176 & w25177) | (w25176 & w36760) | (w25177 & w36760);
assign w36809 = (w25479 & w37448) | (w25479 & w37449) | (w37448 & w37449);
assign w36810 = b_52 & a_32;
assign w36811 = b_46 & a_38;
assign w36812 = ~w12641 & w18801;
assign w36813 = w18801 & ~w34715;
assign w36814 = w18801 & ~w34716;
assign w36815 = (~w25172 & w37450) | (~w25172 & w37451) | (w37450 & w37451);
assign w36816 = (w25171 & w37451) | (w25171 & w37452) | (w37451 & w37452);
assign w36817 = (~w25158 & w37453) | (~w25158 & w37454) | (w37453 & w37454);
assign w36818 = (~w36765 & w37455) | (~w36765 & w37456) | (w37455 & w37456);
assign w36819 = (w25172 & w37457) | (w25172 & w37458) | (w37457 & w37458);
assign w36820 = (~w25171 & w37458) | (~w25171 & w37459) | (w37458 & w37459);
assign w36821 = (w25158 & w37460) | (w25158 & w37461) | (w37460 & w37461);
assign w36822 = (w36765 & w37462) | (w36765 & w37463) | (w37462 & w37463);
assign w36823 = (w25172 & w37464) | (w25172 & w37465) | (w37464 & w37465);
assign w36824 = (~w25171 & w37465) | (~w25171 & w37466) | (w37465 & w37466);
assign w36825 = (w25158 & w37467) | (w25158 & w37468) | (w37467 & w37468);
assign w36826 = (w36765 & w37469) | (w36765 & w37470) | (w37469 & w37470);
assign w36827 = w35283 & ~w18869;
assign w36828 = ~w36827 & ~w18869;
assign w36829 = b_53 & a_32;
assign w36830 = (w18715 & ~w18382) | (w18715 & w37471) | (~w18382 & w37471);
assign w36831 = ~a_62 & w18950;
assign w36832 = a_62 & ~w18950;
assign w36833 = b_47 & a_38;
assign w36834 = (~w25172 & w37472) | (~w25172 & w37473) | (w37472 & w37473);
assign w36835 = (w25171 & w37473) | (w25171 & w37474) | (w37473 & w37474);
assign w36836 = (~w25158 & w37475) | (~w25158 & w37476) | (w37475 & w37476);
assign w36837 = (~w36765 & w37477) | (~w36765 & w37478) | (w37477 & w37478);
assign w36838 = w19197 & w31396;
assign w36839 = (w19197 & w18933) | (w19197 & w37479) | (w18933 & w37479);
assign w36840 = w18933 | ~w18966;
assign w36841 = ~w19197 & ~w31396;
assign w36842 = ~w18933 & w37480;
assign w36843 = b_45 & a_41;
assign w36844 = b_48 & a_38;
assign w36845 = (w25172 & w37481) | (w25172 & w37482) | (w37481 & w37482);
assign w36846 = (~w25171 & w37482) | (~w25171 & w37483) | (w37482 & w37483);
assign w36847 = (w25158 & w37484) | (w25158 & w37485) | (w37484 & w37485);
assign w36848 = (w36765 & w37486) | (w36765 & w37487) | (w37486 & w37487);
assign w36849 = (~w25172 & w37488) | (~w25172 & w37489) | (w37488 & w37489);
assign w36850 = (w25171 & w37489) | (w25171 & w37490) | (w37489 & w37490);
assign w36851 = (~w25158 & w37491) | (~w25158 & w37492) | (w37491 & w37492);
assign w36852 = (~w36765 & w37493) | (~w36765 & w37494) | (w37493 & w37494);
assign w36853 = ~w12641 & w19345;
assign w36854 = w19345 & ~w34715;
assign w36855 = w19345 & ~w34716;
assign w36856 = b_46 & a_41;
assign w36857 = (w25172 & w37495) | (w25172 & w37496) | (w37495 & w37496);
assign w36858 = (~w25171 & w37496) | (~w25171 & w37497) | (w37496 & w37497);
assign w36859 = (w25158 & w37498) | (w25158 & w37499) | (w37498 & w37499);
assign w36860 = (w36765 & w37500) | (w36765 & w37501) | (w37500 & w37501);
assign w36861 = (~w25172 & w37502) | (~w25172 & w37503) | (w37502 & w37503);
assign w36862 = (w25171 & w37503) | (w25171 & w37504) | (w37503 & w37504);
assign w36863 = (~w25158 & w37505) | (~w25158 & w37506) | (w37505 & w37506);
assign w36864 = (~w36765 & w37507) | (~w36765 & w37508) | (w37507 & w37508);
assign w36865 = (w25342 & w37509) | (w25342 & w37510) | (w37509 & w37510);
assign w36866 = (w27076 & w27075) | (w27076 & w25167) | (w27075 & w25167);
assign w36867 = (w25158 & w36869) | (w25158 & w36870) | (w36869 & w36870);
assign w36868 = (w27076 & w27075) | (w27076 & w36765) | (w27075 & w36765);
assign w36869 = (w27076 & w27075) | (w27076 & w36760) | (w27075 & w36760);
assign w36870 = (w25479 & w37511) | (w25479 & w36866) | (w37511 & w36866);
assign w36871 = w35420 & ~w19620;
assign w36872 = ~w35420 & ~w19620;
assign w36873 = b_56 & a_32;
assign w36874 = (w19562 & ~w19288) | (w19562 & w37512) | (~w19288 & w37512);
assign w36875 = (w19403 & ~w19235) | (w19403 & w37513) | (~w19235 & w37513);
assign w36876 = (w19451 & w37514) | (w19451 & w19479) | (w37514 & w19479);
assign w36877 = ~a_62 & w19681;
assign w36878 = a_62 & ~w19681;
assign w36879 = (w19498 & w19214) | (w19498 & w37515) | (w19214 & w37515);
assign w36880 = (~w25172 & w37516) | (~w25172 & w37517) | (w37516 & w37517);
assign w36881 = (w25171 & w37516) | (w25171 & w37518) | (w37516 & w37518);
assign w36882 = (~w25158 & w37519) | (~w25158 & w37520) | (w37519 & w37520);
assign w36883 = (~w36765 & w37521) | (~w36765 & w37522) | (w37521 & w37522);
assign w36884 = (~w25167 & w37521) | (~w25167 & w37522) | (w37521 & w37522);
assign w36885 = (~w25342 & w37523) | (~w25342 & w37524) | (w37523 & w37524);
assign w36886 = (w25172 & w37525) | (w25172 & w37526) | (w37525 & w37526);
assign w36887 = (~w25171 & w37525) | (~w25171 & w37527) | (w37525 & w37527);
assign w36888 = (w25158 & w37528) | (w25158 & w37529) | (w37528 & w37529);
assign w36889 = (w36765 & w37530) | (w36765 & w37531) | (w37530 & w37531);
assign w36890 = (w25167 & w37530) | (w25167 & w37531) | (w37530 & w37531);
assign w36891 = (w25342 & w37532) | (w25342 & w37533) | (w37532 & w37533);
assign w36892 = b_39 & a_50;
assign w36893 = (~w19506 & w37534) | (~w19506 & w37535) | (w37534 & w37535);
assign w36894 = (w19785 & ~w19506) | (w19785 & w37536) | (~w19506 & w37536);
assign w36895 = (~w25172 & w37537) | (~w25172 & w37538) | (w37537 & w37538);
assign w36896 = (w25171 & w37537) | (w25171 & w37539) | (w37537 & w37539);
assign w36897 = (~w25158 & w37540) | (~w25158 & w37541) | (w37540 & w37541);
assign w36898 = (~w36765 & w37542) | (~w36765 & w37543) | (w37542 & w37543);
assign w36899 = (~w25167 & w37542) | (~w25167 & w37543) | (w37542 & w37543);
assign w36900 = (~w25342 & w37544) | (~w25342 & w37545) | (w37544 & w37545);
assign w36901 = (w25172 & w37546) | (w25172 & w37547) | (w37546 & w37547);
assign w36902 = (~w25171 & w37547) | (~w25171 & w37548) | (w37547 & w37548);
assign w36903 = (w25158 & w37549) | (w25158 & w37550) | (w37549 & w37550);
assign w36904 = (w36765 & w37551) | (w36765 & w37552) | (w37551 & w37552);
assign w36905 = b_40 & a_50;
assign w36906 = ~w12641 & w20293;
assign w36907 = w20293 & ~w34715;
assign w36908 = w20293 & ~w34716;
assign w36909 = (~w25172 & w37553) | (~w25172 & w37554) | (w37553 & w37554);
assign w36910 = (w25171 & w37553) | (w25171 & w37555) | (w37553 & w37555);
assign w36911 = (~w25158 & w37556) | (~w25158 & w37557) | (w37556 & w37557);
assign w36912 = (~w36765 & w37558) | (~w36765 & w37559) | (w37558 & w37559);
assign w36913 = (~w25167 & w37558) | (~w25167 & w37559) | (w37558 & w37559);
assign w36914 = (~w25342 & w37560) | (~w25342 & w37561) | (w37560 & w37561);
assign w36915 = (w25172 & w37562) | (w25172 & w37563) | (w37562 & w37563);
assign w36916 = (~w25171 & w37563) | (~w25171 & w37564) | (w37563 & w37564);
assign w36917 = (w25158 & w37565) | (w25158 & w37566) | (w37565 & w37566);
assign w36918 = (w36765 & w37567) | (w36765 & w37568) | (w37567 & w37568);
assign w36919 = (w25172 & w37569) | (w25172 & w37570) | (w37569 & w37570);
assign w36920 = (~w25171 & w37569) | (~w25171 & w37571) | (w37569 & w37571);
assign w36921 = (w25158 & w37572) | (w25158 & w37573) | (w37572 & w37573);
assign w36922 = (w36765 & w37574) | (w36765 & w37575) | (w37574 & w37575);
assign w36923 = (w25167 & w37574) | (w25167 & w37575) | (w37574 & w37575);
assign w36924 = (w25342 & w37576) | (w25342 & w37577) | (w37576 & w37577);
assign w36925 = b_44 & a_47;
assign w36926 = b_50 & a_41;
assign w36927 = (~w25158 & w37578) | (~w25158 & w37579) | (w37578 & w37579);
assign w36928 = (~w36765 & w37580) | (~w36765 & w37581) | (w37580 & w37581);
assign w36929 = (~w25167 & w37580) | (~w25167 & w37581) | (w37580 & w37581);
assign w36930 = (~w25342 & w37582) | (~w25342 & w37583) | (w37582 & w37583);
assign w36931 = b_42 & a_50;
assign w36932 = ~w20704 & w20717;
assign w36933 = w20704 & ~w20717;
assign w36934 = (w25172 & w37584) | (w25172 & w37585) | (w37584 & w37585);
assign w36935 = (~w25171 & w37584) | (~w25171 & w37586) | (w37584 & w37586);
assign w36936 = (w25158 & w37587) | (w25158 & w37588) | (w37587 & w37588);
assign w36937 = (w36765 & w37589) | (w36765 & w37590) | (w37589 & w37590);
assign w36938 = (w25167 & w37589) | (w25167 & w37590) | (w37589 & w37590);
assign w36939 = (w25342 & w37591) | (w25342 & w37592) | (w37591 & w37592);
assign w36940 = (~w25172 & w37593) | (~w25172 & w37594) | (w37593 & w37594);
assign w36941 = (w25171 & w37594) | (w25171 & w37595) | (w37594 & w37595);
assign w36942 = (~w25158 & w37596) | (~w25158 & w37597) | (w37596 & w37597);
assign w36943 = (~w36765 & w37598) | (~w36765 & w37599) | (w37598 & w37599);
assign w36944 = ~w20759 & w37600;
assign w36945 = ~w20759 & w37601;
assign w36946 = ~w20759 & w37602;
assign w36947 = b_43 & a_50;
assign w36948 = b_31 & a_62;
assign w36949 = b_49 & a_44;
assign w36950 = (w25158 & w37603) | (w25158 & w37604) | (w37603 & w37604);
assign w36951 = (w36765 & w36952) | (w36765 & w36953) | (w36952 & w36953);
assign w36952 = (w25172 & w37605) | (w25172 & w37606) | (w37605 & w37606);
assign w36953 = (~w25171 & w37606) | (~w25171 & w37607) | (w37606 & w37607);
assign w36954 = w20950 & ~w20703;
assign w36955 = w20950 & w31798;
assign w36956 = (w20804 & ~w20626) | (w20804 & w37608) | (~w20626 & w37608);
assign w36957 = b_44 & a_50;
assign w36958 = b_50 & a_44;
assign w36959 = (w25172 & w37609) | (w25172 & w37610) | (w37609 & w37610);
assign w36960 = (~w25171 & w37609) | (~w25171 & w37611) | (w37609 & w37611);
assign w36961 = (w25158 & w37612) | (w25158 & w37613) | (w37612 & w37613);
assign w36962 = (w36765 & w37614) | (w36765 & w37615) | (w37614 & w37615);
assign w36963 = (w26934 & w26933) | (w26934 & w36866) | (w26933 & w36866);
assign w36964 = (w26934 & w26933) | (w26934 & w36865) | (w26933 & w36865);
assign w36965 = (w27083 & w27084) | (w27083 & w25176) | (w27084 & w25176);
assign w36966 = (w27083 & w27084) | (w27083 & w25177) | (w27084 & w25177);
assign w36967 = (w27083 & w27084) | (w27083 & w36806) | (w27084 & w36806);
assign w36968 = (w27083 & w27084) | (w27083 & w36807) | (w27084 & w36807);
assign w36969 = b_39 & a_56;
assign w36970 = ~w12641 & w21395;
assign w36971 = w21395 & ~w34715;
assign w36972 = w21395 & ~w34716;
assign w36973 = b_40 & a_56;
assign w36974 = b_34 & a_62;
assign w36975 = b_52 & a_44;
assign w36976 = ~w21549 & w21325;
assign w36977 = ~w21549 & ~w31967;
assign w36978 = w21549 & ~w21325;
assign w36979 = w21549 & w31967;
assign w36980 = (w27085 & w27086) | (w27085 & w25176) | (w27086 & w25176);
assign w36981 = (w27085 & w27086) | (w27085 & w25177) | (w27086 & w25177);
assign w36982 = (w27085 & w27086) | (w27085 & w36806) | (w27086 & w36806);
assign w36983 = (w27085 & w27086) | (w27085 & w36807) | (w27086 & w36807);
assign w36984 = b_56 & a_41;
assign w36985 = b_53 & a_44;
assign w36986 = b_41 & a_56;
assign w36987 = (w26936 & w26935) | (w26936 & w27076) | (w26935 & w27076);
assign w36988 = (w26936 & w26935) | (w26936 & w27075) | (w26935 & w27075);
assign w36989 = (w26936 & w26935) | (w26936 & w36867) | (w26935 & w36867);
assign w36990 = (w26936 & w26935) | (w26936 & w36868) | (w26935 & w36868);
assign w36991 = (w26936 & w26935) | (w26936 & w36866) | (w26935 & w36866);
assign w36992 = (w26936 & w26935) | (w26936 & w36865) | (w26935 & w36865);
assign w36993 = (w26844 & w26843) | (w26844 & w27076) | (w26843 & w27076);
assign w36994 = (w26844 & w26843) | (w26844 & w27075) | (w26843 & w27075);
assign w36995 = (w26844 & w26843) | (w26844 & w36867) | (w26843 & w36867);
assign w36996 = (w26844 & w26843) | (w26844 & w36868) | (w26843 & w36868);
assign w36997 = (w26844 & w26843) | (w26844 & w36866) | (w26843 & w36866);
assign w36998 = (w26844 & w26843) | (w26844 & w36865) | (w26843 & w36865);
assign w36999 = b_39 & a_59;
assign w37000 = b_54 & a_44;
assign w37001 = ~w12641 & w21968;
assign w37002 = w21968 & ~w34715;
assign w37003 = w21968 & ~w34716;
assign w37004 = b_43 & a_56;
assign w37005 = b_49 & a_50;
assign w37006 = (w26938 & w26937) | (w26938 & w27076) | (w26937 & w27076);
assign w37007 = (w26938 & w26937) | (w26938 & w27075) | (w26937 & w27075);
assign w37008 = (w26938 & w26937) | (w26938 & w36867) | (w26937 & w36867);
assign w37009 = (w26938 & w26937) | (w26938 & w36868) | (w26937 & w36868);
assign w37010 = (w26938 & w26937) | (w26938 & w36866) | (w26937 & w36866);
assign w37011 = (w26938 & w26937) | (w26938 & w36865) | (w26937 & w36865);
assign w37012 = (w26940 & w26939) | (w26940 & w27076) | (w26939 & w27076);
assign w37013 = (w26940 & w26939) | (w26940 & w27075) | (w26939 & w27075);
assign w37014 = (w26940 & w26939) | (w26940 & w36867) | (w26939 & w36867);
assign w37015 = (w26940 & w26939) | (w26940 & w36868) | (w26939 & w36868);
assign w37016 = (w26940 & w26939) | (w26940 & w36866) | (w26939 & w36866);
assign w37017 = (w26940 & w26939) | (w26940 & w36865) | (w26939 & w36865);
assign w37018 = w22107 & ~w26715;
assign w37019 = w22107 & w32125;
assign w37020 = b_44 & a_56;
assign w37021 = ~w21848 & w22055;
assign w37022 = (w26942 & w26941) | (w26942 & w27076) | (w26941 & w27076);
assign w37023 = (w26942 & w26941) | (w26942 & w27075) | (w26941 & w27075);
assign w37024 = (w26942 & w26941) | (w26942 & w36867) | (w26941 & w36867);
assign w37025 = (w26942 & w26941) | (w26942 & w36868) | (w26941 & w36868);
assign w37026 = (w26942 & w26941) | (w26942 & w36866) | (w26941 & w36866);
assign w37027 = (w26942 & w26941) | (w26942 & w36865) | (w26941 & w36865);
assign w37028 = ~w12641 & w22501;
assign w37029 = w22501 & ~w34715;
assign w37030 = w22501 & ~w34716;
assign w37031 = w22525 & w32284;
assign w37032 = w22525 & w32283;
assign w37033 = b_55 & a_47;
assign w37034 = (w26944 & w26943) | (w26944 & w27076) | (w26943 & w27076);
assign w37035 = (w26944 & w26943) | (w26944 & w27075) | (w26943 & w27075);
assign w37036 = (w26944 & w26943) | (w26944 & w36867) | (w26943 & w36867);
assign w37037 = (w26944 & w26943) | (w26944 & w36868) | (w26943 & w36868);
assign w37038 = (w26944 & w26943) | (w26944 & w36866) | (w26943 & w36866);
assign w37039 = (w26944 & w26943) | (w26944 & w36865) | (w26943 & w36865);
assign w37040 = (w26946 & w26945) | (w26946 & w27076) | (w26945 & w27076);
assign w37041 = (w26946 & w26945) | (w26946 & w27075) | (w26945 & w27075);
assign w37042 = (w26946 & w26945) | (w26946 & w36867) | (w26945 & w36867);
assign w37043 = (w26946 & w26945) | (w26946 & w36868) | (w26945 & w36868);
assign w37044 = (w26946 & w26945) | (w26946 & w36866) | (w26945 & w36866);
assign w37045 = (w26946 & w26945) | (w26946 & w36865) | (w26945 & w36865);
assign w37046 = w22598 & ~w22409;
assign w37047 = w22598 & w26052;
assign w37048 = ~w22372 & w22563;
assign w37049 = b_50 & a_53;
assign w37050 = ~w22432 & w22635;
assign w37051 = (w27087 & w27088) | (w27087 & w25176) | (w27088 & w25176);
assign w37052 = (w27087 & w27088) | (w27087 & w25177) | (w27088 & w25177);
assign w37053 = (w27087 & w27088) | (w27087 & w36806) | (w27088 & w36806);
assign w37054 = (w27087 & w27088) | (w27087 & w36807) | (w27088 & w36807);
assign w37055 = w22769 & w32336;
assign w37056 = w22769 & ~w22552;
assign w37057 = w22875 & ~w22894;
assign w37058 = ~w22875 & ~w22894;
assign w37059 = ~w22752 & w32332;
assign w37060 = ~w22752 & ~w22534;
assign w37061 = b_57 & a_47;
assign w37062 = w22815 & w32346;
assign w37063 = w22815 & ~w22624;
assign w37064 = ~w12641 & w22987;
assign w37065 = w22987 & ~w34715;
assign w37066 = w22987 & ~w34716;
assign w37067 = ~w22918 & w23099;
assign w37068 = b_51 & a_56;
assign w37069 = ~w12641 & w23420;
assign w37070 = w23420 & ~w34715;
assign w37071 = w23420 & ~w34716;
assign w37072 = w23446 & w32495;
assign w37073 = w23446 & w32496;
assign w37074 = ~w23446 & ~w32495;
assign w37075 = ~w23446 & ~w32496;
assign w37076 = b_49 & a_59;
assign w37077 = b_50 & a_59;
assign w37078 = b_48 & a_62;
assign w37079 = b_51 & a_59;
assign w37080 = ~w12641 & w23804;
assign w37081 = w23804 & ~w34715;
assign w37082 = w23804 & ~w34716;
assign w37083 = b_52 & a_59;
assign w37084 = (w26948 & w26947) | (w26948 & ~w27076) | (w26947 & ~w27076);
assign w37085 = (w26948 & w26947) | (w26948 & ~w27075) | (w26947 & ~w27075);
assign w37086 = (w26948 & w26947) | (w26948 & ~w36867) | (w26947 & ~w36867);
assign w37087 = (w26948 & w26947) | (w26948 & ~w36868) | (w26947 & ~w36868);
assign w37088 = b_56 & a_56;
assign w37089 = w23819 & ~w24011;
assign w37090 = ~w23819 & w24011;
assign w37091 = w12641 & w7616;
assign w37092 = w7616 & w34715;
assign w37093 = w7616 & w34716;
assign w37094 = w24146 & ~w24304;
assign w37095 = ~w24146 & w24304;
assign w37096 = b_57 & a_59;
assign w37097 = b_54 & a_62;
assign w37098 = w24295 & w32679;
assign w37099 = w24295 & ~w24198;
assign w37100 = w12641 & w8529;
assign w37101 = w8529 & w34715;
assign w37102 = w8529 & w34716;
assign w37103 = w12641 & w9537;
assign w37104 = w9537 & w34715;
assign w37105 = w9537 & w34716;
assign w37106 = w12641 & w10565;
assign w37107 = w10565 & w34715;
assign w37108 = w10565 & w34716;
assign w37109 = ~w12641 & w24923;
assign w37110 = (w26500 & w26501) | (w26500 & ~w26076) | (w26501 & ~w26076);
assign w37111 = (w26500 & w26501) | (w26500 & ~w26075) | (w26501 & ~w26075);
assign w37112 = (w26502 & w26503) | (w26502 & ~w26076) | (w26503 & ~w26076);
assign w37113 = (w26502 & w26503) | (w26502 & ~w26075) | (w26503 & ~w26075);
assign w37114 = (w26504 & w26505) | (w26504 & ~w26076) | (w26505 & ~w26076);
assign w37115 = (w26504 & w26505) | (w26504 & ~w26075) | (w26505 & ~w26075);
assign w37116 = (w26506 & w26507) | (w26506 & w26076) | (w26507 & w26076);
assign w37117 = (w26506 & w26507) | (w26506 & w26075) | (w26507 & w26075);
assign w37118 = ~w21779 & ~w21777;
assign w37119 = ~w23131 & w23544;
assign w37120 = w26510 & ~w23543;
assign w37121 = w26747 | w26746;
assign w37122 = w24314 & w24400;
assign w37123 = w26874 & ~w24399;
assign w37124 = (~w24399 & w26874) | (~w24399 & ~w24314) | (w26874 & ~w24314);
assign w37125 = w26982 | w26981;
assign w37126 = (w26981 & w26982) | (w26981 & w24314) | (w26982 & w24314);
assign w37127 = ~w24871 & ~w24905;
assign w37128 = ~w24932 & w24935;
assign w37129 = w25329 | w25328;
assign w37130 = w25333 | w25332;
assign w37131 = ~w14034 & w14021;
assign w37132 = w34954 & w16249;
assign w37133 = w20886 & w21142;
assign w37134 = ~w24548 & ~w24549;
assign w37135 = ~w24548 & ~w33042;
assign w37136 = ~w24548 & ~w33043;
assign w37137 = ~w24548 & ~w33044;
assign w37138 = (w25299 & w25300) | (w25299 & ~w24549) | (w25300 & ~w24549);
assign w37139 = (w25299 & w25300) | (w25299 & ~w33042) | (w25300 & ~w33042);
assign w37140 = (w25299 & w25300) | (w25299 & ~w33043) | (w25300 & ~w33043);
assign w37141 = (w25299 & w25300) | (w25299 & ~w33044) | (w25300 & ~w33044);
assign w37142 = (w25304 & w25303) | (w25304 & ~w24549) | (w25303 & ~w24549);
assign w37143 = (w25304 & w25303) | (w25304 & ~w33042) | (w25303 & ~w33042);
assign w37144 = (w25304 & w25303) | (w25304 & ~w33043) | (w25303 & ~w33043);
assign w37145 = (w25304 & w25303) | (w25304 & ~w33044) | (w25303 & ~w33044);
assign w37146 = (w25308 & w25307) | (w25308 & ~w24549) | (w25307 & ~w24549);
assign w37147 = (w25308 & w25307) | (w25308 & ~w33042) | (w25307 & ~w33042);
assign w37148 = (w25308 & w25307) | (w25308 & ~w33043) | (w25307 & ~w33043);
assign w37149 = (w25308 & w25307) | (w25308 & ~w33044) | (w25307 & ~w33044);
assign w37150 = (w25311 & w25312) | (w25311 & ~w24549) | (w25312 & ~w24549);
assign w37151 = (w25311 & w25312) | (w25311 & ~w33042) | (w25312 & ~w33042);
assign w37152 = (w25311 & w25312) | (w25311 & ~w33043) | (w25312 & ~w33043);
assign w37153 = (w25311 & w25312) | (w25311 & ~w33044) | (w25312 & ~w33044);
assign w37154 = w24980 & ~w24970;
assign w37155 = w24980 & w33076;
assign w37156 = ~w24980 & w24970;
assign w37157 = ~w24980 & ~w33076;
assign w37158 = ~w23909 & ~w33020;
assign w37159 = ~w23909 & ~w33021;
assign w37160 = ~w23909 & ~w23910;
assign w37161 = ~w23909 & ~w26980;
assign w37162 = (w25274 & w25275) | (w25274 & ~w33020) | (w25275 & ~w33020);
assign w37163 = (w25274 & w25275) | (w25274 & ~w33021) | (w25275 & ~w33021);
assign w37164 = (w25274 & w25275) | (w25274 & ~w23910) | (w25275 & ~w23910);
assign w37165 = (w25274 & w25275) | (w25274 & ~w26980) | (w25275 & ~w26980);
assign w37166 = (w25279 & w25278) | (w25279 & ~w33020) | (w25278 & ~w33020);
assign w37167 = (w25279 & w25278) | (w25279 & ~w33021) | (w25278 & ~w33021);
assign w37168 = (w25279 & w25278) | (w25279 & ~w23910) | (w25278 & ~w23910);
assign w37169 = (w25279 & w25278) | (w25279 & ~w26980) | (w25278 & ~w26980);
assign w37170 = (w25282 & w25283) | (w25282 & ~w33020) | (w25283 & ~w33020);
assign w37171 = (w25282 & w25283) | (w25282 & ~w33021) | (w25283 & ~w33021);
assign w37172 = (w25282 & w25283) | (w25282 & ~w23910) | (w25283 & ~w23910);
assign w37173 = (w25282 & w25283) | (w25282 & ~w26980) | (w25283 & ~w26980);
assign w37174 = (w25286 & w25287) | (w25286 & ~w33020) | (w25287 & ~w33020);
assign w37175 = (w25286 & w25287) | (w25286 & ~w33021) | (w25287 & ~w33021);
assign w37176 = (w25286 & w25287) | (w25286 & ~w23910) | (w25287 & ~w23910);
assign w37177 = (w25286 & w25287) | (w25286 & ~w26980) | (w25287 & ~w26980);
assign w37178 = (w25290 & w25291) | (w25290 & ~w33020) | (w25291 & ~w33020);
assign w37179 = (w25290 & w25291) | (w25290 & ~w33021) | (w25291 & ~w33021);
assign w37180 = (w25290 & w25291) | (w25290 & ~w23910) | (w25291 & ~w23910);
assign w37181 = (w25290 & w25291) | (w25290 & ~w26980) | (w25291 & ~w26980);
assign w37182 = (w25294 & w25295) | (w25294 & ~w33020) | (w25295 & ~w33020);
assign w37183 = (w25294 & w25295) | (w25294 & ~w33021) | (w25295 & ~w33021);
assign w37184 = (w25294 & w25295) | (w25294 & ~w23910) | (w25295 & ~w23910);
assign w37185 = (w25294 & w25295) | (w25294 & ~w26980) | (w25295 & ~w26980);
assign w37186 = (w25325 & w25326) | (w25325 & w24549) | (w25326 & w24549);
assign w37187 = (w25325 & w25326) | (w25325 & w33042) | (w25326 & w33042);
assign w37188 = (w25325 & w25326) | (w25325 & w33043) | (w25326 & w33043);
assign w37189 = (w25325 & w25326) | (w25325 & w33044) | (w25326 & w33044);
assign w37190 = w11906 & w11201;
assign w37191 = w11906 & w34663;
assign w37192 = w11211 & w11906;
assign w37193 = ~w11906 & ~w11201;
assign w37194 = ~w11906 & ~w34663;
assign w37195 = ~w11211 & ~w11906;
assign w37196 = (~w22978 & w25246) | (~w22978 & w32993) | (w25246 & w32993);
assign w37197 = (~w22978 & w25246) | (~w22978 & w32994) | (w25246 & w32994);
assign w37198 = (w25250 & w25249) | (w25250 & w32993) | (w25249 & w32993);
assign w37199 = (w25250 & w25249) | (w25250 & w32994) | (w25249 & w32994);
assign w37200 = ~w23126 & w25250;
assign w37201 = (w25254 & w25253) | (w25254 & w32993) | (w25253 & w32993);
assign w37202 = (w25254 & w25253) | (w25254 & w32994) | (w25253 & w32994);
assign w37203 = (w25258 & w25257) | (w25258 & w32993) | (w25257 & w32993);
assign w37204 = (w25258 & w25257) | (w25258 & w32994) | (w25257 & w32994);
assign w37205 = (w25262 & w25261) | (w25262 & w32993) | (w25261 & w32993);
assign w37206 = (w25262 & w25261) | (w25262 & w32994) | (w25261 & w32994);
assign w37207 = (w25266 & w25265) | (w25266 & w32993) | (w25265 & w32993);
assign w37208 = (w25266 & w25265) | (w25266 & w32994) | (w25265 & w32994);
assign w37209 = (w25270 & w25269) | (w25270 & w32993) | (w25269 & w32993);
assign w37210 = (w25270 & w25269) | (w25270 & w32994) | (w25269 & w32994);
assign w37211 = (w26076 & w26075) | (w26076 & ~w32993) | (w26075 & ~w32993);
assign w37212 = (w26076 & w26075) | (w26076 & ~w32994) | (w26075 & ~w32994);
assign w37213 = w3769 & w4023;
assign w37214 = ~w21779 & w32972;
assign w37215 = ~w21779 & w32971;
assign w37216 = ~w21779 & ~w21581;
assign w37217 = ~w21779 & w26870;
assign w37218 = w25225 & ~w21960;
assign w37219 = (~w21960 & w25225) | (~w21960 & ~w21777) | (w25225 & ~w21777);
assign w37220 = (~w21960 & w25225) | (~w21960 & w32976) | (w25225 & w32976);
assign w37221 = (~w21960 & w25225) | (~w21960 & w32977) | (w25225 & w32977);
assign w37222 = w25228 & w25229;
assign w37223 = (w25229 & w25228) | (w25229 & ~w21777) | (w25228 & ~w21777);
assign w37224 = (w25229 & w25228) | (w25229 & w32976) | (w25228 & w32976);
assign w37225 = (w25229 & w25228) | (w25229 & w32977) | (w25228 & w32977);
assign w37226 = w25232 & w25233;
assign w37227 = (w25233 & w25232) | (w25233 & ~w21777) | (w25232 & ~w21777);
assign w37228 = (w25233 & w25232) | (w25233 & w32976) | (w25232 & w32976);
assign w37229 = (w25233 & w25232) | (w25233 & w32977) | (w25232 & w32977);
assign w37230 = w25236 & w25237;
assign w37231 = (w25237 & w25236) | (w25237 & ~w21777) | (w25236 & ~w21777);
assign w37232 = (w25237 & w25236) | (w25237 & w32976) | (w25236 & w32976);
assign w37233 = (w25237 & w25236) | (w25237 & w32977) | (w25236 & w32977);
assign w37234 = w25240 & w25241;
assign w37235 = (w25241 & w25240) | (w25241 & ~w21777) | (w25240 & ~w21777);
assign w37236 = (w25241 & w25240) | (w25241 & w32976) | (w25240 & w32976);
assign w37237 = (w25241 & w25240) | (w25241 & w32977) | (w25240 & w32977);
assign w37238 = w26485 | w26484;
assign w37239 = (w26484 & w26485) | (w26484 & w21777) | (w26485 & w21777);
assign w37240 = (w26484 & w26485) | (w26484 & ~w32976) | (w26485 & ~w32976);
assign w37241 = (w26484 & w26485) | (w26484 & ~w32977) | (w26485 & ~w32977);
assign w37242 = ~w24021 & ~w24125;
assign w37243 = ~w24125 & ~w24022;
assign w37244 = ~w24124 & ~w24222;
assign w37245 = ~w24315 & w33025;
assign w37246 = ~w24315 & w33026;
assign w37247 = ~w24315 & w33027;
assign w37248 = ~w24400 & w33031;
assign w37249 = ~w24400 & w33032;
assign w37250 = ~w24400 & w33033;
assign w37251 = ~w24476 & w33037;
assign w37252 = ~w24476 & w33036;
assign w37253 = ~w24476 & ~w24399;
assign w37254 = ~w24476 & w26874;
assign w37255 = ~w24475 & ~w24549;
assign w37256 = ~w24549 & w33040;
assign w37257 = ~w24549 & w33041;
assign w37258 = w2908 & ~w2727;
assign w37259 = ~w20753 & ~w20754;
assign w37260 = ~w20753 & ~w26972;
assign w37261 = ~w20753 & ~w20305;
assign w37262 = ~w20753 & ~w32962;
assign w37263 = ~w20753 & ~w32963;
assign w37264 = ~w20753 & ~w32964;
assign w37265 = (w25212 & w25211) | (w25212 & ~w20754) | (w25211 & ~w20754);
assign w37266 = (w25212 & w25211) | (w25212 & ~w26972) | (w25211 & ~w26972);
assign w37267 = (w25212 & w25211) | (w25212 & ~w20305) | (w25211 & ~w20305);
assign w37268 = (w25212 & w25211) | (w25212 & ~w32962) | (w25211 & ~w32962);
assign w37269 = (w25212 & w25211) | (w25212 & ~w32963) | (w25211 & ~w32963);
assign w37270 = (w25212 & w25211) | (w25212 & ~w32964) | (w25211 & ~w32964);
assign w37271 = (w25215 & w25216) | (w25215 & ~w20754) | (w25216 & ~w20754);
assign w37272 = (w25215 & w25216) | (w25215 & ~w26972) | (w25216 & ~w26972);
assign w37273 = (w25215 & w25216) | (w25215 & ~w20305) | (w25216 & ~w20305);
assign w37274 = (w25215 & w25216) | (w25215 & ~w32962) | (w25216 & ~w32962);
assign w37275 = (w25215 & w25216) | (w25215 & ~w32963) | (w25216 & ~w32963);
assign w37276 = (w25215 & w25216) | (w25215 & ~w32964) | (w25216 & ~w32964);
assign w37277 = (w26719 & w26718) | (w26719 & ~w26972) | (w26718 & ~w26972);
assign w37278 = (w26719 & w26718) | (w26719 & ~w32964) | (w26718 & ~w32964);
assign w37279 = ~w23126 & ~w23272;
assign w37280 = ~w23413 & ~w23270;
assign w37281 = ~w23413 & w25488;
assign w37282 = ~w23413 & w32996;
assign w37283 = ~w23544 & w33002;
assign w37284 = ~w23544 & w33003;
assign w37285 = ~w23544 & w33001;
assign w37286 = ~w23544 & w33000;
assign w37287 = ~w23676 & w33010;
assign w37288 = ~w23676 & w33011;
assign w37289 = ~w23676 & w33009;
assign w37290 = ~w23676 & w33008;
assign w37291 = ~w23674 & ~w23798;
assign w37292 = ~w23798 & w33016;
assign w37293 = ~w23798 & w33017;
assign w37294 = ~w23910 & w26978;
assign w37295 = ~w23910 & w26979;
assign w37296 = ~w23796 & ~w23910;
assign w37297 = (w24619 & w25298) | (w24619 & w33365) | (w25298 & w33365);
assign w37298 = (w24619 & w25298) | (w24619 & w33364) | (w25298 & w33364);
assign w37299 = (w24619 & w25298) | (w24619 & w33363) | (w25298 & w33363);
assign w37300 = (w24619 & w25298) | (w24619 & w33362) | (w25298 & w33362);
assign w37301 = (w25301 & w25302) | (w25301 & w33365) | (w25302 & w33365);
assign w37302 = (w25301 & w25302) | (w25301 & w33364) | (w25302 & w33364);
assign w37303 = (w25301 & w25302) | (w25301 & w33363) | (w25302 & w33363);
assign w37304 = (w25301 & w25302) | (w25301 & w33362) | (w25302 & w33362);
assign w37305 = (w25305 & w25306) | (w25305 & w33365) | (w25306 & w33365);
assign w37306 = (w25305 & w25306) | (w25305 & w33364) | (w25306 & w33364);
assign w37307 = (w25305 & w25306) | (w25305 & w33363) | (w25306 & w33363);
assign w37308 = (w25305 & w25306) | (w25305 & w33362) | (w25306 & w33362);
assign w37309 = (w25309 & w25310) | (w25309 & w33365) | (w25310 & w33365);
assign w37310 = (w25309 & w25310) | (w25309 & w33364) | (w25310 & w33364);
assign w37311 = (w25309 & w25310) | (w25309 & w33363) | (w25310 & w33363);
assign w37312 = (w25309 & w25310) | (w25309 & w33362) | (w25310 & w33362);
assign w37313 = (w25313 & w25314) | (w25313 & w33365) | (w25314 & w33365);
assign w37314 = (w25313 & w25314) | (w25313 & w33364) | (w25314 & w33364);
assign w37315 = (w25313 & w25314) | (w25313 & w33363) | (w25314 & w33363);
assign w37316 = (w25313 & w25314) | (w25313 & w33362) | (w25314 & w33362);
assign w37317 = (w25318 & w25317) | (w25318 & w33365) | (w25317 & w33365);
assign w37318 = (w25318 & w25317) | (w25318 & w33364) | (w25317 & w33364);
assign w37319 = (w25318 & w25317) | (w25318 & w33363) | (w25317 & w33363);
assign w37320 = (w25318 & w25317) | (w25318 & w33362) | (w25317 & w33362);
assign w37321 = (w25322 & w25321) | (w25322 & w33365) | (w25321 & w33365);
assign w37322 = (w25322 & w25321) | (w25322 & w33364) | (w25321 & w33364);
assign w37323 = (w25322 & w25321) | (w25322 & w33363) | (w25321 & w33363);
assign w37324 = (w25322 & w25321) | (w25322 & w33362) | (w25321 & w33362);
assign w37325 = (w25716 & w25715) | (w25716 & w33365) | (w25715 & w33365);
assign w37326 = (w25716 & w25715) | (w25716 & w33364) | (w25715 & w33364);
assign w37327 = (w25716 & w25715) | (w25716 & w33363) | (w25715 & w33363);
assign w37328 = (w25716 & w25715) | (w25716 & w33362) | (w25715 & w33362);
assign w37329 = (w25718 & w25717) | (w25718 & w33365) | (w25717 & w33365);
assign w37330 = (w25718 & w25717) | (w25718 & w33364) | (w25717 & w33364);
assign w37331 = (w25718 & w25717) | (w25718 & w33363) | (w25717 & w33363);
assign w37332 = (w25718 & w25717) | (w25718 & w33362) | (w25717 & w33362);
assign w37333 = w7312 & ~w7750;
assign w37334 = ~w7529 & ~w7822;
assign w37335 = w5665 & w6056;
assign w37336 = w14190 & w14440;
assign w37337 = w14190 & ~w30187;
assign w37338 = w21197 & w21573;
assign w37339 = ~w1261 & ~w1508;
assign w37340 = w1356 & ~w1508;
assign w37341 = w7822 & w8126;
assign w37342 = w13694 & w13469;
assign w37343 = ~w14468 & ~w14065;
assign w37344 = ~w2604 & ~w2959;
assign w37345 = ~w2959 & w2793;
assign w37346 = w2604 & w2793;
assign w37347 = ~w9094 & w9115;
assign w37348 = w9115 & ~w8466;
assign w37349 = w9115 & w29168;
assign w37350 = w9094 & ~w9115;
assign w37351 = ~w9115 & w8466;
assign w37352 = ~w9115 & ~w29168;
assign w37353 = ~w9094 & ~w9115;
assign w37354 = ~w9115 & ~w8466;
assign w37355 = ~w9115 & w29168;
assign w37356 = w12651 & w12255;
assign w37357 = w12651 & w34698;
assign w37358 = w12242 & w12651;
assign w37359 = a_0 & w12641;
assign w37360 = a_62 & a_2;
assign w37361 = w13645 & w13519;
assign w37362 = w13989 & w13645;
assign w37363 = w13989 & w34789;
assign w37364 = w13631 & w13989;
assign w37365 = ~w14499 & w36469;
assign w37366 = ~w14499 & ~w14454;
assign w37367 = w14555 & ~w14432;
assign w37368 = w14555 & w14432;
assign w37369 = w14374 & w14356;
assign w37370 = ~w13893 & w14331;
assign w37371 = w14667 & w15083;
assign w37372 = ~w15843 & ~w15841;
assign w37373 = ~w15535 & ~w16162;
assign w37374 = ~w16238 & ~w16114;
assign w37375 = w16238 & w16114;
assign w37376 = w15672 & w16007;
assign w37377 = w16773 & ~w16263;
assign w37378 = w25158 | ~w16800;
assign w37379 = w25158 | w16803;
assign w37380 = w16559 & ~w27596;
assign w37381 = w36683 & ~w16848;
assign w37382 = ~w16848 & w36684;
assign w37383 = ~a_62 & w16912;
assign w37384 = a_62 & ~w16912;
assign w37385 = ~w16833 & ~w17057;
assign w37386 = ~w16782 & ~w17088;
assign w37387 = ~w17120 & w16799;
assign w37388 = ~w17120 & ~w30788;
assign w37389 = ~w16802 & ~w17120;
assign w37390 = w17172 & ~w36691;
assign w37391 = w17172 & ~w36690;
assign w37392 = ~w17172 & w36691;
assign w37393 = ~w17172 & w36690;
assign w37394 = w16742 & w16863;
assign w37395 = a_62 & w16912;
assign w37396 = w16692 & w16898;
assign w37397 = ~w17403 & w36696;
assign w37398 = w17417 & ~w25479;
assign w37399 = ~w25162 & w17417;
assign w37400 = ~w17417 & w25479;
assign w37401 = w25162 & ~w17417;
assign w37402 = w17473 & ~w36707;
assign w37403 = w17473 & ~w36708;
assign w37404 = ~w17473 & w36707;
assign w37405 = ~w17473 & w36708;
assign w37406 = w17346 & w16898;
assign w37407 = w17346 & w35118;
assign w37408 = w16698 & w17346;
assign w37409 = (~w17415 & w25164) | (~w17415 & ~w17118) | (w25164 & ~w17118);
assign w37410 = (~w17415 & w25164) | (~w17415 & w25479) | (w25164 & w25479);
assign w37411 = (~w17415 & w25164) | (~w17415 & w32936) | (w25164 & w32936);
assign w37412 = (~w17415 & w25164) | (~w17415 & w32937) | (w25164 & w32937);
assign w37413 = w25164 | ~w17415;
assign w37414 = (~w17415 & w25164) | (~w17415 & w25162) | (w25164 & w25162);
assign w37415 = w25165 & w17118;
assign w37416 = (w17118 & w25165) | (w17118 & w17711) | (w25165 & w17711);
assign w37417 = (w25165 & w25166) | (w25165 & w17118) | (w25166 & w17118);
assign w37418 = w25166 & w25165;
assign w37419 = (w25165 & w25166) | (w25165 & ~w25162) | (w25166 & ~w25162);
assign w37420 = ~w17711 & w37409;
assign w37421 = ~w17711 & w37410;
assign w37422 = ~w17748 & w36735;
assign w37423 = ~w17748 & w36736;
assign w37424 = w17748 & ~w36735;
assign w37425 = w17748 & ~w36736;
assign w37426 = ~w17990 & w25168;
assign w37427 = ~w17990 & w25167;
assign w37428 = (~w17989 & w25169) | (~w17989 & ~w17710) | (w25169 & ~w17710);
assign w37429 = (~w17989 & w25169) | (~w17989 & ~w17711) | (w25169 & ~w17711);
assign w37430 = (~w17989 & w25169) | (~w17989 & w25168) | (w25169 & w25168);
assign w37431 = w17652 & w17964;
assign w37432 = w17884 & w17866;
assign w37433 = ~w31132 & ~w17840;
assign w37434 = ~w31132 & ~w31057;
assign w37435 = w31132 & w17840;
assign w37436 = w31132 & w31057;
assign w37437 = w17551 & w17901;
assign w37438 = w17585 & w17926;
assign w37439 = (w25170 & w25171) | (w25170 & w17710) | (w25171 & w17710);
assign w37440 = (w25170 & w25171) | (w25170 & w17711) | (w25171 & w17711);
assign w37441 = (w25170 & w25171) | (w25170 & ~w25168) | (w25171 & ~w25168);
assign w37442 = (w25172 & w25173) | (w25172 & w25168) | (w25173 & w25168);
assign w37443 = (w25172 & w25173) | (w25172 & w25167) | (w25173 & w25167);
assign w37444 = (w25174 & w25175) | (w25174 & w17710) | (w25175 & w17710);
assign w37445 = (w25174 & w25175) | (w25174 & w17711) | (w25175 & w17711);
assign w37446 = (w25174 & w25175) | (w25174 & ~w25168) | (w25175 & ~w25168);
assign w37447 = ~w18271 & ~w18547;
assign w37448 = (w25176 & w25177) | (w25176 & w25168) | (w25177 & w25168);
assign w37449 = (w25176 & w25177) | (w25176 & w25167) | (w25177 & w25167);
assign w37450 = ~w18816 & w18545;
assign w37451 = ~w18816 & ~w32941;
assign w37452 = ~w18816 & ~w32942;
assign w37453 = ~w18816 & ~w36809;
assign w37454 = ~w18816 & ~w36808;
assign w37455 = ~w18816 & ~w25176;
assign w37456 = ~w18816 & ~w25177;
assign w37457 = ~w18815 & ~w18545;
assign w37458 = ~w18815 & w32941;
assign w37459 = ~w18815 & w32942;
assign w37460 = ~w18815 & w36809;
assign w37461 = ~w18815 & w36808;
assign w37462 = ~w18815 & w25176;
assign w37463 = ~w18815 & w25177;
assign w37464 = (~w18813 & w25178) | (~w18813 & ~w18545) | (w25178 & ~w18545);
assign w37465 = (~w18813 & w25178) | (~w18813 & w32941) | (w25178 & w32941);
assign w37466 = (~w18813 & w25178) | (~w18813 & w32942) | (w25178 & w32942);
assign w37467 = (~w18813 & w25178) | (~w18813 & w36809) | (w25178 & w36809);
assign w37468 = (~w18813 & w25178) | (~w18813 & w36808) | (w25178 & w36808);
assign w37469 = (~w18813 & w25178) | (~w18813 & w25176) | (w25178 & w25176);
assign w37470 = (~w18813 & w25178) | (~w18813 & w25177) | (w25178 & w25177);
assign w37471 = w18392 & w18715;
assign w37472 = (w25179 & w25180) | (w25179 & w18545) | (w25180 & w18545);
assign w37473 = (w25179 & w25180) | (w25179 & ~w32941) | (w25180 & ~w32941);
assign w37474 = (w25179 & w25180) | (w25179 & ~w32942) | (w25180 & ~w32942);
assign w37475 = (w25179 & w25180) | (w25179 & ~w36809) | (w25180 & ~w36809);
assign w37476 = (w25179 & w25180) | (w25179 & ~w36808) | (w25180 & ~w36808);
assign w37477 = (w25179 & w25180) | (w25179 & ~w25176) | (w25180 & ~w25176);
assign w37478 = (w25179 & w25180) | (w25179 & ~w25177) | (w25180 & ~w25177);
assign w37479 = ~w18966 & w19197;
assign w37480 = w18966 & ~w19197;
assign w37481 = (w25181 & w25182) | (w25181 & ~w18545) | (w25182 & ~w18545);
assign w37482 = (w25181 & w25182) | (w25181 & w32941) | (w25182 & w32941);
assign w37483 = (w25181 & w25182) | (w25181 & w32942) | (w25182 & w32942);
assign w37484 = (w25181 & w25182) | (w25181 & w36809) | (w25182 & w36809);
assign w37485 = (w25181 & w25182) | (w25181 & w36808) | (w25182 & w36808);
assign w37486 = (w25181 & w25182) | (w25181 & w25176) | (w25182 & w25176);
assign w37487 = (w25181 & w25182) | (w25181 & w25177) | (w25182 & w25177);
assign w37488 = (w25183 & w25184) | (w25183 & w18545) | (w25184 & w18545);
assign w37489 = (w25183 & w25184) | (w25183 & ~w32941) | (w25184 & ~w32941);
assign w37490 = (w25183 & w25184) | (w25183 & ~w32942) | (w25184 & ~w32942);
assign w37491 = (w25183 & w25184) | (w25183 & ~w36809) | (w25184 & ~w36809);
assign w37492 = (w25183 & w25184) | (w25183 & ~w36808) | (w25184 & ~w36808);
assign w37493 = (w25183 & w25184) | (w25183 & ~w25176) | (w25184 & ~w25176);
assign w37494 = (w25183 & w25184) | (w25183 & ~w25177) | (w25184 & ~w25177);
assign w37495 = (w25185 & w25186) | (w25185 & ~w18545) | (w25186 & ~w18545);
assign w37496 = (w25185 & w25186) | (w25185 & w32941) | (w25186 & w32941);
assign w37497 = (w25185 & w25186) | (w25185 & w32942) | (w25186 & w32942);
assign w37498 = (w25185 & w25186) | (w25185 & w36809) | (w25186 & w36809);
assign w37499 = (w25185 & w25186) | (w25185 & w36808) | (w25186 & w36808);
assign w37500 = (w25185 & w25186) | (w25185 & w25176) | (w25186 & w25176);
assign w37501 = (w25185 & w25186) | (w25185 & w25177) | (w25186 & w25177);
assign w37502 = (w25187 & w25188) | (w25187 & w18545) | (w25188 & w18545);
assign w37503 = (w25187 & w25188) | (w25187 & ~w32941) | (w25188 & ~w32941);
assign w37504 = (w25187 & w25188) | (w25187 & ~w32942) | (w25188 & ~w32942);
assign w37505 = (w25187 & w25188) | (w25187 & ~w36809) | (w25188 & ~w36809);
assign w37506 = (w25187 & w25188) | (w25187 & ~w36808) | (w25188 & ~w36808);
assign w37507 = (w25187 & w25188) | (w25187 & ~w25176) | (w25188 & ~w25176);
assign w37508 = (w25187 & w25188) | (w25187 & ~w25177) | (w25188 & ~w25177);
assign w37509 = (w27076 & w27075) | (w27076 & ~w17710) | (w27075 & ~w17710);
assign w37510 = (w27076 & w27075) | (w27076 & ~w17711) | (w27075 & ~w17711);
assign w37511 = (w27076 & w27075) | (w27076 & w25168) | (w27075 & w25168);
assign w37512 = w19298 & w19562;
assign w37513 = w19245 & w19403;
assign w37514 = w19479 & w19461;
assign w37515 = w19213 & w19498;
assign w37516 = ~w19831 & ~w33753;
assign w37517 = ~w19831 & ~w33755;
assign w37518 = ~w19831 & ~w33754;
assign w37519 = ~w19831 & ~w36870;
assign w37520 = ~w19831 & ~w36869;
assign w37521 = ~w19831 & ~w27076;
assign w37522 = ~w19831 & ~w27075;
assign w37523 = ~w19831 & ~w37510;
assign w37524 = ~w19831 & ~w37509;
assign w37525 = ~w19830 & w33753;
assign w37526 = ~w19830 & w33755;
assign w37527 = ~w19830 & w33754;
assign w37528 = ~w19830 & w36870;
assign w37529 = ~w19830 & w36869;
assign w37530 = ~w19830 & w27076;
assign w37531 = ~w19830 & w27075;
assign w37532 = ~w19830 & w37510;
assign w37533 = ~w19830 & w37509;
assign w37534 = w19785 & w19403;
assign w37535 = w19785 & w35429;
assign w37536 = w19404 & w19785;
assign w37537 = (w25192 & w25193) | (w25192 & ~w33753) | (w25193 & ~w33753);
assign w37538 = (w25192 & w25193) | (w25192 & ~w33755) | (w25193 & ~w33755);
assign w37539 = (w25192 & w25193) | (w25192 & ~w33754) | (w25193 & ~w33754);
assign w37540 = (w25192 & w25193) | (w25192 & ~w36870) | (w25193 & ~w36870);
assign w37541 = (w25192 & w25193) | (w25192 & ~w36869) | (w25193 & ~w36869);
assign w37542 = (w25192 & w25193) | (w25192 & ~w27076) | (w25193 & ~w27076);
assign w37543 = (w25192 & w25193) | (w25192 & ~w27075) | (w25193 & ~w27075);
assign w37544 = (w25192 & w25193) | (w25192 & ~w37510) | (w25193 & ~w37510);
assign w37545 = (w25192 & w25193) | (w25192 & ~w37509) | (w25193 & ~w37509);
assign w37546 = (w27077 & w27078) | (w27077 & ~w18545) | (w27078 & ~w18545);
assign w37547 = (w27077 & w27078) | (w27077 & w32941) | (w27078 & w32941);
assign w37548 = (w27077 & w27078) | (w27077 & w32942) | (w27078 & w32942);
assign w37549 = (w27077 & w27078) | (w27077 & w36809) | (w27078 & w36809);
assign w37550 = (w27077 & w27078) | (w27077 & w36808) | (w27078 & w36808);
assign w37551 = (w27077 & w27078) | (w27077 & w25176) | (w27078 & w25176);
assign w37552 = (w27077 & w27078) | (w27077 & w25177) | (w27078 & w25177);
assign w37553 = (w25196 & w25197) | (w25196 & ~w33753) | (w25197 & ~w33753);
assign w37554 = (w25196 & w25197) | (w25196 & ~w33755) | (w25197 & ~w33755);
assign w37555 = (w25196 & w25197) | (w25196 & ~w33754) | (w25197 & ~w33754);
assign w37556 = (w25196 & w25197) | (w25196 & ~w36870) | (w25197 & ~w36870);
assign w37557 = (w25196 & w25197) | (w25196 & ~w36869) | (w25197 & ~w36869);
assign w37558 = (w25196 & w25197) | (w25196 & ~w27076) | (w25197 & ~w27076);
assign w37559 = (w25196 & w25197) | (w25196 & ~w27075) | (w25197 & ~w27075);
assign w37560 = (w25196 & w25197) | (w25196 & ~w37510) | (w25197 & ~w37510);
assign w37561 = (w25196 & w25197) | (w25196 & ~w37509) | (w25197 & ~w37509);
assign w37562 = (w27079 & w27080) | (w27079 & ~w18545) | (w27080 & ~w18545);
assign w37563 = (w27079 & w27080) | (w27079 & w32941) | (w27080 & w32941);
assign w37564 = (w27079 & w27080) | (w27079 & w32942) | (w27080 & w32942);
assign w37565 = (w27079 & w27080) | (w27079 & w36809) | (w27080 & w36809);
assign w37566 = (w27079 & w27080) | (w27079 & w36808) | (w27080 & w36808);
assign w37567 = (w27079 & w27080) | (w27079 & w25176) | (w27080 & w25176);
assign w37568 = (w27079 & w27080) | (w27079 & w25177) | (w27080 & w25177);
assign w37569 = (w25198 & w25199) | (w25198 & w33753) | (w25199 & w33753);
assign w37570 = (w25198 & w25199) | (w25198 & w33755) | (w25199 & w33755);
assign w37571 = (w25198 & w25199) | (w25198 & w33754) | (w25199 & w33754);
assign w37572 = (w25198 & w25199) | (w25198 & w36870) | (w25199 & w36870);
assign w37573 = (w25198 & w25199) | (w25198 & w36869) | (w25199 & w36869);
assign w37574 = (w25198 & w25199) | (w25198 & w27076) | (w25199 & w27076);
assign w37575 = (w25198 & w25199) | (w25198 & w27075) | (w25199 & w27075);
assign w37576 = (w25198 & w25199) | (w25198 & w37510) | (w25199 & w37510);
assign w37577 = (w25198 & w25199) | (w25198 & w37509) | (w25199 & w37509);
assign w37578 = (w25200 & w25201) | (w25200 & ~w36870) | (w25201 & ~w36870);
assign w37579 = (w25200 & w25201) | (w25200 & ~w36869) | (w25201 & ~w36869);
assign w37580 = (w25200 & w25201) | (w25200 & ~w27076) | (w25201 & ~w27076);
assign w37581 = (w25200 & w25201) | (w25200 & ~w27075) | (w25201 & ~w27075);
assign w37582 = (w25200 & w25201) | (w25200 & ~w37510) | (w25201 & ~w37510);
assign w37583 = (w25200 & w25201) | (w25200 & ~w37509) | (w25201 & ~w37509);
assign w37584 = (w25202 & w25203) | (w25202 & w33753) | (w25203 & w33753);
assign w37585 = (w25202 & w25203) | (w25202 & w33755) | (w25203 & w33755);
assign w37586 = (w25202 & w25203) | (w25202 & w33754) | (w25203 & w33754);
assign w37587 = (w25202 & w25203) | (w25202 & w36870) | (w25203 & w36870);
assign w37588 = (w25202 & w25203) | (w25202 & w36869) | (w25203 & w36869);
assign w37589 = (w25202 & w25203) | (w25202 & w27076) | (w25203 & w27076);
assign w37590 = (w25202 & w25203) | (w25202 & w27075) | (w25203 & w27075);
assign w37591 = (w25202 & w25203) | (w25202 & w37510) | (w25203 & w37510);
assign w37592 = (w25202 & w25203) | (w25202 & w37509) | (w25203 & w37509);
assign w37593 = (w26932 & w26931) | (w26932 & w18545) | (w26931 & w18545);
assign w37594 = (w26932 & w26931) | (w26932 & ~w32941) | (w26931 & ~w32941);
assign w37595 = (w26932 & w26931) | (w26932 & ~w32942) | (w26931 & ~w32942);
assign w37596 = (w26932 & w26931) | (w26932 & ~w36809) | (w26931 & ~w36809);
assign w37597 = (w26932 & w26931) | (w26932 & ~w36808) | (w26931 & ~w36808);
assign w37598 = (w26932 & w26931) | (w26932 & ~w25176) | (w26931 & ~w25176);
assign w37599 = (w26932 & w26931) | (w26932 & ~w25177) | (w26931 & ~w25177);
assign w37600 = ~w20760 & ~w12641;
assign w37601 = ~w20760 & ~w34715;
assign w37602 = ~w20760 & ~w34716;
assign w37603 = (w27081 & w27082) | (w27081 & w36809) | (w27082 & w36809);
assign w37604 = (w27081 & w27082) | (w27081 & w36808) | (w27082 & w36808);
assign w37605 = (w27081 & w27082) | (w27081 & ~w18545) | (w27082 & ~w18545);
assign w37606 = (w27081 & w27082) | (w27081 & w32941) | (w27082 & w32941);
assign w37607 = (w27081 & w27082) | (w27081 & w32942) | (w27082 & w32942);
assign w37608 = w20636 & w20804;
assign w37609 = (w26934 & w26933) | (w26934 & w33753) | (w26933 & w33753);
assign w37610 = (w26934 & w26933) | (w26934 & w33755) | (w26933 & w33755);
assign w37611 = (w26934 & w26933) | (w26934 & w33754) | (w26933 & w33754);
assign w37612 = (w26934 & w26933) | (w26934 & w36870) | (w26933 & w36870);
assign w37613 = (w26934 & w26933) | (w26934 & w36869) | (w26933 & w36869);
assign w37614 = (w26934 & w26933) | (w26934 & w27076) | (w26933 & w27076);
assign w37615 = (w26934 & w26933) | (w26934 & w27075) | (w26933 & w27075);
assign w37616 = ~w7667 & w7579;
assign w37617 = w8008 & ~w8019;
assign w37618 = ~w11841 & w11851;
assign w37619 = w11841 & ~w11851;
assign w37620 = (w13389 & w26837) | (w13389 & ~w13021) | (w26837 & ~w13021);
assign w37621 = (w13389 & w26837) | (w13389 & w26663) | (w26837 & w26663);
assign w37622 = w26838 & w13021;
assign w37623 = w26838 & ~w26663;
assign w37624 = (w30447 & w30448) | (w30447 & ~w30277) | (w30448 & ~w30277);
assign w37625 = (w30528 & w30529) | (w30528 & ~w30277) | (w30529 & ~w30277);
assign w37626 = (w30618 & w30619) | (w30618 & ~w30277) | (w30619 & ~w30277);
assign w37627 = (w30700 & w30701) | (w30700 & ~w30277) | (w30701 & ~w30277);
assign w37628 = (w30793 & w30792) | (w30793 & ~w30277) | (w30792 & ~w30277);
assign w37629 = (w30875 & w30874) | (w30875 & ~w30277) | (w30874 & ~w30277);
assign w37630 = (w31087 & w31086) | (w31087 & ~w30277) | (w31086 & ~w30277);
assign w37631 = (w31166 & w31165) | (w31166 & ~w30277) | (w31165 & ~w30277);
assign w37632 = (w31240 & w31239) | (w31240 & ~w30277) | (w31239 & ~w30277);
assign w37633 = (w31308 & w31307) | (w31308 & ~w30277) | (w31307 & ~w30277);
assign w37634 = (w31310 & w31309) | (w31310 & ~w30277) | (w31309 & ~w30277);
assign w37635 = (w31439 & w31438) | (w31439 & ~w30277) | (w31438 & ~w30277);
assign w37636 = (w31512 & w31511) | (w31512 & ~w30277) | (w31511 & ~w30277);
assign w37637 = (w31574 & w31573) | (w31574 & ~w30277) | (w31573 & ~w30277);
assign w37638 = (w31631 & w31630) | (w31631 & ~w30277) | (w31630 & ~w30277);
assign w37639 = (w31696 & w31695) | (w31696 & ~w30277) | (w31695 & ~w30277);
assign w37640 = (w31698 & w31697) | (w31698 & ~w30277) | (w31697 & ~w30277);
assign w37641 = (w31812 & w31811) | (w31812 & ~w30277) | (w31811 & ~w30277);
assign w37642 = (w31814 & w31813) | (w31814 & w30277) | (w31813 & w30277);
assign w37643 = (w31814 & w31813) | (w31814 & w30278) | (w31813 & w30278);
assign w37644 = (w31870 & w31869) | (w31870 & ~w30277) | (w31869 & ~w30277);
assign w37645 = (w31931 & w31930) | (w31931 & ~w30277) | (w31930 & ~w30277);
assign w37646 = (w31933 & w31932) | (w31933 & ~w30277) | (w31932 & ~w30277);
assign w37647 = (w32039 & w32038) | (w32039 & ~w30277) | (w32038 & ~w30277);
assign w37648 = (w32090 & w32089) | (w32090 & ~w30277) | (w32089 & ~w30277);
assign w37649 = (w32092 & w32091) | (w32092 & ~w30277) | (w32091 & ~w30277);
assign w37650 = (w32194 & w32193) | (w32194 & ~w30277) | (w32193 & ~w30277);
assign w37651 = (w32196 & w32195) | (w32196 & ~w30277) | (w32195 & ~w30277);
assign w37652 = (w32241 & w32240) | (w32241 & ~w30277) | (w32240 & ~w30277);
assign w37653 = (w32311 & w32310) | (w32311 & ~w30277) | (w32310 & ~w30277);
assign w37654 = (w32313 & w32312) | (w32313 & ~w30277) | (w32312 & ~w30277);
assign w37655 = (w32350 & w32349) | (w32350 & ~w30277) | (w32349 & ~w30277);
assign w37656 = (w32599 & w32598) | (w32599 & w30277) | (w32598 & w30277);
assign w37657 = (w32599 & w32598) | (w32599 & w30278) | (w32598 & w30278);
assign w37658 = w13380 & w13367;
assign w37659 = w13380 & ~w26318;
assign w37660 = ~w13414 & ~w25140;
assign w37661 = (w13366 & w37862) | (w13366 & w37863) | (w37862 & w37863);
assign w37662 = w13428 & ~w13334;
assign w37663 = w13428 & w26319;
assign w37664 = ~w13428 & w13334;
assign w37665 = ~w13428 & ~w26319;
assign w37666 = (w13341 & w37864) | (w13341 & w37865) | (w37864 & w37865);
assign w37667 = w13341 & w37866;
assign w37668 = (~w13341 & w37867) | (~w13341 & w37868) | (w37867 & w37868);
assign w37669 = (~w13740 & ~w13341) | (~w13740 & w37869) | (~w13341 & w37869);
assign w37670 = (w25142 & w37870) | (w25142 & w37871) | (w37870 & w37871);
assign w37671 = (w30196 & w30197) | (w30196 & w25141) | (w30197 & w25141);
assign w37672 = (w30198 & w30199) | (w30198 & ~w13755) | (w30199 & ~w13755);
assign w37673 = (w30198 & w30199) | (w30198 & w25141) | (w30199 & w25141);
assign w37674 = (w30277 & w30278) | (w30277 & w13755) | (w30278 & w13755);
assign w37675 = (w30277 & w30278) | (w30277 & ~w25141) | (w30278 & ~w25141);
assign w37676 = ~w15504 & w37624;
assign w37677 = (~w30278 & w37872) | (~w30278 & w37873) | (w37872 & w37873);
assign w37678 = ~w15842 & w37625;
assign w37679 = (~w30278 & w37874) | (~w30278 & w37875) | (w37874 & w37875);
assign w37680 = ~w16172 & w37626;
assign w37681 = (~w30278 & w37876) | (~w30278 & w37877) | (w37876 & w37877);
assign w37682 = ~w16487 & w37627;
assign w37683 = (~w30278 & w37878) | (~w30278 & w37879) | (w37878 & w37879);
assign w37684 = ~w16801 & w37628;
assign w37685 = (~w30278 & w37880) | (~w30278 & w37881) | (w37880 & w37881);
assign w37686 = ~w17119 & w37629;
assign w37687 = (~w30278 & w37882) | (~w30278 & w37883) | (w37882 & w37883);
assign w37688 = w17990 & ~w37630;
assign w37689 = (w30278 & w37884) | (w30278 & w37885) | (w37884 & w37885);
assign w37690 = ~w18272 & w37631;
assign w37691 = (~w30278 & w37886) | (~w30278 & w37887) | (w37886 & w37887);
assign w37692 = ~w18546 & w37632;
assign w37693 = (~w30278 & w37888) | (~w30278 & w37889) | (w37888 & w37889);
assign w37694 = ~w18814 & w37633;
assign w37695 = (~w30278 & w37890) | (~w30278 & w37891) | (w37890 & w37891);
assign w37696 = ~w19079 & w37634;
assign w37697 = (~w30278 & w37892) | (~w30278 & w37893) | (w37892 & w37893);
assign w37698 = ~w19338 & w37635;
assign w37699 = (~w30278 & w37894) | (~w30278 & w37895) | (w37894 & w37895);
assign w37700 = ~w19582 & w37636;
assign w37701 = (~w30278 & w37896) | (~w30278 & w37897) | (w37896 & w37897);
assign w37702 = ~w19829 & w37637;
assign w37703 = (~w30278 & w37898) | (~w30278 & w37899) | (w37898 & w37899);
assign w37704 = ~w20072 & w37638;
assign w37705 = (~w30278 & w37900) | (~w30278 & w37901) | (w37900 & w37901);
assign w37706 = ~w20306 & w37639;
assign w37707 = (~w30278 & w37902) | (~w30278 & w37903) | (w37902 & w37903);
assign w37708 = ~w20535 & w37640;
assign w37709 = (~w30278 & w37904) | (~w30278 & w37905) | (w37904 & w37905);
assign w37710 = ~w20754 & w37641;
assign w37711 = (~w30278 & w37906) | (~w30278 & w37907) | (w37906 & w37907);
assign w37712 = (w20970 & w25206) | (w20970 & w37642) | (w25206 & w37642);
assign w37713 = (w30278 & w37908) | (w30278 & w37909) | (w37908 & w37909);
assign w37714 = (~w30278 & w37910) | (~w30278 & w37911) | (w37910 & w37911);
assign w37715 = ~w20970 & w37644;
assign w37716 = (w25209 & w25210) | (w25209 & w37642) | (w25210 & w37642);
assign w37717 = (w30278 & w37912) | (w30278 & w37913) | (w37912 & w37913);
assign w37718 = ~w21181 & w37645;
assign w37719 = (~w30278 & w37914) | (~w30278 & w37915) | (w37914 & w37915);
assign w37720 = (w25213 & w25214) | (w25213 & w37642) | (w25214 & w37642);
assign w37721 = (w30278 & w37916) | (w30278 & w37917) | (w37916 & w37917);
assign w37722 = ~w21389 & w37646;
assign w37723 = (~w30278 & w37918) | (~w30278 & w37919) | (w37918 & w37919);
assign w37724 = (w25217 & w25218) | (w25217 & w37642) | (w25218 & w37642);
assign w37725 = (w30278 & w37920) | (w30278 & w37921) | (w37920 & w37921);
assign w37726 = w21584 & w37647;
assign w37727 = (~w30278 & w37922) | (~w30278 & w37923) | (w37922 & w37923);
assign w37728 = (w25221 & w25222) | (w25221 & w37642) | (w25222 & w37642);
assign w37729 = (w30278 & w37924) | (w30278 & w37925) | (w37924 & w37925);
assign w37730 = ~w21778 & w37648;
assign w37731 = (~w30278 & w37926) | (~w30278 & w37927) | (w37926 & w37927);
assign w37732 = w21962 & ~w37649;
assign w37733 = (w30278 & w37928) | (w30278 & w37929) | (w37928 & w37929);
assign w37734 = ~w21962 & w37649;
assign w37735 = (~w30278 & w37930) | (~w30278 & w37931) | (w37930 & w37931);
assign w37736 = (w25226 & w25227) | (w25226 & ~w37649) | (w25227 & ~w37649);
assign w37737 = (w30278 & w37932) | (w30278 & w37933) | (w37932 & w37933);
assign w37738 = w22143 & w37650;
assign w37739 = (~w30278 & w37934) | (~w30278 & w37935) | (w37934 & w37935);
assign w37740 = (w25230 & w25231) | (w25230 & ~w37649) | (w25231 & ~w37649);
assign w37741 = (w30278 & w37936) | (w30278 & w37937) | (w37936 & w37937);
assign w37742 = ~w22321 & w37651;
assign w37743 = (~w30278 & w37938) | (~w30278 & w37939) | (w37938 & w37939);
assign w37744 = (w25234 & w25235) | (w25234 & ~w37649) | (w25235 & ~w37649);
assign w37745 = (w30278 & w37940) | (w30278 & w37941) | (w37940 & w37941);
assign w37746 = ~w22494 & w37652;
assign w37747 = (~w30278 & w37942) | (~w30278 & w37943) | (w37942 & w37943);
assign w37748 = (w25238 & w25239) | (w25238 & ~w37649) | (w25239 & ~w37649);
assign w37749 = (w30278 & w37944) | (w30278 & w37945) | (w37944 & w37945);
assign w37750 = ~w22662 & w37653;
assign w37751 = (~w30278 & w37946) | (~w30278 & w37947) | (w37946 & w37947);
assign w37752 = (w25242 & w25243) | (w25242 & ~w37649) | (w25243 & ~w37649);
assign w37753 = (w30278 & w37948) | (w30278 & w37949) | (w37948 & w37949);
assign w37754 = ~w22825 & w37654;
assign w37755 = (~w30278 & w37950) | (~w30278 & w37951) | (w37950 & w37951);
assign w37756 = w22980 & ~w37655;
assign w37757 = (w30278 & w37952) | (w30278 & w37953) | (w37952 & w37953);
assign w37758 = ~w22980 & w37655;
assign w37759 = (~w30278 & w37954) | (~w30278 & w37955) | (w37954 & w37955);
assign w37760 = (w25247 & w25248) | (w25247 & ~w37655) | (w25248 & ~w37655);
assign w37761 = (w30278 & w37956) | (w30278 & w37957) | (w37956 & w37957);
assign w37762 = (w27090 & w27089) | (w27090 & ~w37642) | (w27089 & ~w37642);
assign w37763 = (~w30278 & w37958) | (~w30278 & w37959) | (w37958 & w37959);
assign w37764 = (w25251 & w25252) | (w25251 & ~w37655) | (w25252 & ~w37655);
assign w37765 = (w30278 & w37960) | (w30278 & w37961) | (w37960 & w37961);
assign w37766 = (w27092 & w27091) | (w27092 & ~w37642) | (w27091 & ~w37642);
assign w37767 = (~w30278 & w37962) | (~w30278 & w37963) | (w37962 & w37963);
assign w37768 = (w25255 & w25256) | (w25255 & ~w37655) | (w25256 & ~w37655);
assign w37769 = (w30278 & w37964) | (w30278 & w37965) | (w37964 & w37965);
assign w37770 = (w27094 & w27093) | (w27094 & ~w37642) | (w27093 & ~w37642);
assign w37771 = (~w30278 & w37966) | (~w30278 & w37967) | (w37966 & w37967);
assign w37772 = (w25259 & w25260) | (w25259 & ~w37655) | (w25260 & ~w37655);
assign w37773 = (w30278 & w37968) | (w30278 & w37969) | (w37968 & w37969);
assign w37774 = (w27096 & w27095) | (w27096 & ~w37642) | (w27095 & ~w37642);
assign w37775 = (~w30278 & w37970) | (~w30278 & w37971) | (w37970 & w37971);
assign w37776 = (w25263 & w25264) | (w25263 & ~w37655) | (w25264 & ~w37655);
assign w37777 = (w30278 & w37972) | (w30278 & w37973) | (w37972 & w37973);
assign w37778 = (w27098 & w27097) | (w27098 & ~w37642) | (w27097 & ~w37642);
assign w37779 = (~w30278 & w37974) | (~w30278 & w37975) | (w37974 & w37975);
assign w37780 = (w25268 & w25267) | (w25268 & ~w37655) | (w25267 & ~w37655);
assign w37781 = (w30278 & w37976) | (w30278 & w37977) | (w37976 & w37977);
assign w37782 = (w27100 & w27099) | (w27100 & ~w37642) | (w27099 & ~w37642);
assign w37783 = (~w30278 & w37978) | (~w30278 & w37979) | (w37978 & w37979);
assign w37784 = (w27102 & w27101) | (w27102 & ~w37642) | (w27101 & ~w37642);
assign w37785 = (~w30278 & w37980) | (~w30278 & w37981) | (w37980 & w37981);
assign w37786 = (w24022 & w25273) | (w24022 & w37656) | (w25273 & w37656);
assign w37787 = (w30278 & w37982) | (w30278 & w37983) | (w37982 & w37983);
assign w37788 = (w26949 & w26950) | (w26949 & w37649) | (w26950 & w37649);
assign w37789 = (~w30278 & w37984) | (~w30278 & w37985) | (w37984 & w37985);
assign w37790 = (w25276 & w25277) | (w25276 & w37656) | (w25277 & w37656);
assign w37791 = (w30278 & w37986) | (w30278 & w37987) | (w37986 & w37987);
assign w37792 = (w26951 & w26952) | (w26951 & w37649) | (w26952 & w37649);
assign w37793 = (~w30278 & w37988) | (~w30278 & w37989) | (w37988 & w37989);
assign w37794 = (w25280 & w25281) | (w25280 & w37656) | (w25281 & w37656);
assign w37795 = (w30278 & w37990) | (w30278 & w37991) | (w37990 & w37991);
assign w37796 = (w26953 & w26954) | (w26953 & w37649) | (w26954 & w37649);
assign w37797 = (~w30278 & w37992) | (~w30278 & w37993) | (w37992 & w37993);
assign w37798 = (w25284 & w25285) | (w25284 & w37656) | (w25285 & w37656);
assign w37799 = (w30278 & w37994) | (w30278 & w37995) | (w37994 & w37995);
assign w37800 = (w26955 & w26956) | (w26955 & w37649) | (w26956 & w37649);
assign w37801 = (~w30278 & w37996) | (~w30278 & w37997) | (w37996 & w37997);
assign w37802 = (w25288 & w25289) | (w25288 & w37656) | (w25289 & w37656);
assign w37803 = (w30278 & w37998) | (w30278 & w37999) | (w37998 & w37999);
assign w37804 = (w26957 & w26958) | (w26957 & w37649) | (w26958 & w37649);
assign w37805 = (~w30278 & w38000) | (~w30278 & w38001) | (w38000 & w38001);
assign w37806 = (w25292 & w25293) | (w25292 & w37656) | (w25293 & w37656);
assign w37807 = (w30278 & w38002) | (w30278 & w38003) | (w38002 & w38003);
assign w37808 = (w26959 & w26960) | (w26959 & w37649) | (w26960 & w37649);
assign w37809 = (~w30278 & w38004) | (~w30278 & w38005) | (w38004 & w38005);
assign w37810 = (w26852 & w26853) | (w26852 & w37642) | (w26853 & w37642);
assign w37811 = (w30278 & w38006) | (w30278 & w38007) | (w38006 & w38007);
assign w37812 = (w26961 & w26962) | (w26961 & w37649) | (w26962 & w37649);
assign w37813 = (~w30278 & w38008) | (~w30278 & w38009) | (w38008 & w38009);
assign w37814 = (w27104 & w27103) | (w27104 & w37642) | (w27103 & w37642);
assign w37815 = (w30278 & w38010) | (w30278 & w38011) | (w38010 & w38011);
assign w37816 = (w26855 & w26854) | (w26855 & w37655) | (w26854 & w37655);
assign w37817 = (~w30278 & w38012) | (~w30278 & w38013) | (w38012 & w38013);
assign w37818 = (w27106 & w27105) | (w27106 & w37642) | (w27105 & w37642);
assign w37819 = (w30278 & w38014) | (w30278 & w38015) | (w38014 & w38015);
assign w37820 = (w26857 & w26856) | (w26857 & w37655) | (w26856 & w37655);
assign w37821 = (~w30278 & w38016) | (~w30278 & w38017) | (w38016 & w38017);
assign w37822 = (w27108 & w27107) | (w27108 & w37642) | (w27107 & w37642);
assign w37823 = (w30278 & w38018) | (w30278 & w38019) | (w38018 & w38019);
assign w37824 = (w26859 & w26858) | (w26859 & w37655) | (w26858 & w37655);
assign w37825 = (~w30278 & w38020) | (~w30278 & w38021) | (w38020 & w38021);
assign w37826 = (w27110 & w27109) | (w27110 & w37642) | (w27109 & w37642);
assign w37827 = (w30278 & w38022) | (w30278 & w38023) | (w38022 & w38023);
assign w37828 = (w26861 & w26860) | (w26861 & w37655) | (w26860 & w37655);
assign w37829 = (~w30278 & w38024) | (~w30278 & w38025) | (w38024 & w38025);
assign w37830 = (w27112 & w27111) | (w27112 & w37642) | (w27111 & w37642);
assign w37831 = (w30278 & w38026) | (w30278 & w38027) | (w38026 & w38027);
assign w37832 = (w26863 & w26862) | (w26863 & w37655) | (w26862 & w37655);
assign w37833 = (~w30278 & w38028) | (~w30278 & w38029) | (w38028 & w38029);
assign w37834 = (w27114 & w27113) | (w27114 & w37642) | (w27113 & w37642);
assign w37835 = (w30278 & w38030) | (w30278 & w38031) | (w38030 & w38031);
assign w37836 = (w26736 & w26735) | (w26736 & ~w37656) | (w26735 & ~w37656);
assign w37837 = (~w30278 & w38032) | (~w30278 & w38033) | (w38032 & w38033);
assign w37838 = (w27116 & w27115) | (w27116 & w37642) | (w27115 & w37642);
assign w37839 = (w30278 & w38034) | (w30278 & w38035) | (w38034 & w38035);
assign w37840 = (w26738 & w26737) | (w26738 & ~w37656) | (w26737 & ~w37656);
assign w37841 = (~w30278 & w38036) | (~w30278 & w38037) | (w38036 & w38037);
assign w37842 = (w26739 & w26740) | (w26739 & ~w37655) | (w26740 & ~w37655);
assign w37843 = (w30278 & w38038) | (w30278 & w38039) | (w38038 & w38039);
assign w37844 = (w27118 & w27117) | (w27118 & w37642) | (w27117 & w37642);
assign w37845 = (w30278 & w38040) | (w30278 & w38041) | (w38040 & w38041);
assign w37846 = (w32872 & w32873) | (w32872 & ~w37642) | (w32873 & ~w37642);
assign w37847 = (~w30278 & w38042) | (~w30278 & w38043) | (w38042 & w38043);
assign w37848 = (w27120 & w27119) | (w27120 & w37642) | (w27119 & w37642);
assign w37849 = (w30278 & w38044) | (w30278 & w38045) | (w38044 & w38045);
assign w37850 = (w32880 & w32881) | (w32880 & ~w37642) | (w32881 & ~w37642);
assign w37851 = (~w30278 & w38046) | (~w30278 & w38047) | (w38046 & w38047);
assign w37852 = (w32884 & w32885) | (w32884 & ~w37642) | (w32885 & ~w37642);
assign w37853 = (~w30278 & w38048) | (~w30278 & w38049) | (w38048 & w38049);
assign w37854 = (w32886 & w32887) | (w32886 & w37642) | (w32887 & w37642);
assign w37855 = (w30278 & w38050) | (w30278 & w38051) | (w38050 & w38051);
assign w37856 = (w26079 & w26080) | (w26079 & ~w37656) | (w26080 & ~w37656);
assign w37857 = (~w30278 & w38052) | (~w30278 & w38053) | (w38052 & w38053);
assign w37858 = ~w13718 & ~w13327;
assign w37859 = ~w13718 & w26662;
assign w37860 = (w35275 & w35276) | (w35275 & ~w33965) | (w35276 & ~w33965);
assign w37861 = (w35275 & w35276) | (w35275 & ~w33966) | (w35276 & ~w33966);
assign w37862 = ~w13414 & ~w13367;
assign w37863 = ~w13414 & w26318;
assign w37864 = ~w13740 & ~w13364;
assign w37865 = ~w13740 & ~w33434;
assign w37866 = ~w13351 & ~w13740;
assign w37867 = ~w13740 & w13364;
assign w37868 = ~w13740 & w33434;
assign w37869 = w13351 & ~w13740;
assign w37870 = w30196 & ~w13755;
assign w37871 = (~w13755 & w30196) | (~w13755 & ~w14482) | (w30196 & ~w14482);
assign w37872 = ~w15504 & w30447;
assign w37873 = ~w15504 & w30448;
assign w37874 = ~w15842 & w30528;
assign w37875 = ~w15842 & w30529;
assign w37876 = ~w16172 & w30618;
assign w37877 = ~w16172 & w30619;
assign w37878 = ~w16487 & w30700;
assign w37879 = ~w16487 & w30701;
assign w37880 = ~w16801 & w30793;
assign w37881 = ~w16801 & w30792;
assign w37882 = ~w17119 & w30875;
assign w37883 = ~w17119 & w30874;
assign w37884 = w17990 & ~w31087;
assign w37885 = w17990 & ~w31086;
assign w37886 = ~w18272 & w31166;
assign w37887 = ~w18272 & w31165;
assign w37888 = ~w18546 & w31240;
assign w37889 = ~w18546 & w31239;
assign w37890 = ~w18814 & w31308;
assign w37891 = ~w18814 & w31307;
assign w37892 = ~w19079 & w31310;
assign w37893 = ~w19079 & w31309;
assign w37894 = ~w19338 & w31439;
assign w37895 = ~w19338 & w31438;
assign w37896 = ~w19582 & w31512;
assign w37897 = ~w19582 & w31511;
assign w37898 = ~w19829 & w31574;
assign w37899 = ~w19829 & w31573;
assign w37900 = ~w20072 & w31631;
assign w37901 = ~w20072 & w31630;
assign w37902 = ~w20306 & w31696;
assign w37903 = ~w20306 & w31695;
assign w37904 = ~w20535 & w31698;
assign w37905 = ~w20535 & w31697;
assign w37906 = ~w20754 & w31812;
assign w37907 = ~w20754 & w31811;
assign w37908 = (w20970 & w25206) | (w20970 & w31814) | (w25206 & w31814);
assign w37909 = (w20970 & w25206) | (w20970 & w31813) | (w25206 & w31813);
assign w37910 = ~w20970 & w31870;
assign w37911 = ~w20970 & w31869;
assign w37912 = (w25209 & w25210) | (w25209 & w31814) | (w25210 & w31814);
assign w37913 = (w25209 & w25210) | (w25209 & w31813) | (w25210 & w31813);
assign w37914 = ~w21181 & w31931;
assign w37915 = ~w21181 & w31930;
assign w37916 = (w25213 & w25214) | (w25213 & w31814) | (w25214 & w31814);
assign w37917 = (w25213 & w25214) | (w25213 & w31813) | (w25214 & w31813);
assign w37918 = ~w21389 & w31933;
assign w37919 = ~w21389 & w31932;
assign w37920 = (w25217 & w25218) | (w25217 & w31814) | (w25218 & w31814);
assign w37921 = (w25217 & w25218) | (w25217 & w31813) | (w25218 & w31813);
assign w37922 = w21584 & w32039;
assign w37923 = w21584 & w32038;
assign w37924 = (w25221 & w25222) | (w25221 & w31814) | (w25222 & w31814);
assign w37925 = (w25221 & w25222) | (w25221 & w31813) | (w25222 & w31813);
assign w37926 = ~w21778 & w32090;
assign w37927 = ~w21778 & w32089;
assign w37928 = w21962 & ~w32092;
assign w37929 = w21962 & ~w32091;
assign w37930 = ~w21962 & w32092;
assign w37931 = ~w21962 & w32091;
assign w37932 = (w25226 & w25227) | (w25226 & ~w32092) | (w25227 & ~w32092);
assign w37933 = (w25226 & w25227) | (w25226 & ~w32091) | (w25227 & ~w32091);
assign w37934 = w22143 & w32194;
assign w37935 = w22143 & w32193;
assign w37936 = (w25230 & w25231) | (w25230 & ~w32092) | (w25231 & ~w32092);
assign w37937 = (w25230 & w25231) | (w25230 & ~w32091) | (w25231 & ~w32091);
assign w37938 = ~w22321 & w32196;
assign w37939 = ~w22321 & w32195;
assign w37940 = (w25234 & w25235) | (w25234 & ~w32092) | (w25235 & ~w32092);
assign w37941 = (w25234 & w25235) | (w25234 & ~w32091) | (w25235 & ~w32091);
assign w37942 = ~w22494 & w32241;
assign w37943 = ~w22494 & w32240;
assign w37944 = (w25238 & w25239) | (w25238 & ~w32092) | (w25239 & ~w32092);
assign w37945 = (w25238 & w25239) | (w25238 & ~w32091) | (w25239 & ~w32091);
assign w37946 = ~w22662 & w32311;
assign w37947 = ~w22662 & w32310;
assign w37948 = (w25242 & w25243) | (w25242 & ~w32092) | (w25243 & ~w32092);
assign w37949 = (w25242 & w25243) | (w25242 & ~w32091) | (w25243 & ~w32091);
assign w37950 = ~w22825 & w32313;
assign w37951 = ~w22825 & w32312;
assign w37952 = w22980 & ~w32350;
assign w37953 = w22980 & ~w32349;
assign w37954 = ~w22980 & w32350;
assign w37955 = ~w22980 & w32349;
assign w37956 = (w25247 & w25248) | (w25247 & ~w32350) | (w25248 & ~w32350);
assign w37957 = (w25247 & w25248) | (w25247 & ~w32349) | (w25248 & ~w32349);
assign w37958 = (w27090 & w27089) | (w27090 & ~w31814) | (w27089 & ~w31814);
assign w37959 = (w27090 & w27089) | (w27090 & ~w31813) | (w27089 & ~w31813);
assign w37960 = (w25251 & w25252) | (w25251 & ~w32350) | (w25252 & ~w32350);
assign w37961 = (w25251 & w25252) | (w25251 & ~w32349) | (w25252 & ~w32349);
assign w37962 = (w27092 & w27091) | (w27092 & ~w31814) | (w27091 & ~w31814);
assign w37963 = (w27092 & w27091) | (w27092 & ~w31813) | (w27091 & ~w31813);
assign w37964 = (w25255 & w25256) | (w25255 & ~w32350) | (w25256 & ~w32350);
assign w37965 = (w25255 & w25256) | (w25255 & ~w32349) | (w25256 & ~w32349);
assign w37966 = (w27094 & w27093) | (w27094 & ~w31814) | (w27093 & ~w31814);
assign w37967 = (w27094 & w27093) | (w27094 & ~w31813) | (w27093 & ~w31813);
assign w37968 = (w25259 & w25260) | (w25259 & ~w32350) | (w25260 & ~w32350);
assign w37969 = (w25259 & w25260) | (w25259 & ~w32349) | (w25260 & ~w32349);
assign w37970 = (w27096 & w27095) | (w27096 & ~w31814) | (w27095 & ~w31814);
assign w37971 = (w27096 & w27095) | (w27096 & ~w31813) | (w27095 & ~w31813);
assign w37972 = (w25263 & w25264) | (w25263 & ~w32350) | (w25264 & ~w32350);
assign w37973 = (w25263 & w25264) | (w25263 & ~w32349) | (w25264 & ~w32349);
assign w37974 = (w27098 & w27097) | (w27098 & ~w31814) | (w27097 & ~w31814);
assign w37975 = (w27098 & w27097) | (w27098 & ~w31813) | (w27097 & ~w31813);
assign w37976 = (w25268 & w25267) | (w25268 & ~w32350) | (w25267 & ~w32350);
assign w37977 = (w25268 & w25267) | (w25268 & ~w32349) | (w25267 & ~w32349);
assign w37978 = (w27100 & w27099) | (w27100 & ~w31814) | (w27099 & ~w31814);
assign w37979 = (w27100 & w27099) | (w27100 & ~w31813) | (w27099 & ~w31813);
assign w37980 = (w27102 & w27101) | (w27102 & ~w31814) | (w27101 & ~w31814);
assign w37981 = (w27102 & w27101) | (w27102 & ~w31813) | (w27101 & ~w31813);
assign w37982 = (w24022 & w25273) | (w24022 & w32599) | (w25273 & w32599);
assign w37983 = (w24022 & w25273) | (w24022 & w32598) | (w25273 & w32598);
assign w37984 = (w26949 & w26950) | (w26949 & w32092) | (w26950 & w32092);
assign w37985 = (w26949 & w26950) | (w26949 & w32091) | (w26950 & w32091);
assign w37986 = (w25276 & w25277) | (w25276 & w32599) | (w25277 & w32599);
assign w37987 = (w25276 & w25277) | (w25276 & w32598) | (w25277 & w32598);
assign w37988 = (w26951 & w26952) | (w26951 & w32092) | (w26952 & w32092);
assign w37989 = (w26951 & w26952) | (w26951 & w32091) | (w26952 & w32091);
assign w37990 = (w25280 & w25281) | (w25280 & w32599) | (w25281 & w32599);
assign w37991 = (w25280 & w25281) | (w25280 & w32598) | (w25281 & w32598);
assign w37992 = (w26953 & w26954) | (w26953 & w32092) | (w26954 & w32092);
assign w37993 = (w26953 & w26954) | (w26953 & w32091) | (w26954 & w32091);
assign w37994 = (w25284 & w25285) | (w25284 & w32599) | (w25285 & w32599);
assign w37995 = (w25284 & w25285) | (w25284 & w32598) | (w25285 & w32598);
assign w37996 = (w26955 & w26956) | (w26955 & w32092) | (w26956 & w32092);
assign w37997 = (w26955 & w26956) | (w26955 & w32091) | (w26956 & w32091);
assign w37998 = (w25288 & w25289) | (w25288 & w32599) | (w25289 & w32599);
assign w37999 = (w25288 & w25289) | (w25288 & w32598) | (w25289 & w32598);
assign w38000 = (w26957 & w26958) | (w26957 & w32092) | (w26958 & w32092);
assign w38001 = (w26957 & w26958) | (w26957 & w32091) | (w26958 & w32091);
assign w38002 = (w25292 & w25293) | (w25292 & w32599) | (w25293 & w32599);
assign w38003 = (w25292 & w25293) | (w25292 & w32598) | (w25293 & w32598);
assign w38004 = (w26959 & w26960) | (w26959 & w32092) | (w26960 & w32092);
assign w38005 = (w26959 & w26960) | (w26959 & w32091) | (w26960 & w32091);
assign w38006 = (w26852 & w26853) | (w26852 & w31814) | (w26853 & w31814);
assign w38007 = (w26852 & w26853) | (w26852 & w31813) | (w26853 & w31813);
assign w38008 = (w26961 & w26962) | (w26961 & w32092) | (w26962 & w32092);
assign w38009 = (w26961 & w26962) | (w26961 & w32091) | (w26962 & w32091);
assign w38010 = (w27104 & w27103) | (w27104 & w31814) | (w27103 & w31814);
assign w38011 = (w27104 & w27103) | (w27104 & w31813) | (w27103 & w31813);
assign w38012 = (w26855 & w26854) | (w26855 & w32350) | (w26854 & w32350);
assign w38013 = (w26855 & w26854) | (w26855 & w32349) | (w26854 & w32349);
assign w38014 = (w27106 & w27105) | (w27106 & w31814) | (w27105 & w31814);
assign w38015 = (w27106 & w27105) | (w27106 & w31813) | (w27105 & w31813);
assign w38016 = (w26857 & w26856) | (w26857 & w32350) | (w26856 & w32350);
assign w38017 = (w26857 & w26856) | (w26857 & w32349) | (w26856 & w32349);
assign w38018 = (w27108 & w27107) | (w27108 & w31814) | (w27107 & w31814);
assign w38019 = (w27108 & w27107) | (w27108 & w31813) | (w27107 & w31813);
assign w38020 = (w26859 & w26858) | (w26859 & w32350) | (w26858 & w32350);
assign w38021 = (w26859 & w26858) | (w26859 & w32349) | (w26858 & w32349);
assign w38022 = (w27110 & w27109) | (w27110 & w31814) | (w27109 & w31814);
assign w38023 = (w27110 & w27109) | (w27110 & w31813) | (w27109 & w31813);
assign w38024 = (w26861 & w26860) | (w26861 & w32350) | (w26860 & w32350);
assign w38025 = (w26861 & w26860) | (w26861 & w32349) | (w26860 & w32349);
assign w38026 = (w27112 & w27111) | (w27112 & w31814) | (w27111 & w31814);
assign w38027 = (w27112 & w27111) | (w27112 & w31813) | (w27111 & w31813);
assign w38028 = (w26863 & w26862) | (w26863 & w32350) | (w26862 & w32350);
assign w38029 = (w26863 & w26862) | (w26863 & w32349) | (w26862 & w32349);
assign w38030 = (w27114 & w27113) | (w27114 & w31814) | (w27113 & w31814);
assign w38031 = (w27114 & w27113) | (w27114 & w31813) | (w27113 & w31813);
assign w38032 = (w26736 & w26735) | (w26736 & ~w32599) | (w26735 & ~w32599);
assign w38033 = (w26736 & w26735) | (w26736 & ~w32598) | (w26735 & ~w32598);
assign w38034 = (w27116 & w27115) | (w27116 & w31814) | (w27115 & w31814);
assign w38035 = (w27116 & w27115) | (w27116 & w31813) | (w27115 & w31813);
assign w38036 = (w26738 & w26737) | (w26738 & ~w32599) | (w26737 & ~w32599);
assign w38037 = (w26738 & w26737) | (w26738 & ~w32598) | (w26737 & ~w32598);
assign w38038 = (w26739 & w26740) | (w26739 & ~w32350) | (w26740 & ~w32350);
assign w38039 = (w26739 & w26740) | (w26739 & ~w32349) | (w26740 & ~w32349);
assign w38040 = (w27118 & w27117) | (w27118 & w31814) | (w27117 & w31814);
assign w38041 = (w27118 & w27117) | (w27118 & w31813) | (w27117 & w31813);
assign w38042 = (w32872 & w32873) | (w32872 & ~w31814) | (w32873 & ~w31814);
assign w38043 = (w32872 & w32873) | (w32872 & ~w31813) | (w32873 & ~w31813);
assign w38044 = (w27120 & w27119) | (w27120 & w31814) | (w27119 & w31814);
assign w38045 = (w27120 & w27119) | (w27120 & w31813) | (w27119 & w31813);
assign w38046 = (w32880 & w32881) | (w32880 & ~w31814) | (w32881 & ~w31814);
assign w38047 = (w32880 & w32881) | (w32880 & ~w31813) | (w32881 & ~w31813);
assign w38048 = (w32884 & w32885) | (w32884 & ~w31814) | (w32885 & ~w31814);
assign w38049 = (w32884 & w32885) | (w32884 & ~w31813) | (w32885 & ~w31813);
assign w38050 = (w32886 & w32887) | (w32886 & w31814) | (w32887 & w31814);
assign w38051 = (w32886 & w32887) | (w32886 & w31813) | (w32887 & w31813);
assign w38052 = (w26079 & w26080) | (w26079 & ~w32599) | (w26080 & ~w32599);
assign w38053 = (w26079 & w26080) | (w26079 & ~w32598) | (w26080 & ~w32598);
assign w38054 = ~w13414 & w25140;
assign w38055 = ~w13414 & ~w13369;
assign w38056 = w26670 & ~w13390;
assign w38057 = (~w13390 & w26670) | (~w13390 & ~w13383) | (w26670 & ~w13383);
assign w38058 = (~w13755 & w25141) | (~w13755 & w12665) | (w25141 & w12665);
assign w38059 = (~w13755 & w25141) | (~w13755 & w27785) | (w25141 & w27785);
assign w38060 = ~w14079 & w13719;
assign w38061 = ~w14079 & ~w27566;
assign w38062 = ~w14079 & ~w13719;
assign w38063 = ~w14079 & w27566;
assign w38064 = (w30113 & w30114) | (w30113 & w12665) | (w30114 & w12665);
assign w38065 = (w30113 & w30114) | (w30113 & w27785) | (w30114 & w27785);
assign w38066 = ~w14136 & ~w27796;
assign w38067 = ~w14136 & ~w27797;
assign w38068 = w14139 & w14476;
assign w38069 = ~w14139 & ~w14476;
assign w38070 = ~w14482 & ~w14480;
assign w38071 = ~w27326 & a_2;
assign w38072 = w61 & w66;
assign w38073 = ~w61 & ~w66;
assign w38074 = ~w12 & w27391;
assign w38075 = a_2 & ~w27852;
assign w38076 = a_2 & ~w123;
assign w38077 = a_2 & w27852;
assign w38078 = a_2 & w123;
assign w38079 = a_2 & ~w27855;
assign w38080 = a_2 & ~w184;
assign w38081 = a_2 & w27855;
assign w38082 = a_2 & w184;
assign w38083 = a_2 & ~w27860;
assign w38084 = a_2 & ~w207;
assign w38085 = a_2 & w27860;
assign w38086 = a_2 & w207;
assign w38087 = ~w27014 & a_5;
assign w38088 = ~w306 & w27865;
assign w38089 = ~w306 & w27864;
assign w38090 = w308 & w303;
assign w38091 = w27867 & a_2;
assign w38092 = (a_2 & w27867) | (a_2 & ~w308) | (w27867 & ~w308);
assign w38093 = w308 & w27868;
assign w38094 = a_5 & ~w27870;
assign w38095 = a_5 & ~w326;
assign w38096 = a_5 & w27870;
assign w38097 = a_5 & w326;
assign w38098 = a_2 & ~w27874;
assign w38099 = a_2 & ~w365;
assign w38100 = a_2 & w27874;
assign w38101 = a_2 & w365;
assign w38102 = a_5 & ~w27876;
assign w38103 = a_5 & ~w390;
assign w38104 = a_5 & w27876;
assign w38105 = a_5 & w390;
assign w38106 = a_2 & ~w27884;
assign w38107 = a_2 & ~w448;
assign w38108 = a_2 & w27884;
assign w38109 = a_2 & w448;
assign w38110 = w308 & w472;
assign w38111 = w27888 & a_5;
assign w38112 = (a_5 & w27888) | (a_5 & ~w308) | (w27888 & ~w308);
assign w38113 = ~w26763 & a_8;
assign w38114 = a_2 & ~w27896;
assign w38115 = a_2 & ~w524;
assign w38116 = a_2 & w27896;
assign w38117 = a_2 & w524;
assign w38118 = a_2 & ~w27901;
assign w38119 = a_2 & ~w546;
assign w38120 = a_2 & w27901;
assign w38121 = a_2 & w546;
assign w38122 = a_8 & ~w27903;
assign w38123 = a_8 & ~w562;
assign w38124 = a_8 & w27903;
assign w38125 = a_8 & w562;
assign w38126 = a_5 & ~w27905;
assign w38127 = a_5 & ~w601;
assign w38128 = a_5 & w27905;
assign w38129 = a_5 & w601;
assign w38130 = a_8 & ~w27907;
assign w38131 = a_8 & ~w629;
assign w38132 = a_8 & w27907;
assign w38133 = a_8 & w629;
assign w38134 = a_5 & ~w27912;
assign w38135 = a_5 & ~w687;
assign w38136 = a_5 & w27912;
assign w38137 = a_5 & w687;
assign w38138 = a_2 & ~w27915;
assign w38139 = a_2 & ~w704;
assign w38140 = a_2 & w27915;
assign w38141 = a_2 & w704;
assign w38142 = a_2 & ~w27920;
assign w38143 = a_2 & ~w729;
assign w38144 = a_2 & w27920;
assign w38145 = a_2 & w729;
assign w38146 = a_5 & ~w27922;
assign w38147 = a_5 & ~w745;
assign w38148 = a_5 & w27922;
assign w38149 = a_5 & w745;
assign w38150 = ~w26886 & a_11;
assign w38151 = w308 & w790;
assign w38152 = w27926 & a_8;
assign w38153 = (a_8 & w27926) | (a_8 & ~w308) | (w27926 & ~w308);
assign w38154 = a_2 & ~w27934;
assign w38155 = a_2 & ~w821;
assign w38156 = a_2 & w27934;
assign w38157 = a_2 & w821;
assign w38158 = a_5 & ~w27937;
assign w38159 = a_5 & ~w838;
assign w38160 = a_5 & w27937;
assign w38161 = a_5 & w838;
assign w38162 = a_8 & ~w27939;
assign w38163 = a_8 & ~w849;
assign w38164 = a_8 & w27939;
assign w38165 = a_8 & w849;
assign w38166 = a_11 & ~w27941;
assign w38167 = a_11 & ~w859;
assign w38168 = a_11 & w27941;
assign w38169 = a_11 & w859;
assign w38170 = w923 & ~w27944;
assign w38171 = w923 & ~w27945;
assign w38172 = ~w923 & w27944;
assign w38173 = ~w923 & w27945;
assign w38174 = a_2 & ~w27946;
assign w38175 = a_2 & ~w920;
assign w38176 = a_2 & w27946;
assign w38177 = a_2 & w920;
assign w38178 = a_5 & ~w27949;
assign w38179 = a_5 & ~w937;
assign w38180 = a_5 & w27949;
assign w38181 = a_5 & w937;
assign w38182 = a_8 & ~w27951;
assign w38183 = a_8 & ~w947;
assign w38184 = a_8 & w27951;
assign w38185 = a_8 & w947;
assign w38186 = a_11 & ~w27953;
assign w38187 = a_11 & ~w958;
assign w38188 = a_11 & w27953;
assign w38189 = a_11 & w958;
assign w38190 = (w27960 & w27961) | (w27960 & ~w27944) | (w27961 & ~w27944);
assign w38191 = (w27960 & w27961) | (w27960 & ~w27945) | (w27961 & ~w27945);
assign w38192 = (w27962 & w27963) | (w27962 & w27944) | (w27963 & w27944);
assign w38193 = (w27962 & w27963) | (w27962 & w27945) | (w27963 & w27945);
assign w38194 = a_2 & ~w27964;
assign w38195 = a_2 & ~w1032;
assign w38196 = a_2 & w27964;
assign w38197 = a_2 & w1032;
assign w38198 = a_5 & ~w27966;
assign w38199 = a_5 & ~w1049;
assign w38200 = a_5 & w27966;
assign w38201 = a_5 & w1049;
assign w38202 = a_8 & ~w27968;
assign w38203 = a_8 & ~w1060;
assign w38204 = a_8 & w27968;
assign w38205 = a_8 & w1060;
assign w38206 = ~w26768 & a_14;
assign w38207 = w308 & w1105;
assign w38208 = w27972 & a_11;
assign w38209 = (a_11 & w27972) | (a_11 & ~w308) | (w27972 & ~w308);
assign w38210 = a_5 & ~w27975;
assign w38211 = a_5 & ~w1144;
assign w38212 = a_5 & w27975;
assign w38213 = a_5 & w1144;
assign w38214 = a_8 & ~w27977;
assign w38215 = a_8 & ~w1155;
assign w38216 = a_8 & w27977;
assign w38217 = a_8 & w1155;
assign w38218 = a_14 & ~w27980;
assign w38219 = a_14 & ~w1166;
assign w38220 = a_14 & w27980;
assign w38221 = a_14 & w1166;
assign w38222 = a_11 & ~w27982;
assign w38223 = a_11 & ~w1204;
assign w38224 = a_11 & w27982;
assign w38225 = a_11 & w1204;
assign w38226 = (w27987 & w27988) | (w27987 & ~w27944) | (w27988 & ~w27944);
assign w38227 = (w27987 & w27988) | (w27987 & ~w27945) | (w27988 & ~w27945);
assign w38228 = (w27989 & w27990) | (w27989 & w27944) | (w27990 & w27944);
assign w38229 = (w27989 & w27990) | (w27989 & w27945) | (w27990 & w27945);
assign w38230 = a_2 & ~w27991;
assign w38231 = a_2 & ~w1232;
assign w38232 = a_2 & w27991;
assign w38233 = a_2 & w1232;
assign w38234 = a_5 & ~w27993;
assign w38235 = a_5 & ~w1256;
assign w38236 = a_5 & w27993;
assign w38237 = a_5 & w1256;
assign w38238 = a_14 & ~w27995;
assign w38239 = a_14 & ~w1267;
assign w38240 = a_14 & w27995;
assign w38241 = a_14 & w1267;
assign w38242 = a_11 & ~w28000;
assign w38243 = a_11 & ~w1323;
assign w38244 = a_11 & w28000;
assign w38245 = a_11 & w1323;
assign w38246 = a_8 & ~w28002;
assign w38247 = a_8 & ~w1341;
assign w38248 = a_8 & w28002;
assign w38249 = a_8 & w1341;
assign w38250 = (w28008 & w28007) | (w28008 & ~w27944) | (w28007 & ~w27944);
assign w38251 = (w28008 & w28007) | (w28008 & ~w27945) | (w28007 & ~w27945);
assign w38252 = (w28010 & w28009) | (w28010 & w27944) | (w28009 & w27944);
assign w38253 = (w28010 & w28009) | (w28010 & w27945) | (w28009 & w27945);
assign w38254 = a_2 & ~w1366;
assign w38255 = a_2 & ~w28011;
assign w38256 = a_2 & w1366;
assign w38257 = a_2 & w28011;
assign w38258 = a_5 & ~w28013;
assign w38259 = a_5 & ~w1391;
assign w38260 = a_5 & w28013;
assign w38261 = a_5 & w1391;
assign w38262 = a_8 & ~w28015;
assign w38263 = a_8 & ~w1401;
assign w38264 = a_8 & w28015;
assign w38265 = a_8 & w1401;
assign w38266 = a_11 & ~w28017;
assign w38267 = a_11 & ~w1412;
assign w38268 = a_11 & w28017;
assign w38269 = a_11 & w1412;
assign w38270 = ~w26770 & a_17;
assign w38271 = w308 & w1458;
assign w38272 = w28021 & a_14;
assign w38273 = (a_14 & w28021) | (a_14 & ~w308) | (w28021 & ~w308);
assign w38274 = (w1500 & w28025) | (w1500 & w38251) | (w28025 & w38251);
assign w38275 = (w1500 & w28025) | (w1500 & w38250) | (w28025 & w38250);
assign w38276 = w28026 & ~w38251;
assign w38277 = w28026 & ~w38250;
assign w38278 = a_2 & ~w28027;
assign w38279 = a_2 & ~w1497;
assign w38280 = a_2 & w28027;
assign w38281 = a_2 & w1497;
assign w38282 = ~w27731 & ~w1508;
assign w38283 = a_8 & ~w28030;
assign w38284 = a_8 & ~w1522;
assign w38285 = a_8 & w28030;
assign w38286 = a_8 & w1522;
assign w38287 = a_11 & ~w28032;
assign w38288 = a_11 & ~w1533;
assign w38289 = a_11 & w28032;
assign w38290 = a_11 & w1533;
assign w38291 = a_17 & ~w28035;
assign w38292 = a_17 & ~w1544;
assign w38293 = a_17 & w28035;
assign w38294 = a_17 & w1544;
assign w38295 = a_14 & ~w28037;
assign w38296 = a_14 & ~w1582;
assign w38297 = a_14 & w28037;
assign w38298 = a_14 & w1582;
assign w38299 = a_5 & ~w28039;
assign w38300 = a_5 & ~w1610;
assign w38301 = a_5 & w28039;
assign w38302 = a_5 & w1610;
assign w38303 = (w28045 & w28044) | (w28045 & w38251) | (w28044 & w38251);
assign w38304 = (w28045 & w28044) | (w28045 & w38250) | (w28044 & w38250);
assign w38305 = (w28047 & w28046) | (w28047 & ~w38251) | (w28046 & ~w38251);
assign w38306 = (w28047 & w28046) | (w28047 & ~w38250) | (w28046 & ~w38250);
assign w38307 = a_2 & ~w28048;
assign w38308 = a_2 & ~w1628;
assign w38309 = a_2 & w28048;
assign w38310 = a_2 & w1628;
assign w38311 = a_8 & ~w28051;
assign w38312 = a_8 & ~w1654;
assign w38313 = a_8 & w28051;
assign w38314 = a_8 & w1654;
assign w38315 = a_17 & ~w28054;
assign w38316 = a_17 & ~w1666;
assign w38317 = a_17 & w28054;
assign w38318 = a_17 & w1666;
assign w38319 = a_14 & ~w28059;
assign w38320 = a_14 & ~w1722;
assign w38321 = a_14 & w28059;
assign w38322 = a_14 & w1722;
assign w38323 = a_11 & ~w28061;
assign w38324 = a_11 & ~w1740;
assign w38325 = a_11 & w28061;
assign w38326 = a_11 & w1740;
assign w38327 = a_5 & ~w28063;
assign w38328 = a_5 & ~w1762;
assign w38329 = a_5 & w28063;
assign w38330 = a_5 & w1762;
assign w38331 = (w28069 & w28068) | (w28069 & w38251) | (w28068 & w38251);
assign w38332 = (w28069 & w28068) | (w28069 & w38250) | (w28068 & w38250);
assign w38333 = (w28071 & w28070) | (w28071 & ~w38251) | (w28070 & ~w38251);
assign w38334 = (w28071 & w28070) | (w28071 & ~w38250) | (w28070 & ~w38250);
assign w38335 = a_2 & ~w28072;
assign w38336 = a_2 & ~w1780;
assign w38337 = a_2 & w28072;
assign w38338 = a_2 & w1780;
assign w38339 = a_8 & ~w28075;
assign w38340 = a_8 & ~w1803;
assign w38341 = a_8 & w28075;
assign w38342 = a_8 & w1803;
assign w38343 = a_11 & ~w28077;
assign w38344 = a_11 & ~w1813;
assign w38345 = a_11 & w28077;
assign w38346 = a_11 & w1813;
assign w38347 = a_14 & ~w28079;
assign w38348 = a_14 & ~w1824;
assign w38349 = a_14 & w28079;
assign w38350 = a_14 & w1824;
assign w38351 = ~w26773 & a_20;
assign w38352 = w308 & w1870;
assign w38353 = w28083 & a_17;
assign w38354 = (a_17 & w28083) | (a_17 & ~w308) | (w28083 & ~w308);
assign w38355 = a_5 & ~w28088;
assign w38356 = a_5 & ~w1909;
assign w38357 = a_5 & w28088;
assign w38358 = a_5 & w1909;
assign w38359 = (w28093 & w28092) | (w28093 & w38251) | (w28092 & w38251);
assign w38360 = (w28093 & w28092) | (w28093 & w38250) | (w28092 & w38250);
assign w38361 = (w28094 & w28095) | (w28094 & ~w38251) | (w28095 & ~w38251);
assign w38362 = (w28094 & w28095) | (w28094 & ~w38250) | (w28095 & ~w38250);
assign w38363 = a_2 & ~w28096;
assign w38364 = a_2 & ~w1927;
assign w38365 = a_2 & w28096;
assign w38366 = a_2 & w1927;
assign w38367 = a_5 & ~w28099;
assign w38368 = a_5 & ~w1952;
assign w38369 = a_5 & w28099;
assign w38370 = a_5 & w1952;
assign w38371 = a_11 & ~w28101;
assign w38372 = a_11 & ~w1963;
assign w38373 = a_11 & w28101;
assign w38374 = a_11 & w1963;
assign w38375 = a_14 & ~w28103;
assign w38376 = a_14 & ~w1974;
assign w38377 = a_14 & w28103;
assign w38378 = a_14 & w1974;
assign w38379 = a_20 & ~w28106;
assign w38380 = a_20 & ~w1985;
assign w38381 = a_20 & w28106;
assign w38382 = a_20 & w1985;
assign w38383 = a_17 & ~w28108;
assign w38384 = a_17 & ~w2023;
assign w38385 = a_17 & w28108;
assign w38386 = a_17 & w2023;
assign w38387 = a_8 & ~w28110;
assign w38388 = a_8 & ~w2053;
assign w38389 = a_8 & w28110;
assign w38390 = a_8 & w2053;
assign w38391 = a_2 & ~w28115;
assign w38392 = a_2 & ~w2077;
assign w38393 = a_2 & w28115;
assign w38394 = a_2 & w2077;
assign w38395 = w2070 & ~w2088;
assign w38396 = ~w2070 & ~w2088;
assign w38397 = a_2 & ~w28125;
assign w38398 = a_2 & ~w2102;
assign w38399 = a_2 & w28125;
assign w38400 = a_2 & w2102;
assign w38401 = w1947 & ~w2065;
assign w38402 = a_11 & ~w28127;
assign w38403 = a_11 & ~w2119;
assign w38404 = a_11 & w28127;
assign w38405 = a_11 & w2119;
assign w38406 = a_20 & ~w28129;
assign w38407 = a_20 & ~w2130;
assign w38408 = a_20 & w28129;
assign w38409 = a_20 & w2130;
assign w38410 = a_17 & ~w28134;
assign w38411 = a_17 & ~w2186;
assign w38412 = a_17 & w28134;
assign w38413 = a_17 & w2186;
assign w38414 = a_14 & ~w28136;
assign w38415 = a_14 & ~w2204;
assign w38416 = a_14 & w28136;
assign w38417 = a_14 & w2204;
assign w38418 = a_8 & ~w28139;
assign w38419 = a_8 & ~w2229;
assign w38420 = a_8 & w28139;
assign w38421 = a_8 & w2229;
assign w38422 = a_5 & ~w28141;
assign w38423 = a_5 & ~w2247;
assign w38424 = a_5 & w28141;
assign w38425 = a_5 & w2247;
assign w38426 = w2261 & w2089;
assign w38427 = w2261 & ~w2092;
assign w38428 = ~w2261 & ~w2089;
assign w38429 = ~w2261 & w2092;
assign w38430 = a_14 & ~w28148;
assign w38431 = a_14 & ~w2274;
assign w38432 = a_14 & w28148;
assign w38433 = a_14 & w2274;
assign w38434 = a_17 & ~w28150;
assign w38435 = a_17 & ~w2284;
assign w38436 = a_17 & w28150;
assign w38437 = a_17 & w2284;
assign w38438 = ~w28153 & a_23;
assign w38439 = w308 & w2329;
assign w38440 = w28159 & a_20;
assign w38441 = (a_20 & w28159) | (a_20 & ~w308) | (w28159 & ~w308);
assign w38442 = a_11 & ~w28165;
assign w38443 = a_11 & ~w2359;
assign w38444 = a_11 & w28165;
assign w38445 = a_11 & w2359;
assign w38446 = a_8 & ~w28167;
assign w38447 = a_8 & ~w2375;
assign w38448 = a_8 & w28167;
assign w38449 = a_8 & w2375;
assign w38450 = a_5 & ~w28169;
assign w38451 = a_5 & ~w2393;
assign w38452 = a_5 & w28169;
assign w38453 = a_5 & w2393;
assign w38454 = a_2 & ~w28178;
assign w38455 = a_2 & ~w2410;
assign w38456 = a_2 & w28178;
assign w38457 = a_2 & w2410;
assign w38458 = ~w2424 & ~w2422;
assign w38459 = a_5 & ~w28180;
assign w38460 = a_5 & ~w2433;
assign w38461 = a_5 & w28180;
assign w38462 = a_5 & w2433;
assign w38463 = a_14 & ~w28182;
assign w38464 = a_14 & ~w2443;
assign w38465 = a_14 & w28182;
assign w38466 = a_14 & w2443;
assign w38467 = a_17 & ~w28184;
assign w38468 = a_17 & ~w2454;
assign w38469 = a_17 & w28184;
assign w38470 = a_17 & w2454;
assign w38471 = a_23 & ~w28186;
assign w38472 = a_23 & ~w2465;
assign w38473 = a_23 & w28186;
assign w38474 = a_23 & w2465;
assign w38475 = a_20 & ~w28188;
assign w38476 = a_20 & ~w2503;
assign w38477 = a_20 & w28188;
assign w38478 = a_20 & w2503;
assign w38479 = a_8 & ~w28195;
assign w38480 = a_8 & ~w2551;
assign w38481 = a_8 & w28195;
assign w38482 = a_8 & w2551;
assign w38483 = a_2 & ~w28204;
assign w38484 = a_2 & ~w2576;
assign w38485 = a_2 & w28204;
assign w38486 = a_2 & w2576;
assign w38487 = a_5 & ~w28207;
assign w38488 = a_5 & ~w2599;
assign w38489 = a_5 & w28207;
assign w38490 = a_5 & w2599;
assign w38491 = a_23 & ~w28210;
assign w38492 = a_23 & ~w2611;
assign w38493 = a_23 & w28210;
assign w38494 = a_23 & w2611;
assign w38495 = a_20 & ~w28213;
assign w38496 = a_20 & ~w2667;
assign w38497 = a_20 & w28213;
assign w38498 = a_20 & w2667;
assign w38499 = a_8 & ~w28233;
assign w38500 = a_8 & ~w2740;
assign w38501 = a_8 & w28233;
assign w38502 = a_8 & w2740;
assign w38503 = w2568 & ~w2564;
assign w38504 = w2768 & ~w28238;
assign w38505 = w2768 & ~w28237;
assign w38506 = ~w2768 & w28238;
assign w38507 = ~w2768 & w28237;
assign w38508 = a_2 & ~w28239;
assign w38509 = a_2 & ~w2765;
assign w38510 = a_2 & w28239;
assign w38511 = a_2 & w2765;
assign w38512 = a_5 & ~w28242;
assign w38513 = a_5 & ~w2788;
assign w38514 = a_5 & w28242;
assign w38515 = a_5 & w2788;
assign w38516 = a_17 & ~w28244;
assign w38517 = a_17 & ~w2799;
assign w38518 = a_17 & w28244;
assign w38519 = a_17 & w2799;
assign w38520 = a_20 & ~w28246;
assign w38521 = a_20 & ~w2810;
assign w38522 = a_20 & w28246;
assign w38523 = a_20 & w2810;
assign w38524 = ~w26129 & a_26;
assign w38525 = w308 & w2856;
assign w38526 = w28249 & a_23;
assign w38527 = (a_23 & w28249) | (a_23 & ~w308) | (w28249 & ~w308);
assign w38528 = a_11 & ~w28258;
assign w38529 = a_11 & ~w2905;
assign w38530 = a_11 & w28258;
assign w38531 = a_11 & w2905;
assign w38532 = a_8 & ~w28263;
assign w38533 = a_8 & ~w2922;
assign w38534 = a_8 & w28263;
assign w38535 = a_8 & w2922;
assign w38536 = (w28269 & w28270) | (w28269 & ~w28238) | (w28270 & ~w28238);
assign w38537 = (w28269 & w28270) | (w28269 & ~w28237) | (w28270 & ~w28237);
assign w38538 = (w28271 & w28272) | (w28271 & w28238) | (w28272 & w28238);
assign w38539 = (w28271 & w28272) | (w28271 & w28237) | (w28272 & w28237);
assign w38540 = a_2 & ~w28273;
assign w38541 = a_2 & ~w2948;
assign w38542 = a_2 & w28273;
assign w38543 = a_2 & w2948;
assign w38544 = ~w28274 & ~w2959;
assign w38545 = ~w2779 & ~w2778;
assign w38546 = a_17 & ~w28276;
assign w38547 = a_17 & ~w2973;
assign w38548 = a_17 & w28276;
assign w38549 = a_17 & w2973;
assign w38550 = a_20 & ~w28278;
assign w38551 = a_20 & ~w2984;
assign w38552 = a_20 & w28278;
assign w38553 = a_20 & w2984;
assign w38554 = a_26 & ~w28281;
assign w38555 = a_26 & ~w2995;
assign w38556 = a_26 & w28281;
assign w38557 = a_26 & w2995;
assign w38558 = a_23 & ~w28283;
assign w38559 = a_23 & ~w3033;
assign w38560 = a_23 & w28283;
assign w38561 = a_23 & w3033;
assign w38562 = a_11 & ~w28291;
assign w38563 = a_11 & ~w3081;
assign w38564 = a_11 & w28291;
assign w38565 = a_11 & w3081;
assign w38566 = a_8 & ~w28293;
assign w38567 = a_8 & ~w3098;
assign w38568 = a_8 & w28293;
assign w38569 = a_8 & w3098;
assign w38570 = a_5 & ~w28295;
assign w38571 = a_5 & ~w3114;
assign w38572 = a_5 & w28295;
assign w38573 = a_5 & w3114;
assign w38574 = (w28301 & w28302) | (w28301 & ~w28238) | (w28302 & ~w28238);
assign w38575 = (w28301 & w28302) | (w28301 & ~w28237) | (w28302 & ~w28237);
assign w38576 = (w28303 & w28304) | (w28303 & w28238) | (w28304 & w28238);
assign w38577 = (w28303 & w28304) | (w28303 & w28237) | (w28304 & w28237);
assign w38578 = a_2 & ~w28305;
assign w38579 = a_2 & ~w3132;
assign w38580 = a_2 & w28305;
assign w38581 = a_2 & w3132;
assign w38582 = a_17 & ~w28308;
assign w38583 = a_17 & ~w3156;
assign w38584 = a_17 & w28308;
assign w38585 = a_17 & w3156;
assign w38586 = a_26 & ~w28310;
assign w38587 = a_26 & ~w3167;
assign w38588 = a_26 & w28310;
assign w38589 = a_26 & w3167;
assign w38590 = a_23 & ~w28315;
assign w38591 = a_23 & ~w28316;
assign w38592 = a_20 & ~w28318;
assign w38593 = a_20 & ~w3241;
assign w38594 = a_20 & w28318;
assign w38595 = a_20 & w3241;
assign w38596 = a_8 & ~w28331;
assign w38597 = a_8 & ~w3303;
assign w38598 = a_8 & w28331;
assign w38599 = a_8 & w3303;
assign w38600 = a_5 & ~w28334;
assign w38601 = a_5 & ~w3321;
assign w38602 = a_5 & w28334;
assign w38603 = a_5 & w3321;
assign w38604 = w3124 & ~w3120;
assign w38605 = (w28339 & w28338) | (w28339 & ~w28238) | (w28338 & ~w28238);
assign w38606 = (w28339 & w28338) | (w28339 & ~w28237) | (w28338 & ~w28237);
assign w38607 = (w28341 & w28340) | (w28341 & w28238) | (w28340 & w28238);
assign w38608 = (w28341 & w28340) | (w28341 & w28237) | (w28340 & w28237);
assign w38609 = a_2 & ~w3339;
assign w38610 = a_2 & ~w28342;
assign w38611 = a_2 & w3339;
assign w38612 = a_2 & w28342;
assign w38613 = w3148 & ~w3144;
assign w38614 = w3355 & ~w3351;
assign w38615 = w3331 & ~w3327;
assign w38616 = a_8 & ~w28344;
assign w38617 = a_8 & ~w3365;
assign w38618 = a_8 & w28344;
assign w38619 = a_8 & w3365;
assign w38620 = a_17 & ~w28346;
assign w38621 = a_17 & ~w3377;
assign w38622 = a_17 & w28346;
assign w38623 = a_17 & w3377;
assign w38624 = ~w26540 & a_29;
assign w38625 = w308 & w3424;
assign w38626 = w28349 & a_26;
assign w38627 = (a_26 & w28349) | (a_26 & ~w308) | (w28349 & ~w308);
assign w38628 = a_23 & ~w28355;
assign w38629 = a_23 & ~w3443;
assign w38630 = a_23 & w28355;
assign w38631 = a_23 & w3443;
assign w38632 = a_20 & ~w28358;
assign w38633 = a_20 & ~w3459;
assign w38634 = a_20 & w28358;
assign w38635 = a_20 & w3459;
assign w38636 = a_14 & ~w28362;
assign w38637 = a_14 & ~w3483;
assign w38638 = a_14 & w28362;
assign w38639 = a_14 & w3483;
assign w38640 = w3506 & w3290;
assign w38641 = w3506 & ~w25014;
assign w38642 = ~w3506 & ~w3290;
assign w38643 = ~w3506 & w25014;
assign w38644 = a_5 & ~w28371;
assign w38645 = a_5 & ~w3522;
assign w38646 = a_5 & w28371;
assign w38647 = a_5 & w3522;
assign w38648 = (w28377 & w28378) | (w28377 & ~w28238) | (w28378 & ~w28238);
assign w38649 = (w28377 & w28378) | (w28377 & ~w28237) | (w28378 & ~w28237);
assign w38650 = (w28379 & w28380) | (w28379 & w28238) | (w28380 & w28238);
assign w38651 = (w28379 & w28380) | (w28379 & w28237) | (w28380 & w28237);
assign w38652 = a_2 & ~w28381;
assign w38653 = a_2 & ~w3539;
assign w38654 = a_2 & w28381;
assign w38655 = a_2 & w3539;
assign w38656 = a_8 & ~w28384;
assign w38657 = a_8 & ~w3563;
assign w38658 = a_8 & w28384;
assign w38659 = a_8 & w3563;
assign w38660 = a_20 & ~w28386;
assign w38661 = a_20 & ~w3576;
assign w38662 = a_20 & w28386;
assign w38663 = a_20 & w3576;
assign w38664 = a_29 & ~w28388;
assign w38665 = a_29 & ~w3587;
assign w38666 = a_29 & w28388;
assign w38667 = a_29 & w3587;
assign w38668 = a_26 & ~w28390;
assign w38669 = a_26 & ~w3625;
assign w38670 = a_26 & w28390;
assign w38671 = a_26 & w3625;
assign w38672 = a_23 & ~w28392;
assign w38673 = a_23 & ~w28393;
assign w38674 = a_17 & ~w28395;
assign w38675 = a_17 & ~w3664;
assign w38676 = a_17 & w28395;
assign w38677 = a_17 & w3664;
assign w38678 = a_14 & ~w28397;
assign w38679 = a_14 & ~w3680;
assign w38680 = a_14 & w28397;
assign w38681 = a_14 & w3680;
assign w38682 = a_5 & ~w28404;
assign w38683 = a_5 & ~w3721;
assign w38684 = a_5 & w28404;
assign w38685 = a_5 & w3721;
assign w38686 = (w28408 & w28407) | (w28408 & w28238) | (w28407 & w28238);
assign w38687 = (w28408 & w28407) | (w28408 & w28237) | (w28407 & w28237);
assign w38688 = w3741 & ~w38687;
assign w38689 = w3741 & ~w38686;
assign w38690 = ~w3741 & w38687;
assign w38691 = ~w3741 & w38686;
assign w38692 = a_2 & ~w28409;
assign w38693 = a_2 & ~w3738;
assign w38694 = a_2 & w28409;
assign w38695 = a_2 & w3738;
assign w38696 = w3730 & ~w3727;
assign w38697 = a_26 & ~w28412;
assign w38698 = a_26 & ~w3764;
assign w38699 = a_26 & w28412;
assign w38700 = a_26 & w3764;
assign w38701 = a_29 & ~w28414;
assign w38702 = a_29 & ~w3775;
assign w38703 = a_29 & w28414;
assign w38704 = a_29 & w3775;
assign w38705 = a_23 & ~w28419;
assign w38706 = a_23 & ~w3839;
assign w38707 = a_23 & w28419;
assign w38708 = a_23 & w3839;
assign w38709 = a_20 & ~w28421;
assign w38710 = a_20 & ~w3856;
assign w38711 = a_20 & w28421;
assign w38712 = a_20 & w3856;
assign w38713 = ~w3864 & w3866;
assign w38714 = w3864 & ~w3866;
assign w38715 = ~w3935 & w3936;
assign w38716 = w3935 & ~w3936;
assign w38717 = a_5 & ~w28446;
assign w38718 = a_5 & ~w3944;
assign w38719 = a_5 & w28446;
assign w38720 = a_5 & w3944;
assign w38721 = ~w3951 & w25032;
assign w38722 = (w25032 & ~w3951) | (w25032 & ~w3730) | (~w3951 & ~w3730);
assign w38723 = (w28450 & w28451) | (w28450 & ~w38687) | (w28451 & ~w38687);
assign w38724 = (w28450 & w28451) | (w28450 & ~w38686) | (w28451 & ~w38686);
assign w38725 = (w28452 & w28453) | (w28452 & w38687) | (w28453 & w38687);
assign w38726 = (w28452 & w28453) | (w28452 & w38686) | (w28453 & w38686);
assign w38727 = a_2 & ~w28454;
assign w38728 = a_2 & ~w3961;
assign w38729 = a_2 & w28454;
assign w38730 = a_2 & w3961;
assign w38731 = w3975 & ~w3979;
assign w38732 = a_11 & ~w28464;
assign w38733 = a_11 & ~w3995;
assign w38734 = a_11 & w28464;
assign w38735 = a_11 & w3995;
assign w38736 = a_20 & ~w28466;
assign w38737 = a_20 & ~w4007;
assign w38738 = a_20 & w28466;
assign w38739 = a_20 & w4007;
assign w38740 = a_26 & ~w28468;
assign w38741 = a_26 & ~w4018;
assign w38742 = a_26 & w28468;
assign w38743 = a_26 & w4018;
assign w38744 = ~w26895 & a_32;
assign w38745 = w308 & w4063;
assign w38746 = w28472 & a_29;
assign w38747 = (a_29 & w28472) | (a_29 & ~w308) | (w28472 & ~w308);
assign w38748 = a_23 & ~w28477;
assign w38749 = a_23 & ~w4087;
assign w38750 = a_23 & w28477;
assign w38751 = a_23 & w4087;
assign w38752 = a_17 & ~w28479;
assign w38753 = a_17 & ~w4111;
assign w38754 = a_17 & w28479;
assign w38755 = a_17 & w4111;
assign w38756 = ~w4118 & w4002;
assign w38757 = a_14 & ~w28481;
assign w38758 = a_14 & ~w4128;
assign w38759 = a_14 & w28481;
assign w38760 = a_14 & w4128;
assign w38761 = a_5 & ~w28483;
assign w38762 = a_5 & ~w4158;
assign w38763 = a_5 & w28483;
assign w38764 = a_5 & w4158;
assign w38765 = ~w4164 & w3952;
assign w38766 = ~w4164 & w4165;
assign w38767 = ~w4164 & ~w3952;
assign w38768 = (w28490 & w28491) | (w28490 & ~w38687) | (w28491 & ~w38687);
assign w38769 = (w28490 & w28491) | (w28490 & ~w38686) | (w28491 & ~w38686);
assign w38770 = (w28492 & w28493) | (w28492 & w38687) | (w28493 & w38687);
assign w38771 = (w28492 & w28493) | (w28492 & w38686) | (w28493 & w38686);
assign w38772 = a_2 & ~w28494;
assign w38773 = a_2 & ~w4175;
assign w38774 = a_2 & w28494;
assign w38775 = a_2 & w4175;
assign w38776 = a_5 & ~w28498;
assign w38777 = a_5 & ~w4197;
assign w38778 = a_5 & w28498;
assign w38779 = a_5 & w4197;
assign w38780 = a_11 & ~w28500;
assign w38781 = a_11 & ~w4209;
assign w38782 = a_11 & w28500;
assign w38783 = a_11 & w4209;
assign w38784 = a_23 & ~w28504;
assign w38785 = a_23 & ~w4222;
assign w38786 = a_23 & w28504;
assign w38787 = a_23 & w4222;
assign w38788 = a_32 & ~w28506;
assign w38789 = a_32 & ~w4233;
assign w38790 = a_32 & w28506;
assign w38791 = a_32 & w4233;
assign w38792 = a_29 & ~w28508;
assign w38793 = a_29 & ~w4271;
assign w38794 = a_29 & w28508;
assign w38795 = a_29 & w4271;
assign w38796 = a_26 & ~w28510;
assign w38797 = a_26 & ~w4287;
assign w38798 = a_26 & w28510;
assign w38799 = a_26 & w4287;
assign w38800 = a_20 & ~w28512;
assign w38801 = a_20 & ~w4311;
assign w38802 = a_20 & w28512;
assign w38803 = a_20 & w4311;
assign w38804 = a_17 & ~w28514;
assign w38805 = a_17 & ~w4327;
assign w38806 = a_17 & w28514;
assign w38807 = a_17 & w4327;
assign w38808 = a_14 & ~w28516;
assign w38809 = a_14 & ~w4344;
assign w38810 = a_14 & w28516;
assign w38811 = a_14 & w4344;
assign w38812 = a_8 & ~w28518;
assign w38813 = a_8 & ~w4367;
assign w38814 = a_8 & w28518;
assign w38815 = a_8 & w4367;
assign w38816 = (w28523 & w28522) | (w28523 & ~w38687) | (w28522 & ~w38687);
assign w38817 = (w28523 & w28522) | (w28523 & ~w38686) | (w28522 & ~w38686);
assign w38818 = (w28525 & w28524) | (w28525 & w38687) | (w28524 & w38687);
assign w38819 = (w28525 & w28524) | (w28525 & w38686) | (w28524 & w38686);
assign w38820 = a_2 & ~w4389;
assign w38821 = a_2 & ~w28526;
assign w38822 = a_2 & w4389;
assign w38823 = a_2 & w28526;
assign w38824 = a_5 & ~w28530;
assign w38825 = a_5 & ~w4415;
assign w38826 = a_5 & w28530;
assign w38827 = a_5 & w4415;
assign w38828 = a_8 & ~w28532;
assign w38829 = a_8 & ~w4426;
assign w38830 = a_8 & w28532;
assign w38831 = a_8 & w4426;
assign w38832 = a_23 & ~w28534;
assign w38833 = a_23 & ~w4438;
assign w38834 = a_23 & w28534;
assign w38835 = a_23 & w4438;
assign w38836 = a_26 & ~w28536;
assign w38837 = a_26 & ~w4449;
assign w38838 = a_26 & w28536;
assign w38839 = a_26 & w4449;
assign w38840 = a_29 & ~w28538;
assign w38841 = a_29 & ~w4460;
assign w38842 = a_29 & w28538;
assign w38843 = a_29 & w4460;
assign w38844 = a_32 & ~w28540;
assign w38845 = a_32 & ~w4471;
assign w38846 = a_32 & w28540;
assign w38847 = a_32 & w4471;
assign w38848 = a_20 & ~w28545;
assign w38849 = a_20 & ~w4547;
assign w38850 = a_20 & w28545;
assign w38851 = a_20 & w4547;
assign w38852 = a_17 & ~w28547;
assign w38853 = a_17 & ~w4565;
assign w38854 = a_17 & w28547;
assign w38855 = a_17 & w4565;
assign w38856 = a_14 & ~w28549;
assign w38857 = a_14 & ~w4583;
assign w38858 = a_14 & w28549;
assign w38859 = a_14 & w4583;
assign w38860 = a_11 & ~w28552;
assign w38861 = a_11 & ~w4600;
assign w38862 = a_11 & w28552;
assign w38863 = a_11 & w4600;
assign w38864 = (w28557 & w28558) | (w28557 & ~w38687) | (w28558 & ~w38687);
assign w38865 = (w28557 & w28558) | (w28557 & ~w38686) | (w28558 & ~w38686);
assign w38866 = (w28559 & w28560) | (w28559 & w38687) | (w28560 & w38687);
assign w38867 = (w28559 & w28560) | (w28559 & w38686) | (w28560 & w38686);
assign w38868 = a_2 & ~w28561;
assign w38869 = a_2 & ~w4630;
assign w38870 = a_2 & w28561;
assign w38871 = a_2 & w4630;
assign w38872 = (w28566 & w28565) | (w28566 & ~w38687) | (w28565 & ~w38687);
assign w38873 = (w28566 & w28565) | (w28566 & ~w38686) | (w28565 & ~w38686);
assign w38874 = (w28567 & w28568) | (w28567 & w38687) | (w28568 & w38687);
assign w38875 = (w28567 & w28568) | (w28567 & w38686) | (w28568 & w38686);
assign w38876 = a_2 & ~w28569;
assign w38877 = a_2 & ~w4652;
assign w38878 = a_2 & w28569;
assign w38879 = a_2 & w4652;
assign w38880 = a_5 & ~w28572;
assign w38881 = a_5 & ~w4669;
assign w38882 = a_5 & w28572;
assign w38883 = a_5 & w4669;
assign w38884 = a_8 & ~w28574;
assign w38885 = a_8 & ~w4680;
assign w38886 = a_8 & w28574;
assign w38887 = a_8 & w4680;
assign w38888 = a_11 & ~w28577;
assign w38889 = a_11 & ~w4691;
assign w38890 = a_11 & w28577;
assign w38891 = a_11 & w4691;
assign w38892 = a_23 & ~w28579;
assign w38893 = a_23 & ~w4702;
assign w38894 = a_23 & w28579;
assign w38895 = a_23 & w4702;
assign w38896 = a_29 & ~w28581;
assign w38897 = a_29 & ~w4714;
assign w38898 = a_29 & w28581;
assign w38899 = a_29 & w4714;
assign w38900 = ~w26548 & a_35;
assign w38901 = w308 & w4759;
assign w38902 = w28585 & a_32;
assign w38903 = (a_32 & w28585) | (a_32 & ~w308) | (w28585 & ~w308);
assign w38904 = a_26 & ~w28588;
assign w38905 = a_26 & ~w4782;
assign w38906 = a_26 & w28588;
assign w38907 = a_26 & w4782;
assign w38908 = w4539 & ~w4535;
assign w38909 = a_20 & ~w28590;
assign w38910 = a_20 & ~w4806;
assign w38911 = a_20 & w28590;
assign w38912 = a_20 & w4806;
assign w38913 = w4557 & ~w4553;
assign w38914 = a_17 & ~w28592;
assign w38915 = a_17 & ~w4824;
assign w38916 = a_17 & w28592;
assign w38917 = a_17 & w4824;
assign w38918 = ~w4830 & ~w27340;
assign w38919 = ~w4830 & ~w27339;
assign w38920 = ~w27339 & w27340;
assign w38921 = a_14 & ~w28594;
assign w38922 = a_14 & ~w4840;
assign w38923 = a_14 & w28594;
assign w38924 = a_14 & w4840;
assign w38925 = ~w4835 & w4845;
assign w38926 = w4835 & ~w4845;
assign w38927 = a_2 & ~w28600;
assign w38928 = a_2 & ~w4882;
assign w38929 = a_2 & w28600;
assign w38930 = a_2 & w4882;
assign w38931 = ~w4866 & ~w4865;
assign w38932 = ~w4847 & ~w4848;
assign w38933 = a_14 & ~w28608;
assign w38934 = a_14 & ~w4912;
assign w38935 = a_14 & w28608;
assign w38936 = a_14 & w4912;
assign w38937 = a_26 & ~w28611;
assign w38938 = a_26 & ~w4924;
assign w38939 = a_26 & w28611;
assign w38940 = a_26 & w4924;
assign w38941 = a_35 & ~w28613;
assign w38942 = a_35 & ~w4934;
assign w38943 = a_35 & w28613;
assign w38944 = a_35 & w4934;
assign w38945 = a_32 & ~w28615;
assign w38946 = a_32 & ~w4974;
assign w38947 = a_32 & w28615;
assign w38948 = a_32 & w4974;
assign w38949 = a_29 & ~w28617;
assign w38950 = a_29 & ~w4992;
assign w38951 = a_29 & w28617;
assign w38952 = a_29 & w4992;
assign w38953 = a_23 & ~w28619;
assign w38954 = a_23 & ~w5016;
assign w38955 = a_23 & w28619;
assign w38956 = a_23 & w5016;
assign w38957 = a_20 & ~w28621;
assign w38958 = a_20 & ~w5032;
assign w38959 = a_20 & w28621;
assign w38960 = a_20 & w5032;
assign w38961 = a_17 & ~w28623;
assign w38962 = a_17 & ~w5050;
assign w38963 = a_17 & w28623;
assign w38964 = a_17 & w5050;
assign w38965 = a_11 & ~w28625;
assign w38966 = a_11 & ~w5073;
assign w38967 = a_11 & w28625;
assign w38968 = a_11 & w5073;
assign w38969 = a_5 & ~w28627;
assign w38970 = a_5 & ~w5096;
assign w38971 = a_5 & w28627;
assign w38972 = a_5 & w5096;
assign w38973 = ~w5106 & ~w4893;
assign w38974 = w5106 & ~w4893;
assign w38975 = w5111 & ~w5108;
assign w38976 = a_5 & ~w28631;
assign w38977 = a_5 & ~w5122;
assign w38978 = a_5 & w28631;
assign w38979 = a_5 & w5122;
assign w38980 = a_8 & ~w28634;
assign w38981 = a_8 & ~w5133;
assign w38982 = a_8 & w28634;
assign w38983 = a_8 & w5133;
assign w38984 = a_14 & ~w28636;
assign w38985 = a_14 & ~w5146;
assign w38986 = a_14 & w28636;
assign w38987 = a_14 & w5146;
assign w38988 = a_26 & ~w28638;
assign w38989 = a_26 & ~w5156;
assign w38990 = a_26 & w28638;
assign w38991 = a_26 & w5156;
assign w38992 = a_35 & ~w28640;
assign w38993 = a_35 & ~w5168;
assign w38994 = a_35 & w28640;
assign w38995 = a_35 & w5168;
assign w38996 = a_32 & ~w28645;
assign w38997 = a_32 & ~w5226;
assign w38998 = a_32 & w28645;
assign w38999 = a_32 & w5226;
assign w39000 = a_29 & ~w28647;
assign w39001 = a_29 & ~w5243;
assign w39002 = a_29 & w28647;
assign w39003 = a_29 & w5243;
assign w39004 = a_23 & ~w28650;
assign w39005 = a_23 & ~w5267;
assign w39006 = a_23 & w28650;
assign w39007 = a_23 & w5267;
assign w39008 = a_20 & ~w28652;
assign w39009 = a_20 & ~w5285;
assign w39010 = a_20 & w28652;
assign w39011 = a_20 & w5285;
assign w39012 = a_17 & ~w28654;
assign w39013 = a_17 & ~w5303;
assign w39014 = a_17 & w28654;
assign w39015 = a_17 & w5303;
assign w39016 = a_11 & ~w28656;
assign w39017 = a_11 & ~w5328;
assign w39018 = a_11 & w28656;
assign w39019 = a_11 & w5328;
assign w39020 = ~w5322 & w5333;
assign w39021 = w5322 & ~w5333;
assign w39022 = a_2 & ~w28665;
assign w39023 = a_2 & ~w5357;
assign w39024 = a_2 & w28665;
assign w39025 = a_2 & w5357;
assign w39026 = w5141 & ~w5317;
assign w39027 = a_14 & ~w28680;
assign w39028 = a_14 & ~w5405;
assign w39029 = a_14 & w28680;
assign w39030 = a_14 & w5405;
assign w39031 = w5313 & ~w5309;
assign w39032 = w5295 & ~w5291;
assign w39033 = a_23 & ~w28682;
assign w39034 = a_23 & ~w5417;
assign w39035 = a_23 & w28682;
assign w39036 = a_23 & w5417;
assign w39037 = a_26 & ~w28685;
assign w39038 = a_26 & ~w5428;
assign w39039 = a_26 & w28685;
assign w39040 = a_26 & w5428;
assign w39041 = a_29 & ~w28687;
assign w39042 = a_29 & ~w5439;
assign w39043 = a_29 & w28687;
assign w39044 = a_29 & w5439;
assign w39045 = w308 & w5450;
assign w39046 = w28691 & a_35;
assign w39047 = (a_35 & w28691) | (a_35 & ~w308) | (w28691 & ~w308);
assign w39048 = ~w26552 & a_38;
assign w39049 = a_32 & ~w28694;
assign w39050 = a_32 & ~w5501;
assign w39051 = a_32 & w28694;
assign w39052 = a_32 & w5501;
assign w39053 = a_20 & ~w28696;
assign w39054 = a_20 & ~w5537;
assign w39055 = a_20 & w28696;
assign w39056 = a_20 & w5537;
assign w39057 = a_17 & ~w28701;
assign w39058 = a_17 & ~w5553;
assign w39059 = a_17 & w28701;
assign w39060 = a_17 & w5553;
assign w39061 = a_5 & ~w28709;
assign w39062 = a_5 & ~w5588;
assign w39063 = a_5 & w28709;
assign w39064 = a_5 & w5588;
assign w39065 = a_2 & ~w28718;
assign w39066 = a_2 & ~w5603;
assign w39067 = a_2 & w28718;
assign w39068 = a_2 & w5603;
assign w39069 = a_5 & ~w28724;
assign w39070 = a_5 & ~w5626;
assign w39071 = a_5 & w28724;
assign w39072 = a_5 & w5626;
assign w39073 = a_17 & ~w28732;
assign w39074 = a_17 & ~w5650;
assign w39075 = a_17 & w28732;
assign w39076 = a_17 & w5650;
assign w39077 = a_23 & ~w28734;
assign w39078 = a_23 & ~w5660;
assign w39079 = a_23 & w28734;
assign w39080 = a_23 & w5660;
assign w39081 = a_32 & ~w28737;
assign w39082 = a_32 & ~w5673;
assign w39083 = a_32 & w28737;
assign w39084 = a_32 & w5673;
assign w39085 = a_38 & ~w28739;
assign w39086 = a_38 & ~w5684;
assign w39087 = a_38 & w28739;
assign w39088 = a_38 & w5684;
assign w39089 = a_35 & ~w28741;
assign w39090 = a_35 & ~w5723;
assign w39091 = a_35 & w28741;
assign w39092 = a_35 & w5723;
assign w39093 = a_29 & ~w28743;
assign w39094 = a_29 & ~w5747;
assign w39095 = a_29 & w28743;
assign w39096 = a_29 & w5747;
assign w39097 = a_26 & ~w28745;
assign w39098 = a_26 & ~w5764;
assign w39099 = a_26 & w28745;
assign w39100 = a_26 & w5764;
assign w39101 = a_20 & ~w28747;
assign w39102 = a_20 & ~w5788;
assign w39103 = a_20 & w28747;
assign w39104 = a_20 & w5788;
assign w39105 = a_14 & ~w28749;
assign w39106 = a_14 & ~w5811;
assign w39107 = a_14 & w28749;
assign w39108 = a_14 & w5811;
assign w39109 = a_2 & ~w28762;
assign w39110 = a_2 & ~w5858;
assign w39111 = a_2 & w28762;
assign w39112 = a_2 & w5858;
assign w39113 = w5851 & ~w5869;
assign w39114 = ~w5851 & ~w5869;
assign w39115 = ~w5616 & ~w5617;
assign w39116 = ~w5616 & ~w5372;
assign w39117 = a_2 & ~w28770;
assign w39118 = a_2 & ~w5882;
assign w39119 = a_2 & w28770;
assign w39120 = a_2 & w5882;
assign w39121 = w5621 & ~w5846;
assign w39122 = a_11 & ~w28772;
assign w39123 = a_11 & ~w5900;
assign w39124 = a_11 & w28772;
assign w39125 = a_11 & w5900;
assign w39126 = a_17 & ~w28775;
assign w39127 = a_17 & ~w5912;
assign w39128 = a_17 & w28775;
assign w39129 = a_17 & w5912;
assign w39130 = a_29 & ~w28777;
assign w39131 = a_29 & ~w5922;
assign w39132 = a_29 & w28777;
assign w39133 = a_29 & w5922;
assign w39134 = a_38 & ~w28779;
assign w39135 = a_38 & ~w5934;
assign w39136 = a_38 & w28779;
assign w39137 = a_38 & w5934;
assign w39138 = a_35 & ~w28784;
assign w39139 = a_35 & ~w5992;
assign w39140 = a_35 & w28784;
assign w39141 = a_35 & w5992;
assign w39142 = a_32 & ~w28786;
assign w39143 = a_32 & ~w6009;
assign w39144 = a_32 & w28786;
assign w39145 = a_32 & w6009;
assign w39146 = a_26 & ~w28788;
assign w39147 = a_26 & ~w6033;
assign w39148 = a_26 & w28788;
assign w39149 = a_26 & w6033;
assign w39150 = a_23 & ~w28790;
assign w39151 = a_23 & ~w6051;
assign w39152 = a_23 & w28790;
assign w39153 = a_23 & w6051;
assign w39154 = a_20 & ~w28792;
assign w39155 = a_20 & ~w6069;
assign w39156 = a_20 & w28792;
assign w39157 = a_20 & w6069;
assign w39158 = w6084 & ~w5907;
assign w39159 = a_14 & ~w28794;
assign w39160 = a_14 & ~w6093;
assign w39161 = a_14 & w28794;
assign w39162 = a_14 & w6093;
assign w39163 = a_8 & ~w28796;
assign w39164 = a_8 & ~w6118;
assign w39165 = a_8 & w28796;
assign w39166 = a_8 & w6118;
assign w39167 = a_5 & ~w28799;
assign w39168 = a_5 & ~w6135;
assign w39169 = a_5 & w28799;
assign w39170 = a_5 & w6135;
assign w39171 = a_5 & ~w28802;
assign w39172 = a_5 & ~w6161;
assign w39173 = a_5 & w28802;
assign w39174 = a_5 & w6161;
assign w39175 = a_11 & ~w28804;
assign w39176 = a_11 & ~w6171;
assign w39177 = a_11 & w28804;
assign w39178 = a_11 & w6171;
assign w39179 = a_14 & ~w28806;
assign w39180 = a_14 & ~w6182;
assign w39181 = a_14 & w28806;
assign w39182 = a_14 & w6182;
assign w39183 = a_17 & ~w28808;
assign w39184 = a_17 & ~w6193;
assign w39185 = a_17 & w28808;
assign w39186 = a_17 & w6193;
assign w39187 = a_26 & ~w28810;
assign w39188 = a_26 & ~w6205;
assign w39189 = a_26 & w28810;
assign w39190 = a_26 & w6205;
assign w39191 = a_29 & ~w28812;
assign w39192 = a_29 & ~w6215;
assign w39193 = a_29 & w28812;
assign w39194 = a_29 & w6215;
assign w39195 = a_32 & ~w28814;
assign w39196 = a_32 & ~w6226;
assign w39197 = a_32 & w28814;
assign w39198 = a_32 & w6226;
assign w39199 = w308 & w6237;
assign w39200 = w28818 & a_38;
assign w39201 = (a_38 & w28818) | (a_38 & ~w308) | (w28818 & ~w308);
assign w39202 = ~w26557 & a_41;
assign w39203 = a_35 & ~w28821;
assign w39204 = a_35 & ~w6288;
assign w39205 = a_35 & w28821;
assign w39206 = a_35 & w6288;
assign w39207 = a_23 & ~w28823;
assign w39208 = a_23 & ~w6324;
assign w39209 = a_23 & w28823;
assign w39210 = a_23 & w6324;
assign w39211 = ~w6331 & w6200;
assign w39212 = a_20 & ~w28825;
assign w39213 = a_20 & ~w6341;
assign w39214 = a_20 & w28825;
assign w39215 = a_20 & w6341;
assign w39216 = a_2 & ~w28838;
assign w39217 = a_2 & ~w6402;
assign w39218 = a_2 & w28838;
assign w39219 = a_2 & w6402;
assign w39220 = a_14 & ~w28841;
assign w39221 = a_14 & ~w6428;
assign w39222 = a_14 & w28841;
assign w39223 = a_14 & w6428;
assign w39224 = a_20 & ~w28844;
assign w39225 = a_20 & ~w6440;
assign w39226 = a_20 & w28844;
assign w39227 = a_20 & w6440;
assign w39228 = a_26 & ~w28846;
assign w39229 = a_26 & ~w6450;
assign w39230 = a_26 & w28846;
assign w39231 = a_26 & w6450;
assign w39232 = a_35 & ~w28851;
assign w39233 = a_35 & ~w6463;
assign w39234 = a_35 & w28851;
assign w39235 = a_35 & w6463;
assign w39236 = a_41 & ~w28853;
assign w39237 = a_41 & ~w6474;
assign w39238 = a_41 & w28853;
assign w39239 = a_41 & w6474;
assign w39240 = a_38 & ~w28855;
assign w39241 = a_38 & ~w6513;
assign w39242 = a_38 & w28855;
assign w39243 = a_38 & w6513;
assign w39244 = a_32 & ~w28857;
assign w39245 = a_32 & ~w6537;
assign w39246 = a_32 & w28857;
assign w39247 = a_32 & w6537;
assign w39248 = a_29 & ~w28859;
assign w39249 = a_29 & ~w6554;
assign w39250 = a_29 & w28859;
assign w39251 = a_29 & w6554;
assign w39252 = w6316 & ~w6312;
assign w39253 = a_23 & ~w28861;
assign w39254 = a_23 & ~w6578;
assign w39255 = a_23 & w28861;
assign w39256 = a_23 & w6578;
assign w39257 = a_17 & ~w28863;
assign w39258 = a_17 & ~w6601;
assign w39259 = a_17 & w28863;
assign w39260 = a_17 & w6601;
assign w39261 = a_11 & ~w28865;
assign w39262 = a_11 & ~w6624;
assign w39263 = a_11 & w28865;
assign w39264 = a_11 & w6624;
assign w39265 = a_5 & ~w28872;
assign w39266 = a_5 & ~w6658;
assign w39267 = a_5 & w28872;
assign w39268 = a_5 & w6658;
assign w39269 = (w6679 & w28875) | (w6679 & w28835) | (w28875 & w28835);
assign w39270 = (w6679 & w28875) | (w6679 & w28834) | (w28875 & w28834);
assign w39271 = w28876 & ~w28835;
assign w39272 = w28876 & ~w28834;
assign w39273 = a_2 & ~w28877;
assign w39274 = a_2 & ~w6676;
assign w39275 = a_2 & w28877;
assign w39276 = a_2 & w6676;
assign w39277 = w6649 & ~w6646;
assign w39278 = a_14 & ~w28879;
assign w39279 = a_14 & ~w6699;
assign w39280 = a_14 & w28879;
assign w39281 = a_14 & w6699;
assign w39282 = a_20 & ~w28882;
assign w39283 = a_20 & ~w6711;
assign w39284 = a_20 & w28882;
assign w39285 = a_20 & w6711;
assign w39286 = a_32 & ~w28884;
assign w39287 = a_32 & ~w6721;
assign w39288 = a_32 & w28884;
assign w39289 = a_32 & w6721;
assign w39290 = a_41 & ~w28886;
assign w39291 = a_41 & ~w6733;
assign w39292 = a_41 & w28886;
assign w39293 = a_41 & w6733;
assign w39294 = a_38 & ~w28891;
assign w39295 = a_38 & ~w6791;
assign w39296 = a_38 & w28891;
assign w39297 = a_38 & w6791;
assign w39298 = a_35 & ~w28893;
assign w39299 = a_35 & ~w6808;
assign w39300 = a_35 & w28893;
assign w39301 = a_35 & w6808;
assign w39302 = a_29 & ~w28895;
assign w39303 = a_29 & ~w6832;
assign w39304 = a_29 & w28895;
assign w39305 = a_29 & w6832;
assign w39306 = a_26 & ~w28897;
assign w39307 = a_26 & ~w6850;
assign w39308 = a_26 & w28897;
assign w39309 = a_26 & w6850;
assign w39310 = a_23 & ~w28900;
assign w39311 = a_23 & ~w6868;
assign w39312 = a_23 & w28900;
assign w39313 = a_23 & w6868;
assign w39314 = ~w6586 & ~w6585;
assign w39315 = a_17 & ~w28902;
assign w39316 = a_17 & ~w6892;
assign w39317 = a_17 & w28902;
assign w39318 = a_17 & w6892;
assign w39319 = a_11 & ~w28905;
assign w39320 = a_11 & ~w6916;
assign w39321 = a_11 & w28905;
assign w39322 = a_11 & w6916;
assign w39323 = a_8 & ~w28907;
assign w39324 = a_8 & ~w6934;
assign w39325 = a_8 & w28907;
assign w39326 = a_8 & w6934;
assign w39327 = ~w6694 & ~w25052;
assign w39328 = ~w6694 & ~w6652;
assign w39329 = ~w6940 & ~w25052;
assign w39330 = ~w6940 & ~w6652;
assign w39331 = ~w6652 & w25052;
assign w39332 = a_5 & ~w28910;
assign w39333 = a_5 & ~w6950;
assign w39334 = a_5 & w28910;
assign w39335 = a_5 & w6950;
assign w39336 = w6668 & ~w6664;
assign w39337 = (w28916 & w28915) | (w28916 & w28835) | (w28915 & w28835);
assign w39338 = (w28916 & w28915) | (w28916 & w28834) | (w28915 & w28834);
assign w39339 = (w28918 & w28917) | (w28918 & ~w28835) | (w28917 & ~w28835);
assign w39340 = (w28918 & w28917) | (w28918 & ~w28834) | (w28917 & ~w28834);
assign w39341 = a_2 & ~w28919;
assign w39342 = a_2 & ~w6968;
assign w39343 = a_2 & w28919;
assign w39344 = a_2 & w6968;
assign w39345 = (w28927 & w28926) | (w28927 & w28835) | (w28926 & w28835);
assign w39346 = (w28927 & w28926) | (w28927 & w28834) | (w28926 & w28834);
assign w39347 = (w28929 & w28928) | (w28929 & ~w28835) | (w28928 & ~w28835);
assign w39348 = (w28929 & w28928) | (w28929 & ~w28834) | (w28928 & ~w28834);
assign w39349 = a_2 & ~w28930;
assign w39350 = a_2 & ~w6992;
assign w39351 = a_2 & w28930;
assign w39352 = a_2 & w6992;
assign w39353 = w6960 & ~w6956;
assign w39354 = a_14 & ~w28932;
assign w39355 = a_14 & ~w7009;
assign w39356 = a_14 & w28932;
assign w39357 = a_14 & w7009;
assign w39358 = a_17 & ~w28934;
assign w39359 = a_17 & ~w7020;
assign w39360 = a_17 & w28934;
assign w39361 = a_17 & w7020;
assign w39362 = a_20 & ~w28936;
assign w39363 = a_20 & ~w7031;
assign w39364 = a_20 & w28936;
assign w39365 = a_20 & w7031;
assign w39366 = a_32 & ~w28938;
assign w39367 = a_32 & ~w7044;
assign w39368 = a_32 & w28938;
assign w39369 = a_32 & w7044;
assign w39370 = a_35 & ~w28940;
assign w39371 = a_35 & ~w7055;
assign w39372 = a_35 & w28940;
assign w39373 = a_35 & w7055;
assign w39374 = w308 & w7066;
assign w39375 = w28944 & a_41;
assign w39376 = (a_41 & w28944) | (a_41 & ~w308) | (w28944 & ~w308);
assign w39377 = ~w26789 & a_44;
assign w39378 = a_38 & ~w28947;
assign w39379 = a_38 & ~w7117;
assign w39380 = a_38 & w28947;
assign w39381 = a_38 & w7117;
assign w39382 = a_29 & ~w28949;
assign w39383 = a_29 & ~w7147;
assign w39384 = a_29 & w28949;
assign w39385 = a_29 & w7147;
assign w39386 = a_26 & ~w28952;
assign w39387 = a_26 & ~w7165;
assign w39388 = a_26 & w28952;
assign w39389 = a_26 & w7165;
assign w39390 = a_23 & ~w28955;
assign w39391 = a_23 & ~w7182;
assign w39392 = a_23 & w28955;
assign w39393 = a_23 & w7182;
assign w39394 = a_8 & ~w28962;
assign w39395 = a_8 & ~w7236;
assign w39396 = a_8 & w28962;
assign w39397 = a_8 & w7236;
assign w39398 = ~w7243 & w6943;
assign w39399 = a_5 & ~w28965;
assign w39400 = a_5 & ~w7253;
assign w39401 = a_5 & w28965;
assign w39402 = a_5 & w7253;
assign w39403 = ~w7263 & ~w7003;
assign w39404 = w7263 & ~w7003;
assign w39405 = (w28973 & w28972) | (w28973 & w28835) | (w28972 & w28835);
assign w39406 = (w28973 & w28972) | (w28973 & w28834) | (w28972 & w28834);
assign w39407 = (w28975 & w28974) | (w28975 & ~w28835) | (w28974 & ~w28835);
assign w39408 = (w28975 & w28974) | (w28975 & ~w28834) | (w28974 & ~w28834);
assign w39409 = a_2 & ~w28976;
assign w39410 = a_2 & ~w7278;
assign w39411 = a_2 & w28976;
assign w39412 = a_2 & w7278;
assign w39413 = a_17 & ~w28980;
assign w39414 = a_17 & ~w7296;
assign w39415 = a_17 & w28980;
assign w39416 = a_17 & w7296;
assign w39417 = a_23 & ~w28982;
assign w39418 = a_23 & ~w7307;
assign w39419 = a_23 & w28982;
assign w39420 = a_23 & w7307;
assign w39421 = a_35 & ~w28984;
assign w39422 = a_35 & ~w7318;
assign w39423 = a_35 & w28984;
assign w39424 = a_35 & w7318;
assign w39425 = a_38 & ~w28987;
assign w39426 = a_38 & ~w7329;
assign w39427 = a_38 & w28987;
assign w39428 = a_38 & w7329;
assign w39429 = a_44 & ~w28989;
assign w39430 = a_44 & ~w7340;
assign w39431 = a_44 & w28989;
assign w39432 = a_44 & w7340;
assign w39433 = a_41 & ~w28991;
assign w39434 = a_41 & ~w7379;
assign w39435 = a_41 & w28991;
assign w39436 = a_41 & w7379;
assign w39437 = a_32 & ~w28995;
assign w39438 = a_32 & ~w7408;
assign w39439 = a_32 & w28995;
assign w39440 = a_32 & w7408;
assign w39441 = a_29 & ~w28997;
assign w39442 = a_29 & ~w7426;
assign w39443 = a_29 & w28997;
assign w39444 = a_29 & w7426;
assign w39445 = a_26 & ~w28999;
assign w39446 = a_26 & ~w7444;
assign w39447 = a_26 & w28999;
assign w39448 = a_26 & w7444;
assign w39449 = a_20 & ~w29001;
assign w39450 = a_20 & ~w7467;
assign w39451 = a_20 & w29001;
assign w39452 = a_20 & w7467;
assign w39453 = a_5 & ~w29016;
assign w39454 = a_5 & ~w7541;
assign w39455 = a_5 & w29016;
assign w39456 = a_5 & w7541;
assign w39457 = ~w7552 & ~w7553;
assign w39458 = ~w7552 & ~w7270;
assign w39459 = a_23 & ~w29020;
assign w39460 = a_23 & ~w7563;
assign w39461 = a_23 & w29020;
assign w39462 = a_23 & w7563;
assign w39463 = a_35 & ~w29022;
assign w39464 = a_35 & ~w7573;
assign w39465 = a_35 & w29022;
assign w39466 = a_35 & w7573;
assign w39467 = a_44 & ~w29024;
assign w39468 = a_44 & ~w7585;
assign w39469 = a_44 & w29024;
assign w39470 = a_44 & w7585;
assign w39471 = a_41 & ~w29029;
assign w39472 = a_41 & ~w7643;
assign w39473 = a_41 & w29029;
assign w39474 = a_41 & w7643;
assign w39475 = a_38 & ~w29031;
assign w39476 = a_38 & ~w7660;
assign w39477 = a_38 & w29031;
assign w39478 = a_38 & w7660;
assign w39479 = a_32 & ~w29033;
assign w39480 = a_32 & ~w7684;
assign w39481 = a_32 & w29033;
assign w39482 = a_32 & w7684;
assign w39483 = a_29 & ~w29035;
assign w39484 = a_29 & ~w7702;
assign w39485 = a_29 & w29035;
assign w39486 = a_29 & w7702;
assign w39487 = a_26 & ~w29037;
assign w39488 = a_26 & ~w7720;
assign w39489 = a_26 & w29037;
assign w39490 = a_26 & w7720;
assign w39491 = a_20 & ~w29039;
assign w39492 = a_20 & ~w7745;
assign w39493 = a_20 & w29039;
assign w39494 = a_20 & w7745;
assign w39495 = a_17 & ~w29042;
assign w39496 = a_17 & ~w7763;
assign w39497 = a_17 & w29042;
assign w39498 = a_17 & w7763;
assign w39499 = a_5 & ~w29060;
assign w39500 = a_5 & ~w7835;
assign w39501 = a_5 & w29060;
assign w39502 = a_5 & w7835;
assign w39503 = w7829 & ~w7840;
assign w39504 = (w29067 & w29066) | (w29067 & w28835) | (w29066 & w28835);
assign w39505 = (w29067 & w29066) | (w29067 & w28834) | (w29066 & w28834);
assign w39506 = (w29069 & w29068) | (w29069 & ~w28835) | (w29068 & ~w28835);
assign w39507 = (w29069 & w29068) | (w29069 & ~w28834) | (w29068 & ~w28834);
assign w39508 = a_2 & ~w29070;
assign w39509 = a_2 & ~w7853;
assign w39510 = a_2 & w29070;
assign w39511 = a_2 & w7853;
assign w39512 = a_17 & ~w29072;
assign w39513 = a_17 & ~w7876;
assign w39514 = a_17 & w29072;
assign w39515 = a_17 & w7876;
assign w39516 = a_20 & ~w29074;
assign w39517 = a_20 & ~w7887;
assign w39518 = a_20 & w29074;
assign w39519 = a_20 & w7887;
assign w39520 = a_23 & ~w29076;
assign w39521 = a_23 & ~w7898;
assign w39522 = a_23 & w29076;
assign w39523 = a_23 & w7898;
assign w39524 = w7712 & ~w7708;
assign w39525 = a_35 & ~w29078;
assign w39526 = a_35 & ~w7911;
assign w39527 = a_35 & w29078;
assign w39528 = a_35 & w7911;
assign w39529 = a_38 & ~w29080;
assign w39530 = a_38 & ~w7922;
assign w39531 = a_38 & w29080;
assign w39532 = a_38 & w7922;
assign w39533 = w308 & w7933;
assign w39534 = w29084 & a_44;
assign w39535 = (a_44 & w29084) | (a_44 & ~w308) | (w29084 & ~w308);
assign w39536 = ~w26159 & a_47;
assign w39537 = a_41 & ~w29087;
assign w39538 = a_41 & ~w7983;
assign w39539 = a_41 & w29087;
assign w39540 = a_41 & w7983;
assign w39541 = a_32 & ~w29089;
assign w39542 = a_32 & ~w8014;
assign w39543 = a_32 & w29089;
assign w39544 = a_32 & w8014;
assign w39545 = ~w8008 & ~w8019;
assign w39546 = a_29 & ~w29091;
assign w39547 = a_29 & ~w8032;
assign w39548 = a_29 & w29091;
assign w39549 = a_29 & w8032;
assign w39550 = a_26 & ~w29093;
assign w39551 = a_26 & ~w8049;
assign w39552 = a_26 & w29093;
assign w39553 = a_26 & w8049;
assign w39554 = (w29116 & w29115) | (w29116 & w28835) | (w29115 & w28835);
assign w39555 = (w29116 & w29115) | (w29116 & w28834) | (w29115 & w28834);
assign w39556 = (w29117 & w29118) | (w29117 & ~w28835) | (w29118 & ~w28835);
assign w39557 = (w29117 & w29118) | (w29117 & ~w28834) | (w29118 & ~w28834);
assign w39558 = a_2 & ~w29119;
assign w39559 = a_2 & ~w8156;
assign w39560 = a_2 & w29119;
assign w39561 = a_2 & w8156;
assign w39562 = (w29124 & w29123) | (w29124 & w28835) | (w29123 & w28835);
assign w39563 = (w29124 & w29123) | (w29124 & w28834) | (w29123 & w28834);
assign w39564 = (w29126 & w29125) | (w29126 & ~w28835) | (w29125 & ~w28835);
assign w39565 = (w29126 & w29125) | (w29126 & ~w28834) | (w29125 & ~w28834);
assign w39566 = a_2 & ~w29127;
assign w39567 = a_2 & ~w8180;
assign w39568 = a_2 & w29127;
assign w39569 = a_2 & w8180;
assign w39570 = a_26 & ~w29136;
assign w39571 = a_26 & ~w8220;
assign w39572 = a_26 & w29136;
assign w39573 = a_26 & w8220;
assign w39574 = a_35 & ~w29138;
assign w39575 = a_35 & ~w8231;
assign w39576 = a_35 & w29138;
assign w39577 = a_35 & w8231;
assign w39578 = a_38 & ~w29140;
assign w39579 = a_38 & ~w8242;
assign w39580 = a_38 & w29140;
assign w39581 = a_38 & w8242;
assign w39582 = a_41 & ~w29142;
assign w39583 = a_41 & ~w8253;
assign w39584 = a_41 & w29142;
assign w39585 = a_41 & w8253;
assign w39586 = a_47 & ~w29144;
assign w39587 = a_47 & ~w8263;
assign w39588 = a_47 & w29144;
assign w39589 = a_47 & w8263;
assign w39590 = a_44 & ~w29146;
assign w39591 = a_44 & ~w8302;
assign w39592 = a_44 & w29146;
assign w39593 = a_44 & w8302;
assign w39594 = a_32 & ~w29148;
assign w39595 = a_32 & ~w8337;
assign w39596 = a_32 & w29148;
assign w39597 = a_32 & w8337;
assign w39598 = a_29 & ~w29150;
assign w39599 = a_29 & ~w8355;
assign w39600 = a_29 & w29150;
assign w39601 = a_29 & w8355;
assign w39602 = a_23 & ~w29152;
assign w39603 = a_23 & ~w8378;
assign w39604 = a_23 & w29152;
assign w39605 = a_23 & w8378;
assign w39606 = a_5 & ~w29165;
assign w39607 = a_5 & ~w8459;
assign w39608 = a_5 & w29165;
assign w39609 = a_5 & w8459;
assign w39610 = a_38 & ~w29170;
assign w39611 = a_38 & ~w8486;
assign w39612 = a_38 & w29170;
assign w39613 = a_38 & w8486;
assign w39614 = a_47 & ~w29172;
assign w39615 = a_47 & ~w8498;
assign w39616 = a_47 & w29172;
assign w39617 = a_47 & w8498;
assign w39618 = a_44 & ~w29175;
assign w39619 = a_44 & ~w8556;
assign w39620 = a_44 & w29175;
assign w39621 = a_44 & w8556;
assign w39622 = a_41 & ~w29177;
assign w39623 = a_41 & ~w8572;
assign w39624 = a_41 & w29177;
assign w39625 = a_41 & w8572;
assign w39626 = a_35 & ~w29179;
assign w39627 = a_35 & ~w8596;
assign w39628 = a_35 & w29179;
assign w39629 = a_35 & w8596;
assign w39630 = a_32 & ~w29181;
assign w39631 = a_32 & ~w8613;
assign w39632 = a_32 & w29181;
assign w39633 = a_32 & w8613;
assign w39634 = a_29 & ~w29183;
assign w39635 = a_29 & ~w8631;
assign w39636 = a_29 & w29183;
assign w39637 = a_29 & w8631;
assign w39638 = a_26 & ~w29185;
assign w39639 = a_26 & ~w8648;
assign w39640 = a_26 & w29185;
assign w39641 = a_26 & w8648;
assign w39642 = ~w8757 & w27540;
assign w39643 = ~w8757 & ~w27745;
assign w39644 = a_5 & ~w29210;
assign w39645 = a_5 & ~w8770;
assign w39646 = a_5 & w29210;
assign w39647 = a_5 & w8770;
assign w39648 = (w29215 & w29214) | (w29215 & w28835) | (w29214 & w28835);
assign w39649 = (w29215 & w29214) | (w29215 & w28834) | (w29214 & w28834);
assign w39650 = (w29216 & w29217) | (w29216 & ~w28835) | (w29217 & ~w28835);
assign w39651 = (w29216 & w29217) | (w29216 & ~w28834) | (w29217 & ~w28834);
assign w39652 = a_2 & ~w29218;
assign w39653 = a_2 & ~w8787;
assign w39654 = a_2 & w29218;
assign w39655 = a_2 & w8787;
assign w39656 = a_26 & ~w29232;
assign w39657 = a_26 & ~w8833;
assign w39658 = a_26 & w29232;
assign w39659 = a_26 & w8833;
assign w39660 = w8623 & ~w8619;
assign w39661 = a_32 & ~w29234;
assign w39662 = a_32 & ~w8845;
assign w39663 = a_32 & w29234;
assign w39664 = a_32 & w8845;
assign w39665 = a_38 & ~w29236;
assign w39666 = a_38 & ~w8856;
assign w39667 = a_38 & w29236;
assign w39668 = a_38 & w8856;
assign w39669 = a_41 & ~w29238;
assign w39670 = a_41 & ~w8867;
assign w39671 = a_41 & w29238;
assign w39672 = a_41 & w8867;
assign w39673 = a_44 & ~w29240;
assign w39674 = a_44 & ~w8877;
assign w39675 = a_44 & w29240;
assign w39676 = a_44 & w8877;
assign w39677 = ~w26167 & a_50;
assign w39678 = w308 & w8921;
assign w39679 = w29243 & a_47;
assign w39680 = (a_47 & w29243) | (a_47 & ~w308) | (w29243 & ~w308);
assign w39681 = a_35 & ~w29246;
assign w39682 = a_35 & ~w8959;
assign w39683 = a_35 & w29246;
assign w39684 = a_35 & w8959;
assign w39685 = a_29 & ~w29248;
assign w39686 = a_29 & ~w8982;
assign w39687 = a_29 & w29248;
assign w39688 = a_29 & w8982;
assign w39689 = w9065 & ~w9076;
assign w39690 = ~w9065 & ~w9076;
assign w39691 = ~w8758 & w8762;
assign w39692 = a_5 & ~w29260;
assign w39693 = a_5 & ~w9089;
assign w39694 = a_5 & w29260;
assign w39695 = a_5 & w9089;
assign w39696 = ~w9096 & w29263;
assign w39697 = ~w9096 & w29262;
assign w39698 = (w29267 & w29268) | (w29267 & w28835) | (w29268 & w28835);
assign w39699 = (w29267 & w29268) | (w29267 & w28834) | (w29268 & w28834);
assign w39700 = w9104 | w29271;
assign w39701 = (w29271 & w9104) | (w29271 & w9108) | (w9104 & w9108);
assign w39702 = w8799 & ~w9118;
assign w39703 = ~w8799 & w9118;
assign w39704 = (w29279 & w29278) | (w29279 & w28835) | (w29278 & w28835);
assign w39705 = (w29279 & w29278) | (w29279 & w28834) | (w29278 & w28834);
assign w39706 = (w29281 & w29280) | (w29281 & ~w28835) | (w29280 & ~w28835);
assign w39707 = (w29281 & w29280) | (w29281 & ~w28834) | (w29280 & ~w28834);
assign w39708 = a_2 & ~w29282;
assign w39709 = a_2 & ~w9128;
assign w39710 = a_2 & w29282;
assign w39711 = a_2 & w9128;
assign w39712 = a_26 & ~w29285;
assign w39713 = a_26 & ~w9158;
assign w39714 = a_26 & w29285;
assign w39715 = a_26 & w9158;
assign w39716 = a_29 & ~w29287;
assign w39717 = a_29 & ~w9169;
assign w39718 = a_29 & w29287;
assign w39719 = a_29 & w9169;
assign w39720 = a_32 & ~w29289;
assign w39721 = a_32 & ~w9179;
assign w39722 = a_32 & w29289;
assign w39723 = a_32 & w9179;
assign w39724 = a_35 & ~w29291;
assign w39725 = a_35 & ~w9190;
assign w39726 = a_35 & w29291;
assign w39727 = a_35 & w9190;
assign w39728 = a_41 & ~w29298;
assign w39729 = a_41 & ~w9212;
assign w39730 = a_41 & w29298;
assign w39731 = a_41 & w9212;
assign w39732 = a_44 & ~w29300;
assign w39733 = a_44 & ~w9223;
assign w39734 = a_44 & w29300;
assign w39735 = a_44 & w9223;
assign w39736 = a_47 & ~w29302;
assign w39737 = a_47 & ~w9234;
assign w39738 = a_47 & w29302;
assign w39739 = a_47 & w9234;
assign w39740 = a_50 & ~w29304;
assign w39741 = a_50 & ~w9244;
assign w39742 = a_50 & w29304;
assign w39743 = a_50 & w9244;
assign w39744 = a_5 & ~w29325;
assign w39745 = a_5 & ~w9427;
assign w39746 = a_5 & w29325;
assign w39747 = a_5 & w9427;
assign w39748 = a_5 & ~w29329;
assign w39749 = a_5 & ~w9450;
assign w39750 = a_5 & w29329;
assign w39751 = a_5 & w9450;
assign w39752 = a_41 & ~w29336;
assign w39753 = a_41 & ~w9473;
assign w39754 = a_41 & w29336;
assign w39755 = a_41 & w9473;
assign w39756 = a_44 & ~w29338;
assign w39757 = a_44 & ~w9484;
assign w39758 = a_44 & w29338;
assign w39759 = a_44 & w9484;
assign w39760 = a_47 & ~w29340;
assign w39761 = a_47 & ~w9495;
assign w39762 = a_47 & w29340;
assign w39763 = a_47 & w9495;
assign w39764 = a_50 & ~w29342;
assign w39765 = a_50 & ~w9506;
assign w39766 = a_50 & w29342;
assign w39767 = a_50 & w9506;
assign w39768 = a_38 & ~w29345;
assign w39769 = a_38 & ~w9582;
assign w39770 = a_38 & w29345;
assign w39771 = a_38 & w9582;
assign w39772 = a_35 & ~w29347;
assign w39773 = a_35 & ~w9599;
assign w39774 = a_35 & w29347;
assign w39775 = a_35 & w9599;
assign w39776 = a_32 & ~w29349;
assign w39777 = a_32 & ~w9617;
assign w39778 = a_32 & w29349;
assign w39779 = a_32 & w9617;
assign w39780 = w9773 & ~w29375;
assign w39781 = w9773 & ~w29376;
assign w39782 = ~w9773 & w29375;
assign w39783 = ~w9773 & w29376;
assign w39784 = a_2 & ~w29377;
assign w39785 = a_2 & ~w9769;
assign w39786 = a_2 & w29377;
assign w39787 = a_2 & w9769;
assign w39788 = (w29382 & w29383) | (w29382 & ~w29375) | (w29383 & ~w29375);
assign w39789 = (w29382 & w29383) | (w29382 & ~w29376) | (w29383 & ~w29376);
assign w39790 = (w29384 & w29385) | (w29384 & w29375) | (w29385 & w29375);
assign w39791 = (w29384 & w29385) | (w29384 & w29376) | (w29385 & w29376);
assign w39792 = a_2 & ~w29386;
assign w39793 = a_2 & ~w9792;
assign w39794 = a_2 & w29386;
assign w39795 = a_2 & w9792;
assign w39796 = a_8 & ~w29388;
assign w39797 = a_8 & ~w9810;
assign w39798 = a_8 & w29388;
assign w39799 = a_8 & w9810;
assign w39800 = a_41 & ~w29396;
assign w39801 = a_41 & ~w9845;
assign w39802 = a_41 & w29396;
assign w39803 = a_41 & w9845;
assign w39804 = a_44 & ~w29398;
assign w39805 = a_44 & ~w9856;
assign w39806 = a_44 & w29398;
assign w39807 = a_44 & w9856;
assign w39808 = a_47 & ~w29400;
assign w39809 = a_47 & ~w9867;
assign w39810 = a_47 & w29400;
assign w39811 = a_47 & w9867;
assign w39812 = ~w26175 & a_53;
assign w39813 = w308 & w9911;
assign w39814 = w29403 & a_50;
assign w39815 = (a_50 & w29403) | (a_50 & ~w308) | (w29403 & ~w308);
assign w39816 = a_38 & ~w29406;
assign w39817 = a_38 & ~w9949;
assign w39818 = a_38 & w29406;
assign w39819 = a_38 & w9949;
assign w39820 = a_35 & ~w29408;
assign w39821 = a_35 & ~w9966;
assign w39822 = a_35 & w29408;
assign w39823 = a_35 & w9966;
assign w39824 = a_29 & ~w29415;
assign w39825 = a_29 & ~w9999;
assign w39826 = a_29 & w29415;
assign w39827 = a_29 & w9999;
assign w39828 = w10105 | w29423;
assign w39829 = (w29423 & w10105) | (w29423 & w9108) | (w10105 & w9108);
assign w39830 = a_5 & ~w29425;
assign w39831 = a_5 & ~w10130;
assign w39832 = a_5 & w29425;
assign w39833 = a_5 & w10130;
assign w39834 = a_8 & ~w29427;
assign w39835 = a_8 & ~w10141;
assign w39836 = a_8 & w29427;
assign w39837 = a_8 & w10141;
assign w39838 = a_29 & ~w29431;
assign w39839 = a_29 & ~w10176;
assign w39840 = a_29 & w29431;
assign w39841 = a_29 & w10176;
assign w39842 = a_38 & ~w29433;
assign w39843 = a_38 & ~w10187;
assign w39844 = a_38 & w29433;
assign w39845 = a_38 & w10187;
assign w39846 = a_44 & ~w29440;
assign w39847 = a_44 & ~w10209;
assign w39848 = a_44 & w29440;
assign w39849 = a_44 & w10209;
assign w39850 = a_47 & ~w29442;
assign w39851 = a_47 & ~w10220;
assign w39852 = a_47 & w29442;
assign w39853 = a_47 & w10220;
assign w39854 = a_53 & ~w29444;
assign w39855 = a_53 & ~w10231;
assign w39856 = a_53 & w29444;
assign w39857 = a_53 & w10231;
assign w39858 = a_50 & ~w29446;
assign w39859 = a_50 & ~w10269;
assign w39860 = a_50 & w29446;
assign w39861 = a_50 & w10269;
assign w39862 = a_35 & ~w29448;
assign w39863 = a_35 & ~w10310;
assign w39864 = a_35 & w29448;
assign w39865 = a_35 & w10310;
assign w39866 = a_32 & ~w29450;
assign w39867 = a_32 & ~w10328;
assign w39868 = a_32 & w29450;
assign w39869 = a_32 & w10328;
assign w39870 = (w29466 & w29465) | (w29466 & ~w29375) | (w29465 & ~w29375);
assign w39871 = (w29466 & w29465) | (w29466 & ~w29376) | (w29465 & ~w29376);
assign w39872 = (w29468 & w29467) | (w29468 & w29375) | (w29467 & w29375);
assign w39873 = (w29468 & w29467) | (w29468 & w29376) | (w29467 & w29376);
assign w39874 = a_2 & ~w29469;
assign w39875 = a_2 & ~w10446;
assign w39876 = a_2 & w29469;
assign w39877 = a_2 & w10446;
assign w39878 = ~w25853 & ~w10457;
assign w39879 = (w29475 & w29474) | (w29475 & ~w29375) | (w29474 & ~w29375);
assign w39880 = (w29475 & w29474) | (w29475 & ~w29376) | (w29474 & ~w29376);
assign w39881 = (w29477 & w29476) | (w29477 & w29375) | (w29476 & w29375);
assign w39882 = (w29477 & w29476) | (w29477 & w29376) | (w29476 & w29376);
assign w39883 = a_2 & ~w29478;
assign w39884 = a_2 & ~w10470;
assign w39885 = a_2 & w29478;
assign w39886 = a_2 & w10470;
assign w39887 = a_5 & ~w29480;
assign w39888 = a_5 & ~w10486;
assign w39889 = a_5 & w29480;
assign w39890 = a_5 & w10486;
assign w39891 = a_50 & ~w29490;
assign w39892 = a_50 & ~w10523;
assign w39893 = a_50 & w29490;
assign w39894 = a_50 & w10523;
assign w39895 = a_53 & ~w29492;
assign w39896 = a_53 & ~w10534;
assign w39897 = a_53 & w29492;
assign w39898 = a_53 & w10534;
assign w39899 = a_47 & ~w29495;
assign w39900 = a_47 & ~w10598;
assign w39901 = a_47 & w29495;
assign w39902 = a_47 & w10598;
assign w39903 = a_44 & ~w29497;
assign w39904 = a_44 & ~w10615;
assign w39905 = a_44 & w29497;
assign w39906 = a_44 & w10615;
assign w39907 = a_41 & ~w29499;
assign w39908 = a_41 & ~w10633;
assign w39909 = a_41 & w29499;
assign w39910 = a_41 & w10633;
assign w39911 = a_38 & ~w29501;
assign w39912 = a_38 & ~w10650;
assign w39913 = a_38 & w29501;
assign w39914 = a_38 & w10650;
assign w39915 = ~w10458 & w10462;
assign w39916 = w10835 | w29530;
assign w39917 = (w29530 & w10835) | (w29530 & w9108) | (w10835 & w9108);
assign w39918 = a_50 & ~w29546;
assign w39919 = a_50 & ~w10893;
assign w39920 = a_50 & w29546;
assign w39921 = a_50 & w10893;
assign w39922 = ~w26824 & a_56;
assign w39923 = w308 & w10938;
assign w39924 = w29549 & a_53;
assign w39925 = (a_53 & w29549) | (a_53 & ~w308) | (w29549 & ~w308);
assign w39926 = a_41 & ~w29552;
assign w39927 = a_41 & ~w10976;
assign w39928 = a_41 & w29552;
assign w39929 = a_41 & w10976;
assign w39930 = a_38 & ~w29554;
assign w39931 = a_38 & ~w10993;
assign w39932 = a_38 & w29554;
assign w39933 = a_38 & w10993;
assign w39934 = a_5 & ~w29575;
assign w39935 = a_5 & ~w11150;
assign w39936 = a_5 & w29575;
assign w39937 = a_5 & w11150;
assign w39938 = ~w26220 & ~w11155;
assign w39939 = (w29581 & w29580) | (w29581 & ~w29375) | (w29580 & ~w29375);
assign w39940 = (w29581 & w29580) | (w29581 & ~w29376) | (w29580 & ~w29376);
assign w39941 = (w29583 & w29582) | (w29583 & w29375) | (w29582 & w29375);
assign w39942 = (w29583 & w29582) | (w29583 & w29376) | (w29582 & w29376);
assign w39943 = a_2 & ~w29584;
assign w39944 = a_2 & ~w11163;
assign w39945 = a_2 & w29584;
assign w39946 = a_2 & w11163;
assign w39947 = w11158 & w11174;
assign w39948 = ~w11158 & ~w11174;
assign w39949 = ~w11179 & w10824;
assign w39950 = ~w11179 & w29585;
assign w39951 = ~w11156 & w29588;
assign w39952 = (w29588 & ~w11156) | (w29588 & ~w11158) | (~w11156 & ~w11158);
assign w39953 = (w29592 & w29591) | (w29592 & ~w29375) | (w29591 & ~w29375);
assign w39954 = (w29592 & w29591) | (w29592 & ~w29376) | (w29591 & ~w29376);
assign w39955 = (w29593 & w29594) | (w29593 & w29375) | (w29594 & w29375);
assign w39956 = (w29593 & w29594) | (w29593 & w29376) | (w29594 & w29376);
assign w39957 = a_2 & ~w11190;
assign w39958 = a_2 & ~w29595;
assign w39959 = a_2 & w11190;
assign w39960 = a_2 & w29595;
assign w39961 = a_5 & ~w29597;
assign w39962 = a_5 & ~w11206;
assign w39963 = a_5 & w29597;
assign w39964 = a_5 & w11206;
assign w39965 = a_8 & ~w29599;
assign w39966 = a_8 & ~w11217;
assign w39967 = a_8 & w29599;
assign w39968 = a_8 & w11217;
assign w39969 = a_41 & ~w29607;
assign w39970 = a_41 & ~w11273;
assign w39971 = a_41 & w29607;
assign w39972 = a_41 & w11273;
assign w39973 = a_47 & ~w29612;
assign w39974 = a_47 & ~w11295;
assign w39975 = a_47 & w29612;
assign w39976 = a_47 & w11295;
assign w39977 = a_50 & ~w29614;
assign w39978 = a_50 & ~w11306;
assign w39979 = a_50 & w29614;
assign w39980 = a_50 & w11306;
assign w39981 = a_56 & ~w29616;
assign w39982 = a_56 & ~w11317;
assign w39983 = a_56 & w29616;
assign w39984 = a_56 & w11317;
assign w39985 = a_53 & ~w29618;
assign w39986 = a_53 & ~w11354;
assign w39987 = a_53 & w29618;
assign w39988 = a_53 & w11354;
assign w39989 = ~w11535 & ~w11178;
assign w39990 = ~w11535 & w29587;
assign w39991 = a_8 & ~w29640;
assign w39992 = a_8 & ~w11543;
assign w39993 = a_8 & w29640;
assign w39994 = a_8 & w11543;
assign w39995 = a_53 & ~w29648;
assign w39996 = a_53 & ~w11581;
assign w39997 = a_53 & w29648;
assign w39998 = a_53 & w11581;
assign w39999 = a_56 & ~w29650;
assign w40000 = a_56 & ~w11592;
assign w40001 = a_56 & w29650;
assign w40002 = a_56 & w11592;
assign w40003 = ~w26919 & a_59;
assign w40004 = a_50 & ~w29655;
assign w40005 = a_50 & ~w11656;
assign w40006 = a_50 & w29655;
assign w40007 = a_50 & w11656;
assign w40008 = a_47 & ~w29657;
assign w40009 = a_47 & ~w11673;
assign w40010 = a_47 & w29657;
assign w40011 = a_47 & w11673;
assign w40012 = a_44 & ~w29659;
assign w40013 = a_44 & ~w11691;
assign w40014 = a_44 & w29659;
assign w40015 = a_44 & w11691;
assign w40016 = a_41 & ~w29661;
assign w40017 = a_41 & ~w11707;
assign w40018 = a_41 & w29661;
assign w40019 = a_41 & w11707;
assign w40020 = a_5 & ~w29684;
assign w40021 = a_5 & ~w11882;
assign w40022 = a_5 & w29684;
assign w40023 = a_5 & w11882;
assign w40024 = (w29689 & w29688) | (w29689 & ~w29375) | (w29688 & ~w29375);
assign w40025 = (w29689 & w29688) | (w29689 & ~w29376) | (w29688 & ~w29376);
assign w40026 = (w29690 & w29691) | (w29690 & w29375) | (w29691 & w29375);
assign w40027 = (w29690 & w29691) | (w29690 & w29376) | (w29691 & w29376);
assign w40028 = a_2 & ~w29692;
assign w40029 = a_2 & ~w11895;
assign w40030 = a_2 & w29692;
assign w40031 = a_2 & w11895;
assign w40032 = a_47 & ~w29701;
assign w40033 = a_47 & ~w11939;
assign w40034 = a_47 & w29701;
assign w40035 = a_47 & w11939;
assign w40036 = a_50 & ~w29703;
assign w40037 = a_50 & ~w11949;
assign w40038 = a_50 & w29703;
assign w40039 = a_50 & w11949;
assign w40040 = a_53 & ~w29705;
assign w40041 = a_53 & ~w11960;
assign w40042 = a_53 & w29705;
assign w40043 = a_53 & w11960;
assign w40044 = ~w29707 & a_59;
assign w40045 = w308 & w12005;
assign w40046 = w29710 & a_56;
assign w40047 = (a_56 & w29710) | (a_56 & ~w308) | (w29710 & ~w308);
assign w40048 = a_44 & ~w29713;
assign w40049 = a_44 & ~w12043;
assign w40050 = a_44 & w29713;
assign w40051 = a_44 & w12043;
assign w40052 = a_41 & ~w29715;
assign w40053 = a_41 & ~w12059;
assign w40054 = a_41 & w29715;
assign w40055 = a_41 & w12059;
assign w40056 = w12221 | w29739;
assign w40057 = (w29739 & w12221) | (w29739 & w9108) | (w12221 & w9108);
assign w40058 = a_8 & ~w29741;
assign w40059 = a_8 & ~w12237;
assign w40060 = a_8 & w29741;
assign w40061 = a_8 & w12237;
assign w40062 = (w29749 & w29748) | (w29749 & ~w29375) | (w29748 & ~w29375);
assign w40063 = (w29749 & w29748) | (w29749 & ~w29376) | (w29748 & ~w29376);
assign w40064 = (w29751 & w29750) | (w29751 & w29375) | (w29750 & w29375);
assign w40065 = (w29751 & w29750) | (w29751 & w29376) | (w29750 & w29376);
assign w40066 = a_2 & ~w29752;
assign w40067 = a_2 & ~w12267;
assign w40068 = a_2 & w29752;
assign w40069 = a_2 & w12267;
assign w40070 = a_44 & ~w29767;
assign w40071 = a_44 & ~w12349;
assign w40072 = a_44 & w29767;
assign w40073 = a_44 & w12349;
assign w40074 = a_50 & ~w29769;
assign w40075 = a_50 & ~w12360;
assign w40076 = a_50 & w29769;
assign w40077 = a_50 & w12360;
assign w40078 = a_56 & ~w29772;
assign w40079 = a_56 & ~w12372;
assign w40080 = a_56 & w29772;
assign w40081 = a_56 & w12372;
assign w40082 = a_59 & ~w29774;
assign w40083 = a_59 & ~w12405;
assign w40084 = a_59 & w29774;
assign w40085 = a_59 & w12405;
assign w40086 = a_53 & ~w29776;
assign w40087 = a_53 & ~w12428;
assign w40088 = a_53 & w29776;
assign w40089 = a_53 & w12428;
assign w40090 = a_47 & ~w29778;
assign w40091 = a_47 & ~w12452;
assign w40092 = a_47 & w29778;
assign w40093 = a_47 & w12452;
assign w40094 = a_41 & ~w29780;
assign w40095 = a_41 & ~w12474;
assign w40096 = a_41 & w29780;
assign w40097 = a_41 & w12474;
assign w40098 = a_8 & ~w29803;
assign w40099 = a_8 & ~w12611;
assign w40100 = a_8 & w29803;
assign w40101 = a_8 & w12611;
assign w40102 = (w29814 & w29813) | (w29814 & ~w29375) | (w29813 & ~w29375);
assign w40103 = (w29814 & w29813) | (w29814 & ~w29376) | (w29813 & ~w29376);
assign w40104 = (w29816 & w29815) | (w29816 & w29375) | (w29815 & w29375);
assign w40105 = (w29816 & w29815) | (w29816 & w29376) | (w29815 & w29376);
assign w40106 = a_2 & ~w29817;
assign w40107 = a_2 & ~w12640;
assign w40108 = a_2 & w29817;
assign w40109 = a_2 & w12640;
assign w40110 = (w29821 & w29822) | (w29821 & ~w29375) | (w29822 & ~w29375);
assign w40111 = (w29821 & w29822) | (w29821 & ~w29376) | (w29822 & ~w29376);
assign w40112 = ~w12617 & w12628;
assign w40113 = ~w12617 & ~w27837;
assign w40114 = a_11 & ~w29828;
assign w40115 = a_11 & ~w12685;
assign w40116 = a_11 & w29828;
assign w40117 = a_11 & w12685;
assign w40118 = a_44 & ~w29842;
assign w40119 = a_44 & ~w12739;
assign w40120 = a_44 & w29842;
assign w40121 = a_44 & w12739;
assign w40122 = a_50 & ~w29844;
assign w40123 = a_50 & ~w12749;
assign w40124 = a_50 & w29844;
assign w40125 = a_50 & w12749;
assign w40126 = a_56 & ~w29846;
assign w40127 = a_56 & ~w12759;
assign w40128 = a_56 & w29846;
assign w40129 = a_56 & w12759;
assign w40130 = ~w27251 & a_62;
assign w40131 = w12777 & ~w12768;
assign w40132 = ~w12777 & ~w12768;
assign w40133 = a_59 & ~w29849;
assign w40134 = a_59 & ~w12792;
assign w40135 = a_59 & w29849;
assign w40136 = a_59 & w12792;
assign w40137 = a_53 & ~w29851;
assign w40138 = a_53 & ~w12816;
assign w40139 = a_53 & w29851;
assign w40140 = a_53 & w12816;
assign w40141 = a_47 & ~w29853;
assign w40142 = a_47 & ~w12841;
assign w40143 = a_47 & w29853;
assign w40144 = a_47 & w12841;
assign w40145 = a_41 & ~w29855;
assign w40146 = a_41 & ~w12866;
assign w40147 = a_41 & w29855;
assign w40148 = a_41 & w12866;
assign w40149 = a_8 & ~w29874;
assign w40150 = a_8 & ~w13004;
assign w40151 = a_8 & w29874;
assign w40152 = a_8 & w13004;
assign w40153 = w13041 | w29881;
assign w40154 = (w29881 & w13041) | (w29881 & w9108) | (w13041 & w9108);
assign w40155 = a_53 & ~w29885;
assign w40156 = a_53 & ~w13069;
assign w40157 = a_53 & w29885;
assign w40158 = a_53 & w13069;
assign w40159 = ~w29888 & a_62;
assign w40160 = w13088 & ~w13079;
assign w40161 = ~w13088 & ~w13079;
assign w40162 = w29889 & w27370;
assign w40163 = (w27370 & w29889) | (w27370 & w13094) | (w29889 & w13094);
assign w40164 = w29890 & ~w27370;
assign w40165 = (~w27370 & w29890) | (~w27370 & ~w13094) | (w29890 & ~w13094);
assign w40166 = w308 & w13102;
assign w40167 = w29893 & a_59;
assign w40168 = (a_59 & w29893) | (a_59 & ~w308) | (w29893 & ~w308);
assign w40169 = w12799 & w27252;
assign w40170 = ~w13110 & w27371;
assign w40171 = a_56 & ~w29896;
assign w40172 = a_56 & ~w13120;
assign w40173 = a_56 & w29896;
assign w40174 = a_56 & w13120;
assign w40175 = a_50 & ~w29898;
assign w40176 = a_50 & ~w13143;
assign w40177 = a_50 & w29898;
assign w40178 = a_50 & w13143;
assign w40179 = a_47 & ~w29900;
assign w40180 = a_47 & ~w13159;
assign w40181 = a_47 & w29900;
assign w40182 = a_47 & w13159;
assign w40183 = a_44 & ~w29902;
assign w40184 = a_44 & ~w13176;
assign w40185 = a_44 & w29902;
assign w40186 = a_44 & w13176;
assign w40187 = a_41 & ~w29904;
assign w40188 = a_41 & ~w13192;
assign w40189 = a_41 & w29904;
assign w40190 = a_41 & w13192;
assign w40191 = a_38 & ~w29906;
assign w40192 = a_38 & ~w13210;
assign w40193 = a_38 & w29906;
assign w40194 = a_38 & w13210;
assign w40195 = a_32 & ~w29913;
assign w40196 = a_32 & ~w13245;
assign w40197 = a_32 & w29913;
assign w40198 = a_32 & w13245;
assign w40199 = a_11 & ~w29934;
assign w40200 = a_11 & ~w13346;
assign w40201 = a_11 & w29934;
assign w40202 = a_11 & w13346;
assign w40203 = a_8 & ~w29936;
assign w40204 = a_8 & ~w13359;
assign w40205 = a_8 & w29936;
assign w40206 = a_8 & w13359;
assign w40207 = a_5 & ~w29939;
assign w40208 = a_5 & ~w13375;
assign w40209 = a_5 & w29939;
assign w40210 = a_5 & w13375;
assign w40211 = (w29941 & w29940) | (w29941 & ~w29375) | (w29940 & ~w29375);
assign w40212 = (w29941 & w29940) | (w29941 & ~w29376) | (w29940 & ~w29376);
assign w40213 = a_5 & ~w29945;
assign w40214 = a_5 & ~w13409;
assign w40215 = a_5 & w29945;
assign w40216 = a_5 & w13409;
assign w40217 = a_11 & ~w29947;
assign w40218 = a_11 & ~w13423;
assign w40219 = a_11 & w29947;
assign w40220 = a_11 & w13423;
assign w40221 = a_26 & ~w29961;
assign w40222 = a_26 & ~w13477;
assign w40223 = a_26 & w29961;
assign w40224 = a_26 & w13477;
assign w40225 = a_29 & w13493;
assign w40226 = a_29 & ~w29967;
assign w40227 = a_35 & ~w29971;
assign w40228 = a_35 & ~w13504;
assign w40229 = a_35 & w29971;
assign w40230 = a_35 & w13504;
assign w40231 = a_44 & ~w29973;
assign w40232 = a_44 & ~w13514;
assign w40233 = a_44 & w29973;
assign w40234 = a_44 & w13514;
assign w40235 = a_53 & ~w29975;
assign w40236 = a_53 & ~w13524;
assign w40237 = a_53 & w29975;
assign w40238 = a_53 & w13524;
assign w40239 = a_59 & ~w29983;
assign w40240 = a_59 & ~w13556;
assign w40241 = a_59 & w29983;
assign w40242 = a_59 & w13556;
assign w40243 = a_56 & ~w29985;
assign w40244 = a_56 & ~w13573;
assign w40245 = a_56 & w29985;
assign w40246 = a_56 & w13573;
assign w40247 = a_50 & ~w29990;
assign w40248 = a_50 & ~w13597;
assign w40249 = a_50 & w29990;
assign w40250 = a_50 & w13597;
assign w40251 = a_47 & ~w29993;
assign w40252 = a_47 & ~w13615;
assign w40253 = a_47 & w29993;
assign w40254 = a_47 & w13615;
assign w40255 = ~w13184 & ~w13182;
assign w40256 = a_41 & ~w29996;
assign w40257 = a_41 & ~w13640;
assign w40258 = a_41 & w29996;
assign w40259 = a_41 & w13640;
assign w40260 = a_38 & ~w29998;
assign w40261 = a_38 & ~w13658;
assign w40262 = a_38 & w29998;
assign w40263 = a_38 & w13658;
assign w40264 = a_32 & w13680;
assign w40265 = a_32 & ~w30002;
assign w40266 = a_8 & ~w30016;
assign w40267 = a_8 & ~w13735;
assign w40268 = a_8 & w30016;
assign w40269 = a_8 & w13735;
assign w40270 = a_32 & w13810;
assign w40271 = a_32 & ~w30040;
assign w40272 = a_35 & ~w30044;
assign w40273 = a_35 & ~w13821;
assign w40274 = a_35 & w30044;
assign w40275 = a_35 & w13821;
assign w40276 = a_53 & ~w30047;
assign w40277 = a_53 & ~w13832;
assign w40278 = a_53 & w30047;
assign w40279 = a_53 & w13832;
assign w40280 = a_62 & ~w30049;
assign w40281 = a_62 & ~w13842;
assign w40282 = a_62 & w30049;
assign w40283 = a_62 & w13842;
assign w40284 = a_59 & ~w30054;
assign w40285 = a_59 & ~w13867;
assign w40286 = a_59 & w30054;
assign w40287 = a_59 & w13867;
assign w40288 = a_56 & ~w30057;
assign w40289 = a_56 & ~w13885;
assign w40290 = a_56 & w30057;
assign w40291 = a_56 & w13885;
assign w40292 = a_50 & ~w30061;
assign w40293 = a_50 & ~w13911;
assign w40294 = a_50 & w30061;
assign w40295 = a_50 & w13911;
assign w40296 = a_47 & ~w30064;
assign w40297 = a_47 & ~w13929;
assign w40298 = a_47 & w30064;
assign w40299 = a_47 & w13929;
assign w40300 = a_44 & ~w30067;
assign w40301 = a_44 & ~w13948;
assign w40302 = a_44 & w30067;
assign w40303 = a_44 & w13948;
assign w40304 = ~w13956 & w13958;
assign w40305 = w13956 & ~w13958;
assign w40306 = a_41 & ~w30070;
assign w40307 = a_41 & ~w13966;
assign w40308 = a_41 & w30070;
assign w40309 = a_41 & w13966;
assign w40310 = a_38 & ~w30073;
assign w40311 = a_38 & ~w13984;
assign w40312 = a_38 & w30073;
assign w40313 = a_38 & w13984;
assign w40314 = w13995 & ~w13826;
assign w40315 = ~w13995 & ~w13826;
assign w40316 = a_29 & w14010;
assign w40317 = a_29 & ~w30077;
assign w40318 = w27792 & ~w14057;
assign w40319 = (~w14057 & w27792) | (~w14057 & ~w13702) | (w27792 & ~w13702);
assign w40320 = w13702 & w30088;
assign w40321 = a_5 & w14131;
assign w40322 = a_5 & ~w30116;
assign w40323 = a_5 & ~w14131;
assign w40324 = a_5 & w30116;
assign w40325 = ~w14164 & ~w30122;
assign w40326 = ~w14164 & ~w30121;
assign w40327 = w26336 | w26335;
assign w40328 = (w26335 & w26336) | (w26335 & w9108) | (w26336 & w9108);
assign w40329 = w26338 & w26337;
assign w40330 = (w26337 & w26338) | (w26337 & ~w9108) | (w26338 & ~w9108);
assign w40331 = ~w14190 & ~w25962;
assign w40332 = ~w14190 & w14037;
assign w40333 = ~w14190 & w25962;
assign w40334 = ~w14190 & ~w14037;
assign w40335 = w14190 & ~w25962;
assign w40336 = w14190 & w14037;
assign w40337 = w14000 & w30136;
assign w40338 = w30137 & ~w14218;
assign w40339 = (~w14218 & w30137) | (~w14218 & ~w14000) | (w30137 & ~w14000);
assign w40340 = a_35 & ~w30139;
assign w40341 = a_35 & ~w14226;
assign w40342 = a_35 & w30139;
assign w40343 = a_35 & w14226;
assign w40344 = a_47 & ~w30141;
assign w40345 = a_47 & ~w14236;
assign w40346 = a_47 & w30141;
assign w40347 = a_47 & w14236;
assign w40348 = a_56 & ~w30143;
assign w40349 = a_56 & ~w14246;
assign w40350 = a_56 & w30143;
assign w40351 = a_56 & w14246;
assign w40352 = w308 & w14256;
assign w40353 = w30145 & a_62;
assign w40354 = (a_62 & w30145) | (a_62 & ~w308) | (w30145 & ~w308);
assign w40355 = a_59 & ~w30150;
assign w40356 = a_59 & ~w14282;
assign w40357 = a_59 & w30150;
assign w40358 = a_59 & w14282;
assign w40359 = a_53 & ~w30154;
assign w40360 = a_53 & ~w14308;
assign w40361 = a_53 & w30154;
assign w40362 = a_53 & w14308;
assign w40363 = a_50 & ~w30158;
assign w40364 = a_50 & ~w14326;
assign w40365 = a_50 & w30158;
assign w40366 = a_50 & w14326;
assign w40367 = a_44 & ~w30162;
assign w40368 = a_44 & ~w14351;
assign w40369 = a_44 & w30162;
assign w40370 = a_44 & w14351;
assign w40371 = a_41 & ~w30165;
assign w40372 = a_41 & ~w14369;
assign w40373 = a_41 & w30165;
assign w40374 = a_41 & w14369;
assign w40375 = a_38 & ~w30168;
assign w40376 = a_38 & ~w14387;
assign w40377 = a_38 & w30168;
assign w40378 = a_38 & w14387;
assign w40379 = a_32 & w14409;
assign w40380 = a_32 & ~w30172;
assign w40381 = ~w14432 & ~w30182;
assign w40382 = ~w14432 & ~w30181;
assign w40383 = ~w14435 & ~w14423;
assign w40384 = a_8 & w14465;
assign w40385 = a_8 & ~w30190;
assign w40386 = ~w14468 & ~w27800;
assign w40387 = ~w14468 & ~w27799;
assign w40388 = w14471 & ~w14458;
assign w40389 = a_8 & ~w30203;
assign w40390 = a_8 & ~w14494;
assign w40391 = a_8 & w30203;
assign w40392 = a_8 & w14494;
assign w40393 = ~w14499 & ~w30204;
assign w40394 = ~w14499 & ~w30205;
assign w40395 = a_11 & ~w30207;
assign w40396 = a_11 & ~w14508;
assign w40397 = a_11 & w30207;
assign w40398 = a_11 & w14508;
assign w40399 = w14542 & w27569;
assign w40400 = w14542 & ~w14207;
assign w40401 = ~w14542 & ~w27569;
assign w40402 = ~w14542 & w14207;
assign w40403 = a_29 & ~w30225;
assign w40404 = a_29 & ~w14565;
assign w40405 = a_29 & w30225;
assign w40406 = a_29 & w14565;
assign w40407 = w14570 & ~w14220;
assign w40408 = w14570 & ~w14221;
assign w40409 = ~w14570 & w14220;
assign w40410 = ~w14570 & w14221;
assign w40411 = a_59 & ~w30234;
assign w40412 = a_59 & ~w14584;
assign w40413 = a_59 & w30234;
assign w40414 = a_59 & w14584;
assign w40415 = a_62 & ~w30239;
assign w40416 = a_62 & ~w14606;
assign w40417 = a_62 & w30239;
assign w40418 = a_62 & w14606;
assign w40419 = a_56 & ~w30242;
assign w40420 = a_56 & ~w14627;
assign w40421 = a_56 & w30242;
assign w40422 = a_56 & w14627;
assign w40423 = a_53 & ~w30247;
assign w40424 = a_53 & ~w14644;
assign w40425 = a_53 & w30247;
assign w40426 = a_53 & w14644;
assign w40427 = a_50 & ~w30249;
assign w40428 = a_50 & ~w14662;
assign w40429 = a_50 & w30249;
assign w40430 = a_50 & w14662;
assign w40431 = a_47 & ~w30253;
assign w40432 = a_47 & ~w14678;
assign w40433 = a_47 & w30253;
assign w40434 = a_47 & w14678;
assign w40435 = a_44 & ~w30255;
assign w40436 = a_44 & ~w14694;
assign w40437 = a_44 & w30255;
assign w40438 = a_44 & w14694;
assign w40439 = a_41 & ~w30258;
assign w40440 = a_41 & ~w14712;
assign w40441 = a_41 & w30258;
assign w40442 = a_41 & w14712;
assign w40443 = w30259 & ~w30229;
assign w40444 = w30259 & w14363;
assign w40445 = ~w14719 & w30260;
assign w40446 = a_38 & ~w30262;
assign w40447 = a_38 & ~w14729;
assign w40448 = a_38 & w30262;
assign w40449 = a_38 & w14729;
assign w40450 = a_35 & ~w30264;
assign w40451 = a_35 & ~w14746;
assign w40452 = a_35 & w30264;
assign w40453 = a_35 & w14746;
assign w40454 = a_32 & ~w30266;
assign w40455 = a_32 & ~w14762;
assign w40456 = a_32 & w30266;
assign w40457 = a_32 & w14762;
assign w40458 = w14531 & ~w14802;
assign w40459 = ~w14531 & ~w14802;
assign w40460 = a_14 & ~w30276;
assign w40461 = a_14 & ~w14811;
assign w40462 = a_14 & w30276;
assign w40463 = a_14 & w14811;
assign w40464 = w14502 & w14828;
assign w40465 = ~w14502 & ~w14828;
assign w40466 = ~w14831 & w14137;
assign w40467 = ~w14831 & ~w30200;
assign w40468 = w14831 & ~w14137;
assign w40469 = w14831 & w30200;
assign w40470 = a_11 & ~w30285;
assign w40471 = a_11 & ~w14853;
assign w40472 = a_11 & w30285;
assign w40473 = a_11 & w14853;
assign w40474 = ~w14871 & w14529;
assign w40475 = ~w14871 & ~w27492;
assign w40476 = w14871 & ~w14529;
assign w40477 = w14871 & w27492;
assign w40478 = a_29 & ~w30309;
assign w40479 = a_29 & ~w14935;
assign w40480 = a_29 & w30309;
assign w40481 = a_29 & w14935;
assign w40482 = ~w14940 & ~w30310;
assign w40483 = ~w14940 & w14770;
assign w40484 = a_32 & ~w30312;
assign w40485 = a_32 & ~w14948;
assign w40486 = a_32 & w30312;
assign w40487 = a_32 & w14948;
assign w40488 = a_35 & ~w30316;
assign w40489 = a_35 & ~w14961;
assign w40490 = a_35 & w30316;
assign w40491 = a_35 & w14961;
assign w40492 = a_38 & ~w30319;
assign w40493 = a_38 & ~w14972;
assign w40494 = a_38 & w30319;
assign w40495 = a_38 & w14972;
assign w40496 = a_62 & w14992;
assign w40497 = a_62 & ~w30325;
assign w40498 = a_59 & ~w30331;
assign w40499 = a_59 & ~w15005;
assign w40500 = a_59 & w30331;
assign w40501 = a_59 & w15005;
assign w40502 = a_56 & ~w30333;
assign w40503 = a_56 & ~w15023;
assign w40504 = a_56 & w30333;
assign w40505 = a_56 & w15023;
assign w40506 = a_53 & ~w30335;
assign w40507 = a_53 & ~w15041;
assign w40508 = a_53 & w30335;
assign w40509 = a_53 & w15041;
assign w40510 = a_50 & ~w30338;
assign w40511 = a_50 & ~w15059;
assign w40512 = a_50 & w30338;
assign w40513 = a_50 & w15059;
assign w40514 = a_47 & ~w30341;
assign w40515 = a_47 & ~w15078;
assign w40516 = a_47 & w30341;
assign w40517 = a_47 & w15078;
assign w40518 = a_44 & ~w30346;
assign w40519 = a_44 & ~w15095;
assign w40520 = a_44 & w30346;
assign w40521 = a_44 & w15095;
assign w40522 = a_41 & ~w30351;
assign w40523 = a_41 & ~w15112;
assign w40524 = a_41 & w30351;
assign w40525 = a_41 & w15112;
assign w40526 = w15126 & w14735;
assign w40527 = w15126 & ~w14738;
assign w40528 = ~w15126 & ~w14735;
assign w40529 = ~w15126 & w14738;
assign w40530 = a_8 & w15174;
assign w40531 = a_8 & ~w30361;
assign w40532 = a_8 & ~w15174;
assign w40533 = a_8 & w30361;
assign w40534 = w15192 & w30363;
assign w40535 = w15192 & ~w14901;
assign w40536 = ~w15192 & ~w30363;
assign w40537 = ~w15192 & w14901;
assign w40538 = a_38 & ~w30375;
assign w40539 = a_38 & ~w15244;
assign w40540 = a_38 & w30375;
assign w40541 = a_38 & w15244;
assign w40542 = a_47 & ~w30377;
assign w40543 = a_47 & ~w15254;
assign w40544 = a_47 & w30377;
assign w40545 = a_47 & w15254;
assign w40546 = a_50 & ~w30380;
assign w40547 = a_50 & ~w15265;
assign w40548 = a_50 & w30380;
assign w40549 = a_50 & w15265;
assign w40550 = ~w14984 & ~w14986;
assign w40551 = ~w14984 & ~w14993;
assign w40552 = (w30384 & w30385) | (w30384 & w14986) | (w30385 & w14986);
assign w40553 = (w30384 & w30385) | (w30384 & w14993) | (w30385 & w14993);
assign w40554 = w30388 & ~w14986;
assign w40555 = w30388 & ~w14993;
assign w40556 = a_62 & ~w30390;
assign w40557 = a_62 & ~w15286;
assign w40558 = a_62 & w30390;
assign w40559 = a_62 & w15286;
assign w40560 = a_59 & ~w30394;
assign w40561 = a_59 & ~w15299;
assign w40562 = a_59 & w30394;
assign w40563 = a_59 & w15299;
assign w40564 = a_56 & ~w30396;
assign w40565 = a_56 & ~w15315;
assign w40566 = a_56 & w30396;
assign w40567 = a_56 & w15315;
assign w40568 = a_53 & ~w30399;
assign w40569 = a_53 & ~w15333;
assign w40570 = a_53 & w30399;
assign w40571 = a_53 & w15333;
assign w40572 = ~w15341 & w15270;
assign w40573 = a_44 & ~w30403;
assign w40574 = a_44 & ~w15364;
assign w40575 = a_44 & w30403;
assign w40576 = a_44 & w15364;
assign w40577 = a_41 & ~w30406;
assign w40578 = a_41 & ~w15382;
assign w40579 = a_41 & w30406;
assign w40580 = a_41 & w15382;
assign w40581 = a_35 & ~w30412;
assign w40582 = a_35 & ~w15406;
assign w40583 = a_35 & w30412;
assign w40584 = a_35 & w15406;
assign w40585 = w30413 & ~w15412;
assign w40586 = w30416 | w30415;
assign w40587 = (w30415 & w30416) | (w30415 & ~w30413) | (w30416 & ~w30413);
assign w40588 = w30428 | w30427;
assign w40589 = (w30427 & w30428) | (w30427 & w9108) | (w30428 & w9108);
assign w40590 = w30430 & w30429;
assign w40591 = (w30429 & w30430) | (w30429 & ~w9108) | (w30430 & ~w9108);
assign w40592 = a_11 & w15489;
assign w40593 = a_11 & ~w30439;
assign w40594 = a_11 & ~w30451;
assign w40595 = a_11 & ~w15516;
assign w40596 = a_11 & w30451;
assign w40597 = a_11 & w15516;
assign w40598 = a_14 & ~w30456;
assign w40599 = a_14 & ~w15530;
assign w40600 = a_14 & w30456;
assign w40601 = a_14 & w15530;
assign w40602 = a_17 & ~w30460;
assign w40603 = a_17 & ~w15543;
assign w40604 = a_17 & w30460;
assign w40605 = a_17 & w15543;
assign w40606 = a_20 & ~w30462;
assign w40607 = a_20 & ~w15558;
assign w40608 = a_20 & w30462;
assign w40609 = a_20 & w15558;
assign w40610 = a_26 & ~w30466;
assign w40611 = a_26 & ~w15572;
assign w40612 = a_26 & w30466;
assign w40613 = a_26 & w15572;
assign w40614 = a_32 & ~w30478;
assign w40615 = a_32 & ~w15602;
assign w40616 = a_32 & w30478;
assign w40617 = a_32 & w15602;
assign w40618 = ~w15607 & ~w30476;
assign w40619 = ~w15607 & w15238;
assign w40620 = ~w15607 & w30476;
assign w40621 = ~w15607 & ~w15238;
assign w40622 = a_50 & ~w30483;
assign w40623 = a_50 & ~w15620;
assign w40624 = a_50 & w30483;
assign w40625 = a_50 & w15620;
assign w40626 = a_56 & ~w30485;
assign w40627 = a_56 & ~w15630;
assign w40628 = a_56 & w30485;
assign w40629 = a_56 & w15630;
assign w40630 = w15304 & ~w15636;
assign w40631 = a_62 & ~w30488;
assign w40632 = a_62 & ~w15642;
assign w40633 = a_62 & w30488;
assign w40634 = a_62 & w15642;
assign w40635 = (w30491 & w30490) | (w30491 & w14986) | (w30490 & w14986);
assign w40636 = (w30491 & w30490) | (w30491 & w14993) | (w30490 & w14993);
assign w40637 = (w30493 & w30492) | (w30493 & ~w14986) | (w30492 & ~w14986);
assign w40638 = (w30493 & w30492) | (w30493 & ~w14993) | (w30492 & ~w14993);
assign w40639 = a_59 & ~w30495;
assign w40640 = a_59 & ~w15667;
assign w40641 = a_59 & w30495;
assign w40642 = a_59 & w15667;
assign w40643 = a_53 & ~w30500;
assign w40644 = a_53 & ~w15690;
assign w40645 = a_53 & w30500;
assign w40646 = a_53 & w15690;
assign w40647 = a_47 & ~w30503;
assign w40648 = a_47 & ~w15716;
assign w40649 = a_47 & w30503;
assign w40650 = a_47 & w15716;
assign w40651 = a_44 & ~w30508;
assign w40652 = a_44 & ~w15733;
assign w40653 = a_44 & w30508;
assign w40654 = a_44 & w15733;
assign w40655 = a_41 & ~w30511;
assign w40656 = a_41 & ~w15750;
assign w40657 = a_41 & w30511;
assign w40658 = a_41 & w15750;
assign w40659 = a_38 & ~w30513;
assign w40660 = a_38 & ~w15767;
assign w40661 = a_38 & w30513;
assign w40662 = a_38 & w15767;
assign w40663 = a_35 & ~w30515;
assign w40664 = a_35 & ~w15783;
assign w40665 = a_35 & w30515;
assign w40666 = a_35 & w15783;
assign w40667 = ~w15790 & ~w15793;
assign w40668 = w15595 & w15801;
assign w40669 = ~w15595 & ~w15801;
assign w40670 = a_14 & ~w30533;
assign w40671 = a_14 & ~w15854;
assign w40672 = a_14 & w30533;
assign w40673 = a_14 & w15854;
assign w40674 = w30540 & w30541;
assign w40675 = (w30541 & w30540) | (w30541 & ~w15820) | (w30540 & ~w15820);
assign w40676 = w30542 | w30543;
assign w40677 = (w30543 & w30542) | (w30543 & w15820) | (w30542 & w15820);
assign w40678 = a_23 & ~w30545;
assign w40679 = a_23 & ~w15882;
assign w40680 = a_23 & w30545;
assign w40681 = a_23 & w15882;
assign w40682 = w15887 & w27586;
assign w40683 = w15887 & ~w15580;
assign w40684 = ~w15887 & ~w27586;
assign w40685 = ~w15887 & w15580;
assign w40686 = w15901 & w15593;
assign w40687 = w15901 & ~w25662;
assign w40688 = w30554 & w15793;
assign w40689 = w30554 & ~w15790;
assign w40690 = (~w15916 & w30555) | (~w15916 & ~w15793) | (w30555 & ~w15793);
assign w40691 = (~w15916 & w30555) | (~w15916 & w15790) | (w30555 & w15790);
assign w40692 = a_35 & ~w30557;
assign w40693 = a_35 & ~w15924;
assign w40694 = a_35 & w30557;
assign w40695 = a_35 & w15924;
assign w40696 = a_38 & ~w30560;
assign w40697 = a_38 & ~w15935;
assign w40698 = a_38 & w30560;
assign w40699 = a_38 & w15935;
assign w40700 = a_41 & ~w30563;
assign w40701 = a_41 & ~w15946;
assign w40702 = a_41 & w30563;
assign w40703 = a_41 & w15946;
assign w40704 = a_62 & ~w30565;
assign w40705 = a_62 & ~w15956;
assign w40706 = a_62 & w30565;
assign w40707 = a_62 & w15956;
assign w40708 = a_59 & ~w30571;
assign w40709 = a_59 & ~w15984;
assign w40710 = a_59 & w30571;
assign w40711 = a_59 & w15984;
assign w40712 = w15637 & ~w15673;
assign w40713 = a_56 & ~w30574;
assign w40714 = a_56 & ~w16002;
assign w40715 = a_56 & w30574;
assign w40716 = a_56 & w16002;
assign w40717 = a_53 & ~w30578;
assign w40718 = a_53 & ~w16019;
assign w40719 = a_53 & w30578;
assign w40720 = a_53 & w16019;
assign w40721 = a_50 & ~w30583;
assign w40722 = a_50 & ~w16036;
assign w40723 = a_50 & w30583;
assign w40724 = a_50 & w16036;
assign w40725 = a_47 & ~w30585;
assign w40726 = a_47 & ~w16054;
assign w40727 = a_47 & w30585;
assign w40728 = a_47 & w16054;
assign w40729 = a_44 & ~w30587;
assign w40730 = a_44 & ~w16072;
assign w40731 = a_44 & w30587;
assign w40732 = a_44 & w16072;
assign w40733 = ~w16086 & w15940;
assign w40734 = ~w16114 & ~w30592;
assign w40735 = ~w16114 & ~w30591;
assign w40736 = ~w16116 & ~w16105;
assign w40737 = ~w25664 & ~w16121;
assign w40738 = ~w16126 & w30596;
assign w40739 = a_17 & w16138;
assign w40740 = a_17 & ~w30599;
assign w40741 = ~w16154 | w25666;
assign w40742 = (w25666 & ~w16154) | (w25666 & w15832) | (~w16154 & w15832);
assign w40743 = ~w16162 & ~w30614;
assign w40744 = ~w16162 & ~w30613;
assign w40745 = w16165 & ~w16153;
assign w40746 = a_11 & w16180;
assign w40747 = a_11 & ~w30623;
assign w40748 = a_11 & ~w16180;
assign w40749 = a_11 & w30623;
assign w40750 = a_14 & w16194;
assign w40751 = a_14 & ~w30628;
assign w40752 = a_17 & ~w30636;
assign w40753 = a_17 & ~w16205;
assign w40754 = a_17 & w30636;
assign w40755 = a_17 & w16205;
assign w40756 = ~w16224 & w15890;
assign w40757 = ~w16224 & w15891;
assign w40758 = ~w16224 & ~w15890;
assign w40759 = ~w16224 & ~w15891;
assign w40760 = ~w15918 & w30648;
assign w40761 = a_35 & ~w30656;
assign w40762 = a_35 & ~w16271;
assign w40763 = a_35 & w30656;
assign w40764 = a_35 & w16271;
assign w40765 = a_41 & ~w30658;
assign w40766 = a_41 & ~w16282;
assign w40767 = a_41 & w30658;
assign w40768 = a_41 & w16282;
assign w40769 = a_50 & ~w30661;
assign w40770 = a_50 & ~w16293;
assign w40771 = a_50 & w30661;
assign w40772 = a_50 & w16293;
assign w40773 = a_53 & ~w30664;
assign w40774 = a_53 & ~w16304;
assign w40775 = a_53 & w30664;
assign w40776 = a_53 & w16304;
assign w40777 = a_62 & ~w30670;
assign w40778 = a_62 & ~w16327;
assign w40779 = a_62 & w30670;
assign w40780 = a_62 & w16327;
assign w40781 = a_59 & ~w30673;
assign w40782 = a_59 & ~w16341;
assign w40783 = a_59 & w30673;
assign w40784 = a_59 & w16341;
assign w40785 = a_56 & ~w30677;
assign w40786 = a_56 & ~w16358;
assign w40787 = a_56 & w30677;
assign w40788 = a_56 & w16358;
assign w40789 = a_47 & ~w30681;
assign w40790 = a_47 & ~w16386;
assign w40791 = a_47 & w30681;
assign w40792 = a_47 & w16386;
assign w40793 = a_44 & ~w30684;
assign w40794 = a_44 & ~w16404;
assign w40795 = a_44 & w30684;
assign w40796 = a_44 & w16404;
assign w40797 = a_38 & ~w30688;
assign w40798 = a_38 & ~w16429;
assign w40799 = a_38 & w30688;
assign w40800 = a_38 & w16429;
assign w40801 = w25994 | w25993;
assign w40802 = (w25993 & w25994) | (w25993 & w9108) | (w25994 & w9108);
assign w40803 = w25996 & w25995;
assign w40804 = (w25995 & w25996) | (w25995 & ~w9108) | (w25996 & ~w9108);
assign w40805 = ~w16466 & ~w16454;
assign w40806 = ~w16228 & ~w16472;
assign w40807 = a_14 & ~w30706;
assign w40808 = a_14 & ~w16500;
assign w40809 = a_14 & w30706;
assign w40810 = a_14 & w16500;
assign w40811 = a_17 & ~w30708;
assign w40812 = a_17 & ~w16513;
assign w40813 = a_17 & w30708;
assign w40814 = a_17 & w16513;
assign w40815 = a_20 & ~w30712;
assign w40816 = a_20 & ~w16526;
assign w40817 = a_20 & w30712;
assign w40818 = a_20 & w16526;
assign w40819 = w30713 & w16472;
assign w40820 = w30713 & ~w16228;
assign w40821 = (~w16531 & w30714) | (~w16531 & ~w16472) | (w30714 & ~w16472);
assign w40822 = (~w16531 & w30714) | (~w16531 & w16228) | (w30714 & w16228);
assign w40823 = a_26 & ~w30725;
assign w40824 = a_26 & ~w16554;
assign w40825 = a_26 & w30725;
assign w40826 = a_26 & w16554;
assign w40827 = a_53 & ~w30736;
assign w40828 = a_53 & ~w16588;
assign w40829 = a_53 & w30736;
assign w40830 = a_53 & w16588;
assign w40831 = a_62 & ~w30740;
assign w40832 = a_62 & ~w16599;
assign w40833 = a_62 & w30740;
assign w40834 = a_62 & w16599;
assign w40835 = a_59 & ~w30744;
assign w40836 = a_59 & ~w16626;
assign w40837 = a_59 & w30744;
assign w40838 = a_59 & w16626;
assign w40839 = a_56 & ~w30748;
assign w40840 = a_56 & ~w16644;
assign w40841 = a_56 & w30748;
assign w40842 = a_56 & w16644;
assign w40843 = a_50 & ~w30753;
assign w40844 = a_50 & ~w16669;
assign w40845 = a_50 & w30753;
assign w40846 = a_50 & w16669;
assign w40847 = a_47 & ~w30757;
assign w40848 = a_47 & ~w16687;
assign w40849 = a_47 & w30757;
assign w40850 = a_47 & w16687;
assign w40851 = a_44 & ~w30761;
assign w40852 = a_44 & ~w16705;
assign w40853 = a_44 & w30761;
assign w40854 = a_44 & w16705;
assign w40855 = a_41 & ~w30765;
assign w40856 = a_41 & ~w16721;
assign w40857 = a_41 & w30765;
assign w40858 = a_41 & w16721;
assign w40859 = a_38 & ~w30767;
assign w40860 = a_38 & ~w16737;
assign w40861 = a_38 & w30767;
assign w40862 = a_38 & w16737;
assign w40863 = a_35 & ~w30771;
assign w40864 = a_35 & ~w16753;
assign w40865 = a_35 & w30771;
assign w40866 = a_35 & w16753;
assign w40867 = ~w16791 & w30785;
assign w40868 = a_17 & ~w30797;
assign w40869 = a_17 & ~w16813;
assign w40870 = a_17 & w30797;
assign w40871 = a_17 & w16813;
assign w40872 = ~w16818 & w16533;
assign w40873 = ~w16818 & w16534;
assign w40874 = ~w16818 & ~w16533;
assign w40875 = ~w16818 & ~w16534;
assign w40876 = a_23 & ~w30800;
assign w40877 = a_23 & ~w16828;
assign w40878 = a_23 & w30800;
assign w40879 = a_23 & w16828;
assign w40880 = ~w16776 & ~w16764;
assign w40881 = ~w16776 & ~w30779;
assign w40882 = (~w16848 & w30805) | (~w16848 & w16764) | (w30805 & w16764);
assign w40883 = (~w16848 & w30805) | (~w16848 & w30779) | (w30805 & w30779);
assign w40884 = w30806 & ~w16764;
assign w40885 = w30806 & ~w30779;
assign w40886 = a_35 & ~w30808;
assign w40887 = a_35 & ~w16858;
assign w40888 = a_35 & w30808;
assign w40889 = a_35 & w16858;
assign w40890 = a_38 & ~w30811;
assign w40891 = a_38 & ~w16870;
assign w40892 = a_38 & w30811;
assign w40893 = a_38 & w16870;
assign w40894 = a_41 & ~w30814;
assign w40895 = a_41 & ~w16881;
assign w40896 = a_41 & w30814;
assign w40897 = a_41 & w16881;
assign w40898 = a_44 & ~w30817;
assign w40899 = a_44 & ~w16893;
assign w40900 = a_44 & w30817;
assign w40901 = a_44 & w16893;
assign w40902 = a_47 & ~w30819;
assign w40903 = a_47 & ~w16903;
assign w40904 = a_47 & w30819;
assign w40905 = a_47 & w16903;
assign w40906 = a_62 & ~w30824;
assign w40907 = a_62 & ~w16923;
assign w40908 = a_59 & ~w30829;
assign w40909 = a_59 & ~w16938;
assign w40910 = a_59 & w30829;
assign w40911 = a_59 & w16938;
assign w40912 = a_56 & ~w30832;
assign w40913 = a_56 & ~w16956;
assign w40914 = a_56 & w30832;
assign w40915 = a_56 & w16956;
assign w40916 = a_53 & ~w30834;
assign w40917 = a_53 & ~w16974;
assign w40918 = a_53 & w30834;
assign w40919 = a_53 & w16974;
assign w40920 = a_50 & ~w30837;
assign w40921 = a_50 & ~w16992;
assign w40922 = a_50 & w30837;
assign w40923 = a_50 & w16992;
assign w40924 = ~w30843 & ~w17046;
assign w40925 = ~w16852 & ~w17053;
assign w40926 = a_26 & w17064;
assign w40927 = a_26 & ~w30852;
assign w40928 = ~w17067 & ~w30849;
assign w40929 = ~w17067 & w17058;
assign w40930 = w17067 & w30849;
assign w40931 = w17067 & ~w17058;
assign w40932 = ~w30855 & ~w17074;
assign w40933 = a_20 & w17085;
assign w40934 = a_20 & ~w30859;
assign w40935 = ~w17088 & ~w30863;
assign w40936 = ~w17088 & ~w30862;
assign w40937 = w17091 & ~w17078;
assign w40938 = ~w17091 & ~w17078;
assign w40939 = ~w30784 & ~w17101;
assign w40940 = w17112 & ~w17100;
assign w40941 = w16506 & w17117;
assign w40942 = ~w40941 & w17117;
assign w40943 = a_14 & w17127;
assign w40944 = a_14 & ~w30878;
assign w40945 = a_14 & ~w17127;
assign w40946 = a_14 & w30878;
assign w40947 = a_20 & ~w30882;
assign w40948 = a_20 & ~w17140;
assign w40949 = a_20 & w30882;
assign w40950 = a_20 & w17140;
assign w40951 = w30883 & w17074;
assign w40952 = w30883 & ~w30855;
assign w40953 = (~w17145 & w30884) | (~w17145 & ~w17074) | (w30884 & ~w17074);
assign w40954 = (~w17145 & w30884) | (~w17145 & w30855) | (w30884 & w30855);
assign w40955 = w17167 | w30892;
assign w40956 = (w30892 & w17167) | (w30892 & w9108) | (w17167 & w9108);
assign w40957 = w30893 & w17053;
assign w40958 = w30893 & ~w16852;
assign w40959 = (~w17172 & w30894) | (~w17172 & ~w17053) | (w30894 & ~w17053);
assign w40960 = (~w17172 & w30894) | (~w17172 & w16852) | (w30894 & w16852);
assign w40961 = ~w17184 & ~w30895;
assign w40962 = ~w17184 & w17031;
assign w40963 = w17184 & w30895;
assign w40964 = w17184 & ~w17031;
assign w40965 = a_35 & ~w30899;
assign w40966 = a_35 & ~w17192;
assign w40967 = a_35 & w30899;
assign w40968 = a_35 & w17192;
assign w40969 = a_38 & ~w30902;
assign w40970 = a_38 & ~w17203;
assign w40971 = a_38 & w30902;
assign w40972 = a_38 & w17203;
assign w40973 = a_53 & ~w30907;
assign w40974 = a_53 & ~w17216;
assign w40975 = a_53 & w30907;
assign w40976 = a_53 & w17216;
assign w40977 = a_62 & w17236;
assign w40978 = a_62 & ~w30913;
assign w40979 = a_59 & ~w30918;
assign w40980 = a_59 & ~w17248;
assign w40981 = a_59 & w30918;
assign w40982 = a_59 & w17248;
assign w40983 = a_56 & ~w30921;
assign w40984 = a_56 & ~w17266;
assign w40985 = a_56 & w30921;
assign w40986 = a_56 & w17266;
assign w40987 = a_50 & ~w30923;
assign w40988 = a_50 & ~w17288;
assign w40989 = a_50 & w30923;
assign w40990 = a_50 & w17288;
assign w40991 = a_47 & ~w30926;
assign w40992 = a_47 & ~w17307;
assign w40993 = a_47 & w30926;
assign w40994 = a_47 & w17307;
assign w40995 = a_44 & ~w30928;
assign w40996 = a_44 & ~w17323;
assign w40997 = a_44 & w30928;
assign w40998 = a_44 & w17323;
assign w40999 = a_41 & ~w30931;
assign w41000 = a_41 & ~w17341;
assign w41001 = a_41 & w30931;
assign w41002 = a_41 & w17341;
assign w41003 = a_17 & w17400;
assign w41004 = a_17 & ~w30939;
assign w41005 = a_17 & ~w30953;
assign w41006 = a_17 & ~w17426;
assign w41007 = a_17 & w30953;
assign w41008 = a_17 & w17426;
assign w41009 = a_20 & ~w30957;
assign w41010 = a_20 & ~w17440;
assign w41011 = a_20 & w30957;
assign w41012 = a_20 & w17440;
assign w41013 = a_23 & ~w30961;
assign w41014 = a_23 & ~w17455;
assign w41015 = a_23 & w30961;
assign w41016 = a_23 & w17455;
assign w41017 = a_26 & ~w30963;
assign w41018 = a_26 & ~w17468;
assign w41019 = a_26 & w30963;
assign w41020 = a_26 & w17468;
assign w41021 = w17271 & ~w17260;
assign w41022 = a_62 & ~w30979;
assign w41023 = a_62 & ~w17511;
assign w41024 = a_62 & w30979;
assign w41025 = a_62 & w17511;
assign w41026 = a_59 & ~w30982;
assign w41027 = a_59 & ~w17529;
assign w41028 = a_59 & w30982;
assign w41029 = a_59 & w17529;
assign w41030 = a_56 & ~w30987;
assign w41031 = a_56 & ~w17546;
assign w41032 = a_56 & w30987;
assign w41033 = a_56 & w17546;
assign w41034 = w17495 & ~w17552;
assign w41035 = a_53 & ~w30990;
assign w41036 = a_53 & ~w17563;
assign w41037 = a_53 & w30990;
assign w41038 = a_53 & w17563;
assign w41039 = w17555 & ~w17568;
assign w41040 = ~w17555 & ~w17568;
assign w41041 = a_50 & ~w30995;
assign w41042 = a_50 & ~w17580;
assign w41043 = a_50 & w30995;
assign w41044 = a_50 & w17580;
assign w41045 = a_47 & ~w31000;
assign w41046 = a_47 & ~w17597;
assign w41047 = a_47 & w31000;
assign w41048 = a_47 & w17597;
assign w41049 = a_44 & ~w31002;
assign w41050 = a_44 & ~w17614;
assign w41051 = a_44 & w31002;
assign w41052 = a_44 & w17614;
assign w41053 = a_41 & ~w31004;
assign w41054 = a_41 & ~w17630;
assign w41055 = a_41 & w31004;
assign w41056 = a_41 & w17630;
assign w41057 = a_38 & ~w31006;
assign w41058 = a_38 & ~w17647;
assign w41059 = a_38 & w31006;
assign w41060 = a_38 & w17647;
assign w41061 = ~w17687 & w17185;
assign w41062 = ~w17687 & w17187;
assign w41063 = ~w17722 & w17448;
assign w41064 = ~w17722 & w17449;
assign w41065 = w17722 & ~w17448;
assign w41066 = w17722 & ~w17449;
assign w41067 = a_20 & ~w31029;
assign w41068 = a_20 & ~w17730;
assign w41069 = a_20 & w31029;
assign w41070 = a_20 & w17730;
assign w41071 = w17735 & w31030;
assign w41072 = w17735 & ~w17736;
assign w41073 = ~w17735 & ~w31030;
assign w41074 = ~w17735 & w17736;
assign w41075 = a_23 & w17745;
assign w41076 = a_23 & ~w31033;
assign w41077 = a_26 & ~w31039;
assign w41078 = a_26 & ~w17756;
assign w41079 = a_26 & w31039;
assign w41080 = a_26 & w17756;
assign w41081 = a_38 & ~w31047;
assign w41082 = a_38 & ~w17797;
assign w41083 = a_38 & w31047;
assign w41084 = a_38 & w17797;
assign w41085 = a_41 & ~w31049;
assign w41086 = a_41 & ~w17809;
assign w41087 = a_41 & w31049;
assign w41088 = a_41 & w17809;
assign w41089 = a_44 & ~w31051;
assign w41090 = a_44 & ~w17820;
assign w41091 = a_44 & w31051;
assign w41092 = a_44 & w17820;
assign w41093 = a_50 & ~w31053;
assign w41094 = a_50 & ~w17832;
assign w41095 = a_50 & w31053;
assign w41096 = a_50 & w17832;
assign w41097 = a_62 & w17849;
assign w41098 = a_62 & ~w31060;
assign w41099 = a_59 & ~w31070;
assign w41100 = a_59 & ~w17861;
assign w41101 = a_59 & w31070;
assign w41102 = a_59 & w17861;
assign w41103 = a_56 & ~w31072;
assign w41104 = a_56 & ~w17879;
assign w41105 = a_56 & w31072;
assign w41106 = a_56 & w17879;
assign w41107 = ~w17887 & ~w17556;
assign w41108 = w17887 & w17556;
assign w41109 = a_53 & ~w31074;
assign w41110 = a_53 & ~w17896;
assign w41111 = a_53 & w31074;
assign w41112 = a_53 & w17896;
assign w41113 = ~w17569 & w17572;
assign w41114 = ~w17569 & ~w17570;
assign w41115 = ~w17586 & w17589;
assign w41116 = ~w17586 & ~w17587;
assign w41117 = a_47 & ~w31076;
assign w41118 = a_47 & ~w17921;
assign w41119 = a_47 & w31076;
assign w41120 = a_47 & w17921;
assign w41121 = w17603 & w17929;
assign w41122 = a_35 & ~w31081;
assign w41123 = a_35 & ~w17959;
assign w41124 = a_35 & w31081;
assign w41125 = a_35 & w17959;
assign w41126 = w17987 & ~w17432;
assign w41127 = w17987 & w31085;
assign w41128 = ~w17987 & w17432;
assign w41129 = ~w17987 & ~w31085;
assign w41130 = a_17 & w17996;
assign w41131 = a_17 & ~w31094;
assign w41132 = a_17 & ~w17996;
assign w41133 = a_17 & w31094;
assign w41134 = a_20 & ~w31096;
assign w41135 = a_20 & ~w18009;
assign w41136 = a_20 & w31096;
assign w41137 = a_20 & w18009;
assign w41138 = a_23 & ~w31099;
assign w41139 = a_23 & ~w18023;
assign w41140 = a_23 & w31099;
assign w41141 = a_23 & w18023;
assign w41142 = w18051 | w26002;
assign w41143 = (w26002 & w18051) | (w26002 & w9108) | (w18051 & w9108);
assign w41144 = w26387 & w26386;
assign w41145 = (w26386 & w26387) | (w26386 & ~w9108) | (w26387 & ~w9108);
assign w41146 = w31109 | w31110;
assign w41147 = (w31110 & w31109) | (w31110 & w9108) | (w31109 & w9108);
assign w41148 = w18071 & w31116;
assign w41149 = w18071 & ~w17953;
assign w41150 = ~w18071 & ~w31116;
assign w41151 = ~w18071 & w17953;
assign w41152 = a_38 & ~w31119;
assign w41153 = a_38 & ~w18080;
assign w41154 = a_38 & w31119;
assign w41155 = a_38 & w18080;
assign w41156 = a_41 & ~w31121;
assign w41157 = a_41 & ~w18091;
assign w41158 = a_41 & w31121;
assign w41159 = a_41 & w18091;
assign w41160 = a_56 & ~w31125;
assign w41161 = a_56 & ~w18103;
assign w41162 = a_56 & w31125;
assign w41163 = a_56 & w18103;
assign w41164 = a_62 & ~w31128;
assign w41165 = a_62 & ~w18114;
assign w41166 = a_62 & w31128;
assign w41167 = a_62 & w18114;
assign w41168 = ~w17842 & ~w17843;
assign w41169 = ~w17842 & ~w17850;
assign w41170 = a_59 & ~w31137;
assign w41171 = a_59 & ~w18137;
assign w41172 = a_59 & w31137;
assign w41173 = a_59 & w18137;
assign w41174 = a_53 & ~w31139;
assign w41175 = a_53 & ~w18159;
assign w41176 = a_53 & w31139;
assign w41177 = a_53 & w18159;
assign w41178 = w17887 & ~w17556;
assign w41179 = a_50 & ~w31142;
assign w41180 = a_50 & ~w18179;
assign w41181 = a_50 & w31142;
assign w41182 = a_50 & w18179;
assign w41183 = w18173 & w18184;
assign w41184 = ~w18173 & ~w18184;
assign w41185 = a_47 & ~w31145;
assign w41186 = a_47 & ~w18196;
assign w41187 = a_47 & w31145;
assign w41188 = a_47 & w18196;
assign w41189 = a_44 & ~w31148;
assign w41190 = a_44 & ~w18214;
assign w41191 = a_44 & w31148;
assign w41192 = a_44 & w18214;
assign w41193 = a_20 & ~w31170;
assign w41194 = a_20 & ~w18284;
assign w41195 = a_20 & w31170;
assign w41196 = a_20 & w18284;
assign w41197 = a_23 & ~w31172;
assign w41198 = a_23 & ~w18297;
assign w41199 = a_23 & w31172;
assign w41200 = a_23 & w18297;
assign w41201 = a_29 & ~w31178;
assign w41202 = a_29 & ~w18310;
assign w41203 = a_29 & w31178;
assign w41204 = a_29 & w18310;
assign w41205 = a_56 & ~w31188;
assign w41206 = a_56 & ~w18327;
assign w41207 = a_56 & w31188;
assign w41208 = a_56 & w18327;
assign w41209 = a_62 & ~w31191;
assign w41210 = a_62 & ~w18338;
assign w41211 = a_62 & w31191;
assign w41212 = a_62 & w18338;
assign w41213 = a_59 & ~w31195;
assign w41214 = a_59 & ~w18364;
assign w41215 = a_59 & w31195;
assign w41216 = a_59 & w18364;
assign w41217 = a_53 & ~w31202;
assign w41218 = a_53 & ~w18387;
assign w41219 = a_53 & w31202;
assign w41220 = a_53 & w18387;
assign w41221 = a_50 & ~w31207;
assign w41222 = a_50 & ~w18404;
assign w41223 = a_50 & w31207;
assign w41224 = a_50 & w18404;
assign w41225 = ~w18409 & w18171;
assign w41226 = ~w18409 & ~w31208;
assign w41227 = a_47 & ~w31214;
assign w41228 = a_47 & ~w18418;
assign w41229 = a_47 & w31214;
assign w41230 = a_47 & w18418;
assign w41231 = a_44 & ~w31216;
assign w41232 = a_44 & ~w18434;
assign w41233 = a_44 & w31216;
assign w41234 = a_44 & w18434;
assign w41235 = a_41 & ~w31218;
assign w41236 = a_41 & ~w18451;
assign w41237 = a_41 & w31218;
assign w41238 = a_41 & w18451;
assign w41239 = a_32 & ~w31230;
assign w41240 = a_32 & ~w18502;
assign w41241 = a_32 & w31230;
assign w41242 = a_32 & w18502;
assign w41243 = a_26 & ~w31233;
assign w41244 = a_26 & ~w18524;
assign w41245 = a_26 & w31233;
assign w41246 = a_26 & w18524;
assign w41247 = ~w18045 & ~w18046;
assign w41248 = ~w18278 & ~w18268;
assign w41249 = ~w18278 & w18544;
assign w41250 = ~w18268 & ~w18544;
assign w41251 = a_23 & ~w31244;
assign w41252 = a_23 & ~w18558;
assign w41253 = a_23 & w31244;
assign w41254 = a_23 & w18558;
assign w41255 = a_26 & ~w31247;
assign w41256 = a_26 & ~w18572;
assign w41257 = a_26 & w31247;
assign w41258 = a_26 & w18572;
assign w41259 = a_29 & ~w31251;
assign w41260 = a_29 & ~w18585;
assign w41261 = a_29 & w31251;
assign w41262 = a_29 & w18585;
assign w41263 = w18590 & w31252;
assign w41264 = w18590 & ~w18509;
assign w41265 = ~w18590 & ~w31252;
assign w41266 = ~w18590 & w18509;
assign w41267 = w31258 & w18494;
assign w41268 = w31258 & ~w18492;
assign w41269 = (~w18604 & w31259) | (~w18604 & ~w18494) | (w31259 & ~w18494);
assign w41270 = (~w18604 & w31259) | (~w18604 & w18492) | (w31259 & w18492);
assign w41271 = a_41 & ~w31261;
assign w41272 = a_41 & ~w18612;
assign w41273 = a_41 & w31261;
assign w41274 = a_41 & w18612;
assign w41275 = a_44 & ~w31263;
assign w41276 = a_44 & ~w18624;
assign w41277 = a_44 & w31263;
assign w41278 = a_44 & w18624;
assign w41279 = a_53 & ~w31266;
assign w41280 = a_53 & ~w18635;
assign w41281 = a_53 & w31266;
assign w41282 = a_53 & w18635;
assign w41283 = a_59 & ~w31269;
assign w41284 = a_59 & ~w18646;
assign w41285 = a_59 & w31269;
assign w41286 = a_59 & w18646;
assign w41287 = a_62 & ~w31273;
assign w41288 = a_62 & ~w18663;
assign w41289 = a_56 & ~w31278;
assign w41290 = a_56 & ~w18685;
assign w41291 = a_56 & w31278;
assign w41292 = a_56 & w18685;
assign w41293 = ~w18393 & w18396;
assign w41294 = ~w18393 & ~w18394;
assign w41295 = a_50 & ~w31280;
assign w41296 = a_50 & ~w18710;
assign w41297 = a_50 & w31280;
assign w41298 = a_50 & w18710;
assign w41299 = a_47 & ~w31283;
assign w41300 = a_47 & ~w18729;
assign w41301 = a_47 & w31283;
assign w41302 = a_47 & w18729;
assign w41303 = a_35 & ~w31296;
assign w41304 = a_35 & ~w18776;
assign w41305 = a_35 & w31296;
assign w41306 = a_35 & w18776;
assign w41307 = a_20 & w18822;
assign w41308 = a_20 & ~w31313;
assign w41309 = a_20 & ~w18822;
assign w41310 = a_20 & w31313;
assign w41311 = a_23 & ~w31315;
assign w41312 = a_23 & ~w18835;
assign w41313 = a_23 & w31315;
assign w41314 = a_23 & w18835;
assign w41315 = w18791 & ~w18579;
assign w41316 = w31316 & ~w18840;
assign w41317 = (~w18840 & w31316) | (~w18840 & ~w18791) | (w31316 & ~w18791);
assign w41318 = a_26 & ~w31319;
assign w41319 = a_26 & ~w18850;
assign w41320 = a_26 & w31319;
assign w41321 = a_26 & w18850;
assign w41322 = ~w18607 & ~w18606;
assign w41323 = w31324 & ~w18869;
assign w41324 = (~w18869 & w31324) | (~w18869 & w18607) | (w31324 & w18607);
assign w41325 = ~w18607 & w31325;
assign w41326 = w18879 | w26392;
assign w41327 = (w26392 & w18879) | (w26392 & w9108) | (w18879 & w9108);
assign w41328 = w31328 & w31327;
assign w41329 = (w31327 & w31328) | (w31327 & ~w9108) | (w31328 & ~w9108);
assign w41330 = w31329 | w31330;
assign w41331 = (w31330 & w31329) | (w31330 & w9108) | (w31329 & w9108);
assign w41332 = w18884 & w31331;
assign w41333 = w18884 & ~w18770;
assign w41334 = ~w18884 & ~w31331;
assign w41335 = ~w18884 & w18770;
assign w41336 = a_41 & ~w31334;
assign w41337 = a_41 & ~w18893;
assign w41338 = a_41 & w31334;
assign w41339 = a_41 & w18893;
assign w41340 = a_44 & ~w31336;
assign w41341 = a_44 & ~w18904;
assign w41342 = a_44 & w31336;
assign w41343 = a_44 & w18904;
assign w41344 = a_47 & ~w31339;
assign w41345 = a_47 & ~w18915;
assign w41346 = a_47 & w31339;
assign w41347 = a_47 & w18915;
assign w41348 = a_50 & ~w31342;
assign w41349 = a_50 & ~w18926;
assign w41350 = a_50 & w31342;
assign w41351 = a_50 & w18926;
assign w41352 = a_59 & ~w31346;
assign w41353 = a_59 & ~w18938;
assign w41354 = a_59 & w31346;
assign w41355 = a_59 & w18938;
assign w41356 = a_62 & w18956;
assign w41357 = a_62 & ~w31350;
assign w41358 = a_56 & ~w31355;
assign w41359 = a_56 & ~w18974;
assign w41360 = a_56 & w31355;
assign w41361 = a_56 & w18974;
assign w41362 = a_53 & ~w31358;
assign w41363 = a_53 & ~w18994;
assign w41364 = a_53 & w31358;
assign w41365 = a_53 & w18994;
assign w41366 = a_35 & ~w31366;
assign w41367 = a_35 & ~w19052;
assign w41368 = a_35 & w31366;
assign w41369 = a_35 & w19052;
assign w41370 = a_23 & ~w31374;
assign w41371 = a_23 & ~w19088;
assign w41372 = a_23 & w31374;
assign w41373 = a_23 & w19088;
assign w41374 = ~w19093 & w18842;
assign w41375 = ~w19093 & ~w31372;
assign w41376 = ~w19093 & ~w18842;
assign w41377 = ~w19093 & w31372;
assign w41378 = a_26 & ~w31376;
assign w41379 = a_26 & ~w19102;
assign w41380 = a_26 & w31376;
assign w41381 = a_26 & w19102;
assign w41382 = a_29 & ~w31380;
assign w41383 = a_29 & ~w19117;
assign w41384 = a_29 & w31380;
assign w41385 = a_29 & w19117;
assign w41386 = a_32 & ~w31382;
assign w41387 = a_32 & ~w19130;
assign w41388 = a_32 & w31382;
assign w41389 = a_32 & w19130;
assign w41390 = a_62 & ~w31388;
assign w41391 = a_62 & ~w19155;
assign w41392 = a_62 & w31388;
assign w41393 = a_62 & w19155;
assign w41394 = a_59 & ~w31391;
assign w41395 = a_59 & ~w19174;
assign w41396 = a_59 & w31391;
assign w41397 = a_59 & w19174;
assign w41398 = ~w31392 & ~w19179;
assign w41399 = ~w19182 & w19184;
assign w41400 = w19182 & ~w19184;
assign w41401 = a_56 & ~w31395;
assign w41402 = a_56 & ~w19192;
assign w41403 = a_56 & w31395;
assign w41404 = a_56 & w19192;
assign w41405 = a_53 & ~w31400;
assign w41406 = a_53 & ~w19208;
assign w41407 = a_53 & w31400;
assign w41408 = a_53 & w19208;
assign w41409 = ~w19213 & w18986;
assign w41410 = ~w19213 & ~w31401;
assign w41411 = a_50 & ~w31407;
assign w41412 = a_50 & ~w19224;
assign w41413 = a_50 & w31407;
assign w41414 = a_50 & w19224;
assign w41415 = a_47 & ~w31409;
assign w41416 = a_47 & ~w19240;
assign w41417 = a_47 & w31409;
assign w41418 = a_47 & w19240;
assign w41419 = a_44 & ~w31414;
assign w41420 = a_44 & ~w19257;
assign w41421 = a_44 & w31414;
assign w41422 = a_44 & w19257;
assign w41423 = a_35 & ~w31431;
assign w41424 = a_35 & ~w19310;
assign w41425 = a_35 & w31431;
assign w41426 = a_35 & w19310;
assign w41427 = a_26 & ~w31448;
assign w41428 = a_26 & ~w19357;
assign w41429 = a_26 & w31448;
assign w41430 = a_26 & w19357;
assign w41431 = a_29 & w19374;
assign w41432 = a_29 & ~w31453;
assign w41433 = ~w19377 & ~w31450;
assign w41434 = ~w19377 & w19138;
assign w41435 = w19377 & w31450;
assign w41436 = w19377 & ~w19138;
assign w41437 = a_32 & ~w31457;
assign w41438 = a_32 & ~w19385;
assign w41439 = a_32 & w31457;
assign w41440 = a_32 & w19385;
assign w41441 = a_44 & ~w31461;
assign w41442 = a_44 & ~w19398;
assign w41443 = a_44 & w31461;
assign w41444 = a_44 & w19398;
assign w41445 = a_47 & ~w31463;
assign w41446 = a_47 & ~w19409;
assign w41447 = a_47 & w31463;
assign w41448 = a_47 & w19409;
assign w41449 = a_59 & ~w31467;
assign w41450 = a_59 & ~w19420;
assign w41451 = a_59 & w31467;
assign w41452 = a_59 & w19420;
assign w41453 = a_62 & w19438;
assign w41454 = a_62 & ~w31473;
assign w41455 = a_56 & ~w31487;
assign w41456 = a_56 & ~w19456;
assign w41457 = a_56 & w31487;
assign w41458 = a_56 & w19456;
assign w41459 = ~w19198 & w19200;
assign w41460 = ~w19198 & ~w31398;
assign w41461 = a_53 & ~w31489;
assign w41462 = a_53 & ~w19474;
assign w41463 = a_53 & w31489;
assign w41464 = a_53 & w19474;
assign w41465 = a_50 & ~w31492;
assign w41466 = a_50 & ~w19493;
assign w41467 = a_50 & w31492;
assign w41468 = a_50 & w19493;
assign w41469 = a_38 & ~w31505;
assign w41470 = a_38 & ~w19539;
assign w41471 = a_38 & w31505;
assign w41472 = a_38 & w19539;
assign w41473 = a_35 & ~w31507;
assign w41474 = a_35 & ~w19557;
assign w41475 = a_35 & w31507;
assign w41476 = a_35 & w19557;
assign w41477 = a_23 & w19588;
assign w41478 = a_23 & ~w31519;
assign w41479 = a_23 & ~w19588;
assign w41480 = a_23 & w31519;
assign w41481 = a_26 & ~w31521;
assign w41482 = a_26 & ~w19601;
assign w41483 = a_26 & w31521;
assign w41484 = a_26 & w19601;
assign w41485 = a_29 & ~w31524;
assign w41486 = a_29 & ~w19615;
assign w41487 = a_29 & w31524;
assign w41488 = a_29 & w19615;
assign w41489 = w19393 & ~w19621;
assign w41490 = w31526 & ~w19620;
assign w41491 = (~w19620 & w31526) | (~w19620 & ~w19393) | (w31526 & ~w19393);
assign w41492 = w19393 & w31527;
assign w41493 = w19636 & w31533;
assign w41494 = w19636 & ~w19551;
assign w41495 = ~w19636 & ~w31533;
assign w41496 = ~w19636 & w19551;
assign w41497 = w19644 | w31535;
assign w41498 = (w31535 & w19644) | (w31535 & w9108) | (w19644 & w9108);
assign w41499 = a_44 & ~w31539;
assign w41500 = a_44 & ~w19656;
assign w41501 = a_44 & w31539;
assign w41502 = a_44 & w19656;
assign w41503 = ~w19502 & w19414;
assign w41504 = ~w19502 & ~w31493;
assign w41505 = a_53 & ~w31542;
assign w41506 = a_53 & ~w19668;
assign w41507 = a_53 & w31542;
assign w41508 = a_53 & w19668;
assign w41509 = a_62 & w19687;
assign w41510 = a_62 & ~w31547;
assign w41511 = a_59 & ~w31552;
assign w41512 = a_59 & ~w19699;
assign w41513 = a_59 & w31552;
assign w41514 = a_59 & w19699;
assign w41515 = a_56 & ~w31555;
assign w41516 = a_56 & ~w19717;
assign w41517 = a_56 & w31555;
assign w41518 = a_56 & w19717;
assign w41519 = a_50 & ~w31557;
assign w41520 = a_50 & ~w19739;
assign w41521 = a_50 & w31557;
assign w41522 = a_50 & w19739;
assign w41523 = a_47 & ~w31560;
assign w41524 = a_47 & ~w19758;
assign w41525 = a_47 & w31560;
assign w41526 = a_47 & w19758;
assign w41527 = a_38 & ~w31568;
assign w41528 = a_38 & ~w19797;
assign w41529 = a_38 & w31568;
assign w41530 = a_38 & w19797;
assign w41531 = a_26 & ~w31578;
assign w41532 = a_26 & ~w19842;
assign w41533 = a_26 & w31578;
assign w41534 = a_26 & w19842;
assign w41535 = a_29 & ~w31581;
assign w41536 = a_29 & ~w19856;
assign w41537 = a_29 & w31581;
assign w41538 = a_29 & w19856;
assign w41539 = a_32 & ~w31583;
assign w41540 = a_32 & ~w19869;
assign w41541 = a_32 & w31583;
assign w41542 = a_32 & w19869;
assign w41543 = w19874 & ~w19638;
assign w41544 = w19874 & ~w19639;
assign w41545 = ~w19874 & w19638;
assign w41546 = ~w19874 & w19639;
assign w41547 = a_53 & ~w31590;
assign w41548 = a_53 & ~w19887;
assign w41549 = a_53 & w31590;
assign w41550 = a_53 & w19887;
assign w41551 = a_62 & ~w31594;
assign w41552 = a_62 & ~w19908;
assign w41553 = a_62 & w31594;
assign w41554 = a_62 & w19908;
assign w41555 = a_59 & ~w31597;
assign w41556 = a_59 & ~w19925;
assign w41557 = a_59 & w31597;
assign w41558 = a_59 & w19925;
assign w41559 = a_56 & ~w31599;
assign w41560 = a_56 & ~w19941;
assign w41561 = a_56 & w31599;
assign w41562 = a_56 & w19941;
assign w41563 = a_38 & ~w31619;
assign w41564 = a_38 & ~w20033;
assign w41565 = a_38 & w31619;
assign w41566 = a_38 & w20033;
assign w41567 = ~w31622 & ~w20039;
assign w41568 = a_35 & ~w31624;
assign w41569 = a_35 & ~w20050;
assign w41570 = a_35 & w31624;
assign w41571 = a_35 & w20050;
assign w41572 = ~w20044 & w20055;
assign w41573 = w20044 & ~w20055;
assign w41574 = w19594 & ~w20070;
assign w41575 = ~w19594 & ~w20070;
assign w41576 = a_29 & ~w31634;
assign w41577 = a_29 & ~w20084;
assign w41578 = a_29 & w31634;
assign w41579 = a_29 & w20084;
assign w41580 = a_32 & w20100;
assign w41581 = a_32 & ~w31638;
assign w41582 = w31641 & ~w20103;
assign w41583 = (~w20103 & w31641) | (~w20103 & w20058) | (w31641 & w20058);
assign w41584 = ~w20058 & w31642;
assign w41585 = w19975 & ~w19971;
assign w41586 = a_63 & b_24;
assign w41587 = a_62 & w20141;
assign w41588 = a_62 & ~w31655;
assign w41589 = a_59 & ~w31665;
assign w41590 = a_59 & ~w20153;
assign w41591 = a_59 & w31665;
assign w41592 = a_59 & w20153;
assign w41593 = a_56 & ~w31668;
assign w41594 = a_56 & ~w20171;
assign w41595 = a_56 & w31668;
assign w41596 = a_56 & w20171;
assign w41597 = a_53 & ~w31671;
assign w41598 = a_53 & ~w20189;
assign w41599 = a_53 & w31671;
assign w41600 = a_53 & w20189;
assign w41601 = a_38 & ~w31681;
assign w41602 = a_38 & ~w20257;
assign w41603 = a_38 & w31681;
assign w41604 = a_38 & w20257;
assign w41605 = a_35 & ~w31685;
assign w41606 = a_35 & ~w20273;
assign w41607 = a_35 & w31685;
assign w41608 = a_35 & w20273;
assign w41609 = ~w31686 & w20284;
assign w41610 = ~w20091 & ~w20284;
assign w41611 = ~w20091 & ~w31686;
assign w41612 = a_26 & w20313;
assign w41613 = a_26 & ~w31700;
assign w41614 = a_26 & ~w20313;
assign w41615 = a_26 & w31700;
assign w41616 = (~w20318 & w31701) | (~w20318 & w20284) | (w31701 & w20284);
assign w41617 = (~w20318 & w31701) | (~w20318 & w31686) | (w31701 & w31686);
assign w41618 = a_29 & ~w31704;
assign w41619 = a_29 & ~w20325;
assign w41620 = a_29 & w31704;
assign w41621 = a_29 & w20325;
assign w41622 = a_32 & ~w31707;
assign w41623 = a_32 & ~w20339;
assign w41624 = a_32 & w31707;
assign w41625 = a_32 & w20339;
assign w41626 = a_35 & ~w31710;
assign w41627 = a_35 & ~w20354;
assign w41628 = a_35 & w31710;
assign w41629 = a_35 & w20354;
assign w41630 = w20365 | w31713;
assign w41631 = (w31713 & w20365) | (w31713 & w9108) | (w20365 & w9108);
assign w41632 = a_56 & ~w31724;
assign w41633 = a_56 & ~w20389;
assign w41634 = a_56 & w31724;
assign w41635 = a_56 & w20389;
assign w41636 = a_59 & ~w31727;
assign w41637 = a_59 & ~w20400;
assign w41638 = a_59 & w31727;
assign w41639 = a_59 & w20400;
assign w41640 = a_62 & w20418;
assign w41641 = a_62 & ~w31731;
assign w41642 = a_53 & ~w31737;
assign w41643 = a_53 & ~w20442;
assign w41644 = a_53 & w31737;
assign w41645 = a_53 & w20442;
assign w41646 = a_50 & ~w31740;
assign w41647 = a_50 & ~w20461;
assign w41648 = a_50 & w31740;
assign w41649 = a_50 & w20461;
assign w41650 = w20226 & ~w20215;
assign w41651 = w20298 & w20532;
assign w41652 = ~w20298 & ~w20532;
assign w41653 = a_29 & ~w31756;
assign w41654 = a_29 & ~w20544;
assign w41655 = a_29 & w31756;
assign w41656 = a_29 & w20544;
assign w41657 = a_35 & ~w31760;
assign w41658 = a_35 & ~w20557;
assign w41659 = a_35 & w31760;
assign w41660 = a_35 & w20557;
assign w41661 = a_59 & ~w31765;
assign w41662 = a_59 & ~w20571;
assign w41663 = a_59 & w31765;
assign w41664 = a_59 & w20571;
assign w41665 = a_62 & ~w31771;
assign w41666 = a_62 & ~w20597;
assign w41667 = a_62 & w31771;
assign w41668 = a_62 & w20597;
assign w41669 = a_56 & ~w31773;
assign w41670 = a_56 & ~w20614;
assign w41671 = a_56 & w31773;
assign w41672 = a_56 & w20614;
assign w41673 = a_53 & ~w31778;
assign w41674 = a_53 & ~w20631;
assign w41675 = a_53 & w31778;
assign w41676 = a_53 & w20631;
assign w41677 = a_38 & ~w31800;
assign w41678 = a_38 & ~w20712;
assign w41679 = a_38 & w31800;
assign w41680 = a_38 & w20712;
assign w41681 = a_32 & ~w31805;
assign w41682 = a_32 & ~w20736;
assign w41683 = a_32 & w31805;
assign w41684 = a_32 & w20736;
assign w41685 = w2633 & b_62;
assign w41686 = ~w20766 & ~w31815;
assign w41687 = ~w20766 & w20744;
assign w41688 = w20766 & w31815;
assign w41689 = w20766 & ~w20744;
assign w41690 = a_32 & ~w31821;
assign w41691 = a_32 & ~w20774;
assign w41692 = a_32 & w31821;
assign w41693 = a_32 & w20774;
assign w41694 = a_35 & ~w31824;
assign w41695 = a_35 & ~w20788;
assign w41696 = a_35 & w31824;
assign w41697 = a_35 & w20788;
assign w41698 = ~w20637 & w20640;
assign w41699 = ~w20637 & ~w20638;
assign w41700 = a_53 & ~w31831;
assign w41701 = a_53 & ~w20810;
assign w41702 = a_53 & w31831;
assign w41703 = a_53 & w20810;
assign w41704 = a_59 & ~w31833;
assign w41705 = a_59 & ~w20821;
assign w41706 = a_59 & w31833;
assign w41707 = a_59 & w20821;
assign w41708 = a_56 & ~w31846;
assign w41709 = a_56 & ~w20861;
assign w41710 = a_56 & w31846;
assign w41711 = a_56 & w20861;
assign w41712 = a_41 & ~w31865;
assign w41713 = a_41 & ~w20928;
assign w41714 = a_41 & w31865;
assign w41715 = a_41 & w20928;
assign w41716 = a_38 & ~w31867;
assign w41717 = a_38 & ~w20945;
assign w41718 = a_38 & w31867;
assign w41719 = a_38 & w20945;
assign w41720 = (w31875 & w31874) | (w31875 & ~w29375) | (w31874 & ~w29375);
assign w41721 = (w31875 & w31874) | (w31875 & ~w29376) | (w31874 & ~w29376);
assign w41722 = a_32 & ~w31879;
assign w41723 = a_32 & ~w20990;
assign w41724 = a_32 & w31879;
assign w41725 = a_32 & w20990;
assign w41726 = a_38 & ~w31883;
assign w41727 = a_38 & ~w21006;
assign w41728 = a_38 & w31883;
assign w41729 = a_38 & w21006;
assign w41730 = w21017 | w31886;
assign w41731 = (w31886 & w21017) | (w31886 & w9108) | (w21017 & w9108);
assign w41732 = a_59 & ~w31897;
assign w41733 = a_59 & ~w21041;
assign w41734 = a_59 & w31897;
assign w41735 = a_59 & w21041;
assign w41736 = ~w20832 & ~w20833;
assign w41737 = ~w20832 & ~w31842;
assign w41738 = (w31899 & w31900) | (w31899 & w20833) | (w31900 & w20833);
assign w41739 = (w31899 & w31900) | (w31899 & w31842) | (w31900 & w31842);
assign w41740 = (w31901 & w31902) | (w31901 & ~w20833) | (w31902 & ~w20833);
assign w41741 = (w31901 & w31902) | (w31901 & ~w31842) | (w31902 & ~w31842);
assign w41742 = w31903 & ~w20833;
assign w41743 = w31903 & ~w31842;
assign w41744 = a_62 & ~w31905;
assign w41745 = a_62 & ~w21061;
assign w41746 = a_62 & w31905;
assign w41747 = a_62 & w21061;
assign w41748 = a_56 & ~w31909;
assign w41749 = a_56 & ~w21080;
assign w41750 = a_56 & w31909;
assign w41751 = a_56 & w21080;
assign w41752 = a_53 & ~w31912;
assign w41753 = a_53 & ~w21099;
assign w41754 = a_53 & w31912;
assign w41755 = a_53 & w21099;
assign w41756 = w20899 & ~w20888;
assign w41757 = a_35 & ~w31927;
assign w41758 = a_35 & ~w21164;
assign w41759 = a_35 & w31927;
assign w41760 = a_35 & w21164;
assign w41761 = a_38 & ~w31935;
assign w41762 = a_38 & ~w21192;
assign w41763 = a_38 & w31935;
assign w41764 = a_38 & w21192;
assign w41765 = ~w21146 & w21022;
assign w41766 = ~w21146 & ~w21147;
assign w41767 = w21046 & ~w21213;
assign w41768 = (w31945 & w31946) | (w31945 & w20833) | (w31946 & w20833);
assign w41769 = (w31945 & w31946) | (w31945 & w31842) | (w31946 & w31842);
assign w41770 = (w31947 & w31948) | (w31947 & ~w20833) | (w31948 & ~w20833);
assign w41771 = (w31947 & w31948) | (w31947 & ~w31842) | (w31948 & ~w31842);
assign w41772 = a_62 & ~w31950;
assign w41773 = a_62 & ~w21233;
assign w41774 = a_62 & w31950;
assign w41775 = a_62 & w21233;
assign w41776 = w21227 & w21238;
assign w41777 = ~w21227 & ~w21238;
assign w41778 = a_59 & ~w31952;
assign w41779 = a_59 & ~w21246;
assign w41780 = a_59 & w31952;
assign w41781 = a_59 & w21246;
assign w41782 = ~w21326 & ~w26414;
assign w41783 = ~w21326 & w21131;
assign w41784 = a_41 & ~w31970;
assign w41785 = a_41 & ~w21335;
assign w41786 = a_41 & w31970;
assign w41787 = a_41 & w21335;
assign w41788 = a_35 & ~w31977;
assign w41789 = a_35 & ~w21358;
assign w41790 = a_35 & w31977;
assign w41791 = a_35 & w21358;
assign w41792 = a_32 & ~w31983;
assign w41793 = a_32 & ~w21376;
assign w41794 = a_32 & w31983;
assign w41795 = a_32 & w21376;
assign w41796 = (~w21399 & w31990) | (~w21399 & ~w21367) | (w31990 & ~w21367);
assign w41797 = (~w21399 & w31990) | (~w21399 & w21365) | (w31990 & w21365);
assign w41798 = w31991 & w21367;
assign w41799 = w31991 & ~w21365;
assign w41800 = a_38 & ~w31993;
assign w41801 = a_38 & ~w21407;
assign w41802 = a_38 & w31993;
assign w41803 = a_38 & w21407;
assign w41804 = a_59 & ~w32004;
assign w41805 = a_59 & ~w21440;
assign w41806 = a_59 & w32004;
assign w41807 = a_59 & w21440;
assign w41808 = a_63 & b_30;
assign w41809 = w21464 & w21225;
assign w41810 = w21464 & ~w32005;
assign w41811 = w21464 & ~w21225;
assign w41812 = w21464 & w32005;
assign w41813 = w21278 & ~w21275;
assign w41814 = a_41 & ~w32031;
assign w41815 = a_41 & ~w21544;
assign w41816 = a_41 & w32031;
assign w41817 = a_41 & w21544;
assign w41818 = ~w21347 & w21350;
assign w41819 = ~w21347 & ~w21348;
assign w41820 = a_35 & ~w32035;
assign w41821 = a_35 & ~w21568;
assign w41822 = a_35 & w32035;
assign w41823 = a_35 & w21568;
assign w41824 = ~w21382 & ~w21370;
assign w41825 = ~w21382 & ~w31985;
assign w41826 = ~w32036 & ~w21400;
assign w41827 = a_32 & w21590;
assign w41828 = a_32 & ~w32041;
assign w41829 = a_32 & ~w21590;
assign w41830 = a_32 & w32041;
assign w41831 = ~w21595 & ~w27650;
assign w41832 = ~w21595 & w21562;
assign w41833 = ~w21595 & w27650;
assign w41834 = ~w21595 & ~w21562;
assign w41835 = w21615 | w26432;
assign w41836 = (w26432 & w21615) | (w26432 & w9108) | (w21615 & w9108);
assign w41837 = w32049 & w32048;
assign w41838 = (w32048 & w32049) | (w32048 & ~w9108) | (w32049 & ~w9108);
assign w41839 = w32050 | w32051;
assign w41840 = (w32051 & w32050) | (w32051 & w9108) | (w32050 & w9108);
assign w41841 = ~w21452 & ~w21453;
assign w41842 = ~w21452 & ~w32013;
assign w41843 = (w32062 & w32063) | (w32062 & w21453) | (w32063 & w21453);
assign w41844 = (w32062 & w32063) | (w32062 & w32013) | (w32063 & w32013);
assign w41845 = (w32064 & w32065) | (w32064 & ~w21453) | (w32065 & ~w21453);
assign w41846 = (w32064 & w32065) | (w32064 & ~w32013) | (w32065 & ~w32013);
assign w41847 = w32066 & ~w21453;
assign w41848 = w32066 & ~w32013;
assign w41849 = a_62 & ~w32068;
assign w41850 = a_62 & ~w21660;
assign w41851 = a_62 & w32068;
assign w41852 = a_62 & w21660;
assign w41853 = a_59 & ~w32071;
assign w41854 = a_59 & ~w21674;
assign w41855 = a_59 & w32071;
assign w41856 = a_59 & w21674;
assign w41857 = a_38 & ~w32083;
assign w41858 = a_38 & ~w21746;
assign w41859 = a_38 & w32083;
assign w41860 = a_38 & w21746;
assign w41861 = a_35 & ~w32086;
assign w41862 = a_35 & ~w21764;
assign w41863 = a_35 & w32086;
assign w41864 = a_35 & w21764;
assign w41865 = a_41 & ~w32095;
assign w41866 = a_41 & ~w21789;
assign w41867 = a_41 & w32095;
assign w41868 = a_41 & w21789;
assign w41869 = a_63 & b_32;
assign w41870 = (w32100 & w32101) | (w32100 & w21453) | (w32101 & w21453);
assign w41871 = (w32100 & w32101) | (w32100 & w32013) | (w32101 & w32013);
assign w41872 = (w32102 & w32103) | (w32102 & ~w21453) | (w32103 & ~w21453);
assign w41873 = (w32102 & w32103) | (w32102 & ~w32013) | (w32103 & ~w32013);
assign w41874 = a_62 & ~w32105;
assign w41875 = a_62 & ~w21823;
assign w41876 = a_62 & w32105;
assign w41877 = a_62 & w21823;
assign w41878 = ~w21883 & ~w21884;
assign w41879 = ~w21886 & ~w21898;
assign w41880 = w21886 & w21898;
assign w41881 = ~w21796 & ~w32123;
assign w41882 = ~w21796 & ~w26715;
assign w41883 = ~w21900 & w32125;
assign w41884 = ~w21900 & ~w26715;
assign w41885 = a_38 & ~w32134;
assign w41886 = a_38 & ~w21931;
assign w41887 = a_38 & w32134;
assign w41888 = a_38 & w21931;
assign w41889 = a_35 & ~w32139;
assign w41890 = a_35 & ~w21949;
assign w41891 = a_35 & w32139;
assign w41892 = a_35 & w21949;
assign w41893 = a_41 & ~w32151;
assign w41894 = a_41 & ~w21980;
assign w41895 = a_41 & w32151;
assign w41896 = a_41 & w21980;
assign w41897 = a_59 & ~w32159;
assign w41898 = a_59 & ~w22002;
assign w41899 = a_59 & w32159;
assign w41900 = a_59 & w22002;
assign w41901 = w22008 & w22007;
assign w41902 = a_47 & ~w32186;
assign w41903 = a_47 & ~w22085;
assign w41904 = a_47 & w32186;
assign w41905 = a_47 & w22085;
assign w41906 = a_44 & ~w32188;
assign w41907 = a_44 & ~w22102;
assign w41908 = a_44 & w32188;
assign w41909 = a_44 & w22102;
assign w41910 = ~w21921 & w21923;
assign w41911 = ~w21921 & ~w21922;
assign w41912 = a_38 & ~w32190;
assign w41913 = a_38 & ~w22126;
assign w41914 = a_38 & w32190;
assign w41915 = a_38 & w22126;
assign w41916 = ~w21955 & ~w21943;
assign w41917 = ~w21955 & ~w32141;
assign w41918 = a_35 & w22149;
assign w41919 = a_35 & ~w32200;
assign w41920 = a_35 & ~w22149;
assign w41921 = a_35 & w32200;
assign w41922 = a_44 & ~w32203;
assign w41923 = a_44 & ~w22164;
assign w41924 = a_44 & w32203;
assign w41925 = a_44 & w22164;
assign w41926 = w22175 | w32206;
assign w41927 = (w32206 & w22175) | (w32206 & w9108) | (w22175 & w9108);
assign w41928 = ~w22028 & w22007;
assign w41929 = ~w22028 & ~w22029;
assign w41930 = ~w22015 & ~w22016;
assign w41931 = ~w22015 & ~w32167;
assign w41932 = (w32215 & w32216) | (w32215 & w22016) | (w32216 & w22016);
assign w41933 = (w32215 & w32216) | (w32215 & w32167) | (w32216 & w32167);
assign w41934 = w32219 & ~w22016;
assign w41935 = w32219 & ~w32167;
assign one = 1;
assign f_0 = w3;// level 3
assign f_1 = w22;// level 9
assign f_2 = w44;// level 11
assign f_3 = w72;// level 12
assign f_4 = w118;// level 14
assign f_5 = w156;// level 16
assign f_6 = w201;// level 18
assign f_7 = w264;// level 20
assign f_8 = w321;// level 22
assign f_9 = w384;// level 23
assign f_10 = w465;// level 25
assign f_11 = w541;// level 26
assign f_12 = w622;// level 27
assign f_13 = w722;// level 29
assign f_14 = w814;// level 31
assign f_15 = w914;// level 33
assign f_16 = w1027;// level 34
assign f_17 = w1138;// level 35
assign f_18 = w1251;// level 37
assign f_19 = w1385;// level 39
assign f_20 = w1516;// level 41
assign f_21 = w1647;// level 42
assign f_22 = w1797;// level 44
assign f_23 = w1946;// level 45
assign f_24 = w2096;// level 47
assign f_25 = w2264;// level 48
assign f_26 = w2427;// level 50
assign f_27 = w2593;// level 51
assign f_28 = w2782;// level 53
assign f_29 = w2967;// level 55
assign f_30 = w3151;// level 57
assign f_31 = w3358;// level 59
assign f_32 = w3556;// level 60
assign f_33 = w3755;// level 62
assign f_34 = w3978;// level 63
assign f_35 = w4192;// level 64
assign f_36 = w4409;// level 66
assign f_37 = w4647;// level 67
assign f_38 = w4877;// level 69
assign f_39 = w5115;// level 71
assign f_40 = w5374;// level 72
assign f_41 = w5620;// level 74
assign f_42 = w5877;// level 76
assign f_43 = w6154;// level 77
assign f_44 = w6419;// level 79
assign f_45 = w6693;// level 81
assign f_46 = w6987;// level 83
assign f_47 = w7272;// level 84
assign f_48 = w7556;// level 86
assign f_49 = w7870;// level 88
assign f_50 = w8175;// level 91
assign f_51 = w8476;// level 92
assign f_52 = w8804;// level 93
assign f_53 = w9121;// level 94
assign f_54 = w9444;// level 96
assign f_55 = w9787;// level 97
assign f_56 = w10124;// level 98
assign f_57 = w10465;// level 100
assign f_58 = w10827;// level 101
assign f_59 = w11184;// level 102
assign f_60 = w11538;// level 103
assign f_61 = w11916;// level 105
assign f_62 = w12287;// level 106
assign f_63 = w12664;// level 107
assign f_64 = w13036;// level 108
assign f_65 = w13403;// level 109
assign f_66 = w13760;// level 109
assign f_67 = w14128;// level 110
assign f_68 = w14487;// level 111
assign f_69 = w14837;// level 111
assign f_70 = w15171;// level 111
assign f_71 = w15509;// level 111
assign f_72 = w15847;// level 111
assign f_73 = w16177;// level 111
assign f_74 = w16492;// level 111
assign f_75 = w16806;// level 111
assign f_76 = w17124;// level 111
assign f_77 = w17420;// level 111
assign f_78 = w17714;// level 111
assign f_79 = w17993;// level 111
assign f_80 = w18277;// level 111
assign f_81 = w18551;// level 111
assign f_82 = w18819;// level 111
assign f_83 = w19082;// level 111
assign f_84 = w19341;// level 111
assign f_85 = w19585;// level 111
assign f_86 = w19834;// level 111
assign f_87 = w20077;// level 111
assign f_88 = w20311;// level 111
assign f_89 = w20538;// level 111
assign f_90 = w20757;// level 110
assign f_91 = w20973;// level 110
assign f_92 = w21186;// level 110
assign f_93 = w21392;// level 110
assign f_94 = w21587;// level 110
assign f_95 = w21783;// level 110
assign f_96 = w21965;// level 110
assign f_97 = w22146;// level 110
assign f_98 = w22324;// level 110
assign f_99 = w22497;// level 110
assign f_100 = w22665;// level 110
assign f_101 = w22828;// level 110
assign f_102 = w22983;// level 110
assign f_103 = w23130;// level 110
assign f_104 = w23275;// level 110
assign f_105 = w23416;// level 110
assign f_106 = w23547;// level 110
assign f_107 = w23679;// level 110
assign f_108 = w23801;// level 110
assign f_109 = w23913;// level 110
assign f_110 = w24025;// level 110
assign f_111 = w24128;// level 110
assign f_112 = w24225;// level 110
assign f_113 = w24318;// level 110
assign f_114 = w24403;// level 110
assign f_115 = w24479;// level 110
assign f_116 = w24552;// level 110
assign f_117 = w24622;// level 110
assign f_118 = w24685;// level 110
assign f_119 = w24742;// level 110
assign f_120 = w24794;// level 110
assign f_121 = w24835;// level 110
assign f_122 = w24877;// level 110
assign f_123 = w24911;// level 110
assign f_124 = w24938;// level 110
assign f_125 = w24960;// level 110
assign f_126 = w24975;// level 110
assign f_127 = w24983;// level 110
endmodule

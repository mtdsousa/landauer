module ctrl_best_speed (
        pi0, pi1, pi2, pi3, pi4, pi5, pi6, 
        po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25);
input pi0, pi1, pi2, pi3, pi4, pi5, pi6;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126;
assign w0 = ~pi0 & ~pi2;
assign w1 = pi3 & pi4;
assign w2 = ~w0 & w1;
assign w3 = ~pi3 & ~pi4;
assign w4 = pi2 & w3;
assign w5 = pi1 & w1;
assign w6 = (pi1 & w4) | (pi1 & w5) | (w4 & w5);
assign w7 = ~w2 & ~w6;
assign w8 = ~pi2 & w1;
assign w9 = ~pi0 & ~pi1;
assign w10 = w8 & w9;
assign w11 = pi2 & ~pi4;
assign w12 = ~pi2 & pi4;
assign w13 = ~w11 & ~w12;
assign w14 = pi1 & ~pi3;
assign w15 = ~w13 & w14;
assign w16 = ~w10 & ~w15;
assign w17 = pi3 & ~pi4;
assign w18 = pi1 & w17;
assign w19 = ~pi1 & pi3;
assign w20 = ~w14 & ~w19;
assign w21 = ~pi0 & pi4;
assign w22 = ~w20 & w21;
assign w23 = ~w18 & ~w22;
assign w24 = ~pi2 & ~w23;
assign w25 = ~pi3 & pi4;
assign w26 = ~w17 & ~w21;
assign w27 = ~pi1 & ~pi2;
assign w28 = ~w26 & w27;
assign w29 = ~w25 & ~w28;
assign w30 = pi0 & ~pi6;
assign w31 = pi1 & pi5;
assign w32 = ~w30 & w31;
assign w33 = w8 & w32;
assign w34 = pi1 & ~pi2;
assign w35 = w17 & w34;
assign w36 = pi2 & w25;
assign w37 = ~w35 & ~w36;
assign w38 = pi0 & ~w37;
assign w39 = ~w33 & ~w38;
assign w40 = pi2 & ~pi3;
assign w41 = pi4 & w40;
assign w42 = pi4 & ~pi6;
assign w43 = ~pi2 & pi3;
assign w44 = ~w42 & w43;
assign w45 = ~w41 & ~w44;
assign w46 = pi1 & ~w45;
assign w47 = pi0 & pi1;
assign w48 = pi2 & pi4;
assign w49 = (pi4 & w47) | (pi4 & w48) | (w47 & w48);
assign w50 = pi3 & w49;
assign w51 = ~w17 & ~w25;
assign w52 = ~pi2 & ~w51;
assign w53 = ~w50 & ~w52;
assign w54 = pi1 & w3;
assign w55 = pi0 & w1;
assign w56 = ~w54 & ~w55;
assign w57 = pi2 & ~w56;
assign w58 = ~w10 & ~w57;
assign w59 = w0 & w25;
assign w60 = ~w1 & ~w3;
assign w61 = pi2 & ~w60;
assign w62 = ~w59 & ~w61;
assign w63 = pi1 & ~w62;
assign w64 = w1 & w27;
assign w65 = ~pi0 & w12;
assign w66 = ~pi3 & w11;
assign w67 = (~pi3 & w65) | (~pi3 & w66) | (w65 & w66);
assign w68 = pi1 & w67;
assign w69 = ~w64 & ~w68;
assign w70 = pi0 & pi4;
assign w71 = (pi4 & ~w34) | (pi4 & w70) | (~w34 & w70);
assign w72 = ~pi3 & ~w71;
assign w73 = ~pi1 & pi4;
assign w74 = pi2 & pi3;
assign w75 = (pi3 & w73) | (pi3 & w74) | (w73 & w74);
assign w76 = ~w72 & ~w75;
assign w77 = ~pi2 & w9;
assign w78 = ~pi3 & w77;
assign w79 = ~pi4 & w78;
assign w80 = pi2 & w17;
assign w81 = ~pi1 & ~pi4;
assign w82 = (~pi1 & w0) | (~pi1 & w81) | (w0 & w81);
assign w83 = ~pi2 & ~pi4;
assign w84 = ~pi3 & w83;
assign w85 = (~pi3 & w82) | (~pi3 & w84) | (w82 & w84);
assign w86 = ~w80 & ~w85;
assign w87 = ~pi4 & w40;
assign w88 = pi0 & w87;
assign w89 = ~pi0 & w87;
assign w90 = pi2 & w9;
assign w91 = pi3 & w90;
assign w92 = ~pi4 & w91;
assign w93 = pi0 & ~pi1;
assign w94 = pi2 & w93;
assign w95 = pi3 & w94;
assign w96 = ~pi4 & w95;
assign w97 = pi2 & w47;
assign w98 = pi3 & w97;
assign w99 = ~pi4 & w98;
assign w100 = ~pi0 & pi1;
assign w101 = pi2 & w100;
assign w102 = pi3 & w101;
assign w103 = ~pi4 & w102;
assign w104 = (~pi2 & w31) | (~pi2 & w83) | (w31 & w83);
assign w105 = pi0 & w104;
assign w106 = ~w47 & w48;
assign w107 = ~w105 & ~w106;
assign w108 = pi3 & ~w107;
assign w109 = pi1 & pi4;
assign w110 = pi5 & ~pi6;
assign w111 = w109 & w110;
assign w112 = pi0 & w81;
assign w113 = (pi0 & w111) | (pi0 & w112) | (w111 & w112);
assign w114 = pi3 & w113;
assign w115 = ~pi2 & w114;
assign w116 = pi5 & pi6;
assign w117 = (~pi2 & w83) | (~pi2 & w116) | (w83 & w116);
assign w118 = w47 & w117;
assign w119 = ~w106 & ~w118;
assign w120 = pi3 & ~w119;
assign w121 = ~w9 & ~w47;
assign w122 = w25 & ~w121;
assign w123 = ~pi2 & w122;
assign w124 = ~pi2 & w93;
assign w125 = ~pi3 & w124;
assign w126 = pi4 & w125;
assign one = 1;
assign po00 = ~w7;
assign po01 = ~w16;
assign po02 = w24;
assign po03 = ~w29;
assign po04 = ~w39;
assign po05 = w46;
assign po06 = ~w53;
assign po07 = ~w58;
assign po08 = w63;
assign po09 = ~w69;
assign po10 = w76;
assign po11 = w79;
assign po12 = w86;
assign po13 = w88;
assign po14 = w89;
assign po15 = w92;
assign po16 = w96;
assign po17 = w99;
assign po18 = w103;
assign po19 = w87;
assign po20 = w108;
assign po21 = w115;
assign po22 = w120;
assign po23 = one;
assign po24 = w123;
assign po25 = w126;
endmodule

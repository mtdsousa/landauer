module priority_best_speed (
        pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, 
        po0, po1, po2, po3, po4, po5, po6, po7);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127;
output po0, po1, po2, po3, po4, po5, po6, po7;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497;
assign w0 = pi035 & ~pi036;
assign w1 = pi037 & ~pi038;
assign w2 = (~pi038 & w0) | (~pi038 & w1) | (w0 & w1);
assign w3 = ~pi039 & ~pi041;
assign w4 = ~pi043 & w3;
assign w5 = ~w2 & w4;
assign w6 = ~pi029 & ~pi031;
assign w7 = ~pi033 & w6;
assign w8 = pi025 & ~pi026;
assign w9 = pi027 & ~pi028;
assign w10 = (~pi028 & w8) | (~pi028 & w9) | (w8 & w9);
assign w11 = w7 & ~w10;
assign w12 = pi015 & ~pi016;
assign w13 = pi017 & ~pi018;
assign w14 = (~pi018 & w12) | (~pi018 & w13) | (w12 & w13);
assign w15 = ~pi019 & ~w14;
assign w16 = w11 & w15;
assign w17 = ~pi021 & ~pi023;
assign w18 = w16 & w17;
assign w19 = ~pi006 & ~pi008;
assign w20 = pi001 & ~pi002;
assign w21 = pi003 & ~pi004;
assign w22 = (~pi004 & w20) | (~pi004 & w21) | (w20 & w21);
assign w23 = pi005 & w19;
assign w24 = (w19 & w22) | (w19 & w23) | (w22 & w23);
assign w25 = pi007 & ~pi008;
assign w26 = ~pi011 & ~pi013;
assign w27 = ~w25 & w26;
assign w28 = ~pi009 & w27;
assign w29 = ~w24 & w28;
assign w30 = ~pi014 & ~pi016;
assign w31 = ~pi018 & w30;
assign w32 = pi010 & ~pi011;
assign w33 = pi012 & ~pi013;
assign w34 = (~pi013 & w32) | (~pi013 & w33) | (w32 & w33);
assign w35 = w31 & ~w34;
assign w36 = ~w29 & w35;
assign w37 = w18 & ~w36;
assign w38 = ~pi024 & ~pi026;
assign w39 = ~pi028 & w38;
assign w40 = pi020 & ~pi021;
assign w41 = pi022 & ~pi023;
assign w42 = (~pi023 & w40) | (~pi023 & w41) | (w40 & w41);
assign w43 = w39 & ~w42;
assign w44 = w11 & ~w43;
assign w45 = ~pi034 & ~pi036;
assign w46 = ~pi038 & w45;
assign w47 = pi030 & ~pi031;
assign w48 = pi032 & ~pi033;
assign w49 = (~pi033 & w47) | (~pi033 & w48) | (w47 & w48);
assign w50 = w46 & ~w49;
assign w51 = w5 & ~w50;
assign w52 = (w5 & w44) | (w5 & w51) | (w44 & w51);
assign w53 = (w5 & w37) | (w5 & w52) | (w37 & w52);
assign w54 = pi060 & ~pi061;
assign w55 = pi062 & ~pi063;
assign w56 = (~pi063 & w54) | (~pi063 & w55) | (w54 & w55);
assign w57 = ~pi068 & ~pi069;
assign w58 = ~pi070 & ~pi071;
assign w59 = w57 & w58;
assign w60 = ~pi064 & ~pi065;
assign w61 = ~pi066 & ~pi067;
assign w62 = w60 & w61;
assign w63 = w59 & w62;
assign w64 = ~w56 & w63;
assign w65 = ~pi054 & ~pi056;
assign w66 = ~pi058 & w65;
assign w67 = pi050 & ~pi051;
assign w68 = pi052 & ~pi053;
assign w69 = (~pi053 & w67) | (~pi053 & w68) | (w67 & w68);
assign w70 = w66 & ~w69;
assign w71 = ~pi049 & ~pi051;
assign w72 = ~pi053 & w71;
assign w73 = pi045 & ~pi046;
assign w74 = pi047 & ~pi048;
assign w75 = (~pi048 & w73) | (~pi048 & w74) | (w73 & w74);
assign w76 = w72 & ~w75;
assign w77 = w70 & ~w76;
assign w78 = ~pi059 & ~pi061;
assign w79 = ~pi063 & w78;
assign w80 = pi055 & ~pi056;
assign w81 = pi057 & ~pi058;
assign w82 = (~pi058 & w80) | (~pi058 & w81) | (w80 & w81);
assign w83 = w79 & ~w82;
assign w84 = ~w77 & w83;
assign w85 = w64 & ~w84;
assign w86 = pi040 & ~pi041;
assign w87 = pi042 & ~pi043;
assign w88 = (~pi043 & w86) | (~pi043 & w87) | (w86 & w87);
assign w89 = ~pi044 & ~w88;
assign w90 = w70 & w89;
assign w91 = ~pi046 & ~pi048;
assign w92 = w90 & w91;
assign w93 = w84 & ~w92;
assign w94 = w64 & ~w93;
assign w95 = (~w53 & w85) | (~w53 & w94) | (w85 & w94);
assign w96 = ~pi109 & ~pi111;
assign w97 = ~pi113 & w96;
assign w98 = pi105 & ~pi106;
assign w99 = pi107 & ~pi108;
assign w100 = (~pi108 & w98) | (~pi108 & w99) | (w98 & w99);
assign w101 = w97 & ~w100;
assign w102 = pi115 & ~pi116;
assign w103 = pi117 & ~pi118;
assign w104 = (~pi118 & w102) | (~pi118 & w103) | (w102 & w103);
assign w105 = ~pi119 & ~pi121;
assign w106 = ~pi123 & ~pi125;
assign w107 = w105 & w106;
assign w108 = ~pi127 & w107;
assign w109 = ~w104 & w108;
assign w110 = w101 & w109;
assign w111 = pi090 & ~pi091;
assign w112 = pi092 & ~pi093;
assign w113 = (~pi093 & w111) | (~pi093 & w112) | (w111 & w112);
assign w114 = ~pi094 & ~w113;
assign w115 = pi085 & ~pi086;
assign w116 = pi087 & ~pi088;
assign w117 = (~pi088 & w115) | (~pi088 & w116) | (w115 & w116);
assign w118 = ~pi091 & ~pi093;
assign w119 = ~pi089 & w118;
assign w120 = ~w117 & w119;
assign w121 = w114 & ~w120;
assign w122 = pi097 & ~pi098;
assign w123 = ~pi101 & ~pi103;
assign w124 = ~w122 & w123;
assign w125 = ~pi099 & w124;
assign w126 = ~w121 & w125;
assign w127 = w110 & w126;
assign w128 = ~pi095 & w127;
assign w129 = pi075 & ~pi076;
assign w130 = pi077 & ~pi078;
assign w131 = (~pi078 & w129) | (~pi078 & w130) | (w129 & w130);
assign w132 = ~pi079 & ~pi081;
assign w133 = ~pi083 & w132;
assign w134 = ~w131 & w133;
assign w135 = pi070 & ~pi071;
assign w136 = pi072 & ~pi073;
assign w137 = (~pi073 & w135) | (~pi073 & w136) | (w135 & w136);
assign w138 = ~pi076 & ~pi078;
assign w139 = ~pi074 & w138;
assign w140 = ~w137 & w139;
assign w141 = w134 & ~w140;
assign w142 = pi080 & ~pi081;
assign w143 = pi082 & ~pi083;
assign w144 = (~pi083 & w142) | (~pi083 & w143) | (w142 & w143);
assign w145 = ~pi084 & ~w144;
assign w146 = w114 & w145;
assign w147 = ~pi086 & ~pi088;
assign w148 = w146 & w147;
assign w149 = ~w141 & w148;
assign w150 = w128 & ~w149;
assign w151 = pi065 & ~pi066;
assign w152 = pi067 & ~pi068;
assign w153 = (~pi068 & w151) | (~pi068 & w152) | (w151 & w152);
assign w154 = ~pi069 & ~w153;
assign w155 = w134 & w154;
assign w156 = ~pi071 & ~pi073;
assign w157 = w155 & w156;
assign w158 = w149 & ~w157;
assign w159 = w128 & ~w158;
assign w160 = (~w95 & w150) | (~w95 & w159) | (w150 & w159);
assign w161 = pi100 & ~pi101;
assign w162 = pi102 & ~pi103;
assign w163 = (~pi103 & w161) | (~pi103 & w162) | (w161 & w162);
assign w164 = ~pi104 & ~pi105;
assign w165 = ~pi106 & ~pi107;
assign w166 = w164 & w165;
assign w167 = ~w163 & w166;
assign w168 = ~pi108 & ~pi109;
assign w169 = ~pi110 & ~pi111;
assign w170 = w168 & w169;
assign w171 = w167 & w170;
assign w172 = w101 & ~w171;
assign w173 = ~pi096 & ~pi098;
assign w174 = w97 & ~w173;
assign w175 = ~w100 & w174;
assign w176 = w125 & w175;
assign w177 = ~w172 & ~w176;
assign w178 = pi120 & ~pi121;
assign w179 = pi122 & ~pi123;
assign w180 = (~pi123 & w178) | (~pi123 & w179) | (w178 & w179);
assign w181 = pi125 & ~pi126;
assign w182 = pi124 & ~pi125;
assign w183 = ~pi126 & ~w182;
assign w184 = (~w180 & w181) | (~w180 & w183) | (w181 & w183);
assign w185 = ~pi127 & ~w184;
assign w186 = ~w109 & ~w185;
assign w187 = pi110 & ~pi111;
assign w188 = pi112 & ~pi113;
assign w189 = (~pi113 & w187) | (~pi113 & w188) | (w187 & w188);
assign w190 = ~pi114 & ~pi116;
assign w191 = ~pi118 & w190;
assign w192 = ~w189 & w191;
assign w193 = w109 & ~w192;
assign w194 = ~w185 & ~w193;
assign w195 = (w177 & w186) | (w177 & w194) | (w186 & w194);
assign w196 = ~w160 & w195;
assign w197 = ~pi030 & ~pi031;
assign w198 = ~pi024 & ~pi025;
assign w199 = ~pi026 & ~pi027;
assign w200 = ~w198 & w199;
assign w201 = ~pi028 & ~pi029;
assign w202 = w197 & ~w201;
assign w203 = (w197 & w200) | (w197 & w202) | (w200 & w202);
assign w204 = ~pi032 & ~pi033;
assign w205 = ~pi036 & ~pi037;
assign w206 = w204 & w205;
assign w207 = ~pi040 & ~pi041;
assign w208 = w206 & w207;
assign w209 = ~w203 & w208;
assign w210 = ~pi012 & ~pi013;
assign w211 = ~pi016 & ~pi017;
assign w212 = w210 & w211;
assign w213 = ~pi020 & ~pi021;
assign w214 = w212 & w213;
assign w215 = ~pi002 & ~pi003;
assign w216 = ~pi004 & ~pi005;
assign w217 = ~w215 & w216;
assign w218 = ~pi006 & ~pi007;
assign w219 = ~w217 & w218;
assign w220 = ~pi008 & ~pi009;
assign w221 = ~pi010 & ~pi011;
assign w222 = w220 & w221;
assign w223 = ~pi010 & ~w222;
assign w224 = (~pi010 & w219) | (~pi010 & w223) | (w219 & w223);
assign w225 = pi011 & w213;
assign w226 = w212 & w225;
assign w227 = (w214 & ~w224) | (w214 & w226) | (~w224 & w226);
assign w228 = ~pi014 & ~pi015;
assign w229 = w211 & ~w228;
assign w230 = ~pi018 & ~pi019;
assign w231 = w213 & ~w230;
assign w232 = (w213 & w229) | (w213 & w231) | (w229 & w231);
assign w233 = ~pi022 & ~pi023;
assign w234 = w199 & w233;
assign w235 = w197 & w234;
assign w236 = ~w232 & w235;
assign w237 = w209 & ~w236;
assign w238 = (w209 & w227) | (w209 & w237) | (w227 & w237);
assign w239 = ~pi056 & ~pi057;
assign w240 = ~pi060 & ~pi061;
assign w241 = w239 & w240;
assign w242 = ~pi054 & ~pi055;
assign w243 = w241 & ~w242;
assign w244 = ~pi058 & ~pi059;
assign w245 = w240 & ~w244;
assign w246 = ~w243 & ~w245;
assign w247 = ~pi062 & ~pi063;
assign w248 = w61 & w247;
assign w249 = w58 & w248;
assign w250 = w246 & w249;
assign w251 = ~pi044 & ~pi045;
assign w252 = ~pi046 & ~pi047;
assign w253 = ~w251 & w252;
assign w254 = ~pi048 & ~pi049;
assign w255 = ~pi050 & ~w254;
assign w256 = (~pi050 & w253) | (~pi050 & w255) | (w253 & w255);
assign w257 = ~pi052 & ~pi053;
assign w258 = w241 & w257;
assign w259 = pi051 & ~pi053;
assign w260 = ~pi052 & w259;
assign w261 = w241 & w260;
assign w262 = (~w256 & w258) | (~w256 & w261) | (w258 & w261);
assign w263 = w250 & ~w262;
assign w264 = ~pi034 & ~pi035;
assign w265 = w205 & ~w264;
assign w266 = ~pi038 & ~pi039;
assign w267 = w207 & ~w266;
assign w268 = (w207 & w265) | (w207 & w267) | (w265 & w267);
assign w269 = ~pi042 & ~pi043;
assign w270 = w252 & w269;
assign w271 = ~pi050 & ~pi051;
assign w272 = w270 & w271;
assign w273 = ~w268 & w272;
assign w274 = w262 & ~w273;
assign w275 = w250 & ~w274;
assign w276 = (~w238 & w263) | (~w238 & w275) | (w263 & w275);
assign w277 = ~pi090 & ~pi091;
assign w278 = ~pi094 & ~pi095;
assign w279 = w277 & w278;
assign w280 = ~pi084 & ~pi085;
assign w281 = ~pi086 & ~pi087;
assign w282 = ~w280 & w281;
assign w283 = ~pi088 & ~pi089;
assign w284 = ~w282 & w283;
assign w285 = w279 & ~w284;
assign w286 = ~pi092 & ~pi093;
assign w287 = w278 & ~w286;
assign w288 = ~pi096 & ~pi097;
assign w289 = ~w287 & w288;
assign w290 = ~w285 & w289;
assign w291 = ~pi080 & ~pi081;
assign w292 = ~pi074 & ~pi075;
assign w293 = ~pi076 & ~pi077;
assign w294 = ~w292 & w293;
assign w295 = ~pi078 & ~pi079;
assign w296 = w291 & ~w295;
assign w297 = (w291 & w294) | (w291 & w296) | (w294 & w296);
assign w298 = ~pi082 & ~pi083;
assign w299 = ~pi086 & w298;
assign w300 = w279 & w299;
assign w301 = ~pi087 & w300;
assign w302 = ~w297 & w301;
assign w303 = w290 & ~w302;
assign w304 = ~w60 & w61;
assign w305 = ~w57 & w58;
assign w306 = (w58 & w304) | (w58 & w305) | (w304 & w305);
assign w307 = ~pi072 & ~pi073;
assign w308 = w293 & w307;
assign w309 = w291 & w308;
assign w310 = ~w306 & w309;
assign w311 = w302 & ~w310;
assign w312 = w290 & ~w311;
assign w313 = (~w276 & w303) | (~w276 & w312) | (w303 & w312);
assign w314 = ~pi112 & ~pi113;
assign w315 = ~pi116 & ~pi117;
assign w316 = w314 & w315;
assign w317 = ~w169 & w316;
assign w318 = ~pi114 & ~pi115;
assign w319 = w315 & ~w318;
assign w320 = ~w317 & ~w319;
assign w321 = ~pi118 & ~pi119;
assign w322 = ~pi122 & ~pi123;
assign w323 = w321 & w322;
assign w324 = ~pi126 & ~pi127;
assign w325 = ~pi102 & ~pi103;
assign w326 = w324 & w325;
assign w327 = w323 & w326;
assign w328 = ~pi098 & ~pi099;
assign w329 = w165 & w328;
assign w330 = w327 & w329;
assign w331 = w320 & w330;
assign w332 = ~w313 & w331;
assign w333 = ~pi120 & ~pi121;
assign w334 = w322 & ~w333;
assign w335 = ~pi124 & ~pi125;
assign w336 = w324 & ~w335;
assign w337 = (w324 & w334) | (w324 & w336) | (w334 & w336);
assign w338 = w323 & w324;
assign w339 = w320 & w338;
assign w340 = ~pi100 & ~pi101;
assign w341 = w325 & ~w340;
assign w342 = ~pi106 & ~w164;
assign w343 = (~pi106 & w341) | (~pi106 & w342) | (w341 & w342);
assign w344 = w168 & w316;
assign w345 = pi107 & ~pi109;
assign w346 = ~pi108 & w345;
assign w347 = w316 & w346;
assign w348 = (~w343 & w344) | (~w343 & w347) | (w344 & w347);
assign w349 = ~w337 & w348;
assign w350 = (~w337 & ~w339) | (~w337 & w349) | (~w339 & w349);
assign w351 = ~w332 & w350;
assign w352 = w251 & w252;
assign w353 = w207 & w269;
assign w354 = w352 & ~w353;
assign w355 = w254 & w271;
assign w356 = w292 & w307;
assign w357 = w355 & w356;
assign w358 = ~w354 & w357;
assign w359 = w239 & w244;
assign w360 = w62 & w359;
assign w361 = w358 & w360;
assign w362 = w213 & w233;
assign w363 = w216 & w218;
assign w364 = w222 & ~w363;
assign w365 = w210 & w228;
assign w366 = ~w364 & w365;
assign w367 = w211 & w230;
assign w368 = w213 & w367;
assign w369 = w362 & ~w368;
assign w370 = (w362 & w366) | (w362 & w369) | (w366 & w369);
assign w371 = w205 & w266;
assign w372 = w204 & w264;
assign w373 = w197 & w201;
assign w374 = w372 & ~w373;
assign w375 = w371 & ~w374;
assign w376 = w198 & w199;
assign w377 = w373 & ~w376;
assign w378 = w371 & ~w372;
assign w379 = (w371 & w377) | (w371 & w378) | (w377 & w378);
assign w380 = (w370 & w375) | (w370 & w379) | (w375 & w379);
assign w381 = ~w352 & w360;
assign w382 = w358 & w381;
assign w383 = (w361 & ~w380) | (w361 & w382) | (~w380 & w382);
assign w384 = w278 & w286;
assign w385 = w288 & w328;
assign w386 = ~w384 & w385;
assign w387 = w325 & w340;
assign w388 = w166 & ~w387;
assign w389 = (w166 & w386) | (w166 & w388) | (w386 & w388);
assign w390 = w315 & w321;
assign w391 = w170 & w390;
assign w392 = w280 & w281;
assign w393 = w391 & w392;
assign w394 = ~w389 & w393;
assign w395 = w324 & w335;
assign w396 = w394 & w395;
assign w397 = w291 & w298;
assign w398 = w396 & ~w397;
assign w399 = w242 & w257;
assign w400 = w359 & ~w399;
assign w401 = w240 & w247;
assign w402 = w62 & ~w401;
assign w403 = (w62 & w400) | (w62 & w402) | (w400 & w402);
assign w404 = w293 & w295;
assign w405 = ~w356 & w404;
assign w406 = ~w59 & w356;
assign w407 = w404 & ~w406;
assign w408 = (~w403 & w405) | (~w403 & w407) | (w405 & w407);
assign w409 = w397 & ~w408;
assign w410 = w396 & ~w409;
assign w411 = (~w383 & w398) | (~w383 & w410) | (w398 & w410);
assign w412 = w314 & w318;
assign w413 = w390 & ~w412;
assign w414 = w322 & w333;
assign w415 = ~w413 & w414;
assign w416 = w166 & w385;
assign w417 = w277 & w283;
assign w418 = w416 & w417;
assign w419 = ~w389 & ~w418;
assign w420 = ~w391 & w415;
assign w421 = (w415 & ~w419) | (w415 & w420) | (~w419 & w420);
assign w422 = w395 & ~w421;
assign w423 = ~w411 & ~w422;
assign w424 = w283 & w286;
assign w425 = w279 & w424;
assign w426 = w392 & w397;
assign w427 = w425 & ~w426;
assign w428 = w385 & w387;
assign w429 = w318 & w321;
assign w430 = w316 & w429;
assign w431 = w428 & w430;
assign w432 = ~w427 & w431;
assign w433 = w222 & w365;
assign w434 = w368 & ~w433;
assign w435 = ~w235 & w373;
assign w436 = (w373 & ~w434) | (w373 & w435) | (~w434 & w435);
assign w437 = w352 & w353;
assign w438 = w371 & w372;
assign w439 = w437 & ~w438;
assign w440 = ~w376 & w438;
assign w441 = w437 & ~w440;
assign w442 = (w436 & w439) | (w436 & w441) | (w439 & w441);
assign w443 = ~pi062 & w244;
assign w444 = w241 & w443;
assign w445 = ~pi063 & w444;
assign w446 = w63 & ~w445;
assign w447 = w355 & w399;
assign w448 = w445 & ~w447;
assign w449 = w63 & ~w448;
assign w450 = (~w442 & w446) | (~w442 & w449) | (w446 & w449);
assign w451 = w279 & w356;
assign w452 = w404 & w424;
assign w453 = w451 & w452;
assign w454 = w432 & ~w453;
assign w455 = (w432 & w450) | (w432 & w454) | (w450 & w454);
assign w456 = w166 & w170;
assign w457 = w430 & ~w456;
assign w458 = w395 & w414;
assign w459 = ~w457 & w458;
assign w460 = ~w455 & w459;
assign w461 = w316 & w395;
assign w462 = w414 & w429;
assign w463 = w461 & w462;
assign w464 = w428 & w456;
assign w465 = w235 & w368;
assign w466 = w198 & w201;
assign w467 = w465 & w466;
assign w468 = w437 & w438;
assign w469 = w447 & ~w468;
assign w470 = (w447 & w467) | (w447 & w469) | (w467 & w469);
assign w471 = w445 & w470;
assign w472 = w63 & w426;
assign w473 = w453 & w472;
assign w474 = w463 & w464;
assign w475 = w473 & w474;
assign w476 = w426 & ~w475;
assign w477 = (w426 & w471) | (w426 & w476) | (w471 & w476);
assign w478 = ~w425 & w464;
assign w479 = (w464 & ~w477) | (w464 & w478) | (~w477 & w478);
assign w480 = w463 & ~w479;
assign w481 = w437 & w447;
assign w482 = w438 & w481;
assign w483 = (w63 & w446) | (w63 & ~w482) | (w446 & ~w482);
assign w484 = w426 & w453;
assign w485 = w464 & ~w484;
assign w486 = (w464 & ~w483) | (w464 & w485) | (~w483 & w485);
assign w487 = w463 & w486;
assign w488 = w445 & w482;
assign w489 = w475 & w488;
assign w490 = ~pi000 & ~pi001;
assign w491 = ~pi002 & w490;
assign w492 = w363 & w491;
assign w493 = ~pi003 & w492;
assign w494 = w467 & w493;
assign w495 = w222 & w494;
assign w496 = w489 & w495;
assign w497 = w365 & w496;
assign one = 1;
assign po0 = w196;
assign po1 = w351;
assign po2 = w423;
assign po3 = ~w460;
assign po4 = ~w480;
assign po5 = ~w487;
assign po6 = ~w475;
assign po7 = ~w497;
endmodule

// Benchmark "i9" written by ABC on Sun Apr 22 21:43:05 2018

module i9 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84, pi85, pi86, pi87,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84, pi85, pi86, pi87;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62;
  wire n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n370, n371, n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n548, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039;
  assign n152 = ~pi01 & pi03;
  assign n153 = ~pi02 & n152;
  assign n154 = ~pi01 & pi07;
  assign n155 = ~pi02 & n154;
  assign n156 = ~pi02 & ~pi06;
  assign n157 = ~pi01 & n156;
  assign n158 = ~pi05 & n157;
  assign n159 = pi02 & pi03;
  assign n160 = pi01 & pi03;
  assign n161 = pi00 & pi01;
  assign n162 = pi02 & n161;
  assign n163 = ~pi03 & ~pi04;
  assign n164 = pi07 & n163;
  assign n165 = ~pi05 & n163;
  assign n166 = ~pi03 & ~pi05;
  assign n167 = pi01 & n166;
  assign n168 = ~pi02 & n167;
  assign n169 = ~pi06 & n168;
  assign n170 = pi01 & ~pi03;
  assign n171 = pi08 & n170;
  assign n172 = pi02 & ~pi03;
  assign n173 = pi01 & n172;
  assign n174 = ~pi00 & n173;
  assign n175 = ~pi01 & n166;
  assign n176 = pi04 & n175;
  assign n177 = pi02 & n176;
  assign n178 = ~pi06 & n177;
  assign n179 = ~pi01 & n172;
  assign n180 = pi08 & n179;
  assign n181 = ~n174 & ~n178;
  assign n182 = ~n180 & n181;
  assign n183 = ~n165 & ~n169;
  assign n184 = ~n171 & n183;
  assign n185 = n182 & n184;
  assign n186 = ~n160 & ~n162;
  assign n187 = ~n164 & n186;
  assign n188 = ~n158 & ~n159;
  assign n189 = ~n153 & ~n155;
  assign n190 = n188 & n189;
  assign n191 = n187 & n190;
  assign n192 = n185 & n191;
  assign n193 = ~n155 & ~n158;
  assign n194 = ~n153 & n193;
  assign n195 = ~n164 & ~n171;
  assign n196 = n183 & n195;
  assign n197 = n194 & n196;
  assign n198 = ~n178 & ~n180;
  assign n199 = ~n174 & n198;
  assign n200 = n194 & n199;
  assign n201 = pi09 & n197;
  assign n202 = n200 & n201;
  assign n203 = ~n192 & n202;
  assign n204 = ~n192 & n200;
  assign n205 = ~n197 & n204;
  assign n206 = pi17 & n205;
  assign n207 = pi20 & n197;
  assign n208 = ~n200 & n207;
  assign n209 = ~n192 & n208;
  assign n210 = pi24 & ~n197;
  assign n211 = ~n200 & n210;
  assign n212 = ~n192 & n211;
  assign n213 = ~n209 & ~n212;
  assign n214 = ~n192 & ~n203;
  assign n215 = ~n206 & n214;
  assign po00 = ~n213 | ~n215;
  assign n217 = pi10 & n197;
  assign n218 = n200 & n217;
  assign n219 = ~n192 & n218;
  assign n220 = pi18 & n205;
  assign n221 = pi21 & n197;
  assign n222 = ~n200 & n221;
  assign n223 = ~n192 & n222;
  assign n224 = pi25 & ~n197;
  assign n225 = ~n200 & n224;
  assign n226 = ~n192 & n225;
  assign n227 = ~n223 & ~n226;
  assign n228 = ~n192 & ~n219;
  assign n229 = ~n220 & n228;
  assign po01 = ~n227 | ~n229;
  assign n231 = pi11 & n197;
  assign n232 = n200 & n231;
  assign n233 = ~n192 & n232;
  assign n234 = pi19 & n205;
  assign n235 = pi22 & n197;
  assign n236 = ~n200 & n235;
  assign n237 = ~n192 & n236;
  assign n238 = pi26 & ~n197;
  assign n239 = ~n200 & n238;
  assign n240 = ~n192 & n239;
  assign n241 = ~n237 & ~n240;
  assign n242 = ~n192 & ~n233;
  assign n243 = ~n234 & n242;
  assign po02 = ~n241 | ~n243;
  assign n245 = pi12 & n197;
  assign n246 = n200 & n245;
  assign n247 = ~n192 & n246;
  assign n248 = pi20 & n205;
  assign n249 = pi23 & n197;
  assign n250 = ~n200 & n249;
  assign n251 = ~n192 & n250;
  assign n252 = pi27 & ~n197;
  assign n253 = ~n200 & n252;
  assign n254 = ~n192 & n253;
  assign n255 = ~n251 & ~n254;
  assign n256 = ~n192 & ~n247;
  assign n257 = ~n248 & n256;
  assign po03 = ~n255 | ~n257;
  assign n259 = pi13 & n197;
  assign n260 = n200 & n259;
  assign n261 = ~n192 & n260;
  assign n262 = pi21 & n205;
  assign n263 = pi24 & n197;
  assign n264 = ~n200 & n263;
  assign n265 = ~n192 & n264;
  assign n266 = pi28 & ~n197;
  assign n267 = ~n200 & n266;
  assign n268 = ~n192 & n267;
  assign n269 = ~n265 & ~n268;
  assign n270 = ~n192 & ~n261;
  assign n271 = ~n262 & n270;
  assign po04 = ~n269 | ~n271;
  assign n273 = pi14 & n197;
  assign n274 = n200 & n273;
  assign n275 = ~n192 & n274;
  assign n276 = pi22 & n205;
  assign n277 = pi25 & n197;
  assign n278 = ~n200 & n277;
  assign n279 = ~n192 & n278;
  assign n280 = pi29 & ~n197;
  assign n281 = ~n200 & n280;
  assign n282 = ~n192 & n281;
  assign n283 = ~n279 & ~n282;
  assign n284 = ~n192 & ~n275;
  assign n285 = ~n276 & n284;
  assign po05 = ~n283 | ~n285;
  assign n287 = pi15 & n197;
  assign n288 = n200 & n287;
  assign n289 = ~n192 & n288;
  assign n290 = pi23 & n205;
  assign n291 = pi26 & n197;
  assign n292 = ~n200 & n291;
  assign n293 = ~n192 & n292;
  assign n294 = pi30 & ~n197;
  assign n295 = ~n200 & n294;
  assign n296 = ~n192 & n295;
  assign n297 = ~n293 & ~n296;
  assign n298 = ~n192 & ~n289;
  assign n299 = ~n290 & n298;
  assign po06 = ~n297 | ~n299;
  assign n301 = pi16 & n197;
  assign n302 = n200 & n301;
  assign n303 = ~n192 & n302;
  assign n304 = pi24 & n205;
  assign n305 = pi27 & n197;
  assign n306 = ~n200 & n305;
  assign n307 = ~n192 & n306;
  assign n308 = pi31 & ~n197;
  assign n309 = ~n200 & n308;
  assign n310 = ~n192 & n309;
  assign n311 = ~n307 & ~n310;
  assign n312 = ~n192 & ~n303;
  assign n313 = ~n304 & n312;
  assign po07 = ~n311 | ~n313;
  assign n315 = pi17 & n197;
  assign n316 = n200 & n315;
  assign n317 = ~n192 & n316;
  assign n318 = pi25 & n205;
  assign n319 = pi28 & n197;
  assign n320 = ~n200 & n319;
  assign n321 = ~n192 & n320;
  assign n322 = pi32 & ~n197;
  assign n323 = ~n200 & n322;
  assign n324 = ~n192 & n323;
  assign n325 = ~n321 & ~n324;
  assign n326 = ~n192 & ~n317;
  assign n327 = ~n318 & n326;
  assign po08 = ~n325 | ~n327;
  assign n329 = pi18 & n197;
  assign n330 = n200 & n329;
  assign n331 = ~n192 & n330;
  assign n332 = pi26 & n205;
  assign n333 = pi29 & n197;
  assign n334 = ~n200 & n333;
  assign n335 = ~n192 & n334;
  assign n336 = pi33 & ~n197;
  assign n337 = ~n200 & n336;
  assign n338 = ~n192 & n337;
  assign n339 = ~n335 & ~n338;
  assign n340 = ~n192 & ~n331;
  assign n341 = ~n332 & n340;
  assign po09 = ~n339 | ~n341;
  assign n343 = pi19 & n197;
  assign n344 = n200 & n343;
  assign n345 = ~n192 & n344;
  assign n346 = pi27 & n205;
  assign n347 = pi30 & n197;
  assign n348 = ~n200 & n347;
  assign n349 = ~n192 & n348;
  assign n350 = pi34 & ~n197;
  assign n351 = ~n200 & n350;
  assign n352 = ~n192 & n351;
  assign n353 = ~n349 & ~n352;
  assign n354 = ~n192 & ~n345;
  assign n355 = ~n346 & n354;
  assign po10 = ~n353 | ~n355;
  assign n357 = n200 & n207;
  assign n358 = ~n192 & n357;
  assign n359 = pi28 & n205;
  assign n360 = pi31 & n197;
  assign n361 = ~n200 & n360;
  assign n362 = ~n192 & n361;
  assign n363 = pi35 & ~n197;
  assign n364 = ~n200 & n363;
  assign n365 = ~n192 & n364;
  assign n366 = ~n362 & ~n365;
  assign n367 = ~n192 & ~n358;
  assign n368 = ~n359 & n367;
  assign po11 = ~n366 | ~n368;
  assign n370 = n200 & n221;
  assign n371 = ~n192 & n370;
  assign n372 = pi29 & n205;
  assign n373 = pi32 & n197;
  assign n374 = ~n200 & n373;
  assign n375 = ~n192 & n374;
  assign n376 = pi36 & ~n197;
  assign n377 = ~n200 & n376;
  assign n378 = ~n192 & n377;
  assign n379 = ~n375 & ~n378;
  assign n380 = ~n192 & ~n371;
  assign n381 = ~n372 & n380;
  assign po12 = ~n379 | ~n381;
  assign n383 = n200 & n235;
  assign n384 = ~n192 & n383;
  assign n385 = pi30 & n205;
  assign n386 = pi33 & n197;
  assign n387 = ~n200 & n386;
  assign n388 = ~n192 & n387;
  assign n389 = pi37 & ~n197;
  assign n390 = ~n200 & n389;
  assign n391 = ~n192 & n390;
  assign n392 = ~n388 & ~n391;
  assign n393 = ~n192 & ~n384;
  assign n394 = ~n385 & n393;
  assign po13 = ~n392 | ~n394;
  assign n396 = n200 & n249;
  assign n397 = ~n192 & n396;
  assign n398 = pi31 & n205;
  assign n399 = pi34 & n197;
  assign n400 = ~n200 & n399;
  assign n401 = ~n192 & n400;
  assign n402 = pi38 & ~n197;
  assign n403 = ~n200 & n402;
  assign n404 = ~n192 & n403;
  assign n405 = ~n401 & ~n404;
  assign n406 = ~n192 & ~n397;
  assign n407 = ~n398 & n406;
  assign po14 = ~n405 | ~n407;
  assign n409 = n200 & n263;
  assign n410 = ~n192 & n409;
  assign n411 = pi32 & n205;
  assign n412 = pi35 & n197;
  assign n413 = ~n200 & n412;
  assign n414 = ~n192 & n413;
  assign n415 = pi39 & ~n197;
  assign n416 = ~n200 & n415;
  assign n417 = ~n192 & n416;
  assign n418 = ~n414 & ~n417;
  assign n419 = ~n192 & ~n410;
  assign n420 = ~n411 & n419;
  assign po15 = ~n418 | ~n420;
  assign n422 = n200 & n277;
  assign n423 = ~n192 & n422;
  assign n424 = pi33 & n205;
  assign n425 = pi36 & n197;
  assign n426 = ~n200 & n425;
  assign n427 = ~n192 & n426;
  assign n428 = pi52 & ~n197;
  assign n429 = ~n200 & n428;
  assign n430 = ~n192 & n429;
  assign n431 = ~n427 & ~n430;
  assign n432 = ~n192 & ~n423;
  assign n433 = ~n424 & n432;
  assign po16 = ~n431 | ~n433;
  assign n435 = n200 & n291;
  assign n436 = ~n192 & n435;
  assign n437 = pi34 & n205;
  assign n438 = pi37 & n197;
  assign n439 = ~n200 & n438;
  assign n440 = ~n192 & n439;
  assign n441 = pi53 & ~n197;
  assign n442 = ~n200 & n441;
  assign n443 = ~n192 & n442;
  assign n444 = ~n440 & ~n443;
  assign n445 = ~n192 & ~n436;
  assign n446 = ~n437 & n445;
  assign po17 = ~n444 | ~n446;
  assign n448 = n200 & n305;
  assign n449 = ~n192 & n448;
  assign n450 = pi35 & n205;
  assign n451 = pi38 & n197;
  assign n452 = ~n200 & n451;
  assign n453 = ~n192 & n452;
  assign n454 = pi54 & ~n197;
  assign n455 = ~n200 & n454;
  assign n456 = ~n192 & n455;
  assign n457 = ~n453 & ~n456;
  assign n458 = ~n192 & ~n449;
  assign n459 = ~n450 & n458;
  assign po18 = ~n457 | ~n459;
  assign n461 = n200 & n319;
  assign n462 = ~n192 & n461;
  assign n463 = pi36 & n205;
  assign n464 = pi39 & n197;
  assign n465 = ~n200 & n464;
  assign n466 = ~n192 & n465;
  assign n467 = pi55 & ~n197;
  assign n468 = ~n200 & n467;
  assign n469 = ~n192 & n468;
  assign n470 = ~n466 & ~n469;
  assign n471 = ~n192 & ~n462;
  assign n472 = ~n463 & n471;
  assign po19 = ~n470 | ~n472;
  assign n474 = n200 & n333;
  assign n475 = ~n192 & n474;
  assign n476 = pi37 & n205;
  assign n477 = pi41 & n197;
  assign n478 = ~n200 & n477;
  assign n479 = ~n192 & n478;
  assign n480 = pi56 & ~n197;
  assign n481 = ~n200 & n480;
  assign n482 = ~n192 & n481;
  assign n483 = ~n479 & ~n482;
  assign n484 = ~n192 & ~n475;
  assign n485 = ~n476 & n484;
  assign po20 = ~n483 | ~n485;
  assign n487 = n200 & n347;
  assign n488 = ~n192 & n487;
  assign n489 = pi38 & n205;
  assign n490 = pi42 & n197;
  assign n491 = ~n200 & n490;
  assign n492 = ~n192 & n491;
  assign n493 = pi57 & ~n197;
  assign n494 = ~n200 & n493;
  assign n495 = ~n192 & n494;
  assign n496 = ~n492 & ~n495;
  assign n497 = ~n192 & ~n488;
  assign n498 = ~n489 & n497;
  assign po21 = ~n496 | ~n498;
  assign n500 = n200 & n360;
  assign n501 = ~n192 & n500;
  assign n502 = pi39 & n205;
  assign n503 = pi43 & n197;
  assign n504 = ~n200 & n503;
  assign n505 = ~n192 & n504;
  assign n506 = pi58 & ~n197;
  assign n507 = ~n200 & n506;
  assign n508 = ~n192 & n507;
  assign n509 = ~n505 & ~n508;
  assign n510 = ~n192 & ~n501;
  assign n511 = ~n502 & n510;
  assign po22 = ~n509 | ~n511;
  assign n513 = n200 & n373;
  assign n514 = ~n192 & n513;
  assign n515 = pi40 & n205;
  assign n516 = pi44 & n197;
  assign n517 = ~n200 & n516;
  assign n518 = ~n192 & n517;
  assign n519 = pi59 & ~n197;
  assign n520 = ~n200 & n519;
  assign n521 = ~n192 & n520;
  assign n522 = ~n518 & ~n521;
  assign n523 = ~n192 & ~n514;
  assign n524 = ~n515 & n523;
  assign po23 = ~n522 | ~n524;
  assign n526 = n200 & n386;
  assign n527 = ~n192 & n526;
  assign n528 = pi45 & n197;
  assign n529 = ~n200 & n528;
  assign n530 = ~n192 & n529;
  assign n531 = pi60 & ~n197;
  assign n532 = ~n200 & n531;
  assign n533 = ~n192 & n532;
  assign n534 = ~n530 & ~n533;
  assign n535 = ~n192 & ~n527;
  assign n536 = ~n205 & n535;
  assign po24 = ~n534 | ~n536;
  assign n538 = n200 & n399;
  assign n539 = ~n192 & n538;
  assign n540 = pi46 & n197;
  assign n541 = ~n200 & n540;
  assign n542 = ~n192 & n541;
  assign n543 = pi61 & ~n197;
  assign n544 = ~n200 & n543;
  assign n545 = ~n192 & n544;
  assign n546 = ~n542 & ~n545;
  assign n547 = ~n192 & ~n539;
  assign n548 = ~n205 & n547;
  assign po25 = ~n546 | ~n548;
  assign n550 = n200 & n412;
  assign n551 = ~n192 & n550;
  assign n552 = pi47 & n197;
  assign n553 = ~n200 & n552;
  assign n554 = ~n192 & n553;
  assign n555 = pi62 & ~n197;
  assign n556 = ~n200 & n555;
  assign n557 = ~n192 & n556;
  assign n558 = ~n554 & ~n557;
  assign n559 = ~n192 & ~n551;
  assign n560 = ~n205 & n559;
  assign po26 = ~n558 | ~n560;
  assign n562 = n200 & n425;
  assign n563 = ~n192 & n562;
  assign n564 = pi48 & n197;
  assign n565 = ~n200 & n564;
  assign n566 = ~n192 & n565;
  assign n567 = pi63 & ~n197;
  assign n568 = ~n200 & n567;
  assign n569 = ~n192 & n568;
  assign n570 = ~n566 & ~n569;
  assign n571 = ~n192 & ~n563;
  assign n572 = ~n205 & n571;
  assign po27 = ~n570 | ~n572;
  assign n574 = n200 & n438;
  assign n575 = ~n192 & n574;
  assign n576 = pi49 & n197;
  assign n577 = ~n200 & n576;
  assign n578 = ~n192 & n577;
  assign n579 = pi64 & ~n197;
  assign n580 = ~n200 & n579;
  assign n581 = ~n192 & n580;
  assign n582 = ~n578 & ~n581;
  assign n583 = ~n192 & ~n575;
  assign n584 = ~n205 & n583;
  assign po28 = ~n582 | ~n584;
  assign n586 = n200 & n451;
  assign n587 = ~n192 & n586;
  assign n588 = pi50 & n197;
  assign n589 = ~n200 & n588;
  assign n590 = ~n192 & n589;
  assign n591 = pi65 & ~n197;
  assign n592 = ~n200 & n591;
  assign n593 = ~n192 & n592;
  assign n594 = ~n590 & ~n593;
  assign n595 = ~n192 & ~n587;
  assign n596 = ~n205 & n595;
  assign po29 = ~n594 | ~n596;
  assign n598 = n200 & n464;
  assign n599 = ~n192 & n598;
  assign n600 = pi51 & n197;
  assign n601 = ~n200 & n600;
  assign n602 = ~n192 & n601;
  assign n603 = pi66 & ~n197;
  assign n604 = ~n200 & n603;
  assign n605 = ~n192 & n604;
  assign n606 = ~n602 & ~n605;
  assign n607 = ~n192 & ~n599;
  assign n608 = ~n205 & n607;
  assign po30 = ~n606 | ~n608;
  assign n610 = n192 & n200;
  assign n611 = n197 & n610;
  assign n612 = ~n197 & n610;
  assign n613 = n192 & ~n200;
  assign n614 = n197 & n613;
  assign n615 = ~n197 & n613;
  assign n616 = pi83 & n197;
  assign n617 = n200 & n616;
  assign n618 = ~n192 & n617;
  assign n619 = pi45 & ~n197;
  assign n620 = n200 & n619;
  assign n621 = ~n192 & n620;
  assign n622 = pi87 & ~n197;
  assign n623 = ~n200 & n622;
  assign n624 = ~n192 & n623;
  assign n625 = ~n614 & ~n615;
  assign n626 = ~n611 & ~n612;
  assign n627 = n625 & n626;
  assign n628 = ~n618 & ~n621;
  assign n629 = ~n566 & ~n624;
  assign n630 = n628 & n629;
  assign po31 = ~n627 | ~n630;
  assign n632 = pi84 & n197;
  assign n633 = n200 & n632;
  assign n634 = ~n192 & n633;
  assign n635 = pi46 & ~n197;
  assign n636 = n200 & n635;
  assign n637 = ~n192 & n636;
  assign n638 = pi09 & ~n197;
  assign n639 = ~n200 & n638;
  assign n640 = ~n192 & n639;
  assign n641 = ~n634 & ~n637;
  assign n642 = ~n578 & ~n640;
  assign n643 = n641 & n642;
  assign po32 = ~n627 | ~n643;
  assign n645 = pi85 & n197;
  assign n646 = n200 & n645;
  assign n647 = ~n192 & n646;
  assign n648 = pi47 & ~n197;
  assign n649 = n200 & n648;
  assign n650 = ~n192 & n649;
  assign n651 = pi10 & ~n197;
  assign n652 = ~n200 & n651;
  assign n653 = ~n192 & n652;
  assign n654 = ~n647 & ~n650;
  assign n655 = ~n590 & ~n653;
  assign n656 = n654 & n655;
  assign po33 = ~n627 | ~n656;
  assign n658 = pi86 & n197;
  assign n659 = n200 & n658;
  assign n660 = ~n192 & n659;
  assign n661 = pi48 & ~n197;
  assign n662 = n200 & n661;
  assign n663 = ~n192 & n662;
  assign n664 = pi11 & ~n197;
  assign n665 = ~n200 & n664;
  assign n666 = ~n192 & n665;
  assign n667 = ~n660 & ~n663;
  assign n668 = ~n602 & ~n666;
  assign n669 = n667 & n668;
  assign po34 = ~n627 | ~n669;
  assign n671 = n200 & n477;
  assign n672 = ~n192 & n671;
  assign n673 = pi49 & ~n197;
  assign n674 = n200 & n673;
  assign n675 = ~n192 & n674;
  assign n676 = pi87 & n197;
  assign n677 = ~n200 & n676;
  assign n678 = ~n192 & n677;
  assign n679 = pi12 & ~n197;
  assign n680 = ~n200 & n679;
  assign n681 = ~n192 & n680;
  assign n682 = ~n672 & ~n675;
  assign n683 = ~n678 & ~n681;
  assign n684 = n682 & n683;
  assign po35 = ~n627 | ~n684;
  assign n686 = n200 & n490;
  assign n687 = ~n192 & n686;
  assign n688 = pi50 & ~n197;
  assign n689 = n200 & n688;
  assign n690 = ~n192 & n689;
  assign n691 = ~n200 & n201;
  assign n692 = ~n192 & n691;
  assign n693 = pi13 & ~n197;
  assign n694 = ~n200 & n693;
  assign n695 = ~n192 & n694;
  assign n696 = ~n687 & ~n690;
  assign n697 = ~n692 & ~n695;
  assign n698 = n696 & n697;
  assign po36 = ~n627 | ~n698;
  assign n700 = n200 & n503;
  assign n701 = ~n192 & n700;
  assign n702 = pi51 & ~n197;
  assign n703 = n200 & n702;
  assign n704 = ~n192 & n703;
  assign n705 = ~n200 & n217;
  assign n706 = ~n192 & n705;
  assign n707 = pi14 & ~n197;
  assign n708 = ~n200 & n707;
  assign n709 = ~n192 & n708;
  assign n710 = ~n701 & ~n704;
  assign n711 = ~n706 & ~n709;
  assign n712 = n710 & n711;
  assign po37 = ~n627 | ~n712;
  assign n714 = n200 & n516;
  assign n715 = ~n192 & n714;
  assign n716 = n200 & n622;
  assign n717 = ~n192 & n716;
  assign n718 = ~n200 & n231;
  assign n719 = ~n192 & n718;
  assign n720 = pi15 & ~n197;
  assign n721 = ~n200 & n720;
  assign n722 = ~n192 & n721;
  assign n723 = ~n715 & ~n717;
  assign n724 = ~n719 & ~n722;
  assign n725 = n723 & n724;
  assign po38 = ~n627 | ~n725;
  assign n727 = n200 & n528;
  assign n728 = ~n192 & n727;
  assign n729 = n200 & n638;
  assign n730 = ~n192 & n729;
  assign n731 = ~n200 & n245;
  assign n732 = ~n192 & n731;
  assign n733 = pi16 & ~n197;
  assign n734 = ~n200 & n733;
  assign n735 = ~n192 & n734;
  assign n736 = ~n728 & ~n730;
  assign n737 = ~n732 & ~n735;
  assign n738 = n736 & n737;
  assign po39 = ~n627 | ~n738;
  assign n740 = n200 & n540;
  assign n741 = ~n192 & n740;
  assign n742 = n200 & n651;
  assign n743 = ~n192 & n742;
  assign n744 = ~n200 & n259;
  assign n745 = ~n192 & n744;
  assign n746 = pi17 & ~n197;
  assign n747 = ~n200 & n746;
  assign n748 = ~n192 & n747;
  assign n749 = ~n741 & ~n743;
  assign n750 = ~n745 & ~n748;
  assign n751 = n749 & n750;
  assign po40 = ~n627 | ~n751;
  assign n753 = n200 & n552;
  assign n754 = ~n192 & n753;
  assign n755 = n200 & n664;
  assign n756 = ~n192 & n755;
  assign n757 = ~n200 & n273;
  assign n758 = ~n192 & n757;
  assign n759 = pi18 & ~n197;
  assign n760 = ~n200 & n759;
  assign n761 = ~n192 & n760;
  assign n762 = ~n754 & ~n756;
  assign n763 = ~n758 & ~n761;
  assign n764 = n762 & n763;
  assign po41 = ~n627 | ~n764;
  assign n766 = n200 & n564;
  assign n767 = ~n192 & n766;
  assign n768 = n200 & n679;
  assign n769 = ~n192 & n768;
  assign n770 = ~n200 & n287;
  assign n771 = ~n192 & n770;
  assign n772 = pi19 & ~n197;
  assign n773 = ~n200 & n772;
  assign n774 = ~n192 & n773;
  assign n775 = ~n767 & ~n769;
  assign n776 = ~n771 & ~n774;
  assign n777 = n775 & n776;
  assign po42 = ~n627 | ~n777;
  assign n779 = n200 & n576;
  assign n780 = ~n192 & n779;
  assign n781 = n200 & n693;
  assign n782 = ~n192 & n781;
  assign n783 = ~n200 & n301;
  assign n784 = ~n192 & n783;
  assign n785 = pi20 & ~n197;
  assign n786 = ~n200 & n785;
  assign n787 = ~n192 & n786;
  assign n788 = ~n780 & ~n782;
  assign n789 = ~n784 & ~n787;
  assign n790 = n788 & n789;
  assign po43 = ~n627 | ~n790;
  assign n792 = n200 & n588;
  assign n793 = ~n192 & n792;
  assign n794 = n200 & n707;
  assign n795 = ~n192 & n794;
  assign n796 = ~n200 & n315;
  assign n797 = ~n192 & n796;
  assign n798 = pi21 & ~n197;
  assign n799 = ~n200 & n798;
  assign n800 = ~n192 & n799;
  assign n801 = ~n793 & ~n795;
  assign n802 = ~n797 & ~n800;
  assign n803 = n801 & n802;
  assign po44 = ~n627 | ~n803;
  assign n805 = n200 & n600;
  assign n806 = ~n192 & n805;
  assign n807 = n200 & n720;
  assign n808 = ~n192 & n807;
  assign n809 = ~n200 & n329;
  assign n810 = ~n192 & n809;
  assign n811 = pi22 & ~n197;
  assign n812 = ~n200 & n811;
  assign n813 = ~n192 & n812;
  assign n814 = ~n806 & ~n808;
  assign n815 = ~n810 & ~n813;
  assign n816 = n814 & n815;
  assign po45 = ~n627 | ~n816;
  assign n818 = n200 & n676;
  assign n819 = ~n192 & n818;
  assign n820 = n200 & n733;
  assign n821 = ~n192 & n820;
  assign n822 = ~n200 & n343;
  assign n823 = ~n192 & n822;
  assign n824 = pi23 & ~n197;
  assign n825 = ~n200 & n824;
  assign n826 = ~n192 & n825;
  assign n827 = ~n819 & ~n821;
  assign n828 = ~n823 & ~n826;
  assign n829 = n827 & n828;
  assign po46 = ~n627 | ~n829;
  assign n831 = pi67 & n197;
  assign n832 = n200 & n831;
  assign n833 = ~n192 & n832;
  assign n834 = pi75 & ~n197;
  assign n835 = n200 & n834;
  assign n836 = ~n192 & n835;
  assign n837 = pi78 & n197;
  assign n838 = ~n200 & n837;
  assign n839 = ~n192 & n838;
  assign n840 = pi82 & ~n197;
  assign n841 = ~n200 & n840;
  assign n842 = ~n192 & n841;
  assign n843 = ~n833 & ~n836;
  assign n844 = ~n839 & ~n842;
  assign n845 = n843 & n844;
  assign po47 = ~n627 | ~n845;
  assign n847 = pi68 & n197;
  assign n848 = n200 & n847;
  assign n849 = ~n192 & n848;
  assign n850 = pi76 & ~n197;
  assign n851 = n200 & n850;
  assign n852 = ~n192 & n851;
  assign n853 = pi79 & n197;
  assign n854 = ~n200 & n853;
  assign n855 = ~n192 & n854;
  assign n856 = pi83 & ~n197;
  assign n857 = ~n200 & n856;
  assign n858 = ~n192 & n857;
  assign n859 = ~n849 & ~n852;
  assign n860 = ~n855 & ~n858;
  assign n861 = n859 & n860;
  assign po48 = ~n627 | ~n861;
  assign n863 = pi69 & n197;
  assign n864 = n200 & n863;
  assign n865 = ~n192 & n864;
  assign n866 = pi77 & ~n197;
  assign n867 = n200 & n866;
  assign n868 = ~n192 & n867;
  assign n869 = pi80 & n197;
  assign n870 = ~n200 & n869;
  assign n871 = ~n192 & n870;
  assign n872 = pi84 & ~n197;
  assign n873 = ~n200 & n872;
  assign n874 = ~n192 & n873;
  assign n875 = ~n865 & ~n868;
  assign n876 = ~n871 & ~n874;
  assign n877 = n875 & n876;
  assign po49 = ~n627 | ~n877;
  assign n879 = pi70 & n197;
  assign n880 = n200 & n879;
  assign n881 = ~n192 & n880;
  assign n882 = pi78 & ~n197;
  assign n883 = n200 & n882;
  assign n884 = ~n192 & n883;
  assign n885 = pi81 & n197;
  assign n886 = ~n200 & n885;
  assign n887 = ~n192 & n886;
  assign n888 = pi85 & ~n197;
  assign n889 = ~n200 & n888;
  assign n890 = ~n192 & n889;
  assign n891 = ~n881 & ~n884;
  assign n892 = ~n887 & ~n890;
  assign n893 = n891 & n892;
  assign po50 = ~n627 | ~n893;
  assign n895 = pi71 & n197;
  assign n896 = n200 & n895;
  assign n897 = ~n192 & n896;
  assign n898 = pi79 & ~n197;
  assign n899 = n200 & n898;
  assign n900 = ~n192 & n899;
  assign n901 = pi82 & n197;
  assign n902 = ~n200 & n901;
  assign n903 = ~n192 & n902;
  assign n904 = pi86 & ~n197;
  assign n905 = ~n200 & n904;
  assign n906 = ~n192 & n905;
  assign n907 = ~n897 & ~n900;
  assign n908 = ~n903 & ~n906;
  assign n909 = n907 & n908;
  assign po51 = ~n627 | ~n909;
  assign n911 = pi72 & n197;
  assign n912 = n200 & n911;
  assign n913 = ~n192 & n912;
  assign n914 = pi80 & ~n197;
  assign n915 = n200 & n914;
  assign n916 = ~n192 & n915;
  assign n917 = ~n200 & n616;
  assign n918 = ~n192 & n917;
  assign n919 = pi41 & ~n197;
  assign n920 = ~n200 & n919;
  assign n921 = ~n192 & n920;
  assign n922 = ~n913 & ~n916;
  assign n923 = ~n918 & ~n921;
  assign n924 = n922 & n923;
  assign po52 = ~n627 | ~n924;
  assign n926 = pi73 & n197;
  assign n927 = n200 & n926;
  assign n928 = ~n192 & n927;
  assign n929 = pi81 & ~n197;
  assign n930 = n200 & n929;
  assign n931 = ~n192 & n930;
  assign n932 = ~n200 & n632;
  assign n933 = ~n192 & n932;
  assign n934 = pi42 & ~n197;
  assign n935 = ~n200 & n934;
  assign n936 = ~n192 & n935;
  assign n937 = ~n928 & ~n931;
  assign n938 = ~n933 & ~n936;
  assign n939 = n937 & n938;
  assign po53 = ~n627 | ~n939;
  assign n941 = pi74 & n197;
  assign n942 = n200 & n941;
  assign n943 = ~n192 & n942;
  assign n944 = n200 & n840;
  assign n945 = ~n192 & n944;
  assign n946 = ~n200 & n645;
  assign n947 = ~n192 & n946;
  assign n948 = pi43 & ~n197;
  assign n949 = ~n200 & n948;
  assign n950 = ~n192 & n949;
  assign n951 = ~n943 & ~n945;
  assign n952 = ~n947 & ~n950;
  assign n953 = n951 & n952;
  assign po54 = ~n627 | ~n953;
  assign n955 = pi75 & n197;
  assign n956 = n200 & n955;
  assign n957 = ~n192 & n956;
  assign n958 = n200 & n856;
  assign n959 = ~n192 & n958;
  assign n960 = ~n200 & n658;
  assign n961 = ~n192 & n960;
  assign n962 = pi44 & ~n197;
  assign n963 = ~n200 & n962;
  assign n964 = ~n192 & n963;
  assign n965 = ~n957 & ~n959;
  assign n966 = ~n961 & ~n964;
  assign n967 = n965 & n966;
  assign po55 = ~n627 | ~n967;
  assign n969 = pi76 & n197;
  assign n970 = n200 & n969;
  assign n971 = ~n192 & n970;
  assign n972 = n200 & n872;
  assign n973 = ~n192 & n972;
  assign n974 = ~n200 & n619;
  assign n975 = ~n192 & n974;
  assign n976 = ~n971 & ~n973;
  assign n977 = ~n479 & ~n975;
  assign n978 = n976 & n977;
  assign po56 = ~n627 | ~n978;
  assign n980 = pi77 & n197;
  assign n981 = n200 & n980;
  assign n982 = ~n192 & n981;
  assign n983 = n200 & n888;
  assign n984 = ~n192 & n983;
  assign n985 = ~n200 & n635;
  assign n986 = ~n192 & n985;
  assign n987 = ~n982 & ~n984;
  assign n988 = ~n492 & ~n986;
  assign n989 = n987 & n988;
  assign po57 = ~n627 | ~n989;
  assign n991 = n200 & n837;
  assign n992 = ~n192 & n991;
  assign n993 = n200 & n904;
  assign n994 = ~n192 & n993;
  assign n995 = ~n200 & n648;
  assign n996 = ~n192 & n995;
  assign n997 = ~n992 & ~n994;
  assign n998 = ~n505 & ~n996;
  assign n999 = n997 & n998;
  assign po58 = ~n627 | ~n999;
  assign n1001 = n200 & n853;
  assign n1002 = ~n192 & n1001;
  assign n1003 = n200 & n919;
  assign n1004 = ~n192 & n1003;
  assign n1005 = ~n200 & n661;
  assign n1006 = ~n192 & n1005;
  assign n1007 = ~n1002 & ~n1004;
  assign n1008 = ~n518 & ~n1006;
  assign n1009 = n1007 & n1008;
  assign po59 = ~n627 | ~n1009;
  assign n1011 = n200 & n869;
  assign n1012 = ~n192 & n1011;
  assign n1013 = n200 & n934;
  assign n1014 = ~n192 & n1013;
  assign n1015 = ~n200 & n673;
  assign n1016 = ~n192 & n1015;
  assign n1017 = ~n1012 & ~n1014;
  assign n1018 = ~n530 & ~n1016;
  assign n1019 = n1017 & n1018;
  assign po60 = ~n627 | ~n1019;
  assign n1021 = n200 & n885;
  assign n1022 = ~n192 & n1021;
  assign n1023 = n200 & n948;
  assign n1024 = ~n192 & n1023;
  assign n1025 = ~n200 & n688;
  assign n1026 = ~n192 & n1025;
  assign n1027 = ~n1022 & ~n1024;
  assign n1028 = ~n542 & ~n1026;
  assign n1029 = n1027 & n1028;
  assign po61 = ~n627 | ~n1029;
  assign n1031 = n200 & n901;
  assign n1032 = ~n192 & n1031;
  assign n1033 = n200 & n962;
  assign n1034 = ~n192 & n1033;
  assign n1035 = ~n200 & n702;
  assign n1036 = ~n192 & n1035;
  assign n1037 = ~n1032 & ~n1034;
  assign n1038 = ~n554 & ~n1036;
  assign n1039 = n1037 & n1038;
  assign po62 = ~n627 | ~n1039;
endmodule



module i2c_best_speed (
        pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, 
        po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107;
assign w0 = pi012 & ~pi013;
assign w1 = ~pi012 & pi013;
assign w2 = ~w0 & ~w1;
assign w3 = ~pi009 & ~w2;
assign w4 = ~pi012 & ~pi013;
assign w5 = ~pi007 & pi009;
assign w6 = w4 & w5;
assign w7 = (~pi007 & w3) | (~pi007 & w6) | (w3 & w6);
assign w8 = ~pi009 & w4;
assign w9 = pi006 & ~pi007;
assign w10 = pi006 & ~w9;
assign w11 = (pi006 & ~w8) | (pi006 & w10) | (~w8 & w10);
assign w12 = w8 & w9;
assign w13 = pi007 & ~pi009;
assign w14 = w4 & w13;
assign w15 = ~pi006 & w14;
assign w16 = ~w12 & ~w15;
assign w17 = (~w7 & w11) | (~w7 & w16) | (w11 & w16);
assign w18 = ~pi005 & ~pi011;
assign w19 = ~pi016 & ~pi018;
assign w20 = w18 & w19;
assign w21 = ~pi019 & ~pi022;
assign w22 = w20 & w21;
assign w23 = ~pi008 & ~pi010;
assign w24 = ~pi014 & ~pi021;
assign w25 = w23 & w24;
assign w26 = ~pi017 & w25;
assign w27 = ~pi004 & ~pi007;
assign w28 = ~pi009 & ~pi012;
assign w29 = w27 & w28;
assign w30 = ~pi013 & w29;
assign w31 = w26 & w30;
assign w32 = w22 & w31;
assign w33 = w17 & w32;
assign w34 = ~pi000 & ~pi054;
assign w35 = (~pi000 & w33) | (~pi000 & w34) | (w33 & w34);
assign w36 = pi007 & pi013;
assign w37 = (pi007 & ~w25) | (pi007 & w36) | (~w25 & w36);
assign w38 = ~pi004 & ~pi005;
assign w39 = ~pi006 & ~pi012;
assign w40 = w38 & w39;
assign w41 = ~pi022 & w40;
assign w42 = ~w37 & w41;
assign w43 = ~pi011 & ~pi016;
assign w44 = ~pi017 & ~pi018;
assign w45 = w43 & w44;
assign w46 = ~pi019 & pi054;
assign w47 = ~pi009 & w46;
assign w48 = w45 & w47;
assign w49 = w42 & w48;
assign w50 = pi014 & ~pi021;
assign w51 = ~pi014 & pi021;
assign w52 = ~w50 & ~w51;
assign w53 = ~pi010 & ~w52;
assign w54 = ~pi007 & ~pi010;
assign w55 = w24 & ~w54;
assign w56 = ~pi013 & w55;
assign w57 = (~pi013 & w53) | (~pi013 & w56) | (w53 & w56);
assign w58 = pi008 & ~pi010;
assign w59 = w24 & w58;
assign w60 = pi008 & pi013;
assign w61 = (pi008 & ~w59) | (pi008 & w60) | (~w59 & w60);
assign w62 = ~pi013 & w59;
assign w63 = ~pi010 & pi013;
assign w64 = w24 & w63;
assign w65 = ~pi008 & w64;
assign w66 = ~w62 & ~w65;
assign w67 = (~w57 & w61) | (~w57 & w66) | (w61 & w66);
assign w68 = w49 & ~w67;
assign w69 = ~pi005 & ~pi022;
assign w70 = ~pi009 & ~pi011;
assign w71 = ~w69 & w70;
assign w72 = w69 & ~w70;
assign w73 = ~w71 & ~w72;
assign w74 = pi054 & ~pi056;
assign w75 = ~w73 & w74;
assign w76 = ~w68 & ~w75;
assign w77 = ~w35 & w76;
assign w78 = ~pi003 & ~pi129;
assign w79 = ~w77 & w78;
assign w80 = w22 & w25;
assign w81 = w30 & w80;
assign w82 = w17 & w81;
assign w83 = ~pi001 & w78;
assign w84 = ~pi017 & pi054;
assign w85 = w78 & ~w84;
assign w86 = ~pi001 & w85;
assign w87 = (w82 & w83) | (w82 & w86) | (w83 & w86);
assign w88 = ~pi005 & ~w17;
assign w89 = pi005 & ~pi013;
assign w90 = w29 & w89;
assign w91 = w17 & w90;
assign w92 = ~w88 & ~w91;
assign w93 = w45 & w46;
assign w94 = ~pi003 & ~pi004;
assign w95 = ~pi022 & ~pi129;
assign w96 = w94 & w95;
assign w97 = w25 & w96;
assign w98 = w93 & w97;
assign w99 = ~w92 & w98;
assign w100 = ~w87 & ~w99;
assign w101 = ~pi002 & ~pi015;
assign w102 = ~pi020 & ~pi024;
assign w103 = w101 & w102;
assign w104 = ~pi045 & ~pi049;
assign w105 = w103 & w104;
assign w106 = ~pi043 & ~pi047;
assign w107 = ~pi048 & w106;
assign w108 = w105 & w107;
assign w109 = ~pi038 & ~pi040;
assign w110 = ~pi042 & ~pi044;
assign w111 = w109 & w110;
assign w112 = ~pi046 & ~pi050;
assign w113 = ~pi041 & w112;
assign w114 = w111 & w113;
assign w115 = pi082 & ~w114;
assign w116 = (pi082 & ~w108) | (pi082 & w115) | (~w108 & w115);
assign w117 = pi122 & pi127;
assign w118 = ~pi065 & ~w117;
assign w119 = ~w116 & w118;
assign w120 = ~w116 & w117;
assign w121 = w111 & w112;
assign w122 = ~pi024 & ~pi043;
assign w123 = ~pi045 & ~pi047;
assign w124 = w122 & w123;
assign w125 = ~pi048 & ~pi049;
assign w126 = w124 & w125;
assign w127 = w121 & w126;
assign w128 = ~pi015 & ~pi020;
assign w129 = ~pi041 & pi082;
assign w130 = w128 & w129;
assign w131 = w127 & w130;
assign w132 = w116 & ~w131;
assign w133 = ~w120 & ~w132;
assign w134 = ~pi002 & pi065;
assign w135 = (~pi002 & w117) | (~pi002 & w134) | (w117 & w134);
assign w136 = (~pi002 & w116) | (~pi002 & w135) | (w116 & w135);
assign w137 = (~w119 & w133) | (~w119 & w136) | (w133 & w136);
assign w138 = ~pi129 & ~w137;
assign w139 = pi000 & ~pi113;
assign w140 = ~pi123 & w139;
assign w141 = w25 & w30;
assign w142 = ~pi017 & w21;
assign w143 = w20 & w142;
assign w144 = w141 & w143;
assign w145 = w17 & w144;
assign w146 = ~pi061 & ~pi118;
assign w147 = ~w140 & ~w146;
assign w148 = (~w140 & w145) | (~w140 & w147) | (w145 & w147);
assign w149 = ~pi129 & ~w148;
assign w150 = pi004 & ~pi054;
assign w151 = w41 & w93;
assign w152 = ~pi007 & ~pi009;
assign w153 = ~pi013 & w152;
assign w154 = ~pi008 & pi010;
assign w155 = w24 & w154;
assign w156 = w153 & w155;
assign w157 = ~w150 & ~w156;
assign w158 = (~w150 & ~w151) | (~w150 & w157) | (~w151 & w157);
assign w159 = w78 & ~w158;
assign w160 = ~pi016 & ~pi017;
assign w161 = w18 & w160;
assign w162 = ~pi022 & pi054;
assign w163 = w78 & w162;
assign w164 = w161 & w163;
assign w165 = ~pi018 & ~pi019;
assign w166 = ~pi029 & w165;
assign w167 = ~pi059 & w166;
assign w168 = w164 & w167;
assign w169 = w141 & w168;
assign w170 = w17 & w169;
assign w171 = ~pi025 & pi028;
assign w172 = w170 & w171;
assign w173 = pi005 & ~pi054;
assign w174 = w78 & w173;
assign w175 = ~w172 & ~w174;
assign w176 = pi025 & ~pi028;
assign w177 = w170 & w176;
assign w178 = ~pi054 & w78;
assign w179 = pi006 & w178;
assign w180 = ~w177 & ~w179;
assign w181 = w151 & w153;
assign w182 = w59 & w181;
assign w183 = pi007 & ~pi054;
assign w184 = ~w182 & ~w183;
assign w185 = w78 & ~w184;
assign w186 = pi008 & ~pi054;
assign w187 = ~pi007 & ~pi013;
assign w188 = w23 & w187;
assign w189 = ~pi009 & w188;
assign w190 = w151 & w189;
assign w191 = ~w51 & ~w186;
assign w192 = (~w186 & ~w190) | (~w186 & w191) | (~w190 & w191);
assign w193 = w78 & ~w192;
assign w194 = pi009 & ~pi054;
assign w195 = ~pi005 & ~pi017;
assign w196 = w165 & w195;
assign w197 = w162 & w196;
assign w198 = w141 & w197;
assign w199 = w17 & w198;
assign w200 = pi011 & ~pi016;
assign w201 = ~w194 & ~w200;
assign w202 = (~w194 & ~w199) | (~w194 & w201) | (~w199 & w201);
assign w203 = w78 & ~w202;
assign w204 = pi010 & ~pi054;
assign w205 = ~pi021 & w189;
assign w206 = w151 & w205;
assign w207 = ~pi014 & ~w204;
assign w208 = (~w204 & ~w206) | (~w204 & w207) | (~w206 & w207);
assign w209 = w78 & ~w208;
assign w210 = ~pi005 & w46;
assign w211 = w45 & w210;
assign w212 = pi022 & w211;
assign w213 = w141 & w212;
assign w214 = w17 & w213;
assign w215 = pi011 & ~pi054;
assign w216 = ~w214 & ~w215;
assign w217 = w78 & ~w216;
assign w218 = pi012 & ~pi054;
assign w219 = w161 & w162;
assign w220 = w141 & w219;
assign w221 = w17 & w220;
assign w222 = pi018 & ~pi019;
assign w223 = ~w218 & ~w222;
assign w224 = (~w218 & ~w221) | (~w218 & w223) | (~w221 & w223);
assign w225 = w78 & ~w224;
assign w226 = pi013 & ~pi054;
assign w227 = ~pi025 & ~pi028;
assign w228 = pi029 & pi054;
assign w229 = w227 & w228;
assign w230 = ~pi059 & w229;
assign w231 = ~w226 & ~w230;
assign w232 = (~w145 & ~w226) | (~w145 & w231) | (~w226 & w231);
assign w233 = w78 & ~w232;
assign w234 = (~pi008 & w57) | (~pi008 & w65) | (w57 & w65);
assign w235 = pi013 & w48;
assign w236 = w42 & w235;
assign w237 = w234 & w236;
assign w238 = pi014 & ~pi054;
assign w239 = ~w237 & ~w238;
assign w240 = w78 & ~w239;
assign w241 = ~pi015 & ~pi041;
assign w242 = w127 & w241;
assign w243 = pi015 & pi041;
assign w244 = (pi015 & ~w127) | (pi015 & w243) | (~w127 & w243);
assign w245 = ~w242 & ~w244;
assign w246 = ~pi082 & ~pi129;
assign w247 = (~pi129 & ~w245) | (~pi129 & w246) | (~w245 & w246);
assign w248 = pi070 & ~pi082;
assign w249 = ~w117 & w248;
assign w250 = ~pi020 & pi070;
assign w251 = (~pi020 & w117) | (~pi020 & w250) | (w117 & w250);
assign w252 = ~pi002 & w251;
assign w253 = ~pi082 & w117;
assign w254 = ~pi015 & w253;
assign w255 = (~pi015 & w252) | (~pi015 & w254) | (w252 & w254);
assign w256 = ~w249 & ~w255;
assign w257 = w247 & w256;
assign w258 = pi006 & w98;
assign w259 = ~w92 & w258;
assign w260 = pi016 & ~pi054;
assign w261 = w78 & w260;
assign w262 = ~w259 & ~w261;
assign w263 = pi017 & ~pi054;
assign w264 = ~pi029 & pi059;
assign w265 = w227 & w264;
assign w266 = w84 & w265;
assign w267 = ~w263 & ~w266;
assign w268 = (~w82 & ~w263) | (~w82 & w267) | (~w263 & w267);
assign w269 = w78 & ~w268;
assign w270 = pi018 & ~pi054;
assign w271 = ~pi011 & pi016;
assign w272 = ~w270 & ~w271;
assign w273 = (~w199 & ~w270) | (~w199 & w272) | (~w270 & w272);
assign w274 = w78 & ~w273;
assign w275 = pi019 & ~pi054;
assign w276 = pi017 & pi054;
assign w277 = ~w275 & ~w276;
assign w278 = (~w82 & ~w275) | (~w82 & w277) | (~w275 & w277);
assign w279 = w78 & ~w278;
assign w280 = ~pi020 & w241;
assign w281 = w127 & w280;
assign w282 = pi020 & ~w241;
assign w283 = (pi020 & ~w127) | (pi020 & w282) | (~w127 & w282);
assign w284 = ~w281 & ~w283;
assign w285 = (~pi129 & w246) | (~pi129 & ~w284) | (w246 & ~w284);
assign w286 = pi071 & ~pi082;
assign w287 = ~w117 & w286;
assign w288 = ~pi002 & pi071;
assign w289 = (~pi002 & w117) | (~pi002 & w288) | (w117 & w288);
assign w290 = ~w253 & ~w289;
assign w291 = pi020 & ~w287;
assign w292 = (~w287 & w290) | (~w287 & w291) | (w290 & w291);
assign w293 = w285 & w292;
assign w294 = pi021 & ~pi054;
assign w295 = ~pi018 & pi019;
assign w296 = ~w294 & ~w295;
assign w297 = (~w221 & ~w294) | (~w221 & w296) | (~w294 & w296);
assign w298 = w78 & ~w297;
assign w299 = pi022 & ~pi054;
assign w300 = ~pi022 & w141;
assign w301 = w17 & w300;
assign w302 = pi005 & w46;
assign w303 = w45 & w302;
assign w304 = ~w299 & ~w303;
assign w305 = (~w299 & ~w301) | (~w299 & w304) | (~w301 & w304);
assign w306 = w78 & ~w305;
assign w307 = ~pi023 & pi055;
assign w308 = ~pi129 & ~w307;
assign w309 = pi061 & w308;
assign w310 = ~pi024 & ~pi045;
assign w311 = pi082 & ~w310;
assign w312 = pi082 | w311;
assign w313 = ~pi041 & ~pi048;
assign w314 = w106 & w313;
assign w315 = (pi082 & w311) | (pi082 & ~w314) | (w311 & ~w314);
assign w316 = (~w121 & w312) | (~w121 & w315) | (w312 & w315);
assign w317 = pi082 & ~w104;
assign w318 = (pi082 & ~w103) | (pi082 & w317) | (~w103 & w317);
assign w319 = pi024 & w117;
assign w320 = ~pi063 & ~w117;
assign w321 = ~w319 & ~w320;
assign w322 = ~w318 & w321;
assign w323 = ~w316 & ~w322;
assign w324 = pi045 & ~w322;
assign w325 = pi082 & ~w314;
assign w326 = (pi082 & ~w121) | (pi082 & w325) | (~w121 & w325);
assign w327 = pi024 & w326;
assign w328 = (pi024 & w324) | (pi024 & w327) | (w324 & w327);
assign w329 = ~w323 & ~w328;
assign w330 = ~pi129 & ~w329;
assign w331 = pi058 & ~pi085;
assign w332 = ~pi058 & pi085;
assign w333 = ~w331 & ~w332;
assign w334 = ~pi053 & ~w333;
assign w335 = ~pi058 & ~pi085;
assign w336 = ~pi027 & pi053;
assign w337 = w335 & w336;
assign w338 = (~pi027 & w334) | (~pi027 & w337) | (w334 & w337);
assign w339 = ~pi053 & w335;
assign w340 = pi026 & ~pi027;
assign w341 = pi026 & ~w340;
assign w342 = (pi026 & ~w339) | (pi026 & w341) | (~w339 & w341);
assign w343 = w339 & w340;
assign w344 = pi027 & ~pi053;
assign w345 = w335 & w344;
assign w346 = ~pi026 & w345;
assign w347 = ~w343 & ~w346;
assign w348 = (~w338 & w342) | (~w338 & w347) | (w342 & w347);
assign w349 = ~pi095 & ~pi100;
assign w350 = pi097 & ~pi110;
assign w351 = (~pi110 & ~w349) | (~pi110 & w350) | (~w349 & w350);
assign w352 = ~pi026 & ~pi027;
assign w353 = ~w351 & w352;
assign w354 = pi085 & ~pi116;
assign w355 = w335 & ~w352;
assign w356 = ~pi116 & ~w355;
assign w357 = (~w353 & w354) | (~w353 & w356) | (w354 & w356);
assign w358 = ~w348 & w357;
assign w359 = (~pi085 & w353) | (~pi085 & w355) | (w353 & w355);
assign w360 = ~pi058 & ~pi116;
assign w361 = w352 & w360;
assign w362 = ~pi039 & ~pi051;
assign w363 = ~pi052 & pi116;
assign w364 = w362 & w363;
assign w365 = ~pi026 & ~pi053;
assign w366 = pi026 & pi027;
assign w367 = ~pi053 & ~w366;
assign w368 = (~w364 & w365) | (~w364 & w367) | (w365 & w367);
assign w369 = ~w361 & ~w368;
assign w370 = w359 & ~w369;
assign w371 = w78 & w370;
assign w372 = (w78 & w358) | (w78 & w371) | (w358 & w371);
assign w373 = ~pi025 & ~pi116;
assign w374 = ~pi052 & w362;
assign w375 = pi027 & pi116;
assign w376 = ~w373 & ~w375;
assign w377 = (~w373 & w374) | (~w373 & w376) | (w374 & w376);
assign w378 = pi058 & pi116;
assign w379 = ~pi025 & ~pi027;
assign w380 = (~pi027 & w378) | (~pi027 & w379) | (w378 & w379);
assign w381 = ~pi026 & w380;
assign w382 = w377 & ~w381;
assign w383 = w372 & w382;
assign w384 = ~pi085 & ~pi096;
assign w385 = ~pi110 & w384;
assign w386 = pi085 & pi116;
assign w387 = ~w385 & ~w386;
assign w388 = ~pi003 & ~pi026;
assign w389 = ~pi027 & ~pi053;
assign w390 = w388 & w389;
assign w391 = ~pi058 & ~pi129;
assign w392 = w390 & w391;
assign w393 = ~w387 & w392;
assign w394 = pi100 & w393;
assign w395 = ~w383 & ~w394;
assign w396 = ~pi053 & ~pi058;
assign w397 = ~pi085 & w396;
assign w398 = w340 & w397;
assign w399 = w78 & ~w364;
assign w400 = w398 & w399;
assign w401 = ~w394 & ~w400;
assign w402 = pi027 & ~pi129;
assign w403 = w388 & w402;
assign w404 = w397 & w403;
assign w405 = ~w364 & w404;
assign w406 = ~pi100 & w391;
assign w407 = w390 & w406;
assign w408 = ~pi096 & ~pi110;
assign w409 = ~pi085 & pi095;
assign w410 = w408 & w409;
assign w411 = ~w386 & ~w410;
assign w412 = w407 & ~w411;
assign w413 = ~w405 & ~w412;
assign w414 = ~pi116 & ~w348;
assign w415 = ~w413 & ~w414;
assign w416 = pi028 & ~pi116;
assign w417 = ~w348 & w416;
assign w418 = ~pi026 & pi028;
assign w419 = ~w351 & w418;
assign w420 = pi026 & w364;
assign w421 = ~w419 & ~w420;
assign w422 = ~pi027 & ~pi085;
assign w423 = w396 & w422;
assign w424 = ~w421 & w423;
assign w425 = ~w417 & ~w424;
assign w426 = ~w415 & w425;
assign w427 = w78 & ~w426;
assign w428 = ~pi095 & ~pi096;
assign w429 = pi097 & ~pi100;
assign w430 = w428 & w429;
assign w431 = ~pi053 & pi110;
assign w432 = ~pi058 & w431;
assign w433 = (w396 & ~w430) | (w396 & w432) | (~w430 & w432);
assign w434 = pi053 & pi116;
assign w435 = ~pi085 & ~w434;
assign w436 = ~pi027 & ~pi129;
assign w437 = w388 & w436;
assign w438 = w435 & w437;
assign w439 = ~w433 & w438;
assign w440 = pi097 & pi116;
assign w441 = pi058 & ~w440;
assign w442 = w439 & ~w441;
assign w443 = ~w414 & w442;
assign w444 = ~pi026 & ~pi085;
assign w445 = w396 & w444;
assign w446 = ~pi027 & w445;
assign w447 = pi116 & w351;
assign w448 = (pi116 & ~w446) | (pi116 & w447) | (~w446 & w447);
assign w449 = pi029 & ~w448;
assign w450 = pi029 & ~w351;
assign w451 = w446 & w450;
assign w452 = (~w348 & w449) | (~w348 & w451) | (w449 & w451);
assign w453 = ~w443 & ~w452;
assign w454 = w78 & ~w453;
assign w455 = pi060 & pi109;
assign w456 = pi030 & ~pi109;
assign w457 = ~w455 & ~w456;
assign w458 = ~pi106 & ~w457;
assign w459 = pi088 & pi106;
assign w460 = ~w458 & ~w459;
assign w461 = ~pi129 & ~w460;
assign w462 = pi031 & ~pi109;
assign w463 = pi030 & pi109;
assign w464 = ~w462 & ~w463;
assign w465 = ~pi106 & ~w464;
assign w466 = pi089 & pi106;
assign w467 = ~w465 & ~w466;
assign w468 = ~pi129 & ~w467;
assign w469 = pi032 & ~pi109;
assign w470 = pi031 & pi109;
assign w471 = ~w469 & ~w470;
assign w472 = ~pi106 & ~w471;
assign w473 = pi099 & pi106;
assign w474 = ~w472 & ~w473;
assign w475 = ~pi129 & ~w474;
assign w476 = pi033 & ~pi109;
assign w477 = pi032 & pi109;
assign w478 = ~w476 & ~w477;
assign w479 = ~pi106 & ~w478;
assign w480 = pi090 & pi106;
assign w481 = ~w479 & ~w480;
assign w482 = ~pi129 & ~w481;
assign w483 = pi034 & ~pi109;
assign w484 = pi033 & pi109;
assign w485 = ~w483 & ~w484;
assign w486 = ~pi106 & ~w485;
assign w487 = pi091 & pi106;
assign w488 = ~w486 & ~w487;
assign w489 = ~pi129 & ~w488;
assign w490 = pi035 & ~pi109;
assign w491 = pi034 & pi109;
assign w492 = ~w490 & ~w491;
assign w493 = ~pi106 & ~w492;
assign w494 = pi092 & pi106;
assign w495 = ~w493 & ~w494;
assign w496 = ~pi129 & ~w495;
assign w497 = pi036 & ~pi109;
assign w498 = pi035 & pi109;
assign w499 = ~w497 & ~w498;
assign w500 = ~pi106 & ~w499;
assign w501 = pi098 & pi106;
assign w502 = ~w500 & ~w501;
assign w503 = ~pi129 & ~w502;
assign w504 = pi037 & ~pi109;
assign w505 = pi036 & pi109;
assign w506 = ~w504 & ~w505;
assign w507 = ~pi106 & ~w506;
assign w508 = pi093 & pi106;
assign w509 = ~w507 & ~w508;
assign w510 = ~pi129 & ~w509;
assign w511 = ~pi050 & w104;
assign w512 = w103 & w511;
assign w513 = ~pi041 & ~pi043;
assign w514 = ~pi046 & ~pi047;
assign w515 = w513 & w514;
assign w516 = ~pi038 & ~pi048;
assign w517 = w515 & w516;
assign w518 = w512 & w517;
assign w519 = pi082 & ~w518;
assign w520 = ~pi074 & ~w117;
assign w521 = pi038 & w117;
assign w522 = ~w520 & ~w521;
assign w523 = ~w519 & w522;
assign w524 = ~pi129 & ~w523;
assign w525 = ~pi040 & ~pi042;
assign w526 = ~pi044 & w525;
assign w527 = pi038 & w526;
assign w528 = ~pi038 & ~w526;
assign w529 = ~w527 & ~w528;
assign w530 = pi082 & ~w529;
assign w531 = w524 & ~w530;
assign w532 = ~pi051 & ~pi052;
assign w533 = ~pi039 & pi109;
assign w534 = w532 & w533;
assign w535 = ~pi106 & ~w534;
assign w536 = ~pi052 & pi109;
assign w537 = ~pi051 & w536;
assign w538 = pi039 & ~w537;
assign w539 = w535 & ~w538;
assign w540 = ~pi129 & ~w539;
assign w541 = ~pi073 & ~w117;
assign w542 = w526 & w541;
assign w543 = ~pi082 & ~w541;
assign w544 = w526 & ~w543;
assign w545 = (~w518 & w542) | (~w518 & w544) | (w542 & w544);
assign w546 = ~pi073 & ~pi082;
assign w547 = ~w117 & w546;
assign w548 = pi082 & ~w110;
assign w549 = ~w253 & ~w548;
assign w550 = ~pi040 & ~w547;
assign w551 = (~w547 & w549) | (~w547 & w550) | (w549 & w550);
assign w552 = ~w545 & w551;
assign w553 = ~pi129 & ~w552;
assign w554 = pi041 & w117;
assign w555 = ~pi076 & ~w117;
assign w556 = ~w554 & ~w555;
assign w557 = ~pi048 & w515;
assign w558 = w105 & w557;
assign w559 = pi082 & ~w558;
assign w560 = w556 & ~w559;
assign w561 = pi041 & ~w121;
assign w562 = ~w114 & ~w561;
assign w563 = pi082 & w562;
assign w564 = ~pi129 & ~w563;
assign w565 = ~w560 & w564;
assign w566 = w110 & w116;
assign w567 = pi044 & pi082;
assign w568 = ~w253 & ~w567;
assign w569 = pi042 & ~w568;
assign w570 = ~w117 & ~w548;
assign w571 = ~pi072 & w570;
assign w572 = ~w569 & ~w571;
assign w573 = ~w566 & w572;
assign w574 = ~pi129 & ~w573;
assign w575 = pi077 & ~w117;
assign w576 = ~pi043 & w117;
assign w577 = ~w575 & ~w576;
assign w578 = ~w559 & ~w577;
assign w579 = ~pi129 & ~w578;
assign w580 = pi043 & w114;
assign w581 = ~pi043 & ~w114;
assign w582 = ~w580 & ~w581;
assign w583 = pi082 & ~w582;
assign w584 = w579 & ~w583;
assign w585 = pi044 & w117;
assign w586 = ~w116 & w585;
assign w587 = ~pi044 & w116;
assign w588 = ~w586 & ~w587;
assign w589 = ~pi044 & ~pi067;
assign w590 = ~w117 & w589;
assign w591 = pi044 & ~pi067;
assign w592 = (~pi067 & ~w117) | (~pi067 & w591) | (~w117 & w591);
assign w593 = (~w116 & w590) | (~w116 & w592) | (w590 & w592);
assign w594 = w588 & ~w593;
assign w595 = ~pi129 & ~w594;
assign w596 = ~pi045 & w314;
assign w597 = w121 & w596;
assign w598 = pi045 & ~w314;
assign w599 = (pi045 & ~w121) | (pi045 & w598) | (~w121 & w598);
assign w600 = ~w597 & ~w599;
assign w601 = (~pi129 & w246) | (~pi129 & ~w600) | (w246 & ~w600);
assign w602 = pi068 & ~pi082;
assign w603 = ~w117 & w602;
assign w604 = ~pi068 & ~w117;
assign w605 = ~w253 & w604;
assign w606 = (~w105 & ~w253) | (~w105 & w605) | (~w253 & w605);
assign w607 = pi045 & ~w603;
assign w608 = (~w603 & w606) | (~w603 & w607) | (w606 & w607);
assign w609 = w601 & w608;
assign w610 = pi046 & w117;
assign w611 = ~pi075 & ~w117;
assign w612 = ~w610 & ~w611;
assign w613 = ~w116 & w612;
assign w614 = ~pi038 & ~pi050;
assign w615 = ~pi046 & w526;
assign w616 = w614 & w615;
assign w617 = pi082 & ~w616;
assign w618 = ~pi050 & w526;
assign w619 = ~pi038 & w618;
assign w620 = pi046 & ~w619;
assign w621 = w617 & ~w620;
assign w622 = ~pi129 & ~w621;
assign w623 = ~w613 & w622;
assign w624 = pi082 & ~w106;
assign w625 = (pi082 & ~w114) | (pi082 & w624) | (~w114 & w624);
assign w626 = pi043 & pi047;
assign w627 = (pi047 & ~w114) | (pi047 & w626) | (~w114 & w626);
assign w628 = w625 & ~w627;
assign w629 = ~pi129 & ~w628;
assign w630 = pi064 & ~pi082;
assign w631 = ~w117 & w630;
assign w632 = ~pi064 & ~w117;
assign w633 = w557 & ~w632;
assign w634 = ~w105 & ~w253;
assign w635 = (~w253 & ~w633) | (~w253 & w634) | (~w633 & w634);
assign w636 = pi047 & ~w631;
assign w637 = (~w631 & w635) | (~w631 & w636) | (w635 & w636);
assign w638 = w629 & w637;
assign w639 = ~pi048 & w114;
assign w640 = w106 & w639;
assign w641 = pi082 & ~w640;
assign w642 = w106 & w114;
assign w643 = pi048 & ~w642;
assign w644 = w641 & ~w643;
assign w645 = ~pi062 & ~w117;
assign w646 = ~w318 & ~w645;
assign w647 = ~pi082 & ~w117;
assign w648 = pi048 & ~w647;
assign w649 = w646 & ~w648;
assign w650 = ~pi129 & ~w649;
assign w651 = ~w644 & w650;
assign w652 = ~pi045 & w112;
assign w653 = w111 & w652;
assign w654 = ~pi024 & ~pi048;
assign w655 = w106 & w654;
assign w656 = ~pi041 & w655;
assign w657 = w653 & w656;
assign w658 = pi049 & w253;
assign w659 = ~pi082 & ~w253;
assign w660 = pi049 & ~w659;
assign w661 = (~w657 & w658) | (~w657 & w660) | (w658 & w660);
assign w662 = ~pi069 & ~pi082;
assign w663 = ~w117 & w662;
assign w664 = ~pi069 & ~w117;
assign w665 = ~w318 & ~w664;
assign w666 = ~pi041 & w121;
assign w667 = ~w665 & w666;
assign w668 = ~w126 & ~w663;
assign w669 = (~w663 & ~w667) | (~w663 & w668) | (~w667 & w668);
assign w670 = ~w661 & w669;
assign w671 = ~pi129 & ~w670;
assign w672 = ~pi066 & ~w117;
assign w673 = ~w559 & ~w672;
assign w674 = pi050 & ~w647;
assign w675 = w673 & ~w674;
assign w676 = pi082 & ~w619;
assign w677 = ~pi038 & w526;
assign w678 = pi050 & ~w677;
assign w679 = w676 & ~w678;
assign w680 = ~pi129 & ~w679;
assign w681 = ~w675 & w680;
assign w682 = ~pi051 & pi109;
assign w683 = pi051 & ~pi109;
assign w684 = ~w682 & ~w683;
assign w685 = ~pi106 & w684;
assign w686 = ~pi129 & ~w685;
assign w687 = ~pi106 & ~w537;
assign w688 = pi052 & ~w682;
assign w689 = w687 & ~w688;
assign w690 = ~pi129 & ~w689;
assign w691 = ~w116 & ~w117;
assign w692 = ~pi129 & ~w691;
assign w693 = pi114 & ~pi122;
assign w694 = ~pi123 & w693;
assign w695 = ~pi129 & w694;
assign w696 = pi058 & ~pi116;
assign w697 = pi026 & pi116;
assign w698 = ~w696 & ~w697;
assign w699 = ~pi094 & ~w698;
assign w700 = ~pi026 & ~pi058;
assign w701 = pi026 & ~pi116;
assign w702 = ~w700 & ~w701;
assign w703 = ~pi037 & ~w702;
assign w704 = ~w699 & ~w703;
assign w705 = pi058 & pi085;
assign w706 = ~pi053 & ~w705;
assign w707 = ~pi027 & w335;
assign w708 = (~pi027 & w706) | (~pi027 & w707) | (w706 & w707);
assign w709 = ~pi026 & w339;
assign w710 = (~pi026 & w708) | (~pi026 & w709) | (w708 & w709);
assign w711 = w335 & w389;
assign w712 = w78 & w711;
assign w713 = (w78 & w710) | (w78 & w712) | (w710 & w712);
assign w714 = w704 & w713;
assign w715 = pi060 & w378;
assign w716 = pi057 & ~w378;
assign w717 = ~w715 & ~w716;
assign w718 = w713 & ~w717;
assign w719 = ~pi026 & ~pi116;
assign w720 = ~pi027 & pi058;
assign w721 = w719 & w720;
assign w722 = ~pi026 & pi027;
assign w723 = ~w340 & ~w722;
assign w724 = ~pi058 & ~w723;
assign w725 = w364 & w724;
assign w726 = ~w721 & ~w725;
assign w727 = w713 & ~w726;
assign w728 = pi059 & ~w351;
assign w729 = pi096 & w351;
assign w730 = ~w728 & ~w729;
assign w731 = w446 & ~w730;
assign w732 = pi059 & ~pi116;
assign w733 = ~w348 & w732;
assign w734 = ~w731 & ~w733;
assign w735 = w78 & ~w734;
assign w736 = ~pi117 & ~pi122;
assign w737 = pi123 & w736;
assign w738 = pi060 & ~w736;
assign w739 = ~w737 & ~w738;
assign w740 = ~pi114 & ~pi122;
assign w741 = pi123 & w740;
assign w742 = ~pi129 & w741;
assign w743 = pi131 & pi132;
assign w744 = pi133 & w743;
assign w745 = pi136 & w744;
assign w746 = ~pi137 & w745;
assign w747 = ~pi138 & w746;
assign w748 = ~pi140 & w747;
assign w749 = pi062 & ~w747;
assign w750 = ~w748 & ~w749;
assign w751 = ~pi129 & ~w750;
assign w752 = ~pi142 & w747;
assign w753 = pi063 & ~w747;
assign w754 = ~w752 & ~w753;
assign w755 = ~pi129 & ~w754;
assign w756 = ~pi139 & w747;
assign w757 = pi064 & ~w747;
assign w758 = ~w756 & ~w757;
assign w759 = ~pi129 & ~w758;
assign w760 = ~pi146 & w747;
assign w761 = pi065 & ~w747;
assign w762 = ~w760 & ~w761;
assign w763 = ~pi129 & ~w762;
assign w764 = ~pi136 & w744;
assign w765 = ~pi137 & w764;
assign w766 = ~pi138 & w765;
assign w767 = ~pi143 & w766;
assign w768 = pi066 & ~w766;
assign w769 = ~w767 & ~w768;
assign w770 = ~pi129 & ~w769;
assign w771 = ~pi139 & w766;
assign w772 = pi067 & ~w766;
assign w773 = ~w771 & ~w772;
assign w774 = ~pi129 & ~w773;
assign w775 = ~pi141 & w747;
assign w776 = pi068 & ~w747;
assign w777 = ~w775 & ~w776;
assign w778 = ~pi129 & ~w777;
assign w779 = ~pi143 & w747;
assign w780 = pi069 & ~w747;
assign w781 = ~w779 & ~w780;
assign w782 = ~pi129 & ~w781;
assign w783 = ~pi144 & w747;
assign w784 = pi070 & ~w747;
assign w785 = ~w783 & ~w784;
assign w786 = ~pi129 & ~w785;
assign w787 = ~pi145 & w747;
assign w788 = pi071 & ~w747;
assign w789 = ~w787 & ~w788;
assign w790 = ~pi129 & ~w789;
assign w791 = ~pi140 & w766;
assign w792 = pi072 & ~w766;
assign w793 = ~w791 & ~w792;
assign w794 = ~pi129 & ~w793;
assign w795 = ~pi141 & w766;
assign w796 = pi073 & ~w766;
assign w797 = ~w795 & ~w796;
assign w798 = ~pi129 & ~w797;
assign w799 = ~pi142 & w766;
assign w800 = pi074 & ~w766;
assign w801 = ~w799 & ~w800;
assign w802 = ~pi129 & ~w801;
assign w803 = ~pi144 & w766;
assign w804 = pi075 & ~w766;
assign w805 = ~w803 & ~w804;
assign w806 = ~pi129 & ~w805;
assign w807 = ~pi145 & w766;
assign w808 = pi076 & ~w766;
assign w809 = ~w807 & ~w808;
assign w810 = ~pi129 & ~w809;
assign w811 = ~pi146 & w766;
assign w812 = pi077 & ~w766;
assign w813 = ~w811 & ~w812;
assign w814 = ~pi129 & ~w813;
assign w815 = pi137 & w764;
assign w816 = ~pi138 & w815;
assign w817 = pi142 & w816;
assign w818 = pi078 & ~w816;
assign w819 = ~w817 & ~w818;
assign w820 = ~pi129 & ~w819;
assign w821 = pi143 & w816;
assign w822 = pi079 & ~w816;
assign w823 = ~w821 & ~w822;
assign w824 = ~pi129 & ~w823;
assign w825 = pi144 & w816;
assign w826 = pi080 & ~w816;
assign w827 = ~w825 & ~w826;
assign w828 = ~pi129 & ~w827;
assign w829 = pi145 & w816;
assign w830 = pi081 & ~w816;
assign w831 = ~w829 & ~w830;
assign w832 = ~pi129 & ~w831;
assign w833 = pi146 & w816;
assign w834 = pi082 & ~w816;
assign w835 = ~w833 & ~w834;
assign w836 = ~pi129 & ~w835;
assign w837 = ~pi119 & pi138;
assign w838 = pi072 & ~pi138;
assign w839 = ~w837 & ~w838;
assign w840 = ~pi137 & ~w839;
assign w841 = pi115 & pi138;
assign w842 = ~pi087 & ~pi138;
assign w843 = ~w841 & ~w842;
assign w844 = pi137 & ~w843;
assign w845 = ~w840 & ~w844;
assign w846 = ~pi136 & w845;
assign w847 = pi089 & pi138;
assign w848 = ~pi062 & ~pi138;
assign w849 = ~w847 & ~w848;
assign w850 = ~pi137 & ~w849;
assign w851 = pi137 & ~pi138;
assign w852 = pi031 & w851;
assign w853 = ~w850 & ~w852;
assign w854 = pi136 & ~w853;
assign w855 = ~w846 & ~w854;
assign w856 = pi141 & w816;
assign w857 = pi084 & ~w816;
assign w858 = ~w856 & ~w857;
assign w859 = ~pi129 & ~w858;
assign w860 = ~pi085 & w351;
assign w861 = pi096 & w860;
assign w862 = ~w354 & ~w861;
assign w863 = w392 & ~w862;
assign w864 = pi139 & w816;
assign w865 = pi086 & ~w816;
assign w866 = ~w864 & ~w865;
assign w867 = ~pi129 & ~w866;
assign w868 = pi140 & w816;
assign w869 = pi087 & ~w816;
assign w870 = ~w868 & ~w869;
assign w871 = ~pi129 & ~w870;
assign w872 = pi137 & w745;
assign w873 = ~pi138 & w872;
assign w874 = pi139 & w873;
assign w875 = pi088 & ~w873;
assign w876 = ~w874 & ~w875;
assign w877 = ~pi129 & ~w876;
assign w878 = pi140 & w873;
assign w879 = pi089 & ~w873;
assign w880 = ~w878 & ~w879;
assign w881 = ~pi129 & ~w880;
assign w882 = pi142 & w873;
assign w883 = pi090 & ~w873;
assign w884 = ~w882 & ~w883;
assign w885 = ~pi129 & ~w884;
assign w886 = pi143 & w873;
assign w887 = pi091 & ~w873;
assign w888 = ~w886 & ~w887;
assign w889 = ~pi129 & ~w888;
assign w890 = pi144 & w873;
assign w891 = pi092 & ~w873;
assign w892 = ~w890 & ~w891;
assign w893 = ~pi129 & ~w892;
assign w894 = pi146 & w873;
assign w895 = pi093 & ~w873;
assign w896 = ~w894 & ~w895;
assign w897 = ~pi129 & ~w896;
assign w898 = pi082 & ~pi136;
assign w899 = ~pi137 & w898;
assign w900 = pi138 & w899;
assign w901 = w744 & w900;
assign w902 = pi142 & w901;
assign w903 = pi094 & ~w901;
assign w904 = ~w902 & ~w903;
assign w905 = ~pi129 & ~w904;
assign w906 = pi143 & w901;
assign w907 = ~pi110 & ~w744;
assign w908 = ~pi003 & w907;
assign w909 = w744 & ~w900;
assign w910 = ~w908 & ~w909;
assign w911 = pi095 & ~w910;
assign w912 = ~w906 & ~w911;
assign w913 = ~pi129 & ~w912;
assign w914 = pi146 & w901;
assign w915 = pi096 & ~w910;
assign w916 = ~w914 & ~w915;
assign w917 = ~pi129 & ~w916;
assign w918 = pi145 & w901;
assign w919 = pi097 & ~w910;
assign w920 = ~w918 & ~w919;
assign w921 = ~pi129 & ~w920;
assign w922 = pi145 & w873;
assign w923 = pi098 & ~w873;
assign w924 = ~w922 & ~w923;
assign w925 = ~pi129 & ~w924;
assign w926 = pi141 & w873;
assign w927 = pi099 & ~w873;
assign w928 = ~w926 & ~w927;
assign w929 = ~pi129 & ~w928;
assign w930 = pi144 & w901;
assign w931 = pi100 & ~w910;
assign w932 = ~w930 & ~w931;
assign w933 = ~pi129 & ~w932;
assign w934 = ~pi077 & ~pi138;
assign w935 = pi124 & pi138;
assign w936 = ~w934 & ~w935;
assign w937 = ~pi137 & ~w936;
assign w938 = ~pi136 & w937;
assign w939 = pi037 & pi136;
assign w940 = w851 & w939;
assign w941 = ~w938 & ~w940;
assign w942 = pi136 & ~pi137;
assign w943 = pi093 & w942;
assign w944 = ~pi136 & pi137;
assign w945 = pi096 & w944;
assign w946 = ~w943 & ~w945;
assign w947 = pi138 & ~w946;
assign w948 = ~pi065 & w942;
assign w949 = pi082 & w944;
assign w950 = ~w948 & ~w949;
assign w951 = ~pi138 & ~w950;
assign w952 = ~w947 & ~w951;
assign w953 = w941 & w952;
assign w954 = pi091 & w942;
assign w955 = pi095 & w944;
assign w956 = ~w954 & ~w955;
assign w957 = pi138 & ~w956;
assign w958 = ~pi079 & pi137;
assign w959 = pi066 & ~pi137;
assign w960 = ~w958 & ~w959;
assign w961 = ~pi136 & ~w960;
assign w962 = pi069 & ~pi137;
assign w963 = ~pi034 & pi137;
assign w964 = ~w962 & ~w963;
assign w965 = pi136 & ~w964;
assign w966 = ~w961 & ~w965;
assign w967 = ~pi138 & w966;
assign w968 = ~w957 & ~w967;
assign w969 = pi090 & w942;
assign w970 = pi094 & w944;
assign w971 = ~w969 & ~w970;
assign w972 = pi138 & ~w971;
assign w973 = pi074 & ~pi137;
assign w974 = ~pi078 & pi137;
assign w975 = ~w973 & ~w974;
assign w976 = ~pi136 & ~w975;
assign w977 = ~pi033 & pi137;
assign w978 = pi063 & ~pi137;
assign w979 = ~w977 & ~w978;
assign w980 = pi136 & ~w979;
assign w981 = ~w976 & ~w980;
assign w982 = ~pi138 & w981;
assign w983 = ~w972 & ~w982;
assign w984 = ~pi112 & w944;
assign w985 = pi099 & w942;
assign w986 = ~w984 & ~w985;
assign w987 = pi138 & ~w986;
assign w988 = pi073 & ~pi137;
assign w989 = ~pi084 & pi137;
assign w990 = ~w988 & ~w989;
assign w991 = ~pi136 & ~w990;
assign w992 = ~pi032 & pi137;
assign w993 = pi068 & ~pi137;
assign w994 = ~w992 & ~w993;
assign w995 = pi136 & ~w994;
assign w996 = ~w991 & ~w995;
assign w997 = ~pi138 & w996;
assign w998 = ~w987 & ~w997;
assign w999 = ~pi075 & ~pi138;
assign w1000 = pi125 & pi138;
assign w1001 = ~w999 & ~w1000;
assign w1002 = ~pi137 & ~w1001;
assign w1003 = ~pi136 & w1002;
assign w1004 = pi035 & pi136;
assign w1005 = w851 & w1004;
assign w1006 = ~w1003 & ~w1005;
assign w1007 = pi092 & w942;
assign w1008 = pi100 & w944;
assign w1009 = ~w1007 & ~w1008;
assign w1010 = pi138 & ~w1009;
assign w1011 = ~pi070 & w942;
assign w1012 = pi080 & w944;
assign w1013 = ~w1011 & ~w1012;
assign w1014 = ~pi138 & ~w1013;
assign w1015 = ~w1010 & ~w1014;
assign w1016 = w1006 & w1015;
assign w1017 = w351 & w446;
assign w1018 = ~w386 & ~w1017;
assign w1019 = w78 & ~w1018;
assign w1020 = pi023 & pi138;
assign w1021 = ~pi076 & ~pi138;
assign w1022 = ~w1020 & ~w1021;
assign w1023 = ~pi137 & ~w1022;
assign w1024 = pi081 & ~pi138;
assign w1025 = pi097 & pi138;
assign w1026 = ~w1024 & ~w1025;
assign w1027 = pi137 & ~w1026;
assign w1028 = ~w1023 & ~w1027;
assign w1029 = ~pi136 & ~w1028;
assign w1030 = pi098 & pi138;
assign w1031 = ~pi071 & ~pi138;
assign w1032 = ~w1030 & ~w1031;
assign w1033 = ~pi137 & ~w1032;
assign w1034 = pi036 & w851;
assign w1035 = ~w1033 & ~w1034;
assign w1036 = pi136 & ~w1035;
assign w1037 = ~w1029 & ~w1036;
assign w1038 = ~pi111 & pi138;
assign w1039 = ~pi086 & ~pi138;
assign w1040 = ~w1038 & ~w1039;
assign w1041 = pi137 & ~w1040;
assign w1042 = ~pi120 & pi138;
assign w1043 = pi067 & ~pi138;
assign w1044 = ~w1042 & ~w1043;
assign w1045 = ~pi137 & ~w1044;
assign w1046 = ~w1041 & ~w1045;
assign w1047 = ~pi136 & w1046;
assign w1048 = pi088 & pi138;
assign w1049 = ~pi064 & ~pi138;
assign w1050 = ~w1048 & ~w1049;
assign w1051 = ~pi137 & ~w1050;
assign w1052 = pi030 & w851;
assign w1053 = ~w1051 & ~w1052;
assign w1054 = pi136 & ~w1053;
assign w1055 = ~w1047 & ~w1054;
assign w1056 = ~w374 & w722;
assign w1057 = ~w340 & ~w1056;
assign w1058 = pi116 & ~w1057;
assign w1059 = w78 & w1058;
assign w1060 = ~pi053 & pi058;
assign w1061 = ~pi097 & w1060;
assign w1062 = pi053 & ~pi058;
assign w1063 = ~w1061 & ~w1062;
assign w1064 = pi116 & ~w1063;
assign w1065 = w78 & w1064;
assign w1066 = pi111 & ~w900;
assign w1067 = pi139 & w900;
assign w1068 = ~w1066 & ~w1067;
assign w1069 = ~pi129 & ~w1068;
assign w1070 = w744 & w1069;
assign w1071 = pi141 & w900;
assign w1072 = ~pi112 & ~w900;
assign w1073 = ~w1071 & ~w1072;
assign w1074 = ~pi129 & ~w1073;
assign w1075 = w744 & w1074;
assign w1076 = ~pi011 & ~pi022;
assign w1077 = pi054 & ~w1076;
assign w1078 = ~pi054 & ~pi113;
assign w1079 = ~w1077 & ~w1078;
assign w1080 = w78 & ~w1079;
assign w1081 = ~pi123 & ~pi129;
assign w1082 = pi140 & w900;
assign w1083 = ~pi115 & ~w900;
assign w1084 = ~w1082 & ~w1083;
assign w1085 = ~pi129 & ~w1084;
assign w1086 = w744 & w1085;
assign w1087 = pi054 & ~w29;
assign w1088 = w78 & w1087;
assign w1089 = pi122 & ~pi129;
assign w1090 = ~pi054 & pi118;
assign w1091 = ~w230 & ~w1090;
assign w1092 = ~pi129 & ~w1091;
assign w1093 = ~pi129 & ~w349;
assign w1094 = ~pi003 & ~pi110;
assign w1095 = ~pi120 & w1094;
assign w1096 = ~pi129 & ~w1095;
assign w1097 = ~pi111 & w1096;
assign w1098 = pi081 & pi120;
assign w1099 = ~pi129 & w1098;
assign w1100 = ~pi129 & ~pi134;
assign w1101 = ~pi129 & ~pi135;
assign w1102 = pi057 & ~pi129;
assign w1103 = ~pi096 & pi125;
assign w1104 = ~pi003 & ~w1103;
assign w1105 = ~pi129 & ~w1104;
assign w1106 = ~pi126 & pi132;
assign w1107 = pi133 & w1106;
assign one = 1;
assign po000 = pi108;
assign po001 = pi083;
assign po002 = pi104;
assign po003 = pi103;
assign po004 = pi102;
assign po005 = pi105;
assign po006 = pi107;
assign po007 = pi101;
assign po008 = pi126;
assign po009 = pi121;
assign po010 = pi001;
assign po011 = pi000;
assign po012 = one;
assign po013 = pi130;
assign po014 = pi128;
assign po015 = ~w79;
assign po016 = w100;
assign po017 = w138;
assign po018 = w149;
assign po019 = w159;
assign po020 = ~w175;
assign po021 = ~w180;
assign po022 = w185;
assign po023 = w193;
assign po024 = w203;
assign po025 = w209;
assign po026 = w217;
assign po027 = w225;
assign po028 = w233;
assign po029 = w240;
assign po030 = w257;
assign po031 = ~w262;
assign po032 = w269;
assign po033 = w274;
assign po034 = w279;
assign po035 = w293;
assign po036 = w298;
assign po037 = w306;
assign po038 = w309;
assign po039 = w330;
assign po040 = ~w395;
assign po041 = ~w401;
assign po042 = ~w413;
assign po043 = w427;
assign po044 = w454;
assign po045 = w461;
assign po046 = w468;
assign po047 = w475;
assign po048 = w482;
assign po049 = w489;
assign po050 = w496;
assign po051 = w503;
assign po052 = w510;
assign po053 = w531;
assign po054 = w540;
assign po055 = w553;
assign po056 = w565;
assign po057 = w574;
assign po058 = w584;
assign po059 = w595;
assign po060 = w609;
assign po061 = w623;
assign po062 = w638;
assign po063 = w651;
assign po064 = w671;
assign po065 = w681;
assign po066 = w686;
assign po067 = w690;
assign po068 = w442;
assign po069 = ~w692;
assign po070 = w695;
assign po071 = w714;
assign po072 = w718;
assign po073 = w727;
assign po074 = w735;
assign po075 = ~w739;
assign po076 = w742;
assign po077 = ~w751;
assign po078 = ~w755;
assign po079 = ~w759;
assign po080 = ~w763;
assign po081 = ~w770;
assign po082 = ~w774;
assign po083 = ~w778;
assign po084 = ~w782;
assign po085 = ~w786;
assign po086 = ~w790;
assign po087 = ~w794;
assign po088 = ~w798;
assign po089 = ~w802;
assign po090 = ~w806;
assign po091 = ~w810;
assign po092 = ~w814;
assign po093 = w820;
assign po094 = w824;
assign po095 = w828;
assign po096 = w832;
assign po097 = w836;
assign po098 = ~w855;
assign po099 = w859;
assign po100 = w863;
assign po101 = w867;
assign po102 = w871;
assign po103 = w877;
assign po104 = w881;
assign po105 = w885;
assign po106 = w889;
assign po107 = w893;
assign po108 = w897;
assign po109 = w905;
assign po110 = w913;
assign po111 = w917;
assign po112 = w921;
assign po113 = w925;
assign po114 = w929;
assign po115 = w933;
assign po116 = ~w953;
assign po117 = ~w968;
assign po118 = ~w983;
assign po119 = ~w998;
assign po120 = ~w1016;
assign po121 = w1019;
assign po122 = ~w1037;
assign po123 = ~w1055;
assign po124 = w1059;
assign po125 = w1065;
assign po126 = w1070;
assign po127 = w1075;
assign po128 = w1080;
assign po129 = ~w1081;
assign po130 = w1086;
assign po131 = w1088;
assign po132 = ~w1089;
assign po133 = w1092;
assign po134 = w1093;
assign po135 = w1097;
assign po136 = w1099;
assign po137 = ~w1100;
assign po138 = ~w1101;
assign po139 = w1102;
assign po140 = w1105;
assign po141 = w1107;
endmodule

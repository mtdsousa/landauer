//Written by the Majority Logic Package Thu Jun 18 13:34:09 2015
module top (
            a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27], a[28], a[29], a[30], a[31], a[32], a[33], a[34], a[35], a[36], a[37], a[38], a[39], a[40], a[41], a[42], a[43], a[44], a[45], a[46], a[47], a[48], a[49], a[50], a[51], a[52], a[53], a[54], a[55], a[56], a[57], a[58], a[59], a[60], a[61], a[62], a[63], a[64], a[65], a[66], a[67], a[68], a[69], a[70], a[71], a[72], a[73], a[74], a[75], a[76], a[77], a[78], a[79], a[80], a[81], a[82], a[83], a[84], a[85], a[86], a[87], a[88], a[89], a[90], a[91], a[92], a[93], a[94], a[95], a[96], a[97], a[98], a[99], a[100], a[101], a[102], a[103], a[104], a[105], a[106], a[107], a[108], a[109], a[110], a[111], a[112], a[113], a[114], a[115], a[116], a[117], a[118], a[119], a[120], a[121], a[122], a[123], a[124], a[125], a[126], a[127], 
            asqrt[0], asqrt[1], asqrt[2], asqrt[3], asqrt[4], asqrt[5], asqrt[6], asqrt[7], asqrt[8], asqrt[9], asqrt[10], asqrt[11], asqrt[12], asqrt[13], asqrt[14], asqrt[15], asqrt[16], asqrt[17], asqrt[18], asqrt[19], asqrt[20], asqrt[21], asqrt[22], asqrt[23], asqrt[24], asqrt[25], asqrt[26], asqrt[27], asqrt[28], asqrt[29], asqrt[30], asqrt[31], asqrt[32], asqrt[33], asqrt[34], asqrt[35], asqrt[36], asqrt[37], asqrt[38], asqrt[39], asqrt[40], asqrt[41], asqrt[42], asqrt[43], asqrt[44], asqrt[45], asqrt[46], asqrt[47], asqrt[48], asqrt[49], asqrt[50], asqrt[51], asqrt[52], asqrt[53], asqrt[54], asqrt[55], asqrt[56], asqrt[57], asqrt[58], asqrt[59], asqrt[60], asqrt[61], asqrt[62], asqrt[63]);
input a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27], a[28], a[29], a[30], a[31], a[32], a[33], a[34], a[35], a[36], a[37], a[38], a[39], a[40], a[41], a[42], a[43], a[44], a[45], a[46], a[47], a[48], a[49], a[50], a[51], a[52], a[53], a[54], a[55], a[56], a[57], a[58], a[59], a[60], a[61], a[62], a[63], a[64], a[65], a[66], a[67], a[68], a[69], a[70], a[71], a[72], a[73], a[74], a[75], a[76], a[77], a[78], a[79], a[80], a[81], a[82], a[83], a[84], a[85], a[86], a[87], a[88], a[89], a[90], a[91], a[92], a[93], a[94], a[95], a[96], a[97], a[98], a[99], a[100], a[101], a[102], a[103], a[104], a[105], a[106], a[107], a[108], a[109], a[110], a[111], a[112], a[113], a[114], a[115], a[116], a[117], a[118], a[119], a[120], a[121], a[122], a[123], a[124], a[125], a[126], a[127];
output asqrt[0], asqrt[1], asqrt[2], asqrt[3], asqrt[4], asqrt[5], asqrt[6], asqrt[7], asqrt[8], asqrt[9], asqrt[10], asqrt[11], asqrt[12], asqrt[13], asqrt[14], asqrt[15], asqrt[16], asqrt[17], asqrt[18], asqrt[19], asqrt[20], asqrt[21], asqrt[22], asqrt[23], asqrt[24], asqrt[25], asqrt[26], asqrt[27], asqrt[28], asqrt[29], asqrt[30], asqrt[31], asqrt[32], asqrt[33], asqrt[34], asqrt[35], asqrt[36], asqrt[37], asqrt[38], asqrt[39], asqrt[40], asqrt[41], asqrt[42], asqrt[43], asqrt[44], asqrt[45], asqrt[46], asqrt[47], asqrt[48], asqrt[49], asqrt[50], asqrt[51], asqrt[52], asqrt[53], asqrt[54], asqrt[55], asqrt[56], asqrt[57], asqrt[58], asqrt[59], asqrt[60], asqrt[61], asqrt[62], asqrt[63];
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935, w41936, w41937, w41938, w41939, w41940, w41941, w41942, w41943, w41944, w41945, w41946, w41947, w41948, w41949, w41950, w41951, w41952, w41953, w41954, w41955, w41956, w41957, w41958, w41959, w41960, w41961, w41962, w41963, w41964, w41965, w41966, w41967, w41968, w41969, w41970, w41971, w41972, w41973, w41974, w41975, w41976, w41977, w41978, w41979, w41980, w41981, w41982, w41983, w41984, w41985, w41986, w41987, w41988, w41989, w41990, w41991, w41992, w41993, w41994, w41995, w41996, w41997, w41998, w41999, w42000, w42001, w42002, w42003, w42004, w42005, w42006, w42007, w42008, w42009, w42010, w42011, w42012, w42013, w42014, w42015, w42016, w42017, w42018, w42019, w42020, w42021, w42022, w42023, w42024, w42025, w42026, w42027, w42028, w42029, w42030, w42031, w42032, w42033, w42034, w42035, w42036, w42037, w42038, w42039, w42040, w42041, w42042, w42043, w42044, w42045, w42046, w42047, w42048, w42049, w42050, w42051, w42052, w42053, w42054, w42055, w42056, w42057, w42058, w42059, w42060, w42061, w42062, w42063, w42064, w42065, w42066, w42067, w42068, w42069, w42070, w42071, w42072, w42073, w42074, w42075, w42076, w42077, w42078, w42079, w42080, w42081, w42082, w42083, w42084, w42085, w42086, w42087, w42088, w42089, w42090, w42091, w42092, w42093, w42094, w42095, w42096, w42097, w42098, w42099, w42100, w42101, w42102, w42103, w42104, w42105, w42106, w42107, w42108, w42109, w42110, w42111, w42112, w42113, w42114, w42115, w42116, w42117, w42118, w42119, w42120, w42121, w42122, w42123, w42124, w42125, w42126, w42127, w42128, w42129, w42130, w42131, w42132, w42133, w42134, w42135, w42136, w42137, w42138, w42139, w42140, w42141, w42142, w42143, w42144, w42145, w42146, w42147, w42148, w42149, w42150, w42151, w42152, w42153, w42154, w42155, w42156, w42157, w42158, w42159, w42160, w42161, w42162, w42163, w42164, w42165, w42166, w42167, w42168, w42169, w42170, w42171, w42172, w42173, w42174, w42175, w42176, w42177, w42178, w42179, w42180, w42181, w42182, w42183, w42184, w42185, w42186, w42187, w42188, w42189, w42190, w42191, w42192, w42193, w42194, w42195, w42196, w42197, w42198, w42199, w42200, w42201, w42202, w42203, w42204, w42205, w42206, w42207, w42208, w42209, w42210, w42211, w42212, w42213, w42214, w42215, w42216, w42217, w42218, w42219, w42220, w42221, w42222, w42223, w42224, w42225, w42226, w42227, w42228, w42229, w42230, w42231, w42232, w42233, w42234, w42235, w42236, w42237, w42238, w42239, w42240, w42241, w42242, w42243, w42244, w42245, w42246, w42247, w42248, w42249, w42250, w42251, w42252, w42253, w42254, w42255, w42256, w42257, w42258, w42259, w42260, w42261, w42262, w42263, w42264, w42265, w42266, w42267, w42268, w42269, w42270, w42271, w42272, w42273, w42274, w42275, w42276, w42277, w42278, w42279, w42280, w42281, w42282, w42283, w42284, w42285, w42286, w42287, w42288, w42289, w42290, w42291, w42292, w42293, w42294, w42295, w42296, w42297, w42298, w42299, w42300, w42301, w42302, w42303, w42304, w42305, w42306, w42307, w42308, w42309, w42310, w42311, w42312, w42313, w42314, w42315, w42316, w42317, w42318, w42319, w42320, w42321, w42322, w42323, w42324, w42325, w42326, w42327, w42328, w42329, w42330, w42331, w42332, w42333, w42334, w42335, w42336, w42337, w42338, w42339, w42340, w42341, w42342, w42343, w42344, w42345, w42346, w42347, w42348, w42349, w42350, w42351, w42352, w42353, w42354, w42355, w42356, w42357, w42358, w42359, w42360, w42361, w42362, w42363, w42364, w42365, w42366, w42367, w42368, w42369, w42370, w42371, w42372, w42373, w42374, w42375, w42376, w42377, w42378, w42379, w42380, w42381, w42382, w42383, w42384, w42385, w42386, w42387, w42388, w42389, w42390, w42391, w42392, w42393, w42394, w42395, w42396, w42397, w42398, w42399, w42400, w42401, w42402, w42403, w42404, w42405, w42406, w42407, w42408, w42409, w42410, w42411, w42412, w42413, w42414, w42415, w42416, w42417, w42418, w42419, w42420, w42421, w42422, w42423, w42424, w42425, w42426, w42427, w42428, w42429, w42430, w42431, w42432, w42433, w42434, w42435, w42436, w42437, w42438, w42439, w42440, w42441, w42442, w42443, w42444, w42445, w42446, w42447, w42448, w42449, w42450, w42451, w42452, w42453, w42454, w42455, w42456, w42457, w42458, w42459, w42460, w42461, w42462, w42463, w42464, w42465, w42466, w42467, w42468, w42469, w42470, w42471, w42472, w42473, w42474, w42475, w42476, w42477, w42478, w42479, w42480, w42481, w42482, w42483, w42484, w42485, w42486, w42487, w42488, w42489, w42490, w42491, w42492, w42493, w42494, w42495, w42496, w42497, w42498, w42499, w42500, w42501, w42502, w42503, w42504, w42505, w42506, w42507, w42508, w42509, w42510, w42511, w42512, w42513, w42514, w42515, w42516, w42517, w42518, w42519, w42520, w42521, w42522, w42523, w42524, w42525, w42526, w42527, w42528, w42529, w42530, w42531, w42532, w42533, w42534, w42535, w42536, w42537, w42538, w42539, w42540, w42541, w42542, w42543, w42544, w42545, w42546, w42547, w42548, w42549, w42550, w42551, w42552, w42553, w42554, w42555, w42556, w42557, w42558, w42559, w42560, w42561, w42562, w42563, w42564, w42565, w42566, w42567, w42568, w42569, w42570, w42571, w42572, w42573, w42574, w42575, w42576, w42577, w42578, w42579, w42580, w42581, w42582, w42583, w42584, w42585, w42586, w42587, w42588, w42589, w42590, w42591, w42592, w42593, w42594, w42595, w42596, w42597, w42598, w42599, w42600, w42601, w42602, w42603, w42604, w42605, w42606, w42607, w42608, w42609, w42610, w42611, w42612, w42613, w42614, w42615, w42616, w42617, w42618, w42619, w42620, w42621, w42622, w42623, w42624, w42625, w42626, w42627, w42628, w42629, w42630, w42631, w42632, w42633, w42634, w42635, w42636, w42637, w42638, w42639, w42640, w42641, w42642, w42643, w42644, w42645, w42646, w42647, w42648, w42649, w42650, w42651, w42652, w42653, w42654, w42655, w42656, w42657, w42658, w42659, w42660, w42661, w42662, w42663, w42664, w42665, w42666, w42667, w42668, w42669, w42670, w42671, w42672, w42673, w42674, w42675, w42676, w42677, w42678, w42679, w42680, w42681, w42682, w42683, w42684, w42685, w42686, w42687, w42688, w42689, w42690, w42691, w42692, w42693, w42694, w42695, w42696, w42697, w42698, w42699, w42700, w42701, w42702, w42703, w42704, w42705, w42706, w42707, w42708, w42709, w42710, w42711, w42712, w42713, w42714, w42715, w42716, w42717, w42718, w42719, w42720, w42721, w42722, w42723, w42724, w42725, w42726, w42727, w42728, w42729, w42730, w42731, w42732, w42733, w42734, w42735, w42736, w42737, w42738, w42739, w42740, w42741, w42742, w42743, w42744, w42745, w42746, w42747, w42748, w42749, w42750, w42751, w42752, w42753, w42754, w42755, w42756, w42757, w42758, w42759, w42760, w42761, w42762, w42763, w42764, w42765, w42766, w42767, w42768, w42769, w42770, w42771, w42772, w42773, w42774, w42775, w42776, w42777, w42778, w42779, w42780, w42781, w42782, w42783, w42784, w42785, w42786, w42787, w42788, w42789, w42790, w42791, w42792, w42793, w42794, w42795, w42796, w42797, w42798, w42799, w42800, w42801, w42802, w42803, w42804, w42805, w42806, w42807, w42808, w42809, w42810, w42811, w42812, w42813, w42814, w42815, w42816, w42817, w42818, w42819, w42820, w42821, w42822, w42823, w42824, w42825, w42826, w42827, w42828, w42829, w42830, w42831, w42832, w42833, w42834, w42835, w42836, w42837, w42838, w42839, w42840, w42841, w42842, w42843, w42844, w42845, w42846, w42847, w42848, w42849, w42850, w42851, w42852, w42853, w42854, w42855, w42856, w42857, w42858, w42859, w42860, w42861, w42862, w42863, w42864, w42865, w42866, w42867, w42868, w42869, w42870, w42871, w42872, w42873, w42874, w42875, w42876, w42877, w42878, w42879, w42880, w42881, w42882, w42883, w42884, w42885, w42886, w42887, w42888, w42889, w42890, w42891, w42892, w42893, w42894, w42895, w42896, w42897, w42898, w42899, w42900, w42901, w42902, w42903, w42904, w42905, w42906, w42907, w42908, w42909, w42910, w42911, w42912, w42913, w42914, w42915, w42916, w42917, w42918, w42919, w42920, w42921, w42922, w42923, w42924, w42925, w42926, w42927, w42928, w42929, w42930, w42931, w42932, w42933, w42934, w42935, w42936, w42937, w42938, w42939, w42940, w42941, w42942, w42943, w42944, w42945, w42946, w42947, w42948, w42949, w42950, w42951, w42952, w42953, w42954, w42955, w42956, w42957, w42958, w42959, w42960, w42961, w42962, w42963, w42964, w42965, w42966, w42967, w42968, w42969, w42970, w42971, w42972, w42973, w42974, w42975, w42976, w42977, w42978, w42979, w42980, w42981, w42982, w42983, w42984, w42985, w42986, w42987, w42988, w42989, w42990, w42991, w42992, w42993, w42994, w42995, w42996, w42997, w42998, w42999, w43000, w43001, w43002, w43003, w43004, w43005, w43006, w43007, w43008, w43009, w43010, w43011, w43012, w43013, w43014, w43015, w43016, w43017, w43018, w43019, w43020, w43021, w43022, w43023, w43024, w43025, w43026, w43027, w43028, w43029, w43030, w43031, w43032, w43033, w43034, w43035, w43036, w43037, w43038, w43039, w43040, w43041, w43042, w43043, w43044, w43045, w43046, w43047, w43048, w43049, w43050, w43051, w43052, w43053, w43054, w43055, w43056, w43057, w43058, w43059, w43060, w43061, w43062, w43063, w43064, w43065, w43066, w43067, w43068, w43069, w43070, w43071, w43072, w43073, w43074, w43075, w43076, w43077, w43078, w43079, w43080, w43081, w43082, w43083, w43084, w43085, w43086, w43087, w43088, w43089, w43090, w43091, w43092, w43093, w43094, w43095, w43096, w43097, w43098, w43099, w43100, w43101, w43102, w43103, w43104, w43105, w43106, w43107, w43108, w43109, w43110, w43111, w43112, w43113, w43114, w43115, w43116, w43117, w43118, w43119, w43120, w43121, w43122, w43123, w43124, w43125, w43126, w43127, w43128, w43129, w43130, w43131, w43132, w43133, w43134, w43135, w43136, w43137, w43138, w43139, w43140, w43141, w43142, w43143, w43144, w43145, w43146, w43147, w43148, w43149, w43150, w43151, w43152, w43153, w43154, w43155, w43156, w43157, w43158, w43159, w43160, w43161, w43162, w43163, w43164, w43165, w43166, w43167, w43168, w43169, w43170, w43171, w43172, w43173, w43174, w43175, w43176, w43177, w43178, w43179, w43180, w43181, w43182, w43183, w43184, w43185, w43186, w43187, w43188, w43189, w43190, w43191, w43192, w43193, w43194, w43195, w43196, w43197, w43198, w43199, w43200, w43201, w43202, w43203, w43204, w43205, w43206, w43207, w43208, w43209, w43210, w43211, w43212, w43213, w43214, w43215, w43216, w43217, w43218, w43219, w43220, w43221, w43222, w43223, w43224, w43225, w43226, w43227, w43228, w43229, w43230, w43231, w43232, w43233, w43234, w43235, w43236, w43237, w43238, w43239, w43240, w43241, w43242, w43243, w43244, w43245, w43246, w43247, w43248, w43249, w43250, w43251, w43252, w43253, w43254, w43255, w43256, w43257, w43258, w43259, w43260, w43261, w43262, w43263, w43264, w43265, w43266, w43267, w43268, w43269, w43270, w43271, w43272, w43273, w43274, w43275, w43276, w43277, w43278, w43279, w43280, w43281, w43282, w43283, w43284, w43285, w43286, w43287, w43288, w43289, w43290, w43291, w43292, w43293, w43294, w43295, w43296, w43297, w43298, w43299, w43300, w43301, w43302, w43303, w43304, w43305, w43306, w43307, w43308, w43309, w43310, w43311, w43312, w43313, w43314, w43315, w43316, w43317, w43318, w43319, w43320, w43321, w43322, w43323, w43324, w43325, w43326, w43327, w43328, w43329, w43330, w43331, w43332, w43333, w43334, w43335, w43336, w43337, w43338, w43339, w43340, w43341, w43342, w43343, w43344, w43345, w43346, w43347, w43348, w43349, w43350, w43351, w43352, w43353, w43354, w43355, w43356, w43357, w43358, w43359, w43360, w43361, w43362, w43363, w43364, w43365, w43366, w43367, w43368, w43369, w43370, w43371, w43372, w43373, w43374, w43375, w43376, w43377, w43378, w43379, w43380, w43381, w43382, w43383, w43384, w43385, w43386, w43387, w43388, w43389, w43390, w43391, w43392, w43393, w43394, w43395, w43396, w43397, w43398, w43399, w43400, w43401, w43402, w43403, w43404, w43405, w43406, w43407, w43408, w43409, w43410, w43411, w43412, w43413, w43414, w43415, w43416, w43417, w43418, w43419, w43420, w43421, w43422, w43423, w43424, w43425, w43426, w43427, w43428, w43429, w43430, w43431, w43432, w43433, w43434, w43435, w43436, w43437, w43438, w43439, w43440, w43441, w43442, w43443, w43444, w43445, w43446, w43447, w43448, w43449, w43450, w43451, w43452, w43453, w43454, w43455, w43456, w43457, w43458, w43459, w43460, w43461, w43462, w43463, w43464, w43465, w43466, w43467, w43468, w43469, w43470, w43471, w43472, w43473, w43474, w43475, w43476, w43477, w43478, w43479, w43480, w43481, w43482, w43483, w43484, w43485, w43486, w43487, w43488, w43489, w43490, w43491, w43492, w43493, w43494, w43495, w43496, w43497, w43498, w43499, w43500, w43501, w43502, w43503, w43504, w43505, w43506, w43507, w43508, w43509, w43510, w43511, w43512, w43513, w43514, w43515, w43516, w43517, w43518, w43519, w43520, w43521, w43522, w43523, w43524, w43525, w43526, w43527, w43528, w43529, w43530, w43531, w43532, w43533, w43534, w43535, w43536, w43537, w43538, w43539, w43540, w43541, w43542, w43543, w43544, w43545, w43546, w43547, w43548, w43549, w43550, w43551, w43552, w43553, w43554, w43555, w43556, w43557, w43558, w43559, w43560, w43561, w43562, w43563, w43564, w43565, w43566, w43567, w43568, w43569, w43570, w43571, w43572, w43573, w43574, w43575, w43576, w43577, w43578, w43579, w43580, w43581, w43582, w43583, w43584, w43585, w43586, w43587, w43588, w43589, w43590, w43591, w43592, w43593, w43594, w43595, w43596, w43597, w43598, w43599, w43600, w43601, w43602, w43603, w43604, w43605, w43606, w43607, w43608, w43609, w43610, w43611, w43612, w43613, w43614, w43615, w43616, w43617, w43618, w43619, w43620, w43621, w43622, w43623, w43624, w43625, w43626, w43627, w43628, w43629, w43630, w43631, w43632, w43633, w43634, w43635, w43636, w43637, w43638, w43639, w43640, w43641, w43642, w43643, w43644, w43645, w43646, w43647, w43648, w43649, w43650, w43651, w43652, w43653, w43654, w43655, w43656, w43657, w43658, w43659, w43660, w43661, w43662, w43663, w43664, w43665, w43666, w43667, w43668, w43669, w43670, w43671, w43672, w43673, w43674, w43675, w43676, w43677, w43678, w43679, w43680, w43681, w43682, w43683, w43684, w43685, w43686, w43687, w43688, w43689, w43690, w43691, w43692, w43693, w43694, w43695, w43696, w43697, w43698, w43699, w43700, w43701, w43702, w43703, w43704, w43705, w43706, w43707, w43708, w43709, w43710, w43711, w43712, w43713, w43714, w43715, w43716, w43717, w43718, w43719, w43720, w43721, w43722, w43723, w43724, w43725, w43726, w43727, w43728, w43729, w43730, w43731, w43732, w43733, w43734, w43735, w43736, w43737, w43738, w43739, w43740, w43741, w43742, w43743, w43744, w43745, w43746, w43747, w43748, w43749, w43750, w43751, w43752, w43753, w43754, w43755, w43756, w43757, w43758, w43759, w43760, w43761, w43762, w43763, w43764, w43765, w43766, w43767, w43768, w43769, w43770, w43771, w43772, w43773, w43774, w43775, w43776, w43777, w43778, w43779, w43780, w43781, w43782, w43783, w43784, w43785, w43786, w43787, w43788, w43789, w43790, w43791, w43792, w43793, w43794, w43795, w43796, w43797, w43798, w43799, w43800, w43801, w43802, w43803, w43804, w43805, w43806, w43807, w43808, w43809, w43810, w43811, w43812, w43813, w43814, w43815, w43816, w43817, w43818, w43819, w43820, w43821, w43822, w43823, w43824, w43825, w43826, w43827, w43828, w43829, w43830, w43831, w43832, w43833, w43834, w43835, w43836, w43837, w43838, w43839, w43840, w43841, w43842, w43843, w43844, w43845, w43846, w43847, w43848, w43849, w43850, w43851, w43852, w43853, w43854, w43855, w43856, w43857, w43858, w43859, w43860, w43861, w43862, w43863, w43864, w43865, w43866, w43867, w43868, w43869, w43870, w43871, w43872, w43873, w43874, w43875, w43876, w43877, w43878, w43879, w43880, w43881, w43882, w43883, w43884, w43885, w43886, w43887, w43888, w43889, w43890, w43891, w43892, w43893, w43894, w43895, w43896, w43897, w43898, w43899, w43900, w43901, w43902, w43903, w43904, w43905, w43906, w43907, w43908, w43909, w43910, w43911, w43912, w43913, w43914, w43915, w43916, w43917, w43918, w43919, w43920, w43921, w43922, w43923, w43924, w43925, w43926, w43927, w43928, w43929, w43930, w43931, w43932, w43933, w43934, w43935, w43936, w43937, w43938, w43939, w43940, w43941, w43942, w43943, w43944, w43945, w43946, w43947, w43948, w43949, w43950, w43951, w43952, w43953, w43954, w43955, w43956, w43957, w43958, w43959, w43960, w43961, w43962, w43963, w43964, w43965, w43966, w43967, w43968, w43969, w43970, w43971, w43972, w43973, w43974, w43975, w43976, w43977, w43978, w43979, w43980, w43981, w43982, w43983, w43984, w43985, w43986, w43987, w43988, w43989, w43990, w43991, w43992, w43993, w43994, w43995, w43996, w43997, w43998, w43999, w44000, w44001, w44002, w44003, w44004, w44005, w44006, w44007, w44008, w44009, w44010, w44011, w44012, w44013, w44014, w44015, w44016, w44017, w44018, w44019, w44020, w44021, w44022, w44023, w44024, w44025, w44026, w44027, w44028, w44029, w44030, w44031, w44032, w44033, w44034, w44035, w44036, w44037, w44038, w44039, w44040, w44041, w44042, w44043, w44044, w44045, w44046, w44047, w44048, w44049, w44050, w44051, w44052, w44053, w44054, w44055, w44056, w44057, w44058, w44059, w44060, w44061, w44062, w44063, w44064, w44065, w44066, w44067, w44068, w44069, w44070, w44071, w44072, w44073, w44074, w44075, w44076, w44077, w44078, w44079, w44080, w44081, w44082, w44083, w44084, w44085, w44086, w44087, w44088, w44089, w44090, w44091, w44092, w44093, w44094, w44095, w44096, w44097, w44098, w44099, w44100, w44101, w44102, w44103, w44104, w44105, w44106, w44107, w44108, w44109, w44110, w44111, w44112, w44113, w44114, w44115, w44116, w44117, w44118, w44119, w44120, w44121, w44122, w44123, w44124, w44125, w44126, w44127, w44128, w44129, w44130, w44131, w44132, w44133, w44134, w44135, w44136, w44137, w44138, w44139, w44140, w44141, w44142, w44143, w44144, w44145, w44146, w44147, w44148, w44149, w44150, w44151, w44152, w44153, w44154, w44155, w44156, w44157, w44158, w44159, w44160, w44161, w44162, w44163, w44164, w44165, w44166, w44167, w44168, w44169, w44170, w44171, w44172, w44173, w44174, w44175, w44176, w44177, w44178, w44179, w44180, w44181, w44182, w44183, w44184, w44185, w44186, w44187, w44188, w44189, w44190, w44191, w44192, w44193, w44194, w44195, w44196, w44197, w44198, w44199, w44200, w44201, w44202, w44203, w44204, w44205, w44206, w44207, w44208, w44209, w44210, w44211, w44212, w44213, w44214, w44215, w44216, w44217, w44218, w44219, w44220, w44221, w44222, w44223, w44224, w44225, w44226, w44227, w44228, w44229, w44230, w44231, w44232, w44233, w44234, w44235, w44236, w44237, w44238, w44239, w44240, w44241, w44242, w44243, w44244, w44245, w44246, w44247, w44248, w44249, w44250, w44251, w44252, w44253, w44254, w44255, w44256, w44257, w44258, w44259, w44260, w44261, w44262, w44263, w44264, w44265, w44266, w44267, w44268, w44269, w44270, w44271, w44272, w44273, w44274, w44275, w44276, w44277, w44278, w44279, w44280, w44281, w44282, w44283, w44284, w44285, w44286, w44287, w44288, w44289, w44290, w44291, w44292, w44293, w44294, w44295, w44296, w44297, w44298, w44299, w44300, w44301, w44302, w44303, w44304, w44305, w44306, w44307, w44308, w44309, w44310, w44311, w44312, w44313, w44314, w44315, w44316, w44317, w44318, w44319, w44320, w44321, w44322, w44323, w44324, w44325, w44326, w44327, w44328, w44329, w44330, w44331, w44332, w44333, w44334, w44335, w44336, w44337, w44338, w44339, w44340, w44341, w44342, w44343, w44344, w44345, w44346, w44347, w44348, w44349, w44350, w44351, w44352, w44353, w44354, w44355, w44356, w44357, w44358, w44359, w44360, w44361, w44362, w44363, w44364, w44365, w44366, w44367, w44368, w44369, w44370, w44371, w44372, w44373, w44374, w44375, w44376, w44377, w44378, w44379, w44380, w44381, w44382, w44383, w44384, w44385, w44386, w44387, w44388, w44389, w44390, w44391, w44392, w44393, w44394, w44395, w44396, w44397, w44398, w44399, w44400, w44401, w44402, w44403, w44404, w44405, w44406, w44407, w44408, w44409, w44410, w44411, w44412, w44413, w44414, w44415, w44416, w44417, w44418, w44419, w44420, w44421, w44422, w44423, w44424, w44425, w44426, w44427, w44428, w44429, w44430, w44431, w44432, w44433, w44434, w44435, w44436, w44437, w44438, w44439, w44440, w44441, w44442, w44443, w44444, w44445, w44446, w44447, w44448, w44449, w44450, w44451, w44452, w44453, w44454, w44455, w44456, w44457, w44458, w44459, w44460, w44461, w44462, w44463, w44464, w44465, w44466, w44467, w44468, w44469, w44470, w44471, w44472, w44473, w44474, w44475, w44476, w44477, w44478, w44479, w44480, w44481, w44482, w44483, w44484, w44485, w44486, w44487, w44488, w44489, w44490, w44491, w44492, w44493, w44494, w44495, w44496, w44497, w44498, w44499, w44500, w44501, w44502, w44503, w44504, w44505, w44506, w44507, w44508, w44509, w44510, w44511, w44512, w44513, w44514, w44515, w44516, w44517, w44518, w44519, w44520, w44521, w44522, w44523, w44524, w44525, w44526, w44527, w44528, w44529, w44530, w44531, w44532, w44533, w44534, w44535, w44536, w44537, w44538, w44539, w44540, w44541, w44542, w44543, w44544, w44545, w44546, w44547, w44548, w44549, w44550, w44551, w44552, w44553, w44554, w44555, w44556, w44557, w44558, w44559, w44560, w44561, w44562, w44563, w44564, w44565, w44566, w44567, w44568, w44569, w44570, w44571, w44572, w44573, w44574, w44575, w44576, w44577, w44578, w44579, w44580, w44581, w44582, w44583, w44584, w44585, w44586, w44587, w44588, w44589, w44590, w44591, w44592, w44593, w44594, w44595, w44596, w44597, w44598, w44599, w44600, w44601, w44602, w44603, w44604, w44605, w44606, w44607, w44608, w44609, w44610, w44611, w44612, w44613, w44614, w44615, w44616, w44617, w44618, w44619, w44620, w44621, w44622, w44623, w44624, w44625, w44626, w44627, w44628, w44629, w44630, w44631, w44632, w44633, w44634, w44635, w44636, w44637, w44638, w44639, w44640, w44641, w44642, w44643, w44644, w44645, w44646, w44647, w44648, w44649, w44650, w44651, w44652, w44653, w44654, w44655, w44656, w44657, w44658, w44659, w44660, w44661, w44662, w44663, w44664, w44665, w44666, w44667, w44668, w44669, w44670, w44671, w44672, w44673, w44674, w44675, w44676, w44677, w44678, w44679, w44680, w44681, w44682, w44683, w44684, w44685, w44686, w44687, w44688, w44689, w44690, w44691, w44692, w44693, w44694, w44695, w44696, w44697, w44698, w44699, w44700, w44701, w44702, w44703, w44704, w44705, w44706, w44707, w44708, w44709, w44710, w44711, w44712, w44713, w44714, w44715, w44716, w44717, w44718, w44719, w44720, w44721, w44722, w44723, w44724, w44725, w44726, w44727, w44728, w44729, w44730, w44731, w44732, w44733, w44734, w44735, w44736, w44737, w44738, w44739, w44740, w44741, w44742, w44743, w44744, w44745, w44746, w44747, w44748, w44749, w44750, w44751, w44752, w44753, w44754, w44755, w44756, w44757, w44758, w44759, w44760, w44761, w44762, w44763, w44764, w44765, w44766, w44767, w44768, w44769, w44770, w44771, w44772, w44773, w44774, w44775, w44776, w44777, w44778, w44779, w44780, w44781, w44782, w44783, w44784, w44785, w44786, w44787, w44788, w44789, w44790, w44791, w44792, w44793, w44794, w44795, w44796, w44797, w44798, w44799, w44800, w44801, w44802, w44803, w44804, w44805, w44806, w44807, w44808, w44809, w44810, w44811, w44812, w44813, w44814, w44815, w44816, w44817, w44818, w44819, w44820, w44821, w44822, w44823, w44824, w44825, w44826, w44827, w44828, w44829, w44830, w44831, w44832, w44833, w44834, w44835, w44836, w44837, w44838, w44839, w44840, w44841, w44842, w44843, w44844, w44845, w44846, w44847, w44848, w44849, w44850, w44851, w44852, w44853, w44854, w44855, w44856, w44857, w44858, w44859, w44860, w44861, w44862, w44863, w44864, w44865, w44866, w44867, w44868, w44869, w44870, w44871, w44872, w44873, w44874, w44875, w44876, w44877, w44878, w44879, w44880, w44881, w44882, w44883, w44884, w44885, w44886, w44887, w44888, w44889, w44890, w44891, w44892, w44893, w44894, w44895, w44896, w44897, w44898, w44899, w44900, w44901, w44902, w44903, w44904, w44905, w44906, w44907, w44908, w44909, w44910, w44911, w44912, w44913, w44914, w44915, w44916, w44917, w44918, w44919, w44920, w44921, w44922, w44923, w44924, w44925, w44926, w44927, w44928, w44929, w44930, w44931, w44932, w44933, w44934, w44935, w44936, w44937, w44938, w44939, w44940, w44941, w44942, w44943, w44944, w44945, w44946, w44947, w44948, w44949, w44950, w44951, w44952, w44953, w44954, w44955, w44956, w44957, w44958, w44959, w44960, w44961, w44962, w44963, w44964, w44965, w44966, w44967, w44968, w44969, w44970, w44971, w44972, w44973, w44974, w44975, w44976, w44977, w44978, w44979, w44980, w44981, w44982, w44983, w44984, w44985, w44986, w44987, w44988, w44989, w44990, w44991, w44992, w44993, w44994, w44995, w44996, w44997, w44998, w44999, w45000, w45001, w45002, w45003, w45004, w45005, w45006, w45007, w45008, w45009, w45010, w45011, w45012, w45013, w45014, w45015, w45016, w45017, w45018, w45019, w45020, w45021, w45022, w45023, w45024, w45025, w45026, w45027, w45028, w45029, w45030, w45031, w45032, w45033, w45034, w45035, w45036, w45037, w45038, w45039, w45040, w45041, w45042, w45043, w45044, w45045, w45046, w45047, w45048, w45049, w45050, w45051, w45052, w45053, w45054, w45055, w45056, w45057, w45058, w45059, w45060, w45061, w45062, w45063, w45064, w45065, w45066, w45067, w45068, w45069, w45070, w45071, w45072, w45073, w45074, w45075, w45076, w45077, w45078, w45079, w45080, w45081, w45082, w45083, w45084, w45085, w45086, w45087, w45088, w45089, w45090, w45091, w45092, w45093, w45094, w45095, w45096, w45097, w45098, w45099, w45100, w45101, w45102, w45103, w45104, w45105, w45106, w45107, w45108, w45109, w45110, w45111, w45112, w45113, w45114, w45115, w45116, w45117, w45118, w45119, w45120, w45121, w45122, w45123, w45124, w45125, w45126, w45127, w45128, w45129, w45130, w45131, w45132, w45133, w45134, w45135, w45136, w45137, w45138, w45139, w45140, w45141, w45142, w45143, w45144, w45145, w45146, w45147, w45148, w45149, w45150, w45151, w45152, w45153, w45154, w45155, w45156, w45157, w45158, w45159, w45160, w45161, w45162, w45163, w45164, w45165, w45166, w45167, w45168, w45169, w45170, w45171, w45172, w45173, w45174, w45175, w45176, w45177, w45178, w45179, w45180, w45181, w45182, w45183, w45184, w45185, w45186, w45187, w45188, w45189, w45190, w45191, w45192, w45193, w45194, w45195, w45196, w45197, w45198, w45199, w45200, w45201, w45202, w45203, w45204, w45205, w45206, w45207, w45208, w45209, w45210, w45211, w45212, w45213, w45214, w45215, w45216, w45217, w45218, w45219, w45220, w45221, w45222, w45223, w45224, w45225, w45226, w45227, w45228, w45229, w45230, w45231, w45232, w45233, w45234, w45235, w45236, w45237, w45238, w45239, w45240, w45241, w45242, w45243, w45244, w45245, w45246, w45247, w45248, w45249, w45250, w45251, w45252, w45253, w45254, w45255, w45256, w45257, w45258, w45259, w45260, w45261, w45262, w45263, w45264, w45265, w45266, w45267, w45268, w45269, w45270, w45271, w45272, w45273, w45274, w45275, w45276, w45277, w45278, w45279, w45280, w45281, w45282, w45283, w45284, w45285, w45286, w45287, w45288, w45289, w45290, w45291, w45292, w45293, w45294, w45295, w45296, w45297, w45298, w45299, w45300, w45301, w45302, w45303, w45304, w45305, w45306, w45307, w45308, w45309, w45310, w45311, w45312, w45313, w45314, w45315, w45316, w45317, w45318, w45319, w45320, w45321, w45322, w45323, w45324, w45325, w45326, w45327, w45328, w45329, w45330, w45331, w45332, w45333, w45334, w45335, w45336, w45337, w45338, w45339, w45340, w45341, w45342, w45343, w45344, w45345, w45346, w45347, w45348, w45349, w45350, w45351, w45352, w45353, w45354, w45355, w45356, w45357, w45358, w45359, w45360, w45361, w45362, w45363, w45364, w45365, w45366, w45367, w45368, w45369, w45370, w45371, w45372, w45373, w45374, w45375, w45376, w45377, w45378, w45379, w45380, w45381, w45382, w45383, w45384, w45385, w45386, w45387, w45388, w45389, w45390, w45391, w45392, w45393, w45394, w45395, w45396, w45397, w45398, w45399, w45400, w45401, w45402, w45403, w45404, w45405, w45406, w45407, w45408, w45409, w45410, w45411, w45412, w45413, w45414, w45415, w45416, w45417, w45418, w45419, w45420, w45421, w45422, w45423, w45424, w45425, w45426, w45427, w45428, w45429, w45430, w45431, w45432, w45433, w45434, w45435, w45436, w45437, w45438, w45439, w45440, w45441, w45442, w45443, w45444, w45445, w45446, w45447, w45448, w45449, w45450, w45451, w45452, w45453, w45454, w45455, w45456, w45457, w45458, w45459, w45460, w45461, w45462, w45463, w45464, w45465, w45466, w45467, w45468, w45469, w45470, w45471, w45472, w45473, w45474, w45475, w45476, w45477, w45478, w45479, w45480, w45481, w45482, w45483, w45484, w45485, w45486, w45487, w45488, w45489, w45490, w45491, w45492, w45493, w45494, w45495, w45496, w45497, w45498, w45499, w45500, w45501, w45502, w45503, w45504, w45505, w45506, w45507, w45508, w45509, w45510, w45511, w45512, w45513, w45514, w45515, w45516, w45517, w45518, w45519, w45520, w45521, w45522, w45523, w45524, w45525, w45526, w45527, w45528, w45529, w45530, w45531, w45532, w45533, w45534, w45535, w45536, w45537, w45538, w45539, w45540, w45541, w45542, w45543, w45544, w45545, w45546, w45547, w45548, w45549, w45550, w45551, w45552, w45553, w45554, w45555, w45556, w45557, w45558, w45559, w45560, w45561, w45562, w45563, w45564, w45565, w45566, w45567, w45568, w45569, w45570, w45571, w45572, w45573, w45574, w45575, w45576, w45577, w45578, w45579, w45580, w45581, w45582, w45583, w45584, w45585, w45586, w45587, w45588, w45589, w45590, w45591, w45592, w45593, w45594, w45595, w45596, w45597, w45598, w45599, w45600, w45601, w45602, w45603, w45604, w45605, w45606, w45607, w45608, w45609, w45610, w45611, w45612, w45613, w45614, w45615, w45616, w45617, w45618, w45619, w45620, w45621, w45622, w45623, w45624, w45625, w45626, w45627, w45628, w45629, w45630, w45631, w45632, w45633, w45634, w45635, w45636, w45637, w45638, w45639, w45640, w45641, w45642, w45643, w45644, w45645, w45646, w45647, w45648, w45649, w45650, w45651, w45652, w45653, w45654, w45655, w45656, w45657, w45658, w45659, w45660, w45661, w45662, w45663, w45664, w45665, w45666, w45667, w45668, w45669, w45670, w45671, w45672, w45673, w45674, w45675, w45676, w45677, w45678, w45679, w45680, w45681, w45682, w45683, w45684, w45685, w45686, w45687, w45688, w45689, w45690, w45691, w45692, w45693, w45694, w45695, w45696, w45697, w45698, w45699, w45700, w45701, w45702, w45703, w45704, w45705, w45706, w45707, w45708, w45709, w45710, w45711, w45712, w45713, w45714, w45715, w45716, w45717, w45718, w45719, w45720, w45721, w45722, w45723, w45724, w45725, w45726, w45727, w45728, w45729, w45730, w45731, w45732, w45733, w45734, w45735, w45736, w45737, w45738, w45739, w45740, w45741, w45742, w45743, w45744, w45745, w45746, w45747, w45748, w45749, w45750, w45751, w45752, w45753, w45754, w45755, w45756, w45757, w45758, w45759, w45760, w45761, w45762, w45763, w45764, w45765, w45766, w45767, w45768, w45769, w45770, w45771, w45772, w45773, w45774, w45775, w45776, w45777, w45778, w45779, w45780, w45781, w45782, w45783, w45784, w45785, w45786, w45787, w45788, w45789, w45790, w45791, w45792, w45793, w45794, w45795, w45796, w45797, w45798, w45799, w45800, w45801, w45802, w45803, w45804, w45805, w45806, w45807, w45808, w45809, w45810, w45811, w45812, w45813, w45814, w45815, w45816, w45817, w45818, w45819, w45820, w45821, w45822, w45823, w45824, w45825, w45826, w45827, w45828, w45829, w45830, w45831, w45832, w45833, w45834, w45835, w45836, w45837, w45838, w45839, w45840, w45841, w45842, w45843, w45844, w45845, w45846, w45847, w45848, w45849, w45850, w45851, w45852, w45853, w45854, w45855, w45856, w45857, w45858, w45859, w45860, w45861, w45862, w45863, w45864, w45865, w45866, w45867, w45868, w45869, w45870, w45871, w45872, w45873, w45874, w45875, w45876, w45877, w45878, w45879, w45880, w45881, w45882, w45883, w45884, w45885, w45886, w45887, w45888, w45889, w45890, w45891, w45892, w45893, w45894, w45895, w45896, w45897, w45898, w45899, w45900, w45901, w45902, w45903, w45904, w45905, w45906, w45907, w45908, w45909, w45910, w45911, w45912, w45913, w45914, w45915, w45916, w45917, w45918, w45919, w45920, w45921, w45922, w45923, w45924, w45925, w45926, w45927, w45928, w45929, w45930, w45931, w45932, w45933, w45934, w45935, w45936, w45937, w45938, w45939, w45940, w45941, w45942, w45943, w45944, w45945, w45946, w45947, w45948, w45949, w45950, w45951, w45952, w45953, w45954, w45955, w45956, w45957, w45958, w45959, w45960, w45961, w45962, w45963, w45964, w45965, w45966, w45967, w45968, w45969, w45970, w45971, w45972, w45973, w45974, w45975, w45976, w45977, w45978, w45979, w45980, w45981, w45982, w45983, w45984, w45985, w45986, w45987, w45988, w45989, w45990, w45991, w45992, w45993, w45994, w45995, w45996, w45997, w45998, w45999, w46000, w46001, w46002, w46003, w46004, w46005, w46006, w46007, w46008, w46009, w46010, w46011, w46012, w46013, w46014, w46015, w46016, w46017, w46018, w46019, w46020, w46021, w46022, w46023, w46024, w46025, w46026, w46027, w46028, w46029, w46030, w46031, w46032, w46033, w46034, w46035, w46036, w46037, w46038, w46039, w46040, w46041, w46042, w46043, w46044, w46045, w46046, w46047, w46048, w46049, w46050, w46051, w46052, w46053, w46054, w46055, w46056, w46057, w46058, w46059, w46060, w46061, w46062, w46063, w46064, w46065, w46066, w46067, w46068, w46069, w46070, w46071, w46072, w46073, w46074, w46075, w46076, w46077, w46078, w46079, w46080, w46081, w46082, w46083, w46084, w46085, w46086, w46087, w46088, w46089, w46090, w46091, w46092, w46093, w46094, w46095, w46096, w46097, w46098, w46099, w46100, w46101, w46102, w46103, w46104, w46105, w46106, w46107, w46108, w46109, w46110, w46111, w46112, w46113, w46114, w46115, w46116, w46117, w46118, w46119, w46120, w46121, w46122, w46123, w46124, w46125, w46126, w46127, w46128, w46129, w46130, w46131, w46132, w46133, w46134, w46135, w46136, w46137, w46138, w46139, w46140, w46141, w46142, w46143, w46144, w46145, w46146, w46147, w46148, w46149, w46150, w46151, w46152, w46153, w46154, w46155, w46156, w46157, w46158, w46159, w46160, w46161, w46162, w46163, w46164, w46165, w46166, w46167, w46168, w46169, w46170, w46171, w46172, w46173, w46174, w46175, w46176, w46177, w46178, w46179, w46180, w46181, w46182, w46183, w46184, w46185, w46186, w46187, w46188, w46189, w46190, w46191, w46192, w46193, w46194, w46195, w46196, w46197, w46198, w46199, w46200, w46201, w46202, w46203, w46204, w46205, w46206, w46207, w46208, w46209, w46210, w46211, w46212, w46213, w46214, w46215, w46216, w46217, w46218, w46219, w46220, w46221, w46222, w46223, w46224, w46225, w46226, w46227, w46228, w46229, w46230, w46231, w46232, w46233, w46234, w46235, w46236, w46237, w46238, w46239, w46240, w46241, w46242, w46243, w46244, w46245, w46246, w46247, w46248, w46249, w46250, w46251, w46252, w46253, w46254, w46255, w46256, w46257, w46258, w46259, w46260, w46261, w46262, w46263, w46264, w46265, w46266, w46267, w46268, w46269, w46270, w46271, w46272, w46273, w46274, w46275, w46276, w46277, w46278, w46279, w46280, w46281, w46282, w46283, w46284, w46285, w46286, w46287, w46288, w46289, w46290, w46291, w46292, w46293, w46294, w46295, w46296, w46297, w46298, w46299, w46300, w46301, w46302, w46303, w46304, w46305, w46306, w46307, w46308, w46309, w46310, w46311, w46312, w46313, w46314, w46315, w46316, w46317, w46318, w46319, w46320, w46321, w46322, w46323, w46324, w46325, w46326, w46327, w46328, w46329, w46330, w46331, w46332, w46333, w46334, w46335, w46336, w46337, w46338, w46339, w46340, w46341, w46342, w46343, w46344, w46345, w46346, w46347, w46348, w46349, w46350, w46351, w46352, w46353, w46354, w46355, w46356, w46357, w46358, w46359, w46360, w46361, w46362, w46363, w46364, w46365, w46366, w46367, w46368, w46369, w46370, w46371, w46372, w46373, w46374, w46375, w46376, w46377, w46378, w46379, w46380, w46381, w46382, w46383, w46384, w46385, w46386, w46387, w46388, w46389, w46390, w46391, w46392, w46393, w46394, w46395, w46396, w46397, w46398, w46399, w46400, w46401, w46402, w46403, w46404, w46405, w46406, w46407, w46408, w46409, w46410, w46411, w46412, w46413, w46414, w46415, w46416, w46417, w46418, w46419, w46420, w46421, w46422, w46423, w46424, w46425, w46426, w46427, w46428, w46429, w46430, w46431, w46432, w46433, w46434, w46435, w46436, w46437, w46438, w46439, w46440, w46441, w46442, w46443, w46444, w46445, w46446, w46447, w46448, w46449, w46450, w46451, w46452, w46453, w46454, w46455, w46456, w46457, w46458, w46459, w46460, w46461, w46462, w46463, w46464, w46465, w46466, w46467, w46468, w46469, w46470, w46471, w46472, w46473, w46474, w46475, w46476, w46477, w46478, w46479, w46480, w46481, w46482, w46483, w46484, w46485, w46486, w46487, w46488, w46489, w46490, w46491, w46492, w46493, w46494, w46495, w46496, w46497, w46498, w46499, w46500, w46501, w46502, w46503, w46504, w46505, w46506, w46507, w46508, w46509, w46510, w46511, w46512, w46513, w46514, w46515, w46516, w46517, w46518, w46519, w46520, w46521, w46522, w46523, w46524, w46525, w46526, w46527, w46528, w46529, w46530, w46531, w46532, w46533, w46534, w46535, w46536, w46537, w46538, w46539, w46540, w46541, w46542, w46543, w46544, w46545, w46546, w46547, w46548, w46549, w46550, w46551, w46552, w46553, w46554, w46555, w46556, w46557, w46558, w46559, w46560, w46561, w46562, w46563, w46564, w46565, w46566, w46567, w46568, w46569, w46570, w46571, w46572, w46573, w46574, w46575, w46576, w46577, w46578, w46579, w46580, w46581, w46582, w46583, w46584, w46585, w46586, w46587, w46588, w46589, w46590, w46591, w46592, w46593, w46594, w46595, w46596, w46597, w46598, w46599, w46600, w46601, w46602, w46603, w46604, w46605, w46606, w46607, w46608, w46609, w46610, w46611, w46612, w46613, w46614, w46615, w46616, w46617, w46618, w46619, w46620, w46621, w46622, w46623, w46624, w46625, w46626, w46627, w46628, w46629, w46630, w46631, w46632, w46633, w46634, w46635, w46636, w46637, w46638, w46639, w46640, w46641, w46642, w46643, w46644, w46645, w46646, w46647, w46648, w46649, w46650, w46651, w46652, w46653, w46654, w46655, w46656, w46657, w46658, w46659, w46660, w46661, w46662, w46663, w46664, w46665, w46666, w46667, w46668, w46669, w46670, w46671, w46672, w46673, w46674, w46675, w46676, w46677, w46678, w46679, w46680, w46681, w46682, w46683, w46684, w46685, w46686, w46687, w46688, w46689, w46690, w46691, w46692, w46693, w46694, w46695, w46696, w46697, w46698, w46699, w46700, w46701, w46702, w46703, w46704, w46705, w46706, w46707, w46708, w46709, w46710, w46711, w46712, w46713, w46714, w46715, w46716, w46717, w46718, w46719, w46720, w46721, w46722, w46723, w46724, w46725, w46726, w46727, w46728, w46729, w46730, w46731, w46732, w46733, w46734, w46735, w46736, w46737, w46738, w46739, w46740, w46741, w46742, w46743, w46744, w46745, w46746, w46747, w46748, w46749, w46750, w46751, w46752, w46753, w46754, w46755, w46756, w46757, w46758, w46759, w46760, w46761, w46762, w46763, w46764, w46765, w46766, w46767, w46768, w46769, w46770, w46771, w46772, w46773, w46774, w46775, w46776, w46777, w46778, w46779, w46780, w46781, w46782, w46783, w46784, w46785, w46786, w46787, w46788, w46789, w46790, w46791, w46792, w46793, w46794, w46795, w46796, w46797, w46798, w46799, w46800, w46801, w46802, w46803, w46804, w46805, w46806, w46807, w46808, w46809, w46810, w46811, w46812, w46813, w46814, w46815, w46816, w46817, w46818, w46819, w46820, w46821, w46822, w46823, w46824, w46825, w46826, w46827, w46828, w46829, w46830, w46831, w46832, w46833, w46834, w46835, w46836, w46837, w46838, w46839, w46840, w46841, w46842, w46843, w46844, w46845, w46846, w46847, w46848, w46849, w46850, w46851, w46852, w46853, w46854, w46855, w46856, w46857, w46858, w46859, w46860, w46861, w46862, w46863, w46864, w46865, w46866, w46867, w46868, w46869, w46870, w46871, w46872, w46873, w46874, w46875, w46876, w46877, w46878, w46879, w46880, w46881, w46882, w46883, w46884, w46885, w46886, w46887, w46888, w46889, w46890, w46891, w46892, w46893, w46894, w46895, w46896, w46897, w46898, w46899, w46900, w46901, w46902, w46903, w46904, w46905, w46906, w46907, w46908, w46909, w46910, w46911, w46912, w46913, w46914, w46915, w46916, w46917, w46918, w46919, w46920, w46921, w46922, w46923, w46924, w46925, w46926, w46927, w46928, w46929, w46930, w46931, w46932, w46933, w46934, w46935, w46936, w46937, w46938, w46939, w46940, w46941, w46942, w46943, w46944, w46945, w46946, w46947, w46948, w46949, w46950, w46951, w46952, w46953, w46954, w46955, w46956, w46957, w46958, w46959, w46960, w46961, w46962, w46963, w46964, w46965, w46966, w46967, w46968, w46969, w46970, w46971, w46972, w46973, w46974, w46975, w46976, w46977, w46978, w46979, w46980, w46981, w46982, w46983, w46984, w46985, w46986, w46987, w46988, w46989, w46990, w46991, w46992, w46993, w46994, w46995, w46996, w46997, w46998, w46999, w47000, w47001, w47002, w47003, w47004, w47005, w47006, w47007, w47008, w47009, w47010, w47011, w47012, w47013, w47014, w47015, w47016, w47017, w47018, w47019, w47020, w47021, w47022, w47023, w47024, w47025, w47026, w47027, w47028, w47029, w47030, w47031, w47032, w47033, w47034, w47035, w47036, w47037, w47038, w47039, w47040, w47041, w47042, w47043, w47044, w47045, w47046, w47047, w47048, w47049, w47050, w47051, w47052, w47053, w47054, w47055, w47056, w47057, w47058, w47059, w47060, w47061, w47062, w47063, w47064, w47065, w47066, w47067, w47068, w47069, w47070, w47071, w47072, w47073, w47074, w47075, w47076, w47077, w47078, w47079, w47080, w47081, w47082, w47083, w47084, w47085, w47086, w47087, w47088, w47089, w47090, w47091, w47092, w47093, w47094, w47095, w47096, w47097, w47098, w47099, w47100, w47101, w47102, w47103, w47104, w47105, w47106, w47107, w47108, w47109, w47110, w47111, w47112, w47113, w47114, w47115, w47116, w47117, w47118, w47119, w47120, w47121, w47122, w47123, w47124, w47125, w47126, w47127, w47128, w47129, w47130, w47131, w47132, w47133, w47134, w47135, w47136, w47137, w47138, w47139, w47140, w47141, w47142, w47143, w47144, w47145, w47146, w47147, w47148, w47149, w47150, w47151, w47152, w47153, w47154, w47155, w47156, w47157, w47158, w47159, w47160, w47161, w47162, w47163, w47164, w47165, w47166, w47167, w47168, w47169, w47170, w47171, w47172, w47173, w47174, w47175, w47176, w47177, w47178, w47179, w47180, w47181, w47182, w47183, w47184, w47185, w47186, w47187, w47188, w47189, w47190, w47191, w47192, w47193, w47194, w47195, w47196, w47197, w47198, w47199, w47200, w47201, w47202, w47203, w47204, w47205, w47206, w47207, w47208, w47209, w47210, w47211, w47212, w47213, w47214, w47215, w47216, w47217, w47218, w47219, w47220, w47221, w47222, w47223, w47224, w47225, w47226, w47227, w47228, w47229, w47230, w47231, w47232, w47233, w47234, w47235, w47236, w47237, w47238, w47239, w47240, w47241, w47242, w47243, w47244, w47245, w47246, w47247, w47248, w47249, w47250, w47251, w47252, w47253, w47254, w47255, w47256, w47257, w47258, w47259, w47260, w47261, w47262, w47263, w47264, w47265, w47266, w47267, w47268, w47269, w47270, w47271, w47272, w47273, w47274, w47275, w47276, w47277, w47278, w47279, w47280, w47281, w47282, w47283, w47284, w47285, w47286, w47287, w47288, w47289, w47290, w47291, w47292, w47293, w47294, w47295, w47296, w47297, w47298, w47299, w47300, w47301, w47302, w47303, w47304, w47305, w47306, w47307, w47308, w47309, w47310, w47311, w47312, w47313, w47314, w47315, w47316, w47317, w47318, w47319, w47320, w47321, w47322, w47323, w47324, w47325, w47326, w47327, w47328, w47329, w47330, w47331, w47332, w47333, w47334, w47335, w47336, w47337, w47338, w47339, w47340, w47341, w47342, w47343, w47344, w47345, w47346, w47347, w47348, w47349, w47350, w47351, w47352, w47353, w47354, w47355, w47356, w47357, w47358, w47359, w47360, w47361, w47362, w47363, w47364, w47365, w47366, w47367, w47368, w47369, w47370, w47371, w47372, w47373, w47374, w47375, w47376, w47377, w47378, w47379, w47380, w47381, w47382, w47383, w47384, w47385, w47386, w47387, w47388, w47389, w47390, w47391, w47392, w47393, w47394, w47395, w47396, w47397, w47398, w47399, w47400, w47401, w47402, w47403, w47404, w47405, w47406, w47407, w47408, w47409, w47410, w47411, w47412, w47413, w47414, w47415, w47416, w47417, w47418, w47419, w47420, w47421, w47422, w47423, w47424, w47425, w47426, w47427, w47428, w47429, w47430, w47431, w47432, w47433, w47434, w47435, w47436, w47437, w47438, w47439, w47440, w47441, w47442, w47443, w47444, w47445, w47446, w47447, w47448, w47449, w47450, w47451, w47452, w47453, w47454, w47455, w47456, w47457, w47458, w47459, w47460, w47461, w47462, w47463, w47464, w47465, w47466, w47467, w47468, w47469, w47470, w47471, w47472, w47473, w47474, w47475, w47476, w47477, w47478, w47479, w47480, w47481, w47482, w47483, w47484, w47485, w47486, w47487, w47488, w47489, w47490, w47491, w47492, w47493, w47494, w47495, w47496, w47497, w47498, w47499, w47500, w47501, w47502, w47503, w47504, w47505, w47506, w47507, w47508, w47509, w47510, w47511, w47512, w47513, w47514, w47515, w47516, w47517, w47518, w47519, w47520, w47521, w47522, w47523, w47524, w47525, w47526, w47527, w47528, w47529, w47530, w47531, w47532, w47533, w47534, w47535, w47536, w47537, w47538, w47539, w47540, w47541, w47542, w47543, w47544, w47545, w47546, w47547, w47548, w47549, w47550, w47551, w47552, w47553, w47554, w47555, w47556, w47557, w47558, w47559, w47560, w47561, w47562, w47563, w47564, w47565, w47566, w47567, w47568, w47569, w47570, w47571, w47572, w47573, w47574, w47575, w47576, w47577, w47578, w47579, w47580, w47581, w47582, w47583, w47584, w47585, w47586, w47587, w47588, w47589, w47590, w47591, w47592, w47593, w47594, w47595, w47596, w47597, w47598, w47599, w47600, w47601, w47602, w47603, w47604, w47605, w47606, w47607, w47608, w47609, w47610, w47611, w47612, w47613, w47614, w47615, w47616, w47617, w47618, w47619, w47620, w47621, w47622, w47623, w47624, w47625, w47626, w47627, w47628, w47629, w47630, w47631, w47632, w47633, w47634, w47635, w47636, w47637, w47638, w47639, w47640, w47641, w47642, w47643, w47644, w47645, w47646, w47647, w47648, w47649, w47650, w47651, w47652, w47653, w47654, w47655, w47656, w47657, w47658, w47659, w47660, w47661, w47662, w47663, w47664, w47665, w47666, w47667, w47668, w47669, w47670, w47671, w47672, w47673, w47674, w47675, w47676, w47677, w47678, w47679, w47680, w47681, w47682, w47683, w47684, w47685, w47686, w47687, w47688, w47689, w47690, w47691, w47692, w47693, w47694, w47695, w47696, w47697, w47698, w47699, w47700, w47701, w47702, w47703, w47704, w47705, w47706, w47707, w47708, w47709, w47710, w47711, w47712, w47713, w47714, w47715, w47716, w47717, w47718, w47719, w47720, w47721, w47722, w47723, w47724, w47725, w47726, w47727, w47728, w47729, w47730, w47731, w47732, w47733, w47734, w47735, w47736, w47737, w47738, w47739, w47740, w47741, w47742, w47743, w47744, w47745, w47746, w47747, w47748, w47749, w47750, w47751, w47752, w47753, w47754, w47755, w47756, w47757, w47758, w47759, w47760, w47761, w47762, w47763, w47764, w47765, w47766, w47767, w47768, w47769, w47770, w47771, w47772, w47773, w47774, w47775, w47776, w47777, w47778, w47779, w47780, w47781, w47782, w47783, w47784, w47785, w47786, w47787, w47788, w47789, w47790, w47791, w47792, w47793, w47794, w47795, w47796, w47797, w47798, w47799, w47800, w47801, w47802, w47803, w47804, w47805, w47806, w47807, w47808, w47809, w47810, w47811, w47812, w47813, w47814, w47815, w47816, w47817, w47818, w47819, w47820, w47821, w47822, w47823, w47824, w47825, w47826, w47827, w47828, w47829, w47830, w47831, w47832, w47833, w47834, w47835, w47836, w47837, w47838, w47839, w47840, w47841, w47842, w47843, w47844, w47845, w47846, w47847, w47848, w47849, w47850, w47851, w47852, w47853, w47854, w47855, w47856, w47857, w47858, w47859, w47860, w47861, w47862, w47863, w47864, w47865, w47866, w47867, w47868, w47869, w47870, w47871, w47872, w47873, w47874, w47875, w47876, w47877, w47878, w47879, w47880, w47881, w47882, w47883, w47884, w47885, w47886, w47887, w47888, w47889, w47890, w47891, w47892, w47893, w47894, w47895, w47896, w47897, w47898, w47899, w47900, w47901, w47902, w47903, w47904, w47905, w47906, w47907, w47908, w47909, w47910, w47911, w47912, w47913, w47914, w47915, w47916, w47917, w47918, w47919, w47920, w47921, w47922, w47923, w47924, w47925, w47926, w47927, w47928, w47929, w47930, w47931, w47932, w47933, w47934, w47935, w47936, w47937, w47938, w47939, w47940, w47941, w47942, w47943, w47944, w47945, w47946, w47947, w47948, w47949, w47950, w47951, w47952, w47953, w47954, w47955, w47956, w47957, w47958, w47959, w47960, w47961, w47962, w47963, w47964, w47965, w47966, w47967, w47968, w47969, w47970, w47971, w47972, w47973, w47974, w47975, w47976, w47977, w47978, w47979, w47980, w47981, w47982, w47983, w47984, w47985, w47986, w47987, w47988, w47989, w47990, w47991, w47992, w47993, w47994, w47995, w47996, w47997, w47998, w47999, w48000, w48001, w48002, w48003, w48004, w48005, w48006, w48007, w48008, w48009, w48010, w48011, w48012, w48013, w48014, w48015, w48016, w48017, w48018, w48019, w48020, w48021, w48022, w48023, w48024, w48025, w48026, w48027, w48028, w48029, w48030, w48031, w48032, w48033, w48034, w48035, w48036, w48037, w48038, w48039, w48040, w48041, w48042, w48043, w48044, w48045, w48046, w48047, w48048, w48049, w48050, w48051, w48052, w48053, w48054, w48055, w48056, w48057, w48058, w48059, w48060, w48061, w48062, w48063, w48064, w48065, w48066, w48067, w48068, w48069, w48070, w48071, w48072, w48073, w48074, w48075, w48076, w48077, w48078, w48079, w48080, w48081, w48082, w48083, w48084, w48085, w48086, w48087, w48088, w48089, w48090, w48091, w48092, w48093, w48094, w48095, w48096, w48097, w48098, w48099, w48100, w48101, w48102, w48103, w48104, w48105, w48106, w48107, w48108, w48109, w48110, w48111, w48112, w48113, w48114, w48115, w48116, w48117, w48118, w48119, w48120, w48121, w48122, w48123, w48124, w48125, w48126, w48127, w48128, w48129, w48130, w48131, w48132, w48133, w48134, w48135, w48136, w48137, w48138, w48139, w48140, w48141, w48142, w48143, w48144, w48145, w48146, w48147, w48148, w48149, w48150, w48151, w48152, w48153, w48154, w48155, w48156, w48157, w48158, w48159, w48160, w48161, w48162, w48163, w48164, w48165, w48166, w48167, w48168, w48169, w48170, w48171, w48172, w48173, w48174, w48175, w48176, w48177, w48178, w48179, w48180, w48181, w48182, w48183, w48184, w48185, w48186, w48187, w48188, w48189, w48190, w48191, w48192, w48193, w48194, w48195, w48196, w48197, w48198, w48199, w48200, w48201, w48202, w48203, w48204, w48205, w48206, w48207, w48208, w48209, w48210, w48211, w48212, w48213, w48214, w48215, w48216, w48217, w48218, w48219, w48220, w48221, w48222, w48223, w48224, w48225, w48226, w48227, w48228, w48229, w48230, w48231, w48232, w48233, w48234, w48235, w48236, w48237, w48238, w48239, w48240, w48241, w48242, w48243, w48244, w48245, w48246, w48247, w48248, w48249, w48250, w48251, w48252, w48253, w48254, w48255, w48256, w48257, w48258, w48259, w48260, w48261, w48262, w48263, w48264, w48265, w48266, w48267, w48268, w48269, w48270, w48271, w48272, w48273, w48274, w48275, w48276, w48277, w48278, w48279, w48280, w48281, w48282, w48283, w48284, w48285, w48286, w48287, w48288, w48289, w48290, w48291, w48292, w48293, w48294, w48295, w48296, w48297, w48298, w48299, w48300, w48301, w48302, w48303, w48304, w48305, w48306, w48307, w48308, w48309, w48310, w48311, w48312, w48313, w48314, w48315, w48316, w48317, w48318, w48319, w48320, w48321, w48322, w48323, w48324, w48325, w48326, w48327, w48328, w48329, w48330, w48331, w48332, w48333, w48334, w48335, w48336, w48337, w48338, w48339, w48340, w48341, w48342, w48343, w48344, w48345, w48346, w48347, w48348, w48349, w48350, w48351, w48352, w48353, w48354, w48355, w48356, w48357, w48358, w48359, w48360, w48361, w48362, w48363, w48364, w48365, w48366, w48367, w48368, w48369, w48370, w48371, w48372, w48373, w48374, w48375, w48376, w48377, w48378, w48379, w48380, w48381, w48382, w48383, w48384, w48385, w48386, w48387, w48388, w48389, w48390, w48391, w48392, w48393, w48394, w48395, w48396, w48397, w48398, w48399, w48400, w48401, w48402, w48403, w48404, w48405, w48406, w48407, w48408, w48409, w48410, w48411, w48412, w48413, w48414, w48415, w48416, w48417, w48418, w48419, w48420, w48421, w48422, w48423, w48424, w48425, w48426, w48427, w48428, w48429, w48430, w48431, w48432, w48433, w48434, w48435, w48436, w48437, w48438, w48439, w48440, w48441, w48442, w48443, w48444, w48445, w48446, w48447, w48448, w48449, w48450, w48451, w48452, w48453, w48454, w48455, w48456, w48457, w48458, w48459, w48460, w48461, w48462, w48463, w48464, w48465, w48466, w48467, w48468, w48469, w48470, w48471, w48472, w48473, w48474, w48475, w48476, w48477, w48478, w48479, w48480, w48481, w48482, w48483, w48484, w48485, w48486, w48487, w48488, w48489, w48490, w48491, w48492, w48493, w48494, w48495, w48496, w48497, w48498, w48499, w48500, w48501, w48502, w48503, w48504, w48505, w48506, w48507, w48508, w48509, w48510, w48511, w48512, w48513, w48514, w48515, w48516, w48517, w48518, w48519, w48520, w48521, w48522, w48523, w48524, w48525, w48526, w48527, w48528, w48529, w48530, w48531, w48532, w48533, w48534, w48535, w48536, w48537, w48538, w48539, w48540, w48541, w48542, w48543, w48544, w48545, w48546, w48547, w48548, w48549, w48550, w48551, w48552, w48553, w48554, w48555, w48556, w48557, w48558, w48559, w48560, w48561, w48562, w48563, w48564, w48565, w48566, w48567, w48568, w48569, w48570, w48571, w48572, w48573, w48574, w48575, w48576, w48577, w48578, w48579, w48580, w48581, w48582, w48583, w48584, w48585, w48586, w48587, w48588, w48589, w48590, w48591, w48592, w48593, w48594, w48595, w48596, w48597, w48598, w48599, w48600, w48601, w48602, w48603, w48604, w48605, w48606, w48607, w48608, w48609, w48610, w48611, w48612, w48613, w48614, w48615, w48616, w48617, w48618, w48619, w48620, w48621, w48622, w48623, w48624, w48625, w48626, w48627, w48628, w48629, w48630, w48631, w48632, w48633, w48634, w48635, w48636, w48637, w48638, w48639, w48640, w48641, w48642, w48643, w48644, w48645, w48646, w48647, w48648, w48649, w48650, w48651, w48652, w48653, w48654, w48655, w48656, w48657, w48658, w48659, w48660, w48661, w48662, w48663, w48664, w48665, w48666, w48667, w48668, w48669, w48670, w48671, w48672, w48673, w48674, w48675, w48676, w48677, w48678, w48679, w48680, w48681, w48682, w48683, w48684, w48685, w48686, w48687, w48688, w48689, w48690, w48691, w48692, w48693, w48694, w48695, w48696, w48697, w48698, w48699, w48700, w48701, w48702, w48703, w48704, w48705, w48706, w48707, w48708, w48709, w48710, w48711, w48712, w48713, w48714, w48715, w48716, w48717, w48718, w48719, w48720, w48721, w48722, w48723, w48724, w48725, w48726, w48727, w48728, w48729, w48730, w48731, w48732, w48733, w48734, w48735, w48736, w48737, w48738, w48739, w48740, w48741, w48742, w48743, w48744, w48745, w48746, w48747, w48748, w48749, w48750, w48751, w48752, w48753, w48754, w48755, w48756, w48757, w48758, w48759, w48760, w48761, w48762, w48763, w48764, w48765, w48766, w48767, w48768, w48769, w48770, w48771, w48772, w48773, w48774, w48775, w48776, w48777, w48778, w48779, w48780, w48781, w48782, w48783, w48784, w48785, w48786, w48787, w48788, w48789, w48790, w48791, w48792, w48793, w48794, w48795, w48796, w48797, w48798, w48799, w48800, w48801, w48802, w48803, w48804, w48805, w48806, w48807, w48808, w48809, w48810, w48811, w48812, w48813, w48814, w48815, w48816, w48817, w48818, w48819, w48820, w48821, w48822, w48823, w48824, w48825, w48826, w48827, w48828, w48829, w48830, w48831, w48832, w48833, w48834, w48835, w48836, w48837, w48838, w48839, w48840, w48841, w48842, w48843, w48844, w48845, w48846, w48847, w48848, w48849, w48850, w48851, w48852, w48853, w48854, w48855, w48856, w48857, w48858, w48859, w48860, w48861, w48862, w48863, w48864, w48865, w48866, w48867, w48868, w48869, w48870, w48871, w48872, w48873, w48874, w48875, w48876, w48877, w48878, w48879, w48880, w48881, w48882, w48883, w48884, w48885, w48886, w48887, w48888, w48889, w48890, w48891, w48892, w48893, w48894, w48895, w48896, w48897, w48898, w48899, w48900, w48901, w48902, w48903, w48904, w48905, w48906, w48907, w48908, w48909, w48910, w48911, w48912, w48913, w48914, w48915, w48916, w48917, w48918, w48919, w48920, w48921, w48922, w48923, w48924, w48925, w48926, w48927, w48928, w48929, w48930, w48931, w48932, w48933, w48934, w48935, w48936, w48937, w48938, w48939, w48940, w48941, w48942, w48943, w48944, w48945, w48946, w48947, w48948, w48949, w48950, w48951, w48952, w48953, w48954, w48955, w48956, w48957, w48958, w48959, w48960, w48961, w48962, w48963, w48964, w48965, w48966, w48967, w48968, w48969, w48970, w48971, w48972, w48973, w48974, w48975, w48976, w48977, w48978, w48979, w48980, w48981, w48982, w48983, w48984, w48985, w48986, w48987, w48988, w48989, w48990, w48991, w48992, w48993, w48994, w48995, w48996, w48997, w48998, w48999, w49000, w49001, w49002, w49003, w49004, w49005, w49006, w49007, w49008, w49009, w49010, w49011, w49012, w49013, w49014, w49015, w49016, w49017, w49018, w49019, w49020, w49021, w49022, w49023, w49024, w49025, w49026, w49027, w49028, w49029, w49030, w49031, w49032, w49033, w49034, w49035, w49036, w49037, w49038, w49039, w49040, w49041, w49042, w49043, w49044, w49045, w49046, w49047, w49048, w49049, w49050, w49051, w49052, w49053, w49054, w49055, w49056, w49057, w49058, w49059, w49060, w49061, w49062, w49063, w49064, w49065, w49066, w49067, w49068, w49069, w49070, w49071, w49072, w49073, w49074, w49075, w49076, w49077, w49078, w49079, w49080, w49081, w49082, w49083, w49084, w49085, w49086, w49087, w49088, w49089, w49090, w49091, w49092, w49093, w49094, w49095, w49096, w49097, w49098, w49099, w49100, w49101, w49102, w49103, w49104, w49105, w49106, w49107, w49108, w49109, w49110, w49111, w49112, w49113, w49114, w49115, w49116, w49117, w49118, w49119, w49120, w49121, w49122, w49123, w49124, w49125, w49126, w49127, w49128, w49129, w49130, w49131, w49132, w49133, w49134, w49135, w49136, w49137, w49138, w49139, w49140, w49141, w49142, w49143, w49144, w49145, w49146, w49147, w49148, w49149, w49150, w49151, w49152, w49153, w49154, w49155, w49156, w49157, w49158, w49159, w49160, w49161, w49162, w49163, w49164, w49165, w49166, w49167, w49168, w49169, w49170, w49171, w49172, w49173, w49174, w49175, w49176, w49177, w49178, w49179, w49180, w49181, w49182, w49183, w49184, w49185, w49186, w49187, w49188, w49189, w49190, w49191, w49192, w49193, w49194, w49195, w49196, w49197, w49198, w49199, w49200, w49201, w49202, w49203, w49204, w49205, w49206, w49207, w49208, w49209, w49210, w49211, w49212, w49213, w49214, w49215, w49216, w49217, w49218, w49219, w49220, w49221, w49222, w49223, w49224, w49225, w49226, w49227, w49228, w49229, w49230, w49231, w49232, w49233, w49234, w49235, w49236, w49237, w49238, w49239, w49240, w49241, w49242, w49243, w49244, w49245, w49246, w49247, w49248, w49249, w49250, w49251, w49252, w49253, w49254, w49255, w49256, w49257, w49258, w49259, w49260, w49261, w49262, w49263, w49264, w49265, w49266, w49267, w49268, w49269, w49270, w49271, w49272, w49273, w49274, w49275, w49276, w49277, w49278, w49279, w49280, w49281, w49282, w49283, w49284, w49285, w49286, w49287, w49288, w49289, w49290, w49291, w49292, w49293, w49294, w49295, w49296, w49297, w49298, w49299, w49300, w49301, w49302, w49303, w49304, w49305, w49306, w49307, w49308, w49309, w49310, w49311, w49312, w49313, w49314, w49315, w49316, w49317, w49318, w49319, w49320, w49321, w49322, w49323, w49324, w49325, w49326, w49327, w49328, w49329, w49330, w49331, w49332, w49333, w49334, w49335, w49336, w49337, w49338, w49339, w49340, w49341, w49342, w49343, w49344, w49345, w49346, w49347, w49348, w49349, w49350, w49351, w49352, w49353, w49354, w49355, w49356, w49357, w49358, w49359, w49360, w49361, w49362, w49363, w49364, w49365, w49366, w49367, w49368, w49369, w49370, w49371, w49372, w49373, w49374, w49375, w49376, w49377, w49378, w49379, w49380, w49381, w49382, w49383, w49384, w49385, w49386, w49387, w49388, w49389, w49390, w49391, w49392, w49393, w49394, w49395, w49396, w49397, w49398, w49399, w49400, w49401, w49402, w49403, w49404, w49405, w49406, w49407, w49408, w49409, w49410, w49411, w49412, w49413, w49414, w49415, w49416, w49417, w49418, w49419, w49420, w49421, w49422, w49423, w49424, w49425, w49426, w49427, w49428, w49429, w49430, w49431, w49432, w49433, w49434, w49435, w49436, w49437, w49438, w49439, w49440, w49441, w49442, w49443, w49444, w49445, w49446, w49447, w49448, w49449, w49450, w49451, w49452, w49453, w49454, w49455, w49456, w49457, w49458, w49459, w49460, w49461, w49462, w49463, w49464, w49465, w49466, w49467, w49468, w49469, w49470, w49471, w49472, w49473, w49474, w49475, w49476, w49477, w49478, w49479, w49480, w49481, w49482, w49483, w49484, w49485, w49486, w49487, w49488, w49489, w49490, w49491, w49492, w49493, w49494, w49495, w49496, w49497, w49498, w49499, w49500, w49501, w49502, w49503, w49504, w49505, w49506, w49507, w49508, w49509, w49510, w49511, w49512, w49513, w49514, w49515, w49516, w49517, w49518, w49519, w49520, w49521, w49522, w49523, w49524, w49525, w49526, w49527, w49528, w49529, w49530, w49531, w49532, w49533, w49534, w49535, w49536, w49537, w49538, w49539, w49540, w49541, w49542, w49543, w49544, w49545, w49546, w49547, w49548, w49549, w49550, w49551, w49552, w49553, w49554, w49555, w49556, w49557, w49558, w49559, w49560, w49561, w49562, w49563, w49564, w49565, w49566, w49567, w49568, w49569, w49570, w49571, w49572, w49573, w49574, w49575, w49576, w49577, w49578, w49579, w49580, w49581, w49582, w49583, w49584, w49585, w49586, w49587, w49588, w49589, w49590, w49591, w49592, w49593, w49594, w49595, w49596, w49597, w49598, w49599, w49600, w49601, w49602, w49603, w49604, w49605, w49606, w49607, w49608, w49609, w49610, w49611, w49612, w49613, w49614, w49615, w49616, w49617, w49618, w49619, w49620, w49621, w49622, w49623, w49624, w49625, w49626, w49627, w49628, w49629, w49630, w49631, w49632, w49633, w49634, w49635, w49636, w49637, w49638, w49639, w49640, w49641, w49642, w49643, w49644, w49645, w49646, w49647, w49648, w49649, w49650, w49651, w49652, w49653, w49654, w49655, w49656, w49657, w49658, w49659, w49660, w49661, w49662, w49663, w49664, w49665, w49666, w49667, w49668, w49669, w49670, w49671, w49672, w49673, w49674, w49675, w49676, w49677, w49678, w49679, w49680, w49681, w49682, w49683, w49684, w49685, w49686, w49687, w49688, w49689, w49690, w49691, w49692, w49693, w49694, w49695, w49696, w49697, w49698, w49699, w49700, w49701, w49702, w49703, w49704, w49705, w49706, w49707, w49708, w49709, w49710, w49711, w49712, w49713, w49714, w49715, w49716, w49717, w49718, w49719, w49720, w49721, w49722, w49723, w49724, w49725, w49726, w49727, w49728, w49729, w49730, w49731, w49732, w49733, w49734, w49735, w49736, w49737, w49738, w49739, w49740, w49741, w49742, w49743, w49744, w49745, w49746, w49747, w49748, w49749, w49750, w49751, w49752, w49753, w49754, w49755, w49756, w49757, w49758, w49759, w49760, w49761, w49762, w49763, w49764, w49765, w49766, w49767, w49768, w49769, w49770, w49771, w49772, w49773, w49774, w49775, w49776, w49777, w49778, w49779, w49780, w49781, w49782, w49783, w49784, w49785, w49786, w49787, w49788, w49789, w49790, w49791, w49792, w49793, w49794, w49795, w49796, w49797, w49798, w49799, w49800, w49801, w49802, w49803, w49804, w49805, w49806, w49807, w49808, w49809, w49810, w49811, w49812, w49813, w49814, w49815, w49816, w49817, w49818, w49819, w49820, w49821, w49822, w49823, w49824, w49825, w49826, w49827, w49828, w49829, w49830, w49831, w49832, w49833, w49834, w49835, w49836, w49837, w49838, w49839, w49840, w49841, w49842, w49843, w49844, w49845, w49846, w49847, w49848, w49849, w49850, w49851, w49852, w49853, w49854, w49855, w49856, w49857, w49858, w49859, w49860, w49861, w49862, w49863, w49864, w49865, w49866, w49867, w49868, w49869, w49870, w49871, w49872, w49873, w49874, w49875, w49876, w49877, w49878, w49879, w49880, w49881, w49882, w49883, w49884, w49885, w49886, w49887, w49888, w49889, w49890, w49891, w49892, w49893, w49894, w49895, w49896, w49897, w49898, w49899, w49900, w49901, w49902, w49903, w49904, w49905, w49906, w49907, w49908, w49909, w49910, w49911, w49912, w49913, w49914, w49915, w49916, w49917, w49918, w49919, w49920, w49921, w49922, w49923, w49924, w49925, w49926, w49927, w49928, w49929, w49930, w49931, w49932, w49933, w49934, w49935, w49936, w49937, w49938, w49939, w49940, w49941, w49942, w49943, w49944, w49945, w49946, w49947, w49948, w49949, w49950, w49951, w49952, w49953, w49954, w49955, w49956, w49957, w49958, w49959, w49960, w49961, w49962, w49963, w49964, w49965, w49966, w49967, w49968, w49969, w49970, w49971, w49972, w49973, w49974, w49975, w49976, w49977, w49978, w49979, w49980, w49981, w49982, w49983, w49984, w49985, w49986, w49987, w49988, w49989, w49990, w49991, w49992, w49993, w49994, w49995, w49996, w49997, w49998, w49999, w50000, w50001, w50002, w50003, w50004, w50005, w50006, w50007, w50008, w50009, w50010, w50011, w50012, w50013, w50014, w50015, w50016, w50017, w50018, w50019, w50020, w50021, w50022, w50023, w50024, w50025, w50026, w50027, w50028, w50029, w50030, w50031, w50032, w50033, w50034, w50035, w50036, w50037, w50038, w50039, w50040, w50041, w50042, w50043, w50044, w50045, w50046, w50047, w50048, w50049, w50050, w50051, w50052, w50053, w50054, w50055, w50056, w50057, w50058, w50059, w50060, w50061, w50062, w50063, w50064, w50065, w50066, w50067, w50068, w50069, w50070, w50071, w50072, w50073, w50074, w50075, w50076, w50077, w50078, w50079, w50080, w50081, w50082, w50083, w50084, w50085, w50086, w50087, w50088, w50089, w50090, w50091, w50092, w50093, w50094, w50095, w50096, w50097, w50098, w50099, w50100, w50101, w50102, w50103, w50104, w50105, w50106, w50107, w50108, w50109, w50110, w50111, w50112, w50113, w50114, w50115, w50116, w50117, w50118, w50119, w50120, w50121, w50122, w50123, w50124, w50125, w50126, w50127, w50128, w50129, w50130, w50131, w50132, w50133, w50134, w50135, w50136, w50137, w50138, w50139, w50140, w50141, w50142, w50143, w50144, w50145, w50146, w50147, w50148, w50149, w50150, w50151, w50152, w50153, w50154, w50155, w50156, w50157, w50158, w50159, w50160, w50161, w50162, w50163, w50164, w50165, w50166, w50167, w50168, w50169, w50170, w50171, w50172, w50173, w50174, w50175, w50176, w50177, w50178, w50179, w50180, w50181, w50182, w50183, w50184, w50185, w50186, w50187, w50188, w50189, w50190, w50191, w50192, w50193, w50194, w50195, w50196, w50197, w50198, w50199, w50200, w50201, w50202, w50203, w50204, w50205, w50206, w50207, w50208, w50209, w50210, w50211, w50212, w50213, w50214, w50215, w50216, w50217, w50218, w50219, w50220, w50221, w50222, w50223, w50224, w50225, w50226, w50227, w50228, w50229, w50230, w50231, w50232, w50233, w50234, w50235, w50236, w50237, w50238, w50239, w50240, w50241, w50242, w50243, w50244, w50245, w50246, w50247, w50248, w50249, w50250, w50251, w50252, w50253, w50254, w50255, w50256, w50257, w50258, w50259, w50260, w50261, w50262, w50263, w50264, w50265, w50266, w50267, w50268, w50269, w50270, w50271, w50272, w50273, w50274, w50275, w50276, w50277, w50278, w50279, w50280, w50281, w50282, w50283, w50284, w50285, w50286, w50287, w50288, w50289, w50290, w50291, w50292, w50293, w50294, w50295, w50296, w50297, w50298, w50299, w50300, w50301, w50302, w50303, w50304, w50305, w50306, w50307, w50308, w50309, w50310, w50311, w50312, w50313, w50314, w50315, w50316, w50317, w50318, w50319, w50320, w50321, w50322, w50323, w50324, w50325, w50326, w50327, w50328, w50329, w50330, w50331, w50332, w50333, w50334, w50335, w50336, w50337, w50338, w50339, w50340, w50341, w50342, w50343, w50344, w50345, w50346, w50347, w50348, w50349, w50350, w50351, w50352, w50353, w50354, w50355, w50356, w50357, w50358, w50359, w50360, w50361, w50362, w50363, w50364, w50365, w50366, w50367, w50368, w50369, w50370, w50371, w50372, w50373, w50374, w50375, w50376, w50377, w50378, w50379, w50380, w50381, w50382, w50383, w50384, w50385, w50386, w50387, w50388, w50389, w50390, w50391, w50392, w50393, w50394, w50395, w50396, w50397, w50398, w50399, w50400, w50401, w50402, w50403, w50404, w50405, w50406, w50407, w50408, w50409, w50410, w50411, w50412, w50413, w50414, w50415, w50416, w50417, w50418, w50419, w50420, w50421, w50422, w50423, w50424, w50425, w50426, w50427, w50428, w50429, w50430, w50431, w50432, w50433, w50434, w50435, w50436, w50437, w50438, w50439, w50440, w50441, w50442, w50443, w50444, w50445, w50446, w50447, w50448, w50449, w50450, w50451, w50452, w50453, w50454, w50455, w50456, w50457, w50458, w50459, w50460, w50461, w50462, w50463, w50464, w50465, w50466, w50467, w50468, w50469, w50470, w50471, w50472, w50473, w50474, w50475, w50476, w50477, w50478, w50479, w50480, w50481, w50482, w50483, w50484, w50485, w50486, w50487, w50488, w50489, w50490, w50491, w50492, w50493, w50494, w50495, w50496, w50497, w50498, w50499, w50500, w50501, w50502, w50503, w50504, w50505, w50506, w50507, w50508, w50509, w50510, w50511, w50512, w50513, w50514, w50515, w50516, w50517, w50518, w50519, w50520, w50521, w50522, w50523, w50524, w50525, w50526, w50527, w50528, w50529, w50530, w50531, w50532, w50533, w50534, w50535, w50536, w50537, w50538, w50539, w50540, w50541, w50542, w50543, w50544, w50545, w50546, w50547, w50548, w50549, w50550, w50551, w50552, w50553, w50554, w50555, w50556, w50557, w50558, w50559, w50560, w50561, w50562, w50563, w50564, w50565, w50566, w50567, w50568, w50569, w50570, w50571, w50572, w50573, w50574, w50575, w50576, w50577, w50578, w50579, w50580, w50581, w50582, w50583, w50584, w50585, w50586, w50587, w50588, w50589, w50590, w50591, w50592, w50593, w50594, w50595, w50596, w50597, w50598, w50599, w50600, w50601, w50602, w50603, w50604, w50605, w50606, w50607, w50608, w50609, w50610, w50611, w50612, w50613, w50614, w50615, w50616, w50617, w50618, w50619, w50620, w50621, w50622, w50623, w50624, w50625, w50626, w50627, w50628, w50629, w50630, w50631, w50632, w50633, w50634, w50635, w50636, w50637, w50638, w50639, w50640, w50641, w50642, w50643, w50644, w50645, w50646, w50647, w50648, w50649, w50650, w50651, w50652, w50653, w50654, w50655, w50656, w50657, w50658, w50659, w50660, w50661, w50662, w50663, w50664, w50665, w50666, w50667, w50668, w50669, w50670, w50671, w50672, w50673, w50674, w50675, w50676, w50677, w50678, w50679, w50680, w50681, w50682, w50683, w50684, w50685, w50686, w50687, w50688, w50689, w50690, w50691, w50692, w50693, w50694, w50695, w50696, w50697, w50698, w50699, w50700, w50701, w50702, w50703, w50704, w50705, w50706, w50707, w50708, w50709, w50710, w50711, w50712, w50713, w50714, w50715, w50716, w50717, w50718, w50719, w50720, w50721, w50722, w50723, w50724, w50725, w50726, w50727, w50728, w50729, w50730, w50731, w50732, w50733, w50734, w50735, w50736, w50737, w50738, w50739, w50740, w50741, w50742, w50743, w50744, w50745, w50746, w50747, w50748, w50749, w50750, w50751, w50752, w50753, w50754, w50755, w50756, w50757, w50758, w50759, w50760, w50761, w50762, w50763, w50764, w50765, w50766, w50767, w50768, w50769, w50770, w50771, w50772, w50773, w50774, w50775, w50776, w50777, w50778, w50779, w50780, w50781, w50782, w50783, w50784, w50785, w50786, w50787, w50788, w50789, w50790, w50791, w50792, w50793, w50794, w50795, w50796, w50797, w50798, w50799, w50800, w50801, w50802, w50803, w50804, w50805, w50806, w50807, w50808, w50809, w50810, w50811, w50812, w50813, w50814, w50815, w50816, w50817, w50818, w50819, w50820, w50821, w50822, w50823, w50824, w50825, w50826, w50827, w50828, w50829, w50830, w50831, w50832, w50833, w50834, w50835, w50836, w50837, w50838, w50839, w50840, w50841, w50842, w50843, w50844, w50845, w50846, w50847, w50848, w50849, w50850, w50851, w50852, w50853, w50854, w50855, w50856, w50857, w50858, w50859, w50860, w50861, w50862, w50863, w50864, w50865, w50866, w50867, w50868, w50869, w50870, w50871, w50872, w50873, w50874, w50875, w50876, w50877, w50878, w50879, w50880, w50881, w50882, w50883, w50884, w50885, w50886, w50887, w50888, w50889, w50890, w50891, w50892, w50893, w50894, w50895, w50896, w50897, w50898, w50899, w50900, w50901, w50902, w50903, w50904, w50905, w50906, w50907, w50908, w50909, w50910, w50911, w50912, w50913, w50914, w50915, w50916, w50917, w50918, w50919, w50920, w50921, w50922, w50923, w50924, w50925, w50926, w50927, w50928, w50929, w50930, w50931, w50932, w50933, w50934, w50935, w50936, w50937, w50938, w50939, w50940, w50941, w50942, w50943, w50944, w50945, w50946, w50947, w50948, w50949, w50950, w50951, w50952, w50953, w50954, w50955, w50956, w50957, w50958, w50959, w50960, w50961, w50962, w50963, w50964, w50965, w50966, w50967, w50968, w50969, w50970, w50971, w50972, w50973, w50974, w50975, w50976, w50977, w50978, w50979, w50980, w50981, w50982, w50983, w50984, w50985, w50986, w50987, w50988, w50989, w50990, w50991, w50992, w50993, w50994, w50995, w50996, w50997, w50998, w50999, w51000, w51001, w51002, w51003, w51004, w51005, w51006, w51007, w51008, w51009, w51010, w51011, w51012, w51013, w51014, w51015, w51016, w51017, w51018, w51019, w51020, w51021, w51022, w51023, w51024, w51025, w51026, w51027, w51028, w51029, w51030, w51031, w51032, w51033, w51034, w51035, w51036, w51037, w51038, w51039, w51040, w51041, w51042, w51043, w51044, w51045, w51046, w51047, w51048, w51049, w51050, w51051, w51052, w51053, w51054, w51055, w51056, w51057, w51058, w51059, w51060, w51061, w51062, w51063, w51064, w51065, w51066, w51067, w51068, w51069, w51070, w51071, w51072, w51073, w51074, w51075, w51076, w51077, w51078, w51079, w51080, w51081, w51082, w51083, w51084, w51085, w51086, w51087, w51088, w51089, w51090, w51091, w51092, w51093, w51094, w51095, w51096, w51097, w51098, w51099, w51100, w51101, w51102, w51103, w51104, w51105, w51106, w51107, w51108, w51109, w51110, w51111, w51112, w51113, w51114, w51115, w51116, w51117, w51118, w51119, w51120, w51121, w51122, w51123, w51124, w51125, w51126, w51127, w51128, w51129, w51130, w51131, w51132, w51133, w51134, w51135, w51136, w51137, w51138, w51139, w51140, w51141, w51142, w51143, w51144, w51145, w51146, w51147, w51148, w51149, w51150, w51151, w51152, w51153, w51154, w51155, w51156, w51157, w51158, w51159, w51160, w51161, w51162, w51163, w51164, w51165, w51166, w51167, w51168, w51169, w51170, w51171, w51172, w51173, w51174, w51175, w51176, w51177, w51178, w51179, w51180, w51181, w51182, w51183, w51184, w51185, w51186, w51187, w51188, w51189, w51190, w51191, w51192, w51193, w51194, w51195, w51196, w51197, w51198, w51199, w51200, w51201, w51202, w51203, w51204, w51205, w51206, w51207, w51208, w51209, w51210, w51211, w51212, w51213, w51214, w51215, w51216, w51217, w51218, w51219, w51220, w51221, w51222, w51223, w51224, w51225, w51226, w51227, w51228, w51229, w51230, w51231, w51232, w51233, w51234, w51235, w51236, w51237, w51238, w51239, w51240, w51241, w51242, w51243, w51244, w51245, w51246, w51247, w51248, w51249, w51250, w51251, w51252, w51253, w51254, w51255, w51256, w51257, w51258, w51259, w51260, w51261, w51262, w51263, w51264, w51265, w51266, w51267, w51268, w51269, w51270, w51271, w51272, w51273, w51274, w51275, w51276, w51277, w51278, w51279, w51280, w51281, w51282, w51283, w51284, w51285, w51286, w51287, w51288, w51289, w51290, w51291, w51292, w51293, w51294, w51295, w51296, w51297, w51298, w51299, w51300, w51301, w51302, w51303, w51304, w51305, w51306, w51307, w51308, w51309, w51310, w51311, w51312, w51313, w51314, w51315, w51316, w51317, w51318, w51319, w51320, w51321, w51322, w51323, w51324, w51325, w51326, w51327, w51328, w51329, w51330, w51331, w51332, w51333, w51334, w51335, w51336, w51337, w51338, w51339, w51340, w51341, w51342, w51343, w51344, w51345, w51346, w51347, w51348, w51349, w51350, w51351, w51352, w51353, w51354, w51355, w51356, w51357, w51358, w51359, w51360, w51361, w51362, w51363, w51364, w51365, w51366, w51367, w51368, w51369, w51370, w51371, w51372, w51373, w51374, w51375, w51376, w51377, w51378, w51379, w51380, w51381, w51382, w51383, w51384, w51385, w51386, w51387, w51388, w51389, w51390, w51391, w51392, w51393, w51394, w51395, w51396, w51397, w51398, w51399, w51400, w51401, w51402, w51403, w51404, w51405, w51406, w51407, w51408, w51409, w51410, w51411, w51412, w51413, w51414, w51415, w51416, w51417, w51418, w51419, w51420, w51421, w51422, w51423, w51424, w51425, w51426, w51427, w51428, w51429, w51430, w51431, w51432, w51433, w51434, w51435, w51436, w51437, w51438, w51439, w51440, w51441, w51442, w51443, w51444, w51445, w51446, w51447, w51448, w51449, w51450, w51451, w51452, w51453, w51454, w51455, w51456, w51457, w51458, w51459, w51460, w51461, w51462, w51463, w51464, w51465, w51466, w51467, w51468, w51469, w51470, w51471, w51472, w51473, w51474, w51475, w51476, w51477, w51478, w51479, w51480, w51481, w51482, w51483, w51484, w51485, w51486, w51487, w51488, w51489, w51490, w51491, w51492, w51493, w51494, w51495, w51496, w51497, w51498, w51499, w51500, w51501, w51502, w51503, w51504, w51505, w51506, w51507, w51508, w51509, w51510, w51511, w51512, w51513, w51514, w51515, w51516, w51517, w51518, w51519, w51520, w51521, w51522, w51523, w51524, w51525, w51526, w51527, w51528, w51529, w51530, w51531, w51532, w51533, w51534, w51535, w51536, w51537, w51538, w51539, w51540, w51541, w51542, w51543, w51544, w51545, w51546, w51547, w51548, w51549, w51550, w51551, w51552, w51553, w51554, w51555, w51556, w51557, w51558, w51559, w51560, w51561, w51562, w51563, w51564, w51565, w51566, w51567, w51568, w51569, w51570, w51571, w51572, w51573, w51574, w51575, w51576, w51577, w51578, w51579, w51580, w51581, w51582, w51583, w51584, w51585, w51586, w51587, w51588, w51589, w51590, w51591, w51592, w51593, w51594, w51595, w51596, w51597, w51598, w51599, w51600, w51601, w51602, w51603, w51604, w51605, w51606, w51607, w51608, w51609, w51610, w51611, w51612, w51613, w51614, w51615, w51616, w51617, w51618, w51619, w51620, w51621, w51622, w51623, w51624, w51625, w51626, w51627, w51628, w51629, w51630, w51631, w51632, w51633, w51634, w51635, w51636, w51637, w51638, w51639, w51640, w51641, w51642, w51643, w51644, w51645, w51646, w51647, w51648, w51649, w51650, w51651, w51652, w51653, w51654, w51655, w51656, w51657, w51658, w51659, w51660, w51661, w51662, w51663, w51664, w51665, w51666, w51667, w51668, w51669, w51670, w51671, w51672, w51673, w51674, w51675, w51676, w51677, w51678, w51679, w51680, w51681, w51682, w51683, w51684, w51685, w51686, w51687, w51688, w51689, w51690, w51691, w51692, w51693, w51694, w51695, w51696, w51697, w51698, w51699, w51700, w51701, w51702, w51703, w51704, w51705, w51706, w51707, w51708, w51709, w51710, w51711, w51712, w51713, w51714, w51715, w51716, w51717, w51718, w51719, w51720, w51721, w51722, w51723, w51724, w51725, w51726, w51727, w51728, w51729, w51730, w51731, w51732, w51733, w51734, w51735, w51736, w51737, w51738, w51739, w51740, w51741, w51742, w51743, w51744, w51745, w51746, w51747, w51748, w51749, w51750, w51751, w51752, w51753, w51754, w51755, w51756, w51757, w51758, w51759, w51760, w51761, w51762, w51763, w51764, w51765, w51766, w51767, w51768, w51769, w51770, w51771, w51772, w51773, w51774, w51775, w51776, w51777, w51778, w51779, w51780, w51781, w51782, w51783, w51784, w51785, w51786, w51787, w51788, w51789, w51790, w51791, w51792, w51793, w51794, w51795, w51796, w51797, w51798, w51799, w51800, w51801, w51802, w51803, w51804, w51805, w51806, w51807, w51808, w51809, w51810, w51811, w51812, w51813, w51814, w51815, w51816, w51817, w51818, w51819, w51820, w51821, w51822, w51823, w51824, w51825, w51826, w51827, w51828, w51829, w51830, w51831, w51832, w51833, w51834, w51835, w51836, w51837, w51838, w51839, w51840, w51841, w51842, w51843, w51844, w51845, w51846, w51847, w51848, w51849, w51850, w51851, w51852, w51853, w51854, w51855, w51856, w51857, w51858, w51859, w51860, w51861, w51862, w51863, w51864, w51865, w51866, w51867, w51868, w51869, w51870, w51871, w51872, w51873, w51874, w51875, w51876, w51877, w51878, w51879, w51880, w51881, w51882, w51883, w51884, w51885, w51886, w51887, w51888, w51889, w51890, w51891, w51892, w51893, w51894, w51895, w51896, w51897, w51898, w51899, w51900, w51901, w51902, w51903, w51904, w51905, w51906, w51907, w51908, w51909, w51910, w51911, w51912, w51913, w51914, w51915, w51916, w51917, w51918, w51919, w51920, w51921, w51922, w51923, w51924, w51925, w51926, w51927, w51928, w51929, w51930, w51931, w51932, w51933, w51934, w51935, w51936, w51937, w51938, w51939, w51940, w51941, w51942, w51943, w51944, w51945, w51946, w51947, w51948, w51949, w51950, w51951, w51952, w51953, w51954, w51955, w51956, w51957, w51958, w51959, w51960, w51961, w51962, w51963, w51964, w51965, w51966, w51967, w51968, w51969, w51970, w51971, w51972, w51973, w51974, w51975, w51976, w51977, w51978, w51979, w51980, w51981, w51982, w51983, w51984, w51985, w51986, w51987, w51988, w51989, w51990, w51991, w51992, w51993, w51994, w51995, w51996, w51997, w51998, w51999, w52000, w52001, w52002, w52003, w52004, w52005, w52006, w52007, w52008, w52009, w52010, w52011, w52012, w52013, w52014, w52015, w52016, w52017, w52018, w52019, w52020, w52021, w52022, w52023, w52024, w52025, w52026, w52027, w52028, w52029, w52030, w52031, w52032, w52033, w52034, w52035, w52036, w52037, w52038, w52039, w52040, w52041, w52042, w52043, w52044, w52045, w52046, w52047, w52048, w52049, w52050, w52051, w52052, w52053, w52054, w52055, w52056, w52057, w52058, w52059, w52060, w52061, w52062, w52063, w52064, w52065, w52066, w52067, w52068, w52069, w52070, w52071, w52072, w52073, w52074, w52075, w52076, w52077, w52078, w52079, w52080, w52081, w52082, w52083, w52084, w52085, w52086, w52087, w52088, w52089, w52090, w52091, w52092, w52093, w52094, w52095, w52096, w52097, w52098, w52099, w52100, w52101, w52102, w52103, w52104, w52105, w52106, w52107, w52108, w52109, w52110, w52111, w52112, w52113, w52114, w52115, w52116, w52117, w52118, w52119, w52120, w52121, w52122, w52123, w52124, w52125, w52126, w52127, w52128, w52129, w52130, w52131, w52132, w52133, w52134, w52135, w52136, w52137, w52138, w52139, w52140, w52141, w52142, w52143, w52144, w52145, w52146, w52147, w52148, w52149, w52150, w52151, w52152, w52153, w52154, w52155, w52156, w52157, w52158, w52159, w52160, w52161, w52162, w52163, w52164, w52165, w52166, w52167, w52168, w52169, w52170, w52171, w52172, w52173, w52174, w52175, w52176, w52177, w52178, w52179, w52180, w52181, w52182, w52183, w52184, w52185, w52186, w52187, w52188, w52189, w52190, w52191, w52192, w52193, w52194, w52195, w52196, w52197, w52198, w52199, w52200, w52201, w52202, w52203, w52204, w52205, w52206, w52207, w52208, w52209, w52210, w52211, w52212, w52213, w52214, w52215, w52216, w52217, w52218, w52219, w52220, w52221, w52222, w52223, w52224, w52225, w52226, w52227, w52228, w52229, w52230, w52231, w52232, w52233, w52234, w52235, w52236, w52237, w52238, w52239, w52240, w52241, w52242, w52243, w52244, w52245, w52246, w52247, w52248, w52249, w52250, w52251, w52252, w52253, w52254, w52255, w52256, w52257, w52258, w52259, w52260, w52261, w52262, w52263, w52264, w52265, w52266, w52267, w52268, w52269, w52270, w52271, w52272, w52273, w52274, w52275, w52276, w52277, w52278, w52279, w52280, w52281, w52282, w52283, w52284, w52285, w52286, w52287, w52288, w52289, w52290, w52291, w52292, w52293, w52294, w52295, w52296, w52297, w52298, w52299, w52300, w52301, w52302, w52303, w52304, w52305, w52306, w52307, w52308, w52309, w52310, w52311, w52312, w52313, w52314, w52315, w52316, w52317, w52318, w52319, w52320, w52321, w52322, w52323, w52324, w52325, w52326, w52327, w52328, w52329, w52330, w52331, w52332, w52333, w52334, w52335, w52336, w52337, w52338, w52339, w52340, w52341, w52342, w52343;
assign w0 = a[126] & a[127];
assign w1 = ~a[124] & ~a[125];
assign w2 = ~a[126] & ~w1;
assign w3 = ~w0 & ~w2;
assign w4 = a[124] & ~a[125];
assign w5 = a[126] & ~w4;
assign w6 = a[123] & ~a[125];
assign w7 = ~a[123] & ~a[126];
assign w8 = a[125] & w7;
assign w9 = ~w6 & ~w8;
assign w10 = ~a[125] & a[126];
assign w11 = a[126] & ~a[127];
assign w12 = ~a[126] & a[127];
assign w13 = ~w11 & ~w12;
assign w14 = ~a[124] & ~w13;
assign w15 = ~w8 & ~w10;
assign w16 = w14 & ~w15;
assign w17 = (~w9 & w16) | (~w9 & w39641) | (w16 & w39641);
assign w18 = ~a[120] & ~a[121];
assign w19 = ~a[122] & ~w18;
assign w20 = a[123] & a[126];
assign w21 = ~w10 & ~w20;
assign w22 = w14 & ~w21;
assign w23 = a[124] & a[126];
assign w24 = a[125] & ~a[127];
assign w25 = a[123] & a[124];
assign w26 = w24 & ~w25;
assign w27 = ~a[123] & ~w23;
assign w28 = w26 & ~w27;
assign w29 = ~a[127] & ~w7;
assign w30 = w4 & ~w29;
assign w31 = ~w28 & ~w30;
assign w32 = ~w22 & w31;
assign w33 = w19 & w32;
assign w34 = ~w17 & w33;
assign w35 = ~a[122] & ~a[123];
assign w36 = a[125] & ~a[126];
assign w37 = ~a[125] & a[127];
assign w38 = ~w24 & ~w37;
assign w39 = a[126] & w38;
assign w40 = w38 & w39642;
assign w41 = a[124] & w36;
assign w42 = ~a[126] & ~a[127];
assign w43 = ~a[124] & ~a[127];
assign w44 = a[123] & ~w43;
assign w45 = w6 & w42;
assign w46 = ~w37 & w44;
assign w47 = a[124] & a[125];
assign w48 = ~w12 & ~w35;
assign w49 = ~a[124] & ~w48;
assign w50 = w38 & w47;
assign w51 = ~w38 & w49;
assign w52 = ~w50 & ~w51;
assign w53 = (a[122] & w46) | (a[122] & w39643) | (w46 & w39643);
assign w54 = w52 & ~w53;
assign w55 = (~w35 & w40) | (~w35 & w43865) | (w40 & w43865);
assign w56 = w52 & w46985;
assign w57 = ~w34 & w56;
assign w58 = ~w10 & ~w36;
assign w59 = ~a[123] & a[124];
assign w60 = ~w0 & w59;
assign w61 = w58 & w60;
assign w62 = a[122] & ~a[125];
assign w63 = w7 & w62;
assign w64 = ~a[127] & w63;
assign w65 = a[120] & ~a[121];
assign w66 = ~w61 & ~w64;
assign w67 = w65 & w66;
assign w68 = ~w38 & ~w47;
assign w69 = ~w49 & w68;
assign w70 = ~w16 & ~w69;
assign w71 = w67 & w70;
assign w72 = ~a[118] & ~a[119];
assign w73 = ~a[120] & w72;
assign w74 = ~a[126] & w1;
assign w75 = ~w0 & ~w24;
assign w76 = ~w74 & w75;
assign w77 = ~w1 & ~w43;
assign w78 = ~w12 & w35;
assign w79 = ~w77 & w78;
assign w80 = ~w76 & ~w79;
assign w81 = (a[121] & ~w72) | (a[121] & w39644) | (~w72 & w39644);
assign w82 = w18 & w72;
assign w83 = ~w81 & ~w82;
assign w84 = w80 & ~w83;
assign w85 = w72 & w50622;
assign w86 = (~w85 & ~w80) | (~w85 & w39645) | (~w80 & w39645);
assign w87 = ~w71 & w86;
assign w88 = ~w57 & ~w87;
assign w89 = ~w80 & w83;
assign w90 = (~w81 & w80) | (~w81 & w39646) | (w80 & w39646);
assign w91 = ~w71 & ~w90;
assign w92 = w57 & ~w91;
assign w93 = ~w88 & ~w92;
assign w94 = ~a[123] & ~a[127];
assign w95 = a[125] & a[126];
assign w96 = a[122] & w95;
assign w97 = ~w74 & ~w96;
assign w98 = ~a[124] & ~w58;
assign w99 = a[124] & ~a[126];
assign w100 = ~w94 & ~w99;
assign w101 = ~w13 & w98;
assign w102 = (~a[122] & w101) | (~a[122] & w39647) | (w101 & w39647);
assign w103 = w94 & ~w97;
assign w104 = ~w102 & ~w103;
assign w105 = ~w34 & w104;
assign w106 = ~a[126] & ~w24;
assign w107 = w68 & ~w106;
assign w108 = (~w18 & ~w68) | (~w18 & w50623) | (~w68 & w50623);
assign w109 = a[122] & ~w108;
assign w110 = (~w3 & w34) | (~w3 & w39649) | (w34 & w39649);
assign w111 = ~w108 & w50624;
assign w112 = (w111 & ~w54) | (w111 & w50625) | (~w54 & w50625);
assign w113 = ~w110 & ~w112;
assign w114 = w93 & w113;
assign w115 = w6 & w11;
assign w116 = ~w19 & ~w115;
assign w117 = (a[123] & w106) | (a[123] & w39650) | (w106 & w39650);
assign w118 = ~a[122] & w116;
assign w119 = ~w76 & w116;
assign w120 = ~w117 & w119;
assign w121 = ~w118 & ~w120;
assign w122 = ~w95 & ~w99;
assign w123 = ~w38 & w122;
assign w124 = ~w13 & w47;
assign w125 = ~w123 & ~w124;
assign w126 = ~w2 & ~w13;
assign w127 = w35 & w126;
assign w128 = ~w125 & w127;
assign w129 = (~w1 & w75) | (~w1 & w39651) | (w75 & w39651);
assign w130 = ~w11 & w52128;
assign w131 = (~a[123] & w58) | (~a[123] & w59) | (w58 & w59);
assign w132 = ~w129 & w131;
assign w133 = w130 & ~w132;
assign w134 = (~w35 & ~w58) | (~w35 & w39653) | (~w58 & w39653);
assign w135 = ~w24 & w35;
assign w136 = ~a[124] & ~w135;
assign w137 = ~w134 & w136;
assign w138 = a[127] & w35;
assign w139 = (w47 & w138) | (w47 & w39654) | (w138 & w39654);
assign w140 = ~w42 & ~w139;
assign w141 = ~w137 & w140;
assign w142 = ~w133 & ~w141;
assign w143 = ~w121 & ~w128;
assign w144 = w142 & ~w143;
assign w145 = (~a[127] & w4) | (~a[127] & w42) | (w4 & w42);
assign w146 = w23 & ~w35;
assign w147 = ~w145 & ~w146;
assign w148 = (~a[124] & w138) | (~a[124] & w39655) | (w138 & w39655);
assign w149 = w147 & ~w148;
assign w150 = w133 & ~w149;
assign w151 = ~w128 & ~w149;
assign w152 = ~w121 & w151;
assign w153 = ~w150 & ~w152;
assign w154 = ~w144 & w153;
assign w155 = (w109 & ~w54) | (w109 & w50626) | (~w54 & w50626);
assign w156 = w105 & ~w155;
assign w157 = w105 & w50627;
assign w158 = (~w157 & ~w93) | (~w157 & w50628) | (~w93 & w50628);
assign w159 = ~w42 & ~w154;
assign w160 = (w159 & w114) | (w159 & w39656) | (w114 & w39656);
assign w161 = (a[127] & ~w1) | (a[127] & w0) | (~w1 & w0);
assign w162 = w105 & w50786;
assign w163 = ~w1 & w42;
assign w164 = ~w7 & ~w20;
assign w165 = (a[123] & w24) | (a[123] & w20) | (w24 & w20);
assign w166 = a[126] & w47;
assign w167 = w165 & ~w166;
assign w168 = ~w2 & ~w164;
assign w169 = a[127] & w168;
assign w170 = ~w167 & ~w169;
assign w171 = a[124] & a[127];
assign w172 = (w171 & w8) | (w171 & w50788) | (w8 & w50788);
assign w173 = ~w11 & ~w77;
assign w174 = w44 & w106;
assign w175 = w18 & ~w174;
assign w176 = ~a[123] & ~w75;
assign w177 = ~w173 & w176;
assign w178 = w175 & ~w177;
assign w179 = ~a[122] & ~w178;
assign w180 = a[123] & w16;
assign w181 = ~w179 & ~w180;
assign w182 = (a[122] & ~w170) | (a[122] & w39657) | (~w170 & w39657);
assign w183 = w181 & ~w182;
assign w184 = ~w38 & w99;
assign w185 = ~w39 & ~w184;
assign w186 = (w19 & w185) | (w19 & w50789) | (w185 & w50789);
assign w187 = ~a[123] & ~w125;
assign w188 = w186 & ~w187;
assign w189 = (~w188 & ~w181) | (~w188 & w50790) | (~w181 & w50790);
assign w190 = (w163 & w71) | (w163 & w50791) | (w71 & w50791);
assign w191 = w57 & w190;
assign w192 = w189 & ~w191;
assign w193 = ~w57 & w50792;
assign w194 = w192 & ~w193;
assign w195 = (~w162 & ~w93) | (~w162 & w50787) | (~w93 & w50787);
assign w196 = w194 & w195;
assign w197 = ~w160 & ~w196;
assign w198 = (w42 & w183) | (w42 & w39658) | (w183 & w39658);
assign w199 = ~w154 & ~w198;
assign w200 = (~w3 & w71) | (~w3 & w39659) | (w71 & w39659);
assign w201 = ~w57 & w200;
assign w202 = (~w3 & w71) | (~w3 & w39660) | (w71 & w39660);
assign w203 = w57 & w202;
assign w204 = ~w201 & ~w203;
assign w205 = w154 & ~w189;
assign w206 = w3 & w93;
assign w207 = w204 & ~w205;
assign w208 = ~w206 & w207;
assign w209 = w156 & ~w208;
assign w210 = w199 & w204;
assign w211 = w158 & w210;
assign w212 = ~w209 & ~w211;
assign w213 = ~w209 & w50629;
assign w214 = (~w205 & w114) | (~w205 & w39661) | (w114 & w39661);
assign w215 = (~a[120] & w34) | (~a[120] & w50698) | (w34 & w50698);
assign w216 = w18 & ~w56;
assign w217 = (a[121] & w39644) | (a[121] & w57) | (w39644 & w57);
assign w218 = ~w216 & ~w217;
assign w219 = ~w84 & ~w89;
assign w220 = (w219 & w34) | (w219 & w46986) | (w34 & w46986);
assign w221 = ~w34 & w46987;
assign w222 = ~w220 & ~w221;
assign w223 = ~w205 & ~w222;
assign w224 = w199 & ~w222;
assign w225 = (~w224 & w158) | (~w224 & w39662) | (w158 & w39662);
assign w226 = ~w199 & w218;
assign w227 = ~w214 & w226;
assign w228 = w225 & ~w227;
assign w229 = ~w204 & w43866;
assign w230 = (~w3 & w204) | (~w3 & w50699) | (w204 & w50699);
assign w231 = w197 & w213;
assign w232 = ~w196 & w43867;
assign w233 = ~w228 & w232;
assign w234 = ~w231 & ~w233;
assign w235 = ~a[116] & ~a[117];
assign w236 = ~a[118] & w235;
assign w237 = ~w34 & w50793;
assign w238 = ~a[119] & ~w237;
assign w239 = ~w199 & w238;
assign w240 = ~w214 & w239;
assign w241 = ~w34 & w50700;
assign w242 = ~w72 & ~w241;
assign w243 = ~w205 & w242;
assign w244 = ~w158 & w243;
assign w245 = (w236 & w34) | (w236 & w50794) | (w34 & w50794);
assign w246 = (~w245 & ~w199) | (~w245 & w50701) | (~w199 & w50701);
assign w247 = ~w244 & w246;
assign w248 = ~w240 & w247;
assign w249 = (w80 & ~w247) | (w80 & w39664) | (~w247 & w39664);
assign w250 = w247 & w39665;
assign w251 = ~w249 & ~w250;
assign w252 = ~w199 & ~w214;
assign w253 = a[120] & ~w72;
assign w254 = ~w73 & ~w253;
assign w255 = ~w34 & w50702;
assign w256 = ~w215 & ~w255;
assign w257 = (w254 & w214) | (w254 & w50795) | (w214 & w50795);
assign w258 = ~w214 & w50796;
assign w259 = ~w257 & ~w258;
assign w260 = (w3 & w217) | (w3 & w50797) | (w217 & w50797);
assign w261 = ~w199 & ~w260;
assign w262 = w3 & w222;
assign w263 = ~w205 & ~w262;
assign w264 = w199 & ~w262;
assign w265 = (~w264 & w158) | (~w264 & w46988) | (w158 & w46988);
assign w266 = ~w214 & w261;
assign w267 = w265 & ~w266;
assign w268 = ~w196 & w39666;
assign w269 = ~w267 & w268;
assign w270 = (w259 & ~w234) | (w259 & w39667) | (~w234 & w39667);
assign w271 = ~w259 & ~w269;
assign w272 = w234 & w46989;
assign w273 = ~w270 & ~w272;
assign w274 = ~w272 & w39668;
assign w275 = w80 & w256;
assign w276 = ~w275 & w39669;
assign w277 = ~w214 & w276;
assign w278 = w80 & w254;
assign w279 = (w3 & ~w80) | (w3 & w50798) | (~w80 & w50798);
assign w280 = w199 & w279;
assign w281 = (w279 & ~w154) | (w279 & w50799) | (~w154 & w50799);
assign w282 = (~w280 & w158) | (~w280 & w39670) | (w158 & w39670);
assign w283 = ~w277 & w282;
assign w284 = w248 & ~w283;
assign w285 = ~w80 & ~w256;
assign w286 = ~w80 & ~w254;
assign w287 = ~w80 & w50798;
assign w288 = (w287 & w214) | (w287 & w50800) | (w214 & w50800);
assign w289 = w277 & w285;
assign w290 = ~w288 & ~w289;
assign w291 = ~w284 & w290;
assign w292 = w199 & w278;
assign w293 = (w278 & ~w154) | (w278 & w50801) | (~w154 & w50801);
assign w294 = (~w292 & w158) | (~w292 & w39671) | (w158 & w39671);
assign w295 = ~w199 & w275;
assign w296 = ~w214 & w295;
assign w297 = w294 & ~w296;
assign w298 = w248 & w297;
assign w299 = (~w3 & w80) | (~w3 & w50802) | (w80 & w50802);
assign w300 = (w299 & w214) | (w299 & w50803) | (w214 & w50803);
assign w301 = (~w3 & w256) | (~w3 & w536) | (w256 & w536);
assign w302 = ~w214 & w50804;
assign w303 = ~w300 & ~w302;
assign w304 = ~w298 & ~w303;
assign w305 = w291 & ~w304;
assign w306 = w305 & w39672;
assign w307 = ~w214 & w50703;
assign w308 = (w286 & w214) | (w286 & w50704) | (w214 & w50704);
assign w309 = ~w307 & ~w308;
assign w310 = ~w298 & w309;
assign w311 = w212 & w268;
assign w312 = w161 & ~w311;
assign w313 = ~w42 & ~w228;
assign w314 = (~w313 & w310) | (~w313 & w39673) | (w310 & w39673);
assign w315 = w126 & ~w311;
assign w316 = w310 & w315;
assign w317 = w314 & ~w316;
assign w318 = ~w306 & ~w317;
assign w319 = w163 & ~w228;
assign w320 = ~w213 & ~w319;
assign w321 = ~w42 & ~w197;
assign w322 = ~w3 & ~w228;
assign w323 = w321 & ~w322;
assign w324 = ~w298 & w43868;
assign w325 = w323 & ~w324;
assign w326 = w304 & w320;
assign w327 = ~w325 & ~w326;
assign w328 = w305 & w43869;
assign w329 = w327 & ~w328;
assign w330 = (w329 & w318) | (w329 & w50705) | (w318 & w50705);
assign w331 = (w3 & w272) | (w3 & w43870) | (w272 & w43870);
assign w332 = w329 & ~w331;
assign w333 = ~w298 & w46990;
assign w334 = ~a[114] & ~a[115];
assign w335 = ~a[116] & w334;
assign w336 = (w335 & w214) | (w335 & w50706) | (w214 & w50706);
assign w337 = w235 & ~w336;
assign w338 = ~w231 & w43871;
assign w339 = a[117] & ~w336;
assign w340 = (~w339 & w231) | (~w339 & w43872) | (w231 & w43872);
assign w341 = w269 & ~w339;
assign w342 = w310 & w341;
assign w343 = ~w340 & ~w342;
assign w344 = ~w333 & w338;
assign w345 = w343 & ~w344;
assign w346 = ~w214 & w50805;
assign w347 = ~w231 & w43873;
assign w348 = ~w333 & w347;
assign w349 = (w346 & w333) | (w346 & w43874) | (w333 & w43874);
assign w350 = ~w345 & ~w349;
assign w351 = w234 & ~w333;
assign w352 = a[118] & ~w235;
assign w353 = ~w236 & ~w352;
assign w354 = ~w34 & w50806;
assign w355 = (a[118] & w214) | (a[118] & w50707) | (w214 & w50707);
assign w356 = ~w214 & w50708;
assign w357 = ~w355 & ~w356;
assign w358 = w57 & w357;
assign w359 = ~w333 & w39674;
assign w360 = (w358 & w333) | (w358 & w39675) | (w333 & w39675);
assign w361 = ~w359 & ~w360;
assign w362 = (~w357 & w231) | (~w357 & w43875) | (w231 & w43875);
assign w363 = w269 & ~w357;
assign w364 = w310 & w363;
assign w365 = ~w362 & ~w364;
assign w366 = ~w57 & ~w365;
assign w367 = (w353 & w34) | (w353 & w50807) | (w34 & w50807);
assign w368 = ~w333 & w39676;
assign w369 = ~w366 & w39677;
assign w370 = w350 & w361;
assign w371 = w369 & ~w370;
assign w372 = (~w213 & w298) | (~w213 & w39678) | (w298 & w39678);
assign w373 = ~w284 & w39679;
assign w374 = w372 & ~w373;
assign w375 = w39666 & w50808;
assign w376 = (~w57 & w214) | (~w57 & w50709) | (w214 & w50709);
assign w377 = ~w214 & w50710;
assign w378 = ~w376 & ~w377;
assign w379 = ~w235 & ~w378;
assign w380 = (a[118] & w333) | (a[118] & w43877) | (w333 & w43877);
assign w381 = w236 & w378;
assign w382 = w234 & w381;
assign w383 = ~w333 & w382;
assign w384 = w365 & ~w383;
assign w385 = ~w380 & w384;
assign w386 = (a[119] & ~w385) | (a[119] & w39680) | (~w385 & w39680);
assign w387 = w385 & w39681;
assign w388 = ~w386 & ~w387;
assign w389 = w80 & ~w354;
assign w390 = ~w333 & w39682;
assign w391 = (w80 & ~w357) | (w80 & w33829) | (~w357 & w33829);
assign w392 = (w391 & w333) | (w391 & w39683) | (w333 & w39683);
assign w393 = ~w390 & ~w392;
assign w394 = (w80 & w366) | (w80 & w39684) | (w366 & w39684);
assign w395 = w350 & ~w393;
assign w396 = ~w394 & ~w395;
assign w397 = (~w330 & w371) | (~w330 & w39685) | (w371 & w39685);
assign w398 = ~w330 & w396;
assign w399 = ~w388 & w398;
assign w400 = ~w397 & ~w399;
assign w401 = ~a[112] & ~a[113];
assign w402 = ~a[114] & w401;
assign w403 = (~w402 & w333) | (~w402 & w50809) | (w333 & w50809);
assign w404 = ~a[115] & ~w403;
assign w405 = ~w399 & w39686;
assign w406 = a[115] & ~w403;
assign w407 = (w406 & w399) | (w406 & w39687) | (w399 & w39687);
assign w408 = ~w405 & ~w407;
assign w409 = a[114] & ~a[115];
assign w410 = ~w333 & w50810;
assign w411 = (~w252 & ~w408) | (~w252 & w50632) | (~w408 & w50632);
assign w412 = ~w333 & w50811;
assign w413 = (a[116] & w333) | (a[116] & w50812) | (w333 & w50812);
assign w414 = a[116] & ~w334;
assign w415 = ~w335 & ~w414;
assign w416 = ~w412 & ~w413;
assign w417 = ~w399 & w43878;
assign w418 = (w415 & w399) | (w415 & w43879) | (w399 & w43879);
assign w419 = ~w417 & ~w418;
assign w420 = w252 & ~w410;
assign w421 = (~w39688 & w50633) | (~w39688 & w50634) | (w50633 & w50634);
assign w422 = w408 & w421;
assign w423 = ~w419 & ~w422;
assign w424 = ~w411 & ~w423;
assign w425 = ~w345 & w50813;
assign w426 = (w57 & w345) | (w57 & w50814) | (w345 & w50814);
assign w427 = ~w425 & ~w426;
assign w428 = (w427 & w399) | (w427 & w39689) | (w399 & w39689);
assign w429 = ~w333 & w50815;
assign w430 = w365 & ~w429;
assign w431 = w80 & ~w430;
assign w432 = (~w39689 & w50635) | (~w39689 & w50636) | (w50635 & w50636);
assign w433 = w80 & w430;
assign w434 = (w39689 & w50637) | (w39689 & w50638) | (w50637 & w50638);
assign w435 = ~w432 & ~w434;
assign w436 = ~w330 & ~w371;
assign w437 = w396 & w436;
assign w438 = (~w388 & ~w436) | (~w388 & w43880) | (~w436 & w43880);
assign w439 = ~w332 & w388;
assign w440 = w437 & w439;
assign w441 = ~w438 & ~w440;
assign w442 = ~w440 & w43881;
assign w443 = w435 & ~w442;
assign w444 = ~w336 & ~w346;
assign w445 = (a[117] & w333) | (a[117] & w50762) | (w333 & w50762);
assign w446 = ~w348 & ~w445;
assign w447 = w444 & ~w446;
assign w448 = ~w444 & w446;
assign w449 = ~w447 & ~w448;
assign w450 = a[117] & ~w412;
assign w451 = ~a[117] & w412;
assign w452 = ~w450 & ~w451;
assign w453 = (w449 & w399) | (w449 & w39690) | (w399 & w39690);
assign w454 = ~w399 & w39691;
assign w455 = ~w453 & ~w454;
assign w456 = ~w57 & w455;
assign w457 = w443 & ~w456;
assign w458 = w424 & w457;
assign w459 = w57 & ~w455;
assign w460 = ~w80 & ~w430;
assign w461 = (w39689 & w50639) | (w39689 & w50640) | (w50639 & w50640);
assign w462 = ~w80 & w430;
assign w463 = (~w39689 & w50641) | (~w39689 & w50642) | (w50641 & w50642);
assign w464 = ~w461 & ~w463;
assign w465 = ~w459 & w464;
assign w466 = ~w388 & w396;
assign w467 = (~w331 & w370) | (~w331 & w39692) | (w370 & w39692);
assign w468 = (~w274 & w466) | (~w274 & w39693) | (w466 & w39693);
assign w469 = (w42 & w466) | (w42 & w50711) | (w466 & w50711);
assign w470 = (w329 & w466) | (w329 & w50816) | (w466 & w50816);
assign w471 = ~w468 & ~w469;
assign w472 = ~w470 & ~w471;
assign w473 = (w3 & w440) | (w3 & w43882) | (w440 & w43882);
assign w474 = (w228 & ~w351) | (w228 & w50817) | (~w351 & w50817);
assign w475 = ~w306 & ~w474;
assign w476 = ~w468 & ~w475;
assign w477 = ~w468 & w50712;
assign w478 = ~w473 & ~w477;
assign w479 = ~w472 & w478;
assign w480 = (w479 & w465) | (w479 & w50643) | (w465 & w50643);
assign w481 = ~w458 & w480;
assign w482 = ~w466 & w39695;
assign w483 = (w3 & w466) | (w3 & w39696) | (w466 & w39696);
assign w484 = ~w482 & ~w483;
assign w485 = (w273 & ~w484) | (w273 & w43883) | (~w484 & w43883);
assign w486 = ~w273 & ~w330;
assign w487 = w484 & w486;
assign w488 = ~w485 & ~w487;
assign w489 = ~w329 & w468;
assign w490 = ~w476 & ~w489;
assign w491 = ~w42 & w490;
assign w492 = ~w488 & w491;
assign w493 = (~w492 & w458) | (~w492 & w50644) | (w458 & w50644);
assign w494 = w435 & ~w456;
assign w495 = (w494 & w424) | (w494 & w39697) | (w424 & w39697);
assign w496 = w464 & ~w495;
assign w497 = (w3 & w458) | (w3 & w50645) | (w458 & w50645);
assign w498 = w496 & w497;
assign w499 = (~w3 & w458) | (~w3 & w50646) | (w458 & w50646);
assign w500 = ~w496 & w499;
assign w501 = ~w498 & ~w500;
assign w502 = w441 & w501;
assign w503 = ~w495 & w50647;
assign w504 = ~w492 & w50713;
assign w505 = (w504 & w495) | (w504 & w50648) | (w495 & w50648);
assign w506 = ~w503 & ~w505;
assign w507 = (~w473 & w465) | (~w473 & w50763) | (w465 & w50763);
assign w508 = (w458 & w50764) | (w458 & w50765) | (w50764 & w50765);
assign w509 = (w490 & w458) | (w490 & w50766) | (w458 & w50766);
assign w510 = w508 & ~w509;
assign w511 = w42 & w506;
assign w512 = (~w510 & w502) | (~w510 & w39698) | (w502 & w39698);
assign w513 = ~w423 & w50649;
assign w514 = (w57 & w423) | (w57 & w50650) | (w423 & w50650);
assign w515 = ~w513 & ~w514;
assign w516 = w80 & ~w455;
assign w517 = w493 & w39699;
assign w518 = w80 & w455;
assign w519 = (w518 & ~w493) | (w518 & w39700) | (~w493 & w39700);
assign w520 = ~w517 & ~w519;
assign w521 = w3 & w520;
assign w522 = w428 & ~w430;
assign w523 = ~w428 & w430;
assign w524 = ~w522 & ~w523;
assign w525 = w80 & ~w524;
assign w526 = w464 & w52129;
assign w527 = (w424 & w43885) | (w424 & w43886) | (w43885 & w43886);
assign w528 = w493 & w39702;
assign w529 = ~w435 & w52129;
assign w530 = ~w80 & w524;
assign w531 = (w424 & w43887) | (w424 & w43888) | (w43887 & w43888);
assign w532 = ~w529 & ~w531;
assign w533 = (~w458 & w50651) | (~w458 & w50652) | (w50651 & w50652);
assign w534 = w532 & ~w533;
assign w535 = ~w528 & w534;
assign w536 = ~w3 & w80;
assign w537 = ~w455 & w536;
assign w538 = w493 & w39704;
assign w539 = w455 & w536;
assign w540 = (w539 & ~w493) | (w539 & w39705) | (~w493 & w39705);
assign w541 = ~w538 & ~w540;
assign w542 = w535 & w541;
assign w543 = ~w521 & ~w542;
assign w544 = (w506 & ~w501) | (w506 & w39706) | (~w501 & w39706);
assign w545 = ~w42 & ~w544;
assign w546 = ~w543 & ~w545;
assign w547 = (w512 & w543) | (w512 & w50714) | (w543 & w50714);
assign w548 = ~w411 & ~w422;
assign w549 = (~w458 & w50653) | (~w458 & w50654) | (w50653 & w50654);
assign w550 = (w39708 & w458) | (w39708 & w50655) | (w458 & w50655);
assign w551 = ~w549 & ~w550;
assign w552 = w57 & ~w551;
assign w553 = ~w80 & ~w455;
assign w554 = (w553 & ~w493) | (w553 & w39709) | (~w493 & w39709);
assign w555 = ~w80 & w455;
assign w556 = w493 & w39710;
assign w557 = ~w554 & ~w556;
assign w558 = ~w552 & w557;
assign w559 = w534 & w50715;
assign w560 = w558 & ~w559;
assign w561 = w512 & w560;
assign w562 = ~a[110] & ~a[111];
assign w563 = (w562 & w399) | (w562 & w50767) | (w399 & w50767);
assign w564 = ~a[112] & w562;
assign w565 = ~w399 & w43889;
assign w566 = (~w401 & ~w565) | (~w401 & w50818) | (~w565 & w50818);
assign w567 = ~a[112] & w563;
assign w568 = ~a[113] & ~w565;
assign w569 = ~w567 & ~w568;
assign w570 = (w351 & w566) | (w351 & w50819) | (w566 & w50819);
assign w571 = ~w481 & w39711;
assign w572 = w351 & ~w569;
assign w573 = (~w458 & w50656) | (~w458 & w50657) | (w50656 & w50657);
assign w574 = ~w571 & ~w573;
assign w575 = (a[114] & w399) | (a[114] & w50820) | (w399 & w50820);
assign w576 = ~w399 & w50821;
assign w577 = ~w575 & ~w576;
assign w578 = a[114] & ~w401;
assign w579 = (~w458 & w50658) | (~w458 & w50659) | (w50658 & w50659);
assign w580 = ~w402 & ~w578;
assign w581 = (w39714 & w458) | (w39714 & w50660) | (w458 & w50660);
assign w582 = ~w579 & ~w581;
assign w583 = w574 & w582;
assign w584 = ~w566 & w50822;
assign w585 = ~w481 & w39715;
assign w586 = ~w351 & w569;
assign w587 = (~w458 & w50661) | (~w458 & w50662) | (w50661 & w50662);
assign w588 = ~w585 & ~w587;
assign w589 = ~w403 & ~w410;
assign w590 = (a[115] & w399) | (a[115] & w43890) | (w399 & w43890);
assign w591 = ~w399 & w43891;
assign w592 = ~w590 & ~w591;
assign w593 = w589 & w592;
assign w594 = ~w589 & ~w592;
assign w595 = ~w593 & ~w594;
assign w596 = (~w409 & w592) | (~w409 & w50823) | (w592 & w50823);
assign w597 = w252 & w595;
assign w598 = ~w481 & w39717;
assign w599 = (w592 & w50824) | (w592 & w50825) | (w50824 & w50825);
assign w600 = (w599 & w481) | (w599 & w39718) | (w481 & w39718);
assign w601 = ~w598 & ~w600;
assign w602 = w588 & w601;
assign w603 = ~w583 & w602;
assign w604 = (w39719 & w458) | (w39719 & w50663) | (w458 & w50663);
assign w605 = (~w458 & w50664) | (~w458 & w50665) | (w50664 & w50665);
assign w606 = ~w604 & ~w605;
assign w607 = ~w252 & w606;
assign w608 = ~w57 & w551;
assign w609 = ~w607 & ~w608;
assign w610 = ~w603 & w609;
assign w611 = w561 & ~w610;
assign w612 = ~w547 & ~w611;
assign w613 = a[113] & ~w493;
assign w614 = ~w565 & ~w567;
assign w615 = ~a[113] & w493;
assign w616 = ~w613 & ~w615;
assign w617 = w614 & ~w616;
assign w618 = ~w614 & w616;
assign w619 = ~w617 & ~w618;
assign w620 = (w619 & w39721) | (w619 & w612) | (w39721 & w612);
assign w621 = ~a[112] & w493;
assign w622 = (a[113] & ~w493) | (a[113] & w50826) | (~w493 & w50826);
assign w623 = w493 & w401;
assign w624 = ~w622 & ~w623;
assign w625 = (~w624 & w611) | (~w624 & w50827) | (w611 & w50827);
assign w626 = (w351 & w39722) | (w351 & w612) | (w39722 & w612);
assign w627 = ~w620 & w626;
assign w628 = w574 & w588;
assign w629 = ~w611 & w50828;
assign w630 = w252 & w582;
assign w631 = (w611 & w50768) | (w611 & w50769) | (w50768 & w50769);
assign w632 = w252 & ~w582;
assign w633 = ~w611 & w50770;
assign w634 = ~w631 & ~w633;
assign w635 = ~w583 & w39725;
assign w636 = (w252 & w583) | (w252 & w39726) | (w583 & w39726);
assign w637 = ~w635 & ~w636;
assign w638 = ~w561 & w637;
assign w639 = ~w606 & w637;
assign w640 = ~w611 & w50716;
assign w641 = (w606 & ~w638) | (w606 & w50717) | (~w638 & w50717);
assign w642 = ~w640 & ~w641;
assign w643 = ~w57 & ~w642;
assign w644 = ~w252 & ~w582;
assign w645 = (w611 & w50771) | (w611 & w50772) | (w50771 & w50772);
assign w646 = ~w252 & w582;
assign w647 = ~w611 & w50773;
assign w648 = ~w645 & ~w647;
assign w649 = ~w643 & w648;
assign w650 = w627 & w634;
assign w651 = w649 & ~w650;
assign w652 = a[110] & ~a[111];
assign w653 = ~a[108] & ~a[109];
assign w654 = ~a[110] & w653;
assign w655 = ~w493 & ~w654;
assign w656 = (a[111] & w493) | (a[111] & w50829) | (w493 & w50829);
assign w657 = (w493 & w50832) | (w493 & w50833) | (w50832 & w50833);
assign w658 = (~a[111] & w493) | (~a[111] & w50843) | (w493 & w50843);
assign w659 = w493 & w654;
assign w660 = (w50834 & w493) | (w50834 & w50844) | (w493 & w50844);
assign w661 = w493 & w50835;
assign w662 = (~w611 & w50718) | (~w611 & w50719) | (w50718 & w50719);
assign w663 = ~w611 & w50720;
assign w664 = w662 & ~w663;
assign w665 = a[112] & ~w493;
assign w666 = a[112] & ~w562;
assign w667 = ~w564 & ~w666;
assign w668 = ~w621 & ~w665;
assign w669 = (w668 & w611) | (w668 & w50721) | (w611 & w50721);
assign w670 = ~w611 & w50722;
assign w671 = ~w669 & ~w670;
assign w672 = w664 & w671;
assign w673 = w658 & ~w659;
assign w674 = (w673 & w611) | (w673 & w50723) | (w611 & w50723);
assign w675 = w656 & ~w659;
assign w676 = ~w611 & w50724;
assign w677 = ~w674 & ~w676;
assign w678 = (w400 & ~w493) | (w400 & w50836) | (~w493 & w50836);
assign w679 = (w611 & w50774) | (w611 & w50775) | (w50774 & w50775);
assign w680 = w677 & w679;
assign w681 = (w39731 & w611) | (w39731 & w50776) | (w611 & w50776);
assign w682 = ~w351 & w619;
assign w683 = (w682 & w39732) | (w682 & w612) | (w39732 & w612);
assign w684 = ~w681 & ~w683;
assign w685 = ~w680 & w684;
assign w686 = ~w672 & w685;
assign w687 = ~w634 & ~w643;
assign w688 = w686 & ~w687;
assign w689 = w651 & ~w688;
assign w690 = w57 & w642;
assign w691 = ~w603 & w39733;
assign w692 = (w57 & w603) | (w57 & w39734) | (w603 & w39734);
assign w693 = ~w691 & ~w692;
assign w694 = (~w551 & w547) | (~w551 & w39735) | (w547 & w39735);
assign w695 = ~w551 & w52130;
assign w696 = w612 & w39736;
assign w697 = ~w695 & ~w696;
assign w698 = ~w690 & w697;
assign w699 = w560 & ~w610;
assign w700 = ~w42 & ~w510;
assign w701 = ~w699 & w39737;
assign w702 = (w545 & w699) | (w545 & w39738) | (w699 & w39738);
assign w703 = ~w701 & ~w702;
assign w704 = (w455 & ~w493) | (w455 & w43892) | (~w493 & w43892);
assign w705 = w493 & w43893;
assign w706 = ~w704 & ~w705;
assign w707 = w80 & ~w706;
assign w708 = w557 & ~w707;
assign w709 = ~w708 & w52131;
assign w710 = ~w546 & w39739;
assign w711 = w709 & ~w710;
assign w712 = (~w80 & ~w560) | (~w80 & w50725) | (~w560 & w50725);
assign w713 = ~w547 & w712;
assign w714 = ~w706 & ~w713;
assign w715 = (w558 & w603) | (w558 & w50667) | (w603 & w50667);
assign w716 = ~w547 & ~w715;
assign w717 = ~w710 & w50778;
assign w718 = (w3 & w547) | (w3 & w723) | (w547 & w723);
assign w719 = ~w714 & w718;
assign w720 = ~w717 & ~w719;
assign w721 = ~w521 & w541;
assign w722 = (~w50667 & w50726) | (~w50667 & w50727) | (w50726 & w50727);
assign w723 = ~w610 & w39740;
assign w724 = ~w722 & ~w723;
assign w725 = (w42 & ~w534) | (w42 & w50837) | (~w534 & w50837);
assign w726 = (w725 & ~w612) | (w725 & w50728) | (~w612 & w50728);
assign w727 = w534 & w50838;
assign w728 = (w727 & w546) | (w727 & w39741) | (w546 & w39741);
assign w729 = ~w724 & w728;
assign w730 = w703 & ~w729;
assign w731 = ~w726 & w730;
assign w732 = w720 & ~w731;
assign w733 = w698 & w732;
assign w734 = (w733 & w688) | (w733 & w39742) | (w688 & w39742);
assign w735 = (~w711 & w714) | (~w711 & w39743) | (w714 & w39743);
assign w736 = (~w535 & ~w612) | (~w535 & w50729) | (~w612 & w50729);
assign w737 = (w535 & w546) | (w535 & w43894) | (w546 & w43894);
assign w738 = ~w724 & w737;
assign w739 = ~w736 & ~w738;
assign w740 = (~w703 & w736) | (~w703 & w39744) | (w736 & w39744);
assign w741 = ~w699 & w43895;
assign w742 = (w544 & w699) | (w544 & w43896) | (w699 & w43896);
assign w743 = ~w741 & ~w742;
assign w744 = w161 & w743;
assign w745 = w735 & w744;
assign w746 = ~w740 & ~w745;
assign w747 = ~w739 & w39745;
assign w748 = w746 & ~w747;
assign w749 = w612 & w39746;
assign w750 = ~w694 & ~w749;
assign w751 = ~w749 & w43897;
assign w752 = w732 & w751;
assign w753 = w748 & ~w752;
assign w754 = ~w734 & w753;
assign w755 = ~w651 & w698;
assign w756 = ~w687 & w698;
assign w757 = w686 & w756;
assign w758 = ~w755 & ~w757;
assign w759 = (~w750 & ~w758) | (~w750 & w39747) | (~w758 & w39747);
assign w760 = ~w643 & ~w690;
assign w761 = (w760 & w688) | (w760 & w39748) | (w688 & w39748);
assign w762 = ~w732 & ~w740;
assign w763 = ~w732 & w39749;
assign w764 = (~w643 & w763) | (~w643 & w43898) | (w763 & w43898);
assign w765 = ~w761 & w764;
assign w766 = ~w759 & ~w765;
assign w767 = (w42 & w736) | (w42 & w50839) | (w736 & w50839);
assign w768 = ~w80 & ~w767;
assign w769 = w762 & w768;
assign w770 = ~w758 & w769;
assign w771 = (w3 & ~w766) | (w3 & w43899) | (~w766 & w43899);
assign w772 = ~w711 & w52132;
assign w773 = ~w751 & ~w772;
assign w774 = ~w736 & w50841;
assign w775 = w774 & w52133;
assign w776 = ~w42 & ~w743;
assign w777 = (w758 & w50845) | (w758 & w50846) | (w50845 & w50846);
assign w778 = ~w775 & ~w777;
assign w779 = w43897 & w50668;
assign w780 = (w3 & ~w43897) | (w3 & w50669) | (~w43897 & w50669);
assign w781 = ~w779 & ~w780;
assign w782 = w3 & ~w758;
assign w783 = w758 & w781;
assign w784 = ~w782 & ~w783;
assign w785 = w42 & ~w735;
assign w786 = w784 & w785;
assign w787 = w735 & w739;
assign w788 = w42 & w787;
assign w789 = ~w784 & w788;
assign w790 = ~w786 & ~w789;
assign w791 = w778 & w790;
assign w792 = w790 & w43900;
assign w793 = w735 & ~w781;
assign w794 = ~w735 & ~w740;
assign w795 = w781 & w794;
assign w796 = ~w793 & ~w795;
assign w797 = ~w720 & ~w740;
assign w798 = ~w772 & ~w797;
assign w799 = ~w711 & w52134;
assign w800 = (~w799 & w758) | (~w799 & w43901) | (w758 & w43901);
assign w801 = (~w796 & w758) | (~w796 & w46991) | (w758 & w46991);
assign w802 = w800 & ~w801;
assign w803 = (w758 & w43902) | (w758 & w43903) | (w43902 & w43903);
assign w804 = (~w42 & w736) | (~w42 & w50848) | (w736 & w50848);
assign w805 = w804 & w52133;
assign w806 = ~w803 & ~w805;
assign w807 = ~w802 & ~w806;
assign w808 = (~w627 & ~w685) | (~w627 & w39752) | (~w685 & w39752);
assign w809 = w634 & w648;
assign w810 = ~w808 & w809;
assign w811 = w648 & ~w760;
assign w812 = ~w810 & w811;
assign w813 = ~w761 & ~w812;
assign w814 = w754 & ~w813;
assign w815 = (w642 & ~w748) | (w642 & w50779) | (~w748 & w50779);
assign w816 = w642 & w733;
assign w817 = ~w689 & w816;
assign w818 = ~w815 & ~w817;
assign w819 = ~w814 & w818;
assign w820 = ~w80 & ~w819;
assign w821 = w582 & ~w629;
assign w822 = ~w582 & w629;
assign w823 = ~w821 & ~w822;
assign w824 = w808 & ~w809;
assign w825 = ~w810 & ~w824;
assign w826 = (~w57 & ~w754) | (~w57 & w43904) | (~w754 & w43904);
assign w827 = ~w754 & ~w823;
assign w828 = w826 & ~w827;
assign w829 = ~w820 & w828;
assign w830 = ~w817 & w39753;
assign w831 = ~w814 & w830;
assign w832 = (~w3 & w758) | (~w3 & w43905) | (w758 & w43905);
assign w833 = w766 & w832;
assign w834 = ~w831 & ~w833;
assign w835 = (~w807 & ~w791) | (~w807 & w39754) | (~w791 & w39754);
assign w836 = ~w807 & w834;
assign w837 = ~w829 & w836;
assign w838 = ~w835 & ~w837;
assign w839 = ~w620 & ~w625;
assign w840 = ~w672 & ~w680;
assign w841 = w351 & ~w840;
assign w842 = ~w351 & w840;
assign w843 = ~w841 & ~w842;
assign w844 = w753 & ~w843;
assign w845 = (w839 & ~w844) | (w839 & w50730) | (~w844 & w50730);
assign w846 = w844 & w50731;
assign w847 = ~w845 & ~w846;
assign w848 = ~w252 & ~w847;
assign w849 = w664 & ~w680;
assign w850 = w748 & w50732;
assign w851 = ~w734 & w850;
assign w852 = ~w351 & w671;
assign w853 = ~w851 & w852;
assign w854 = ~w351 & ~w671;
assign w855 = w851 & w854;
assign w856 = ~w853 & ~w855;
assign w857 = w252 & ~w839;
assign w858 = (w857 & ~w844) | (w857 & w50733) | (~w844 & w50733);
assign w859 = w252 & w839;
assign w860 = w844 & w50734;
assign w861 = ~w858 & ~w860;
assign w862 = w856 & w861;
assign w863 = ~w655 & ~w659;
assign w864 = (a[111] & w611) | (a[111] & w50849) | (w611 & w50849);
assign w865 = ~w611 & w50850;
assign w866 = ~w864 & ~w865;
assign w867 = ~w863 & ~w866;
assign w868 = w677 & ~w867;
assign w869 = ~w863 & w864;
assign w870 = (~w652 & ~w866) | (~w652 & w50851) | (~w866 & w50851);
assign w871 = (w870 & ~w748) | (w870 & w50735) | (~w748 & w50735);
assign w872 = w733 & w870;
assign w873 = ~w689 & w872;
assign w874 = ~w871 & ~w873;
assign w875 = ~w873 & w39755;
assign w876 = ~w734 & w43906;
assign w877 = w875 & ~w876;
assign w878 = (w400 & ~w875) | (w400 & w43907) | (~w875 & w43907);
assign w879 = ~a[106] & ~a[107];
assign w880 = ~a[108] & w879;
assign w881 = (~w880 & w611) | (~w880 & w50852) | (w611 & w50852);
assign w882 = (~w653 & ~w881) | (~w653 & w50853) | (~w881 & w50853);
assign w883 = w748 & w50736;
assign w884 = ~w734 & w883;
assign w885 = ~a[109] & ~w881;
assign w886 = ~w611 & w50854;
assign w887 = (~w886 & ~w733) | (~w886 & w39756) | (~w733 & w39756);
assign w888 = w649 & w50855;
assign w889 = ~w688 & w888;
assign w890 = ~w887 & ~w889;
assign w891 = (w885 & ~w748) | (w885 & w50856) | (~w748 & w50856);
assign w892 = ~w890 & ~w891;
assign w893 = (w493 & ~w892) | (w493 & w39757) | (~w892 & w39757);
assign w894 = ~w752 & ~w868;
assign w895 = (~w400 & ~w864) | (~w400 & w50857) | (~w864 & w50857);
assign w896 = (w895 & ~w894) | (w895 & w39758) | (~w894 & w39758);
assign w897 = w733 & w895;
assign w898 = ~w689 & w897;
assign w899 = ~w896 & ~w898;
assign w900 = w874 & ~w899;
assign w901 = a[109] & ~a[110];
assign w902 = a[110] & w653;
assign w903 = ~w879 & ~w901;
assign w904 = ~w611 & w50858;
assign w905 = ~w901 & ~w902;
assign w906 = (a[109] & ~w879) | (a[109] & w50869) | (~w879 & w50869);
assign w907 = ~a[110] & ~w653;
assign w908 = ~w906 & w907;
assign w909 = ~w908 & w52135;
assign w910 = (a[110] & w611) | (a[110] & w51480) | (w611 & w51480);
assign w911 = ~w611 & w50860;
assign w912 = ~w910 & ~w911;
assign w913 = w879 & w653;
assign w914 = (a[110] & w880) | (a[110] & w50861) | (w880 & w50861);
assign w915 = ~w913 & ~w914;
assign w916 = ~w493 & w915;
assign w917 = ~w910 & w50862;
assign w918 = (w917 & ~w748) | (w917 & w50737) | (~w748 & w50737);
assign w919 = w733 & w917;
assign w920 = ~w689 & w919;
assign w921 = ~w918 & ~w920;
assign w922 = w748 & w50738;
assign w923 = ~w734 & w922;
assign w924 = w921 & ~w923;
assign w925 = ~w900 & w924;
assign w926 = ~w893 & w925;
assign w927 = (~w878 & ~w925) | (~w878 & w43908) | (~w925 & w43908);
assign w928 = w671 & ~w851;
assign w929 = ~w671 & w851;
assign w930 = ~w928 & ~w929;
assign w931 = w351 & w930;
assign w932 = ~w848 & ~w862;
assign w933 = ~w848 & ~w931;
assign w934 = (~w932 & w927) | (~w932 & w39759) | (w927 & w39759);
assign w935 = ~w838 & ~w934;
assign w936 = w57 & ~w823;
assign w937 = (w936 & w734) | (w936 & w43909) | (w734 & w43909);
assign w938 = w57 & ~w825;
assign w939 = w754 & w938;
assign w940 = ~w937 & ~w939;
assign w941 = ~w831 & ~w940;
assign w942 = ~w820 & ~w941;
assign w943 = w792 & w942;
assign w944 = ~w838 & ~w943;
assign w945 = ~w935 & ~w944;
assign w946 = (w940 & w848) | (w940 & w43910) | (w848 & w43910);
assign w947 = (~w931 & w926) | (~w931 & w39760) | (w926 & w39760);
assign w948 = w862 & w940;
assign w949 = (~w946 & w947) | (~w946 & w43911) | (w947 & w43911);
assign w950 = ~w820 & ~w831;
assign w951 = w949 & ~w950;
assign w952 = ~w949 & w950;
assign w953 = ~w951 & ~w952;
assign w954 = ~w819 & w945;
assign w955 = ~w945 & ~w953;
assign w956 = ~w954 & ~w955;
assign w957 = w3 & ~w956;
assign w958 = ~w820 & w946;
assign w959 = ~w820 & w948;
assign w960 = ~w947 & w959;
assign w961 = ~w958 & ~w960;
assign w962 = ~w960 & w43912;
assign w963 = ~w42 & ~w802;
assign w964 = ~w962 & w50863;
assign w965 = (~w806 & w962) | (~w806 & w50864) | (w962 & w50864);
assign w966 = ~w964 & ~w965;
assign w967 = ~w771 & ~w833;
assign w968 = ~w831 & ~w838;
assign w969 = w961 & w968;
assign w970 = w3 & w838;
assign w971 = w792 & w39761;
assign w972 = w934 & w971;
assign w973 = ~w970 & ~w972;
assign w974 = ~w969 & w973;
assign w975 = w967 & ~w974;
assign w976 = ~w967 & w974;
assign w977 = ~w975 & ~w976;
assign w978 = ~w966 & ~w977;
assign w979 = w957 & ~w978;
assign w980 = ~w967 & w969;
assign w981 = w967 & w974;
assign w982 = ~w981 & w43913;
assign w983 = w966 & ~w982;
assign w984 = ~w979 & ~w983;
assign w985 = ~a[104] & ~a[105];
assign w986 = ~a[106] & w985;
assign w987 = ~w754 & ~w986;
assign w988 = w754 & w986;
assign w989 = w934 & w943;
assign w990 = (~w879 & w754) | (~w879 & w50866) | (w754 & w50866);
assign w991 = ~w838 & w990;
assign w992 = ~w989 & w991;
assign w993 = ~w988 & ~w992;
assign w994 = (~a[107] & w754) | (~a[107] & w50867) | (w754 & w50867);
assign w995 = w945 & w994;
assign w996 = w993 & ~w995;
assign w997 = ~a[108] & w754;
assign w998 = a[108] & ~w754;
assign w999 = ~w997 & ~w998;
assign w1000 = a[108] & ~w879;
assign w1001 = ~w880 & ~w1000;
assign w1002 = ~w612 & ~w999;
assign w1003 = w945 & w1002;
assign w1004 = (~w1001 & w611) | (~w1001 & w50868) | (w611 & w50868);
assign w1005 = ~w945 & w1004;
assign w1006 = ~w1003 & ~w1005;
assign w1007 = ~w996 & w1006;
assign w1008 = ~w612 & ~w754;
assign w1009 = w612 & w754;
assign w1010 = ~w1008 & ~w1009;
assign w1011 = ~w906 & ~w913;
assign w1012 = w1010 & ~w1011;
assign w1013 = ~w1010 & w1011;
assign w1014 = ~w1012 & ~w1013;
assign w1015 = (a[109] & ~w754) | (a[109] & w50869) | (~w754 & w50869);
assign w1016 = w754 & w653;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = w493 & w1017;
assign w1019 = w945 & w1018;
assign w1020 = w493 & ~w1014;
assign w1021 = ~w945 & w1020;
assign w1022 = ~w1019 & ~w1021;
assign w1023 = w612 & w999;
assign w1024 = w945 & w1023;
assign w1025 = ~w611 & w50870;
assign w1026 = ~w945 & w1025;
assign w1027 = ~w1024 & ~w1026;
assign w1028 = w1022 & w1027;
assign w1029 = ~w1007 & w1028;
assign w1030 = w892 & w50871;
assign w1031 = ~w893 & ~w1030;
assign w1032 = ~w838 & w1031;
assign w1033 = ~w989 & w1032;
assign w1034 = ~w754 & ~w912;
assign w1035 = ~w902 & ~w907;
assign w1036 = w754 & w1035;
assign w1037 = ~w1034 & ~w1036;
assign w1038 = w400 & ~w1037;
assign w1039 = ~w1033 & w1038;
assign w1040 = w400 & w1037;
assign w1041 = w1033 & w1040;
assign w1042 = ~w1039 & ~w1041;
assign w1043 = ~w493 & w1014;
assign w1044 = ~w945 & w1043;
assign w1045 = ~w493 & ~w1017;
assign w1046 = w945 & w1045;
assign w1047 = ~w1044 & ~w1046;
assign w1048 = w1042 & w1047;
assign w1049 = (w351 & w926) | (w351 & w39762) | (w926 & w39762);
assign w1050 = ~w926 & w39763;
assign w1051 = ~w1049 & ~w1050;
assign w1052 = ~w838 & ~w1051;
assign w1053 = ~w989 & w1052;
assign w1054 = w252 & ~w930;
assign w1055 = ~w1053 & w1054;
assign w1056 = w252 & w930;
assign w1057 = w1053 & w1056;
assign w1058 = ~w1055 & ~w1057;
assign w1059 = ~w893 & w924;
assign w1060 = ~w878 & ~w900;
assign w1061 = w1059 & ~w1060;
assign w1062 = ~w1059 & w1060;
assign w1063 = ~w1061 & ~w1062;
assign w1064 = w875 & w50872;
assign w1065 = w945 & w1064;
assign w1066 = w351 & w1063;
assign w1067 = ~w945 & w1066;
assign w1068 = ~w1065 & ~w1067;
assign w1069 = ~w252 & w930;
assign w1070 = ~w1053 & w1069;
assign w1071 = ~w252 & ~w930;
assign w1072 = w1053 & w1071;
assign w1073 = ~w1070 & ~w1072;
assign w1074 = w1058 & ~w1068;
assign w1075 = w1073 & ~w1074;
assign w1076 = (~w400 & w1033) | (~w400 & w39764) | (w1033 & w39764);
assign w1077 = w1033 & w1037;
assign w1078 = w1076 & ~w1077;
assign w1079 = (w252 & w947) | (w252 & w39765) | (w947 & w39765);
assign w1080 = ~w252 & w856;
assign w1081 = ~w947 & w1080;
assign w1082 = ~w838 & ~w1081;
assign w1083 = (~w847 & ~w792) | (~w847 & w39766) | (~w792 & w39766);
assign w1084 = (w847 & ~w1082) | (w847 & w39767) | (~w1082 & w39767);
assign w1085 = w1082 & w39768;
assign w1086 = ~w1084 & ~w1085;
assign w1087 = ~w57 & w1086;
assign w1088 = ~w1078 & ~w1087;
assign w1089 = w1075 & w1088;
assign w1090 = ~w1029 & w1048;
assign w1091 = w1089 & ~w1090;
assign w1092 = ~w828 & w940;
assign w1093 = (w57 & w838) | (w57 & w43914) | (w838 & w43914);
assign w1094 = (w1092 & w1093) | (w1092 & w39769) | (w1093 & w39769);
assign w1095 = ~w1093 & w39770;
assign w1096 = ~w1094 & ~w1095;
assign w1097 = ~w80 & w1096;
assign w1098 = (~w351 & ~w875) | (~w351 & w50873) | (~w875 & w50873);
assign w1099 = w945 & w1098;
assign w1100 = ~w351 & ~w1063;
assign w1101 = ~w945 & w1100;
assign w1102 = ~w1099 & ~w1101;
assign w1103 = w1073 & ~w1102;
assign w1104 = w57 & w847;
assign w1105 = (w1104 & ~w1082) | (w1104 & w39771) | (~w1082 & w39771);
assign w1106 = ~w847 & w52136;
assign w1107 = w1082 & w50875;
assign w1108 = ~w1105 & ~w1107;
assign w1109 = w1058 & w1108;
assign w1110 = ~w1103 & w1109;
assign w1111 = ~w1087 & ~w1110;
assign w1112 = (~w1097 & w1110) | (~w1097 & w39772) | (w1110 & w39772);
assign w1113 = ~w1091 & w1112;
assign w1114 = ~w955 & w39773;
assign w1115 = ~w42 & ~w977;
assign w1116 = (~w1114 & w977) | (~w1114 & w43915) | (w977 & w43915);
assign w1117 = w80 & ~w1096;
assign w1118 = ~w1115 & w39774;
assign w1119 = (w1118 & w1091) | (w1118 & w39775) | (w1091 & w39775);
assign w1120 = w984 & ~w1119;
assign w1121 = w984 & w1113;
assign w1122 = w984 & ~w1118;
assign w1123 = w1068 & w1102;
assign w1124 = ~w1078 & w1123;
assign w1125 = ~w1090 & w1124;
assign w1126 = w1078 & ~w1123;
assign w1127 = w1048 & ~w1123;
assign w1128 = ~w1029 & w1127;
assign w1129 = ~w1126 & ~w1128;
assign w1130 = ~w1125 & w1129;
assign w1131 = w877 & w945;
assign w1132 = ~w945 & w1063;
assign w1133 = ~w1131 & ~w1132;
assign w1134 = ~w979 & w43916;
assign w1135 = ~w1119 & w1134;
assign w1136 = ~w1122 & w1130;
assign w1137 = ~w1121 & w1136;
assign w1138 = ~w1135 & ~w1137;
assign w1139 = (w252 & w1137) | (w252 & w39776) | (w1137 & w39776);
assign w1140 = w1058 & w1073;
assign w1141 = w1048 & w1102;
assign w1142 = ~w1029 & w1141;
assign w1143 = (w1102 & ~w1123) | (w1102 & w39777) | (~w1123 & w39777);
assign w1144 = (~w1140 & w1142) | (~w1140 & w39778) | (w1142 & w39778);
assign w1145 = ~w1142 & w39779;
assign w1146 = ~w1144 & ~w1145;
assign w1147 = ~w930 & ~w1053;
assign w1148 = w930 & w1053;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = w57 & w1146;
assign w1151 = ~w1120 & w1150;
assign w1152 = w57 & ~w1149;
assign w1153 = ~w1119 & w43917;
assign w1154 = ~w1151 & ~w1153;
assign w1155 = ~w1139 & w1154;
assign w1156 = ~w1137 & w43918;
assign w1157 = ~w1029 & w1047;
assign w1158 = (~w1157 & ~w984) | (~w1157 & w39780) | (~w984 & w39780);
assign w1159 = ~w1121 & w1158;
assign w1160 = ~w979 & w43919;
assign w1161 = w1042 & ~w1078;
assign w1162 = w351 & w1161;
assign w1163 = (w1162 & w1159) | (w1162 & w39781) | (w1159 & w39781);
assign w1164 = w351 & ~w1161;
assign w1165 = ~w1159 & w39782;
assign w1166 = ~w1163 & ~w1165;
assign w1167 = ~w1156 & w1166;
assign w1168 = w1155 & ~w1167;
assign w1169 = ~w1097 & ~w1117;
assign w1170 = (w1169 & w1091) | (w1169 & w39783) | (w1091 & w39783);
assign w1171 = ~w1111 & ~w1169;
assign w1172 = ~w1091 & w1171;
assign w1173 = ~w979 & w43920;
assign w1174 = ~w1172 & ~w1173;
assign w1175 = ~w983 & ~w1116;
assign w1176 = w1096 & w1175;
assign w1177 = (~w1176 & ~w1174) | (~w1176 & w39784) | (~w1174 & w39784);
assign w1178 = ~w3 & w1177;
assign w1179 = (~w1117 & w1091) | (~w1117 & w39785) | (w1091 & w39785);
assign w1180 = (w956 & w982) | (w956 & w50876) | (w982 & w50876);
assign w1181 = (~w1114 & w978) | (~w1114 & w50252) | (w978 & w50252);
assign w1182 = ~w979 & w39786;
assign w1183 = ~w1180 & w1181;
assign w1184 = ~w1179 & w1183;
assign w1185 = ~w1180 & ~w1182;
assign w1186 = w1179 & w1185;
assign w1187 = ~w1184 & ~w1186;
assign w1188 = ~w42 & w1187;
assign w1189 = ~w1178 & ~w1188;
assign w1190 = w3 & ~w1177;
assign w1191 = ~w1087 & w1108;
assign w1192 = w1058 & ~w1191;
assign w1193 = ~w1058 & w1191;
assign w1194 = ~w1192 & ~w1193;
assign w1195 = w1145 & w1191;
assign w1196 = ~w1145 & ~w1194;
assign w1197 = ~w1195 & ~w1196;
assign w1198 = ~w1120 & ~w1197;
assign w1199 = ~w979 & w43921;
assign w1200 = ~w1119 & w1199;
assign w1201 = (~w80 & w1119) | (~w80 & w43922) | (w1119 & w43922);
assign w1202 = ~w1198 & w1201;
assign w1203 = ~w1190 & ~w1202;
assign w1204 = w80 & ~w1197;
assign w1205 = ~w57 & ~w1146;
assign w1206 = w80 & w1086;
assign w1207 = ~w57 & w1149;
assign w1208 = ~w1206 & ~w1207;
assign w1209 = ~w1119 & w50877;
assign w1210 = ~w1120 & ~w1205;
assign w1211 = ~w1204 & w1210;
assign w1212 = ~w1209 & ~w1211;
assign w1213 = w1203 & w1212;
assign w1214 = w1189 & ~w1213;
assign w1215 = ~w1168 & w1214;
assign w1216 = ~w42 & w966;
assign w1217 = (w1179 & w50878) | (w1179 & w50879) | (w50878 & w50879);
assign w1218 = ~w42 & w977;
assign w1219 = w1218 & w52137;
assign w1220 = ~w1217 & ~w1219;
assign w1221 = w42 & ~w1187;
assign w1222 = w1220 & ~w1221;
assign w1223 = w1189 & ~w1203;
assign w1224 = w1222 & ~w1223;
assign w1225 = ~a[102] & ~a[103];
assign w1226 = ~a[104] & w1225;
assign w1227 = (a[105] & ~w1225) | (a[105] & w50880) | (~w1225 & w50880);
assign w1228 = ~w985 & ~w1227;
assign w1229 = w985 & ~w1225;
assign w1230 = (~w1229 & ~w945) | (~w1229 & w50881) | (~w945 & w50881);
assign w1231 = w985 & w1225;
assign w1232 = (~w1231 & w945) | (~w1231 & w50882) | (w945 & w50882);
assign w1233 = ~w979 & w51481;
assign w1234 = ~w1119 & w1233;
assign w1235 = (w1230 & ~w984) | (w1230 & w39787) | (~w984 & w39787);
assign w1236 = ~w1121 & w1235;
assign w1237 = ~w1234 & ~w1236;
assign w1238 = a[106] & ~w945;
assign w1239 = ~a[106] & w945;
assign w1240 = ~w1238 & ~w1239;
assign w1241 = ~w754 & w1240;
assign w1242 = ~w979 & w50883;
assign w1243 = a[106] & ~w985;
assign w1244 = ~w986 & ~w1243;
assign w1245 = ~w754 & ~w1244;
assign w1246 = (~w1245 & ~w984) | (~w1245 & w39788) | (~w984 & w39788);
assign w1247 = ~w1121 & w1246;
assign w1248 = ~w1119 & w1242;
assign w1249 = ~w1247 & ~w1248;
assign w1250 = w754 & ~w1240;
assign w1251 = ~w1119 & w50884;
assign w1252 = w754 & w1244;
assign w1253 = (w1252 & w1119) | (w1252 & w50885) | (w1119 & w50885);
assign w1254 = ~w1251 & ~w1253;
assign w1255 = ~w1237 & ~w1249;
assign w1256 = w1254 & ~w1255;
assign w1257 = a[106] & a[107];
assign w1258 = ~w979 & w50886;
assign w1259 = ~w987 & ~w988;
assign w1260 = a[107] & ~w945;
assign w1261 = ~a[107] & w945;
assign w1262 = ~w1260 & ~w1261;
assign w1263 = w1259 & ~w1262;
assign w1264 = (~w1263 & ~w984) | (~w1263 & w39789) | (~w984 & w39789);
assign w1265 = ~w1121 & w1264;
assign w1266 = ~w1119 & w1258;
assign w1267 = ~w1265 & ~w1266;
assign w1268 = ~w1259 & w1262;
assign w1269 = (w1268 & ~w984) | (w1268 & w39790) | (~w984 & w39790);
assign w1270 = ~w1121 & w1269;
assign w1271 = ~w1238 & w1262;
assign w1272 = ~w979 & w50887;
assign w1273 = ~w1119 & w1272;
assign w1274 = ~w1270 & ~w1273;
assign w1275 = ~w1267 & w1274;
assign w1276 = w612 & w1275;
assign w1277 = ~w612 & ~w1275;
assign w1278 = w612 & ~w996;
assign w1279 = ~w612 & w996;
assign w1280 = ~w1278 & ~w1279;
assign w1281 = (w1280 & ~w984) | (w1280 & w39791) | (~w984 & w39791);
assign w1282 = w945 & w999;
assign w1283 = ~w945 & w1001;
assign w1284 = ~w1282 & ~w1283;
assign w1285 = ~w1121 & w39792;
assign w1286 = (~w1284 & w1121) | (~w1284 & w39793) | (w1121 & w39793);
assign w1287 = ~w1285 & ~w1286;
assign w1288 = ~w493 & w1287;
assign w1289 = ~w1277 & ~w1288;
assign w1290 = w1256 & ~w1276;
assign w1291 = w1289 & ~w1290;
assign w1292 = w493 & ~w1287;
assign w1293 = ~w1007 & w1027;
assign w1294 = (w1022 & w1121) | (w1022 & w39794) | (w1121 & w39794);
assign w1295 = ~w1293 & ~w1294;
assign w1296 = w1029 & w1047;
assign w1297 = (w1296 & ~w984) | (w1296 & w39795) | (~w984 & w39795);
assign w1298 = ~w1121 & w1297;
assign w1299 = ~w945 & ~w1014;
assign w1300 = w945 & w1017;
assign w1301 = ~w1299 & ~w1300;
assign w1302 = ~w979 & w43923;
assign w1303 = ~w1119 & w1302;
assign w1304 = ~w1298 & ~w1303;
assign w1305 = ~w1295 & w1304;
assign w1306 = ~w400 & ~w1305;
assign w1307 = ~w1292 & ~w1306;
assign w1308 = ~w1291 & w1307;
assign w1309 = ~w1159 & w39796;
assign w1310 = (w1161 & w1159) | (w1161 & w39797) | (w1159 & w39797);
assign w1311 = ~w1309 & ~w1310;
assign w1312 = ~w351 & w1311;
assign w1313 = ~w1298 & w39798;
assign w1314 = ~w1295 & w1313;
assign w1315 = w1155 & ~w1314;
assign w1316 = ~w1312 & w1315;
assign w1317 = ~w1215 & w1224;
assign w1318 = w1224 & w1316;
assign w1319 = ~w1308 & w1318;
assign w1320 = ~w1317 & ~w1319;
assign w1321 = ~w1120 & w1146;
assign w1322 = ~w1119 & w50888;
assign w1323 = ~w1321 & ~w1322;
assign w1324 = (w1291 & w43924) | (w1291 & w43925) | (w43924 & w43925);
assign w1325 = w1166 & ~w1324;
assign w1326 = ~w1321 & w50889;
assign w1327 = w1154 & ~w1326;
assign w1328 = (w1316 & w1291) | (w1316 & w39800) | (w1291 & w39800);
assign w1329 = w1156 & ~w1327;
assign w1330 = ~w1319 & w39801;
assign w1331 = ~w1328 & w43926;
assign w1332 = ~w1139 & ~w1327;
assign w1333 = (w1332 & w1324) | (w1332 & w50890) | (w1324 & w50890);
assign w1334 = w1330 & w50891;
assign w1335 = (~w1323 & w1319) | (~w1323 & w50254) | (w1319 & w50254);
assign w1336 = ~w1334 & ~w1335;
assign w1337 = (~a[104] & w1119) | (~a[104] & w50892) | (w1119 & w50892);
assign w1338 = a[105] & ~w1337;
assign w1339 = ~a[105] & w1337;
assign w1340 = ~w1338 & ~w1339;
assign w1341 = ~w1227 & ~w1231;
assign w1342 = ~w1119 & w50893;
assign w1343 = (w945 & w1119) | (w945 & w50894) | (w1119 & w50894);
assign w1344 = ~w1342 & ~w1343;
assign w1345 = w1341 & w1344;
assign w1346 = ~w1341 & ~w1344;
assign w1347 = ~w1345 & ~w1346;
assign w1348 = (~w1340 & w1319) | (~w1340 & w39802) | (w1319 & w39802);
assign w1349 = ~w1319 & w39803;
assign w1350 = ~w1348 & ~w1349;
assign w1351 = ~a[100] & ~a[101];
assign w1352 = w1225 & w1351;
assign w1353 = ~a[102] & w1351;
assign w1354 = (a[103] & ~w1351) | (a[103] & w50895) | (~w1351 & w50895);
assign w1355 = (~w1354 & w1119) | (~w1354 & w50896) | (w1119 & w50896);
assign w1356 = ~w1225 & ~w1354;
assign w1357 = ~w1119 & w50897;
assign w1358 = w1225 & ~w1351;
assign w1359 = (w945 & w1357) | (w945 & w50898) | (w1357 & w50898);
assign w1360 = ~w1319 & w39804;
assign w1361 = ~w1355 & w50899;
assign w1362 = (w1361 & w1319) | (w1361 & w39805) | (w1319 & w39805);
assign w1363 = ~w1360 & ~w1362;
assign w1364 = ~w1119 & w50900;
assign w1365 = a[104] & ~w1225;
assign w1366 = ~w1226 & ~w1365;
assign w1367 = ~w1337 & ~w1364;
assign w1368 = (w1367 & w1319) | (w1367 & w39806) | (w1319 & w39806);
assign w1369 = ~w1319 & w39807;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = w1363 & ~w1370;
assign w1372 = (~w945 & w1355) | (~w945 & w50901) | (w1355 & w50901);
assign w1373 = (w1372 & w1319) | (w1372 & w39808) | (w1319 & w39808);
assign w1374 = ~w1357 & w50902;
assign w1375 = ~w1319 & w39809;
assign w1376 = ~w1373 & ~w1375;
assign w1377 = ~w754 & ~w1350;
assign w1378 = ~w1350 & w1376;
assign w1379 = ~w1371 & w1378;
assign w1380 = ~w1377 & ~w1379;
assign w1381 = ~w1249 & w1254;
assign w1382 = w1237 & ~w1381;
assign w1383 = ~w1237 & w1381;
assign w1384 = ~w1382 & ~w1383;
assign w1385 = ~w1119 & w50903;
assign w1386 = (w1244 & w1119) | (w1244 & w50904) | (w1119 & w50904);
assign w1387 = ~w1385 & ~w1386;
assign w1388 = ~w1319 & w39810;
assign w1389 = (~w1387 & w1319) | (~w1387 & w39811) | (w1319 & w39811);
assign w1390 = ~w1388 & ~w1389;
assign w1391 = ~w612 & w1390;
assign w1392 = ~w754 & w1376;
assign w1393 = ~w1371 & w1392;
assign w1394 = ~w1391 & ~w1393;
assign w1395 = w1380 & w1394;
assign w1396 = ~w1256 & ~w1277;
assign w1397 = ~w1396 & w39812;
assign w1398 = (~w493 & w1396) | (~w493 & w50905) | (w1396 & w50905);
assign w1399 = ~w1397 & ~w1398;
assign w1400 = w400 & w1287;
assign w1401 = ~w493 & w1275;
assign w1402 = (~w1401 & w1396) | (~w1401 & w39813) | (w1396 & w39813);
assign w1403 = ~w1397 & w1402;
assign w1404 = ~w1255 & w50906;
assign w1405 = w493 & w1275;
assign w1406 = w1404 & ~w1405;
assign w1407 = w1275 & ~w1400;
assign w1408 = (~w1407 & ~w1320) | (~w1407 & w39814) | (~w1320 & w39814);
assign w1409 = (w612 & w1255) | (w612 & w50907) | (w1255 & w50907);
assign w1410 = ~w1404 & ~w1409;
assign w1411 = ~w1319 & w39815;
assign w1412 = w1275 & w1411;
assign w1413 = ~w1408 & ~w1412;
assign w1414 = w400 & ~w1287;
assign w1415 = w1320 & w43927;
assign w1416 = w1413 & ~w1415;
assign w1417 = w1413 & w43928;
assign w1418 = w612 & ~w1390;
assign w1419 = ~w400 & ~w1287;
assign w1420 = (w1419 & ~w1320) | (w1419 & w39816) | (~w1320 & w39816);
assign w1421 = ~w400 & w1287;
assign w1422 = w1320 & w39817;
assign w1423 = ~w1420 & ~w1422;
assign w1424 = ~w351 & w1423;
assign w1425 = ~w1418 & w1424;
assign w1426 = ~w1417 & w1425;
assign w1427 = ~w1395 & w1426;
assign w1428 = ~w1306 & ~w1314;
assign w1429 = (~w1428 & w1291) | (~w1428 & w50908) | (w1291 & w50908);
assign w1430 = (~w1314 & ~w1320) | (~w1314 & w50909) | (~w1320 & w50909);
assign w1431 = (w1305 & w1319) | (w1305 & w50910) | (w1319 & w50910);
assign w1432 = (~w1431 & w1430) | (~w1431 & w50911) | (w1430 & w50911);
assign w1433 = (w1287 & ~w1320) | (w1287 & w39818) | (~w1320 & w39818);
assign w1434 = w1320 & w39819;
assign w1435 = ~w1433 & ~w1434;
assign w1436 = ~w1416 & w1424;
assign w1437 = (w493 & w1435) | (w493 & w19000) | (w1435 & w19000);
assign w1438 = w1436 & ~w1437;
assign w1439 = (w1432 & ~w1436) | (w1432 & w50912) | (~w1436 & w50912);
assign w1440 = ~w1427 & w1439;
assign w1441 = (w351 & w1435) | (w351 & w43929) | (w1435 & w43929);
assign w1442 = ~w493 & ~w1275;
assign w1443 = ~w1411 & w1442;
assign w1444 = w1401 & w1411;
assign w1445 = ~w1443 & ~w1444;
assign w1446 = w1423 & ~w1445;
assign w1447 = w1441 & ~w1446;
assign w1448 = w1395 & w1447;
assign w1449 = w1418 & w1445;
assign w1450 = w1405 & ~w1411;
assign w1451 = w493 & ~w1275;
assign w1452 = w1411 & w1451;
assign w1453 = ~w1450 & ~w1452;
assign w1454 = w1423 & w1453;
assign w1455 = ~w1449 & w1454;
assign w1456 = w1441 & ~w1455;
assign w1457 = (~w1291 & w50255) | (~w1291 & w50256) | (w50255 & w50256);
assign w1458 = (w1291 & w43930) | (w1291 & w43931) | (w43930 & w43931);
assign w1459 = (w1311 & ~w1320) | (w1311 & w43932) | (~w1320 & w43932);
assign w1460 = w1320 & w43933;
assign w1461 = ~w1459 & ~w1460;
assign w1462 = ~w252 & w1461;
assign w1463 = (~w1462 & w1455) | (~w1462 & w43934) | (w1455 & w43934);
assign w1464 = ~w1448 & w1463;
assign w1465 = ~w1440 & w1464;
assign w1466 = ~w1139 & ~w1156;
assign w1467 = (w1138 & w1319) | (w1138 & w50913) | (w1319 & w50913);
assign w1468 = ~w1319 & w39821;
assign w1469 = ~w1325 & w1468;
assign w1470 = ~w1319 & w39822;
assign w1471 = w1325 & w1470;
assign w1472 = ~w1469 & ~w1471;
assign w1473 = ~w1467 & w1472;
assign w1474 = (~w57 & ~w1472) | (~w57 & w43935) | (~w1472 & w43935);
assign w1475 = ~w1334 & w43936;
assign w1476 = ~w1474 & ~w1475;
assign w1477 = w1465 & w1476;
assign w1478 = (~w80 & w1334) | (~w80 & w46992) | (w1334 & w46992);
assign w1479 = w252 & ~w1461;
assign w1480 = w1472 & w43937;
assign w1481 = ~w1479 & ~w1480;
assign w1482 = w1476 & ~w1481;
assign w1483 = ~w1478 & ~w1482;
assign w1484 = ~w1328 & w43938;
assign w1485 = ~w1198 & ~w1200;
assign w1486 = (w80 & w1198) | (w80 & w50914) | (w1198 & w50914);
assign w1487 = (~w1202 & w1319) | (~w1202 & w46993) | (w1319 & w46993);
assign w1488 = (~w1202 & w1328) | (~w1202 & w50257) | (w1328 & w50257);
assign w1489 = (~w1485 & w1319) | (~w1485 & w46994) | (w1319 & w46994);
assign w1490 = w1320 & ~w1488;
assign w1491 = ~w1489 & ~w1490;
assign w1492 = w1484 & ~w1487;
assign w1493 = ~w1491 & ~w1492;
assign w1494 = ~w1328 & w43941;
assign w1495 = (w1328 & w51482) | (w1328 & w51483) | (w51482 & w51483);
assign w1496 = w50916 & w52138;
assign w1497 = ~w1495 & ~w1496;
assign w1498 = ~w42 & w1497;
assign w1499 = ~w1178 & ~w1190;
assign w1500 = ~w1319 & w39823;
assign w1501 = ~w1494 & w1500;
assign w1502 = (w1499 & w1501) | (w1499 & w39825) | (w1501 & w39825);
assign w1503 = ~w1501 & w39826;
assign w1504 = ~w1502 & ~w1503;
assign w1505 = w42 & w1504;
assign w1506 = (~w1498 & ~w1504) | (~w1498 & w50917) | (~w1504 & w50917);
assign w1507 = (w1493 & w1505) | (w1493 & w46996) | (w1505 & w46996);
assign w1508 = w1483 & w1507;
assign w1509 = (w1508 & ~w1465) | (w1508 & w43942) | (~w1465 & w43942);
assign w1510 = (w3 & w1491) | (w3 & w46997) | (w1491 & w46997);
assign w1511 = ~w1478 & ~w1510;
assign w1512 = w1481 & w1511;
assign w1513 = ~w1491 & w46998;
assign w1514 = (~w1513 & ~w1511) | (~w1513 & w39827) | (~w1511 & w39827);
assign w1515 = ~w1474 & ~w1481;
assign w1516 = (~w3 & w536) | (~w3 & w1336) | (w536 & w1336);
assign w1517 = ~w1515 & w50918;
assign w1518 = ~w1475 & ~w1493;
assign w1519 = w163 & w1504;
assign w1520 = ~w1518 & w1519;
assign w1521 = ~w1498 & ~w1520;
assign w1522 = w1504 & w50919;
assign w1523 = w1474 & w1522;
assign w1524 = ~w1517 & w1521;
assign w1525 = w1521 & ~w1523;
assign w1526 = (~w1524 & ~w1465) | (~w1524 & w50920) | (~w1465 & w50920);
assign w1527 = ~w1504 & w1514;
assign w1528 = (w1527 & w1465) | (w1527 & w43943) | (w1465 & w43943);
assign w1529 = w1526 & ~w1528;
assign w1530 = ~w1474 & w1481;
assign w1531 = (w80 & w1481) | (w80 & w46999) | (w1481 & w46999);
assign w1532 = ~w1481 & w47000;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = w1465 & w39828;
assign w1535 = (~w1533 & ~w1465) | (~w1533 & w43944) | (~w1465 & w43944);
assign w1536 = ~w1534 & ~w1535;
assign w1537 = (~w1336 & w1529) | (~w1336 & w43945) | (w1529 & w43945);
assign w1538 = (w1465 & w48589) | (w1465 & w48590) | (w48589 & w48590);
assign w1539 = ~w1529 & w43946;
assign w1540 = ~w1537 & ~w1539;
assign w1541 = (~w1509 & ~w1526) | (~w1509 & w43947) | (~w1526 & w43947);
assign w1542 = ~w1465 & w47001;
assign w1543 = (w57 & w1465) | (w57 & w47002) | (w1465 & w47002);
assign w1544 = ~w1542 & ~w1543;
assign w1545 = (w80 & ~w1472) | (w80 & w50921) | (~w1472 & w50921);
assign w1546 = (w1545 & ~w1541) | (w1545 & w39829) | (~w1541 & w39829);
assign w1547 = w1472 & w50922;
assign w1548 = w1541 & w39830;
assign w1549 = ~w1546 & ~w1548;
assign w1550 = ~a[98] & ~a[99];
assign w1551 = ~a[100] & w1550;
assign w1552 = (~w1551 & w1319) | (~w1551 & w50923) | (w1319 & w50923);
assign w1553 = a[101] & w1552;
assign w1554 = (~w1351 & ~w1552) | (~w1351 & w50924) | (~w1552 & w50924);
assign w1555 = ~w1319 & w50925;
assign w1556 = a[101] & ~w1555;
assign w1557 = ~w1552 & ~w1556;
assign w1558 = ~w1529 & w39833;
assign w1559 = ~w1556 & w50926;
assign w1560 = (w1559 & w1529) | (w1559 & w39834) | (w1529 & w39834);
assign w1561 = ~w1558 & ~w1560;
assign w1562 = a[102] & ~w1351;
assign w1563 = ~w1319 & w50927;
assign w1564 = (a[102] & w1319) | (a[102] & w50928) | (w1319 & w50928);
assign w1565 = ~w1563 & ~w1564;
assign w1566 = (w1565 & w1529) | (w1565 & w39835) | (w1529 & w39835);
assign w1567 = ~w1353 & ~w1562;
assign w1568 = ~w1529 & w39836;
assign w1569 = ~w1566 & ~w1568;
assign w1570 = w1561 & w1569;
assign w1571 = (w1120 & w1529) | (w1120 & w39837) | (w1529 & w39837);
assign w1572 = (w1557 & w1529) | (w1557 & w43948) | (w1529 & w43948);
assign w1573 = w1571 & ~w1572;
assign w1574 = a[103] & ~w1563;
assign w1575 = ~a[103] & w1563;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = ~w1352 & ~w1354;
assign w1578 = (w1577 & w1119) | (w1577 & w50929) | (w1119 & w50929);
assign w1579 = ~w1119 & w50930;
assign w1580 = ~w1578 & ~w1579;
assign w1581 = ~w1319 & w50931;
assign w1582 = (w1580 & w1319) | (w1580 & w50932) | (w1319 & w50932);
assign w1583 = ~w1581 & ~w1582;
assign w1584 = w945 & w1583;
assign w1585 = ~w1529 & w39838;
assign w1586 = w945 & ~w1576;
assign w1587 = (w1586 & w1529) | (w1586 & w39839) | (w1529 & w39839);
assign w1588 = ~w1585 & ~w1587;
assign w1589 = ~w1573 & w1588;
assign w1590 = w1363 & w1376;
assign w1591 = (w1465 & w51461) | (w1465 & w51462) | (w51461 & w51462);
assign w1592 = (~w1529 & w47003) | (~w1529 & w47004) | (w47003 & w47004);
assign w1593 = ~w1529 & w43949;
assign w1594 = w1592 & ~w1593;
assign w1595 = w1589 & w39841;
assign w1596 = (~w1576 & w1529) | (~w1576 & w39842) | (w1529 & w39842);
assign w1597 = ~w1529 & w39843;
assign w1598 = ~w1596 & ~w1597;
assign w1599 = ~w945 & w1598;
assign w1600 = ~w1594 & w1599;
assign w1601 = (w754 & w1371) | (w754 & w50933) | (w1371 & w50933);
assign w1602 = ~w1393 & ~w1601;
assign w1603 = w612 & w1350;
assign w1604 = (w1603 & w1529) | (w1603 & w39845) | (w1529 & w39845);
assign w1605 = w612 & ~w1350;
assign w1606 = ~w1529 & w39846;
assign w1607 = ~w1604 & ~w1606;
assign w1608 = w754 & ~w1370;
assign w1609 = (w1608 & w1529) | (w1608 & w39847) | (w1529 & w39847);
assign w1610 = w754 & w1370;
assign w1611 = ~w1529 & w39848;
assign w1612 = ~w1609 & ~w1611;
assign w1613 = ~w1391 & ~w1418;
assign w1614 = w1380 & w50934;
assign w1615 = (w1613 & ~w1380) | (w1613 & w50935) | (~w1380 & w50935);
assign w1616 = ~w1614 & ~w1615;
assign w1617 = w493 & ~w1390;
assign w1618 = (w1617 & w1529) | (w1617 & w39849) | (w1529 & w39849);
assign w1619 = w493 & ~w1616;
assign w1620 = ~w1529 & w39850;
assign w1621 = ~w1618 & ~w1620;
assign w1622 = w1607 & w1612;
assign w1623 = w1621 & w1622;
assign w1624 = ~w1600 & w1623;
assign w1625 = ~w1595 & w1624;
assign w1626 = w1445 & w1453;
assign w1627 = ~w1395 & w50936;
assign w1628 = (w1626 & w1395) | (w1626 & w50937) | (w1395 & w50937);
assign w1629 = ~w1627 & ~w1628;
assign w1630 = w1275 & ~w1411;
assign w1631 = ~w1275 & w1411;
assign w1632 = ~w1630 & ~w1631;
assign w1633 = (w43947 & w50938) | (w43947 & w50939) | (w50938 & w50939);
assign w1634 = (~w43947 & w50940) | (~w43947 & w50941) | (w50940 & w50941);
assign w1635 = ~w1633 & ~w1634;
assign w1636 = w400 & w1635;
assign w1637 = (w1390 & w1529) | (w1390 & w39851) | (w1529 & w39851);
assign w1638 = ~w1529 & w39852;
assign w1639 = ~w1637 & ~w1638;
assign w1640 = ~w493 & ~w1639;
assign w1641 = ~w612 & ~w1350;
assign w1642 = (w1641 & w1529) | (w1641 & w39853) | (w1529 & w39853);
assign w1643 = ~w612 & w1350;
assign w1644 = ~w1529 & w39854;
assign w1645 = ~w1642 & ~w1644;
assign w1646 = w1621 & ~w1645;
assign w1647 = ~w1640 & ~w1646;
assign w1648 = ~w1636 & w1647;
assign w1649 = ~w1625 & w1648;
assign w1650 = ~w1448 & ~w1456;
assign w1651 = ~w1427 & ~w1438;
assign w1652 = w1650 & w1651;
assign w1653 = (w1652 & w1477) | (w1652 & w39855) | (w1477 & w39855);
assign w1654 = ~w1529 & w1653;
assign w1655 = ~w252 & w1432;
assign w1656 = (w1655 & w1529) | (w1655 & w39856) | (w1529 & w39856);
assign w1657 = ~w252 & ~w1432;
assign w1658 = ~w1529 & w39857;
assign w1659 = ~w1656 & ~w1658;
assign w1660 = ~w1462 & ~w1479;
assign w1661 = ~w1440 & w1650;
assign w1662 = w1660 & ~w1661;
assign w1663 = ~w1660 & w1661;
assign w1664 = ~w1662 & ~w1663;
assign w1665 = ~w57 & w1461;
assign w1666 = (w1665 & w1529) | (w1665 & w39858) | (w1529 & w39858);
assign w1667 = ~w57 & w1664;
assign w1668 = w1541 & w1667;
assign w1669 = ~w1666 & ~w1668;
assign w1670 = w1659 & w1669;
assign w1671 = ~w400 & ~w1635;
assign w1672 = ~w400 & w52139;
assign w1673 = (w1395 & w50942) | (w1395 & w50943) | (w50942 & w50943);
assign w1674 = ~w1672 & ~w1673;
assign w1675 = (w1465 & w50944) | (w1465 & w50945) | (w50944 & w50945);
assign w1676 = w351 & w1435;
assign w1677 = (w1676 & w1529) | (w1676 & w43950) | (w1529 & w43950);
assign w1678 = w351 & ~w1435;
assign w1679 = ~w1529 & w43951;
assign w1680 = ~w1677 & ~w1679;
assign w1681 = w1670 & w50946;
assign w1682 = (w1681 & w1625) | (w1681 & w43952) | (w1625 & w43952);
assign w1683 = ~w1461 & ~w1541;
assign w1684 = w1541 & ~w1664;
assign w1685 = ~w1683 & ~w1684;
assign w1686 = (w57 & w1684) | (w57 & w50947) | (w1684 & w50947);
assign w1687 = ~w351 & ~w1435;
assign w1688 = (w1687 & w1529) | (w1687 & w43953) | (w1529 & w43953);
assign w1689 = ~w351 & w1435;
assign w1690 = ~w1529 & w43954;
assign w1691 = ~w1688 & ~w1690;
assign w1692 = w252 & ~w1432;
assign w1693 = (w1692 & w1529) | (w1692 & w39859) | (w1529 & w39859);
assign w1694 = w252 & w1432;
assign w1695 = ~w1529 & w39860;
assign w1696 = ~w1693 & ~w1695;
assign w1697 = w1691 & w1696;
assign w1698 = w1670 & ~w1697;
assign w1699 = ~w1686 & ~w1698;
assign w1700 = w1472 & w50948;
assign w1701 = (w1700 & ~w1541) | (w1700 & w39861) | (~w1541 & w39861);
assign w1702 = (~w80 & ~w1472) | (~w80 & w50949) | (~w1472 & w50949);
assign w1703 = w1541 & w39862;
assign w1704 = ~w1701 & ~w1703;
assign w1705 = ~w1698 & w50950;
assign w1706 = (w1549 & w1682) | (w1549 & w47005) | (w1682 & w47005);
assign w1707 = w126 & ~w1497;
assign w1708 = ~w1491 & w51484;
assign w1709 = (w1465 & w50951) | (w1465 & w50952) | (w50951 & w50952);
assign w1710 = ~w1510 & ~w1708;
assign w1711 = w1710 & w52140;
assign w1712 = ~w1709 & ~w1711;
assign w1713 = (w1465 & w50953) | (w1465 & w50954) | (w50953 & w50954);
assign w1714 = ~w1529 & w1713;
assign w1715 = w1712 & ~w1714;
assign w1716 = ~w1493 & w1529;
assign w1717 = w1715 & ~w1716;
assign w1718 = ~w1504 & w52141;
assign w1719 = (w1465 & w50956) | (w1465 & w50957) | (w50956 & w50957);
assign w1720 = w50958 & w52141;
assign w1721 = ~w1719 & ~w1720;
assign w1722 = (w1715 & w50959) | (w1715 & w50960) | (w50959 & w50960);
assign w1723 = w3 & ~w1540;
assign w1724 = ~w1723 & w50961;
assign w1725 = w1699 & w1724;
assign w1726 = w1699 & w50962;
assign w1727 = ~w3 & w1540;
assign w1728 = (w1465 & w50963) | (w1465 & w50964) | (w50963 & w50964);
assign w1729 = ~w42 & ~w1728;
assign w1730 = w1715 & w39865;
assign w1731 = ~w1727 & ~w1730;
assign w1732 = ~w1549 & ~w1723;
assign w1733 = w1731 & ~w1732;
assign w1734 = w1722 & ~w1733;
assign w1735 = ~w1726 & ~w1734;
assign w1736 = w1699 & w50965;
assign w1737 = w1725 & w1649;
assign w1738 = w1735 & ~w1737;
assign w1739 = w39866 & w50966;
assign w1740 = w39867 & w50967;
assign w1741 = ~w1739 & ~w1740;
assign w1742 = w42 & w1540;
assign w1743 = ~w1741 & w1742;
assign w1744 = w42 & ~w1540;
assign w1745 = w1741 & w1744;
assign w1746 = ~w1743 & ~w1745;
assign w1747 = ~w1682 & w47006;
assign w1748 = w1549 & w1704;
assign w1749 = (~w1748 & w1682) | (~w1748 & w47007) | (w1682 & w47007);
assign w1750 = (w1473 & ~w1541) | (w1473 & w50968) | (~w1541 & w50968);
assign w1751 = w1541 & w50969;
assign w1752 = ~w1750 & ~w1751;
assign w1753 = ~w1738 & w1752;
assign w1754 = ~w1747 & ~w1749;
assign w1755 = w1738 & w1754;
assign w1756 = ~w1753 & ~w1755;
assign w1757 = w3 & w1756;
assign w1758 = w1561 & ~w1573;
assign w1759 = (w1758 & w1733) | (w1758 & w39868) | (w1733 & w39868);
assign w1760 = ~w1726 & w1759;
assign w1761 = ~w1737 & w1760;
assign w1762 = ~w945 & ~w1569;
assign w1763 = (w1762 & ~w1760) | (w1762 & w39869) | (~w1760 & w39869);
assign w1764 = ~w945 & w1569;
assign w1765 = w1760 & w39870;
assign w1766 = ~w1763 & ~w1765;
assign w1767 = ~w1509 & w52142;
assign w1768 = a[101] & ~w1767;
assign w1769 = ~a[101] & w1767;
assign w1770 = ~w1768 & ~w1769;
assign w1771 = ~a[101] & w1555;
assign w1772 = (~w1553 & ~w1557) | (~w1553 & w50971) | (~w1557 & w50971);
assign w1773 = ~w1509 & w52143;
assign w1774 = w1772 & ~w1541;
assign w1775 = ~w1773 & ~w1774;
assign w1776 = w1120 & ~w1770;
assign w1777 = (w1776 & ~w1735) | (w1776 & w39871) | (~w1735 & w39871);
assign w1778 = ~w1773 & w50972;
assign w1779 = w1735 & w39872;
assign w1780 = ~w1777 & ~w1779;
assign w1781 = w1766 & ~w1780;
assign w1782 = w945 & w1569;
assign w1783 = (w1782 & ~w1760) | (w1782 & w39873) | (~w1760 & w39873);
assign w1784 = w945 & ~w1569;
assign w1785 = w1760 & w39874;
assign w1786 = ~w1783 & ~w1785;
assign w1787 = w1588 & ~w1599;
assign w1788 = ~w1570 & ~w1573;
assign w1789 = w1787 & ~w1788;
assign w1790 = ~w1787 & w1788;
assign w1791 = ~w1789 & ~w1790;
assign w1792 = ~w754 & ~w1598;
assign w1793 = (w1792 & ~w1735) | (w1792 & w39875) | (~w1735 & w39875);
assign w1794 = ~w754 & w1791;
assign w1795 = w1735 & w39876;
assign w1796 = ~w1793 & ~w1795;
assign w1797 = w1786 & w1796;
assign w1798 = ~w1781 & w1797;
assign w1799 = (~w1770 & ~w1735) | (~w1770 & w39877) | (~w1735 & w39877);
assign w1800 = w1735 & w39878;
assign w1801 = ~w1799 & ~w1800;
assign w1802 = ~w1120 & w1801;
assign w1803 = w1766 & ~w1802;
assign w1804 = ~a[96] & ~a[97];
assign w1805 = ~a[98] & w1804;
assign w1806 = ~w1509 & w52144;
assign w1807 = a[98] & ~a[99];
assign w1808 = (w1807 & w1733) | (w1807 & w39879) | (w1733 & w39879);
assign w1809 = ~w1726 & w1808;
assign w1810 = (~w1806 & ~w1809) | (~w1806 & w39880) | (~w1809 & w39880);
assign w1811 = ~w1805 & ~w1541;
assign w1812 = ~a[99] & ~w1811;
assign w1813 = (w1812 & ~w1735) | (w1812 & w39881) | (~w1735 & w39881);
assign w1814 = a[99] & ~w1811;
assign w1815 = w1735 & w39882;
assign w1816 = ~w1813 & ~w1815;
assign w1817 = (w1320 & ~w1816) | (w1320 & w43955) | (~w1816 & w43955);
assign w1818 = (w39880 & w50974) | (w39880 & w50975) | (w50974 & w50975);
assign w1819 = w1816 & w1818;
assign w1820 = a[100] & ~w1550;
assign w1821 = a[100] & ~w1541;
assign w1822 = ~w1767 & ~w1821;
assign w1823 = ~w1738 & w1822;
assign w1824 = ~w1551 & ~w1820;
assign w1825 = w1738 & w1824;
assign w1826 = ~w1823 & ~w1825;
assign w1827 = ~w1819 & ~w1826;
assign w1828 = ~w1817 & ~w1827;
assign w1829 = w1803 & w1828;
assign w1830 = (w1798 & ~w1828) | (w1798 & w43956) | (~w1828 & w43956);
assign w1831 = (w1659 & w1680) | (w1659 & w39883) | (w1680 & w39883);
assign w1832 = ~w1697 & w1831;
assign w1833 = w1648 & ~w1832;
assign w1834 = w1671 & w1697;
assign w1835 = w1831 & ~w1834;
assign w1836 = ~w1625 & w1833;
assign w1837 = w1669 & ~w1686;
assign w1838 = ~w1836 & w43957;
assign w1839 = (w1837 & w1836) | (w1837 & w43958) | (w1836 & w43958);
assign w1840 = ~w1838 & ~w1839;
assign w1841 = w1685 & ~w1738;
assign w1842 = w1738 & w1840;
assign w1843 = ~w1841 & ~w1842;
assign w1844 = (w80 & w1842) | (w80 & w50976) | (w1842 & w50976);
assign w1845 = ~w1636 & ~w1671;
assign w1846 = (w1845 & w1625) | (w1845 & w47008) | (w1625 & w47008);
assign w1847 = ~w1625 & w47009;
assign w1848 = ~w1846 & ~w1847;
assign w1849 = w1635 & ~w1738;
assign w1850 = w1738 & w1848;
assign w1851 = ~w1849 & ~w1850;
assign w1852 = w351 & w1851;
assign w1853 = w1621 & ~w1640;
assign w1854 = (w1612 & ~w1599) | (w1612 & w47010) | (~w1599 & w47010);
assign w1855 = ~w1595 & w1854;
assign w1856 = (w47012 & w50977) | (w47012 & w50978) | (w50977 & w50978);
assign w1857 = w1853 & w52145;
assign w1858 = ~w1639 & ~w1738;
assign w1859 = w1738 & w39884;
assign w1860 = ~w1858 & ~w1859;
assign w1861 = ~w400 & w1860;
assign w1862 = ~w1852 & ~w1861;
assign w1863 = ~w1844 & w1862;
assign w1864 = w1598 & ~w1738;
assign w1865 = w1738 & ~w1791;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = w754 & ~w1866;
assign w1868 = (~w1599 & ~w1589) | (~w1599 & w50979) | (~w1589 & w50979);
assign w1869 = w1623 & w1868;
assign w1870 = w1736 & ~w1869;
assign w1871 = w1735 & ~w1870;
assign w1872 = w754 & ~w1871;
assign w1873 = (~w1868 & w1733) | (~w1868 & w50980) | (w1733 & w50980);
assign w1874 = ~w1726 & w1873;
assign w1875 = ~w1737 & w1874;
assign w1876 = ~w1594 & w1612;
assign w1877 = (w612 & w1594) | (w612 & w50981) | (w1594 & w50981);
assign w1878 = (w1877 & w1872) | (w1877 & w39885) | (w1872 & w39885);
assign w1879 = ~w1594 & w50982;
assign w1880 = ~w1872 & w39886;
assign w1881 = ~w1878 & ~w1880;
assign w1882 = ~w1867 & w1881;
assign w1883 = ~w1595 & w47013;
assign w1884 = w1736 & ~w1883;
assign w1885 = w1735 & ~w1884;
assign w1886 = ~w612 & ~w1885;
assign w1887 = ~w1734 & w1855;
assign w1888 = ~w1726 & w1887;
assign w1889 = ~w1737 & w1888;
assign w1890 = ~w1886 & ~w1889;
assign w1891 = w1607 & w1645;
assign w1892 = w493 & w1891;
assign w1893 = (w1892 & w1886) | (w1892 & w39887) | (w1886 & w39887);
assign w1894 = w493 & ~w1891;
assign w1895 = ~w1886 & w39888;
assign w1896 = ~w1893 & ~w1895;
assign w1897 = w1882 & w1896;
assign w1898 = w1863 & w1897;
assign w1899 = ~w1830 & w1898;
assign w1900 = ~w1842 & w50983;
assign w1901 = w1680 & w1691;
assign w1902 = ~w1671 & w1901;
assign w1903 = (w1902 & w1625) | (w1902 & w47014) | (w1625 & w47014);
assign w1904 = w1691 & ~w1903;
assign w1905 = ~w252 & w1691;
assign w1906 = ~w1903 & w1905;
assign w1907 = w1738 & ~w1906;
assign w1908 = w1432 & ~w1654;
assign w1909 = ~w1432 & w1654;
assign w1910 = ~w1908 & ~w1909;
assign w1911 = w57 & w1910;
assign w1912 = (w1911 & w39889) | (w1911 & ~w1907) | (w39889 & ~w1907);
assign w1913 = w57 & ~w1910;
assign w1914 = w1738 & w47015;
assign w1915 = ~w1912 & ~w1914;
assign w1916 = ~w1900 & w1915;
assign w1917 = ~w351 & ~w1851;
assign w1918 = (~w1671 & w1625) | (~w1671 & w43960) | (w1625 & w43960);
assign w1919 = ~w1901 & ~w1918;
assign w1920 = ~w1903 & ~w1919;
assign w1921 = w1735 & ~w1920;
assign w1922 = ~w1529 & w50984;
assign w1923 = (~w1435 & w1529) | (~w1435 & w50985) | (w1529 & w50985);
assign w1924 = ~w1922 & ~w1923;
assign w1925 = (w1924 & ~w1738) | (w1924 & w39891) | (~w1738 & w39891);
assign w1926 = ~w1921 & ~w1925;
assign w1927 = ~w1925 & w47016;
assign w1928 = ~w1917 & ~w1927;
assign w1929 = w1916 & w1928;
assign w1930 = w400 & ~w1860;
assign w1931 = ~w493 & w1891;
assign w1932 = (w1931 & ~w1888) | (w1931 & w39892) | (~w1888 & w39892);
assign w1933 = ~w1886 & w1932;
assign w1934 = ~w493 & ~w1891;
assign w1935 = ~w1891 & w50986;
assign w1936 = ~w1885 & w1935;
assign w1937 = w1888 & w39893;
assign w1938 = ~w1936 & ~w1937;
assign w1939 = ~w1933 & w1938;
assign w1940 = (~w612 & w1594) | (~w612 & w50987) | (w1594 & w50987);
assign w1941 = (w1940 & ~w1874) | (w1940 & w39894) | (~w1874 & w39894);
assign w1942 = ~w1872 & w1941;
assign w1943 = ~w1594 & w50988;
assign w1944 = w50988 & w51486;
assign w1945 = ~w1871 & w1944;
assign w1946 = w1874 & w39895;
assign w1947 = ~w1945 & ~w1946;
assign w1948 = ~w1942 & w1947;
assign w1949 = w1939 & w1948;
assign w1950 = w1896 & ~w1949;
assign w1951 = (~w1930 & w1949) | (~w1930 & w39896) | (w1949 & w39896);
assign w1952 = w1863 & ~w1951;
assign w1953 = w1929 & ~w1952;
assign w1954 = ~w1899 & w1953;
assign w1955 = ~w3 & ~w1756;
assign w1956 = (~w252 & w1925) | (~w252 & w47017) | (w1925 & w47017);
assign w1957 = ~w57 & ~w1910;
assign w1958 = (w1957 & ~w1907) | (w1957 & w39897) | (~w1907 & w39897);
assign w1959 = ~w57 & w1910;
assign w1960 = w1907 & w39898;
assign w1961 = ~w1958 & ~w1960;
assign w1962 = ~w1956 & w1961;
assign w1963 = w1916 & ~w1962;
assign w1964 = ~w1963 & w50989;
assign w1965 = ~w1746 & w52146;
assign w1966 = ~w1540 & ~w1741;
assign w1967 = w1540 & w1741;
assign w1968 = ~w1966 & ~w1967;
assign w1969 = (w1954 & w50990) | (w1954 & w50991) | (w50990 & w50991);
assign w1970 = ~w1718 & ~w1728;
assign w1971 = w1715 & w50993;
assign w1972 = ~w3 & ~w1706;
assign w1973 = w1540 & ~w1717;
assign w1974 = (w1973 & ~w1738) | (w1973 & w51487) | (~w1738 & w51487);
assign w1975 = (w1682 & w51544) | (w1682 & w51545) | (w51544 & w51545);
assign w1976 = (~w1974 & w1968) | (~w1974 & w50994) | (w1968 & w50994);
assign w1977 = w1746 & w1976;
assign w1978 = ~w1977 & w52146;
assign w1979 = w42 & ~w1965;
assign w1980 = ~w1969 & ~w1978;
assign w1981 = ~w1979 & ~w1980;
assign w1982 = ~w42 & ~w1540;
assign w1983 = ~w1741 & w1982;
assign w1984 = ~w42 & w1540;
assign w1985 = w1741 & w1984;
assign w1986 = ~w1983 & ~w1985;
assign w1987 = ~w1955 & w1986;
assign w1988 = ~w1963 & w1987;
assign w1989 = ~w1844 & ~w1929;
assign w1990 = w1988 & w1989;
assign w1991 = (~w42 & ~w1715) | (~w42 & w50995) | (~w1715 & w50995);
assign w1992 = w1991 & w52342;
assign w1993 = ~w42 & w1971;
assign w1994 = (w1682 & w51488) | (w1682 & w51489) | (w51488 & w51489);
assign w1995 = ~w1992 & ~w1994;
assign w1996 = w1746 & w1995;
assign w1997 = w1746 & w50996;
assign w1998 = ~w1990 & w1997;
assign w1999 = ~w1899 & ~w1952;
assign w2000 = w1998 & w1999;
assign w2001 = w1844 & w1929;
assign w2002 = w1988 & ~w2001;
assign w2003 = w1757 & w1986;
assign w2004 = w1996 & ~w2003;
assign w2005 = ~w2002 & w2004;
assign w2006 = ~w2000 & ~w2005;
assign w2007 = ~w3 & w1929;
assign w2008 = ~w1952 & w2007;
assign w2009 = ~w1899 & w2008;
assign w2010 = ~w1963 & w50997;
assign w2011 = ~w1954 & w2010;
assign w2012 = (~w3 & w1963) | (~w3 & w50998) | (w1963 & w50998);
assign w2013 = ~w2009 & ~w2012;
assign w2014 = ~w2011 & w2013;
assign w2015 = w2006 & w2014;
assign w2016 = w42 & w1756;
assign w2017 = (w2016 & ~w2006) | (w2016 & w43961) | (~w2006 & w43961);
assign w2018 = ~w1746 & ~w1756;
assign w2019 = w2006 & w43962;
assign w2020 = ~w2017 & ~w2019;
assign w2021 = ~w1981 & w2020;
assign w2022 = ~w1927 & ~w1956;
assign w2023 = ~w1861 & w1896;
assign w2024 = w1882 & w2023;
assign w2025 = ~w1852 & ~w1917;
assign w2026 = w2024 & w2025;
assign w2027 = ~w1830 & w2026;
assign w2028 = (~w1917 & w1951) | (~w1917 & w47019) | (w1951 & w47019);
assign w2029 = (w2022 & w2027) | (w2022 & w47020) | (w2027 & w47020);
assign w2030 = ~w2027 & w47021;
assign w2031 = ~w2029 & ~w2030;
assign w2032 = w2006 & w2031;
assign w2033 = (w1926 & w2000) | (w1926 & w50999) | (w2000 & w50999);
assign w2034 = ~w2032 & ~w2033;
assign w2035 = (w57 & w2032) | (w57 & w51000) | (w2032 & w51000);
assign w2036 = ~w1897 & ~w1950;
assign w2037 = (w1798 & w1949) | (w1798 & w39899) | (w1949 & w39899);
assign w2038 = ~w1829 & w2037;
assign w2039 = ~w1861 & ~w1930;
assign w2040 = ~w2038 & w43963;
assign w2041 = (w2039 & w2038) | (w2039 & w43964) | (w2038 & w43964);
assign w2042 = ~w2040 & ~w2041;
assign w2043 = ~w351 & ~w1860;
assign w2044 = (w2043 & w2000) | (w2043 & w39900) | (w2000 & w39900);
assign w2045 = ~w351 & ~w2042;
assign w2046 = w2006 & w2045;
assign w2047 = ~w2044 & ~w2046;
assign w2048 = ~w1830 & w2024;
assign w2049 = (~w2025 & w1951) | (~w2025 & w39901) | (w1951 & w39901);
assign w2050 = ~w2048 & w2049;
assign w2051 = ~w1951 & w39902;
assign w2052 = ~w2027 & ~w2051;
assign w2053 = ~w2050 & w2052;
assign w2054 = w252 & ~w1851;
assign w2055 = (w2054 & w2000) | (w2054 & w39903) | (w2000 & w39903);
assign w2056 = w252 & w2053;
assign w2057 = w2006 & w2056;
assign w2058 = ~w2055 & ~w2057;
assign w2059 = w2047 & w2058;
assign w2060 = (~w57 & w1925) | (~w57 & w51001) | (w1925 & w51001);
assign w2061 = (~w57 & w2002) | (~w57 & w39904) | (w2002 & w39904);
assign w2062 = (~w2060 & w2000) | (~w2060 & w39905) | (w2000 & w39905);
assign w2063 = ~w2032 & ~w2062;
assign w2064 = ~w252 & w1851;
assign w2065 = (w2064 & w2000) | (w2064 & w39906) | (w2000 & w39906);
assign w2066 = ~w252 & ~w2053;
assign w2067 = w2006 & w2066;
assign w2068 = ~w2065 & ~w2067;
assign w2069 = ~w2063 & w2068;
assign w2070 = ~w2059 & w2069;
assign w2071 = ~w2035 & ~w2070;
assign w2072 = ~w1844 & ~w1900;
assign w2073 = w1862 & ~w1956;
assign w2074 = w1897 & w2073;
assign w2075 = ~w1830 & w2074;
assign w2076 = ~w1951 & w2073;
assign w2077 = (~w1956 & w1917) | (~w1956 & w51002) | (w1917 & w51002);
assign w2078 = (w1915 & w1928) | (w1915 & w39907) | (w1928 & w39907);
assign w2079 = ~w2076 & w2078;
assign w2080 = ~w2075 & w2079;
assign w2081 = (~w2072 & w2080) | (~w2072 & w39908) | (w2080 & w39908);
assign w2082 = w2006 & w2081;
assign w2083 = (~w1843 & w2000) | (~w1843 & w39909) | (w2000 & w39909);
assign w2084 = ~w2080 & w39910;
assign w2085 = ~w2000 & w43965;
assign w2086 = ~w2083 & ~w2085;
assign w2087 = (w3 & ~w2006) | (w3 & w39911) | (~w2006 & w39911);
assign w2088 = w2086 & w2087;
assign w2089 = w1915 & w1961;
assign w2090 = ~w2076 & ~w2077;
assign w2091 = ~w2075 & w2090;
assign w2092 = w2089 & ~w2091;
assign w2093 = ~w2089 & w2091;
assign w2094 = (w1915 & ~w1961) | (w1915 & w51003) | (~w1961 & w51003);
assign w2095 = (~w2094 & w2000) | (~w2094 & w39912) | (w2000 & w39912);
assign w2096 = ~w80 & w2095;
assign w2097 = (~w80 & ~w2091) | (~w80 & w51004) | (~w2091 & w51004);
assign w2098 = w43966 & w51005;
assign w2099 = ~w2096 & ~w2098;
assign w2100 = ~w2088 & w2099;
assign w2101 = w2021 & w2100;
assign w2102 = w2071 & w2101;
assign w2103 = (~w3 & ~w2086) | (~w3 & w39913) | (~w2086 & w39913);
assign w2104 = w1756 & ~w2015;
assign w2105 = ~w1756 & w2015;
assign w2106 = ~w2104 & ~w2105;
assign w2107 = ~w42 & w2106;
assign w2108 = ~w2103 & ~w2107;
assign w2109 = w80 & ~w2095;
assign w2110 = w43966 & w47022;
assign w2111 = w2109 & ~w2110;
assign w2112 = ~w2088 & w2111;
assign w2113 = w2108 & ~w2112;
assign w2114 = w1890 & ~w1891;
assign w2115 = ~w1890 & w1891;
assign w2116 = ~w2114 & ~w2115;
assign w2117 = w1896 & w1939;
assign w2118 = w1803 & ~w1867;
assign w2119 = w1828 & w2118;
assign w2120 = (w1948 & w1798) | (w1948 & w43967) | (w1798 & w43967);
assign w2121 = (~w2119 & w43968) | (~w2119 & w43969) | (w43968 & w43969);
assign w2122 = (w39915 & w2119) | (w39915 & w43970) | (w2119 & w43970);
assign w2123 = ~w2121 & ~w2122;
assign w2124 = (w2116 & w2000) | (w2116 & w39916) | (w2000 & w39916);
assign w2125 = ~w2000 & w39917;
assign w2126 = ~w2124 & ~w2125;
assign w2127 = ~w400 & w2126;
assign w2128 = (w1860 & w2000) | (w1860 & w39918) | (w2000 & w39918);
assign w2129 = ~w2000 & w43971;
assign w2130 = ~w2128 & ~w2129;
assign w2131 = (w351 & w2129) | (w351 & w39919) | (w2129 & w39919);
assign w2132 = ~w2127 & ~w2131;
assign w2133 = w2069 & w2132;
assign w2134 = (w2021 & ~w2108) | (w2021 & w39920) | (~w2108 & w39920);
assign w2135 = w2071 & w43972;
assign w2136 = ~w2134 & ~w2135;
assign w2137 = a[99] & ~w1738;
assign w2138 = ~a[99] & w1738;
assign w2139 = ~w2137 & ~w2138;
assign w2140 = a[98] & w1738;
assign w2141 = (w2140 & w2000) | (w2140 & w39921) | (w2000 & w39921);
assign w2142 = ~w1806 & ~w1811;
assign w2143 = ~w2000 & w39922;
assign w2144 = ~w2141 & ~w2143;
assign w2145 = ~w2139 & ~w2144;
assign w2146 = w2139 & w2144;
assign w2147 = ~w2145 & ~w2146;
assign w2148 = ~w1320 & w2147;
assign w2149 = (~a[97] & w2002) | (~a[97] & w39923) | (w2002 & w39923);
assign w2150 = ~w2000 & w2149;
assign w2151 = a[97] & ~w1952;
assign w2152 = ~w1899 & w2151;
assign w2153 = w1998 & w2152;
assign w2154 = a[97] & w2004;
assign w2155 = ~w2002 & w2154;
assign w2156 = ~a[94] & ~a[95];
assign w2157 = ~a[96] & w2156;
assign w2158 = ~w1738 & ~w2157;
assign w2159 = ~w2155 & ~w2158;
assign w2160 = ~w2153 & w2159;
assign w2161 = ~w2150 & w2160;
assign w2162 = w1738 & w2157;
assign w2163 = a[96] & ~a[97];
assign w2164 = (w2163 & w2002) | (w2163 & w39924) | (w2002 & w39924);
assign w2165 = (~w2162 & w2000) | (~w2162 & w39925) | (w2000 & w39925);
assign w2166 = (w1541 & w2161) | (w1541 & w39926) | (w2161 & w39926);
assign w2167 = (~w1541 & ~w1738) | (~w1541 & w51006) | (~w1738 & w51006);
assign w2168 = (w2167 & w2000) | (w2167 & w39927) | (w2000 & w39927);
assign w2169 = ~w2161 & w2168;
assign w2170 = ~a[98] & ~w1738;
assign w2171 = a[98] & ~w1804;
assign w2172 = ~w1805 & ~w2171;
assign w2173 = ~w2140 & ~w2170;
assign w2174 = (w2173 & w2000) | (w2173 & w39928) | (w2000 & w39928);
assign w2175 = ~w2000 & w39929;
assign w2176 = ~w2174 & ~w2175;
assign w2177 = ~w2169 & w2176;
assign w2178 = ~w2166 & ~w2177;
assign w2179 = w1320 & ~w2139;
assign w2180 = ~w2144 & w2179;
assign w2181 = w1320 & w2139;
assign w2182 = w2144 & w2181;
assign w2183 = ~w2180 & ~w2182;
assign w2184 = w2178 & w2183;
assign w2185 = ~w2148 & ~w2184;
assign w2186 = (w612 & w2119) | (w612 & w39930) | (w2119 & w39930);
assign w2187 = ~w2119 & w39931;
assign w2188 = ~w2186 & ~w2187;
assign w2189 = ~w2005 & ~w2188;
assign w2190 = ~w2000 & w2189;
assign w2191 = ~w1872 & w51007;
assign w2192 = (w1876 & w1872) | (w1876 & w51008) | (w1872 & w51008);
assign w2193 = ~w2191 & ~w2192;
assign w2194 = w493 & w2193;
assign w2195 = ~w2190 & w2194;
assign w2196 = w493 & ~w2193;
assign w2197 = w2190 & w2196;
assign w2198 = ~w2195 & ~w2197;
assign w2199 = w400 & ~w2123;
assign w2200 = ~w2000 & w43973;
assign w2201 = w400 & w2116;
assign w2202 = (w2201 & w2000) | (w2201 & w39932) | (w2000 & w39932);
assign w2203 = ~w2200 & ~w2202;
assign w2204 = ~w2198 & w2203;
assign w2205 = w1780 & ~w1802;
assign w2206 = ~w1828 & w2205;
assign w2207 = (~w1802 & w1828) | (~w1802 & w39933) | (w1828 & w39933);
assign w2208 = ~w945 & w2207;
assign w2209 = w945 & ~w2207;
assign w2210 = ~w2208 & ~w2209;
assign w2211 = ~w2005 & ~w2210;
assign w2212 = ~w2000 & w2211;
assign w2213 = w1569 & ~w1761;
assign w2214 = ~w1569 & w1761;
assign w2215 = ~w2213 & ~w2214;
assign w2216 = w754 & w2215;
assign w2217 = ~w2212 & w2216;
assign w2218 = w754 & ~w2215;
assign w2219 = w2212 & w2218;
assign w2220 = ~w2217 & ~w2219;
assign w2221 = w1796 & ~w1867;
assign w2222 = ~w1781 & w1786;
assign w2223 = (w2222 & ~w1828) | (w2222 & w51009) | (~w1828 & w51009);
assign w2224 = w2221 & ~w2223;
assign w2225 = ~w2221 & w2223;
assign w2226 = ~w2224 & ~w2225;
assign w2227 = w612 & ~w1866;
assign w2228 = (w2227 & w2000) | (w2227 & w39934) | (w2000 & w39934);
assign w2229 = w612 & ~w2226;
assign w2230 = ~w2000 & w51463;
assign w2231 = ~w2228 & ~w2230;
assign w2232 = w2220 & w2231;
assign w2233 = w1828 & ~w2205;
assign w2234 = ~w2206 & ~w2233;
assign w2235 = ~w945 & w1801;
assign w2236 = (w2235 & w2000) | (w2235 & w39935) | (w2000 & w39935);
assign w2237 = ~w945 & w2234;
assign w2238 = ~w2000 & w39936;
assign w2239 = ~w2236 & ~w2238;
assign w2240 = ~w1817 & ~w1819;
assign w2241 = (w2240 & w2002) | (w2240 & w39937) | (w2002 & w39937);
assign w2242 = ~w2000 & w39938;
assign w2243 = ~w1120 & ~w2242;
assign w2244 = (w1826 & w2000) | (w1826 & w47023) | (w2000 & w47023);
assign w2245 = w2243 & ~w2244;
assign w2246 = w2239 & ~w2245;
assign w2247 = w2232 & w2246;
assign w2248 = ~w2204 & w2247;
assign w2249 = ~w2185 & w2248;
assign w2250 = w1120 & w1826;
assign w2251 = (w2250 & w2000) | (w2250 & w39939) | (w2000 & w39939);
assign w2252 = w1120 & ~w1826;
assign w2253 = ~w2000 & w39940;
assign w2254 = ~w2251 & ~w2253;
assign w2255 = ~w754 & ~w2215;
assign w2256 = ~w2212 & w2255;
assign w2257 = ~w754 & w2215;
assign w2258 = w2212 & w2257;
assign w2259 = ~w2256 & ~w2258;
assign w2260 = w945 & ~w1801;
assign w2261 = (w2260 & w2000) | (w2260 & w39941) | (w2000 & w39941);
assign w2262 = w945 & ~w2234;
assign w2263 = ~w2000 & w39942;
assign w2264 = ~w2261 & ~w2263;
assign w2265 = w2259 & w2264;
assign w2266 = w2239 & ~w2254;
assign w2267 = w2265 & ~w2266;
assign w2268 = ~w493 & ~w2193;
assign w2269 = ~w2190 & w2268;
assign w2270 = ~w493 & w2193;
assign w2271 = w2190 & w2270;
assign w2272 = ~w2269 & ~w2271;
assign w2273 = ~w612 & w1866;
assign w2274 = (w2273 & w2000) | (w2273 & w39943) | (w2000 & w39943);
assign w2275 = ~w612 & w2226;
assign w2276 = ~w2000 & w51464;
assign w2277 = ~w2274 & ~w2276;
assign w2278 = w2272 & w2277;
assign w2279 = (w2203 & w2278) | (w2203 & w2204) | (w2278 & w2204);
assign w2280 = ~w2204 & w2232;
assign w2281 = ~w2267 & w2280;
assign w2282 = w2279 & ~w2281;
assign w2283 = w2102 & w2282;
assign w2284 = ~w2249 & w2283;
assign w2285 = w2136 & ~w2284;
assign w2286 = (w1851 & w2000) | (w1851 & w51010) | (w2000 & w51010);
assign w2287 = w2006 & ~w2053;
assign w2288 = ~w2286 & ~w2287;
assign w2289 = w2132 & ~w2204;
assign w2290 = (w2289 & w2281) | (w2289 & w39944) | (w2281 & w39944);
assign w2291 = w2247 & w2289;
assign w2292 = ~w2185 & w2291;
assign w2293 = ~w2292 & w39945;
assign w2294 = w2068 & w2293;
assign w2295 = w2058 & w2068;
assign w2296 = ~w2292 & w39946;
assign w2297 = ~w2295 & ~w2296;
assign w2298 = ~w2285 & ~w2288;
assign w2299 = ~w2294 & ~w2297;
assign w2300 = w2285 & w2299;
assign w2301 = ~w2298 & ~w2300;
assign w2302 = ~w2000 & w51011;
assign w2303 = (a[96] & w2000) | (a[96] & w51012) | (w2000 & w51012);
assign w2304 = ~w2302 & ~w2303;
assign w2305 = a[96] & ~w2156;
assign w2306 = ~w2157 & ~w2305;
assign w2307 = w1738 & w2304;
assign w2308 = ~w2285 & w2307;
assign w2309 = w1738 & w2306;
assign w2310 = w2285 & w2309;
assign w2311 = ~w2308 & ~w2310;
assign w2312 = ~a[92] & ~a[93];
assign w2313 = ~a[94] & w2312;
assign w2314 = ~w2000 & w51013;
assign w2315 = (~w2313 & w2000) | (~w2313 & w51014) | (w2000 & w51014);
assign w2316 = (~w2156 & ~w2315) | (~w2156 & w51015) | (~w2315 & w51015);
assign w2317 = ~a[95] & ~w2315;
assign w2318 = ~w2314 & ~w2317;
assign w2319 = ~w2285 & w2318;
assign w2320 = ~w2314 & ~w2316;
assign w2321 = w2285 & w2320;
assign w2322 = ~w2319 & ~w2321;
assign w2323 = ~w1738 & ~w2304;
assign w2324 = ~w2285 & w2323;
assign w2325 = ~w1738 & ~w2306;
assign w2326 = w2285 & w2325;
assign w2327 = ~w2324 & ~w2326;
assign w2328 = w2322 & w2327;
assign w2329 = (w1541 & w2328) | (w1541 & w39947) | (w2328 & w39947);
assign w2330 = ~w2166 & ~w2169;
assign w2331 = (w2176 & ~w2285) | (w2176 & w39948) | (~w2285 & w39948);
assign w2332 = w2285 & w39949;
assign w2333 = ~w2331 & ~w2332;
assign w2334 = w1320 & ~w2333;
assign w2335 = (w2133 & w2249) | (w2133 & w39950) | (w2249 & w39950);
assign w2336 = w2071 & ~w2335;
assign w2337 = w2020 & w51016;
assign w2338 = (w2337 & ~w2108) | (w2337 & w51017) | (~w2108 & w51017);
assign w2339 = (~w1738 & w2000) | (~w1738 & w51490) | (w2000 & w51490);
assign w2340 = ~w2000 & w51018;
assign w2341 = ~w2339 & ~w2340;
assign w2342 = (w2157 & w2339) | (w2157 & w51019) | (w2339 & w51019);
assign w2343 = ~w2339 & w51020;
assign w2344 = ~w2342 & ~w2343;
assign w2345 = ~w2284 & w43974;
assign w2346 = (a[97] & ~w2338) | (a[97] & w47024) | (~w2338 & w47024);
assign w2347 = ~w2345 & w2346;
assign w2348 = w2336 & w2338;
assign w2349 = w2347 & ~w2348;
assign w2350 = w2285 & w39951;
assign w2351 = ~w2070 & w51021;
assign w2352 = w2338 & w2351;
assign w2353 = ~w2335 & w2352;
assign w2354 = w2338 & w47025;
assign w2355 = ~w2353 & ~w2354;
assign w2356 = ~w2350 & w2355;
assign w2357 = ~w2349 & w2356;
assign w2358 = ~w2334 & ~w2357;
assign w2359 = ~w2329 & w2358;
assign w2360 = ~w1320 & w2333;
assign w2361 = ~w1541 & w2311;
assign w2362 = ~w2328 & w2361;
assign w2363 = ~w2334 & w2362;
assign w2364 = (~w2360 & ~w2362) | (~w2360 & w39952) | (~w2362 & w39952);
assign w2365 = ~w2359 & w2364;
assign w2366 = ~w2245 & w2254;
assign w2367 = ~w2284 & w43975;
assign w2368 = (w1120 & w2284) | (w1120 & w43976) | (w2284 & w43976);
assign w2369 = ~w2367 & ~w2368;
assign w2370 = w2366 & ~w2369;
assign w2371 = ~w2366 & w2369;
assign w2372 = ~w2370 & ~w2371;
assign w2373 = ~w945 & ~w2372;
assign w2374 = w2148 & w2178;
assign w2375 = w2285 & w39953;
assign w2376 = ~w2178 & ~w2183;
assign w2377 = (~w2376 & w2285) | (~w2376 & w39954) | (w2285 & w39954);
assign w2378 = ~w2375 & w2377;
assign w2379 = ~w1120 & ~w2378;
assign w2380 = ~w2373 & ~w2379;
assign w2381 = ~w2365 & w2380;
assign w2382 = w1120 & w2378;
assign w2383 = w945 & w2372;
assign w2384 = ~w2184 & w39955;
assign w2385 = (~w945 & w2384) | (~w945 & w47026) | (w2384 & w47026);
assign w2386 = ~w2384 & w47027;
assign w2387 = (w1801 & w2000) | (w1801 & w51022) | (w2000 & w51022);
assign w2388 = ~w2000 & w51023;
assign w2389 = ~w2387 & ~w2388;
assign w2390 = w2285 & w47028;
assign w2391 = (~w2389 & ~w2285) | (~w2389 & w47029) | (~w2285 & w47029);
assign w2392 = ~w2390 & ~w2391;
assign w2393 = ~w754 & w2392;
assign w2394 = ~w2383 & ~w2393;
assign w2395 = (w2382 & w2372) | (w2382 & w39957) | (w2372 & w39957);
assign w2396 = w2394 & ~w2395;
assign w2397 = ~w2127 & w2203;
assign w2398 = (w2247 & w2184) | (w2247 & w39958) | (w2184 & w39958);
assign w2399 = (w2278 & w2267) | (w2278 & w47030) | (w2267 & w47030);
assign w2400 = (w2198 & w2398) | (w2198 & w47031) | (w2398 & w47031);
assign w2401 = w2397 & ~w2400;
assign w2402 = ~w2397 & w2400;
assign w2403 = ~w2401 & ~w2402;
assign w2404 = w2285 & w2403;
assign w2405 = w2126 & ~w2285;
assign w2406 = (~w351 & w2285) | (~w351 & w47032) | (w2285 & w47032);
assign w2407 = ~w2404 & w2406;
assign w2408 = (w2277 & w2267) | (w2277 & w51024) | (w2267 & w51024);
assign w2409 = ~w2398 & w2408;
assign w2410 = ~w2284 & w43977;
assign w2411 = ~w2070 & w43978;
assign w2412 = w2282 & w2411;
assign w2413 = ~w2249 & w2412;
assign w2414 = (~w493 & w2135) | (~w493 & w39959) | (w2135 & w39959);
assign w2415 = w2020 & w51025;
assign w2416 = w2413 & w2415;
assign w2417 = ~w2414 & ~w2416;
assign w2418 = ~w2410 & w2417;
assign w2419 = w2198 & w2272;
assign w2420 = w400 & w2419;
assign w2421 = w2417 & w43979;
assign w2422 = w400 & ~w2419;
assign w2423 = (w2422 & ~w2417) | (w2422 & w43980) | (~w2417 & w43980);
assign w2424 = ~w2421 & ~w2423;
assign w2425 = ~w2407 & w2424;
assign w2426 = w2254 & w2264;
assign w2427 = ~w2184 & w39960;
assign w2428 = (w2264 & w2245) | (w2264 & w51026) | (w2245 & w51026);
assign w2429 = w2220 & ~w2428;
assign w2430 = (w2259 & w2427) | (w2259 & w47033) | (w2427 & w47033);
assign w2431 = (w612 & w2284) | (w612 & w43981) | (w2284 & w43981);
assign w2432 = w2285 & w2430;
assign w2433 = w2231 & w2277;
assign w2434 = w493 & w2433;
assign w2435 = ~w2432 & w43982;
assign w2436 = w493 & ~w2433;
assign w2437 = (w2436 & w2432) | (w2436 & w43983) | (w2432 & w43983);
assign w2438 = ~w2435 & ~w2437;
assign w2439 = ~w400 & w2419;
assign w2440 = (w2439 & ~w2417) | (w2439 & w43984) | (~w2417 & w43984);
assign w2441 = ~w400 & ~w2419;
assign w2442 = w2417 & w43985;
assign w2443 = ~w2440 & ~w2442;
assign w2444 = w2438 & w2443;
assign w2445 = w2425 & ~w2444;
assign w2446 = (~w754 & w2135) | (~w754 & w39961) | (w2135 & w39961);
assign w2447 = w2020 & w51027;
assign w2448 = w2413 & w2447;
assign w2449 = ~w2446 & ~w2448;
assign w2450 = ~w2427 & ~w2428;
assign w2451 = w2220 & w2259;
assign w2452 = ~w612 & ~w2451;
assign w2453 = (w2452 & ~w2449) | (w2452 & w43987) | (~w2449 & w43987);
assign w2454 = ~w612 & w2451;
assign w2455 = w2449 & w43988;
assign w2456 = ~w2453 & ~w2455;
assign w2457 = ~w2433 & ~w2430;
assign w2458 = (w2427 & w51028) | (w2427 & w51029) | (w51028 & w51029);
assign w2459 = w2285 & w47034;
assign w2460 = (w1866 & w2000) | (w1866 & w51030) | (w2000 & w51030);
assign w2461 = ~w2000 & w51031;
assign w2462 = ~w2460 & ~w2461;
assign w2463 = (~w493 & w2285) | (~w493 & w47035) | (w2285 & w47035);
assign w2464 = ~w2459 & w2463;
assign w2465 = w2456 & ~w2464;
assign w2466 = w2425 & w2465;
assign w2467 = ~w2445 & ~w2466;
assign w2468 = w2396 & ~w2467;
assign w2469 = ~w2381 & w2468;
assign w2470 = w2449 & w43989;
assign w2471 = (w2451 & ~w2449) | (w2451 & w43990) | (~w2449 & w43990);
assign w2472 = ~w2470 & ~w2471;
assign w2473 = w612 & ~w2472;
assign w2474 = w754 & ~w2392;
assign w2475 = ~w2473 & ~w2474;
assign w2476 = w2466 & ~w2475;
assign w2477 = (~w2127 & w2249) | (~w2127 & w43991) | (w2249 & w43991);
assign w2478 = ~w2292 & w39962;
assign w2479 = w2047 & ~w2478;
assign w2480 = ~w2477 & ~w2479;
assign w2481 = w2285 & ~w2480;
assign w2482 = w2477 & w2479;
assign w2483 = w2481 & ~w2482;
assign w2484 = (w2130 & ~w2285) | (w2130 & w47036) | (~w2285 & w47036);
assign w2485 = ~w252 & ~w2484;
assign w2486 = ~w2483 & w2485;
assign w2487 = ~w2404 & ~w2405;
assign w2488 = w351 & ~w2487;
assign w2489 = ~w2486 & ~w2488;
assign w2490 = ~w2445 & w2489;
assign w2491 = ~w2476 & w2490;
assign w2492 = ~w2469 & w2491;
assign w2493 = (~w2484 & ~w2481) | (~w2484 & w51032) | (~w2481 & w51032);
assign w2494 = (w252 & w2483) | (w252 & w43992) | (w2483 & w43992);
assign w2495 = (~w2494 & w2469) | (~w2494 & w39963) | (w2469 & w39963);
assign w2496 = ~w2300 & w47037;
assign w2497 = ~w2494 & ~w2496;
assign w2498 = (w2497 & w2469) | (w2497 & w39964) | (w2469 & w39964);
assign w2499 = (~w57 & w2300) | (~w57 & w43993) | (w2300 & w43993);
assign w2500 = ~w2111 & ~w2336;
assign w2501 = ~w3 & ~w2285;
assign w2502 = ~w2284 & w43994;
assign w2503 = ~w2500 & w2502;
assign w2504 = ~w2501 & ~w2503;
assign w2505 = ~w2088 & ~w2103;
assign w2506 = w42 & ~w2505;
assign w2507 = w2504 & w2506;
assign w2508 = w42 & w2505;
assign w2509 = ~w2504 & w2508;
assign w2510 = ~w2507 & ~w2509;
assign w2511 = ~w1965 & w2106;
assign w2512 = w2020 & ~w2511;
assign w2513 = (w2336 & w51036) | (w2336 & w51037) | (w51036 & w51037);
assign w2514 = ~w2021 & ~w2512;
assign w2515 = w2514 & w52147;
assign w2516 = ~w2513 & ~w2515;
assign w2517 = w2510 & w2516;
assign w2518 = w2068 & ~w2293;
assign w2519 = ~w2035 & ~w2063;
assign w2520 = ~w2284 & w43995;
assign w2521 = ~w2518 & w2520;
assign w2522 = ~w2284 & w43996;
assign w2523 = w2518 & w2522;
assign w2524 = ~w2521 & ~w2523;
assign w2525 = (w80 & ~w2524) | (w80 & w39965) | (~w2524 & w39965);
assign w2526 = ~w2499 & ~w2525;
assign w2527 = w2524 & w39966;
assign w2528 = (w80 & w2284) | (w80 & w43997) | (w2284 & w43997);
assign w2529 = w2285 & w2336;
assign w2530 = w2099 & ~w2111;
assign w2531 = w3 & ~w2530;
assign w2532 = ~w2529 & w43998;
assign w2533 = w3 & w2530;
assign w2534 = (w2533 & w2529) | (w2533 & w43999) | (w2529 & w43999);
assign w2535 = ~w2532 & ~w2534;
assign w2536 = ~w2527 & w2535;
assign w2537 = ~w2526 & w2536;
assign w2538 = ~w3 & w2530;
assign w2539 = ~w2529 & w44000;
assign w2540 = ~w3 & ~w2530;
assign w2541 = (w2540 & w2529) | (w2540 & w44001) | (w2529 & w44001);
assign w2542 = ~w2539 & ~w2541;
assign w2543 = ~w42 & w2505;
assign w2544 = w2504 & w2543;
assign w2545 = ~w42 & ~w2505;
assign w2546 = ~w2504 & w2545;
assign w2547 = w2542 & ~w2546;
assign w2548 = ~w2544 & w2547;
assign w2549 = ~w2537 & w2548;
assign w2550 = w2517 & ~w2549;
assign w2551 = (~w2499 & w2549) | (~w2499 & w51038) | (w2549 & w51038);
assign w2552 = ~w2498 & w2551;
assign w2553 = w2497 & w2536;
assign w2554 = w2549 & ~w2553;
assign w2555 = w2517 & ~w2554;
assign w2556 = w2491 & w2549;
assign w2557 = ~w2469 & w2556;
assign w2558 = w2555 & ~w2557;
assign w2559 = (~w57 & w2557) | (~w57 & w39967) | (w2557 & w39967);
assign w2560 = ~w2552 & w2559;
assign w2561 = ~w2301 & w2495;
assign w2562 = w2560 & ~w2561;
assign w2563 = ~w2495 & w2496;
assign w2564 = (~w2554 & w51039) | (~w2554 & w51040) | (w51039 & w51040);
assign w2565 = (~w2564 & w2498) | (~w2564 & w51041) | (w2498 & w51041);
assign w2566 = ~w2563 & ~w2565;
assign w2567 = (~w80 & w2562) | (~w80 & w51042) | (w2562 & w51042);
assign w2568 = (w80 & w2495) | (w80 & w44003) | (w2495 & w44003);
assign w2569 = ~w2565 & w2568;
assign w2570 = ~w2562 & w2569;
assign w2571 = ~w2567 & ~w2570;
assign w2572 = w2527 & ~w2535;
assign w2573 = w2527 & ~w2542;
assign w2574 = (~w2572 & w2517) | (~w2572 & w51043) | (w2517 & w51043);
assign w2575 = w2526 & w52148;
assign w2576 = w2497 & w2574;
assign w2577 = (w2576 & w2469) | (w2576 & w51044) | (w2469 & w51044);
assign w2578 = w2574 & ~w2575;
assign w2579 = (~w2578 & w2492) | (~w2578 & w44005) | (w2492 & w44005);
assign w2580 = (w2553 & w2469) | (w2553 & w39968) | (w2469 & w39968);
assign w2581 = ~w2537 & w52149;
assign w2582 = ~w2580 & w2581;
assign w2583 = (~w2530 & w2529) | (~w2530 & w51045) | (w2529 & w51045);
assign w2584 = ~w2529 & w51046;
assign w2585 = ~w2583 & ~w2584;
assign w2586 = w2510 & w51047;
assign w2587 = (w2542 & w2557) | (w2542 & w39969) | (w2557 & w39969);
assign w2588 = ~w2582 & w2587;
assign w2589 = ~w2579 & ~w2588;
assign w2590 = ~w2588 & w44006;
assign w2591 = ~w2537 & w2542;
assign w2592 = w2504 & ~w2505;
assign w2593 = ~w2504 & w2505;
assign w2594 = ~w2592 & ~w2593;
assign w2595 = ~w1976 & w52146;
assign w2596 = ~w1969 & ~w2595;
assign w2597 = w2106 & ~w2596;
assign w2598 = ~w2597 & w52147;
assign w2599 = (w2336 & w51048) | (w2336 & w51049) | (w51048 & w51049);
assign w2600 = ~w2598 & ~w2599;
assign w2601 = w2594 & w2600;
assign w2602 = w2594 & w51050;
assign w2603 = w2510 & ~w2602;
assign w2604 = ~w2020 & w52147;
assign w2605 = (w2336 & w51051) | (w2336 & w51052) | (w51051 & w51052);
assign w2606 = w2594 & w51053;
assign w2607 = ~w2580 & w44007;
assign w2608 = w2510 & ~w2606;
assign w2609 = (w2608 & w2580) | (w2608 & w44008) | (w2580 & w44008);
assign w2610 = ~w2607 & ~w2609;
assign w2611 = w2590 & w2610;
assign w2612 = ~w2557 & w39970;
assign w2613 = ~w2552 & ~w2612;
assign w2614 = ~w2525 & ~w2527;
assign w2615 = w3 & ~w2614;
assign w2616 = ~w2613 & w2615;
assign w2617 = w3 & w2614;
assign w2618 = w2613 & w2617;
assign w2619 = ~w2616 & ~w2618;
assign w2620 = w42 & w2542;
assign w2621 = (w2620 & w2557) | (w2620 & w39971) | (w2557 & w39971);
assign w2622 = ~w2582 & w2621;
assign w2623 = ~w2577 & w39972;
assign w2624 = ~w2622 & ~w2623;
assign w2625 = w2610 & w2624;
assign w2626 = w2619 & w2625;
assign w2627 = ~w2611 & ~w2626;
assign w2628 = w2613 & ~w2614;
assign w2629 = ~w2613 & w2614;
assign w2630 = ~w2628 & ~w2629;
assign w2631 = ~w3 & ~w2630;
assign w2632 = ~w2611 & ~w2631;
assign w2633 = ~w2486 & ~w2494;
assign w2634 = ~w2445 & ~w2488;
assign w2635 = ~w2476 & w2634;
assign w2636 = ~w2469 & w39973;
assign w2637 = ~w2550 & ~w2636;
assign w2638 = (w2633 & w2469) | (w2633 & w44009) | (w2469 & w44009);
assign w2639 = ~w2554 & w51054;
assign w2640 = (~w2639 & ~w2637) | (~w2639 & w44010) | (~w2637 & w44010);
assign w2641 = ~w57 & ~w2640;
assign w2642 = ~w2570 & ~w2641;
assign w2643 = ~w2567 & ~w2642;
assign w2644 = w2632 & ~w2643;
assign w2645 = ~w2627 & ~w2644;
assign w2646 = w57 & w2640;
assign w2647 = ~w2569 & w2646;
assign w2648 = ~w2567 & ~w2647;
assign w2649 = ~w2627 & w2648;
assign w2650 = w2438 & ~w2465;
assign w2651 = w2396 & ~w2650;
assign w2652 = w2465 & ~w2475;
assign w2653 = ~w2381 & w2651;
assign w2654 = (~w400 & w2653) | (~w400 & w39974) | (w2653 & w39974);
assign w2655 = ~w2653 & w39975;
assign w2656 = w2418 & ~w2419;
assign w2657 = ~w2418 & w2419;
assign w2658 = ~w2656 & ~w2657;
assign w2659 = (~w2658 & w2653) | (~w2658 & w51055) | (w2653 & w51055);
assign w2660 = ~w2558 & w51056;
assign w2661 = ~w2557 & w44011;
assign w2662 = ~w2407 & ~w2488;
assign w2663 = ~w2660 & w39976;
assign w2664 = (w2662 & w2660) | (w2662 & w39977) | (w2660 & w39977);
assign w2665 = ~w2663 & ~w2664;
assign w2666 = w252 & w2665;
assign w2667 = ~w2558 & w39978;
assign w2668 = w2658 & ~w2667;
assign w2669 = ~w2658 & w2667;
assign w2670 = ~w2668 & ~w2669;
assign w2671 = w351 & w2670;
assign w2672 = ~w2488 & w51057;
assign w2673 = (w2672 & w2660) | (w2672 & w39979) | (w2660 & w39979);
assign w2674 = (~w252 & w2488) | (~w252 & w51058) | (w2488 & w51058);
assign w2675 = ~w2660 & w39980;
assign w2676 = ~w2673 & ~w2675;
assign w2677 = ~w2671 & w2676;
assign w2678 = ~w2666 & ~w2677;
assign w2679 = w2649 & w2678;
assign w2680 = ~w2645 & ~w2679;
assign w2681 = ~w2381 & w2396;
assign w2682 = ~w2360 & ~w2382;
assign w2683 = ~w2363 & w2682;
assign w2684 = ~w2359 & w2683;
assign w2685 = ~w2373 & ~w2383;
assign w2686 = ~w2379 & w2685;
assign w2687 = ~w2684 & w2686;
assign w2688 = w754 & w2392;
assign w2689 = (~w2688 & w39981) | (~w2688 & w2687) | (w39981 & w2687);
assign w2690 = w2510 & w51059;
assign w2691 = ~w2554 & w2690;
assign w2692 = ~w2557 & w2691;
assign w2693 = ~w754 & ~w2392;
assign w2694 = (w39982 & w2684) | (w39982 & w44012) | (w2684 & w44012);
assign w2695 = (w2693 & w39983) | (w2693 & w2687) | (w39983 & w2687);
assign w2696 = ~w2694 & ~w2695;
assign w2697 = ~w2692 & w2696;
assign w2698 = ~w2681 & ~w2689;
assign w2699 = ~w2558 & w2698;
assign w2700 = w2697 & ~w2699;
assign w2701 = w612 & ~w2700;
assign w2702 = (~w2379 & ~w2683) | (~w2379 & w51060) | (~w2683 & w51060);
assign w2703 = ~w2685 & ~w2702;
assign w2704 = ~w2557 & w39984;
assign w2705 = ~w2687 & ~w2703;
assign w2706 = ~w2558 & w2705;
assign w2707 = ~w2706 & w39985;
assign w2708 = ~w2701 & ~w2707;
assign w2709 = w2456 & ~w2473;
assign w2710 = w2396 & w2709;
assign w2711 = ~w2381 & w2710;
assign w2712 = (~w2474 & w2473) | (~w2474 & w51061) | (w2473 & w51061);
assign w2713 = (w2712 & w2381) | (w2712 & w39986) | (w2381 & w39986);
assign w2714 = ~w2473 & w51062;
assign w2715 = ~w2711 & ~w2714;
assign w2716 = ~w2713 & w2715;
assign w2717 = ~w2557 & w39987;
assign w2718 = ~w2558 & w2716;
assign w2719 = ~w2717 & ~w2718;
assign w2720 = ~w2718 & w39988;
assign w2721 = ~w612 & w2700;
assign w2722 = ~w2720 & ~w2721;
assign w2723 = (w493 & w2718) | (w493 & w51063) | (w2718 & w51063);
assign w2724 = (~w2433 & w2432) | (~w2433 & w51064) | (w2432 & w51064);
assign w2725 = ~w2432 & w51065;
assign w2726 = ~w2724 & ~w2725;
assign w2727 = w2438 & ~w2464;
assign w2728 = w2394 & w39989;
assign w2729 = (w2456 & w2473) | (w2456 & w51062) | (w2473 & w51062);
assign w2730 = ~w2727 & ~w50181;
assign w2731 = w2727 & w50181;
assign w2732 = ~w2557 & w51066;
assign w2733 = ~w2558 & w39991;
assign w2734 = ~w2732 & ~w2733;
assign w2735 = (~w400 & w2733) | (~w400 & w51067) | (w2733 & w51067);
assign w2736 = ~w2723 & ~w2735;
assign w2737 = ~w2708 & w2722;
assign w2738 = w2736 & ~w2737;
assign w2739 = ~w2379 & ~w2382;
assign w2740 = w2365 & ~w2739;
assign w2741 = ~w2365 & w2739;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = w945 & w2378;
assign w2744 = ~w2557 & w39992;
assign w2745 = w945 & w2742;
assign w2746 = ~w2558 & w2745;
assign w2747 = ~w2744 & ~w2746;
assign w2748 = ~w2334 & ~w2360;
assign w2749 = ~w2329 & ~w2357;
assign w2750 = (w2748 & w2749) | (w2748 & w44013) | (w2749 & w44013);
assign w2751 = ~w2749 & w44014;
assign w2752 = ~w2750 & ~w2751;
assign w2753 = w1120 & w2333;
assign w2754 = ~w2557 & w39993;
assign w2755 = w1120 & w2752;
assign w2756 = (w2755 & w2557) | (w2755 & w39994) | (w2557 & w39994);
assign w2757 = ~w2754 & ~w2756;
assign w2758 = w2747 & w2757;
assign w2759 = ~w945 & ~w2378;
assign w2760 = ~w2557 & w39995;
assign w2761 = ~w945 & ~w2742;
assign w2762 = ~w2558 & w2761;
assign w2763 = ~w2760 & ~w2762;
assign w2764 = ~w2329 & ~w2362;
assign w2765 = ~w2357 & w2764;
assign w2766 = (w2765 & w2557) | (w2765 & w39996) | (w2557 & w39996);
assign w2767 = w2357 & ~w2764;
assign w2768 = (w2557 & w51068) | (w2557 & w51069) | (w51068 & w51069);
assign w2769 = w1320 & w2357;
assign w2770 = (~w2557 & w51070) | (~w2557 & w51071) | (w51070 & w51071);
assign w2771 = ~w2768 & ~w2770;
assign w2772 = ~w1120 & ~w2333;
assign w2773 = ~w2557 & w39998;
assign w2774 = ~w1120 & ~w2752;
assign w2775 = (w2774 & w2557) | (w2774 & w39999) | (w2557 & w39999);
assign w2776 = ~w2773 & ~w2775;
assign w2777 = ~w2758 & w2763;
assign w2778 = w2763 & w51072;
assign w2779 = ~w2777 & ~w2778;
assign w2780 = (~w754 & w2706) | (~w754 & w40000) | (w2706 & w40000);
assign w2781 = ~w2701 & w2780;
assign w2782 = w2722 & ~w2781;
assign w2783 = w2779 & w2782;
assign w2784 = w2738 & ~w2783;
assign w2785 = ~w2733 & w51073;
assign w2786 = (~w2785 & w2670) | (~w2785 & w51074) | (w2670 & w51074);
assign w2787 = w1738 & w2322;
assign w2788 = ~w1738 & ~w2322;
assign w2789 = ~w2787 & ~w2788;
assign w2790 = ~w2285 & w2304;
assign w2791 = w2285 & w2306;
assign w2792 = ~w2790 & ~w2791;
assign w2793 = (w2557 & w44015) | (w2557 & w44016) | (w44015 & w44016);
assign w2794 = (~w2557 & w44017) | (~w2557 & w44018) | (w44017 & w44018);
assign w2795 = ~w2793 & ~w2794;
assign w2796 = w1541 & ~w2795;
assign w2797 = ~w2006 & ~w2285;
assign w2798 = w2006 & w2285;
assign w2799 = ~w2797 & ~w2798;
assign w2800 = ~a[94] & w2285;
assign w2801 = ~w2557 & w40001;
assign w2802 = ~w2313 & w2799;
assign w2803 = (w2802 & w2557) | (w2802 & w40002) | (w2557 & w40002);
assign w2804 = ~w2801 & ~w2803;
assign w2805 = w2285 & w51075;
assign w2806 = ~w2285 & w51076;
assign w2807 = ~w2557 & w40003;
assign w2808 = w2313 & ~w2799;
assign w2809 = (~a[95] & ~w2804) | (~a[95] & w44022) | (~w2804 & w44022);
assign w2810 = w2804 & w44023;
assign w2811 = ~w2809 & ~w2810;
assign w2812 = a[94] & ~w2285;
assign w2813 = ~w2800 & ~w2812;
assign w2814 = w2510 & w51077;
assign w2815 = ~w2554 & w2814;
assign w2816 = ~w2557 & w2815;
assign w2817 = a[94] & ~w2312;
assign w2818 = ~w2313 & ~w2817;
assign w2819 = ~w2557 & w40004;
assign w2820 = ~w2000 & w51078;
assign w2821 = (w2820 & w2557) | (w2820 & w40005) | (w2557 & w40005);
assign w2822 = ~w2819 & ~w2821;
assign w2823 = (w2818 & w2557) | (w2818 & w40006) | (w2557 & w40006);
assign w2824 = ~a[90] & ~a[91];
assign w2825 = ~a[92] & w2824;
assign w2826 = ~w2285 & ~w2825;
assign w2827 = (~w2312 & w2285) | (~w2312 & w51080) | (w2285 & w51080);
assign w2828 = w2285 & w2825;
assign w2829 = (~a[93] & w2285) | (~a[93] & w51081) | (w2285 & w51081);
assign w2830 = ~w2827 & ~w2828;
assign w2831 = (w2830 & w2557) | (w2830 & w40007) | (w2557 & w40007);
assign w2832 = ~w2828 & ~w2829;
assign w2833 = ~w2557 & w40008;
assign w2834 = ~w2831 & ~w2833;
assign w2835 = (~w2006 & w2557) | (~w2006 & w40009) | (w2557 & w40009);
assign w2836 = ~w2823 & w2835;
assign w2837 = w2834 & ~w2836;
assign w2838 = (w1738 & w2837) | (w1738 & w44024) | (w2837 & w44024);
assign w2839 = ~w2811 & ~w2838;
assign w2840 = ~w1738 & w2822;
assign w2841 = ~w2837 & w2840;
assign w2842 = ~w1541 & w2795;
assign w2843 = ~w2841 & ~w2842;
assign w2844 = ~w2839 & w2843;
assign w2845 = ~w2796 & ~w2844;
assign w2846 = (~w2557 & w44025) | (~w2557 & w44026) | (w44025 & w44026);
assign w2847 = (~w2557 & w44027) | (~w2557 & w44028) | (w44027 & w44028);
assign w2848 = ~w2846 & w2847;
assign w2849 = w2776 & w2848;
assign w2850 = w2758 & ~w2849;
assign w2851 = w2782 & w2850;
assign w2852 = w2782 & w51082;
assign w2853 = ~w2784 & w2786;
assign w2854 = ~w2845 & w2852;
assign w2855 = ~w2853 & ~w2854;
assign w2856 = ~w2631 & ~w2648;
assign w2857 = w2626 & ~w2666;
assign w2858 = ~w2856 & w2857;
assign w2859 = ~w2645 & ~w2858;
assign w2860 = (w2763 & ~w2758) | (w2763 & w51083) | (~w2758 & w51083);
assign w2861 = ~w2737 & w51084;
assign w2862 = w2845 & w2861;
assign w2863 = ~w2859 & ~w2862;
assign w2864 = ~w2855 & w2863;
assign w2865 = w2680 & ~w2864;
assign w2866 = ~w2666 & w2786;
assign w2867 = (~w2678 & w2784) | (~w2678 & w40010) | (w2784 & w40010);
assign w2868 = w2851 & w2866;
assign w2869 = ~w2845 & w2868;
assign w2870 = w2867 & ~w2869;
assign w2871 = (~w2646 & ~w40011) | (~w2646 & w44029) | (~w40011 & w44029);
assign w2872 = w2865 & w2871;
assign w2873 = ~w2872 & w47039;
assign w2874 = (~w2571 & w2872) | (~w2571 & w47040) | (w2872 & w47040);
assign w2875 = ~w2873 & ~w2874;
assign w2876 = ~w3 & ~w2875;
assign w2877 = (~w2862 & w2853) | (~w2862 & w51085) | (w2853 & w51085);
assign w2878 = w2648 & ~w2666;
assign w2879 = ~w2677 & w2878;
assign w2880 = ~w2643 & ~w2879;
assign w2881 = (w2880 & w2855) | (w2880 & w48591) | (w2855 & w48591);
assign w2882 = ~w3 & ~w2881;
assign w2883 = ~w2879 & w51086;
assign w2884 = (w2883 & w2855) | (w2883 & w51087) | (w2855 & w51087);
assign w2885 = w2865 & ~w2884;
assign w2886 = ~w42 & ~w2630;
assign w2887 = (w2886 & ~w2885) | (w2886 & w48592) | (~w2885 & w48592);
assign w2888 = ~w42 & w2630;
assign w2889 = w2885 & w48593;
assign w2890 = ~w2887 & ~w2889;
assign w2891 = ~w2876 & w2890;
assign w2892 = ~w2845 & w2851;
assign w2893 = w2784 & ~w2892;
assign w2894 = w2649 & w2866;
assign w2895 = ~w2893 & w2894;
assign w2896 = w2680 & ~w2895;
assign w2897 = w2632 & ~w2648;
assign w2898 = ~w2680 & ~w2897;
assign w2899 = ~w2895 & ~w2898;
assign w2900 = ~w2631 & ~w2643;
assign w2901 = w2589 & w2619;
assign w2902 = ~w2643 & w51088;
assign w2903 = (w2902 & w2870) | (w2902 & w51089) | (w2870 & w51089);
assign w2904 = w2630 & ~w2899;
assign w2905 = w2903 & ~w2904;
assign w2906 = w2589 & ~w2610;
assign w2907 = w2631 & ~w2906;
assign w2908 = (w2589 & w2897) | (w2589 & w44031) | (w2897 & w44031);
assign w2909 = (w2897 & w51090) | (w2897 & w51091) | (w51090 & w51091);
assign w2910 = (w2870 & w51465) | (w2870 & w51466) | (w51465 & w51466);
assign w2911 = (~w2630 & w2895) | (~w2630 & w51094) | (w2895 & w51094);
assign w2912 = ~w2884 & w2911;
assign w2913 = ~w2905 & w51095;
assign w2914 = w2619 & ~w2856;
assign w2915 = (w2594 & w2580) | (w2594 & w51491) | (w2580 & w51491);
assign w2916 = ~w2580 & w51097;
assign w2917 = ~w2915 & ~w2916;
assign w2918 = w2589 & w2917;
assign w2919 = (w2870 & w51098) | (w2870 & w51099) | (w51098 & w51099);
assign w2920 = (w2870 & w51492) | (w2870 & w51493) | (w51492 & w51493);
assign w2921 = ~w2919 & w2920;
assign w2922 = ~w2913 & ~w2921;
assign w2923 = (~w2671 & w2855) | (~w2671 & w44032) | (w2855 & w44032);
assign w2924 = ~w2666 & w2676;
assign w2925 = (w2924 & w2644) | (w2924 & w51102) | (w2644 & w51102);
assign w2926 = (~w2665 & w2645) | (~w2665 & w51103) | (w2645 & w51103);
assign w2927 = ~w2925 & ~w2926;
assign w2928 = w252 & ~w2665;
assign w2929 = ~w2895 & w51104;
assign w2930 = (w252 & w2644) | (w252 & w51105) | (w2644 & w51105);
assign w2931 = w2665 & ~w2930;
assign w2932 = w2923 & ~w2927;
assign w2933 = (~w2855 & w51106) | (~w2855 & w51107) | (w51106 & w51107);
assign w2934 = ~w2929 & w2933;
assign w2935 = ~w2932 & ~w2934;
assign w2936 = ~w57 & ~w2935;
assign w2937 = ~w2869 & w40012;
assign w2938 = (w57 & w2869) | (w57 & w40013) | (w2869 & w40013);
assign w2939 = ~w2937 & ~w2938;
assign w2940 = w2865 & ~w2939;
assign w2941 = w2640 & ~w2940;
assign w2942 = ~w2640 & w2940;
assign w2943 = ~w2941 & ~w2942;
assign w2944 = w80 & w2943;
assign w2945 = (~w2936 & ~w2943) | (~w2936 & w51108) | (~w2943 & w51108);
assign w2946 = w57 & w2935;
assign w2947 = (w351 & w2893) | (w351 & w47042) | (w2893 & w47042);
assign w2948 = ~w2893 & w47043;
assign w2949 = ~w2947 & ~w2948;
assign w2950 = ~w2895 & w47044;
assign w2951 = ~w2949 & w2950;
assign w2952 = (w2670 & ~w2865) | (w2670 & w47045) | (~w2865 & w47045);
assign w2953 = ~w2951 & ~w2952;
assign w2954 = ~w2952 & w51109;
assign w2955 = ~w2946 & ~w2954;
assign w2956 = w2945 & ~w2955;
assign w2957 = ~w80 & ~w2943;
assign w2958 = w3 & ~w2571;
assign w2959 = ~w2872 & w47046;
assign w2960 = w3 & w2571;
assign w2961 = (w2960 & w2872) | (w2960 & w47047) | (w2872 & w47047);
assign w2962 = ~w2959 & ~w2961;
assign w2963 = ~w2957 & w2962;
assign w2964 = (w2922 & w2876) | (w2922 & w51110) | (w2876 & w51110);
assign w2965 = ~w2957 & w51111;
assign w2966 = ~w2956 & w2965;
assign w2967 = ~w2964 & ~w2966;
assign w2968 = ~w2557 & w51112;
assign w2969 = (w2742 & w2557) | (w2742 & w51113) | (w2557 & w51113);
assign w2970 = ~w2968 & ~w2969;
assign w2971 = w2796 & ~w2848;
assign w2972 = ~w2841 & w44033;
assign w2973 = ~w2839 & w2972;
assign w2974 = ~w2971 & ~w2973;
assign w2975 = ~w2973 & w51114;
assign w2976 = w2747 & w2763;
assign w2977 = (w2976 & w2975) | (w2976 & w51115) | (w2975 & w51115);
assign w2978 = ~w2975 & w51116;
assign w2979 = (~w2970 & w2895) | (~w2970 & w51494) | (w2895 & w51494);
assign w2980 = ~w2895 & w51117;
assign w2981 = ~w2979 & ~w2980;
assign w2982 = ~w2979 & w51118;
assign w2983 = ~w2557 & w51119;
assign w2984 = (w2752 & w2557) | (w2752 & w51120) | (w2557 & w51120);
assign w2985 = ~w2983 & ~w2984;
assign w2986 = (~w2776 & w2973) | (~w2776 & w51121) | (w2973 & w51121);
assign w2987 = ~w2899 & w2985;
assign w2988 = (~w2986 & w2899) | (~w2986 & w51122) | (w2899 & w51122);
assign w2989 = (w2645 & w2869) | (w2645 & w40014) | (w2869 & w40014);
assign w2990 = ~w2895 & ~w2989;
assign w2991 = (~w2757 & w2973) | (~w2757 & w51123) | (w2973 & w51123);
assign w2992 = (w2991 & w2680) | (w2991 & w51495) | (w2680 & w51495);
assign w2993 = ~w2989 & w51496;
assign w2994 = w2757 & w2975;
assign w2995 = w2899 & w2994;
assign w2996 = ~w2993 & ~w2995;
assign w2997 = ~w2993 & w51124;
assign w2998 = (~w945 & ~w2996) | (~w945 & w44034) | (~w2996 & w44034);
assign w2999 = (w2996 & w51125) | (w2996 & w51126) | (w51125 & w51126);
assign w3000 = (~w754 & w2979) | (~w754 & w51127) | (w2979 & w51127);
assign w3001 = w2843 & w2850;
assign w3002 = ~w2839 & w3001;
assign w3003 = w2758 & w51128;
assign w3004 = (~w3003 & ~w3001) | (~w3003 & w51129) | (~w3001 & w51129);
assign w3005 = (~w754 & w2895) | (~w754 & w47050) | (w2895 & w47050);
assign w3006 = ~w2779 & w3004;
assign w3007 = ~w2895 & w47051;
assign w3008 = ~w3005 & ~w3007;
assign w3009 = ~w2707 & ~w2780;
assign w3010 = ~w612 & ~w3009;
assign w3011 = ~w3008 & w3010;
assign w3012 = ~w612 & w3009;
assign w3013 = w3008 & w3012;
assign w3014 = ~w3011 & ~w3013;
assign w3015 = ~w3000 & w3014;
assign w3016 = ~w2999 & w3015;
assign w3017 = ~w2816 & ~w2823;
assign w3018 = w2006 & ~w2834;
assign w3019 = ~w2006 & w2834;
assign w3020 = ~w3018 & ~w3019;
assign w3021 = (~w3020 & w2680) | (~w3020 & w44035) | (w2680 & w44035);
assign w3022 = ~w2895 & w3021;
assign w3023 = w3017 & ~w3020;
assign w3024 = w2680 & w3023;
assign w3025 = ~w2864 & w3024;
assign w3026 = ~w3017 & ~w3022;
assign w3027 = ~w3025 & ~w3026;
assign w3028 = ~w1738 & w3027;
assign w3029 = ~w2838 & ~w2841;
assign w3030 = (w3029 & w2680) | (w3029 & w51130) | (w2680 & w51130);
assign w3031 = ~w2989 & w51131;
assign w3032 = w1541 & w2811;
assign w3033 = (w3032 & ~w2990) | (w3032 & w44036) | (~w2990 & w44036);
assign w3034 = w1541 & ~w2811;
assign w3035 = w2990 & w44037;
assign w3036 = ~w3033 & ~w3035;
assign w3037 = (w1541 & w2839) | (w1541 & w51132) | (w2839 & w51132);
assign w3038 = ~w2839 & w51133;
assign w3039 = ~w3037 & ~w3038;
assign w3040 = (w2795 & ~w2680) | (w2795 & w44038) | (~w2680 & w44038);
assign w3041 = w2649 & w51134;
assign w3042 = ~w2893 & w3041;
assign w3043 = ~w3040 & ~w3042;
assign w3044 = ~w2795 & ~w3039;
assign w3045 = (w3044 & w2680) | (w3044 & w51135) | (w2680 & w51135);
assign w3046 = ~w1320 & ~w3043;
assign w3047 = ~w2898 & w44039;
assign w3048 = w2990 & w3047;
assign w3049 = ~w3046 & ~w3048;
assign w3050 = ~w1541 & w2811;
assign w3051 = w3031 & w3050;
assign w3052 = ~w1541 & ~w2811;
assign w3053 = (w3052 & ~w2990) | (w3052 & w44040) | (~w2990 & w44040);
assign w3054 = w3049 & w51136;
assign w3055 = w3028 & w3036;
assign w3056 = w3054 & ~w3055;
assign w3057 = ~w2844 & w51137;
assign w3058 = ~w2844 & w51138;
assign w3059 = (~w3058 & ~w2990) | (~w3058 & w44041) | (~w2990 & w44041);
assign w3060 = ~w2766 & ~w2846;
assign w3061 = (w3060 & w2864) | (w3060 & w44042) | (w2864 & w44042);
assign w3062 = (~w1320 & w2973) | (~w1320 & w47052) | (w2973 & w47052);
assign w3063 = (w3062 & w2680) | (w3062 & w44043) | (w2680 & w44043);
assign w3064 = ~w2895 & w3063;
assign w3065 = ~w1120 & ~w3064;
assign w3066 = ~w3061 & w3065;
assign w3067 = w3059 & w3066;
assign w3068 = w1320 & ~w2795;
assign w3069 = w2680 & w44044;
assign w3070 = ~w2895 & w3069;
assign w3071 = ~w3068 & ~w3070;
assign w3072 = ~w2989 & w51139;
assign w3073 = ~w3071 & ~w3072;
assign w3074 = ~w3067 & ~w3073;
assign w3075 = (w3074 & ~w3054) | (w3074 & w44045) | (~w3054 & w44045);
assign w3076 = ~w3061 & ~w3064;
assign w3077 = w3059 & w3076;
assign w3078 = w1120 & ~w3077;
assign w3079 = w2996 & w44046;
assign w3080 = ~w3078 & ~w3079;
assign w3081 = w3015 & w3080;
assign w3082 = ~w3075 & w3081;
assign w3083 = ~w3016 & ~w3082;
assign w3084 = (~a[92] & w2557) | (~a[92] & w51140) | (w2557 & w51140);
assign w3085 = (w2828 & w2557) | (w2828 & w51141) | (w2557 & w51141);
assign w3086 = a[93] & ~w3085;
assign w3087 = (w3084 & ~w2632) | (w3084 & w51142) | (~w2632 & w51142);
assign w3088 = (w3086 & w2859) | (w3086 & w47053) | (w2859 & w47053);
assign w3089 = (a[93] & ~w2285) | (a[93] & w51143) | (~w2285 & w51143);
assign w3090 = (w3089 & w2588) | (w3089 & w51497) | (w2588 & w51497);
assign w3091 = ~w2671 & w51144;
assign w3092 = w2900 & w3091;
assign w3093 = (w3092 & w2855) | (w3092 & w44047) | (w2855 & w44047);
assign w3094 = ~w3088 & ~w3093;
assign w3095 = (w2285 & w2557) | (w2285 & w51145) | (w2557 & w51145);
assign w3096 = ~w2807 & ~w3095;
assign w3097 = ~w2825 & w3096;
assign w3098 = ~w2557 & w51146;
assign w3099 = (~w3098 & ~w3096) | (~w3098 & w51147) | (~w3096 & w51147);
assign w3100 = w2826 & w3084;
assign w3101 = (~w3100 & w2864) | (~w3100 & w44048) | (w2864 & w44048);
assign w3102 = ~w2285 & w2824;
assign w3103 = (w3102 & w2644) | (w3102 & w44049) | (w2644 & w44049);
assign w3104 = ~w2645 & w51148;
assign w3105 = w2558 & ~w3104;
assign w3106 = (w2677 & w3103) | (w2677 & w51149) | (w3103 & w51149);
assign w3107 = ~w2877 & w3106;
assign w3108 = w3105 & ~w3107;
assign w3109 = w2285 & ~w2824;
assign w3110 = (~w3109 & ~w3096) | (~w3109 & w51150) | (~w3096 & w51150);
assign w3111 = (~w3110 & w2644) | (~w3110 & w44050) | (w2644 & w44050);
assign w3112 = (w2677 & w3111) | (w2677 & w51151) | (w3111 & w51151);
assign w3113 = (w2312 & ~w3111) | (w2312 & w51152) | (~w3111 & w51152);
assign w3114 = (w3113 & w2877) | (w3113 & w44051) | (w2877 & w44051);
assign w3115 = ~w3094 & w3101;
assign w3116 = ~w3108 & w3114;
assign w3117 = w2834 & w3097;
assign w3118 = ~w2895 & w47054;
assign w3119 = ~a[88] & ~a[89];
assign w3120 = (w3119 & w2557) | (w3119 & w51153) | (w2557 & w51153);
assign w3121 = w2824 & ~w3120;
assign w3122 = ~a[90] & w3119;
assign w3123 = a[90] & ~a[91];
assign w3124 = ~w3122 & ~w3123;
assign w3125 = ~w2557 & w51154;
assign w3126 = (~w3125 & ~w2680) | (~w3125 & w44052) | (~w2680 & w44052);
assign w3127 = w2649 & w51155;
assign w3128 = ~w2893 & w3127;
assign w3129 = ~w3126 & ~w3128;
assign w3130 = (a[91] & ~w3119) | (a[91] & w51156) | (~w3119 & w51156);
assign w3131 = ~w2557 & w51157;
assign w3132 = ~w3130 & ~w3131;
assign w3133 = ~w2680 & w44053;
assign w3134 = w2649 & w51158;
assign w3135 = ~w2893 & w3134;
assign w3136 = ~w3133 & ~w3135;
assign w3137 = ~w3129 & w3136;
assign w3138 = ~w2285 & ~w3137;
assign w3139 = w2285 & w3137;
assign w3140 = w2649 & w51159;
assign w3141 = (a[92] & w2680) | (a[92] & w44054) | (w2680 & w44054);
assign w3142 = ~w2893 & w3140;
assign w3143 = w3141 & ~w3142;
assign w3144 = (~w2824 & w2680) | (~w2824 & w44055) | (w2680 & w44055);
assign w3145 = ~w2895 & w3144;
assign w3146 = w3143 & ~w3145;
assign w3147 = ~a[92] & ~w2824;
assign w3148 = (w3147 & w2680) | (w3147 & w44056) | (w2680 & w44056);
assign w3149 = ~w2895 & w3148;
assign w3150 = ~w2680 & w44057;
assign w3151 = w2649 & w51160;
assign w3152 = ~w2893 & w3151;
assign w3153 = ~w3150 & ~w3152;
assign w3154 = ~w3149 & w3153;
assign w3155 = ~w3146 & w3154;
assign w3156 = ~w3139 & w3155;
assign w3157 = (~w3138 & ~w3155) | (~w3138 & w44058) | (~w3155 & w44058);
assign w3158 = w2006 & ~w3118;
assign w3159 = ~w3116 & w44059;
assign w3160 = ~w3157 & ~w3159;
assign w3161 = ~w3116 & w44060;
assign w3162 = (~w2006 & ~w44060) | (~w2006 & w51161) | (~w44060 & w51161);
assign w3163 = ~w3160 & ~w3162;
assign w3164 = ~w3036 & w3049;
assign w3165 = ~w2864 & w44061;
assign w3166 = w1738 & ~w3017;
assign w3167 = ~w3022 & w3166;
assign w3168 = ~w3165 & ~w3167;
assign w3169 = ~w3073 & w3168;
assign w3170 = ~w3067 & w3169;
assign w3171 = ~w3164 & w3170;
assign w3172 = w2999 & w3171;
assign w3173 = ~w3163 & w3172;
assign w3174 = ~w2779 & w51162;
assign w3175 = ~w2721 & ~w2781;
assign w3176 = (~w40015 & w51163) | (~w40015 & w51164) | (w51163 & w51164);
assign w3177 = ~w2720 & w3176;
assign w3178 = ~w2864 & w51165;
assign w3179 = w3175 & w52150;
assign w3180 = ~w2898 & w3179;
assign w3181 = ~w2895 & w3180;
assign w3182 = ~w2680 & ~w2719;
assign w3183 = w3175 & w52151;
assign w3184 = ~w3182 & ~w3183;
assign w3185 = w2649 & w51168;
assign w3186 = ~w2893 & w3185;
assign w3187 = w3184 & ~w3186;
assign w3188 = ~w3181 & w3187;
assign w3189 = ~w3178 & w3188;
assign w3190 = (~w400 & ~w3188) | (~w400 & w51169) | (~w3188 & w51169);
assign w3191 = w3188 & w51170;
assign w3192 = ~w2701 & ~w2721;
assign w3193 = (~w2707 & w2777) | (~w2707 & w51171) | (w2777 & w51171);
assign w3194 = w2780 & ~w3192;
assign w3195 = ~w2779 & w40016;
assign w3196 = (~w3194 & ~w3004) | (~w3194 & w40017) | (~w3004 & w40017);
assign w3197 = w2680 & w3196;
assign w3198 = (w2700 & w2895) | (w2700 & w40018) | (w2895 & w40018);
assign w3199 = w2680 & ~w3196;
assign w3200 = ~w2864 & w3199;
assign w3201 = ~w2780 & w3192;
assign w3202 = (w3201 & ~w3004) | (w3201 & w40019) | (~w3004 & w40019);
assign w3203 = (w3202 & w2680) | (w3202 & w51172) | (w2680 & w51172);
assign w3204 = ~w2895 & w3203;
assign w3205 = ~w3200 & ~w3204;
assign w3206 = ~w3198 & w3205;
assign w3207 = (~w493 & ~w3205) | (~w493 & w40020) | (~w3205 & w40020);
assign w3208 = ~w3191 & ~w3207;
assign w3209 = ~w3190 & ~w3208;
assign w3210 = (w40015 & w51173) | (w40015 & w51174) | (w51173 & w51174);
assign w3211 = ~w2735 & ~w2785;
assign w3212 = ~w3210 & w3211;
assign w3213 = (~w400 & w2895) | (~w400 & w40022) | (w2895 & w40022);
assign w3214 = w3212 & ~w3213;
assign w3215 = (w40015 & w51175) | (w40015 & w51176) | (w51175 & w51176);
assign w3216 = ~w2895 & w51498;
assign w3217 = (~w2734 & w2895) | (~w2734 & w40023) | (w2895 & w40023);
assign w3218 = ~w3216 & ~w3217;
assign w3219 = ~w3214 & w3218;
assign w3220 = w3218 & w47055;
assign w3221 = (~w3220 & w3208) | (~w3220 & w44062) | (w3208 & w44062);
assign w3222 = (w3221 & ~w3172) | (w3221 & w44063) | (~w3172 & w44063);
assign w3223 = ~w3083 & w3222;
assign w3224 = (w351 & ~w3218) | (w351 & w40024) | (~w3218 & w40024);
assign w3225 = ~w252 & w2951;
assign w3226 = ~w252 & w2670;
assign w3227 = (w3226 & w2949) | (w3226 & w40025) | (w2949 & w40025);
assign w3228 = ~w3225 & ~w3227;
assign w3229 = ~w3224 & w3228;
assign w3230 = w612 & ~w3009;
assign w3231 = w3008 & w3230;
assign w3232 = w612 & w3009;
assign w3233 = ~w3008 & w3232;
assign w3234 = ~w3231 & ~w3233;
assign w3235 = w3205 & w40026;
assign w3236 = ~w3190 & w47056;
assign w3237 = (w3229 & ~w3221) | (w3229 & w40027) | (~w3221 & w40027);
assign w3238 = ~w2945 & w2963;
assign w3239 = (w2922 & w3238) | (w2922 & w2964) | (w3238 & w2964);
assign w3240 = w3237 & ~w3239;
assign w3241 = ~w3223 & w3240;
assign w3242 = (~w2967 & ~w3240) | (~w2967 & w44064) | (~w3240 & w44064);
assign w3243 = ~a[86] & ~a[87];
assign w3244 = ~a[88] & w3243;
assign w3245 = (~w3244 & w2895) | (~w3244 & w51177) | (w2895 & w51177);
assign w3246 = (~w3119 & ~w3245) | (~w3119 & w51178) | (~w3245 & w51178);
assign w3247 = ~w2895 & w51499;
assign w3248 = ~a[89] & ~w3245;
assign w3249 = (w3248 & w2966) | (w3248 & w40028) | (w2966 & w40028);
assign w3250 = (~w3247 & w3241) | (~w3247 & w40029) | (w3241 & w40029);
assign w3251 = (~w44064 & w50260) | (~w44064 & w50261) | (w50260 & w50261);
assign w3252 = w3250 & ~w3251;
assign w3253 = ~w2895 & w51179;
assign w3254 = (a[90] & w2895) | (a[90] & w51180) | (w2895 & w51180);
assign w3255 = ~w3253 & ~w3254;
assign w3256 = a[90] & ~w3119;
assign w3257 = ~w3122 & ~w3256;
assign w3258 = w2558 & ~w3255;
assign w3259 = ~w3241 & w40030;
assign w3260 = ~w2557 & w51181;
assign w3261 = (w3260 & w3241) | (w3260 & w40031) | (w3241 & w40031);
assign w3262 = ~w3259 & ~w3261;
assign w3263 = ~w3252 & w3262;
assign w3264 = ~w3252 & w40032;
assign w3265 = ~w3138 & ~w3139;
assign w3266 = w2006 & w3155;
assign w3267 = w3265 & w3266;
assign w3268 = (w3267 & w3241) | (w3267 & w40033) | (w3241 & w40033);
assign w3269 = w2006 & ~w3155;
assign w3270 = ~w3265 & w3269;
assign w3271 = (w3269 & w2966) | (w3269 & w40034) | (w2966 & w40034);
assign w3272 = (~w3270 & w3241) | (~w3270 & w40035) | (w3241 & w40035);
assign w3273 = ~w3268 & w3272;
assign w3274 = a[91] & ~w3253;
assign w3275 = ~a[91] & w3253;
assign w3276 = ~w3274 & ~w3275;
assign w3277 = ~w2895 & w51182;
assign w3278 = (w2558 & w2895) | (w2558 & w51183) | (w2895 & w51183);
assign w3279 = ~w3277 & ~w3278;
assign w3280 = w3119 & w2824;
assign w3281 = ~w3130 & ~w3280;
assign w3282 = w3279 & ~w3281;
assign w3283 = ~w3279 & w3281;
assign w3284 = ~w3282 & ~w3283;
assign w3285 = ~w3241 & w40036;
assign w3286 = (w3284 & w3241) | (w3284 & w40037) | (w3241 & w40037);
assign w3287 = ~w3285 & ~w3286;
assign w3288 = (w3257 & w2557) | (w3257 & w51184) | (w2557 & w51184);
assign w3289 = w2285 & w3288;
assign w3290 = (w3289 & w3241) | (w3289 & w40038) | (w3241 & w40038);
assign w3291 = w3255 & w51185;
assign w3292 = ~w3241 & w40039;
assign w3293 = ~w3290 & ~w3292;
assign w3294 = ~w3287 & w3293;
assign w3295 = (~w2285 & ~w3255) | (~w2285 & w51186) | (~w3255 & w51186);
assign w3296 = ~w3241 & w40040;
assign w3297 = ~w2285 & ~w3288;
assign w3298 = (w3297 & w3241) | (w3297 & w40041) | (w3241 & w40041);
assign w3299 = ~w3296 & ~w3298;
assign w3300 = w3273 & ~w3299;
assign w3301 = ~w3263 & w3300;
assign w3302 = w3155 & w52152;
assign w3303 = (w3241 & w51187) | (w3241 & w51188) | (w51187 & w51188);
assign w3304 = ~w3302 & ~w3303;
assign w3305 = ~w2006 & ~w3304;
assign w3306 = ~w3301 & ~w3305;
assign w3307 = w3273 & w3294;
assign w3308 = ~w3264 & w3307;
assign w3309 = w3306 & ~w3308;
assign w3310 = (~w2006 & w3156) | (~w2006 & w40043) | (w3156 & w40043);
assign w3311 = ~w3156 & w40044;
assign w3312 = ~w1541 & ~w3311;
assign w3313 = (w3028 & w3312) | (w3028 & w51189) | (w3312 & w51189);
assign w3314 = (w3168 & w3160) | (w3168 & w51500) | (w3160 & w51500);
assign w3315 = w1738 & w3027;
assign w3316 = ~w3160 & w51190;
assign w3317 = ~w1541 & ~w3316;
assign w3318 = ~w3313 & w3314;
assign w3319 = ~w3161 & w3313;
assign w3320 = (~w3319 & w3318) | (~w3319 & w51191) | (w3318 & w51191);
assign w3321 = (~w44064 & w51378) | (~w44064 & w51379) | (w51378 & w51379);
assign w3322 = w3027 & w52153;
assign w3323 = ~w3241 & w40045;
assign w3324 = ~w3321 & ~w3323;
assign w3325 = ~w3310 & ~w3311;
assign w3326 = ~w3161 & w3325;
assign w3327 = w3161 & ~w3325;
assign w3328 = (w3116 & w47057) | (w3116 & w47058) | (w47057 & w47058);
assign w3329 = (~w47058 & w51193) | (~w47058 & w51194) | (w51193 & w51194);
assign w3330 = (~w1738 & w3312) | (~w1738 & w51195) | (w3312 & w51195);
assign w3331 = ~w3325 & w51380;
assign w3332 = w3330 & ~w3331;
assign w3333 = ~w3331 & w51196;
assign w3334 = ~w2967 & w3332;
assign w3335 = (~w3333 & w3241) | (~w3333 & w44065) | (w3241 & w44065);
assign w3336 = w3160 & ~w3328;
assign w3337 = (~w3328 & w2966) | (~w3328 & w40047) | (w2966 & w40047);
assign w3338 = (~w3336 & w3241) | (~w3336 & w40048) | (w3241 & w40048);
assign w3339 = ~w3335 & w3338;
assign w3340 = w3324 & ~w3339;
assign w3341 = (w3163 & w51198) | (w3163 & w51199) | (w51198 & w51199);
assign w3342 = (~w3163 & w51200) | (~w3163 & w51201) | (w51200 & w51201);
assign w3343 = ~w3341 & ~w3342;
assign w3344 = w3343 & ~w3242;
assign w3345 = w2811 & ~w3031;
assign w3346 = ~w2811 & w3031;
assign w3347 = ~w3345 & ~w3346;
assign w3348 = ~w1320 & ~w3347;
assign w3349 = (~w44064 & w51202) | (~w44064 & w51203) | (w51202 & w51203);
assign w3350 = ~w1320 & w3347;
assign w3351 = (w44064 & w51204) | (w44064 & w51205) | (w51204 & w51205);
assign w3352 = ~w3349 & ~w3351;
assign w3353 = w3324 & w51206;
assign w3354 = w3306 & w40051;
assign w3355 = w3049 & ~w3073;
assign w3356 = ~w3241 & w40052;
assign w3357 = (w3341 & w3241) | (w3341 & w40053) | (w3241 & w40053);
assign w3358 = ~w3356 & ~w3357;
assign w3359 = w40054 & ~w3242;
assign w3360 = w3358 & ~w3359;
assign w3361 = (~w1120 & ~w3049) | (~w1120 & w51207) | (~w3049 & w51207);
assign w3362 = (w3361 & ~w3358) | (w3361 & w51208) | (~w3358 & w51208);
assign w3363 = w3049 & w51209;
assign w3364 = w3358 & w51210;
assign w3365 = ~w3362 & ~w3364;
assign w3366 = ~w3241 & w40055;
assign w3367 = ~w3326 & ~w3327;
assign w3368 = (w3367 & w3241) | (w3367 & w40056) | (w3241 & w40056);
assign w3369 = ~w3366 & ~w3368;
assign w3370 = (w1738 & w3160) | (w1738 & w51211) | (w3160 & w51211);
assign w3371 = ~w3160 & w51212;
assign w3372 = ~w3370 & ~w3371;
assign w3373 = w1541 & ~w3027;
assign w3374 = w3373 & w52154;
assign w3375 = w1541 & w3027;
assign w3376 = (w3241 & w51213) | (w3241 & w51214) | (w51213 & w51214);
assign w3377 = ~w3374 & ~w3376;
assign w3378 = w1738 & w3369;
assign w3379 = w3377 & ~w3378;
assign w3380 = w3353 & ~w3379;
assign w3381 = w3344 & w3347;
assign w3382 = ~w3344 & ~w3347;
assign w3383 = ~w3381 & ~w3382;
assign w3384 = w1320 & ~w3383;
assign w3385 = ~w3067 & ~w3078;
assign w3386 = ~w2895 & w51215;
assign w3387 = ~w3071 & ~w3386;
assign w3388 = (~w3387 & w3036) | (~w3387 & w40058) | (w3036 & w40058);
assign w3389 = ~w3387 & w52155;
assign w3390 = ~w3163 & w3389;
assign w3391 = (w3385 & w3390) | (w3385 & w40059) | (w3390 & w40059);
assign w3392 = ~w3390 & w40060;
assign w3393 = ~w3391 & ~w3392;
assign w3394 = ~w945 & w3077;
assign w3395 = ~w3241 & w40061;
assign w3396 = ~w945 & ~w3393;
assign w3397 = ~w3242 & w3396;
assign w3398 = ~w3395 & ~w3397;
assign w3399 = w3365 & ~w3380;
assign w3400 = ~w3384 & w3398;
assign w3401 = w3399 & w3400;
assign w3402 = ~w3354 & w3401;
assign w3403 = w3049 & w51217;
assign w3404 = ~w3397 & w40062;
assign w3405 = ~w3360 & w3404;
assign w3406 = (w1120 & ~w3049) | (w1120 & w51218) | (~w3049 & w51218);
assign w3407 = ~w3397 & w40063;
assign w3408 = w3360 & w3407;
assign w3409 = ~w3405 & ~w3408;
assign w3410 = ~w3163 & w3171;
assign w3411 = ~w3075 & w3080;
assign w3412 = ~w3410 & w3411;
assign w3413 = w3014 & w3234;
assign w3414 = ~w3000 & ~w3413;
assign w3415 = (w3414 & w3412) | (w3414 & w40064) | (w3412 & w40064);
assign w3416 = (w3234 & w2999) | (w3234 & w47059) | (w2999 & w47059);
assign w3417 = ~w3082 & w3416;
assign w3418 = w3172 & w44066;
assign w3419 = (w3014 & w3417) | (w3014 & w51467) | (w3417 & w51467);
assign w3420 = ~w3415 & ~w3419;
assign w3421 = ~w3242 & w3420;
assign w3422 = ~w3008 & ~w3009;
assign w3423 = w3008 & w3009;
assign w3424 = ~w3422 & ~w3423;
assign w3425 = (~w3424 & w2966) | (~w3424 & w40065) | (w2966 & w40065);
assign w3426 = ~w3241 & w3425;
assign w3427 = ~w3421 & ~w3426;
assign w3428 = (~w493 & w3421) | (~w493 & w40066) | (w3421 & w40066);
assign w3429 = ~w3207 & ~w3235;
assign w3430 = ~w3417 & w51468;
assign w3431 = (~w3429 & w3417) | (~w3429 & w51469) | (w3417 & w51469);
assign w3432 = ~w3430 & ~w3431;
assign w3433 = ~w3242 & w3432;
assign w3434 = (w3206 & w2966) | (w3206 & w40067) | (w2966 & w40067);
assign w3435 = ~w3241 & w3434;
assign w3436 = (w400 & w3241) | (w400 & w40068) | (w3241 & w40068);
assign w3437 = ~w3433 & w3436;
assign w3438 = ~w2982 & ~w3000;
assign w3439 = (w3438 & w3412) | (w3438 & w40069) | (w3412 & w40069);
assign w3440 = ~w3412 & w40070;
assign w3441 = ~w3439 & ~w3440;
assign w3442 = ~w3242 & w3441;
assign w3443 = (w2981 & w2966) | (w2981 & w40071) | (w2966 & w40071);
assign w3444 = ~w3241 & w3443;
assign w3445 = (~w612 & w3241) | (~w612 & w40072) | (w3241 & w40072);
assign w3446 = ~w3442 & w3445;
assign w3447 = ~w3437 & ~w3446;
assign w3448 = ~w3428 & w3447;
assign w3449 = ~w3241 & w40073;
assign w3450 = (w3393 & w3241) | (w3393 & w40074) | (w3241 & w40074);
assign w3451 = ~w3449 & ~w3450;
assign w3452 = w945 & ~w3451;
assign w3453 = ~w2998 & ~w3079;
assign w3454 = (~w3078 & w3163) | (~w3078 & w40075) | (w3163 & w40075);
assign w3455 = w3074 & w52156;
assign w3456 = (w3453 & ~w3454) | (w3453 & w51220) | (~w3454 & w51220);
assign w3457 = w3454 & w51221;
assign w3458 = ~w3456 & ~w3457;
assign w3459 = w3458 & ~w3242;
assign w3460 = (~w754 & w3459) | (~w754 & w40077) | (w3459 & w40077);
assign w3461 = ~w3452 & ~w3460;
assign w3462 = w3448 & w3461;
assign w3463 = w3409 & w3462;
assign w3464 = (w3463 & ~w3401) | (w3463 & w40078) | (~w3401 & w40078);
assign w3465 = ~w3442 & ~w3444;
assign w3466 = (w612 & w3442) | (w612 & w40079) | (w3442 & w40079);
assign w3467 = ~w3459 & w40080;
assign w3468 = ~w3466 & ~w3467;
assign w3469 = w3448 & ~w3468;
assign w3470 = (~w400 & w3433) | (~w400 & w40081) | (w3433 & w40081);
assign w3471 = (w493 & w3241) | (w493 & w44067) | (w3241 & w44067);
assign w3472 = ~w3421 & w3471;
assign w3473 = ~w3437 & w3472;
assign w3474 = ~w3470 & ~w3473;
assign w3475 = ~w3469 & w3474;
assign w3476 = w3475 & ~w3464;
assign w3477 = (w3417 & w51501) | (w3417 & w51502) | (w51501 & w51502);
assign w3478 = (~w44064 & w51538) | (~w44064 & w51539) | (w51538 & w51539);
assign w3479 = ~w3190 & ~w3191;
assign w3480 = (w400 & w2966) | (w400 & w40083) | (w2966 & w40083);
assign w3481 = ~w3209 & ~w3236;
assign w3482 = (~w3209 & ~w3172) | (~w3209 & w47060) | (~w3172 & w47060);
assign w3483 = ~w3083 & w3482;
assign w3484 = ~w3483 & w40084;
assign w3485 = ~w3242 & w3484;
assign w3486 = ~w3241 & w40085;
assign w3487 = ~w3485 & ~w3486;
assign w3488 = (~w3479 & w3241) | (~w3479 & w40086) | (w3241 & w40086);
assign w3489 = ~w3478 & w3488;
assign w3490 = w3487 & ~w3489;
assign w3491 = w3487 & w51546;
assign w3492 = ~w2954 & w3221;
assign w3493 = ~w3173 & w3492;
assign w3494 = ~w3083 & w3493;
assign w3495 = ~w2954 & ~w3237;
assign w3496 = ~w3494 & ~w3495;
assign w3497 = (w3493 & w50262) | (w3493 & w50263) | (w50262 & w50263);
assign w3498 = (~w2936 & w3241) | (~w2936 & w40088) | (w3241 & w40088);
assign w3499 = ~w3497 & w3498;
assign w3500 = ~w3241 & w40089;
assign w3501 = ~w2944 & ~w2957;
assign w3502 = ~w3 & w3501;
assign w3503 = (w3502 & w3499) | (w3502 & w51222) | (w3499 & w51222);
assign w3504 = ~w3 & ~w3501;
assign w3505 = ~w3499 & w51223;
assign w3506 = ~w3503 & ~w3505;
assign w3507 = ~w2954 & ~w3229;
assign w3508 = w2945 & ~w3507;
assign w3509 = (~w2954 & ~w47056) | (~w2954 & w51224) | (~w47056 & w51224);
assign w3510 = w3221 & w3509;
assign w3511 = w3508 & ~w3510;
assign w3512 = (~w2946 & w2943) | (~w2946 & w51225) | (w2943 & w51225);
assign w3513 = ~w2944 & ~w3512;
assign w3514 = (~w3513 & w3494) | (~w3513 & w40091) | (w3494 & w40091);
assign w3515 = ~w3242 & ~w3514;
assign w3516 = ~w2876 & w2962;
assign w3517 = ~w3515 & w40092;
assign w3518 = (w3516 & w3515) | (w3516 & w40093) | (w3515 & w40093);
assign w3519 = ~w3517 & ~w3518;
assign w3520 = ~w42 & ~w3519;
assign w3521 = w3506 & ~w3520;
assign w3522 = (~w2630 & ~w2885) | (~w2630 & w51226) | (~w2885 & w51226);
assign w3523 = w2885 & w51227;
assign w3524 = ~w3522 & ~w3523;
assign w3525 = ~w3 & w3524;
assign w3526 = w42 & ~w2875;
assign w3527 = ~w3515 & w40095;
assign w3528 = (w3494 & w3534) | (w3494 & w47061) | (w3534 & w47061);
assign w3529 = ~w2876 & w51228;
assign w3530 = ~w3512 & w47062;
assign w3531 = w3529 & ~w3530;
assign w3532 = ~w3510 & w44068;
assign w3533 = (w3531 & w3494) | (w3531 & w44069) | (w3494 & w44069);
assign w3534 = w2962 & ~w3513;
assign w3535 = (~w2876 & w3513) | (~w2876 & w51229) | (w3513 & w51229);
assign w3536 = ~w2876 & w3511;
assign w3537 = (~w3535 & w3494) | (~w3535 & w51230) | (w3494 & w51230);
assign w3538 = w2921 & ~w3524;
assign w3539 = (w40096 & w3494) | (w40096 & w51231) | (w3494 & w51231);
assign w3540 = (~w42 & w3524) | (~w42 & w51232) | (w3524 & w51232);
assign w3541 = (w3540 & w40097) | (w3540 & w52157) | (w40097 & w52157);
assign w3542 = ~w3539 & ~w3541;
assign w3543 = ~w3242 & w51233;
assign w3544 = w3542 & ~w3543;
assign w3545 = ~w3527 & w3544;
assign w3546 = (~w3545 & w3520) | (~w3545 & w51234) | (w3520 & w51234);
assign w3547 = ~w3242 & w3496;
assign w3548 = ~w2936 & ~w2946;
assign w3549 = ~w80 & ~w3548;
assign w3550 = (w3549 & w3547) | (w3549 & w40099) | (w3547 & w40099);
assign w3551 = ~w80 & w3548;
assign w3552 = ~w3547 & w40100;
assign w3553 = ~w3550 & ~w3552;
assign w3554 = w80 & w3548;
assign w3555 = w3548 & w51235;
assign w3556 = ~w3241 & w40101;
assign w3557 = (w40102 & ~w3493) | (w40102 & w47063) | (~w3493 & w47063);
assign w3558 = ~w3242 & w3557;
assign w3559 = ~w3556 & ~w3558;
assign w3560 = w80 & ~w3548;
assign w3561 = (w3493 & w47064) | (w3493 & w47065) | (w47064 & w47065);
assign w3562 = ~w2935 & w33829;
assign w3563 = ~w3241 & w40104;
assign w3564 = ~w3242 & w3561;
assign w3565 = ~w3563 & ~w3564;
assign w3566 = w3559 & w3565;
assign w3567 = ~w3241 & w40105;
assign w3568 = w3229 & w52158;
assign w3569 = ~w3223 & w3568;
assign w3570 = ~w2954 & w3228;
assign w3571 = w3221 & ~w3570;
assign w3572 = ~w3173 & w3571;
assign w3573 = ~w3570 & w52159;
assign w3574 = (~w3573 & ~w3572) | (~w3573 & w47066) | (~w3572 & w47066);
assign w3575 = ~w3569 & w3574;
assign w3576 = ~w3242 & w3575;
assign w3577 = (w57 & w3576) | (w57 & w40107) | (w3576 & w40107);
assign w3578 = w3566 & w3577;
assign w3579 = w3553 & ~w3578;
assign w3580 = w3 & w3501;
assign w3581 = (w3580 & w3241) | (w3580 & w44070) | (w3241 & w44070);
assign w3582 = ~w3499 & w3581;
assign w3583 = w3 & ~w3501;
assign w3584 = w3583 & ~w3497;
assign w3585 = w3498 & w3584;
assign w3586 = ~w3241 & w44071;
assign w3587 = ~w3585 & ~w3586;
assign w3588 = ~w3582 & w3587;
assign w3589 = ~w3545 & w3588;
assign w3590 = w3579 & w3589;
assign w3591 = ~w3220 & ~w3224;
assign w3592 = ~w3483 & w40108;
assign w3593 = (w3591 & w3483) | (w3591 & w40109) | (w3483 & w40109);
assign w3594 = ~w3592 & ~w3593;
assign w3595 = ~w2967 & w52160;
assign w3596 = ~w3242 & ~w3594;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = ~w3596 & w51238;
assign w3599 = ~w3238 & w47067;
assign w3600 = w3237 & w3599;
assign w3601 = ~w3223 & w3600;
assign w3602 = ~w57 & ~w3601;
assign w3603 = ~w3567 & w3602;
assign w3604 = w2967 & w3575;
assign w3605 = w3603 & ~w3604;
assign w3606 = w3566 & ~w3605;
assign w3607 = w3566 & w51239;
assign w3608 = w3579 & w51240;
assign w3609 = ~w3608 & w40111;
assign w3610 = (w3491 & w3608) | (w3491 & w47068) | (w3608 & w47068);
assign w3611 = w3476 & w3610;
assign w3612 = (w3491 & w3608) | (w3491 & w47069) | (w3608 & w47069);
assign w3613 = ~w3476 & w3612;
assign w3614 = ~w3611 & ~w3613;
assign w3615 = (w252 & w3596) | (w252 & w51241) | (w3596 & w51241);
assign w3616 = w3487 & w51540;
assign w3617 = (~w3615 & ~w3490) | (~w3615 & w51242) | (~w3490 & w51242);
assign w3618 = w3607 & ~w3617;
assign w3619 = w3590 & ~w3618;
assign w3620 = (~w3546 & ~w3590) | (~w3546 & w51243) | (~w3590 & w51243);
assign w3621 = (w351 & ~w3487) | (w351 & w51541) | (~w3487 & w51541);
assign w3622 = ~w3619 & w40112;
assign w3623 = (~w351 & ~w3487) | (~w351 & w51547) | (~w3487 & w51547);
assign w3624 = ~w3619 & w40113;
assign w3625 = ~w3619 & w47070;
assign w3626 = w3476 & w3625;
assign w3627 = ~w3619 & w47071;
assign w3628 = ~w3476 & w3627;
assign w3629 = ~w3626 & ~w3628;
assign w3630 = w3614 & w3629;
assign w3631 = (w3490 & w3608) | (w3490 & w47072) | (w3608 & w47072);
assign w3632 = w3476 & ~w3622;
assign w3633 = w3490 & ~w3609;
assign w3634 = w3632 & ~w3633;
assign w3635 = ~w3476 & w47073;
assign w3636 = ~w3634 & ~w3635;
assign w3637 = (~w252 & w3634) | (~w252 & w47074) | (w3634 & w47074);
assign w3638 = w3630 & ~w3637;
assign w3639 = ~w3578 & w40114;
assign w3640 = w3474 & ~w3621;
assign w3641 = ~w3469 & w3640;
assign w3642 = w3521 & w3641;
assign w3643 = ~w3607 & w3639;
assign w3644 = w3642 & ~w3643;
assign w3645 = ~w3464 & w3644;
assign w3646 = (~w3620 & w3464) | (~w3620 & w44072) | (w3464 & w44072);
assign w3647 = w3409 & w3461;
assign w3648 = ~w3442 & w51244;
assign w3649 = w3409 & w44073;
assign w3650 = (w493 & w3442) | (w493 & w51245) | (w3442 & w51245);
assign w3651 = ~w3427 & ~w3650;
assign w3652 = w3649 & ~w3651;
assign w3653 = ~w3468 & w51246;
assign w3654 = ~w3472 & ~w3653;
assign w3655 = (w3654 & w3402) | (w3654 & w40115) | (w3402 & w40115);
assign w3656 = w3655 & ~w3646;
assign w3657 = w400 & ~w3620;
assign w3658 = ~w3437 & ~w3470;
assign w3659 = ~w3656 & w47075;
assign w3660 = (w3658 & w3656) | (w3658 & w47076) | (w3656 & w47076);
assign w3661 = ~w3659 & ~w3660;
assign w3662 = ~w351 & w3661;
assign w3663 = ~w3468 & w3650;
assign w3664 = w3409 & w44074;
assign w3665 = (~w40117 & w44075) | (~w40117 & w44076) | (w44075 & w44076);
assign w3666 = (~w493 & w3468) | (~w493 & w51247) | (w3468 & w51247);
assign w3667 = (~w40116 & w44077) | (~w40116 & w44078) | (w44077 & w44078);
assign w3668 = w3665 & ~w3667;
assign w3669 = (w400 & w3421) | (w400 & w51248) | (w3421 & w51248);
assign w3670 = (w3669 & w3646) | (w3669 & w48594) | (w3646 & w48594);
assign w3671 = ~w3421 & w51249;
assign w3672 = ~w3646 & w48595;
assign w3673 = ~w3670 & ~w3672;
assign w3674 = ~w3446 & ~w3466;
assign w3675 = w3467 & ~w3674;
assign w3676 = w3409 & w44079;
assign w3677 = (~w40119 & w44080) | (~w40119 & w44081) | (w44080 & w44081);
assign w3678 = w3468 & w52161;
assign w3679 = w3677 & ~w3678;
assign w3680 = w3446 & ~w3467;
assign w3681 = (~w40118 & w51250) | (~w40118 & w51251) | (w51250 & w51251);
assign w3682 = (w3465 & w3619) | (w3465 & w48596) | (w3619 & w48596);
assign w3683 = (~w3681 & w3645) | (~w3681 & w51252) | (w3645 & w51252);
assign w3684 = ~w3646 & w3679;
assign w3685 = w3683 & ~w3684;
assign w3686 = ~w3684 & w51253;
assign w3687 = w3673 & w3686;
assign w3688 = ~w754 & ~w3620;
assign w3689 = ~w3645 & w3688;
assign w3690 = w3409 & ~w3452;
assign w3691 = ~w3402 & w3690;
assign w3692 = ~w3691 & ~w3646;
assign w3693 = ~w3460 & ~w3467;
assign w3694 = ~w612 & ~w3693;
assign w3695 = (w3694 & w3692) | (w3694 & w48597) | (w3692 & w48597);
assign w3696 = ~w612 & w3693;
assign w3697 = ~w3692 & w48598;
assign w3698 = ~w3695 & ~w3697;
assign w3699 = (~w493 & w3684) | (~w493 & w51254) | (w3684 & w51254);
assign w3700 = w3673 & ~w3699;
assign w3701 = w3698 & w3700;
assign w3702 = w612 & w3693;
assign w3703 = (w3702 & w3692) | (w3702 & w48599) | (w3692 & w48599);
assign w3704 = w612 & ~w3693;
assign w3705 = (w3704 & w3645) | (w3704 & w44082) | (w3645 & w44082);
assign w3706 = ~w3692 & w3705;
assign w3707 = (w3355 & ~w3358) | (w3355 & w51255) | (~w3358 & w51255);
assign w3708 = w3358 & w51256;
assign w3709 = ~w3707 & ~w3708;
assign w3710 = (~w945 & w3451) | (~w945 & w51257) | (w3451 & w51257);
assign w3711 = w754 & w3451;
assign w3712 = (~w3711 & ~w3709) | (~w3711 & w51258) | (~w3709 & w51258);
assign w3713 = ~w3380 & ~w3384;
assign w3714 = ~w3354 & w3713;
assign w3715 = w1120 & ~w3709;
assign w3716 = w3365 & ~w3715;
assign w3717 = (w3716 & w3354) | (w3716 & w51259) | (w3354 & w51259);
assign w3718 = w3398 & ~w3452;
assign w3719 = ~w3365 & ~w3718;
assign w3720 = w3365 & w3718;
assign w3721 = ~w3719 & ~w3720;
assign w3722 = w754 & ~w3718;
assign w3723 = ~w3714 & w44083;
assign w3724 = w754 & ~w3721;
assign w3725 = ~w3717 & w3724;
assign w3726 = ~w3723 & ~w3725;
assign w3727 = w3712 & w3646;
assign w3728 = ~w3646 & w3726;
assign w3729 = ~w3727 & ~w3728;
assign w3730 = ~w3706 & ~w3729;
assign w3731 = ~w3703 & w3730;
assign w3732 = ~w3354 & w51260;
assign w3733 = ~w3717 & ~w3732;
assign w3734 = (~w44072 & w51261) | (~w44072 & w51262) | (w51261 & w51262);
assign w3735 = w3709 & w3646;
assign w3736 = ~w3734 & ~w3735;
assign w3737 = ~w3734 & w48600;
assign w3738 = ~w3714 & w44084;
assign w3739 = (w3721 & w3714) | (w3721 & w44085) | (w3714 & w44085);
assign w3740 = ~w3738 & ~w3739;
assign w3741 = ~w3451 & w3646;
assign w3742 = ~w3646 & ~w3740;
assign w3743 = ~w3741 & ~w3742;
assign w3744 = (~w754 & w3742) | (~w754 & w48601) | (w3742 & w48601);
assign w3745 = ~w3737 & ~w3744;
assign w3746 = w3731 & ~w3745;
assign w3747 = w3701 & ~w3746;
assign w3748 = (~w3687 & w3746) | (~w3687 & w51263) | (w3746 & w51263);
assign w3749 = ~a[84] & ~a[85];
assign w3750 = ~a[86] & w3749;
assign w3751 = w3750 & ~w3242;
assign w3752 = ~w2967 & w52162;
assign w3753 = ~w3751 & ~w3752;
assign w3754 = ~a[87] & w3753;
assign w3755 = (~w3751 & ~w3753) | (~w3751 & w51265) | (~w3753 & w51265);
assign w3756 = (w3755 & w3619) | (w3755 & w48602) | (w3619 & w48602);
assign w3757 = ~w3645 & w3756;
assign w3758 = a[86] & ~a[87];
assign w3759 = ~w3751 & ~w3758;
assign w3760 = w3642 & w40121;
assign w3761 = ~w3464 & w3760;
assign w3762 = w3759 & w52163;
assign w3763 = ~w3761 & ~w3762;
assign w3764 = ~w3757 & w3763;
assign w3765 = a[87] & w3753;
assign w3766 = w3620 & w3765;
assign w3767 = w3642 & w40122;
assign w3768 = ~w3464 & w3767;
assign w3769 = (w2896 & w3764) | (w2896 & w44086) | (w3764 & w44086);
assign w3770 = ~w2967 & w52164;
assign w3771 = ~a[88] & ~w3242;
assign w3772 = a[88] & ~w3243;
assign w3773 = ~w3244 & ~w3772;
assign w3774 = ~w3770 & ~w3771;
assign w3775 = ~w3620 & w52165;
assign w3776 = w3773 & ~w3646;
assign w3777 = ~w3775 & ~w3776;
assign w3778 = ~w3769 & w3777;
assign w3779 = ~a[89] & w52166;
assign w3780 = w3642 & w40124;
assign w3781 = ~w3464 & w3780;
assign w3782 = ~w3779 & ~w3781;
assign w3783 = ~w3245 & ~w3247;
assign w3784 = w3783 & ~w3242;
assign w3785 = ~w2967 & w52167;
assign w3786 = ~w3784 & ~w3785;
assign w3787 = w3786 & w52168;
assign w3788 = w3642 & w40126;
assign w3789 = ~w3464 & w3788;
assign w3790 = ~w3787 & ~w3789;
assign w3791 = ~w3782 & w3790;
assign w3792 = a[89] & w3786;
assign w3793 = w3792 & w52168;
assign w3794 = w3642 & w40127;
assign w3795 = ~w3464 & w3794;
assign w3796 = ~w3793 & ~w3795;
assign w3797 = a[89] & w3771;
assign w3798 = (w3797 & w3619) | (w3797 & w40128) | (w3619 & w40128);
assign w3799 = (w3798 & w3464) | (w3798 & w44087) | (w3464 & w44087);
assign w3800 = w3796 & ~w3799;
assign w3801 = ~w3791 & w3800;
assign w3802 = w3095 & ~w3801;
assign w3803 = w3778 & ~w3802;
assign w3804 = ~w3768 & w44088;
assign w3805 = ~w3764 & w3804;
assign w3806 = (~w2558 & w3764) | (~w2558 & w44089) | (w3764 & w44089);
assign w3807 = w3801 & ~w3806;
assign w3808 = (w2285 & w3764) | (w2285 & w51269) | (w3764 & w51269);
assign w3809 = ~w3807 & w3808;
assign w3810 = ~w3803 & w3809;
assign w3811 = ~w2558 & w3252;
assign w3812 = w2558 & ~w3252;
assign w3813 = ~w3811 & ~w3812;
assign w3814 = w3642 & w40129;
assign w3815 = ~w3464 & w3814;
assign w3816 = ~w2967 & w52169;
assign w3817 = w3257 & ~w3242;
assign w3818 = ~w3816 & ~w3817;
assign w3819 = ~w3815 & w44091;
assign w3820 = (~w3818 & w3815) | (~w3818 & w44092) | (w3815 & w44092);
assign w3821 = ~w3819 & ~w3820;
assign w3822 = w2558 & ~w3798;
assign w3823 = w3642 & w40130;
assign w3824 = ~w3464 & w3823;
assign w3825 = ~w3822 & ~w3824;
assign w3826 = w3796 & ~w3825;
assign w3827 = ~w3791 & w3826;
assign w3828 = ~w3805 & ~w3827;
assign w3829 = ~w2285 & w3801;
assign w3830 = ~w2807 & w3821;
assign w3831 = ~w3263 & ~w3299;
assign w3832 = ~w3264 & ~w3831;
assign w3833 = w3293 & w3832;
assign w3834 = (w44072 & w51470) | (w44072 & w51471) | (w51470 & w51471);
assign w3835 = (~w44072 & w51472) | (~w44072 & w51473) | (w51472 & w51473);
assign w3836 = ~w3834 & ~w3835;
assign w3837 = w2006 & ~w3836;
assign w3838 = (~w3837 & w3829) | (~w3837 & w51474) | (w3829 & w51474);
assign w3839 = w3821 & w3828;
assign w3840 = ~w3778 & w3839;
assign w3841 = w3838 & ~w3840;
assign w3842 = ~w3810 & w3841;
assign w3843 = w3306 & w40131;
assign w3844 = ~w1738 & ~w3309;
assign w3845 = ~w3843 & ~w3844;
assign w3846 = w3369 & w3845;
assign w3847 = (~w44072 & w47077) | (~w44072 & w47078) | (w47077 & w47078);
assign w3848 = (~w44072 & w50266) | (~w44072 & w50267) | (w50266 & w50267);
assign w3849 = ~w1541 & w3847;
assign w3850 = ~w1541 & ~w3369;
assign w3851 = ~w3848 & w3850;
assign w3852 = ~w3849 & ~w3851;
assign w3853 = (~w3369 & ~w40131) | (~w3369 & w44093) | (~w40131 & w44093);
assign w3854 = ~w3844 & ~w3853;
assign w3855 = w1541 & ~w3854;
assign w3856 = ~w1541 & w3854;
assign w3857 = ~w3855 & ~w3856;
assign w3858 = w3027 & w52154;
assign w3859 = (w3241 & w51271) | (w3241 & w51272) | (w51271 & w51272);
assign w3860 = ~w3858 & ~w3859;
assign w3861 = ~w1320 & ~w3860;
assign w3862 = (w3861 & w3646) | (w3861 & w47079) | (w3646 & w47079);
assign w3863 = ~w1320 & w3860;
assign w3864 = ~w3646 & w47080;
assign w3865 = ~w3862 & ~w3864;
assign w3866 = w3852 & w3865;
assign w3867 = ~w2006 & w3836;
assign w3868 = ~w3294 & ~w3831;
assign w3869 = (w2006 & w3868) | (w2006 & w51273) | (w3868 & w51273);
assign w3870 = ~w3868 & w51274;
assign w3871 = ~w3869 & ~w3870;
assign w3872 = ~w3620 & w3871;
assign w3873 = w3304 & ~w3871;
assign w3874 = ~w3304 & w3871;
assign w3875 = ~w3873 & ~w3874;
assign w3876 = (~w3875 & w3645) | (~w3875 & w51275) | (w3645 & w51275);
assign w3877 = ~w3645 & w44094;
assign w3878 = ~w3876 & ~w3877;
assign w3879 = ~w1738 & w3878;
assign w3880 = ~w3867 & ~w3879;
assign w3881 = w3866 & w3880;
assign w3882 = w1320 & w52170;
assign w3883 = (w3309 & w51277) | (w3309 & w51278) | (w51277 & w51278);
assign w3884 = ~w3882 & ~w3883;
assign w3885 = (w44072 & w51503) | (w44072 & w51504) | (w51503 & w51504);
assign w3886 = (~w44072 & w51505) | (~w44072 & w51506) | (w51505 & w51506);
assign w3887 = ~w3885 & ~w3886;
assign w3888 = w1120 & w3887;
assign w3889 = w3880 & w51279;
assign w3890 = (w3889 & ~w3841) | (w3889 & w51280) | (~w3841 & w51280);
assign w3891 = ~w3748 & w3890;
assign w3892 = w1541 & ~w3847;
assign w3893 = ~w3369 & ~w3848;
assign w3894 = w3892 & ~w3893;
assign w3895 = (w1738 & w3876) | (w1738 & w44095) | (w3876 & w44095);
assign w3896 = ~w3894 & ~w3895;
assign w3897 = w3866 & ~w3896;
assign w3898 = ~w1120 & ~w3887;
assign w3899 = ~w3646 & w47083;
assign w3900 = (w3860 & w3646) | (w3860 & w47084) | (w3646 & w47084);
assign w3901 = ~w3899 & ~w3900;
assign w3902 = w1320 & ~w3901;
assign w3903 = ~w3898 & ~w3902;
assign w3904 = ~w3897 & w3903;
assign w3905 = ~w3888 & ~w3904;
assign w3906 = ~w3748 & w3905;
assign w3907 = w351 & ~w3658;
assign w3908 = (w3907 & w3645) | (w3907 & w44096) | (w3645 & w44096);
assign w3909 = ~w3656 & w3908;
assign w3910 = w351 & w3658;
assign w3911 = (w3402 & w47085) | (w3402 & w47086) | (w47085 & w47086);
assign w3912 = ~w3646 & w3911;
assign w3913 = ~w3645 & w44097;
assign w3914 = ~w3912 & ~w3913;
assign w3915 = ~w3909 & w3914;
assign w3916 = (~w3427 & w3646) | (~w3427 & w51281) | (w3646 & w51281);
assign w3917 = ~w400 & ~w3916;
assign w3918 = ~w3646 & w51282;
assign w3919 = w3917 & ~w3918;
assign w3920 = ~w3687 & ~w3919;
assign w3921 = ~w754 & ~w3740;
assign w3922 = w3734 & w48603;
assign w3923 = w3730 & w44098;
assign w3924 = w3701 & ~w3923;
assign w3925 = w3920 & ~w3924;
assign w3926 = ~w3924 & w44099;
assign w3927 = ~w3906 & w3926;
assign w3928 = ~w3891 & w3927;
assign w3929 = ~w3662 & ~w3928;
assign w3930 = (w3638 & w3928) | (w3638 & w44100) | (w3928 & w44100);
assign w3931 = (w3881 & ~w3841) | (w3881 & w44101) | (~w3841 & w44101);
assign w3932 = w3904 & ~w3931;
assign w3933 = (~w3746 & w51283) | (~w3746 & w51284) | (w51283 & w51284);
assign w3934 = (~w3598 & w3616) | (~w3598 & w40132) | (w3616 & w40132);
assign w3935 = w3462 & w51542;
assign w3936 = ~w3402 & w3935;
assign w3937 = (w3607 & w3641) | (w3607 & w3618) | (w3641 & w3618);
assign w3938 = (w3937 & w3402) | (w3937 & w40133) | (w3402 & w40133);
assign w3939 = ~w3619 & w48604;
assign w3940 = w3642 & w40134;
assign w3941 = ~w3464 & w3940;
assign w3942 = ~w3939 & ~w3941;
assign w3943 = (~w3938 & w3941) | (~w3938 & w44102) | (w3941 & w44102);
assign w3944 = w3506 & w3588;
assign w3945 = w3944 & ~w3938;
assign w3946 = ~w3942 & w3945;
assign w3947 = (~w3944 & w3645) | (~w3944 & w44103) | (w3645 & w44103);
assign w3948 = ~w3943 & w3947;
assign w3949 = ~w3645 & w44104;
assign w3950 = ~w3946 & ~w3949;
assign w3951 = ~w3948 & w3950;
assign w3952 = w3506 & ~w3639;
assign w3953 = (~w3952 & w3936) | (~w3952 & w40135) | (w3936 & w40135);
assign w3954 = w3519 & w3620;
assign w3955 = w3642 & w40136;
assign w3956 = ~w3464 & w3955;
assign w3957 = ~w3954 & ~w3956;
assign w3958 = (w42 & w3957) | (w42 & w44105) | (w3957 & w44105);
assign w3959 = ~w3646 & w51285;
assign w3960 = w3958 & ~w3959;
assign w3961 = w3524 & w3537;
assign w3962 = ~w3537 & w3538;
assign w3963 = ~w3961 & ~w3962;
assign w3964 = (w3936 & w47087) | (w3936 & w47088) | (w47087 & w47088);
assign w3965 = ~w3519 & ~w3963;
assign w3966 = (~w3936 & w50268) | (~w3936 & w50269) | (w50268 & w50269);
assign w3967 = ~w3964 & ~w3966;
assign w3968 = ~w42 & w3967;
assign w3969 = (~w3968 & ~w3951) | (~w3968 & w44106) | (~w3951 & w44106);
assign w3970 = w3951 & w3968;
assign w3971 = ~w3577 & ~w3605;
assign w3972 = w3463 & w40137;
assign w3973 = ~w3402 & w3972;
assign w3974 = w3598 & w3971;
assign w3975 = ~w3616 & w40138;
assign w3976 = (~w3974 & w3641) | (~w3974 & w40139) | (w3641 & w40139);
assign w3977 = ~w3605 & w3976;
assign w3978 = ~w3973 & w3977;
assign w3979 = ~w3646 & ~w3978;
assign w3980 = w80 & ~w3620;
assign w3981 = ~w3645 & w3980;
assign w3982 = w3553 & w3566;
assign w3983 = w3 & ~w3982;
assign w3984 = (w3983 & w3645) | (w3983 & w44107) | (w3645 & w44107);
assign w3985 = ~w3979 & w3984;
assign w3986 = w3 & w3982;
assign w3987 = ~w3645 & w44108;
assign w3988 = (w3986 & w3973) | (w3986 & w40140) | (w3973 & w40140);
assign w3989 = ~w3646 & w3988;
assign w3990 = ~w3987 & ~w3989;
assign w3991 = ~w3985 & w3990;
assign w3992 = (~w3991 & ~w3951) | (~w3991 & w44109) | (~w3951 & w44109);
assign w3993 = ~w3969 & ~w3992;
assign w3994 = ~w57 & ~w3605;
assign w3995 = ~w3577 & ~w3994;
assign w3996 = ~w3598 & ~w3971;
assign w3997 = (w3996 & w3641) | (w3996 & w51286) | (w3641 & w51286);
assign w3998 = ~w3936 & w3997;
assign w3999 = (w3976 & w3402) | (w3976 & w40141) | (w3402 & w40141);
assign w4000 = ~w3998 & w3999;
assign w4001 = ~w3620 & w52171;
assign w4002 = ~w3646 & w4000;
assign w4003 = ~w4001 & ~w4002;
assign w4004 = ~w4002 & w40142;
assign w4005 = ~w3616 & ~w3641;
assign w4006 = w3462 & w47089;
assign w4007 = (~w4005 & w3402) | (~w4005 & w40143) | (w3402 & w40143);
assign w4008 = ~w3598 & ~w3615;
assign w4009 = ~w4008 & w52172;
assign w4010 = ~w4007 & w4009;
assign w4011 = w4008 & w52172;
assign w4012 = w4007 & w4011;
assign w4013 = ~w4010 & ~w4012;
assign w4014 = w3597 & ~w3620;
assign w4015 = (w57 & w3645) | (w57 & w44110) | (w3645 & w44110);
assign w4016 = w4013 & w4015;
assign w4017 = w3630 & ~w4016;
assign w4018 = ~w4004 & w4017;
assign w4019 = ~w3662 & w4018;
assign w4020 = ~w3637 & w3915;
assign w4021 = w4018 & ~w4020;
assign w4022 = (w80 & w4002) | (w80 & w47090) | (w4002 & w47090);
assign w4023 = (~w57 & ~w4013) | (~w57 & w47091) | (~w4013 & w47091);
assign w4024 = ~w4004 & w4023;
assign w4025 = ~w4022 & ~w4024;
assign w4026 = ~w4021 & w4025;
assign w4027 = ~w4019 & w4026;
assign w4028 = ~w4027 & w51288;
assign w4029 = ~w3932 & w4028;
assign w4030 = ~w3 & w3982;
assign w4031 = (w4030 & w3645) | (w4030 & w44111) | (w3645 & w44111);
assign w4032 = ~w3979 & w4031;
assign w4033 = ~w3 & ~w3982;
assign w4034 = ~w3645 & w44112;
assign w4035 = (w4033 & w3973) | (w4033 & w40145) | (w3973 & w40145);
assign w4036 = ~w3646 & w4035;
assign w4037 = ~w4034 & ~w4036;
assign w4038 = ~w4032 & w4037;
assign w4039 = (w4038 & ~w3951) | (w4038 & w44113) | (~w3951 & w44113);
assign w4040 = (w3630 & w4039) | (w3630 & w51289) | (w4039 & w51289);
assign w4041 = (w4019 & w3924) | (w4019 & w44114) | (w3924 & w44114);
assign w4042 = ~w3993 & w4040;
assign w4043 = w4026 & w4040;
assign w4044 = ~w4041 & w4043;
assign w4045 = ~w4042 & ~w4044;
assign w4046 = ~w4029 & ~w4045;
assign w4047 = ~w3930 & w4046;
assign w4048 = ~w3991 & w4038;
assign w4049 = ~w3970 & w4048;
assign w4050 = ~w3969 & ~w4049;
assign w4051 = w4026 & w4039;
assign w4052 = w4019 & w4050;
assign w4053 = ~w3925 & w4052;
assign w4054 = w4050 & ~w4051;
assign w4055 = ~w4053 & ~w4054;
assign w4056 = ~w4029 & w4055;
assign w4057 = (~w57 & w4029) | (~w57 & w40146) | (w4029 & w40146);
assign w4058 = ~w4016 & ~w4023;
assign w4059 = w80 & w4058;
assign w4060 = w4059 & ~w4057;
assign w4061 = ~w4047 & w4060;
assign w4062 = w80 & ~w4058;
assign w4063 = w4046 & w4062;
assign w4064 = ~w3930 & w4063;
assign w4065 = (w40146 & w51290) | (w40146 & w51291) | (w51290 & w51291);
assign w4066 = ~w4064 & ~w4065;
assign w4067 = ~w4061 & w4066;
assign w4068 = w4018 & w51507;
assign w4069 = ~w4004 & ~w4022;
assign w4070 = w3637 & ~w4016;
assign w4071 = ~w4023 & ~w4070;
assign w4072 = w4069 & ~w4071;
assign w4073 = (~w4072 & w3928) | (~w4072 & w40147) | (w3928 & w40147);
assign w4074 = (~w3888 & w4021) | (~w3888 & w51292) | (w4021 & w51292);
assign w4075 = w4018 & w51475;
assign w4076 = (~w44115 & w51293) | (~w44115 & w51294) | (w51293 & w51294);
assign w4077 = ~w3904 & w3993;
assign w4078 = ~w3992 & w51476;
assign w4079 = (~w4077 & w3842) | (~w4077 & w44116) | (w3842 & w44116);
assign w4080 = ~w4076 & ~w4079;
assign w4081 = (~w4003 & w4080) | (~w4003 & w40149) | (w4080 & w40149);
assign w4082 = ~w4073 & ~w4081;
assign w4083 = ~w4069 & w4071;
assign w4084 = ~w4053 & w44117;
assign w4085 = ~w4029 & w4084;
assign w4086 = ~w3662 & w4017;
assign w4087 = ~w3928 & w4086;
assign w4088 = w4085 & ~w4087;
assign w4089 = (w4003 & w4029) | (w4003 & w40150) | (w4029 & w40150);
assign w4090 = ~w4088 & ~w4089;
assign w4091 = ~w4082 & w4090;
assign w4092 = w4090 & w40151;
assign w4093 = w4067 & ~w4092;
assign w4094 = ~w80 & ~w4058;
assign w4095 = w4094 & ~w4057;
assign w4096 = ~w4047 & w4095;
assign w4097 = ~w80 & w4058;
assign w4098 = w4046 & w4097;
assign w4099 = ~w3930 & w4098;
assign w4100 = (w40146 & w51295) | (w40146 & w51296) | (w51295 & w51296);
assign w4101 = ~w4099 & ~w4100;
assign w4102 = ~w4096 & w4101;
assign w4103 = ~w4053 & w44118;
assign w4104 = w252 & ~w3636;
assign w4105 = (~w4104 & w4080) | (~w4104 & w51297) | (w4080 & w51297);
assign w4106 = ~w3638 & ~w3662;
assign w4107 = ~w3928 & w4106;
assign w4108 = (w3636 & w4029) | (w3636 & w40152) | (w4029 & w40152);
assign w4109 = w4056 & ~w4107;
assign w4110 = ~w4108 & ~w4109;
assign w4111 = ~w4110 & w44119;
assign w4112 = w4102 & ~w4111;
assign w4113 = w4093 & ~w4112;
assign w4114 = (w3 & ~w4090) | (w3 & w40153) | (~w4090 & w40153);
assign w4115 = w3991 & w4038;
assign w4116 = ~w3932 & ~w4076;
assign w4117 = (w4026 & w3925) | (w4026 & w4027) | (w3925 & w4027);
assign w4118 = (w4115 & w4116) | (w4115 & w40154) | (w4116 & w40154);
assign w4119 = w4026 & w52173;
assign w4120 = ~w4116 & w4119;
assign w4121 = (w3982 & w3979) | (w3982 & w51299) | (w3979 & w51299);
assign w4122 = ~w3979 & w51300;
assign w4123 = ~w4121 & ~w4122;
assign w4124 = ~w4056 & w4123;
assign w4125 = w4056 & ~w4120;
assign w4126 = ~w4118 & w4125;
assign w4127 = ~w4124 & ~w4126;
assign w4128 = (~w42 & w4126) | (~w42 & w40155) | (w4126 & w40155);
assign w4129 = ~w42 & w3951;
assign w4130 = w42 & ~w3951;
assign w4131 = ~w4129 & ~w4130;
assign w4132 = ~w3960 & w4131;
assign w4133 = w4132 & w52174;
assign w4134 = ~w3968 & ~w4131;
assign w4135 = (w50271 & w51301) | (w50271 & w51302) | (w51301 & w51302);
assign w4136 = ~w4133 & ~w4135;
assign w4137 = ~w4126 & w40156;
assign w4138 = w4136 & ~w4137;
assign w4139 = w4114 & ~w4128;
assign w4140 = w4138 & ~w4139;
assign w4141 = ~w4113 & w4140;
assign w4142 = ~w3906 & w3925;
assign w4143 = ~w3891 & w4142;
assign w4144 = ~w3662 & w3915;
assign w4145 = w4143 & ~w4144;
assign w4146 = ~w4143 & w4144;
assign w4147 = ~w3661 & ~w4056;
assign w4148 = w4056 & ~w4145;
assign w4149 = ~w4146 & w4148;
assign w4150 = ~w4147 & ~w4149;
assign w4151 = (w40157 & ~w4148) | (w40157 & w44120) | (~w4148 & w44120);
assign w4152 = (w3923 & w3904) | (w3923 & w40158) | (w3904 & w40158);
assign w4153 = (w4152 & w3842) | (w4152 & w44121) | (w3842 & w44121);
assign w4154 = (w3698 & ~w3731) | (w3698 & w51303) | (~w3731 & w51303);
assign w4155 = ~w3699 & w4154;
assign w4156 = (w4155 & w3890) | (w4155 & w40159) | (w3890 & w40159);
assign w4157 = (~w3686 & w4039) | (~w3686 & w51304) | (w4039 & w51304);
assign w4158 = ~w3993 & w4157;
assign w4159 = w4026 & w4157;
assign w4160 = ~w4041 & w4159;
assign w4161 = ~w4158 & ~w4160;
assign w4162 = ~w4029 & ~w4156;
assign w4163 = ~w4161 & w4162;
assign w4164 = (~w351 & w3919) | (~w351 & w51305) | (w3919 & w51305);
assign w4165 = (w4164 & w4163) | (w4164 & w40161) | (w4163 & w40161);
assign w4166 = ~w3919 & w51306;
assign w4167 = ~w4163 & w40162;
assign w4168 = ~w4165 & ~w4167;
assign w4169 = ~w4151 & w4168;
assign w4170 = ~w3919 & w51307;
assign w4171 = (w4170 & w4163) | (w4170 & w40163) | (w4163 & w40163);
assign w4172 = (w351 & w3919) | (w351 & w51308) | (w3919 & w51308);
assign w4173 = ~w4163 & w40164;
assign w4174 = ~w4171 & ~w4173;
assign w4175 = ~w3686 & ~w3699;
assign w4176 = ~w4175 & w50182;
assign w4177 = w4154 & w4175;
assign w4178 = ~w4153 & w4177;
assign w4179 = (w3685 & w4029) | (w3685 & w48605) | (w4029 & w48605);
assign w4180 = w4056 & w40166;
assign w4181 = ~w4179 & ~w4180;
assign w4182 = ~w4180 & w48606;
assign w4183 = w4174 & w4182;
assign w4184 = w4169 & ~w4183;
assign w4185 = ~w4113 & w47092;
assign w4186 = ~w3742 & w51309;
assign w4187 = ~w3744 & ~w4186;
assign w4188 = ~w945 & ~w3736;
assign w4189 = (~w3842 & w44122) | (~w3842 & w44123) | (w44122 & w44123);
assign w4190 = w4187 & w4189;
assign w4191 = (~w612 & w4029) | (~w612 & w48607) | (w4029 & w48607);
assign w4192 = ~w4029 & w48608;
assign w4193 = ~w4191 & ~w4192;
assign w4194 = ~w3703 & ~w3706;
assign w4195 = w3698 & w4194;
assign w4196 = w4193 & ~w4195;
assign w4197 = ~w4193 & w4195;
assign w4198 = ~w4196 & ~w4197;
assign w4199 = w493 & ~w4198;
assign w4200 = ~w4187 & ~w4189;
assign w4201 = (w3743 & w4029) | (w3743 & w48609) | (w4029 & w48609);
assign w4202 = w4056 & w40169;
assign w4203 = ~w4201 & ~w4202;
assign w4204 = (w612 & w4202) | (w612 & w48610) | (w4202 & w48610);
assign w4205 = (~w493 & ~w4194) | (~w493 & w51508) | (~w4194 & w51508);
assign w4206 = ~w4193 & w4205;
assign w4207 = w4194 & w51509;
assign w4208 = w4193 & w4207;
assign w4209 = ~w4206 & ~w4208;
assign w4210 = w4204 & w4209;
assign w4211 = ~w4199 & ~w4210;
assign w4212 = ~a[82] & ~a[83];
assign w4213 = ~a[84] & w4212;
assign w4214 = ~w3620 & w52175;
assign w4215 = ~a[85] & ~w4214;
assign w4216 = (w4215 & w4080) | (w4215 & w40170) | (w4080 & w40170);
assign w4217 = (~w3749 & ~w4214) | (~w3749 & w51311) | (~w4214 & w51311);
assign w4218 = (w4217 & w4039) | (w4217 & w51381) | (w4039 & w51381);
assign w4219 = ~w3993 & w4218;
assign w4220 = w4026 & w4218;
assign w4221 = ~w4041 & w4220;
assign w4222 = ~w4219 & ~w4221;
assign w4223 = w4213 & ~w3646;
assign w4224 = (~w4223 & w4080) | (~w4223 & w51510) | (w4080 & w51510);
assign w4225 = (~w3242 & ~w4224) | (~w3242 & w40171) | (~w4224 & w40171);
assign w4226 = w3242 & ~w4223;
assign w4227 = (w4226 & w4080) | (w4226 & w51382) | (w4080 & w51382);
assign w4228 = ~w4216 & w4227;
assign w4229 = ~a[86] & ~w3646;
assign w4230 = ~w3620 & w52176;
assign w4231 = a[86] & ~w3749;
assign w4232 = ~w3750 & ~w4231;
assign w4233 = ~w4229 & ~w4230;
assign w4234 = (w4233 & w4080) | (w4233 & w40172) | (w4080 & w40172);
assign w4235 = ~w4080 & w40173;
assign w4236 = ~w4234 & ~w4235;
assign w4237 = ~w4228 & ~w4236;
assign w4238 = ~w4225 & ~w4237;
assign w4239 = a[87] & ~w3753;
assign w4240 = ~w3754 & ~w4239;
assign w4241 = w4240 & ~w3646;
assign w4242 = ~w3620 & w52177;
assign w4243 = ~w4241 & ~w4242;
assign w4244 = a[87] & ~w4229;
assign w4245 = ~a[87] & w4229;
assign w4246 = ~w4244 & ~w4245;
assign w4247 = ~w4029 & w40174;
assign w4248 = (~w4246 & w4029) | (~w4246 & w40175) | (w4029 & w40175);
assign w4249 = ~w4247 & ~w4248;
assign w4250 = ~w2896 & ~w4249;
assign w4251 = ~w3769 & ~w3805;
assign w4252 = (w4251 & w4039) | (w4251 & w51314) | (w4039 & w51314);
assign w4253 = ~w3993 & w4252;
assign w4254 = w4026 & w4252;
assign w4255 = ~w4041 & w4254;
assign w4256 = ~w4253 & ~w4255;
assign w4257 = ~w4029 & ~w4256;
assign w4258 = w2558 & w3777;
assign w4259 = ~w4257 & w4258;
assign w4260 = w2558 & ~w3777;
assign w4261 = w4257 & w4260;
assign w4262 = ~w4259 & ~w4261;
assign w4263 = ~w4250 & w4262;
assign w4264 = ~w4238 & w4263;
assign w4265 = w3777 & ~w4257;
assign w4266 = ~w3777 & w4257;
assign w4267 = ~w4265 & ~w4266;
assign w4268 = ~w2558 & w4267;
assign w4269 = w2896 & w4243;
assign w4270 = ~w4080 & w40176;
assign w4271 = w2896 & w4246;
assign w4272 = (w4271 & w4080) | (w4271 & w40177) | (w4080 & w40177);
assign w4273 = ~w4270 & ~w4272;
assign w4274 = w4262 & ~w4273;
assign w4275 = ~w4268 & ~w4274;
assign w4276 = ~w3778 & w3828;
assign w4277 = (~w2807 & ~w3801) | (~w2807 & w51315) | (~w3801 & w51315);
assign w4278 = ~w4276 & ~w4277;
assign w4279 = ~w3810 & ~w4278;
assign w4280 = w2006 & w3821;
assign w4281 = (w4280 & ~w40178) | (w4280 & w51316) | (~w40178 & w51316);
assign w4282 = w2006 & ~w3821;
assign w4283 = w40178 & w51317;
assign w4284 = ~w4281 & ~w4283;
assign w4285 = ~w3778 & w51318;
assign w4286 = (w2558 & w3778) | (w2558 & w51319) | (w3778 & w51319);
assign w4287 = ~w4285 & ~w4286;
assign w4288 = w2285 & ~w3801;
assign w4289 = (w4288 & ~w40179) | (w4288 & w51320) | (~w40179 & w51320);
assign w4290 = w2285 & w3801;
assign w4291 = w40179 & w51321;
assign w4292 = ~w4289 & ~w4291;
assign w4293 = w4284 & w4292;
assign w4294 = w4275 & w4293;
assign w4295 = ~w4264 & w4294;
assign w4296 = ~w2285 & ~w3801;
assign w4297 = (w3829 & ~w40179) | (w3829 & w51322) | (~w40179 & w51322);
assign w4298 = w40179 & w51323;
assign w4299 = ~w4297 & ~w4298;
assign w4300 = ~w2006 & ~w3821;
assign w4301 = (w4300 & ~w40178) | (w4300 & w51324) | (~w40178 & w51324);
assign w4302 = ~w2006 & w3821;
assign w4303 = w40178 & w51325;
assign w4304 = ~w4301 & ~w4303;
assign w4305 = w4299 & w4304;
assign w4306 = w4284 & ~w4305;
assign w4307 = (w3841 & w51326) | (w3841 & w51327) | (w51326 & w51327);
assign w4308 = (w40181 & ~w3841) | (w40181 & w51328) | (~w3841 & w51328);
assign w4309 = ~w4307 & ~w4308;
assign w4310 = (w4080 & w51329) | (w4080 & w51330) | (w51329 & w51330);
assign w4311 = (~w3878 & ~w40182) | (~w3878 & w51331) | (~w40182 & w51331);
assign w4312 = w4310 & ~w4311;
assign w4313 = (w3880 & ~w3841) | (w3880 & w44124) | (~w3841 & w44124);
assign w4314 = ~w3895 & ~w4313;
assign w4315 = ~w4029 & w40184;
assign w4316 = ~w3992 & w51332;
assign w4317 = ~w4027 & w51333;
assign w4318 = ~w3932 & w4317;
assign w4319 = (w1541 & w4053) | (w1541 & w44125) | (w4053 & w44125);
assign w4320 = ~w4318 & ~w4319;
assign w4321 = w3852 & ~w3894;
assign w4322 = ~w1320 & ~w4321;
assign w4323 = ~w4318 & w48611;
assign w4324 = ~w4315 & w4323;
assign w4325 = ~w1320 & w4321;
assign w4326 = (w4325 & w4318) | (w4325 & w48612) | (w4318 & w48612);
assign w4327 = (w4325 & w4313) | (w4325 & w51334) | (w4313 & w51334);
assign w4328 = ~w4029 & w47093;
assign w4329 = ~w4326 & ~w4328;
assign w4330 = ~w4324 & w4329;
assign w4331 = ~w4312 & w4330;
assign w4332 = (w3821 & w4276) | (w3821 & w51335) | (w4276 & w51335);
assign w4333 = ~w3810 & ~w4332;
assign w4334 = w2006 & ~w4333;
assign w4335 = ~w2006 & w4333;
assign w4336 = ~w4334 & ~w4335;
assign w4337 = (w3836 & ~w4056) | (w3836 & w40185) | (~w4056 & w40185);
assign w4338 = w4056 & w40186;
assign w4339 = ~w4337 & ~w4338;
assign w4340 = ~w1738 & ~w4339;
assign w4341 = w4331 & ~w4340;
assign w4342 = ~w4306 & w4341;
assign w4343 = ~w4295 & w4342;
assign w4344 = ~w3897 & ~w3902;
assign w4345 = ~w3888 & ~w3898;
assign w4346 = (~w4345 & w3931) | (~w4345 & w51336) | (w3931 & w51336);
assign w4347 = ~w3932 & ~w4346;
assign w4348 = w4056 & w4347;
assign w4349 = (w4029 & w48613) | (w4029 & w48614) | (w48613 & w48614);
assign w4350 = ~w4348 & ~w4349;
assign w4351 = ~w4348 & w48615;
assign w4352 = (w945 & w4029) | (w945 & w40188) | (w4029 & w40188);
assign w4353 = (~w3905 & w3842) | (~w3905 & w44126) | (w3842 & w44126);
assign w4354 = ~w4029 & w40189;
assign w4355 = ~w3737 & ~w4188;
assign w4356 = w754 & w4355;
assign w4357 = (w4356 & w4354) | (w4356 & w51337) | (w4354 & w51337);
assign w4358 = w754 & ~w4355;
assign w4359 = ~w4354 & w51338;
assign w4360 = ~w4357 & ~w4359;
assign w4361 = ~w4351 & w4360;
assign w4362 = ~w4080 & w51339;
assign w4363 = w1541 & ~w3878;
assign w4364 = (w4363 & ~w40182) | (w4363 & w51340) | (~w40182 & w51340);
assign w4365 = ~w4362 & ~w4364;
assign w4366 = w1738 & ~w3836;
assign w4367 = (w4366 & ~w4056) | (w4366 & w40191) | (~w4056 & w40191);
assign w4368 = w1738 & w3836;
assign w4369 = w4056 & w40192;
assign w4370 = ~w4367 & ~w4369;
assign w4371 = w4365 & w4370;
assign w4372 = w4331 & ~w4371;
assign w4373 = w1320 & ~w4321;
assign w4374 = (w4373 & w4315) | (w4373 & w44127) | (w4315 & w44127);
assign w4375 = w1320 & w4321;
assign w4376 = ~w4315 & w44128;
assign w4377 = ~w4374 & ~w4376;
assign w4378 = w3865 & ~w3902;
assign w4379 = (w3841 & w51341) | (w3841 & w51342) | (w51341 & w51342);
assign w4380 = w3852 & ~w4379;
assign w4381 = (~w3901 & w4029) | (~w3901 & w40195) | (w4029 & w40195);
assign w4382 = ~w4379 & w51343;
assign w4383 = w4056 & w4382;
assign w4384 = ~w4381 & ~w4383;
assign w4385 = (w4378 & w4379) | (w4378 & w51344) | (w4379 & w51344);
assign w4386 = w4385 & w52178;
assign w4387 = w4384 & ~w4386;
assign w4388 = (~w1120 & ~w4384) | (~w1120 & w40196) | (~w4384 & w40196);
assign w4389 = w4377 & ~w4388;
assign w4390 = ~w4372 & w40197;
assign w4391 = (w4390 & w4295) | (w4390 & w51345) | (w4295 & w51345);
assign w4392 = w4384 & w40198;
assign w4393 = (w945 & w4348) | (w945 & w48616) | (w4348 & w48616);
assign w4394 = ~w4392 & ~w4393;
assign w4395 = w4361 & ~w4394;
assign w4396 = ~w4202 & w48617;
assign w4397 = ~w754 & ~w4355;
assign w4398 = (w4397 & w4354) | (w4397 & w51346) | (w4354 & w51346);
assign w4399 = ~w754 & w4355;
assign w4400 = ~w4354 & w51347;
assign w4401 = ~w4398 & ~w4400;
assign w4402 = ~w4396 & w4401;
assign w4403 = w4209 & w4402;
assign w4404 = ~w4395 & w4403;
assign w4405 = (~w40199 & w44129) | (~w40199 & w44130) | (w44129 & w44130);
assign w4406 = (~w44130 & w47094) | (~w44130 & w47095) | (w47094 & w47095);
assign w4407 = w4128 & w4136;
assign w4408 = (~w252 & w4149) | (~w252 & w51348) | (w4149 & w51348);
assign w4409 = (~w400 & w4180) | (~w400 & w48618) | (w4180 & w48618);
assign w4410 = w4174 & ~w4409;
assign w4411 = w4169 & ~w4410;
assign w4412 = ~w4408 & ~w4411;
assign w4413 = (~w57 & w4110) | (~w57 & w44131) | (w4110 & w44131);
assign w4414 = w4067 & w48619;
assign w4415 = (~w4407 & w4113) | (~w4407 & w40200) | (w4113 & w40200);
assign w4416 = w4093 & w40201;
assign w4417 = w4412 & w4416;
assign w4418 = ~w4415 & ~w4417;
assign w4419 = (w4273 & w4268) | (w4273 & w51349) | (w4268 & w51349);
assign w4420 = (w4419 & w4238) | (w4419 & w51350) | (w4238 & w51350);
assign w4421 = (~w4268 & w4264) | (~w4268 & w48620) | (w4264 & w48620);
assign w4422 = ~w4420 & ~w4421;
assign w4423 = ~w4418 & ~w4422;
assign w4424 = ~w4406 & w4423;
assign w4425 = ~w4267 & w4418;
assign w4426 = w4185 & ~w4267;
assign w4427 = ~w4405 & w4426;
assign w4428 = ~w4425 & ~w4427;
assign w4429 = ~w4424 & w4428;
assign w4430 = ~w4406 & ~w4418;
assign w4431 = ~w4184 & ~w4408;
assign w4432 = w4414 & w4431;
assign w4433 = w4141 & ~w4432;
assign w4434 = ~a[80] & ~a[81];
assign w4435 = ~a[82] & w4434;
assign w4436 = ~w4056 & ~w4435;
assign w4437 = ~w4405 & w4433;
assign w4438 = (~w4436 & w4437) | (~w4436 & w47096) | (w4437 & w47096);
assign w4439 = a[83] & w52179;
assign w4440 = ~w4430 & w4439;
assign w4441 = w4438 & ~w4440;
assign w4442 = w4056 & w4435;
assign w4443 = w4211 & w4412;
assign w4444 = ~w4431 & ~w4443;
assign w4445 = w4404 & ~w4431;
assign w4446 = ~w4391 & w4445;
assign w4447 = a[82] & ~a[83];
assign w4448 = (w4447 & ~w4128) | (w4447 & w51351) | (~w4128 & w51351);
assign w4449 = (w4141 & w4446) | (w4141 & w47097) | (w4446 & w47097);
assign w4450 = (~w4442 & w4449) | (~w4442 & w48621) | (w4449 & w48621);
assign w4451 = ~w4441 & w4450;
assign w4452 = (~w4114 & ~w4113) | (~w4114 & w40203) | (~w4113 & w40203);
assign w4453 = w4412 & w4414;
assign w4454 = w4452 & ~w4453;
assign w4455 = ~a[84] & w4056;
assign w4456 = a[84] & ~w4056;
assign w4457 = ~w4455 & ~w4456;
assign w4458 = w4457 & w52179;
assign w4459 = ~w4128 & ~w4454;
assign w4460 = w4405 & w4459;
assign w4461 = w4458 & ~w4460;
assign w4462 = a[84] & ~w4212;
assign w4463 = ~w4213 & ~w4462;
assign w4464 = ~w4418 & w4463;
assign w4465 = ~w4406 & w4464;
assign w4466 = (~w3646 & w4461) | (~w3646 & w48622) | (w4461 & w48622);
assign w4467 = w4451 & ~w4466;
assign w4468 = ~w4461 & w44133;
assign w4469 = ~w4214 & ~w4223;
assign w4470 = a[85] & ~w4056;
assign w4471 = ~w4080 & w51352;
assign w4472 = ~w4470 & ~w4471;
assign w4473 = w4469 & ~w4472;
assign w4474 = ~w4469 & w4472;
assign w4475 = ~w4473 & ~w4474;
assign w4476 = (a[85] & ~w4056) | (a[85] & w51353) | (~w4056 & w51353);
assign w4477 = w4056 & w3749;
assign w4478 = ~w4476 & ~w4477;
assign w4479 = w3242 & w4475;
assign w4480 = ~w4406 & w48623;
assign w4481 = w3242 & ~w4478;
assign w4482 = (w4481 & w4406) | (w4481 & w48624) | (w4406 & w48624);
assign w4483 = ~w4480 & ~w4482;
assign w4484 = ~w4468 & w4483;
assign w4485 = ~w4467 & w4484;
assign w4486 = ~w4225 & ~w4228;
assign w4487 = ~w4418 & w4486;
assign w4488 = ~w4406 & w4487;
assign w4489 = w4236 & ~w4488;
assign w4490 = ~w4236 & w4488;
assign w4491 = ~w4489 & ~w4490;
assign w4492 = w2896 & w4491;
assign w4493 = ~w4406 & w48625;
assign w4494 = (~w4478 & w4406) | (~w4478 & w48626) | (w4406 & w48626);
assign w4495 = ~w4493 & ~w4494;
assign w4496 = ~w3242 & w4495;
assign w4497 = ~w4492 & ~w4496;
assign w4498 = ~w4485 & w4497;
assign w4499 = ~w2896 & w4236;
assign w4500 = ~w4488 & w4499;
assign w4501 = ~w2896 & ~w4236;
assign w4502 = w4488 & w4501;
assign w4503 = ~w4500 & ~w4502;
assign w4504 = (w2896 & w4237) | (w2896 & w51354) | (w4237 & w51354);
assign w4505 = ~w4237 & w51355;
assign w4506 = ~w4504 & ~w4505;
assign w4507 = ~w4418 & w4506;
assign w4508 = ~w4406 & w4507;
assign w4509 = ~w4080 & w51356;
assign w4510 = (~w4246 & w4080) | (~w4246 & w51357) | (w4080 & w51357);
assign w4511 = ~w4509 & ~w4510;
assign w4512 = w2558 & ~w4249;
assign w4513 = ~w4508 & w4512;
assign w4514 = w2558 & w4511;
assign w4515 = w4508 & w4514;
assign w4516 = ~w4513 & ~w4515;
assign w4517 = w4503 & w4516;
assign w4518 = (~w2285 & ~w4428) | (~w2285 & w47098) | (~w4428 & w47098);
assign w4519 = w4292 & w4299;
assign w4520 = ~w4264 & w48627;
assign w4521 = (w4519 & w4264) | (w4519 & w48628) | (w4264 & w48628);
assign w4522 = ~w4520 & ~w4521;
assign w4523 = (w3801 & ~w40179) | (w3801 & w51358) | (~w40179 & w51358);
assign w4524 = w40179 & w51359;
assign w4525 = ~w4523 & ~w4524;
assign w4526 = w4185 & w4525;
assign w4527 = ~w4405 & w4526;
assign w4528 = w4418 & w4525;
assign w4529 = ~w4527 & ~w4528;
assign w4530 = ~w4418 & w4522;
assign w4531 = ~w4406 & w4530;
assign w4532 = w4529 & ~w4531;
assign w4533 = (w2006 & ~w4529) | (w2006 & w47099) | (~w4529 & w47099);
assign w4534 = w4518 & ~w4533;
assign w4535 = w4517 & ~w4534;
assign w4536 = (w4535 & w4485) | (w4535 & w48629) | (w4485 & w48629);
assign w4537 = (~w4264 & w51360) | (~w4264 & w51361) | (w51360 & w51361);
assign w4538 = (w40204 & w4264) | (w40204 & w51362) | (w4264 & w51362);
assign w4539 = (~w4264 & w51363) | (~w4264 & w51364) | (w51363 & w51364);
assign w4540 = ~w4537 & ~w4539;
assign w4541 = w4330 & w4377;
assign w4542 = ~w4312 & ~w4541;
assign w4543 = w4540 & w4542;
assign w4544 = ~w4365 & ~w4541;
assign w4545 = ~w4544 & w52180;
assign w4546 = (w4321 & w4315) | (w4321 & w51365) | (w4315 & w51365);
assign w4547 = ~w4315 & w51366;
assign w4548 = ~w4546 & ~w4547;
assign w4549 = (~w4548 & w4406) | (~w4548 & w48631) | (w4406 & w48631);
assign w4550 = ~w4543 & w4545;
assign w4551 = w4430 & w4550;
assign w4552 = ~w4549 & ~w4551;
assign w4553 = ~w1541 & w4185;
assign w4554 = ~w4405 & w4553;
assign w4555 = ~w1541 & w4418;
assign w4556 = ~w4554 & ~w4555;
assign w4557 = ~w4418 & ~w4540;
assign w4558 = ~w4406 & w4557;
assign w4559 = ~w4312 & w4365;
assign w4560 = w1320 & w4559;
assign w4561 = (w4560 & ~w4556) | (w4560 & w48632) | (~w4556 & w48632);
assign w4562 = w1320 & ~w4559;
assign w4563 = w4556 & w48633;
assign w4564 = ~w4561 & ~w4563;
assign w4565 = ~w4551 & w51367;
assign w4566 = w4564 & ~w4565;
assign w4567 = ~w4537 & ~w4538;
assign w4568 = ~w4418 & w4567;
assign w4569 = ~w4406 & w4568;
assign w4570 = w1541 & w4339;
assign w4571 = ~w4569 & w4570;
assign w4572 = w1541 & ~w4339;
assign w4573 = w4569 & w4572;
assign w4574 = ~w4571 & ~w4573;
assign w4575 = w4284 & w4304;
assign w4576 = (w4292 & w48634) | (w4292 & w4295) | (w48634 & w4295);
assign w4577 = (~w4575 & w48635) | (~w4575 & w52181) | (w48635 & w52181);
assign w4578 = ~w4418 & ~w4577;
assign w4579 = w4575 & ~w4576;
assign w4580 = w4578 & ~w4579;
assign w4581 = (w3821 & ~w40178) | (w3821 & w51368) | (~w40178 & w51368);
assign w4582 = w40178 & w51369;
assign w4583 = ~w4581 & ~w4582;
assign w4584 = w4185 & ~w4583;
assign w4585 = ~w4405 & w4584;
assign w4586 = w4418 & ~w4583;
assign w4587 = ~w4585 & ~w4586;
assign w4588 = ~w4406 & w4580;
assign w4589 = w4587 & ~w4588;
assign w4590 = (w1738 & w4588) | (w1738 & w44134) | (w4588 & w44134);
assign w4591 = w4574 & ~w4590;
assign w4592 = (w2285 & ~w4418) | (w2285 & w44135) | (~w4418 & w44135);
assign w4593 = ~w4427 & w4592;
assign w4594 = ~w4424 & w4593;
assign w4595 = ~w2558 & ~w4511;
assign w4596 = ~w4418 & w44136;
assign w4597 = ~w2558 & w4249;
assign w4598 = (~w4597 & w4418) | (~w4597 & w44137) | (w4418 & w44137);
assign w4599 = w4185 & ~w4597;
assign w4600 = ~w4405 & w4599;
assign w4601 = ~w4598 & ~w4600;
assign w4602 = ~w4406 & w4596;
assign w4603 = w4601 & ~w4602;
assign w4604 = ~w4594 & ~w4603;
assign w4605 = ~w4518 & ~w4604;
assign w4606 = (~w4533 & w4604) | (~w4533 & w4534) | (w4604 & w4534);
assign w4607 = w4591 & w4606;
assign w4608 = w4566 & w4607;
assign w4609 = ~w4536 & w4608;
assign w4610 = ~w4588 & w44138;
assign w4611 = w4529 & w47102;
assign w4612 = ~w4610 & ~w4611;
assign w4613 = w4591 & ~w4612;
assign w4614 = (~w1541 & w4569) | (~w1541 & w48636) | (w4569 & w48636);
assign w4615 = ~w4339 & w4569;
assign w4616 = w4614 & ~w4615;
assign w4617 = ~w1320 & ~w4559;
assign w4618 = (w4617 & ~w4556) | (w4617 & w47103) | (~w4556 & w47103);
assign w4619 = ~w1320 & w4559;
assign w4620 = w4556 & w47104;
assign w4621 = ~w4618 & ~w4620;
assign w4622 = ~w4616 & w4621;
assign w4623 = ~w4613 & w4622;
assign w4624 = w4566 & ~w4623;
assign w4625 = (~w4351 & w4392) | (~w4351 & w51511) | (w4392 & w51511);
assign w4626 = ~w4372 & w40206;
assign w4627 = w4360 & w4401;
assign w4628 = (w4343 & w49480) | (w4343 & w49481) | (w49480 & w49481);
assign w4629 = (~w4343 & w49482) | (~w4343 & w49483) | (w49482 & w49483);
assign w4630 = ~w4628 & ~w4629;
assign w4631 = ~w4354 & w51370;
assign w4632 = (w4355 & w4354) | (w4355 & w51371) | (w4354 & w51371);
assign w4633 = ~w4631 & ~w4632;
assign w4634 = w4430 & w4630;
assign w4635 = (w4633 & w4406) | (w4633 & w48637) | (w4406 & w48637);
assign w4636 = ~w4634 & ~w4635;
assign w4637 = ~w4634 & w48638;
assign w4638 = ~w4395 & w4401;
assign w4639 = (w4343 & w51372) | (w4343 & w51373) | (w51372 & w51373);
assign w4640 = ~w612 & w4360;
assign w4641 = (~w4343 & w51374) | (~w4343 & w51375) | (w51374 & w51375);
assign w4642 = ~w4639 & ~w4641;
assign w4643 = w4430 & w4642;
assign w4644 = w493 & ~w4203;
assign w4645 = ~w4643 & w4644;
assign w4646 = w493 & w4203;
assign w4647 = w4643 & w4646;
assign w4648 = ~w4645 & ~w4647;
assign w4649 = ~w4637 & w4648;
assign w4650 = (w4343 & w51376) | (w4343 & w51377) | (w51376 & w51377);
assign w4651 = ~w4351 & ~w4393;
assign w4652 = w4392 & ~w4651;
assign w4653 = ~w4372 & w40208;
assign w4654 = (~w4652 & w4343) | (~w4652 & w40209) | (w4343 & w40209);
assign w4655 = ~w4418 & w4654;
assign w4656 = ~w4650 & w4655;
assign w4657 = ~w4406 & w4656;
assign w4658 = w4185 & w4350;
assign w4659 = ~w4405 & w4658;
assign w4660 = w4350 & w4418;
assign w4661 = ~w4659 & ~w4660;
assign w4662 = ~w4657 & w4661;
assign w4663 = ~w4657 & w44139;
assign w4664 = ~w612 & w4630;
assign w4665 = w4430 & w4664;
assign w4666 = ~w612 & w4633;
assign w4667 = (w4666 & w4406) | (w4666 & w51512) | (w4406 & w51512);
assign w4668 = ~w4665 & ~w4667;
assign w4669 = ~w4663 & w4668;
assign w4670 = (w754 & w4657) | (w754 & w44140) | (w4657 & w44140);
assign w4671 = (w40210 & w4295) | (w40210 & w48639) | (w4295 & w48639);
assign w4672 = w4185 & w4387;
assign w4673 = ~w4405 & w4672;
assign w4674 = w4387 & w4418;
assign w4675 = ~w4673 & ~w4674;
assign w4676 = ~w4418 & w44141;
assign w4677 = ~w4406 & w4676;
assign w4678 = w4675 & ~w4677;
assign w4679 = (w1120 & w40211) | (w1120 & w4343) | (w40211 & w4343);
assign w4680 = ~w4418 & w44142;
assign w4681 = ~w4406 & w4680;
assign w4682 = ~w4671 & ~w4679;
assign w4683 = w4387 & w4682;
assign w4684 = ~w4681 & ~w4683;
assign w4685 = w4678 & w4684;
assign w4686 = (w945 & ~w4678) | (w945 & w47106) | (~w4678 & w47106);
assign w4687 = ~w4670 & w4686;
assign w4688 = w4669 & ~w4687;
assign w4689 = (~w4182 & w4418) | (~w4182 & w51513) | (w4418 & w51513);
assign w4690 = w400 & ~w4185;
assign w4691 = ~w4418 & w4690;
assign w4692 = ~w4181 & ~w4691;
assign w4693 = ~w4182 & ~w4211;
assign w4694 = ~w4182 & w4404;
assign w4695 = ~w4391 & w4694;
assign w4696 = w400 & w4185;
assign w4697 = ~w4695 & ~w4696;
assign w4698 = ~w4418 & ~w4693;
assign w4699 = w4697 & w4698;
assign w4700 = ~w4692 & ~w4699;
assign w4701 = w4405 & ~w4689;
assign w4702 = (~w4701 & w4699) | (~w4701 & w51514) | (w4699 & w51514);
assign w4703 = ~w4700 & w47107;
assign w4704 = ~w4199 & w4209;
assign w4705 = (~w4204 & w40212) | (~w4204 & w52182) | (w40212 & w52182);
assign w4706 = w4704 & ~w4705;
assign w4707 = ~w4704 & w4705;
assign w4708 = ~w4706 & ~w4707;
assign w4709 = (~w4198 & w4406) | (~w4198 & w48640) | (w4406 & w48640);
assign w4710 = w4430 & w4708;
assign w4711 = ~w4710 & w48641;
assign w4712 = (~w351 & w4700) | (~w351 & w47108) | (w4700 & w47108);
assign w4713 = ~w351 & w4168;
assign w4714 = w4174 & ~w4713;
assign w4715 = w4168 & w4174;
assign w4716 = (~w4715 & w40213) | (~w4715 & w4695) | (w40213 & w4695);
assign w4717 = ~w4409 & w4715;
assign w4718 = (w4717 & w4211) | (w4717 & w51383) | (w4211 & w51383);
assign w4719 = (w4718 & w4391) | (w4718 & w48642) | (w4391 & w48642);
assign w4720 = ~w4716 & ~w4719;
assign w4721 = w4430 & w4720;
assign w4722 = (w252 & w4721) | (w252 & w47109) | (w4721 & w47109);
assign w4723 = ~w4712 & ~w4722;
assign w4724 = (w1120 & w4551) | (w1120 & w48643) | (w4551 & w48643);
assign w4725 = ~w493 & w4203;
assign w4726 = ~w4643 & w4725;
assign w4727 = ~w493 & ~w4203;
assign w4728 = w4643 & w4727;
assign w4729 = ~w4726 & ~w4728;
assign w4730 = ~w4724 & w4729;
assign w4731 = w4723 & w4730;
assign w4732 = ~w4703 & w4711;
assign w4733 = w4731 & ~w4732;
assign w4734 = w4649 & ~w4688;
assign w4735 = w4733 & ~w4734;
assign w4736 = ~w4624 & w4735;
assign w4737 = ~w4609 & w4736;
assign w4738 = (~w400 & w4710) | (~w400 & w48644) | (w4710 & w48644);
assign w4739 = ~w4703 & ~w4738;
assign w4740 = (~w945 & ~w4682) | (~w945 & w47110) | (~w4682 & w47110);
assign w4741 = ~w4681 & w4740;
assign w4742 = w4678 & w4741;
assign w4743 = ~w4670 & ~w4742;
assign w4744 = w4669 & ~w4743;
assign w4745 = w4649 & ~w4744;
assign w4746 = ~w4744 & w47111;
assign w4747 = ~w4711 & w4729;
assign w4748 = w4739 & ~w4747;
assign w4749 = w4723 & ~w4748;
assign w4750 = ~w4746 & w4749;
assign w4751 = w4067 & w4102;
assign w4752 = ~w4413 & w4751;
assign w4753 = (w4102 & ~w4751) | (w4102 & w51515) | (~w4751 & w51515);
assign w4754 = ~w4753 & w52183;
assign w4755 = ~w4113 & ~w4114;
assign w4756 = ~w4113 & w51516;
assign w4757 = ~w4113 & w47112;
assign w4758 = (w42 & w4113) | (w42 & w47113) | (w4113 & w47113);
assign w4759 = ~w4757 & ~w4758;
assign w4760 = w40215 & w44143;
assign w4761 = (w4759 & ~w40215) | (w4759 & w44144) | (~w40215 & w44144);
assign w4762 = ~w4760 & ~w4761;
assign w4763 = (w4136 & w4091) | (w4136 & w51517) | (w4091 & w51517);
assign w4764 = (w4755 & w4446) | (w4755 & w48645) | (w4446 & w48645);
assign w4765 = w163 & w4091;
assign w4766 = (w4127 & w4754) | (w4127 & w48646) | (w4754 & w48646);
assign w4767 = ~w42 & ~w4764;
assign w4768 = w4766 & ~w4767;
assign w4769 = ~w4127 & ~w4763;
assign w4770 = (w4769 & ~w4762) | (w4769 & w47114) | (~w4762 & w47114);
assign w4771 = ~w4768 & ~w4770;
assign w4772 = ~w4092 & ~w4114;
assign w4773 = (~w4091 & w4406) | (~w4091 & w51518) | (w4406 & w51518);
assign w4774 = w4430 & ~w4754;
assign w4775 = (~w4773 & ~w4774) | (~w4773 & w51519) | (~w4774 & w51519);
assign w4776 = w4430 & w4754;
assign w4777 = ~w4772 & w4776;
assign w4778 = (~w4446 & w47115) | (~w4446 & w47116) | (w47115 & w47116);
assign w4779 = w4430 & ~w4778;
assign w4780 = ~w4111 & ~w4751;
assign w4781 = (w4780 & w4446) | (w4780 & w51520) | (w4446 & w51520);
assign w4782 = ~w4047 & ~w4057;
assign w4783 = w4058 & ~w4782;
assign w4784 = ~w4058 & w4782;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = (~w4785 & w4406) | (~w4785 & w51521) | (w4406 & w51521);
assign w4787 = ~w3 & ~w4786;
assign w4788 = w4779 & ~w4781;
assign w4789 = w4787 & ~w4788;
assign w4790 = (~w42 & ~w4776) | (~w42 & w48647) | (~w4776 & w48647);
assign w4791 = w4775 & w4790;
assign w4792 = ~w4789 & ~w4791;
assign w4793 = w4771 & ~w4792;
assign w4794 = ~w4151 & ~w4408;
assign w4795 = (w4168 & w4695) | (w4168 & w40217) | (w4695 & w40217);
assign w4796 = (~w4695 & w47117) | (~w4695 & w47118) | (w47117 & w47118);
assign w4797 = (w4695 & w47119) | (w4695 & w47120) | (w47119 & w47120);
assign w4798 = ~w4796 & ~w4797;
assign w4799 = (w4150 & w4406) | (w4150 & w48648) | (w4406 & w48648);
assign w4800 = ~w57 & ~w4799;
assign w4801 = w4430 & w4798;
assign w4802 = w4800 & ~w4801;
assign w4803 = ~w57 & w4185;
assign w4804 = ~w4405 & w4803;
assign w4805 = (~w4418 & w4446) | (~w4418 & w40218) | (w4446 & w40218);
assign w4806 = ~w4406 & w4805;
assign w4807 = ~w4111 & ~w4413;
assign w4808 = w80 & ~w4807;
assign w4809 = (w4808 & w4806) | (w4808 & w44145) | (w4806 & w44145);
assign w4810 = w80 & w4807;
assign w4811 = ~w4806 & w44146;
assign w4812 = ~w4809 & ~w4811;
assign w4813 = ~w4802 & w4812;
assign w4814 = ~w4721 & w47121;
assign w4815 = (~w4150 & w4406) | (~w4150 & w40219) | (w4406 & w40219);
assign w4816 = w57 & ~w4815;
assign w4817 = w4430 & ~w4798;
assign w4818 = w4816 & ~w4817;
assign w4819 = w4814 & ~w4818;
assign w4820 = w4813 & ~w4819;
assign w4821 = (w40220 & w4406) | (w40220 & w51522) | (w4406 & w51522);
assign w4822 = (w3 & w40221) | (w3 & w52184) | (w40221 & w52184);
assign w4823 = (~w4821 & ~w4779) | (~w4821 & w51523) | (~w4779 & w51523);
assign w4824 = ~w80 & ~w4807;
assign w4825 = ~w4806 & w44147;
assign w4826 = ~w80 & w4807;
assign w4827 = (w4826 & w4806) | (w4826 & w44148) | (w4806 & w44148);
assign w4828 = ~w4825 & ~w4827;
assign w4829 = w4823 & w4828;
assign w4830 = w4771 & w4829;
assign w4831 = ~w4820 & w4830;
assign w4832 = ~w4793 & ~w4831;
assign w4833 = ~w4750 & w4832;
assign w4834 = w4812 & w4818;
assign w4835 = w4829 & ~w4834;
assign w4836 = w4771 & w4835;
assign w4837 = ~w4793 & ~w4836;
assign w4838 = (~w4837 & w4737) | (~w4837 & w4968) | (w4737 & w4968);
assign w4839 = ~w4518 & ~w4594;
assign w4840 = ~w4497 & w4517;
assign w4841 = w4484 & w4517;
assign w4842 = ~w4467 & w4841;
assign w4843 = ~w4840 & ~w4842;
assign w4844 = (w4839 & ~w4843) | (w4839 & w51524) | (~w4843 & w51524);
assign w4845 = w4843 & w51525;
assign w4846 = ~w4844 & ~w4845;
assign w4847 = w4429 & w4838;
assign w4848 = ~w4838 & w4846;
assign w4849 = ~w4847 & ~w4848;
assign w4850 = ~w4606 & ~w4611;
assign w4851 = ~w4518 & ~w4611;
assign w4852 = (w4843 & w44149) | (w4843 & w44150) | (w44149 & w44150);
assign w4853 = ~w4610 & ~w4852;
assign w4854 = w1541 & w4838;
assign w4855 = ~w4838 & w4853;
assign w4856 = ~w4854 & ~w4855;
assign w4857 = w4574 & ~w4616;
assign w4858 = ~w1320 & ~w4857;
assign w4859 = w4856 & w4858;
assign w4860 = ~w4590 & ~w4610;
assign w4861 = (w4843 & w44151) | (w4843 & w44152) | (w44151 & w44152);
assign w4862 = w4860 & w52185;
assign w4863 = ~w4861 & ~w4862;
assign w4864 = ~w1541 & w4589;
assign w4865 = w4838 & w4864;
assign w4866 = ~w1541 & ~w4863;
assign w4867 = ~w4838 & w4866;
assign w4868 = ~w4865 & ~w4867;
assign w4869 = ~w1320 & w4857;
assign w4870 = w4857 & w51526;
assign w4871 = w4838 & w4870;
assign w4872 = ~w4852 & w51527;
assign w4873 = ~w4838 & w4872;
assign w4874 = ~w4871 & ~w4873;
assign w4875 = w4868 & w4874;
assign w4876 = ~w4859 & w4875;
assign w4877 = ~w2006 & w4849;
assign w4878 = (~w4518 & ~w4843) | (~w4518 & w4605) | (~w4843 & w4605);
assign w4879 = w2006 & w4838;
assign w4880 = ~w4838 & w4878;
assign w4881 = ~w4879 & ~w4880;
assign w4882 = ~w4533 & ~w4611;
assign w4883 = ~w1738 & ~w4882;
assign w4884 = w4881 & w4883;
assign w4885 = ~w1738 & w4882;
assign w4886 = ~w4881 & w4885;
assign w4887 = ~w4884 & ~w4886;
assign w4888 = ~w4877 & w4887;
assign w4889 = w4876 & w4888;
assign w4890 = w2006 & ~w4849;
assign w4891 = (~w2558 & w4836) | (~w2558 & w51528) | (w4836 & w51528);
assign w4892 = (w4891 & w4737) | (w4891 & w40223) | (w4737 & w40223);
assign w4893 = (w4503 & w4485) | (w4503 & w51529) | (w4485 & w51529);
assign w4894 = w4833 & w4893;
assign w4895 = ~w4737 & w4894;
assign w4896 = w4837 & w4893;
assign w4897 = ~w4895 & ~w4896;
assign w4898 = w4516 & ~w4603;
assign w4899 = w2285 & ~w4898;
assign w4900 = (w4899 & ~w4897) | (w4899 & w40224) | (~w4897 & w40224);
assign w4901 = w2285 & w4898;
assign w4902 = w4897 & w40225;
assign w4903 = ~w4900 & ~w4902;
assign w4904 = ~w4890 & w4903;
assign w4905 = ~w4492 & w4503;
assign w4906 = (~w4496 & w4467) | (~w4496 & w51530) | (w4467 & w51530);
assign w4907 = w4905 & ~w4906;
assign w4908 = ~w4905 & w4906;
assign w4909 = ~w4907 & ~w4908;
assign w4910 = ~w2558 & w4909;
assign w4911 = ~w4838 & w4910;
assign w4912 = w4491 & w4892;
assign w4913 = ~w4911 & ~w4912;
assign w4914 = (~w4468 & ~w4451) | (~w4468 & w51531) | (~w4451 & w51531);
assign w4915 = ~w3242 & w4914;
assign w4916 = w3242 & ~w4914;
assign w4917 = ~w4915 & ~w4916;
assign w4918 = w4833 & w4917;
assign w4919 = ~w4737 & w4918;
assign w4920 = w4837 & w4917;
assign w4921 = w2896 & ~w4495;
assign w4922 = (w4921 & w4919) | (w4921 & w40226) | (w4919 & w40226);
assign w4923 = w2896 & w4495;
assign w4924 = ~w4919 & w40227;
assign w4925 = ~w4922 & ~w4924;
assign w4926 = w4913 & w4925;
assign w4927 = ~w2896 & w4495;
assign w4928 = (w4927 & w4919) | (w4927 & w40228) | (w4919 & w40228);
assign w4929 = ~w2896 & ~w4495;
assign w4930 = ~w4919 & w40229;
assign w4931 = ~w4928 & ~w4930;
assign w4932 = ~w4441 & w51532;
assign w4933 = (w3646 & w4441) | (w3646 & w51533) | (w4441 & w51533);
assign w4934 = ~w4932 & ~w4933;
assign w4935 = ~w4836 & w51534;
assign w4936 = w4833 & ~w4934;
assign w4937 = ~w4737 & w4936;
assign w4938 = (w3242 & w4461) | (w3242 & w51535) | (w4461 & w51535);
assign w4939 = (w4938 & w4937) | (w4938 & w40230) | (w4937 & w40230);
assign w4940 = ~w4461 & w51536;
assign w4941 = ~w4937 & w40231;
assign w4942 = ~w4939 & ~w4941;
assign w4943 = w4931 & w4942;
assign w4944 = w4926 & ~w4943;
assign w4945 = w4491 & w4838;
assign w4946 = ~w4838 & w4909;
assign w4947 = ~w4945 & ~w4946;
assign w4948 = w2558 & w4947;
assign w4949 = ~w2285 & ~w4898;
assign w4950 = w4897 & w40232;
assign w4951 = ~w2285 & w4898;
assign w4952 = (w4951 & ~w4897) | (w4951 & w40233) | (~w4897 & w40233);
assign w4953 = ~w4950 & ~w4952;
assign w4954 = ~w4948 & w4953;
assign w4955 = ~w4944 & w4954;
assign w4956 = ~w4406 & w51537;
assign w4957 = (w4956 & w4836) | (w4956 & w51548) | (w4836 & w51548);
assign w4958 = ~a[83] & ~w4957;
assign w4959 = ~a[83] & w4833;
assign w4960 = ~w4737 & w4959;
assign w4961 = ~w4958 & ~w4960;
assign w4962 = w4608 & w4843;
assign w4963 = w4735 & ~w4962;
assign w4964 = w4534 & w4591;
assign w4965 = w4564 & ~w4964;
assign w4966 = w4623 & w4965;
assign w4967 = w4566 & ~w4966;
assign w4968 = ~w4833 & ~w4837;
assign w4969 = ~w4837 & ~w4967;
assign w4970 = w4963 & w4969;
assign w4971 = ~w4968 & ~w4970;
assign w4972 = ~w4436 & ~w4442;
assign w4973 = ~w4406 & w51549;
assign w4974 = (w4972 & w4406) | (w4972 & w51550) | (w4406 & w51550);
assign w4975 = ~w4973 & ~w4974;
assign w4976 = w4971 & ~w4975;
assign w4977 = ~w4961 & ~w4976;
assign w4978 = (w40234 & w4836) | (w40234 & w51551) | (w4836 & w51551);
assign w4979 = a[83] & ~w4975;
assign w4980 = w4833 & w4979;
assign w4981 = ~w4737 & w4980;
assign w4982 = ~w4836 & w51552;
assign w4983 = ~w4981 & ~w4982;
assign w4984 = (w4978 & w4737) | (w4978 & w44153) | (w4737 & w44153);
assign w4985 = w4983 & ~w4984;
assign w4986 = ~w4977 & w4985;
assign w4987 = ~w3646 & ~w4986;
assign w4988 = ~a[78] & ~a[79];
assign w4989 = ~a[80] & w4988;
assign w4990 = ~w4406 & w51553;
assign w4991 = (~w4990 & w4836) | (~w4990 & w51554) | (w4836 & w51554);
assign w4992 = (w4991 & w4737) | (w4991 & w40235) | (w4737 & w40235);
assign w4993 = (~w4989 & w4406) | (~w4989 & w51555) | (w4406 & w51555);
assign w4994 = ~a[81] & ~w4990;
assign w4995 = ~w4993 & ~w4994;
assign w4996 = w4434 & w4971;
assign w4997 = (w4993 & w4836) | (w4993 & w51556) | (w4836 & w51556);
assign w4998 = ~a[81] & ~w4997;
assign w4999 = ~a[81] & w4833;
assign w5000 = ~w4737 & w4999;
assign w5001 = ~w4998 & ~w5000;
assign w5002 = ~w4992 & w4995;
assign w5003 = ~w4996 & ~w5001;
assign w5004 = ~w5002 & ~w5003;
assign w5005 = ~a[82] & w4056;
assign w5006 = (w4430 & w4836) | (w4430 & w51557) | (w4836 & w51557);
assign w5007 = w4833 & w5005;
assign w5008 = ~w4737 & w5007;
assign w5009 = w5005 & ~w5006;
assign w5010 = ~w5008 & ~w5009;
assign w5011 = a[82] & w4056;
assign w5012 = w5006 & w5011;
assign w5013 = (w5012 & w4737) | (w5012 & w51558) | (w4737 & w51558);
assign w5014 = w4056 & w51559;
assign w5015 = w4971 & w5014;
assign w5016 = ~w5013 & ~w5015;
assign w5017 = ~w4996 & ~w5010;
assign w5018 = w5016 & ~w5017;
assign w5019 = w5004 & w5018;
assign w5020 = a[82] & ~w4056;
assign w5021 = ~w5006 & w5020;
assign w5022 = w4833 & w5020;
assign w5023 = ~w4737 & w5022;
assign w5024 = ~w5021 & ~w5023;
assign w5025 = ~w4056 & w4957;
assign w5026 = (w5025 & w4737) | (w5025 & w51560) | (w4737 & w51560);
assign w5027 = ~w4056 & w4435;
assign w5028 = w4971 & w5027;
assign w5029 = ~w5026 & ~w5028;
assign w5030 = ~w4996 & ~w5024;
assign w5031 = w5029 & ~w5030;
assign w5032 = w3646 & ~w4978;
assign w5033 = w3646 & w4833;
assign w5034 = ~w4737 & w5033;
assign w5035 = ~w5032 & ~w5034;
assign w5036 = w4983 & ~w5035;
assign w5037 = ~w4977 & w5036;
assign w5038 = w5031 & ~w5037;
assign w5039 = ~w5019 & w5038;
assign w5040 = ~w4987 & ~w5039;
assign w5041 = ~w4461 & w51561;
assign w5042 = (w5041 & w4937) | (w5041 & w40236) | (w4937 & w40236);
assign w5043 = (~w3242 & w4461) | (~w3242 & w51562) | (w4461 & w51562);
assign w5044 = ~w4937 & w40237;
assign w5045 = ~w5042 & ~w5044;
assign w5046 = w4931 & ~w5045;
assign w5047 = w4926 & ~w5046;
assign w5048 = w4904 & ~w4955;
assign w5049 = w4904 & w5047;
assign w5050 = w5040 & w5049;
assign w5051 = ~w5050 & w40238;
assign w5052 = ~w4663 & ~w4670;
assign w5053 = ~w4686 & ~w4724;
assign w5054 = (w5053 & w4623) | (w5053 & w40239) | (w4623 & w40239);
assign w5055 = w4607 & w40240;
assign w5056 = ~w4536 & w5055;
assign w5057 = (~w5052 & w5056) | (~w5052 & w40241) | (w5056 & w40241);
assign w5058 = ~w5056 & w40242;
assign w5059 = ~w5057 & ~w5058;
assign w5060 = ~w4838 & w5059;
assign w5061 = (~w4662 & w4836) | (~w4662 & w51563) | (w4836 & w51563);
assign w5062 = (w5061 & w4737) | (w5061 & w40243) | (w4737 & w40243);
assign w5063 = ~w612 & ~w5062;
assign w5064 = ~w5060 & w5063;
assign w5065 = (~w4685 & w4836) | (~w4685 & w51564) | (w4836 & w51564);
assign w5066 = (w5065 & w4737) | (w5065 & w40244) | (w4737 & w40244);
assign w5067 = ~w4686 & ~w4742;
assign w5068 = ~w5067 & w50183;
assign w5069 = w4607 & w40246;
assign w5070 = ~w4536 & w5069;
assign w5071 = ~w5068 & ~w5070;
assign w5072 = w5067 & ~w50183;
assign w5073 = ~w4609 & w5072;
assign w5074 = w5071 & ~w5073;
assign w5075 = ~w754 & w5066;
assign w5076 = ~w754 & ~w5074;
assign w5077 = ~w4838 & w5076;
assign w5078 = ~w5075 & ~w5077;
assign w5079 = ~w5064 & w5078;
assign w5080 = ~w4838 & ~w5074;
assign w5081 = w754 & ~w5066;
assign w5082 = ~w5080 & w5081;
assign w5083 = w4607 & w4966;
assign w5084 = ~w4536 & w5083;
assign w5085 = ~w1120 & ~w4564;
assign w5086 = w1120 & w4564;
assign w5087 = ~w5085 & ~w5086;
assign w5088 = ~w1120 & w4966;
assign w5089 = ~w4966 & ~w5087;
assign w5090 = ~w5088 & ~w5089;
assign w5091 = w5084 & ~w5090;
assign w5092 = ~w5084 & w5090;
assign w5093 = ~w5091 & ~w5092;
assign w5094 = (~w945 & w4551) | (~w945 & w51565) | (w4551 & w51565);
assign w5095 = ~w5093 & w5094;
assign w5096 = ~w4838 & w5095;
assign w5097 = ~w4551 & w51566;
assign w5098 = (w5097 & w4836) | (w5097 & w51567) | (w4836 & w51567);
assign w5099 = (w5098 & w4737) | (w5098 & w40247) | (w4737 & w40247);
assign w5100 = w5093 & w5097;
assign w5101 = ~w5099 & ~w5100;
assign w5102 = ~w5096 & w5101;
assign w5103 = ~w5082 & w5102;
assign w5104 = ~w4551 & w51568;
assign w5105 = ~w5093 & w5104;
assign w5106 = ~w4838 & w5105;
assign w5107 = (w945 & w4551) | (w945 & w51569) | (w4551 & w51569);
assign w5108 = (w5107 & w4836) | (w5107 & w51570) | (w4836 & w51570);
assign w5109 = (w5108 & w4737) | (w5108 & w40248) | (w4737 & w40248);
assign w5110 = w5093 & w5107;
assign w5111 = ~w5109 & ~w5110;
assign w5112 = ~w5106 & w5111;
assign w5113 = w4556 & w51571;
assign w5114 = (w4559 & ~w4556) | (w4559 & w51572) | (~w4556 & w51572);
assign w5115 = ~w5113 & ~w5114;
assign w5116 = w4564 & w4621;
assign w5117 = ~w4613 & ~w4616;
assign w5118 = ~w4607 & w5117;
assign w5119 = w4535 & w5117;
assign w5120 = ~w4498 & w5119;
assign w5121 = (w5116 & w5120) | (w5116 & w40249) | (w5120 & w40249);
assign w5122 = ~w5120 & w40250;
assign w5123 = ~w5121 & ~w5122;
assign w5124 = ~w1120 & ~w5115;
assign w5125 = w4838 & w5124;
assign w5126 = ~w1120 & w5123;
assign w5127 = ~w4838 & w5126;
assign w5128 = ~w5125 & ~w5127;
assign w5129 = w5112 & ~w5128;
assign w5130 = w5103 & ~w5129;
assign w5131 = w5079 & ~w5130;
assign w5132 = ~w5060 & ~w5062;
assign w5133 = (w612 & w5060) | (w612 & w44154) | (w5060 & w44154);
assign w5134 = ~w4637 & w4668;
assign w5135 = w4566 & w4743;
assign w5136 = ~w4623 & w5135;
assign w5137 = w4607 & w5135;
assign w5138 = ~w4536 & w5137;
assign w5139 = (w5134 & w5138) | (w5134 & w40252) | (w5138 & w40252);
assign w5140 = ~w5138 & w40253;
assign w5141 = ~w5139 & ~w5140;
assign w5142 = w4636 & w4838;
assign w5143 = ~w4838 & ~w5141;
assign w5144 = ~w5142 & ~w5143;
assign w5145 = w493 & ~w5144;
assign w5146 = ~w5133 & ~w5145;
assign w5147 = (w5146 & w5130) | (w5146 & w40254) | (w5130 & w40254);
assign w5148 = ~w4589 & w4838;
assign w5149 = ~w4838 & w4863;
assign w5150 = ~w5148 & ~w5149;
assign w5151 = w1541 & ~w5150;
assign w5152 = ~w4882 & w4878;
assign w5153 = (w4843 & w51573) | (w4843 & w51574) | (w51573 & w51574);
assign w5154 = ~w5152 & ~w5153;
assign w5155 = (w1738 & w4838) | (w1738 & w44155) | (w4838 & w44155);
assign w5156 = w4532 & w4838;
assign w5157 = w5155 & ~w5156;
assign w5158 = ~w5151 & ~w5157;
assign w5159 = ~w4856 & ~w4857;
assign w5160 = w4856 & w4857;
assign w5161 = ~w5159 & ~w5160;
assign w5162 = w4876 & ~w5158;
assign w5163 = w1320 & ~w5161;
assign w5164 = ~w5162 & ~w5163;
assign w5165 = w5147 & w5164;
assign w5166 = ~w5051 & w5165;
assign w5167 = ~w4687 & w51575;
assign w5168 = (w5167 & w4966) | (w5167 & w49484) | (w4966 & w49484);
assign w5169 = ~w4712 & ~w4748;
assign w5170 = w5169 & w52186;
assign w5171 = ~w4838 & w5170;
assign w5172 = ~w4703 & ~w4712;
assign w5173 = ~w4738 & ~w5172;
assign w5174 = ~w4747 & w5173;
assign w5175 = w4745 & w5173;
assign w5176 = ~w5174 & w52187;
assign w5177 = w4702 & w4838;
assign w5178 = ~w4838 & w5176;
assign w5179 = ~w5177 & ~w5178;
assign w5180 = ~w4838 & w49485;
assign w5181 = ~w5179 & ~w5180;
assign w5182 = (w252 & w5179) | (w252 & w49486) | (w5179 & w49486);
assign w5183 = ~w252 & w4838;
assign w5184 = ~w5171 & ~w5183;
assign w5185 = ~w4722 & ~w4814;
assign w5186 = w57 & ~w5185;
assign w5187 = w5184 & w5186;
assign w5188 = w57 & w5185;
assign w5189 = ~w5184 & w5188;
assign w5190 = ~w5187 & ~w5189;
assign w5191 = ~w5182 & w5190;
assign w5192 = ~w5179 & w49487;
assign w5193 = ~w4710 & w51576;
assign w5194 = (w351 & w4710) | (w351 & w51577) | (w4710 & w51577);
assign w5195 = w4203 & ~w4643;
assign w5196 = ~w4203 & w4643;
assign w5197 = ~w5195 & ~w5196;
assign w5198 = (~w5194 & ~w5197) | (~w5194 & w51578) | (~w5197 & w51578);
assign w5199 = (w4729 & w4744) | (w4729 & w51384) | (w4744 & w51384);
assign w5200 = w4729 & ~w4962;
assign w5201 = ~w4711 & ~w4738;
assign w5202 = ~w351 & w5201;
assign w5203 = (w5200 & w49488) | (w5200 & w49489) | (w49488 & w49489);
assign w5204 = ~w351 & ~w5201;
assign w5205 = (w40258 & ~w5200) | (w40258 & w49490) | (~w5200 & w49490);
assign w5206 = ~w5203 & ~w5205;
assign w5207 = ~w4838 & w5206;
assign w5208 = w351 & ~w5201;
assign w5209 = (w5200 & w49491) | (w5200 & w49492) | (w49491 & w49492);
assign w5210 = w351 & w5201;
assign w5211 = (w40260 & ~w5200) | (w40260 & w49493) | (~w5200 & w49493);
assign w5212 = ~w5209 & ~w5211;
assign w5213 = (~w4637 & w4743) | (~w4637 & w51579) | (w4743 & w51579);
assign w5214 = w4648 & w4729;
assign w5215 = ~w400 & ~w5214;
assign w5216 = w5215 & w52188;
assign w5217 = ~w400 & w5214;
assign w5218 = w5213 & w52189;
assign w5219 = ~w5216 & ~w5218;
assign w5220 = w5212 & w5219;
assign w5221 = w4838 & w51580;
assign w5222 = w5207 & ~w5220;
assign w5223 = ~w5221 & ~w5222;
assign w5224 = ~w5192 & w5223;
assign w5225 = w4963 & ~w4967;
assign w5226 = w4828 & ~w4834;
assign w5227 = (w5226 & w5225) | (w5226 & w40263) | (w5225 & w40263);
assign w5228 = ~w3 & w4838;
assign w5229 = ~w4838 & w5227;
assign w5230 = ~w5228 & ~w5229;
assign w5231 = ~w4789 & w4823;
assign w5232 = (~w42 & w4789) | (~w42 & w51581) | (w4789 & w51581);
assign w5233 = ~w5230 & w5232;
assign w5234 = ~w4789 & w51582;
assign w5235 = w5230 & w5234;
assign w5236 = ~w5233 & ~w5235;
assign w5237 = (~w4818 & w5225) | (~w4818 & w40265) | (w5225 & w40265);
assign w5238 = w80 & w4838;
assign w5239 = ~w4838 & w5237;
assign w5240 = ~w5238 & ~w5239;
assign w5241 = w4812 & w4828;
assign w5242 = ~w3 & ~w5241;
assign w5243 = ~w5240 & w5242;
assign w5244 = ~w3 & w5241;
assign w5245 = w5240 & w5244;
assign w5246 = ~w5243 & ~w5245;
assign w5247 = w5236 & w5246;
assign w5248 = ~w4802 & ~w4818;
assign w5249 = ~w4814 & w4833;
assign w5250 = ~w5225 & w5249;
assign w5251 = w5248 & w5250;
assign w5252 = ~w5248 & ~w5250;
assign w5253 = (w252 & w4406) | (w252 & w51583) | (w4406 & w51583);
assign w5254 = w4430 & ~w4795;
assign w5255 = ~w5254 & w51584;
assign w5256 = (~w4794 & w5254) | (~w4794 & w51585) | (w5254 & w51585);
assign w5257 = ~w5255 & ~w5256;
assign w5258 = w4838 & ~w5257;
assign w5259 = ~w4838 & ~w5251;
assign w5260 = (~w5258 & ~w5259) | (~w5258 & w40266) | (~w5259 & w40266);
assign w5261 = w80 & w5260;
assign w5262 = ~w57 & ~w5185;
assign w5263 = ~w5184 & w5262;
assign w5264 = ~w57 & w5185;
assign w5265 = w5184 & w5264;
assign w5266 = ~w5263 & ~w5265;
assign w5267 = ~w5261 & w5266;
assign w5268 = w5247 & w5267;
assign w5269 = w5191 & ~w5224;
assign w5270 = w5268 & ~w5269;
assign w5271 = w4838 & w51586;
assign w5272 = w5207 & w5212;
assign w5273 = w5213 & w52190;
assign w5274 = w5214 & w52188;
assign w5275 = w4838 & w5197;
assign w5276 = ~w4838 & w51588;
assign w5277 = ~w5275 & ~w5276;
assign w5278 = ~w5276 & w44156;
assign w5279 = ~w493 & w5144;
assign w5280 = ~w5278 & ~w5279;
assign w5281 = ~w5272 & w44157;
assign w5282 = w5280 & ~w5281;
assign w5283 = w5191 & w5282;
assign w5284 = w5270 & ~w5283;
assign w5285 = w1120 & w5115;
assign w5286 = w4838 & w5285;
assign w5287 = w1120 & ~w5123;
assign w5288 = ~w4838 & w5287;
assign w5289 = ~w5286 & ~w5288;
assign w5290 = w5112 & w5289;
assign w5291 = w5079 & w5290;
assign w5292 = w5146 & ~w5291;
assign w5293 = ~w5131 & w5292;
assign w5294 = ~w80 & ~w5260;
assign w5295 = w3 & ~w5241;
assign w5296 = w5240 & w5295;
assign w5297 = w3 & w5241;
assign w5298 = ~w5240 & w5297;
assign w5299 = ~w5296 & ~w5298;
assign w5300 = ~w5294 & w5299;
assign w5301 = ~w4789 & w52191;
assign w5302 = w4775 & ~w4777;
assign w5303 = w4127 & ~w4764;
assign w5304 = ~w4127 & w4764;
assign w5305 = ~w5303 & ~w5304;
assign w5306 = ~w5301 & ~w5302;
assign w5307 = ~w4407 & w5305;
assign w5308 = w5302 & w5307;
assign w5309 = w5301 & w5308;
assign w5310 = ~w5306 & ~w5309;
assign w5311 = w4430 & ~w5305;
assign w5312 = w5301 & ~w5302;
assign w5313 = w5302 & w5311;
assign w5314 = ~w5301 & w5313;
assign w5315 = ~w5312 & ~w5314;
assign w5316 = w42 & w5315;
assign w5317 = ~w42 & w5310;
assign w5318 = ~w5316 & ~w5317;
assign w5319 = w5230 & ~w5231;
assign w5320 = ~w5230 & w5231;
assign w5321 = ~w5319 & ~w5320;
assign w5322 = w42 & ~w5321;
assign w5323 = ~w5318 & ~w5322;
assign w5324 = w5247 & ~w5300;
assign w5325 = w5323 & ~w5324;
assign w5326 = ~w5293 & w5325;
assign w5327 = ~w5284 & w5326;
assign w5328 = ~w5166 & w5327;
assign w5329 = ~w5270 & w5325;
assign w5330 = ~w5328 & ~w5329;
assign w5331 = ~w4877 & ~w4890;
assign w5332 = ~w5039 & w40268;
assign w5333 = (w4903 & w5332) | (w4903 & w44158) | (w5332 & w44158);
assign w5334 = w5331 & ~w5333;
assign w5335 = ~w5331 & w5333;
assign w5336 = ~w5334 & ~w5335;
assign w5337 = (w4849 & w5328) | (w4849 & w44159) | (w5328 & w44159);
assign w5338 = ~w5328 & w44160;
assign w5339 = ~w5337 & ~w5338;
assign w5340 = (a[79] & w5328) | (a[79] & w44161) | (w5328 & w44161);
assign w5341 = ~a[79] & ~w5329;
assign w5342 = ~w5328 & w5341;
assign w5343 = ~a[76] & ~a[77];
assign w5344 = ~a[78] & w5343;
assign w5345 = w4838 & ~w5344;
assign w5346 = (w4430 & ~w4838) | (w4430 & w51589) | (~w4838 & w51589);
assign w5347 = (w5346 & w5328) | (w5346 & w44162) | (w5328 & w44162);
assign w5348 = ~w5340 & w5347;
assign w5349 = ~w4838 & w5344;
assign w5350 = ~w4838 & w51589;
assign w5351 = ~w4406 & w51590;
assign w5352 = (~w5350 & w5328) | (~w5350 & w47122) | (w5328 & w47122);
assign w5353 = ~w5348 & w5352;
assign w5354 = ~a[80] & ~w4838;
assign w5355 = a[80] & w4838;
assign w5356 = a[80] & ~w4988;
assign w5357 = ~w4989 & ~w5356;
assign w5358 = ~w5354 & ~w5355;
assign w5359 = (w5358 & w5328) | (w5358 & w44164) | (w5328 & w44164);
assign w5360 = ~w5328 & w44165;
assign w5361 = ~w5359 & ~w5360;
assign w5362 = ~w5345 & ~w5349;
assign w5363 = (w5362 & w5328) | (w5362 & w44166) | (w5328 & w44166);
assign w5364 = ~w5340 & w5363;
assign w5365 = (~w4430 & w4838) | (~w4430 & w51591) | (w4838 & w51591);
assign w5366 = (w5365 & w5328) | (w5365 & w47123) | (w5328 & w47123);
assign w5367 = ~w5364 & w5366;
assign w5368 = (w4056 & w5364) | (w4056 & w47124) | (w5364 & w47124);
assign w5369 = w5353 & w5361;
assign w5370 = w5368 & ~w5369;
assign w5371 = (w5354 & w5328) | (w5354 & w47125) | (w5328 & w47125);
assign w5372 = w4430 & ~w4838;
assign w5373 = ~w4430 & w4838;
assign w5374 = ~w5372 & ~w5373;
assign w5375 = w4989 & w5374;
assign w5376 = ~w5328 & w47126;
assign w5377 = ~w5371 & ~w5376;
assign w5378 = ~w4838 & w51592;
assign w5379 = (~w5001 & w5328) | (~w5001 & w51593) | (w5328 & w51593);
assign w5380 = ~w4989 & ~w5374;
assign w5381 = ~w5328 & w51594;
assign w5382 = a[81] & w52192;
assign w5383 = ~w5377 & w5379;
assign w5384 = ~w5381 & w5382;
assign w5385 = ~w5383 & ~w5384;
assign w5386 = ~w5370 & ~w5385;
assign w5387 = ~w5364 & w47129;
assign w5388 = ~w4056 & w5361;
assign w5389 = w5353 & w5388;
assign w5390 = ~w5387 & ~w5389;
assign w5391 = w5018 & w5031;
assign w5392 = (~w4056 & w5328) | (~w4056 & w44170) | (w5328 & w44170);
assign w5393 = ~w5328 & w44171;
assign w5394 = ~w5392 & ~w5393;
assign w5395 = w5391 & ~w5394;
assign w5396 = ~w5391 & w5394;
assign w5397 = ~w5395 & ~w5396;
assign w5398 = w3646 & w5397;
assign w5399 = w5390 & ~w5398;
assign w5400 = ~w5386 & w5399;
assign w5401 = ~w3646 & ~w5397;
assign w5402 = ~w3242 & w5045;
assign w5403 = w4942 & ~w5402;
assign w5404 = w4942 & w5045;
assign w5405 = ~w5039 & w51595;
assign w5406 = (w5404 & w5039) | (w5404 & w51596) | (w5039 & w51596);
assign w5407 = ~w5405 & ~w5406;
assign w5408 = (w5403 & w5328) | (w5403 & w44172) | (w5328 & w44172);
assign w5409 = ~w5328 & w44173;
assign w5410 = ~w5408 & ~w5409;
assign w5411 = w2896 & ~w5410;
assign w5412 = ~w4987 & ~w5037;
assign w5413 = ~w5019 & w5031;
assign w5414 = w5412 & ~w5413;
assign w5415 = ~w5412 & w5413;
assign w5416 = ~w5414 & ~w5415;
assign w5417 = (w4986 & w5328) | (w4986 & w44174) | (w5328 & w44174);
assign w5418 = ~w5328 & w44175;
assign w5419 = ~w5417 & ~w5418;
assign w5420 = ~w3242 & w5419;
assign w5421 = ~w5411 & ~w5420;
assign w5422 = ~w5401 & w5421;
assign w5423 = ~w5400 & w5422;
assign w5424 = w4913 & ~w4948;
assign w5425 = w4925 & w4931;
assign w5426 = ~w4942 & w5425;
assign w5427 = w5045 & w5425;
assign w5428 = ~w5039 & w40269;
assign w5429 = ~w5426 & ~w5428;
assign w5430 = ~w5428 & w44176;
assign w5431 = ~w4948 & w51597;
assign w5432 = ~w5428 & w44177;
assign w5433 = (~w5424 & w5428) | (~w5424 & w51598) | (w5428 & w51598);
assign w5434 = ~w5329 & w51599;
assign w5435 = (~w2285 & w5328) | (~w2285 & w51600) | (w5328 & w51600);
assign w5436 = (~w4947 & w5328) | (~w4947 & w44178) | (w5328 & w44178);
assign w5437 = w5435 & ~w5436;
assign w5438 = w4897 & w51601;
assign w5439 = (w4898 & ~w4897) | (w4898 & w51602) | (~w4897 & w51602);
assign w5440 = ~w5438 & ~w5439;
assign w5441 = w4903 & w4953;
assign w5442 = ~w4944 & ~w4948;
assign w5443 = (w5441 & w5332) | (w5441 & w51603) | (w5332 & w51603);
assign w5444 = ~w5332 & w51604;
assign w5445 = ~w5443 & ~w5444;
assign w5446 = ~w2006 & ~w5440;
assign w5447 = (w5446 & w5328) | (w5446 & w44179) | (w5328 & w44179);
assign w5448 = ~w2006 & w5445;
assign w5449 = ~w5328 & w51605;
assign w5450 = ~w5447 & ~w5449;
assign w5451 = ~w5437 & w5450;
assign w5452 = w1738 & ~w4849;
assign w5453 = (w5452 & w5328) | (w5452 & w44180) | (w5328 & w44180);
assign w5454 = w1738 & w5336;
assign w5455 = w5330 & w5454;
assign w5456 = ~w5453 & ~w5455;
assign w5457 = w2006 & w5440;
assign w5458 = (w5457 & w5328) | (w5457 & w44181) | (w5328 & w44181);
assign w5459 = w2006 & ~w5445;
assign w5460 = ~w5328 & w51606;
assign w5461 = ~w5458 & ~w5460;
assign w5462 = w5456 & w5461;
assign w5463 = ~w5451 & w5462;
assign w5464 = ~w1738 & ~w5339;
assign w5465 = ~w5050 & w40270;
assign w5466 = w4887 & ~w5157;
assign w5467 = ~w1738 & w4887;
assign w5468 = (w5467 & w5328) | (w5467 & w44182) | (w5328 & w44182);
assign w5469 = (w5466 & w5050) | (w5466 & w51607) | (w5050 & w51607);
assign w5470 = ~w5328 & w44183;
assign w5471 = ~w5468 & ~w5470;
assign w5472 = (w5157 & w5328) | (w5157 & w44184) | (w5328 & w44184);
assign w5473 = ~w5329 & w5465;
assign w5474 = ~w5466 & w5473;
assign w5475 = ~w5328 & w5474;
assign w5476 = ~w1541 & ~w5475;
assign w5477 = ~w5472 & w5476;
assign w5478 = w5471 & w5477;
assign w5479 = ~w5464 & ~w5478;
assign w5480 = ~w5463 & w5479;
assign w5481 = ~w5472 & ~w5475;
assign w5482 = w5471 & w5481;
assign w5483 = w1541 & ~w5482;
assign w5484 = (w4868 & w5151) | (w4868 & w51608) | (w5151 & w51608);
assign w5485 = w4887 & w44185;
assign w5486 = ~w5050 & w40271;
assign w5487 = ~w5484 & ~w5486;
assign w5488 = ~w1320 & w5161;
assign w5489 = ~w5163 & ~w5488;
assign w5490 = ~w5329 & w5489;
assign w5491 = w5487 & w5490;
assign w5492 = ~w5328 & w5491;
assign w5493 = ~w1320 & w5325;
assign w5494 = ~w5284 & w5493;
assign w5495 = w5147 & ~w5329;
assign w5496 = w5494 & ~w5495;
assign w5497 = (~w5489 & w5486) | (~w5489 & w44186) | (w5486 & w44186);
assign w5498 = ~w5496 & w5497;
assign w5499 = ~w5492 & ~w5498;
assign w5500 = (~w5161 & w5328) | (~w5161 & w44187) | (w5328 & w44187);
assign w5501 = w5499 & ~w5500;
assign w5502 = (~w1120 & ~w5499) | (~w1120 & w44188) | (~w5499 & w44188);
assign w5503 = w5128 & w5289;
assign w5504 = ~w5051 & w5164;
assign w5505 = ~w5051 & w44189;
assign w5506 = (~w5503 & w5051) | (~w5503 & w47130) | (w5051 & w47130);
assign w5507 = w4838 & ~w5115;
assign w5508 = ~w4838 & w5123;
assign w5509 = ~w5507 & ~w5508;
assign w5510 = ~w945 & w52193;
assign w5511 = ~w5505 & ~w5506;
assign w5512 = w5330 & w5511;
assign w5513 = w5510 & ~w5512;
assign w5514 = ~w5502 & ~w5513;
assign w5515 = w5499 & w44191;
assign w5516 = ~w5050 & w40272;
assign w5517 = w4868 & ~w5151;
assign w5518 = ~w5516 & w44192;
assign w5519 = (w5517 & w5516) | (w5517 & w44193) | (w5516 & w44193);
assign w5520 = ~w5518 & ~w5519;
assign w5521 = (w5150 & w5328) | (w5150 & w44194) | (w5328 & w44194);
assign w5522 = w5330 & ~w5520;
assign w5523 = ~w5521 & ~w5522;
assign w5524 = ~w5522 & w44195;
assign w5525 = ~w5515 & w5524;
assign w5526 = w5514 & ~w5525;
assign w5527 = ~w5483 & w5526;
assign w5528 = ~w5480 & w5527;
assign w5529 = w3242 & ~w5419;
assign w5530 = ~w5411 & w5529;
assign w5531 = ~w5039 & w51609;
assign w5532 = w4942 & ~w5425;
assign w5533 = ~w5531 & w5532;
assign w5534 = w5429 & ~w5533;
assign w5535 = (w4495 & w4919) | (w4495 & w51610) | (w4919 & w51610);
assign w5536 = ~w4919 & w51611;
assign w5537 = ~w5535 & ~w5536;
assign w5538 = ~w5328 & w44196;
assign w5539 = (~w5537 & w5328) | (~w5537 & w44197) | (w5328 & w44197);
assign w5540 = ~w5538 & ~w5539;
assign w5541 = ~w2896 & w5410;
assign w5542 = w2558 & ~w5540;
assign w5543 = ~w5541 & ~w5542;
assign w5544 = ~w5530 & w5543;
assign w5545 = (~w1320 & w5522) | (~w1320 & w44198) | (w5522 & w44198);
assign w5546 = ~w5515 & ~w5545;
assign w5547 = w5514 & ~w5546;
assign w5548 = w5102 & w5112;
assign w5549 = (w5289 & w5051) | (w5289 & w51612) | (w5051 & w51612);
assign w5550 = ~w5548 & ~w5549;
assign w5551 = w5128 & w5164;
assign w5552 = (w5290 & ~w5164) | (w5290 & w51613) | (~w5164 & w51613);
assign w5553 = w4888 & w51614;
assign w5554 = ~w5050 & w51615;
assign w5555 = (w5102 & w5554) | (w5102 & w44199) | (w5554 & w44199);
assign w5556 = ~w4838 & ~w5093;
assign w5557 = w4552 & ~w5556;
assign w5558 = ~w4552 & w5556;
assign w5559 = ~w5557 & ~w5558;
assign w5560 = (~w5559 & w5328) | (~w5559 & w51616) | (w5328 & w51616);
assign w5561 = ~w5328 & w51617;
assign w5562 = ~w5550 & w5561;
assign w5563 = ~w5560 & ~w5562;
assign w5564 = ~w5562 & w44200;
assign w5565 = (w1120 & w5328) | (w1120 & w44201) | (w5328 & w44201);
assign w5566 = ~w5328 & w44202;
assign w5567 = ~w5565 & ~w5566;
assign w5568 = w945 & w5503;
assign w5569 = w5567 & w5568;
assign w5570 = w945 & ~w5503;
assign w5571 = ~w5567 & w5570;
assign w5572 = ~w5569 & ~w5571;
assign w5573 = ~w5564 & w5572;
assign w5574 = ~w5547 & w5573;
assign w5575 = w5544 & w5574;
assign w5576 = ~w5528 & w5575;
assign w5577 = ~w5423 & w5576;
assign w5578 = (w2558 & w5328) | (w2558 & w44203) | (w5328 & w44203);
assign w5579 = ~w5328 & w44204;
assign w5580 = ~w5578 & ~w5579;
assign w5581 = ~w4948 & w51618;
assign w5582 = ~w5580 & w5581;
assign w5583 = (w2285 & w4948) | (w2285 & w51619) | (w4948 & w51619);
assign w5584 = w5580 & w5583;
assign w5585 = ~w5582 & ~w5584;
assign w5586 = ~w2558 & w5540;
assign w5587 = w5462 & ~w5586;
assign w5588 = w5585 & w5587;
assign w5589 = w5480 & ~w5588;
assign w5590 = w5527 & ~w5589;
assign w5591 = (w5574 & w5589) | (w5574 & w5772) | (w5589 & w5772);
assign w5592 = (~w5133 & w5328) | (~w5133 & w44205) | (w5328 & w44205);
assign w5593 = (w5078 & ~w5102) | (w5078 & w51620) | (~w5102 & w51620);
assign w5594 = w5103 & ~w5290;
assign w5595 = w5078 & ~w5594;
assign w5596 = w5164 & w44206;
assign w5597 = (w5595 & w5051) | (w5595 & w44207) | (w5051 & w44207);
assign w5598 = w5597 & ~w5592;
assign w5599 = ~w5133 & ~w5329;
assign w5600 = ~w5328 & w5599;
assign w5601 = ~w5064 & ~w5597;
assign w5602 = w5600 & w5601;
assign w5603 = (~w5132 & w5328) | (~w5132 & w44208) | (w5328 & w44208);
assign w5604 = ~w5602 & ~w5603;
assign w5605 = (w493 & ~w5604) | (w493 & w44209) | (~w5604 & w44209);
assign w5606 = ~w5060 & w51621;
assign w5607 = ~w493 & ~w5329;
assign w5608 = (~w5606 & w5328) | (~w5606 & w44210) | (w5328 & w44210);
assign w5609 = ~w5602 & w51622;
assign w5610 = w5078 & ~w5082;
assign w5611 = ~w5554 & w40273;
assign w5612 = ~w5554 & w44211;
assign w5613 = w5610 & ~w5611;
assign w5614 = w5330 & w51623;
assign w5615 = ~w5066 & ~w5080;
assign w5616 = ~w612 & w52194;
assign w5617 = ~w5614 & w5616;
assign w5618 = ~w5609 & ~w5617;
assign w5619 = ~w5605 & ~w5618;
assign w5620 = ~w5064 & w5597;
assign w5621 = w5600 & ~w5620;
assign w5622 = ~w5145 & ~w5279;
assign w5623 = ~w5621 & w44214;
assign w5624 = (w5622 & w5621) | (w5622 & w44215) | (w5621 & w44215);
assign w5625 = ~w5623 & ~w5624;
assign w5626 = w400 & w5625;
assign w5627 = ~w5619 & ~w5626;
assign w5628 = (w754 & w5562) | (w754 & w48649) | (w5562 & w48649);
assign w5629 = ~w5605 & ~w5628;
assign w5630 = ~w5619 & w48650;
assign w5631 = ~w400 & ~w5277;
assign w5632 = ~w5278 & ~w5631;
assign w5633 = ~w5279 & ~w5293;
assign w5634 = ~w5166 & w5633;
assign w5635 = w5330 & ~w5634;
assign w5636 = (w5632 & w5635) | (w5632 & w44217) | (w5635 & w44217);
assign w5637 = ~w5635 & w44218;
assign w5638 = ~w5636 & ~w5637;
assign w5639 = w351 & ~w5638;
assign w5640 = ~w400 & ~w5625;
assign w5641 = ~w5639 & ~w5640;
assign w5642 = (w754 & w5328) | (w754 & w48651) | (w5328 & w48651);
assign w5643 = ~w5328 & w51624;
assign w5644 = (w5610 & w5643) | (w5610 & w48652) | (w5643 & w48652);
assign w5645 = ~w5643 & w48653;
assign w5646 = ~w5644 & ~w5645;
assign w5647 = w612 & w5646;
assign w5648 = w5641 & ~w5647;
assign w5649 = ~w5630 & w5648;
assign w5650 = ~w5591 & w5649;
assign w5651 = ~w5577 & w5650;
assign w5652 = (~w5631 & w5166) | (~w5631 & w44219) | (w5166 & w44219);
assign w5653 = (w351 & w5328) | (w351 & w51625) | (w5328 & w51625);
assign w5654 = w5330 & w44220;
assign w5655 = ~w5272 & w51626;
assign w5656 = (w5655 & w5654) | (w5655 & w51627) | (w5654 & w51627);
assign w5657 = (~w252 & w5272) | (~w252 & w51628) | (w5272 & w51628);
assign w5658 = ~w5654 & w51629;
assign w5659 = ~w5656 & ~w5658;
assign w5660 = w5165 & w5224;
assign w5661 = ~w5051 & w5660;
assign w5662 = ~w5182 & w52195;
assign w5663 = ~w5661 & w5662;
assign w5664 = w5190 & w5266;
assign w5665 = ~w5328 & w5663;
assign w5666 = ~w5329 & ~w5664;
assign w5667 = w5665 & w5666;
assign w5668 = ~w5328 & ~w5663;
assign w5669 = ~w5329 & w5664;
assign w5670 = w5668 & w5669;
assign w5671 = w5184 & ~w5185;
assign w5672 = ~w5184 & w5185;
assign w5673 = ~w5671 & ~w5672;
assign w5674 = (w5673 & w5328) | (w5673 & w40275) | (w5328 & w40275);
assign w5675 = ~w5670 & ~w5674;
assign w5676 = (w80 & ~w5675) | (w80 & w40276) | (~w5675 & w40276);
assign w5677 = (~w80 & ~w5665) | (~w80 & w44221) | (~w5665 & w44221);
assign w5678 = w5675 & w5677;
assign w5679 = ~w5182 & ~w5192;
assign w5680 = w5165 & w5223;
assign w5681 = ~w5051 & w5680;
assign w5682 = (w5223 & w5293) | (w5223 & w40277) | (w5293 & w40277);
assign w5683 = (w5679 & w5681) | (w5679 & w40278) | (w5681 & w40278);
assign w5684 = w5330 & ~w5683;
assign w5685 = ~w5681 & w40279;
assign w5686 = w5330 & w44222;
assign w5687 = (~w5181 & w5328) | (~w5181 & w40280) | (w5328 & w40280);
assign w5688 = ~w57 & ~w5687;
assign w5689 = ~w5686 & w5688;
assign w5690 = ~w5678 & w5689;
assign w5691 = ~w5690 & w51630;
assign w5692 = w5191 & w52195;
assign w5693 = (w5266 & w5661) | (w5266 & w51631) | (w5661 & w51631);
assign w5694 = ~w5261 & ~w5294;
assign w5695 = (w5260 & w5328) | (w5260 & w51632) | (w5328 & w51632);
assign w5696 = w5330 & w51633;
assign w5697 = w5330 & w51634;
assign w5698 = ~w5696 & ~w5697;
assign w5699 = ~w5695 & w5698;
assign w5700 = w5698 & w40281;
assign w5701 = (w5328 & w51635) | (w5328 & w51636) | (w51635 & w51636);
assign w5702 = w57 & ~w5685;
assign w5703 = (~w5701 & ~w5684) | (~w5701 & w51637) | (~w5684 & w51637);
assign w5704 = ~w5678 & w5703;
assign w5705 = (~w5700 & w5704) | (~w5700 & w51638) | (w5704 & w51638);
assign w5706 = (w5267 & w5661) | (w5267 & w49495) | (w5661 & w49495);
assign w5707 = w5246 & w5299;
assign w5708 = (w5707 & w5706) | (w5707 & w51639) | (w5706 & w51639);
assign w5709 = w5330 & ~w5708;
assign w5710 = ~w5706 & w51640;
assign w5711 = w5240 & ~w5241;
assign w5712 = ~w5240 & w5241;
assign w5713 = ~w5711 & ~w5712;
assign w5714 = (~w5713 & w5328) | (~w5713 & w51641) | (w5328 & w51641);
assign w5715 = ~w42 & ~w5714;
assign w5716 = (w5715 & ~w5709) | (w5715 & w51642) | (~w5709 & w51642);
assign w5717 = (~w3 & ~w5698) | (~w3 & w51643) | (~w5698 & w51643);
assign w5718 = ~w5716 & ~w5717;
assign w5719 = ~w5691 & w5705;
assign w5720 = w5718 & ~w5719;
assign w5721 = w5650 & w44223;
assign w5722 = ~w5627 & w5641;
assign w5723 = ~w351 & w5638;
assign w5724 = (w252 & w5272) | (w252 & w51644) | (w5272 & w51644);
assign w5725 = (w5724 & w5654) | (w5724 & w40282) | (w5654 & w40282);
assign w5726 = ~w5272 & w51645;
assign w5727 = ~w5654 & w40283;
assign w5728 = ~w5725 & ~w5727;
assign w5729 = ~w5723 & w5728;
assign w5730 = w5705 & w5729;
assign w5731 = ~w5722 & w5730;
assign w5732 = w5720 & ~w5731;
assign w5733 = (w5246 & w5706) | (w5246 & w51646) | (w5706 & w51646);
assign w5734 = w5236 & ~w5316;
assign w5735 = ~w5322 & w5734;
assign w5736 = ~w5735 & ~w5733;
assign w5737 = ~w5236 & ~w5310;
assign w5738 = ~w5322 & ~w5737;
assign w5739 = (w5706 & w51647) | (w5706 & w51648) | (w51647 & w51648);
assign w5740 = ~w5736 & ~w5739;
assign w5741 = (~w5714 & ~w5709) | (~w5714 & w51649) | (~w5709 & w51649);
assign w5742 = w42 & ~w5741;
assign w5743 = (~w5740 & w5741) | (~w5740 & w51650) | (w5741 & w51650);
assign w5744 = ~w5732 & w5743;
assign w5745 = ~w5721 & w5744;
assign w5746 = w5456 & ~w5464;
assign w5747 = ~w5451 & w5461;
assign w5748 = w5461 & ~w5586;
assign w5749 = w5585 & w5748;
assign w5750 = ~w5747 & ~w5749;
assign w5751 = w5422 & ~w5750;
assign w5752 = ~w5544 & w5749;
assign w5753 = ~w5400 & w5751;
assign w5754 = (w5746 & w5753) | (w5746 & w40284) | (w5753 & w40284);
assign w5755 = ~w5753 & w40285;
assign w5756 = ~w5754 & ~w5755;
assign w5757 = ~w5721 & w40286;
assign w5758 = (w5756 & w5721) | (w5756 & w40287) | (w5721 & w40287);
assign w5759 = ~w5757 & ~w5758;
assign w5760 = ~w5625 & w5743;
assign w5761 = ~w5732 & w5760;
assign w5762 = w612 & ~w5609;
assign w5763 = (w5762 & w5577) | (w5762 & w40289) | (w5577 & w40289);
assign w5764 = w5422 & ~w5589;
assign w5765 = ~w5400 & w5764;
assign w5766 = ~w5544 & w5588;
assign w5767 = w5480 & ~w5766;
assign w5768 = ~w5609 & w5646;
assign w5769 = w5574 & w5768;
assign w5770 = ~w5765 & w40290;
assign w5771 = ~w612 & ~w5628;
assign w5772 = ~w5527 & w5574;
assign w5773 = ~w5626 & ~w5640;
assign w5774 = ~w5605 & ~w5773;
assign w5775 = (w5768 & w5772) | (w5768 & w40291) | (w5772 & w40291);
assign w5776 = w5774 & ~w5775;
assign w5777 = ~w5770 & w5776;
assign w5778 = ~w5721 & w5761;
assign w5779 = w5629 & ~w5647;
assign w5780 = (w5779 & w5590) | (w5779 & w40292) | (w5590 & w40292);
assign w5781 = (w5627 & w5577) | (w5627 & w40293) | (w5577 & w40293);
assign w5782 = ~w5745 & ~w5781;
assign w5783 = (~w5640 & w5732) | (~w5640 & w40294) | (w5732 & w40294);
assign w5784 = ~w5719 & w51651;
assign w5785 = w5651 & w5784;
assign w5786 = ~w5783 & ~w5785;
assign w5787 = ~w5778 & w40295;
assign w5788 = (~w351 & w5785) | (~w351 & w40296) | (w5785 & w40296);
assign w5789 = ~w5782 & w5788;
assign w5790 = ~w5787 & ~w5789;
assign w5791 = (w612 & w5577) | (w612 & w40297) | (w5577 & w40297);
assign w5792 = (w5646 & w5772) | (w5646 & w51652) | (w5772 & w51652);
assign w5793 = w5574 & w5646;
assign w5794 = ~w5765 & w40298;
assign w5795 = ~w5792 & ~w5794;
assign w5796 = ~w5791 & w5795;
assign w5797 = ~w5745 & w5796;
assign w5798 = (~w400 & w5605) | (~w400 & w51653) | (w5605 & w51653);
assign w5799 = (w5798 & w5721) | (w5798 & w40300) | (w5721 & w40300);
assign w5800 = ~w5797 & w5799;
assign w5801 = ~w5745 & ~w5796;
assign w5802 = ~w5605 & w51654;
assign w5803 = (w5802 & w5721) | (w5802 & w40302) | (w5721 & w40302);
assign w5804 = ~w5801 & w5803;
assign w5805 = ~w5800 & ~w5804;
assign w5806 = (w351 & w5778) | (w351 & w40303) | (w5778 & w40303);
assign w5807 = ~w5782 & ~w5786;
assign w5808 = w5806 & ~w5807;
assign w5809 = w5805 & ~w5808;
assign w5810 = w5790 & ~w5809;
assign w5811 = ~w5605 & w51655;
assign w5812 = (w5811 & w5721) | (w5811 & w40304) | (w5721 & w40304);
assign w5813 = ~w5797 & w5812;
assign w5814 = (w400 & w5605) | (w400 & w51656) | (w5605 & w51656);
assign w5815 = (w5814 & w5721) | (w5814 & w40305) | (w5721 & w40305);
assign w5816 = ~w5801 & w5815;
assign w5817 = ~w5813 & ~w5816;
assign w5818 = w5790 & w5817;
assign w5819 = ~w5547 & w5572;
assign w5820 = w5480 & w5544;
assign w5821 = (w5819 & w5589) | (w5819 & w48654) | (w5589 & w48654);
assign w5822 = w5819 & w5820;
assign w5823 = ~w5423 & w5822;
assign w5824 = ~w5564 & ~w5628;
assign w5825 = (w5824 & w5823) | (w5824 & w40306) | (w5823 & w40306);
assign w5826 = ~w5745 & w40307;
assign w5827 = ~w493 & ~w5646;
assign w5828 = (w5827 & ~w40307) | (w5827 & w50272) | (~w40307 & w50272);
assign w5829 = ~w493 & w5646;
assign w5830 = w40307 & w50273;
assign w5831 = ~w5828 & ~w5830;
assign w5832 = w5818 & w5831;
assign w5833 = ~w5810 & ~w5832;
assign w5834 = w5659 & w5728;
assign w5835 = ~w5722 & ~w5723;
assign w5836 = ~w5651 & w40308;
assign w5837 = (w5834 & w5651) | (w5834 & w51657) | (w5651 & w51657);
assign w5838 = w252 & w5728;
assign w5839 = w5659 & ~w5838;
assign w5840 = ~w5721 & w51658;
assign w5841 = ~w5745 & w51659;
assign w5842 = ~w5840 & ~w5841;
assign w5843 = (w57 & w5841) | (w57 & w48655) | (w5841 & w48655);
assign w5844 = ~w5841 & w40309;
assign w5845 = ~w5721 & w40310;
assign w5846 = ~w5640 & ~w5781;
assign w5847 = ~w5745 & w5846;
assign w5848 = ~w5639 & ~w5723;
assign w5849 = w252 & ~w5848;
assign w5850 = (w5849 & w5847) | (w5849 & w40311) | (w5847 & w40311);
assign w5851 = w252 & w5848;
assign w5852 = ~w5847 & w40312;
assign w5853 = ~w5850 & ~w5852;
assign w5854 = (~w5843 & w5853) | (~w5843 & w51660) | (w5853 & w51660);
assign w5855 = ~w5833 & w5854;
assign w5856 = ~w5386 & w5390;
assign w5857 = ~w5398 & ~w5401;
assign w5858 = (~w3242 & w5856) | (~w3242 & w51661) | (w5856 & w51661);
assign w5859 = w5856 & w5857;
assign w5860 = w5858 & ~w5859;
assign w5861 = ~w3242 & ~w5397;
assign w5862 = ~w5721 & w40313;
assign w5863 = (w5860 & w5721) | (w5860 & w40314) | (w5721 & w40314);
assign w5864 = ~w5862 & ~w5863;
assign w5865 = ~w5420 & ~w5529;
assign w5866 = ~w5400 & w51662;
assign w5867 = (w5865 & w5400) | (w5865 & w51663) | (w5400 & w51663);
assign w5868 = ~w5866 & ~w5867;
assign w5869 = w2896 & w5419;
assign w5870 = ~w5721 & w40315;
assign w5871 = w2896 & w5868;
assign w5872 = (w5871 & w5721) | (w5871 & w51664) | (w5721 & w51664);
assign w5873 = ~w5870 & ~w5872;
assign w5874 = w5864 & w5873;
assign w5875 = ~w5370 & w5390;
assign w5876 = (w5875 & w5732) | (w5875 & w40316) | (w5732 & w40316);
assign w5877 = ~w5719 & w51665;
assign w5878 = w5651 & w5877;
assign w5879 = w3242 & w5397;
assign w5880 = ~w5732 & w40317;
assign w5881 = ~w5721 & w5880;
assign w5882 = w3242 & ~w5857;
assign w5883 = ~w5856 & w5882;
assign w5884 = w3242 & w5857;
assign w5885 = w5856 & w5884;
assign w5886 = ~w5883 & ~w5885;
assign w5887 = (~w5886 & w5732) | (~w5886 & w44224) | (w5732 & w44224);
assign w5888 = w5720 & ~w5886;
assign w5889 = w5651 & w5888;
assign w5890 = ~w5887 & ~w5889;
assign w5891 = ~w5881 & w5890;
assign w5892 = (w3646 & w5383) | (w3646 & w51666) | (w5383 & w51666);
assign w5893 = ~w5878 & w51667;
assign w5894 = w3646 & w5385;
assign w5895 = (w5894 & w5878) | (w5894 & w40318) | (w5878 & w40318);
assign w5896 = w5891 & w51668;
assign w5897 = w5874 & ~w5896;
assign w5898 = ~w5732 & w40319;
assign w5899 = ~w5721 & w5898;
assign w5900 = (~w5420 & w5397) | (~w5420 & w51669) | (w5397 & w51669);
assign w5901 = (~w5529 & w5400) | (~w5529 & w40320) | (w5400 & w40320);
assign w5902 = (~w5901 & w5732) | (~w5901 & w44225) | (w5732 & w44225);
assign w5903 = w5720 & ~w5901;
assign w5904 = w5651 & w5903;
assign w5905 = ~w5902 & ~w5904;
assign w5906 = ~w5411 & ~w5541;
assign w5907 = w2558 & ~w5906;
assign w5908 = (w5907 & ~w5905) | (w5907 & w44226) | (~w5905 & w44226);
assign w5909 = w2558 & w5906;
assign w5910 = w5905 & w44227;
assign w5911 = ~w5908 & ~w5910;
assign w5912 = ~w2896 & ~w5868;
assign w5913 = (w5912 & w5721) | (w5912 & w51670) | (w5721 & w51670);
assign w5914 = ~w5721 & w51671;
assign w5915 = ~w5913 & ~w5914;
assign w5916 = w5911 & w5915;
assign w5917 = ~w5897 & w5916;
assign w5918 = w5424 & ~w5580;
assign w5919 = ~w5424 & w5580;
assign w5920 = ~w5918 & ~w5919;
assign w5921 = ~w5437 & w5585;
assign w5922 = w5585 & w40321;
assign w5923 = ~w5544 & w5922;
assign w5924 = w5422 & w5922;
assign w5925 = ~w5400 & w5924;
assign w5926 = (w5586 & ~w5585) | (w5586 & w51672) | (~w5585 & w51672);
assign w5927 = ~w5925 & w40322;
assign w5928 = w5544 & ~w5921;
assign w5929 = (w5928 & w5400) | (w5928 & w51673) | (w5400 & w51673);
assign w5930 = w5927 & ~w5929;
assign w5931 = ~w5721 & w40323;
assign w5932 = (w5930 & w5721) | (w5930 & w40324) | (w5721 & w40324);
assign w5933 = ~w5931 & ~w5932;
assign w5934 = (~w2006 & w5932) | (~w2006 & w47131) | (w5932 & w47131);
assign w5935 = w5450 & w5461;
assign w5936 = (~w5935 & w5925) | (~w5935 & w40325) | (w5925 & w40325);
assign w5937 = w5437 & ~w5935;
assign w5938 = ~w5437 & w5935;
assign w5939 = ~w5937 & ~w5938;
assign w5940 = ~w5925 & w40326;
assign w5941 = ~w5936 & ~w5940;
assign w5942 = (w5941 & w5721) | (w5941 & w40327) | (w5721 & w40327);
assign w5943 = (w5440 & w5328) | (w5440 & w51674) | (w5328 & w51674);
assign w5944 = ~w5328 & w51675;
assign w5945 = ~w5943 & ~w5944;
assign w5946 = (~w1738 & w5721) | (~w1738 & w40329) | (w5721 & w40329);
assign w5947 = ~w5942 & w5946;
assign w5948 = ~w5530 & ~w5541;
assign w5949 = (w5948 & w5400) | (w5948 & w40330) | (w5400 & w40330);
assign w5950 = w3096 & w5540;
assign w5951 = ~w3096 & ~w5540;
assign w5952 = ~w5950 & ~w5951;
assign w5953 = w5949 & w5952;
assign w5954 = ~w5949 & ~w5952;
assign w5955 = ~w5953 & ~w5954;
assign w5956 = ~w2285 & ~w5540;
assign w5957 = ~w5721 & w40331;
assign w5958 = ~w2285 & ~w5955;
assign w5959 = ~w5745 & w5958;
assign w5960 = ~w5957 & ~w5959;
assign w5961 = ~w5947 & w5960;
assign w5962 = ~w5934 & w5961;
assign w5963 = (~w1541 & w5758) | (~w1541 & w49496) | (w5758 & w49496);
assign w5964 = ~w5478 & ~w5483;
assign w5965 = (~w5464 & ~w5462) | (~w5464 & w51676) | (~w5462 & w51676);
assign w5966 = ~w5588 & w5965;
assign w5967 = w5544 & w5965;
assign w5968 = ~w5966 & w52196;
assign w5969 = w5964 & w5968;
assign w5970 = ~w5964 & ~w5968;
assign w5971 = ~w5969 & ~w5970;
assign w5972 = ~w5745 & w5971;
assign w5973 = (~w1320 & w5972) | (~w1320 & w40334) | (w5972 & w40334);
assign w5974 = ~w5963 & ~w5973;
assign w5975 = w5962 & w5974;
assign w5976 = w5917 & w5975;
assign w5977 = ~a[74] & ~a[75];
assign w5978 = ~a[76] & w5977;
assign w5979 = ~w5328 & w51677;
assign w5980 = a[76] & ~a[77];
assign w5981 = (~w5980 & w5328) | (~w5980 & w51678) | (w5328 & w51678);
assign w5982 = ~w5719 & w51679;
assign w5983 = w5651 & w5982;
assign w5984 = (~w5978 & w5328) | (~w5978 & w51680) | (w5328 & w51680);
assign w5985 = w5743 & ~w5984;
assign w5986 = a[77] & ~w5984;
assign w5987 = (~w5986 & w5732) | (~w5986 & w40336) | (w5732 & w40336);
assign w5988 = ~w5719 & w49497;
assign w5989 = w5651 & w5988;
assign w5990 = ~w5987 & ~w5989;
assign w5991 = a[77] & w5743;
assign w5992 = ~w5732 & w5991;
assign w5993 = (~w4838 & w5732) | (~w4838 & w40337) | (w5732 & w40337);
assign w5994 = ~w5719 & w49498;
assign w5995 = w5651 & w5994;
assign w5996 = ~w5993 & ~w5995;
assign w5997 = (~w4838 & w5983) | (~w4838 & w40338) | (w5983 & w40338);
assign w5998 = w5990 & ~w5996;
assign w5999 = ~w5997 & ~w5998;
assign w6000 = ~w5328 & w51681;
assign w6001 = (a[78] & w5328) | (a[78] & w51682) | (w5328 & w51682);
assign w6002 = ~w6000 & ~w6001;
assign w6003 = ~w5732 & w40339;
assign w6004 = ~w5721 & w6003;
assign w6005 = a[78] & ~w5343;
assign w6006 = ~w5344 & ~w6005;
assign w6007 = (w6006 & w5732) | (w6006 & w40340) | (w5732 & w40340);
assign w6008 = ~w5719 & w51683;
assign w6009 = w5651 & w6008;
assign w6010 = ~w6007 & ~w6009;
assign w6011 = ~w6004 & w6010;
assign w6012 = ~w5721 & w5992;
assign w6013 = w5990 & ~w6012;
assign w6014 = ~w5983 & w40341;
assign w6015 = ~w6013 & w6014;
assign w6016 = (w4430 & w6013) | (w4430 & w40342) | (w6013 & w40342);
assign w6017 = w5999 & w6011;
assign w6018 = w6016 & ~w6017;
assign w6019 = (a[79] & w5328) | (a[79] & w51684) | (w5328 & w51684);
assign w6020 = ~w5328 & w51685;
assign w6021 = ~w6019 & ~w6020;
assign w6022 = ~w5340 & ~w5342;
assign w6023 = ~w5362 & ~w6022;
assign w6024 = w4988 & ~w5343;
assign w6025 = w4838 & w6024;
assign w6026 = ~w5364 & ~w6025;
assign w6027 = (w4838 & w5328) | (w4838 & w51686) | (w5328 & w51686);
assign w6028 = ~w6023 & w6026;
assign w6029 = (w5328 & w6025) | (w5328 & w51687) | (w6025 & w51687);
assign w6030 = ~w6028 & ~w6029;
assign w6031 = ~w5721 & w51688;
assign w6032 = (w6030 & w5721) | (w6030 & w51689) | (w5721 & w51689);
assign w6033 = ~w6031 & ~w6032;
assign w6034 = (~w6033 & w6017) | (~w6033 & w40343) | (w6017 & w40343);
assign w6035 = w6010 & w44228;
assign w6036 = w5999 & w6035;
assign w6037 = ~w5983 & w40344;
assign w6038 = ~w6013 & w6037;
assign w6039 = w5353 & ~w5367;
assign w6040 = (w6039 & w5732) | (w6039 & w40345) | (w5732 & w40345);
assign w6041 = ~w5719 & w51690;
assign w6042 = w5651 & w6041;
assign w6043 = ~w4056 & ~w5361;
assign w6044 = (w6043 & w6042) | (w6043 & w40346) | (w6042 & w40346);
assign w6045 = ~w6042 & w40347;
assign w6046 = ~w6044 & ~w6045;
assign w6047 = ~w6038 & w6046;
assign w6048 = ~w6036 & w6047;
assign w6049 = ~w6034 & w6048;
assign w6050 = (w5361 & w6042) | (w5361 & w40348) | (w6042 & w40348);
assign w6051 = ~w6042 & w40349;
assign w6052 = ~w6050 & ~w6051;
assign w6053 = w4056 & ~w6052;
assign w6054 = (w5385 & w5878) | (w5385 & w40350) | (w5878 & w40350);
assign w6055 = ~w5878 & w40351;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = w5890 & w44229;
assign w6058 = w6056 & w6057;
assign w6059 = ~w6058 & w51691;
assign w6060 = ~w6049 & w6059;
assign w6061 = w5976 & ~w6060;
assign w6062 = ~w5766 & w40352;
assign w6063 = ~w5524 & ~w5545;
assign w6064 = w5483 & ~w6063;
assign w6065 = ~w5483 & w6063;
assign w6066 = ~w6064 & ~w6065;
assign w6067 = ~w5765 & w40353;
assign w6068 = (w6066 & w5765) | (w6066 & w40354) | (w5765 & w40354);
assign w6069 = ~w6067 & ~w6068;
assign w6070 = ~w5732 & w40355;
assign w6071 = ~w5721 & w6070;
assign w6072 = (~w6069 & w5721) | (~w6069 & w40356) | (w5721 & w40356);
assign w6073 = ~w6071 & ~w6072;
assign w6074 = ~w6072 & w44230;
assign w6075 = ~w5972 & w40357;
assign w6076 = ~w6074 & ~w6075;
assign w6077 = ~w5974 & w6076;
assign w6078 = ~w2558 & ~w5906;
assign w6079 = (w5400 & w51692) | (w5400 & w51693) | (w51692 & w51693);
assign w6080 = ~w5410 & w51694;
assign w6081 = ~w5721 & w40358;
assign w6082 = (w6079 & w5721) | (w6079 & w40359) | (w5721 & w40359);
assign w6083 = ~w6081 & ~w6082;
assign w6084 = ~w2558 & w5906;
assign w6085 = (w6084 & ~w5905) | (w6084 & w44231) | (~w5905 & w44231);
assign w6086 = w6083 & ~w6085;
assign w6087 = w2285 & w5540;
assign w6088 = (w5955 & w5721) | (w5955 & w51695) | (w5721 & w51695);
assign w6089 = ~w5956 & ~w6087;
assign w6090 = ~w5721 & w51696;
assign w6091 = ~w6088 & ~w6090;
assign w6092 = ~w6085 & w51697;
assign w6093 = w5962 & ~w6092;
assign w6094 = (w2006 & ~w5927) | (w2006 & w51698) | (~w5927 & w51698);
assign w6095 = (w6094 & w5721) | (w6094 & w51699) | (w5721 & w51699);
assign w6096 = w2006 & ~w5920;
assign w6097 = ~w5721 & w40360;
assign w6098 = ~w6095 & ~w6097;
assign w6099 = ~w5947 & ~w6098;
assign w6100 = ~w5721 & w40361;
assign w6101 = w1738 & w5941;
assign w6102 = ~w5745 & w6101;
assign w6103 = ~w6100 & ~w6102;
assign w6104 = w1541 & w5339;
assign w6105 = ~w5721 & w40362;
assign w6106 = w1541 & ~w5756;
assign w6107 = ~w5745 & w6106;
assign w6108 = ~w6105 & ~w6107;
assign w6109 = w6103 & w6108;
assign w6110 = ~w6099 & w6109;
assign w6111 = w6076 & w6110;
assign w6112 = ~w6093 & w6111;
assign w6113 = ~w6077 & ~w6112;
assign w6114 = ~w6061 & ~w6113;
assign w6115 = ~w5689 & w5703;
assign w6116 = ~w5722 & w5729;
assign w6117 = (~w5651 & w51700) | (~w5651 & w51701) | (w51700 & w51701);
assign w6118 = w5659 & ~w6115;
assign w6119 = (w6118 & w5651) | (w6118 & w40364) | (w5651 & w40364);
assign w6120 = ~w5686 & ~w5687;
assign w6121 = ~w5721 & w51702;
assign w6122 = ~w5745 & w51703;
assign w6123 = ~w6122 & w40365;
assign w6124 = ~w5676 & ~w5678;
assign w6125 = (~w5689 & w5659) | (~w5689 & w51704) | (w5659 & w51704);
assign w6126 = (w6125 & w5651) | (w6125 & w40366) | (w5651 & w40366);
assign w6127 = ~w5721 & w51705;
assign w6128 = ~w5745 & w6126;
assign w6129 = w3 & ~w6124;
assign w6130 = (w6129 & w6128) | (w6129 & w51706) | (w6128 & w51706);
assign w6131 = w3 & w6124;
assign w6132 = ~w6128 & w51707;
assign w6133 = ~w6130 & ~w6132;
assign w6134 = ~w6123 & w6133;
assign w6135 = (w5651 & w51708) | (w5651 & w51709) | (w51708 & w51709);
assign w6136 = w5321 & ~w5733;
assign w6137 = ~w5739 & ~w6136;
assign w6138 = w5716 & w6137;
assign w6139 = w6135 & ~w6138;
assign w6140 = (w5706 & w51710) | (w5706 & w51711) | (w51710 & w51711);
assign w6141 = ~w5733 & w51712;
assign w6142 = ~w6140 & ~w6141;
assign w6143 = ~w5716 & ~w5742;
assign w6144 = w5741 & w6142;
assign w6145 = w6143 & ~w6144;
assign w6146 = w6135 & w51713;
assign w6147 = ~w6135 & ~w6145;
assign w6148 = ~w6146 & ~w6147;
assign w6149 = w5716 & ~w5740;
assign w6150 = (~w6149 & w5704) | (~w6149 & w51714) | (w5704 & w51714);
assign w6151 = (~w5651 & w51715) | (~w5651 & w51716) | (w51715 & w51716);
assign w6152 = w5700 & ~w6151;
assign w6153 = ~w5721 & w51717;
assign w6154 = w6135 & ~w6153;
assign w6155 = (~w3 & w5704) | (~w3 & w51718) | (w5704 & w51718);
assign w6156 = (w5651 & w51719) | (w5651 & w51720) | (w51719 & w51720);
assign w6157 = ~w5699 & ~w6156;
assign w6158 = (w42 & w6156) | (w42 & w51721) | (w6156 & w51721);
assign w6159 = (w6158 & ~w6154) | (w6158 & w51722) | (~w6154 & w51722);
assign w6160 = ~w6148 & ~w6159;
assign w6161 = (w6124 & w6128) | (w6124 & w51723) | (w6128 & w51723);
assign w6162 = ~w6128 & w51724;
assign w6163 = ~w6161 & ~w6162;
assign w6164 = ~w3 & ~w6163;
assign w6165 = ~w6134 & ~w6164;
assign w6166 = w6160 & ~w6165;
assign w6167 = w493 & w5646;
assign w6168 = (w6167 & ~w40307) | (w6167 & w50274) | (~w40307 & w50274);
assign w6169 = w493 & ~w5646;
assign w6170 = w40307 & w50275;
assign w6171 = ~w6168 & ~w6170;
assign w6172 = w5818 & ~w6171;
assign w6173 = ~w5810 & ~w6172;
assign w6174 = ~w5823 & w40368;
assign w6175 = ~w5825 & ~w6174;
assign w6176 = ~w5721 & w40369;
assign w6177 = ~w5745 & w6175;
assign w6178 = ~w6176 & ~w6177;
assign w6179 = (w612 & w6177) | (w612 & w40370) | (w6177 & w40370);
assign w6180 = ~w5513 & w5572;
assign w6181 = (~w754 & ~w5572) | (~w754 & w51725) | (~w5572 & w51725);
assign w6182 = ~w5589 & w6065;
assign w6183 = w5480 & w51726;
assign w6184 = ~w5423 & w6183;
assign w6185 = ~w6184 & w40371;
assign w6186 = w945 & w6181;
assign w6187 = ~w5721 & w40372;
assign w6188 = w6181 & w6185;
assign w6189 = ~w5745 & w6188;
assign w6190 = ~w6187 & ~w6189;
assign w6191 = w5572 & w51727;
assign w6192 = ~w6185 & w6191;
assign w6193 = ~w5745 & w6192;
assign w6194 = ~w945 & w6191;
assign w6195 = ~w5721 & w40373;
assign w6196 = ~w6193 & ~w6195;
assign w6197 = w6190 & w6196;
assign w6198 = ~w6177 & w40374;
assign w6199 = w6197 & ~w6198;
assign w6200 = (~w6179 & ~w6197) | (~w6179 & w40375) | (~w6197 & w40375);
assign w6201 = ~w5502 & ~w5515;
assign w6202 = (w5820 & w5400) | (w5820 & w40376) | (w5400 & w40376);
assign w6203 = w5545 & ~w6201;
assign w6204 = ~w5589 & w48656;
assign w6205 = (~w6203 & w6202) | (~w6203 & w48657) | (w6202 & w48657);
assign w6206 = (~w5502 & w6184) | (~w5502 & w40377) | (w6184 & w40377);
assign w6207 = w6205 & ~w6206;
assign w6208 = ~w5745 & w6207;
assign w6209 = ~w5732 & w40378;
assign w6210 = ~w5721 & w6209;
assign w6211 = ~w6208 & ~w6210;
assign w6212 = (~w945 & w6208) | (~w945 & w40379) | (w6208 & w40379);
assign w6213 = w5572 & w51728;
assign w6214 = w945 & w6213;
assign w6215 = ~w5721 & w40380;
assign w6216 = w6185 & w6213;
assign w6217 = ~w5745 & w6216;
assign w6218 = ~w6215 & ~w6217;
assign w6219 = (w754 & ~w5572) | (w754 & w51729) | (~w5572 & w51729);
assign w6220 = ~w6185 & w6219;
assign w6221 = ~w5745 & w6220;
assign w6222 = ~w945 & w6219;
assign w6223 = ~w5721 & w40381;
assign w6224 = ~w6221 & ~w6223;
assign w6225 = w6218 & w6224;
assign w6226 = ~w6212 & w6225;
assign w6227 = w6225 & w40382;
assign w6228 = ~w6200 & ~w6227;
assign w6229 = w6173 & ~w6228;
assign w6230 = w6166 & ~w6229;
assign w6231 = ~w5721 & w40383;
assign w6232 = w1120 & ~w6069;
assign w6233 = ~w5745 & w6232;
assign w6234 = ~w6231 & ~w6233;
assign w6235 = (w945 & w5721) | (w945 & w40384) | (w5721 & w40384);
assign w6236 = ~w6208 & w6235;
assign w6237 = w6234 & ~w6236;
assign w6238 = ~w6179 & ~w6237;
assign w6239 = w6226 & w6238;
assign w6240 = ~w6200 & ~w6239;
assign w6241 = w6240 & w40385;
assign w6242 = ~w6230 & ~w6241;
assign w6243 = ~w6242 & w40386;
assign w6244 = (~w6157 & ~w6154) | (~w6157 & w49499) | (~w6154 & w49499);
assign w6245 = w5741 & ~w6135;
assign w6246 = ~w6139 & ~w6245;
assign w6247 = ~w42 & ~w6246;
assign w6248 = ~w6244 & w6247;
assign w6249 = (~w6248 & w6165) | (~w6248 & w40387) | (w6165 & w40387);
assign w6250 = ~w252 & w5848;
assign w6251 = (w6250 & w5847) | (w6250 & w40388) | (w5847 & w40388);
assign w6252 = ~w252 & ~w5848;
assign w6253 = ~w5847 & w40389;
assign w6254 = ~w6251 & ~w6253;
assign w6255 = ~w5844 & w6254;
assign w6256 = (~w5843 & ~w6254) | (~w5843 & w51660) | (~w6254 & w51660);
assign w6257 = ~w6255 & w48658;
assign w6258 = (w80 & w6122) | (w80 & w51730) | (w6122 & w51730);
assign w6259 = ~w6164 & ~w6258;
assign w6260 = w6259 & w48659;
assign w6261 = w5855 & w6230;
assign w6262 = ~w6249 & ~w6260;
assign w6263 = (~w6262 & ~w6230) | (~w6262 & w52106) | (~w6230 & w52106);
assign w6264 = ~w6243 & w6263;
assign w6265 = (w6092 & ~w5916) | (w6092 & w51731) | (~w5916 & w51731);
assign w6266 = w6059 & w6092;
assign w6267 = ~w6049 & w6266;
assign w6268 = (~w5963 & ~w6109) | (~w5963 & w51732) | (~w6109 & w51732);
assign w6269 = w5961 & w49500;
assign w6270 = (~w6268 & w6267) | (~w6268 & w49501) | (w6267 & w49501);
assign w6271 = ~w6099 & w6103;
assign w6272 = ~w5963 & w6108;
assign w6273 = w6271 & ~w6272;
assign w6274 = ~w6267 & w49502;
assign w6275 = w6273 & ~w6274;
assign w6276 = (~w49501 & w51733) | (~w49501 & w51734) | (w51733 & w51734);
assign w6277 = ~w6275 & ~w6276;
assign w6278 = (w5759 & w6243) | (w5759 & w52107) | (w6243 & w52107);
assign w6279 = ~w6243 & w52108;
assign w6280 = ~w6278 & ~w6279;
assign w6281 = w6163 & ~w6264;
assign w6282 = w6133 & ~w6164;
assign w6283 = w5833 & ~w6228;
assign w6284 = ~w6229 & ~w6283;
assign w6285 = w6114 & ~w6284;
assign w6286 = w6173 & ~w6240;
assign w6287 = ~w5833 & ~w6286;
assign w6288 = (~w6256 & w6285) | (~w6256 & w44232) | (w6285 & w44232);
assign w6289 = (~w6285 & w6257) | (~w6285 & w47135) | (w6257 & w47135);
assign w6290 = ~w6258 & ~w6289;
assign w6291 = w6264 & w6282;
assign w6292 = ~w6290 & w6291;
assign w6293 = w6264 & ~w6282;
assign w6294 = w6290 & w6293;
assign w6295 = ~w6292 & ~w6294;
assign w6296 = ~w6281 & w6295;
assign w6297 = ~w6257 & w6259;
assign w6298 = w6244 & w52197;
assign w6299 = (w47137 & w48660) | (w47137 & w48661) | (w48660 & w48661);
assign w6300 = ~w6298 & ~w6299;
assign w6301 = ~w6248 & w6300;
assign w6302 = w42 & w6264;
assign w6303 = ~w6300 & w6302;
assign w6304 = w6300 & w51735;
assign w6305 = ~w6303 & ~w6304;
assign w6306 = (w42 & ~w6295) | (w42 & w48662) | (~w6295 & w48662);
assign w6307 = w6305 & ~w6306;
assign w6308 = (~w42 & w6264) | (~w42 & w51736) | (w6264 & w51736);
assign w6309 = w6295 & w48663;
assign w6310 = ~w6123 & ~w6258;
assign w6311 = (w80 & w6243) | (w80 & w52109) | (w6243 & w52109);
assign w6312 = w6264 & ~w6288;
assign w6313 = (w6310 & w6312) | (w6310 & w52110) | (w6312 & w52110);
assign w6314 = ~w6312 & w52111;
assign w6315 = ~w6313 & ~w6314;
assign w6316 = w3 & ~w6315;
assign w6317 = ~w6309 & w6316;
assign w6318 = w6307 & ~w6317;
assign w6319 = ~a[72] & ~a[73];
assign w6320 = ~a[74] & w6319;
assign w6321 = ~w5721 & w51737;
assign w6322 = a[75] & ~w6249;
assign w6323 = ~w6321 & ~w6322;
assign w6324 = w6199 & w6237;
assign w6325 = ~w5833 & w51738;
assign w6326 = ~w6114 & w6325;
assign w6327 = w5855 & ~w6173;
assign w6328 = w6260 & ~w6327;
assign w6329 = ~w5833 & w40391;
assign w6330 = ~w6321 & ~w6329;
assign w6331 = w6328 & w6330;
assign w6332 = (~w6323 & ~w6331) | (~w6323 & w40392) | (~w6331 & w40392);
assign w6333 = ~w6261 & w48664;
assign w6334 = ~w6243 & w6333;
assign w6335 = ~w6332 & ~w6334;
assign w6336 = ~w6061 & w44234;
assign w6337 = ~w5855 & w6297;
assign w6338 = w6166 & w6240;
assign w6339 = ~w6337 & w6338;
assign w6340 = ~w6336 & w6339;
assign w6341 = (~w6249 & w6327) | (~w6249 & w6262) | (w6327 & w6262);
assign w6342 = a[74] & ~a[75];
assign w6343 = (w6342 & w40393) | (w6342 & w6328) | (w40393 & w6328);
assign w6344 = ~w6340 & w6343;
assign w6345 = (w6320 & w5721) | (w6320 & w51739) | (w5721 & w51739);
assign w6346 = (w5330 & w6335) | (w5330 & w40394) | (w6335 & w40394);
assign w6347 = ~w5330 & ~w6345;
assign w6348 = (w6347 & w6340) | (w6347 & w51740) | (w6340 & w51740);
assign w6349 = ~w6335 & w6348;
assign w6350 = (~a[76] & w5721) | (~a[76] & w51741) | (w5721 & w51741);
assign w6351 = ~w5721 & w51742;
assign w6352 = a[76] & ~w5977;
assign w6353 = ~w5978 & ~w6352;
assign w6354 = ~w6341 & w6353;
assign w6355 = ~w6340 & w6354;
assign w6356 = ~w6350 & ~w6351;
assign w6357 = ~w6264 & w6356;
assign w6358 = ~w6355 & ~w6357;
assign w6359 = ~w6349 & ~w6358;
assign w6360 = ~w6346 & ~w6359;
assign w6361 = a[77] & w6350;
assign w6362 = ~w5979 & ~w5984;
assign w6363 = ~w5721 & w51743;
assign w6364 = (w6362 & w5721) | (w6362 & w51744) | (w5721 & w51744);
assign w6365 = a[77] & ~w6364;
assign w6366 = ~a[77] & w6364;
assign w6367 = ~w6365 & ~w6366;
assign w6368 = ~w6363 & ~w6367;
assign w6369 = ~w6261 & w48665;
assign w6370 = (~w4838 & ~w6369) | (~w4838 & w40395) | (~w6369 & w40395);
assign w6371 = (~w6361 & w6243) | (~w6361 & w44235) | (w6243 & w44235);
assign w6372 = w6370 & ~w6371;
assign w6373 = ~a[77] & ~w6350;
assign w6374 = ~w6350 & w51745;
assign w6375 = (w6374 & ~w44236) | (w6374 & w48666) | (~w44236 & w48666);
assign w6376 = ~w6372 & ~w6375;
assign w6377 = ~w6359 & w40396;
assign w6378 = w5999 & ~w6015;
assign w6379 = ~w6261 & w48667;
assign w6380 = (w6011 & ~w6379) | (w6011 & w40397) | (~w6379 & w40397);
assign w6381 = w6379 & w40398;
assign w6382 = ~w6380 & ~w6381;
assign w6383 = ~w4430 & ~w6382;
assign w6384 = ~w6363 & w6367;
assign w6385 = (w6384 & w40399) | (w6384 & w6328) | (w40399 & w6328);
assign w6386 = a[77] & w6363;
assign w6387 = (~w6386 & w6340) | (~w6386 & w51746) | (w6340 & w51746);
assign w6388 = ~w6361 & ~w6373;
assign w6389 = ~w6264 & w6388;
assign w6390 = w6387 & ~w6389;
assign w6391 = (w4838 & w6389) | (w4838 & w51747) | (w6389 & w51747);
assign w6392 = ~w6383 & ~w6391;
assign w6393 = ~w6377 & w6392;
assign w6394 = ~w6048 & ~w6053;
assign w6395 = ~w6033 & ~w6053;
assign w6396 = ~w6018 & w6395;
assign w6397 = ~w6394 & ~w6396;
assign w6398 = ~w3646 & w6397;
assign w6399 = w3646 & ~w6397;
assign w6400 = ~w6398 & ~w6399;
assign w6401 = ~w6261 & w48668;
assign w6402 = ~w3242 & w6056;
assign w6403 = (w6402 & ~w6401) | (w6402 & w40400) | (~w6401 & w40400);
assign w6404 = ~w3242 & ~w6056;
assign w6405 = w6401 & w40401;
assign w6406 = ~w6403 & ~w6405;
assign w6407 = ~w6036 & ~w6038;
assign w6408 = ~w6034 & w6407;
assign w6409 = w6046 & ~w6053;
assign w6410 = w6408 & ~w6409;
assign w6411 = ~w6408 & w6409;
assign w6412 = ~w6410 & ~w6411;
assign w6413 = ~w3646 & ~w6052;
assign w6414 = (w6413 & w6243) | (w6413 & w44237) | (w6243 & w44237);
assign w6415 = ~w3646 & ~w6412;
assign w6416 = ~w6243 & w44238;
assign w6417 = ~w6414 & ~w6416;
assign w6418 = w6406 & w6417;
assign w6419 = w6034 & w6407;
assign w6420 = ~w6261 & w48669;
assign w6421 = ~w6243 & w6420;
assign w6422 = ~w6018 & w6407;
assign w6423 = ~w6261 & w48670;
assign w6424 = (w6033 & ~w6423) | (w6033 & w40402) | (~w6423 & w40402);
assign w6425 = ~w6421 & ~w6424;
assign w6426 = (w4056 & w6424) | (w4056 & w44239) | (w6424 & w44239);
assign w6427 = w4430 & w6382;
assign w6428 = w6418 & ~w6426;
assign w6429 = ~w6427 & w6428;
assign w6430 = (w6056 & ~w6401) | (w6056 & w47138) | (~w6401 & w47138);
assign w6431 = w6401 & w47139;
assign w6432 = ~w6430 & ~w6431;
assign w6433 = w3242 & w6432;
assign w6434 = (~w4056 & ~w6420) | (~w4056 & w40403) | (~w6420 & w40403);
assign w6435 = ~w6424 & w6434;
assign w6436 = w3646 & w6052;
assign w6437 = (w6436 & w6243) | (w6436 & w44240) | (w6243 & w44240);
assign w6438 = w3646 & w6412;
assign w6439 = ~w6243 & w44241;
assign w6440 = ~w6437 & ~w6439;
assign w6441 = ~w6435 & w6440;
assign w6442 = w6418 & ~w6441;
assign w6443 = ~w6433 & ~w6442;
assign w6444 = w5864 & w5891;
assign w6445 = (~w6056 & ~w6397) | (~w6056 & w40404) | (~w6397 & w40404);
assign w6446 = ~w6399 & ~w6445;
assign w6447 = w6444 & ~w6446;
assign w6448 = ~w6444 & w6446;
assign w6449 = ~w6447 & ~w6448;
assign w6450 = ~w3242 & w5864;
assign w6451 = w5891 & ~w6450;
assign w6452 = w6264 & ~w6449;
assign w6453 = (w6451 & w6243) | (w6451 & w52112) | (w6243 & w52112);
assign w6454 = ~w6452 & ~w6453;
assign w6455 = ~w6452 & w52113;
assign w6456 = ~w6442 & w44242;
assign w6457 = (w6456 & w6393) | (w6456 & w44243) | (w6393 & w44243);
assign w6458 = ~w6267 & w47140;
assign w6459 = w2006 & ~w6458;
assign w6460 = ~w2006 & w6458;
assign w6461 = ~w6459 & ~w6460;
assign w6462 = ~w1738 & ~w5933;
assign w6463 = (w6462 & ~w6264) | (w6462 & w44244) | (~w6264 & w44244);
assign w6464 = ~w1738 & w5933;
assign w6465 = w6264 & w44245;
assign w6466 = ~w6463 & ~w6465;
assign w6467 = (w6086 & w6060) | (w6086 & w49503) | (w6060 & w49503);
assign w6468 = (w2285 & w6261) | (w2285 & w48671) | (w6261 & w48671);
assign w6469 = ~w5833 & w49504;
assign w6470 = ~w6242 & w40405;
assign w6471 = ~w6468 & ~w6470;
assign w6472 = ~w6261 & w48672;
assign w6473 = ~w6243 & w6472;
assign w6474 = w6471 & ~w6473;
assign w6475 = w2006 & w6091;
assign w6476 = ~w6474 & w6475;
assign w6477 = w2006 & ~w6091;
assign w6478 = w6474 & w6477;
assign w6479 = ~w6476 & ~w6478;
assign w6480 = ~w5897 & w5915;
assign w6481 = (w6480 & w6049) | (w6480 & w51748) | (w6049 & w51748);
assign w6482 = ~w6261 & w48673;
assign w6483 = (w2558 & w6261) | (w2558 & w48674) | (w6261 & w48674);
assign w6484 = ~w5833 & w49505;
assign w6485 = ~w6242 & w40406;
assign w6486 = ~w6483 & ~w6485;
assign w6487 = ~w6243 & w6482;
assign w6488 = w6486 & ~w6487;
assign w6489 = w5911 & w6086;
assign w6490 = w2285 & w6489;
assign w6491 = ~w6488 & w6490;
assign w6492 = w2285 & ~w6489;
assign w6493 = w6488 & w6492;
assign w6494 = ~w6491 & ~w6493;
assign w6495 = w1738 & w5933;
assign w6496 = (w6495 & ~w6264) | (w6495 & w44246) | (~w6264 & w44246);
assign w6497 = w1738 & ~w5933;
assign w6498 = w6264 & w44247;
assign w6499 = ~w6496 & ~w6498;
assign w6500 = w6494 & w6499;
assign w6501 = w6466 & ~w6479;
assign w6502 = w6500 & ~w6501;
assign w6503 = ~w5934 & w5960;
assign w6504 = ~w6267 & w40407;
assign w6505 = w6098 & ~w6504;
assign w6506 = (~w1738 & w6261) | (~w1738 & w48675) | (w6261 & w48675);
assign w6507 = ~w5833 & w49506;
assign w6508 = ~w6242 & w40408;
assign w6509 = ~w6506 & ~w6508;
assign w6510 = ~w6261 & w51749;
assign w6511 = ~w6243 & w6510;
assign w6512 = w6509 & ~w6511;
assign w6513 = ~w5947 & w6103;
assign w6514 = w6103 & w51750;
assign w6515 = (w6514 & w6511) | (w6514 & w48676) | (w6511 & w48676);
assign w6516 = (w1541 & ~w6103) | (w1541 & w51751) | (~w6103 & w51751);
assign w6517 = ~w6511 & w48677;
assign w6518 = ~w6515 & ~w6517;
assign w6519 = w1320 & ~w6280;
assign w6520 = w6518 & ~w6519;
assign w6521 = w2896 & ~w6454;
assign w6522 = (w5891 & w6397) | (w5891 & w6057) | (w6397 & w6057);
assign w6523 = ~w6445 & w6522;
assign w6524 = w5864 & ~w6523;
assign w6525 = (~w2896 & w6261) | (~w2896 & w48678) | (w6261 & w48678);
assign w6526 = ~w5833 & w49507;
assign w6527 = ~w6242 & w40409;
assign w6528 = ~w6525 & ~w6527;
assign w6529 = w6263 & w6524;
assign w6530 = ~w6243 & w6529;
assign w6531 = w5873 & w5915;
assign w6532 = ~w6530 & w48679;
assign w6533 = (w6531 & w6530) | (w6531 & w48680) | (w6530 & w48680);
assign w6534 = ~w6532 & ~w6533;
assign w6535 = ~w2558 & ~w6534;
assign w6536 = (~w6521 & w6534) | (~w6521 & w40410) | (w6534 & w40410);
assign w6537 = w6502 & w40411;
assign w6538 = ~w6457 & w6537;
assign w6539 = ~w2006 & ~w6091;
assign w6540 = ~w6474 & w6539;
assign w6541 = ~w2006 & w6091;
assign w6542 = w6474 & w6541;
assign w6543 = ~w6540 & ~w6542;
assign w6544 = w6499 & ~w6543;
assign w6545 = (~w1541 & ~w6103) | (~w1541 & w51752) | (~w6103 & w51752);
assign w6546 = (w6545 & w6511) | (w6545 & w48681) | (w6511 & w48681);
assign w6547 = w6103 & w51753;
assign w6548 = ~w6511 & w48682;
assign w6549 = ~w6546 & ~w6548;
assign w6550 = w6466 & w6549;
assign w6551 = ~w6544 & w6550;
assign w6552 = w2558 & ~w6531;
assign w6553 = (w6552 & w6530) | (w6552 & w48683) | (w6530 & w48683);
assign w6554 = w2558 & w6531;
assign w6555 = ~w6530 & w48684;
assign w6556 = ~w6553 & ~w6555;
assign w6557 = ~w2285 & ~w6489;
assign w6558 = ~w6488 & w6557;
assign w6559 = ~w2285 & w6489;
assign w6560 = w6488 & w6559;
assign w6561 = ~w6558 & ~w6560;
assign w6562 = w6556 & w6561;
assign w6563 = w6520 & ~w6551;
assign w6564 = w6520 & ~w6562;
assign w6565 = w6502 & w6564;
assign w6566 = ~w6563 & ~w6565;
assign w6567 = w5976 & w6234;
assign w6568 = ~w6060 & w6567;
assign w6569 = ~w6112 & w40412;
assign w6570 = ~w6568 & ~w6569;
assign w6571 = (~w945 & w6568) | (~w945 & w40413) | (w6568 & w40413);
assign w6572 = w6263 & ~w6571;
assign w6573 = ~w6568 & w51754;
assign w6574 = w6263 & w51755;
assign w6575 = (w6211 & ~w6572) | (w6211 & w40414) | (~w6572 & w40414);
assign w6576 = ~w6211 & ~w6243;
assign w6577 = w6574 & w6576;
assign w6578 = ~w6575 & ~w6577;
assign w6579 = (~w754 & w6577) | (~w754 & w40415) | (w6577 & w40415);
assign w6580 = (w6261 & w50276) | (w6261 & w50277) | (w50276 & w50277);
assign w6581 = (w5974 & w6093) | (w5974 & w40417) | (w6093 & w40417);
assign w6582 = ~w6075 & ~w6581;
assign w6583 = ~w6061 & w6582;
assign w6584 = ~w6580 & ~w6583;
assign w6585 = w6114 & w6234;
assign w6586 = w6073 & w6243;
assign w6587 = (w6073 & w6261) | (w6073 & w48685) | (w6261 & w48685);
assign w6588 = w6263 & w6585;
assign w6589 = ~w6587 & ~w6588;
assign w6590 = ~w6586 & w6589;
assign w6591 = w6589 & w51756;
assign w6592 = w6589 & w50278;
assign w6593 = ~w6579 & ~w6592;
assign w6594 = ~w1320 & w6280;
assign w6595 = ~w5973 & ~w6075;
assign w6596 = (~w1320 & w6261) | (~w1320 & w48686) | (w6261 & w48686);
assign w6597 = ~w5833 & w50279;
assign w6598 = ~w6242 & w40419;
assign w6599 = ~w6596 & ~w6598;
assign w6600 = ~w6261 & w50280;
assign w6601 = ~w6243 & w6600;
assign w6602 = w6599 & ~w6601;
assign w6603 = w6595 & ~w6602;
assign w6604 = ~w6595 & w6602;
assign w6605 = ~w6603 & ~w6604;
assign w6606 = w1120 & w6605;
assign w6607 = (~w6594 & ~w6605) | (~w6594 & w47141) | (~w6605 & w47141);
assign w6608 = ~w6594 & w52198;
assign w6609 = w6566 & w6608;
assign w6610 = w5853 & w6254;
assign w6611 = ~w6284 & ~w6610;
assign w6612 = ~w6286 & w51758;
assign w6613 = ~w6285 & w6612;
assign w6614 = (~w6610 & w6286) | (~w6610 & w51759) | (w6286 & w51759);
assign w6615 = (~w6614 & ~w6611) | (~w6614 & w51760) | (~w6611 & w51760);
assign w6616 = ~w6613 & w6615;
assign w6617 = ~w5847 & w51761;
assign w6618 = (w5848 & w5847) | (w5848 & w51762) | (w5847 & w51762);
assign w6619 = ~w6617 & ~w6618;
assign w6620 = w6264 & w6616;
assign w6621 = ~w6264 & ~w6619;
assign w6622 = ~w6620 & ~w6621;
assign w6623 = (~w57 & w6620) | (~w57 & w40420) | (w6620 & w40420);
assign w6624 = w5817 & ~w6171;
assign w6625 = w5805 & ~w6624;
assign w6626 = ~w6239 & w40421;
assign w6627 = (w6625 & ~w6626) | (w6625 & w51763) | (~w6626 & w51763);
assign w6628 = ~w6228 & w6625;
assign w6629 = ~w6113 & w6628;
assign w6630 = (~w6627 & ~w6629) | (~w6627 & w51764) | (~w6629 & w51764);
assign w6631 = w6263 & ~w6630;
assign w6632 = (~w351 & w6261) | (~w351 & w48687) | (w6261 & w48687);
assign w6633 = ~w5833 & w49508;
assign w6634 = ~w6242 & w40422;
assign w6635 = ~w6632 & ~w6634;
assign w6636 = ~w6243 & w6631;
assign w6637 = w5790 & ~w5808;
assign w6638 = ~w252 & w6637;
assign w6639 = (w6638 & w6636) | (w6638 & w48688) | (w6636 & w48688);
assign w6640 = ~w252 & ~w6637;
assign w6641 = ~w6636 & w48689;
assign w6642 = ~w6639 & ~w6641;
assign w6643 = ~w6623 & w6642;
assign w6644 = ~w6620 & w40423;
assign w6645 = ~w6286 & w51765;
assign w6646 = ~w6285 & w6645;
assign w6647 = (w6254 & w6285) | (w6254 & w47142) | (w6285 & w47142);
assign w6648 = ~w5843 & ~w5844;
assign w6649 = ~w6261 & w48690;
assign w6650 = ~w6243 & w6649;
assign w6651 = ~w6647 & w6650;
assign w6652 = (w5842 & w6243) | (w5842 & w52114) | (w6243 & w52114);
assign w6653 = ~w6651 & ~w6652;
assign w6654 = ~w6261 & w49509;
assign w6655 = ~w6243 & w6654;
assign w6656 = w6647 & w6655;
assign w6657 = (~w80 & ~w6655) | (~w80 & w40424) | (~w6655 & w40424);
assign w6658 = w6653 & w6657;
assign w6659 = ~w6644 & ~w6658;
assign w6660 = w252 & ~w6637;
assign w6661 = (w6660 & w6636) | (w6660 & w48691) | (w6636 & w48691);
assign w6662 = w252 & w6637;
assign w6663 = ~w6636 & w48692;
assign w6664 = ~w6661 & ~w6663;
assign w6665 = ~w400 & w5805;
assign w6666 = w5817 & ~w6665;
assign w6667 = (~w351 & w6665) | (~w351 & w51766) | (w6665 & w51766);
assign w6668 = ~w6261 & w49510;
assign w6669 = (~w6667 & ~w6668) | (~w6667 & w40425) | (~w6668 & w40425);
assign w6670 = w5805 & w5817;
assign w6671 = w6076 & w6171;
assign w6672 = ~w6228 & w6671;
assign w6673 = ~w6581 & w6672;
assign w6674 = w6171 & ~w6626;
assign w6675 = w6670 & w52199;
assign w6676 = ~w6670 & ~w52199;
assign w6677 = ~w6675 & ~w6676;
assign w6678 = w6264 & ~w6677;
assign w6679 = ~w6669 & ~w6678;
assign w6680 = w6664 & ~w6679;
assign w6681 = w6643 & ~w6680;
assign w6682 = w6659 & ~w6681;
assign w6683 = w5831 & w6171;
assign w6684 = w6336 & ~w6683;
assign w6685 = ~w6179 & ~w6198;
assign w6686 = w6226 & w6685;
assign w6687 = w6240 & w6686;
assign w6688 = (w6683 & w6239) | (w6683 & w51767) | (w6239 & w51767);
assign w6689 = ~w6239 & w51768;
assign w6690 = ~w6688 & ~w6689;
assign w6691 = (w6690 & ~w44248) | (w6690 & w51769) | (~w44248 & w51769);
assign w6692 = w5646 & ~w5826;
assign w6693 = ~w5646 & w5826;
assign w6694 = ~w6692 & ~w6693;
assign w6695 = (~w6694 & w6243) | (~w6694 & w44249) | (w6243 & w44249);
assign w6696 = ~w6684 & ~w6691;
assign w6697 = w6264 & w6696;
assign w6698 = ~w6695 & ~w6697;
assign w6699 = ~w6697 & w44250;
assign w6700 = w5917 & w44251;
assign w6701 = ~w6060 & w6700;
assign w6702 = (w6237 & w5974) | (w6237 & w44252) | (w5974 & w44252);
assign w6703 = (w6226 & w6112) | (w6226 & w40426) | (w6112 & w40426);
assign w6704 = ~w6685 & w52200;
assign w6705 = w6240 & w6685;
assign w6706 = ~w6336 & w6705;
assign w6707 = ~w6704 & ~w6706;
assign w6708 = (w6178 & w6243) | (w6178 & w44253) | (w6243 & w44253);
assign w6709 = w6264 & ~w6707;
assign w6710 = ~w6708 & ~w6709;
assign w6711 = (~w493 & w6709) | (~w493 & w44254) | (w6709 & w44254);
assign w6712 = ~w6699 & ~w6711;
assign w6713 = (~w400 & w6697) | (~w400 & w49511) | (w6697 & w49511);
assign w6714 = (w6666 & w6243) | (w6666 & w52115) | (w6243 & w52115);
assign w6715 = ~w6678 & ~w6714;
assign w6716 = (w351 & w6678) | (w351 & w52116) | (w6678 & w52116);
assign w6717 = ~w6713 & ~w6716;
assign w6718 = ~w6712 & w6717;
assign w6719 = w6643 & w6718;
assign w6720 = w6682 & ~w6719;
assign w6721 = ~w5721 & w51770;
assign w6722 = (w6185 & w5721) | (w6185 & w51771) | (w5721 & w51771);
assign w6723 = ~w6721 & ~w6722;
assign w6724 = w6180 & w6723;
assign w6725 = ~w6180 & ~w6723;
assign w6726 = ~w6724 & ~w6725;
assign w6727 = w6197 & w6225;
assign w6728 = ~w6701 & w40429;
assign w6729 = (w6727 & w6701) | (w6727 & w40430) | (w6701 & w40430);
assign w6730 = ~w6728 & ~w6729;
assign w6731 = ~w612 & ~w6726;
assign w6732 = (w6731 & w6243) | (w6731 & w52117) | (w6243 & w52117);
assign w6733 = ~w612 & ~w6730;
assign w6734 = w6264 & w6733;
assign w6735 = ~w6732 & ~w6734;
assign w6736 = w6682 & w40431;
assign w6737 = w6609 & w47144;
assign w6738 = ~w6577 & w48693;
assign w6739 = (~w945 & ~w6590) | (~w945 & w40432) | (~w6590 & w40432);
assign w6740 = ~w1120 & w6595;
assign w6741 = (w6740 & w6601) | (w6740 & w48694) | (w6601 & w48694);
assign w6742 = ~w1120 & ~w6595;
assign w6743 = ~w6601 & w48695;
assign w6744 = ~w6741 & ~w6743;
assign w6745 = ~w6739 & w6744;
assign w6746 = (~w6738 & w6745) | (~w6738 & w40433) | (w6745 & w40433);
assign w6747 = ~w6679 & w6735;
assign w6748 = w6664 & w6747;
assign w6749 = w6659 & w6748;
assign w6750 = ~w6718 & w6749;
assign w6751 = ~w6746 & w6750;
assign w6752 = (w6726 & w6243) | (w6726 & w44255) | (w6243 & w44255);
assign w6753 = ~w6243 & w44256;
assign w6754 = ~w6752 & ~w6753;
assign w6755 = (w612 & w6753) | (w612 & w49512) | (w6753 & w49512);
assign w6756 = ~w6709 & w44257;
assign w6757 = ~w6755 & ~w6756;
assign w6758 = w6712 & ~w6757;
assign w6759 = w6643 & w6717;
assign w6760 = ~w6758 & w6759;
assign w6761 = w6682 & ~w6760;
assign w6762 = ~w6751 & ~w6761;
assign w6763 = w6653 & ~w6656;
assign w6764 = (w80 & ~w6653) | (w80 & w51772) | (~w6653 & w51772);
assign w6765 = ~w3 & w6315;
assign w6766 = ~w6309 & ~w6765;
assign w6767 = ~w6765 & w49513;
assign w6768 = w6762 & w6767;
assign w6769 = (w6318 & w6737) | (w6318 & w40434) | (w6737 & w40434);
assign w6770 = w6479 & w6500;
assign w6771 = w6518 & ~w6551;
assign w6772 = w6518 & ~w6562;
assign w6773 = w6770 & w6772;
assign w6774 = ~w6771 & ~w6773;
assign w6775 = w6770 & w40435;
assign w6776 = ~w6457 & w6775;
assign w6777 = ~w6519 & ~w6594;
assign w6778 = ~w1120 & w6777;
assign w6779 = (w6778 & w6776) | (w6778 & w48696) | (w6776 & w48696);
assign w6780 = ~w1120 & ~w6777;
assign w6781 = ~w6776 & w48697;
assign w6782 = ~w6779 & ~w6781;
assign w6783 = ~w6769 & ~w6782;
assign w6784 = ~w1120 & ~w6280;
assign w6785 = (w6737 & w48698) | (w6737 & w48699) | (w48698 & w48699);
assign w6786 = ~w6783 & ~w6785;
assign w6787 = w1120 & ~w6777;
assign w6788 = (w6787 & w6776) | (w6787 & w48700) | (w6776 & w48700);
assign w6789 = w1120 & w6777;
assign w6790 = ~w6776 & w48701;
assign w6791 = ~w6788 & ~w6790;
assign w6792 = ~w6769 & ~w6791;
assign w6793 = w1120 & w6280;
assign w6794 = (w6737 & w48702) | (w6737 & w48703) | (w48702 & w48703);
assign w6795 = ~w6792 & ~w6794;
assign w6796 = w6786 & w6795;
assign w6797 = w6512 & ~w6513;
assign w6798 = ~w6512 & w6513;
assign w6799 = ~w6797 & ~w6798;
assign w6800 = ~w6456 & w6536;
assign w6801 = w6429 & w6536;
assign w6802 = ~w6393 & w6801;
assign w6803 = ~w6800 & ~w6802;
assign w6804 = ~w6802 & w44258;
assign w6805 = (w6466 & w6543) | (w6466 & w40436) | (w6543 & w40436);
assign w6806 = w6770 & w6805;
assign w6807 = w6518 & w6549;
assign w6808 = w6805 & ~w6807;
assign w6809 = ~w6805 & w6807;
assign w6810 = ~w6808 & ~w6809;
assign w6811 = ~w6806 & ~w6810;
assign w6812 = w6562 & ~w6810;
assign w6813 = (~w6811 & ~w6803) | (~w6811 & w44259) | (~w6803 & w44259);
assign w6814 = w6770 & w51773;
assign w6815 = (w6814 & w6802) | (w6814 & w51774) | (w6802 & w51774);
assign w6816 = w6813 & ~w6815;
assign w6817 = ~w1320 & w6799;
assign w6818 = (w6737 & w48704) | (w6737 & w48705) | (w48704 & w48705);
assign w6819 = w6813 & w47145;
assign w6820 = ~w6769 & w6819;
assign w6821 = ~w6818 & ~w6820;
assign w6822 = (w6319 & w6317) | (w6319 & w49514) | (w6317 & w49514);
assign w6823 = (~w6822 & w6737) | (~w6822 & w40438) | (w6737 & w40438);
assign w6824 = ~w6317 & w51775;
assign w6825 = (w6824 & w6737) | (w6824 & w40439) | (w6737 & w40439);
assign w6826 = w6823 & ~w6825;
assign w6827 = ~a[71] & ~a[72];
assign w6828 = ~a[70] & w6827;
assign w6829 = w6264 & w6828;
assign w6830 = ~w6826 & ~w6829;
assign w6831 = ~w6264 & ~w6828;
assign w6832 = ~w6317 & w51776;
assign w6833 = (w6832 & w6737) | (w6832 & w40440) | (w6737 & w40440);
assign w6834 = ~w6264 & w7547;
assign w6835 = (~w40440 & w47146) | (~w40440 & w47147) | (w47146 & w47147);
assign w6836 = (w6835 & w6826) | (w6835 & w47148) | (w6826 & w47148);
assign w6837 = w5745 & ~w6836;
assign w6838 = ~w5745 & w6835;
assign w6839 = ~w6830 & w6838;
assign w6840 = ~w6317 & w49515;
assign w6841 = (w6840 & w6737) | (w6840 & w40441) | (w6737 & w40441);
assign w6842 = w6823 & ~w6841;
assign w6843 = a[74] & ~w6842;
assign w6844 = ~a[74] & w6842;
assign w6845 = ~w6843 & ~w6844;
assign w6846 = ~w6839 & w6845;
assign w6847 = ~w6837 & ~w6846;
assign w6848 = ~w6321 & ~w6345;
assign w6849 = w6264 & ~w6848;
assign w6850 = ~w6264 & w6848;
assign w6851 = ~w6849 & ~w6850;
assign w6852 = ~w6851 & ~w6769;
assign w6853 = ~a[74] & w6840;
assign w6854 = ~w5328 & w51777;
assign w6855 = (~w40442 & w47149) | (~w40442 & w47150) | (w47149 & w47150);
assign w6856 = ~w6852 & w6855;
assign w6857 = ~w5328 & w51778;
assign w6858 = (w47151 & w50281) | (w47151 & w40442) | (w50281 & w40442);
assign w6859 = ~w6851 & w6857;
assign w6860 = w6859 & ~w6769;
assign w6861 = ~w6858 & ~w6860;
assign w6862 = ~w6856 & w6861;
assign w6863 = ~w6346 & ~w6349;
assign w6864 = ~w6317 & w49516;
assign w6865 = w6358 & ~w6863;
assign w6866 = ~w6358 & w6863;
assign w6867 = ~w6865 & ~w6866;
assign w6868 = ~w6864 & w6867;
assign w6869 = w6762 & w40443;
assign w6870 = (~w6868 & w6737) | (~w6868 & w40444) | (w6737 & w40444);
assign w6871 = ~w6358 & w6864;
assign w6872 = (w6871 & w6737) | (w6871 & w40445) | (w6737 & w40445);
assign w6873 = w6870 & ~w6872;
assign w6874 = ~w4838 & ~w6873;
assign w6875 = ~w6359 & w51779;
assign w6876 = (w4838 & w6359) | (w4838 & w51780) | (w6359 & w51780);
assign w6877 = ~w6875 & ~w6876;
assign w6878 = (~w6877 & w6317) | (~w6877 & w51781) | (w6317 & w51781);
assign w6879 = w6762 & w40446;
assign w6880 = (w4430 & w6389) | (w4430 & w51782) | (w6389 & w51782);
assign w6881 = (~w40447 & w47152) | (~w40447 & w47153) | (w47152 & w47153);
assign w6882 = ~w6389 & w51783;
assign w6883 = ~w6878 & w6882;
assign w6884 = (w6883 & w6737) | (w6883 & w40448) | (w6737 & w40448);
assign w6885 = ~w6881 & ~w6884;
assign w6886 = ~w6874 & w6885;
assign w6887 = w6862 & w6886;
assign w6888 = ~w6847 & w6887;
assign w6889 = ~a[75] & ~w6851;
assign w6890 = w6889 & ~w6769;
assign w6891 = (~w40442 & w47154) | (~w40442 & w47155) | (w47154 & w47155);
assign w6892 = ~w6852 & w6891;
assign w6893 = (w47156 & w50282) | (w47156 & w40442) | (w50282 & w40442);
assign w6894 = ~w6890 & ~w6893;
assign w6895 = ~w6892 & w6894;
assign w6896 = (~w40448 & w47157) | (~w40448 & w47158) | (w47157 & w47158);
assign w6897 = ~w6881 & w6896;
assign w6898 = ~w6874 & w6897;
assign w6899 = (~w40447 & w47159) | (~w40447 & w47160) | (w47159 & w47160);
assign w6900 = (w47161 & w50283) | (w47161 & w40447) | (w50283 & w40447);
assign w6901 = ~w6899 & ~w6900;
assign w6902 = ~w4430 & ~w6901;
assign w6903 = w4838 & w6873;
assign w6904 = w6885 & w6903;
assign w6905 = ~w6902 & ~w6904;
assign w6906 = ~w6895 & w6898;
assign w6907 = w6905 & ~w6906;
assign w6908 = ~w6392 & ~w6427;
assign w6909 = w6376 & ~w6427;
assign w6910 = w6360 & w6909;
assign w6911 = ~w6908 & ~w6910;
assign w6912 = w6425 & ~w6911;
assign w6913 = ~w6911 & w51784;
assign w6914 = ~w6913 & ~w6769;
assign w6915 = (w3646 & w6424) | (w3646 & w51785) | (w6424 & w51785);
assign w6916 = w6427 & ~w6915;
assign w6917 = ~w6377 & w51786;
assign w6918 = (~w6391 & ~w40396) | (~w6391 & w51787) | (~w40396 & w51787);
assign w6919 = ~w6383 & ~w6427;
assign w6920 = ~w6918 & ~w6919;
assign w6921 = ~w6917 & ~w6920;
assign w6922 = ~w6424 & w51788;
assign w6923 = ~w4430 & ~w6922;
assign w6924 = ~w6918 & w6923;
assign w6925 = w6921 & ~w6924;
assign w6926 = w6912 & ~w6925;
assign w6927 = ~w6425 & w6911;
assign w6928 = (~w3646 & ~w6911) | (~w3646 & w51789) | (~w6911 & w51789);
assign w6929 = ~w6921 & ~w6928;
assign w6930 = w6929 & ~w6769;
assign w6931 = ~w6926 & ~w6930;
assign w6932 = ~w6382 & ~w6914;
assign w6933 = w6931 & ~w6932;
assign w6934 = (w6737 & w48706) | (w6737 & w48707) | (w48706 & w48707);
assign w6935 = w3646 & ~w6934;
assign w6936 = ~w6912 & ~w6927;
assign w6937 = w4056 & w6936;
assign w6938 = ~w6937 & ~w6769;
assign w6939 = ~w4056 & ~w6933;
assign w6940 = w6935 & ~w6938;
assign w6941 = ~w6939 & ~w6940;
assign w6942 = w6907 & w6941;
assign w6943 = ~w6888 & w6942;
assign w6944 = w4430 & ~w6918;
assign w6945 = ~w4430 & w6918;
assign w6946 = ~w6944 & ~w6945;
assign w6947 = ~w6946 & ~w6769;
assign w6948 = ~w6936 & w51790;
assign w6949 = ~w6911 & ~w6915;
assign w6950 = ~w6924 & w6949;
assign w6951 = ~w6948 & ~w6950;
assign w6952 = w6911 & w51791;
assign w6953 = (~w6952 & w6769) | (~w6952 & w51792) | (w6769 & w51792);
assign w6954 = w6382 & ~w6947;
assign w6955 = ~w6935 & w6954;
assign w6956 = w6936 & w6938;
assign w6957 = ~w6934 & ~w6956;
assign w6958 = (w4056 & w6955) | (w4056 & w51793) | (w6955 & w51793);
assign w6959 = ~w3646 & ~w6957;
assign w6960 = ~w6958 & ~w6959;
assign w6961 = w6406 & ~w6433;
assign w6962 = (~w6426 & w6910) | (~w6426 & w40449) | (w6910 & w40449);
assign w6963 = w6417 & w52201;
assign w6964 = w6961 & ~w6963;
assign w6965 = ~w6961 & w6963;
assign w6966 = ~w6964 & ~w6965;
assign w6967 = w2896 & w6966;
assign w6968 = ~w6769 & w6967;
assign w6969 = ~w6317 & w49517;
assign w6970 = (w6969 & w6737) | (w6969 & w40450) | (w6737 & w40450);
assign w6971 = (w40450 & w47164) | (w40450 & w47165) | (w47164 & w47165);
assign w6972 = ~w6968 & ~w6971;
assign w6973 = w6417 & w6440;
assign w6974 = (w6973 & w6962) | (w6973 & w51794) | (w6962 & w51794);
assign w6975 = ~w6962 & w51795;
assign w6976 = ~w6974 & ~w6975;
assign w6977 = w6052 & ~w6264;
assign w6978 = w6264 & w6412;
assign w6979 = ~w6977 & ~w6978;
assign w6980 = w6976 & ~w6769;
assign w6981 = (w6737 & w51796) | (w6737 & w51797) | (w51796 & w51797);
assign w6982 = ~w6980 & ~w6981;
assign w6983 = ~w3242 & w6982;
assign w6984 = w6972 & ~w6983;
assign w6985 = w6960 & w6984;
assign w6986 = ~w6943 & w6985;
assign w6987 = w6091 & ~w6474;
assign w6988 = ~w6091 & w6474;
assign w6989 = ~w6987 & ~w6988;
assign w6990 = w6479 & w6543;
assign w6991 = (w6494 & w6802) | (w6494 & w48708) | (w6802 & w48708);
assign w6992 = w6990 & ~w6991;
assign w6993 = ~w6990 & w6991;
assign w6994 = ~w6992 & ~w6993;
assign w6995 = (w6737 & w48709) | (w6737 & w48710) | (w48709 & w48710);
assign w6996 = ~w6769 & w6994;
assign w6997 = ~w6995 & ~w6996;
assign w6998 = ~w6996 & w48711;
assign w6999 = (w5933 & ~w6264) | (w5933 & w51798) | (~w6264 & w51798);
assign w7000 = w6264 & w51799;
assign w7001 = ~w6999 & ~w7000;
assign w7002 = w6466 & w6499;
assign w7003 = w6479 & w6494;
assign w7004 = (w7003 & w6802) | (w7003 & w48712) | (w6802 & w48712);
assign w7005 = (w7002 & w7004) | (w7002 & w49518) | (w7004 & w49518);
assign w7006 = ~w7004 & w49519;
assign w7007 = (w6737 & w49999) | (w6737 & w50000) | (w49999 & w50000);
assign w7008 = ~w6769 & w48713;
assign w7009 = ~w7007 & ~w7008;
assign w7010 = (~w1541 & w7008) | (~w1541 & w50001) | (w7008 & w50001);
assign w7011 = ~w6998 & ~w7010;
assign w7012 = (w6443 & w6393) | (w6443 & w44260) | (w6393 & w44260);
assign w7013 = ~w6318 & w7012;
assign w7014 = (~w7013 & w6737) | (~w7013 & w40452) | (w6737 & w40452);
assign w7015 = ~w6970 & w7014;
assign w7016 = ~w6455 & ~w6521;
assign w7017 = ~w2558 & ~w7016;
assign w7018 = ~w7015 & w7017;
assign w7019 = ~w2558 & w7016;
assign w7020 = w7015 & w7019;
assign w7021 = ~w7018 & ~w7020;
assign w7022 = ~w6535 & w6556;
assign w7023 = (w7022 & w6457) | (w7022 & w48714) | (w6457 & w48714);
assign w7024 = ~w6457 & w48715;
assign w7025 = ~w7023 & ~w7024;
assign w7026 = w2285 & ~w6534;
assign w7027 = (w6737 & w49520) | (w6737 & w49521) | (w49520 & w49521);
assign w7028 = w2285 & w7025;
assign w7029 = ~w6769 & w7028;
assign w7030 = ~w7027 & ~w7029;
assign w7031 = w7021 & w7030;
assign w7032 = (w2558 & w7015) | (w2558 & w47166) | (w7015 & w47166);
assign w7033 = w7015 & w7016;
assign w7034 = w7032 & ~w7033;
assign w7035 = ~w2285 & w6534;
assign w7036 = (w6737 & w48716) | (w6737 & w48717) | (w48716 & w48717);
assign w7037 = ~w2285 & ~w7025;
assign w7038 = ~w6769 & w7037;
assign w7039 = ~w7036 & ~w7038;
assign w7040 = w6494 & w6561;
assign w7041 = ~w6802 & w48718;
assign w7042 = (w7040 & w6802) | (w7040 & w48719) | (w6802 & w48719);
assign w7043 = ~w7041 & ~w7042;
assign w7044 = w6488 & ~w6489;
assign w7045 = ~w6488 & w6489;
assign w7046 = ~w7044 & ~w7045;
assign w7047 = ~w2006 & w7043;
assign w7048 = ~w6769 & w7047;
assign w7049 = ~w2006 & w7046;
assign w7050 = (w6737 & w44262) | (w6737 & w44263) | (w44262 & w44263);
assign w7051 = ~w7048 & ~w7050;
assign w7052 = w7039 & w7051;
assign w7053 = (w6737 & w44264) | (w6737 & w44265) | (w44264 & w44265);
assign w7054 = w6966 & ~w6769;
assign w7055 = ~w7053 & ~w7054;
assign w7056 = w3242 & w6976;
assign w7057 = w7056 & ~w6769;
assign w7058 = w3242 & ~w6979;
assign w7059 = (w6737 & w44266) | (w6737 & w44267) | (w44266 & w44267);
assign w7060 = ~w7057 & ~w7059;
assign w7061 = ~w7054 & w44268;
assign w7062 = w6972 & ~w7060;
assign w7063 = ~w7061 & ~w7062;
assign w7064 = w7052 & w7063;
assign w7065 = w7031 & w7034;
assign w7066 = w7064 & ~w7065;
assign w7067 = ~w7065 & w47167;
assign w7068 = (w7067 & w6943) | (w7067 & w47168) | (w6943 & w47168);
assign w7069 = ~w7008 & w44269;
assign w7070 = w2006 & ~w7043;
assign w7071 = ~w6769 & w7070;
assign w7072 = w2006 & ~w7046;
assign w7073 = (w6737 & w44270) | (w6737 & w44271) | (w44270 & w44271);
assign w7074 = ~w7071 & ~w7073;
assign w7075 = ~w7052 & w7074;
assign w7076 = w7030 & w7074;
assign w7077 = w7021 & w7076;
assign w7078 = ~w7075 & ~w7077;
assign w7079 = (w1738 & w6996) | (w1738 & w48720) | (w6996 & w48720);
assign w7080 = (~w7069 & w7010) | (~w7069 & w44272) | (w7010 & w44272);
assign w7081 = ~w7069 & ~w7079;
assign w7082 = (~w47169 & w48721) | (~w47169 & w48722) | (w48721 & w48722);
assign w7083 = (w6737 & w49522) | (w6737 & w49523) | (w49522 & w49523);
assign w7084 = ~w6769 & w6816;
assign w7085 = ~w7083 & ~w7084;
assign w7086 = ~w7084 & w49524;
assign w7087 = ~w7082 & ~w7086;
assign w7088 = w6566 & ~w6594;
assign w7089 = ~w6538 & w7088;
assign w7090 = ~w6606 & w6744;
assign w7091 = ~w6606 & w51800;
assign w7092 = (w7091 & ~w7088) | (w7091 & w47170) | (~w7088 & w47170);
assign w7093 = (~w945 & w6606) | (~w945 & w51801) | (w6606 & w51801);
assign w7094 = w7088 & w47171;
assign w7095 = ~w7092 & ~w7094;
assign w7096 = ~w6769 & ~w7095;
assign w7097 = ~w945 & ~w6605;
assign w7098 = (w6737 & w44274) | (w6737 & w44275) | (w44274 & w44275);
assign w7099 = ~w7096 & ~w7098;
assign w7100 = w6786 & w7099;
assign w7101 = ~w7086 & w7100;
assign w7102 = ~w6519 & w6744;
assign w7103 = ~w6606 & ~w7102;
assign w7104 = (~w7103 & ~w6774) | (~w7103 & w40453) | (~w6774 & w40453);
assign w7105 = w6775 & ~w7103;
assign w7106 = ~w6457 & w7105;
assign w7107 = ~w7104 & ~w7106;
assign w7108 = ~w6592 & ~w6739;
assign w7109 = ~w7107 & w7108;
assign w7110 = w7107 & ~w7108;
assign w7111 = (w6737 & w44276) | (w6737 & w44277) | (w44276 & w44277);
assign w7112 = ~w7109 & ~w7110;
assign w7113 = ~w6769 & w7112;
assign w7114 = ~w7111 & ~w7113;
assign w7115 = ~w7113 & w44278;
assign w7116 = ~w6579 & ~w6738;
assign w7117 = w7116 & w52202;
assign w7118 = ~w6592 & ~w7116;
assign w7119 = (w7118 & w7107) | (w7118 & w44280) | (w7107 & w44280);
assign w7120 = ~w6769 & w51802;
assign w7121 = (w6737 & w44281) | (w6737 & w44282) | (w44281 & w44282);
assign w7122 = w612 & ~w7121;
assign w7123 = ~w7120 & w7122;
assign w7124 = ~w7115 & ~w7123;
assign w7125 = (w6746 & ~w6566) | (w6746 & w40454) | (~w6566 & w40454);
assign w7126 = w6537 & w6746;
assign w7127 = ~w6457 & w7126;
assign w7128 = ~w7125 & ~w7127;
assign w7129 = w612 & ~w7128;
assign w7130 = ~w612 & w7128;
assign w7131 = ~w7129 & ~w7130;
assign w7132 = (w6754 & w7131) | (w6754 & w47172) | (w7131 & w47172);
assign w7133 = ~w7131 & w47173;
assign w7134 = ~w7132 & ~w7133;
assign w7135 = ~w7133 & w50284;
assign w7136 = w7124 & ~w7135;
assign w7137 = w7101 & w7136;
assign w7138 = ~w7082 & w7137;
assign w7139 = (~w47168 & w48723) | (~w47168 & w48724) | (w48723 & w48724);
assign w7140 = ~w6317 & w48725;
assign w7141 = (w7140 & w6737) | (w7140 & w40455) | (w6737 & w40455);
assign w7142 = w6717 & ~w6758;
assign w7143 = (w6680 & w6758) | (w6680 & w48726) | (w6758 & w48726);
assign w7144 = ~w6718 & w6748;
assign w7145 = ~w7143 & ~w7144;
assign w7146 = w6609 & ~w7145;
assign w7147 = w6609 & w47174;
assign w7148 = (w6642 & w7142) | (w6642 & w44283) | (w7142 & w44283);
assign w7149 = ~w6746 & w7144;
assign w7150 = w7148 & ~w7149;
assign w7151 = ~w6623 & ~w6644;
assign w7152 = (~w7146 & w47175) | (~w7146 & w47176) | (w47175 & w47176);
assign w7153 = ~w6720 & w6767;
assign w7154 = ~w6658 & w51803;
assign w7155 = ~w6317 & w51804;
assign w7156 = (w7128 & w51805) | (w7128 & w51806) | (w51805 & w51806);
assign w7157 = (~w7156 & w7141) | (~w7156 & w52124) | (w7141 & w52124);
assign w7158 = (w7146 & w47177) | (w7146 & w47178) | (w47177 & w47178);
assign w7159 = ~w6769 & w7158;
assign w7160 = ~w7157 & ~w7159;
assign w7161 = (~w80 & w7157) | (~w80 & w51807) | (w7157 & w51807);
assign w7162 = (w6737 & w44284) | (w6737 & w44285) | (w44284 & w44285);
assign w7163 = ~w6758 & w51808;
assign w7164 = w6712 & w6735;
assign w7165 = (~w6715 & w6758) | (~w6715 & w51809) | (w6758 & w51809);
assign w7166 = w6712 & w51810;
assign w7167 = (~w7165 & ~w7128) | (~w7165 & w44286) | (~w7128 & w44286);
assign w7168 = (w351 & w6758) | (w351 & w51811) | (w6758 & w51811);
assign w7169 = w351 & w7164;
assign w7170 = (~w7168 & ~w7128) | (~w7168 & w44287) | (~w7128 & w44287);
assign w7171 = ~w6769 & w7170;
assign w7172 = ~w6769 & w44288;
assign w7173 = w6642 & w6664;
assign w7174 = w57 & ~w7173;
assign w7175 = (w7174 & w7172) | (w7174 & w51812) | (w7172 & w51812);
assign w7176 = w57 & w7173;
assign w7177 = ~w7172 & w51813;
assign w7178 = ~w7175 & ~w7177;
assign w7179 = ~w7161 & w7178;
assign w7180 = ~w6755 & w6746;
assign w7181 = (w7180 & ~w6566) | (w7180 & w40456) | (~w6566 & w40456);
assign w7182 = w6537 & w7180;
assign w7183 = ~w6457 & w7182;
assign w7184 = ~w7181 & ~w7183;
assign w7185 = w6735 & w7184;
assign w7186 = ~w6699 & ~w6713;
assign w7187 = ~w6756 & ~w7186;
assign w7188 = (w7187 & ~w7184) | (w7187 & w51814) | (~w7184 & w51814);
assign w7189 = ~w6713 & w7164;
assign w7190 = w6756 & w7186;
assign w7191 = (~w7190 & ~w7184) | (~w7190 & w44290) | (~w7184 & w44290);
assign w7192 = (w6737 & w49525) | (w6737 & w49526) | (w49525 & w49526);
assign w7193 = ~w6769 & w51815;
assign w7194 = ~w7192 & ~w7193;
assign w7195 = ~w7193 & w44291;
assign w7196 = w7128 & w7164;
assign w7197 = w252 & w6715;
assign w7198 = (w7197 & ~w7171) | (w7197 & w44292) | (~w7171 & w44292);
assign w7199 = w252 & ~w6715;
assign w7200 = w7171 & w44293;
assign w7201 = ~w7198 & ~w7200;
assign w7202 = ~w7195 & w7201;
assign w7203 = ~w57 & ~w7173;
assign w7204 = ~w7162 & w7203;
assign w7205 = ~w7172 & w7204;
assign w7206 = ~w57 & w7173;
assign w7207 = w7162 & w7206;
assign w7208 = w7206 & w7167;
assign w7209 = ~w6769 & w51816;
assign w7210 = ~w7207 & ~w7209;
assign w7211 = ~w7205 & w7210;
assign w7212 = ~w252 & ~w6715;
assign w7213 = (w7212 & ~w7171) | (w7212 & w44294) | (~w7171 & w44294);
assign w7214 = ~w252 & w6715;
assign w7215 = w7171 & w44295;
assign w7216 = ~w7213 & ~w7215;
assign w7217 = w7211 & w7216;
assign w7218 = ~w7202 & w7217;
assign w7219 = (w80 & w6769) | (w80 & w52125) | (w6769 & w52125);
assign w7220 = ~w7157 & w7219;
assign w7221 = ~w7149 & w44296;
assign w7222 = w80 & ~w6644;
assign w7223 = ~w80 & w6644;
assign w7224 = ~w7222 & ~w7223;
assign w7225 = (w40457 & ~w47174) | (w40457 & w52118) | (~w47174 & w52118);
assign w7226 = (w47174 & w52119) | (w47174 & w52120) | (w52119 & w52120);
assign w7227 = ~w7225 & ~w7226;
assign w7228 = ~w6765 & w51817;
assign w7229 = w6318 & ~w7228;
assign w7230 = (w7229 & w6737) | (w7229 & w40459) | (w6737 & w40459);
assign w7231 = w6653 & w51818;
assign w7232 = (~w40459 & w47179) | (~w40459 & w47180) | (w47179 & w47180);
assign w7233 = ~w7227 & w7232;
assign w7234 = (w7224 & w6317) | (w7224 & w51819) | (w6317 & w51819);
assign w7235 = (w7234 & w7147) | (w7234 & w40460) | (w7147 & w40460);
assign w7236 = (w80 & w6317) | (w80 & w51820) | (w6317 & w51820);
assign w7237 = ~w7147 & w40461;
assign w7238 = ~w7235 & ~w7237;
assign w7239 = (~w3 & ~w6653) | (~w3 & w51821) | (~w6653 & w51821);
assign w7240 = w7238 & w7239;
assign w7241 = ~w7233 & ~w7240;
assign w7242 = ~w7220 & w7241;
assign w7243 = w6643 & ~w6659;
assign w7244 = (w6735 & w7143) | (w6735 & w51822) | (w7143 & w51822);
assign w7245 = (w7153 & ~w7128) | (w7153 & w44297) | (~w7128 & w44297);
assign w7246 = ~w6316 & ~w6765;
assign w7247 = ~w6737 & w44298;
assign w7248 = ~w6306 & w51823;
assign w7249 = ~w7245 & w7248;
assign w7250 = w7247 & ~w7249;
assign w7251 = (~w6316 & w6737) | (~w6316 & w40462) | (w6737 & w40462);
assign w7252 = w6307 & w6315;
assign w7253 = ~w6765 & w52203;
assign w7254 = ~w6769 & ~w7251;
assign w7255 = w7253 & ~w7254;
assign w7256 = ~w7250 & ~w7255;
assign w7257 = ~w7255 & w44299;
assign w7258 = ~w6765 & ~w7251;
assign w7259 = w6295 & w51824;
assign w7260 = ~w6306 & ~w7259;
assign w7261 = w6296 & w6305;
assign w7262 = (w6737 & w51825) | (w6737 & w51826) | (w51825 & w51826);
assign w7263 = w40465 & ~w7251;
assign w7264 = ~w7262 & ~w7263;
assign w7265 = ~w7261 & w7264;
assign w7266 = w7257 & ~w7265;
assign w7267 = w7242 & ~w7266;
assign w7268 = (w7267 & w7218) | (w7267 & w44300) | (w7218 & w44300);
assign w7269 = w6795 & w6821;
assign w7270 = w7100 & ~w7269;
assign w7271 = w7089 & ~w7090;
assign w7272 = ~w7089 & w7090;
assign w7273 = ~w7271 & ~w7272;
assign w7274 = (w6737 & w44301) | (w6737 & w44302) | (w44301 & w44302);
assign w7275 = ~w6769 & ~w7273;
assign w7276 = ~w7274 & ~w7275;
assign w7277 = ~w7275 & w44303;
assign w7278 = (~w754 & w7113) | (~w754 & w44304) | (w7113 & w44304);
assign w7279 = ~w7277 & ~w7278;
assign w7280 = ~w7270 & w7279;
assign w7281 = (~w493 & w7133) | (~w493 & w51827) | (w7133 & w51827);
assign w7282 = (~w612 & w7120) | (~w612 & w40466) | (w7120 & w40466);
assign w7283 = ~w7135 & w7282;
assign w7284 = ~w7281 & ~w7283;
assign w7285 = w7136 & ~w7280;
assign w7286 = w7284 & ~w7285;
assign w7287 = ~w6763 & w7238;
assign w7288 = w6763 & ~w7230;
assign w7289 = ~w7227 & w7288;
assign w7290 = ~w7287 & ~w7289;
assign w7291 = w3 & w7290;
assign w7292 = (w42 & w7255) | (w42 & w44305) | (w7255 & w44305);
assign w7293 = ~w7265 & ~w7292;
assign w7294 = ~w7257 & w7291;
assign w7295 = w7293 & ~w7294;
assign w7296 = ~w6711 & ~w6756;
assign w7297 = (w7296 & ~w7184) | (w7296 & w40467) | (~w7184 & w40467);
assign w7298 = w7184 & w51828;
assign w7299 = (w6737 & w49527) | (w6737 & w49528) | (w49527 & w49528);
assign w7300 = ~w6769 & w51829;
assign w7301 = (w400 & w7300) | (w400 & w51830) | (w7300 & w51830);
assign w7302 = ~w7294 & w44306;
assign w7303 = w7286 & w7302;
assign w7304 = ~w7268 & w7303;
assign w7305 = ~w7139 & w7304;
assign w7306 = ~w7300 & w40468;
assign w7307 = (w351 & w7193) | (w351 & w40469) | (w7193 & w40469);
assign w7308 = ~w7306 & ~w7307;
assign w7309 = w7202 & ~w7308;
assign w7310 = w7242 & ~w7257;
assign w7311 = w7217 & w7310;
assign w7312 = ~w7309 & w7311;
assign w7313 = w7295 & ~w7312;
assign w7314 = ~w7268 & w7313;
assign w7315 = (~w7314 & w7139) | (~w7314 & w40470) | (w7139 & w40470);
assign w7316 = (~w47168 & w48727) | (~w47168 & w48728) | (w48727 & w48728);
assign w7317 = (w40470 & w47181) | (w40470 & w47182) | (w47181 & w47182);
assign w7318 = (w7068 & w49529) | (w7068 & w49530) | (w49529 & w49530);
assign w7319 = w7317 & ~w7318;
assign w7320 = ~w6776 & w51831;
assign w7321 = (w6777 & w6776) | (w6777 & w51832) | (w6776 & w51832);
assign w7322 = ~w7320 & ~w7321;
assign w7323 = (w6737 & w51833) | (w6737 & w51834) | (w51833 & w51834);
assign w7324 = ~w6769 & w7322;
assign w7325 = ~w7323 & ~w7324;
assign w7326 = ~w7325 & ~w7315;
assign w7327 = (w40470 & w49531) | (w40470 & w49532) | (w49531 & w49532);
assign w7328 = ~w7319 & w7327;
assign w7329 = ~w7085 & ~w7315;
assign w7330 = (w40470 & w49533) | (w40470 & w49534) | (w49533 & w49534);
assign w7331 = ~w6998 & ~w7079;
assign w7332 = (w7331 & w7077) | (w7331 & w47183) | (w7077 & w47183);
assign w7333 = w7066 & w7332;
assign w7334 = ~w6986 & w7333;
assign w7335 = (w1541 & w6996) | (w1541 & w52126) | (w6996 & w52126);
assign w7336 = ~w6996 & w52127;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = ~w7078 & w40472;
assign w7339 = (~w47183 & w48729) | (~w47183 & w48730) | (w48729 & w48730);
assign w7340 = ~w7338 & ~w7339;
assign w7341 = ~w6986 & w47184;
assign w7342 = (w7340 & w6986) | (w7340 & w47185) | (w6986 & w47185);
assign w7343 = ~w7341 & ~w7342;
assign w7344 = ~w7008 & w51835;
assign w7345 = w7315 & w47186;
assign w7346 = (~w7082 & w6986) | (~w7082 & w44311) | (w6986 & w44311);
assign w7347 = (~w40470 & w47187) | (~w40470 & w47188) | (w47187 & w47188);
assign w7348 = w7085 & ~w7346;
assign w7349 = (w6986 & w50177) | (w6986 & w50178) | (w50177 & w50178);
assign w7350 = ~w7348 & ~w7349;
assign w7351 = ~w7347 & ~w7350;
assign w7352 = ~w7345 & ~w7351;
assign w7353 = (~w7009 & ~w7315) | (~w7009 & w47189) | (~w7315 & w47189);
assign w7354 = ~w7330 & w7353;
assign w7355 = w7352 & ~w7354;
assign w7356 = ~w7339 & w40473;
assign w7357 = ~w7334 & w7356;
assign w7358 = ~w6986 & w40474;
assign w7359 = ~w7357 & ~w7358;
assign w7360 = (~w1120 & w7357) | (~w1120 & w40475) | (w7357 & w40475);
assign w7361 = w7315 & w7360;
assign w7362 = ~w1320 & ~w7361;
assign w7363 = ~w7008 & w51836;
assign w7364 = (w7363 & ~w7315) | (w7363 & w47190) | (~w7315 & w47190);
assign w7365 = w7362 & ~w7364;
assign w7366 = ~w7328 & w7365;
assign w7367 = ~w7355 & w7366;
assign w7368 = (w40470 & w47191) | (w40470 & w47192) | (w47191 & w47192);
assign w7369 = ~w7347 & ~w7368;
assign w7370 = w1120 & w7329;
assign w7371 = w1120 & w7350;
assign w7372 = ~w7369 & w7371;
assign w7373 = ~w7370 & ~w7372;
assign w7374 = ~w7328 & ~w7373;
assign w7375 = ~w7367 & ~w7374;
assign w7376 = w7066 & w40476;
assign w7377 = ~w6986 & w7376;
assign w7378 = (w7280 & w7082) | (w7280 & w40477) | (w7082 & w40477);
assign w7379 = (~w7378 & w6986) | (~w7378 & w47193) | (w6986 & w47193);
assign w7380 = (~w7115 & ~w7313) | (~w7115 & w44312) | (~w7313 & w44312);
assign w7381 = w7379 & w7380;
assign w7382 = ~w7305 & w7381;
assign w7383 = w7313 & w49535;
assign w7384 = w7303 & w44313;
assign w7385 = ~w7139 & w7384;
assign w7386 = ~w7383 & ~w7385;
assign w7387 = ~w7382 & w7386;
assign w7388 = ~w7123 & ~w7282;
assign w7389 = ~w493 & ~w7388;
assign w7390 = ~w7387 & w7389;
assign w7391 = ~w493 & w7388;
assign w7392 = w7387 & w7391;
assign w7393 = ~w7390 & ~w7392;
assign w7394 = ~w7270 & ~w7277;
assign w7395 = (w7394 & w7082) | (w7394 & w40478) | (w7082 & w40478);
assign w7396 = w7066 & w44314;
assign w7397 = ~w6986 & w7396;
assign w7398 = (~w6986 & w47194) | (~w6986 & w47195) | (w47194 & w47195);
assign w7399 = (w754 & w7113) | (w754 & w51837) | (w7113 & w51837);
assign w7400 = (w40480 & w6986) | (w40480 & w47196) | (w6986 & w47196);
assign w7401 = ~w7398 & ~w7400;
assign w7402 = w7313 & w49536;
assign w7403 = ~w7113 & w51838;
assign w7404 = ~w7397 & w40481;
assign w7405 = ~w7402 & ~w7404;
assign w7406 = w7303 & w44315;
assign w7407 = ~w7139 & w7406;
assign w7408 = (w7115 & w7397) | (w7115 & w40482) | (w7397 & w40482);
assign w7409 = ~w7407 & ~w7408;
assign w7410 = w7405 & w7409;
assign w7411 = w7315 & ~w7401;
assign w7412 = w7410 & ~w7411;
assign w7413 = w7410 & w40483;
assign w7414 = w7393 & ~w7413;
assign w7415 = w7099 & ~w7277;
assign w7416 = ~w6786 & w7415;
assign w7417 = w7269 & w7415;
assign w7418 = (~w47168 & w48731) | (~w47168 & w48732) | (w48731 & w48732);
assign w7419 = (w40470 & w47199) | (w40470 & w47200) | (w47199 & w47200);
assign w7420 = w6786 & ~w7415;
assign w7421 = w7420 & w52204;
assign w7422 = w754 & w52205;
assign w7423 = (w7068 & w49537) | (w7068 & w49538) | (w49537 & w49538);
assign w7424 = w7419 & w7423;
assign w7425 = ~w7422 & ~w7424;
assign w7426 = (w612 & ~w7410) | (w612 & w40485) | (~w7410 & w40485);
assign w7427 = w7425 & ~w7426;
assign w7428 = w7414 & ~w7427;
assign w7429 = (~w7282 & w7377) | (~w7282 & w51839) | (w7377 & w51839);
assign w7430 = ~w7135 & ~w7281;
assign w7431 = (w7430 & ~w7313) | (w7430 & w51840) | (~w7313 & w51840);
assign w7432 = ~w7305 & w7431;
assign w7433 = ~w7429 & w7432;
assign w7434 = w7134 & ~w7315;
assign w7435 = ~w7433 & ~w7434;
assign w7436 = w7315 & w7429;
assign w7437 = w7315 & w51841;
assign w7438 = w7435 & ~w7437;
assign w7439 = (~w400 & ~w7435) | (~w400 & w40487) | (~w7435 & w40487);
assign w7440 = (w493 & w7387) | (w493 & w40488) | (w7387 & w40488);
assign w7441 = w7387 & w7388;
assign w7442 = w7440 & ~w7441;
assign w7443 = ~w7439 & ~w7442;
assign w7444 = ~w7428 & w7443;
assign w7445 = ~w7319 & ~w7326;
assign w7446 = (w945 & w7319) | (w945 & w44320) | (w7319 & w44320);
assign w7447 = (w40470 & w51842) | (w40470 & w51843) | (w51842 & w51843);
assign w7448 = w7419 & ~w7421;
assign w7449 = w7447 & ~w7448;
assign w7450 = ~w7446 & ~w7449;
assign w7451 = w7414 & w7450;
assign w7452 = w7375 & w7451;
assign w7453 = w7078 & ~w7331;
assign w7454 = ~w7332 & ~w7453;
assign w7455 = w7051 & w7074;
assign w7456 = ~w7034 & w7063;
assign w7457 = w7021 & w7491;
assign w7458 = w7456 & w7457;
assign w7459 = (w7454 & w6986) | (w7454 & w49539) | (w6986 & w49539);
assign w7460 = ~w6986 & w49540;
assign w7461 = ~w7459 & ~w7460;
assign w7462 = w7315 & w7461;
assign w7463 = w7313 & w49541;
assign w7464 = w7303 & w49541;
assign w7465 = ~w7139 & w7464;
assign w7466 = ~w7463 & ~w7465;
assign w7467 = ~w7465 & w40490;
assign w7468 = ~w7462 & w7467;
assign w7469 = (w7063 & w6943) | (w7063 & w49542) | (w6943 & w49542);
assign w7470 = w7303 & w44321;
assign w7471 = ~w7139 & w7470;
assign w7472 = w7313 & w49543;
assign w7473 = ~w7471 & ~w7472;
assign w7474 = ~w7314 & w7469;
assign w7475 = ~w7305 & w7474;
assign w7476 = w7473 & ~w7475;
assign w7477 = w7021 & ~w7034;
assign w7478 = w2285 & ~w7477;
assign w7479 = ~w7476 & w7478;
assign w7480 = w2285 & w7477;
assign w7481 = w7476 & w7480;
assign w7482 = ~w7479 & ~w7481;
assign w7483 = (w7021 & w40491) | (w7021 & w6986) | (w40491 & w6986);
assign w7484 = w7303 & w44322;
assign w7485 = ~w7139 & w7484;
assign w7486 = w7313 & w49544;
assign w7487 = ~w7485 & ~w7486;
assign w7488 = ~w7314 & ~w7483;
assign w7489 = ~w7305 & w7488;
assign w7490 = w7487 & ~w7489;
assign w7491 = w7030 & w7039;
assign w7492 = w2006 & ~w7491;
assign w7493 = ~w7490 & w7492;
assign w7494 = w2006 & w7491;
assign w7495 = w7490 & w7494;
assign w7496 = ~w7493 & ~w7495;
assign w7497 = w7482 & w7496;
assign w7498 = ~w2006 & ~w7491;
assign w7499 = w7490 & w7498;
assign w7500 = ~w2006 & w7491;
assign w7501 = ~w7490 & w7500;
assign w7502 = ~w7499 & ~w7501;
assign w7503 = w7043 & ~w6769;
assign w7504 = (w6737 & w51844) | (w6737 & w51845) | (w51844 & w51845);
assign w7505 = ~w7503 & ~w7504;
assign w7506 = (w7039 & ~w7021) | (w7039 & w49545) | (~w7021 & w49545);
assign w7507 = w7455 & ~w7506;
assign w7508 = ~w7455 & w7506;
assign w7509 = ~w7507 & ~w7508;
assign w7510 = ~w6986 & w40492;
assign w7511 = (w7509 & w6986) | (w7509 & w40493) | (w6986 & w40493);
assign w7512 = ~w7510 & ~w7511;
assign w7513 = ~w1738 & ~w7505;
assign w7514 = w7513 & ~w7315;
assign w7515 = ~w1738 & ~w7512;
assign w7516 = w7315 & w7515;
assign w7517 = ~w7514 & ~w7516;
assign w7518 = w7502 & w7517;
assign w7519 = ~w7497 & w7518;
assign w7520 = ~w7505 & ~w7315;
assign w7521 = w7315 & ~w7512;
assign w7522 = ~w7520 & ~w7521;
assign w7523 = ~w7521 & w49546;
assign w7524 = ~w7462 & w7466;
assign w7525 = (w1541 & w7462) | (w1541 & w49547) | (w7462 & w49547);
assign w7526 = ~w7523 & ~w7525;
assign w7527 = (~w7468 & w7519) | (~w7468 & w40494) | (w7519 & w40494);
assign w7528 = ~w1120 & ~w7350;
assign w7529 = ~w7369 & w7528;
assign w7530 = ~w1120 & w7350;
assign w7531 = w7369 & w7530;
assign w7532 = ~w7529 & ~w7531;
assign w7533 = ~w7008 & w51846;
assign w7534 = (w7533 & ~w7315) | (w7533 & w47201) | (~w7315 & w47201);
assign w7535 = ~w7359 & w7368;
assign w7536 = ~w7534 & ~w7535;
assign w7537 = ~w7328 & w7536;
assign w7538 = w7532 & w7537;
assign w7539 = ~w7374 & ~w7538;
assign w7540 = w7444 & ~w7452;
assign w7541 = w7444 & ~w7539;
assign w7542 = ~w7527 & w7541;
assign w7543 = ~w7540 & ~w7542;
assign w7544 = w6264 & ~w6769;
assign w7545 = (w6737 & w51847) | (w6737 & w51848) | (w51847 & w51848);
assign w7546 = ~w7544 & ~w7545;
assign w7547 = (a[73] & ~w6827) | (a[73] & w51849) | (~w6827 & w51849);
assign w7548 = w6827 & w51850;
assign w7549 = ~w7547 & ~w7548;
assign w7550 = w7546 & ~w7549;
assign w7551 = ~w7546 & w7549;
assign w7552 = ~w7550 & ~w7551;
assign w7553 = ~a[72] & ~w6769;
assign w7554 = a[73] & ~w7553;
assign w7555 = w6823 & ~w7554;
assign w7556 = w7303 & w44323;
assign w7557 = ~w7139 & w7556;
assign w7558 = w7313 & w49548;
assign w7559 = ~w7557 & ~w7558;
assign w7560 = (~w7552 & ~w7313) | (~w7552 & w49549) | (~w7313 & w49549);
assign w7561 = ~w7305 & w7560;
assign w7562 = w7559 & ~w7561;
assign w7563 = ~a[72] & w6264;
assign w7564 = (w6737 & w49550) | (w6737 & w49551) | (w49550 & w49551);
assign w7565 = a[72] & ~w6264;
assign w7566 = ~a[68] & ~a[69];
assign w7567 = ~a[71] & ~w6769;
assign w7568 = ~a[70] & w7566;
assign w7569 = ~w6827 & w7568;
assign w7570 = (w7569 & w7567) | (w7569 & w51851) | (w7567 & w51851);
assign w7571 = w7544 & w7566;
assign w7572 = ~w7570 & ~w7571;
assign w7573 = (~w6828 & w6264) | (~w6828 & w51852) | (w6264 & w51852);
assign w7574 = (w7573 & ~w7564) | (w7573 & w51853) | (~w7564 & w51853);
assign w7575 = (~w5745 & ~w7572) | (~w5745 & w51854) | (~w7572 & w51854);
assign w7576 = (~w7575 & ~w7313) | (~w7575 & w49552) | (~w7313 & w49552);
assign w7577 = (a[71] & ~w7566) | (a[71] & w51855) | (~w7566 & w51855);
assign w7578 = (w7577 & w7553) | (w7577 & w51856) | (w7553 & w51856);
assign w7579 = (w6737 & w49553) | (w6737 & w49554) | (w49553 & w49554);
assign w7580 = ~w7553 & ~w7564;
assign w7581 = ~w6833 & ~w7579;
assign w7582 = w7580 & w7581;
assign w7583 = (~w7578 & w7582) | (~w7578 & w51857) | (w7582 & w51857);
assign w7584 = ~w5745 & w7583;
assign w7585 = w7313 & w49555;
assign w7586 = w7303 & w44324;
assign w7587 = ~w7139 & w7586;
assign w7588 = ~w7585 & ~w7587;
assign w7589 = ~w7305 & w7576;
assign w7590 = w7588 & ~w7589;
assign w7591 = w7562 & ~w7590;
assign w7592 = w7572 & w51858;
assign w7593 = (w7592 & ~w7313) | (w7592 & w49556) | (~w7313 & w49556);
assign w7594 = ~w7305 & w7593;
assign w7595 = w5745 & ~w7583;
assign w7596 = w7303 & w44325;
assign w7597 = ~w7139 & w7596;
assign w7598 = w7313 & w49557;
assign w7599 = ~w7597 & ~w7598;
assign w7600 = ~w7594 & w7599;
assign w7601 = ~w6837 & ~w6839;
assign w7602 = (w7601 & ~w7313) | (w7601 & w51859) | (~w7313 & w51859);
assign w7603 = ~w5330 & ~w6845;
assign w7604 = (w40495 & ~w7313) | (w40495 & w49558) | (~w7313 & w49558);
assign w7605 = ~w7305 & w7604;
assign w7606 = ~w5330 & w6845;
assign w7607 = (w7313 & w49559) | (w7313 & w49560) | (w49559 & w49560);
assign w7608 = w7303 & w44326;
assign w7609 = ~w7139 & w7608;
assign w7610 = ~w7607 & ~w7609;
assign w7611 = ~w7605 & w7610;
assign w7612 = w7600 & w7611;
assign w7613 = ~w7591 & w7612;
assign w7614 = w5330 & w6845;
assign w7615 = (w40497 & ~w7313) | (w40497 & w49561) | (~w7313 & w49561);
assign w7616 = ~w7305 & w7615;
assign w7617 = w5330 & ~w6845;
assign w7618 = (w7313 & w49562) | (w7313 & w49563) | (w49562 & w49563);
assign w7619 = w7303 & w44327;
assign w7620 = ~w7139 & w7619;
assign w7621 = ~w7618 & ~w7620;
assign w7622 = ~w7616 & w7621;
assign w7623 = (w5330 & w6846) | (w5330 & w51860) | (w6846 & w51860);
assign w7624 = ~w6846 & w51861;
assign w7625 = ~w7623 & ~w7624;
assign w7626 = (~w7625 & ~w7313) | (~w7625 & w51862) | (~w7313 & w51862);
assign w7627 = ~w4838 & ~w6895;
assign w7628 = (w40499 & ~w7313) | (w40499 & w51863) | (~w7313 & w51863);
assign w7629 = ~w7305 & w7628;
assign w7630 = ~w4838 & w6895;
assign w7631 = (w7313 & w51864) | (w7313 & w51865) | (w51864 & w51865);
assign w7632 = w7303 & w44328;
assign w7633 = ~w7139 & w7632;
assign w7634 = ~w7631 & ~w7633;
assign w7635 = ~w7629 & w7634;
assign w7636 = w7622 & w7635;
assign w7637 = ~w5330 & ~w6895;
assign w7638 = (w6847 & w49564) | (w6847 & w49565) | (w49564 & w49565);
assign w7639 = (~w6847 & w49566) | (~w6847 & w49567) | (w49566 & w49567);
assign w7640 = ~w7638 & ~w7639;
assign w7641 = (w7640 & ~w7313) | (w7640 & w51866) | (~w7313 & w51866);
assign w7642 = w4430 & ~w6873;
assign w7643 = (w7642 & w7305) | (w7642 & w40502) | (w7305 & w40502);
assign w7644 = w4430 & w6873;
assign w7645 = ~w7305 & w40503;
assign w7646 = ~w7643 & ~w7645;
assign w7647 = w7636 & w7646;
assign w7648 = ~w7613 & w7647;
assign w7649 = w4838 & w6895;
assign w7650 = (w40504 & ~w7313) | (w40504 & w51867) | (~w7313 & w51867);
assign w7651 = ~w7305 & w7650;
assign w7652 = w4838 & ~w6895;
assign w7653 = (w7313 & w51868) | (w7313 & w51869) | (w51868 & w51869);
assign w7654 = w7303 & w44329;
assign w7655 = ~w7139 & w7654;
assign w7656 = ~w7653 & ~w7655;
assign w7657 = ~w7651 & w7656;
assign w7658 = ~w4430 & ~w6873;
assign w7659 = ~w7314 & w40506;
assign w7660 = ~w4430 & w6873;
assign w7661 = (~w7660 & w7314) | (~w7660 & w40507) | (w7314 & w40507);
assign w7662 = w7303 & w44330;
assign w7663 = ~w7139 & w7662;
assign w7664 = ~w7661 & ~w7663;
assign w7665 = ~w7305 & w7659;
assign w7666 = w7664 & ~w7665;
assign w7667 = w7657 & ~w7666;
assign w7668 = w7646 & ~w7667;
assign w7669 = w4056 & w6907;
assign w7670 = ~w6888 & w7669;
assign w7671 = ~w4056 & ~w6907;
assign w7672 = w6886 & w47202;
assign w7673 = ~w6847 & w7672;
assign w7674 = ~w7671 & ~w7673;
assign w7675 = ~w7670 & w7674;
assign w7676 = ~w6382 & w6947;
assign w7677 = ~w6954 & ~w7676;
assign w7678 = w3646 & ~w7677;
assign w7679 = ~w7305 & w40508;
assign w7680 = w3646 & w7677;
assign w7681 = (w7680 & w7305) | (w7680 & w40509) | (w7305 & w40509);
assign w7682 = ~w7679 & ~w7681;
assign w7683 = w6885 & ~w6902;
assign w7684 = (~w6903 & ~w40510) | (~w6903 & w49568) | (~w40510 & w49568);
assign w7685 = w6862 & ~w6874;
assign w7686 = (w7685 & w6846) | (w7685 & w49569) | (w6846 & w49569);
assign w7687 = (w7683 & w7686) | (w7683 & w40511) | (w7686 & w40511);
assign w7688 = ~w7686 & w40512;
assign w7689 = ~w7687 & ~w7688;
assign w7690 = ~w4056 & ~w6901;
assign w7691 = w7690 & ~w7315;
assign w7692 = ~w4056 & w7689;
assign w7693 = w7692 & w7315;
assign w7694 = ~w7691 & ~w7693;
assign w7695 = w7682 & w7694;
assign w7696 = ~w7668 & w7695;
assign w7697 = ~w7648 & w7696;
assign w7698 = ~w6958 & w40513;
assign w7699 = (w6982 & w6943) | (w6982 & w40514) | (w6943 & w40514);
assign w7700 = (~w3242 & w6943) | (~w3242 & w40515) | (w6943 & w40515);
assign w7701 = (w6943 & w51870) | (w6943 & w51871) | (w51870 & w51871);
assign w7702 = ~w7699 & ~w7700;
assign w7703 = (~w7701 & ~w7702) | (~w7701 & w51872) | (~w7702 & w51872);
assign w7704 = (w6943 & w51873) | (w6943 & w51874) | (w51873 & w51874);
assign w7705 = (~w7704 & ~w7702) | (~w7704 & w51875) | (~w7702 & w51875);
assign w7706 = (~w2558 & ~w7315) | (~w2558 & w51876) | (~w7315 & w51876);
assign w7707 = (w7055 & ~w7315) | (w7055 & w51877) | (~w7315 & w51877);
assign w7708 = w7706 & ~w7707;
assign w7709 = ~w6943 & w40516;
assign w7710 = ~w7314 & w40517;
assign w7711 = (w6982 & w7305) | (w6982 & w40518) | (w7305 & w40518);
assign w7712 = ~w7305 & w40519;
assign w7713 = ~w7711 & ~w7712;
assign w7714 = w2896 & ~w7713;
assign w7715 = ~w7708 & ~w7714;
assign w7716 = w4056 & ~w7689;
assign w7717 = ~w7314 & ~w7716;
assign w7718 = w4056 & w6901;
assign w7719 = w7313 & w49570;
assign w7720 = w7303 & w44331;
assign w7721 = ~w7139 & w7720;
assign w7722 = ~w7719 & ~w7721;
assign w7723 = ~w7305 & w7717;
assign w7724 = w7722 & ~w7723;
assign w7725 = ~w3646 & w7677;
assign w7726 = ~w7314 & w40520;
assign w7727 = ~w7305 & w7726;
assign w7728 = ~w3646 & ~w7677;
assign w7729 = (w7728 & w7314) | (w7728 & w40521) | (w7314 & w40521);
assign w7730 = w7303 & w44332;
assign w7731 = ~w7139 & w7730;
assign w7732 = ~w7729 & ~w7731;
assign w7733 = ~w7727 & w7732;
assign w7734 = ~w7724 & w7733;
assign w7735 = w3646 & ~w7670;
assign w7736 = w7674 & ~w7677;
assign w7737 = w7735 & ~w7736;
assign w7738 = ~w3646 & w7670;
assign w7739 = w7674 & w7728;
assign w7740 = ~w7738 & ~w7739;
assign w7741 = ~w7314 & ~w7737;
assign w7742 = w7740 & w7741;
assign w7743 = w4056 & w6938;
assign w7744 = w6957 & ~w7743;
assign w7745 = (~w3242 & ~w6957) | (~w3242 & w51878) | (~w6957 & w51878);
assign w7746 = (w7745 & ~w7742) | (w7745 & w47203) | (~w7742 & w47203);
assign w7747 = w6957 & w51879;
assign w7748 = w7742 & w47204;
assign w7749 = ~w7746 & ~w7748;
assign w7750 = ~w2896 & ~w6982;
assign w7751 = (w7750 & w7305) | (w7750 & w40522) | (w7305 & w40522);
assign w7752 = ~w2896 & w6982;
assign w7753 = ~w7305 & w40523;
assign w7754 = ~w7751 & ~w7753;
assign w7755 = w7682 & ~w7734;
assign w7756 = ~w7749 & w7754;
assign w7757 = ~w7755 & ~w7756;
assign w7758 = w7715 & w7757;
assign w7759 = ~w7697 & w7758;
assign w7760 = w7742 & w49571;
assign w7761 = (w7744 & ~w7742) | (w7744 & w49572) | (~w7742 & w49572);
assign w7762 = ~w7760 & ~w7761;
assign w7763 = w3242 & ~w7762;
assign w7764 = (w7754 & w7762) | (w7754 & w40524) | (w7762 & w40524);
assign w7765 = w7715 & ~w7764;
assign w7766 = w2558 & w7055;
assign w7767 = (w7766 & ~w7315) | (w7766 & w51880) | (~w7315 & w51880);
assign w7768 = w7315 & w52083;
assign w7769 = ~w7767 & ~w7768;
assign w7770 = ~w2285 & ~w7477;
assign w7771 = w7476 & w7770;
assign w7772 = ~w2285 & w7477;
assign w7773 = ~w7476 & w7772;
assign w7774 = ~w7771 & ~w7773;
assign w7775 = w7769 & w7774;
assign w7776 = ~w7468 & w7517;
assign w7777 = w7502 & w7776;
assign w7778 = w7775 & w7777;
assign w7779 = ~w7765 & w7778;
assign w7780 = ~w7759 & w7779;
assign w7781 = w7375 & w7780;
assign w7782 = ~w7543 & ~w7781;
assign w7783 = w7435 & w51881;
assign w7784 = ~w7138 & w7286;
assign w7785 = w7067 & w7286;
assign w7786 = ~w6986 & w7785;
assign w7787 = ~w7784 & ~w7786;
assign w7788 = (~w7301 & w7786) | (~w7301 & w47205) | (w7786 & w47205);
assign w7789 = ~w351 & ~w7306;
assign w7790 = (~w7789 & ~w7313) | (~w7789 & w51882) | (~w7313 & w51882);
assign w7791 = ~w7788 & ~w7790;
assign w7792 = (~w351 & ~w7303) | (~w351 & w49573) | (~w7303 & w49573);
assign w7793 = (w7786 & w49574) | (w7786 & w49575) | (w49574 & w49575);
assign w7794 = w7788 & ~w7792;
assign w7795 = w7793 & ~w7794;
assign w7796 = ~w7195 & w7306;
assign w7797 = ~w7307 & w7796;
assign w7798 = (w7797 & ~w7313) | (w7797 & w44333) | (~w7313 & w44333);
assign w7799 = (w7313 & w44334) | (w7313 & w44335) | (w44334 & w44335);
assign w7800 = ~w7798 & ~w7799;
assign w7801 = ~w7193 & w51883;
assign w7802 = w7306 & w7801;
assign w7803 = (~w7802 & ~w7788) | (~w7802 & w40527) | (~w7788 & w40527);
assign w7804 = ~w7788 & ~w7800;
assign w7805 = w7803 & ~w7804;
assign w7806 = ~w7791 & w7795;
assign w7807 = w7805 & ~w7806;
assign w7808 = (w252 & w7806) | (w252 & w40528) | (w7806 & w40528);
assign w7809 = (~w7195 & ~w7313) | (~w7195 & w49576) | (~w7313 & w49576);
assign w7810 = ~w7305 & w7809;
assign w7811 = (w7308 & w40529) | (w7308 & w7787) | (w40529 & w7787);
assign w7812 = w7810 & ~w7811;
assign w7813 = w7201 & w7216;
assign w7814 = w57 & ~w7813;
assign w7815 = ~w7812 & w40530;
assign w7816 = w57 & w7813;
assign w7817 = (w7816 & w7812) | (w7816 & w40531) | (w7812 & w40531);
assign w7818 = ~w7815 & ~w7817;
assign w7819 = ~w7808 & w7818;
assign w7820 = ~w7806 & w40532;
assign w7821 = ~w7786 & w47206;
assign w7822 = (w400 & w7786) | (w400 & w47207) | (w7786 & w47207);
assign w7823 = ~w7821 & ~w7822;
assign w7824 = (w6737 & w51884) | (w6737 & w51885) | (w51884 & w51885);
assign w7825 = ~w6769 & w7185;
assign w7826 = ~w7825 & w51886;
assign w7827 = (~w7296 & w7825) | (~w7296 & w51887) | (w7825 & w51887);
assign w7828 = ~w7826 & ~w7827;
assign w7829 = ~w7823 & w40533;
assign w7830 = (w7828 & w7823) | (w7828 & w40534) | (w7823 & w40534);
assign w7831 = ~w7829 & ~w7830;
assign w7832 = ~w351 & ~w7831;
assign w7833 = ~w7820 & w7832;
assign w7834 = w7819 & ~w7833;
assign w7835 = ~w57 & ~w7813;
assign w7836 = (w7835 & w7812) | (w7835 & w40535) | (w7812 & w40535);
assign w7837 = ~w57 & w7813;
assign w7838 = ~w7812 & w40536;
assign w7839 = ~w7836 & ~w7838;
assign w7840 = (w7839 & w7833) | (w7839 & w50286) | (w7833 & w50286);
assign w7841 = (~w7783 & w7834) | (~w7783 & w44336) | (w7834 & w44336);
assign w7842 = w7444 & ~w7451;
assign w7843 = w7201 & w51888;
assign w7844 = w7217 & ~w7309;
assign w7845 = (w7786 & w49577) | (w7786 & w49578) | (w49577 & w49578);
assign w7846 = ~w7161 & ~w7220;
assign w7847 = w7846 & w7315;
assign w7848 = ~w7845 & w7847;
assign w7849 = w7160 & ~w7315;
assign w7850 = (w40470 & w47208) | (w40470 & w47209) | (w47208 & w47209);
assign w7851 = w7845 & w7850;
assign w7852 = ~w7849 & ~w7851;
assign w7853 = (w3 & ~w7847) | (w3 & w44339) | (~w7847 & w44339);
assign w7854 = w7852 & w7853;
assign w7855 = ~w7309 & w51889;
assign w7856 = (w40538 & w7855) | (w40538 & w7787) | (w7855 & w7787);
assign w7857 = ~w7179 & ~w7220;
assign w7858 = ~w7856 & ~w7857;
assign w7859 = w7303 & w44340;
assign w7860 = ~w7139 & w7859;
assign w7861 = w7313 & w49579;
assign w7862 = ~w7860 & ~w7861;
assign w7863 = w7241 & ~w7291;
assign w7864 = (~w7863 & ~w7313) | (~w7863 & w49580) | (~w7313 & w49580);
assign w7865 = ~w7305 & w7864;
assign w7866 = (w7863 & ~w7313) | (w7863 & w49581) | (~w7313 & w49581);
assign w7867 = ~w7305 & w7866;
assign w7868 = w7862 & ~w7867;
assign w7869 = w7858 & w7868;
assign w7870 = w7862 & ~w7865;
assign w7871 = ~w7858 & w7870;
assign w7872 = ~w7869 & ~w7871;
assign w7873 = w42 & w7872;
assign w7874 = ~w7291 & ~w7857;
assign w7875 = ~w6296 & ~w7258;
assign w7876 = w6295 & w51890;
assign w7877 = w7258 & w7876;
assign w7878 = ~w7875 & ~w7877;
assign w7879 = w7256 & ~w7878;
assign w7880 = w7256 & w51891;
assign w7881 = ~w7292 & ~w7880;
assign w7882 = w7256 & ~w7265;
assign w7883 = (w7787 & w51892) | (w7787 & w51893) | (w51892 & w51893);
assign w7884 = w7881 & ~w7882;
assign w7885 = w7884 & w52206;
assign w7886 = ~w7883 & ~w7885;
assign w7887 = ~w7873 & w40539;
assign w7888 = (w7216 & ~w7202) | (w7216 & w51894) | (~w7202 & w51894);
assign w7889 = (~w7786 & w47212) | (~w7786 & w47213) | (w47212 & w47213);
assign w7890 = w7178 & w7211;
assign w7891 = ~w7889 & w7890;
assign w7892 = w7315 & ~w7891;
assign w7893 = w7889 & ~w7890;
assign w7894 = w7892 & ~w7893;
assign w7895 = ~w7172 & w51895;
assign w7896 = (w7173 & w7172) | (w7173 & w51896) | (w7172 & w51896);
assign w7897 = ~w7895 & ~w7896;
assign w7898 = ~w7897 & ~w7315;
assign w7899 = ~w80 & ~w7898;
assign w7900 = ~w7894 & w7899;
assign w7901 = w7887 & ~w7900;
assign w7902 = ~w7842 & w7901;
assign w7903 = ~w7842 & w44343;
assign w7904 = (w7903 & w7543) | (w7903 & w44344) | (w7543 & w44344);
assign w7905 = ~w42 & ~w7872;
assign w7906 = w7256 & w52206;
assign w7907 = (w7787 & w49582) | (w7787 & w49583) | (w49582 & w49583);
assign w7908 = ~w7906 & ~w7907;
assign w7909 = ~w7872 & w44345;
assign w7910 = ~w7887 & ~w7909;
assign w7911 = w351 & w7831;
assign w7912 = ~w7820 & ~w7911;
assign w7913 = w7819 & ~w7912;
assign w7914 = ~w7912 & w47214;
assign w7915 = (~w7898 & ~w7892) | (~w7898 & w49584) | (~w7892 & w49584);
assign w7916 = w80 & ~w7915;
assign w7917 = ~w7839 & ~w7900;
assign w7918 = ~w7916 & ~w7917;
assign w7919 = ~w7848 & w7852;
assign w7920 = (~w3 & ~w7852) | (~w3 & w49585) | (~w7852 & w49585);
assign w7921 = ~w7909 & ~w7920;
assign w7922 = w7918 & w7921;
assign w7923 = (~w7910 & ~w7922) | (~w7910 & w40541) | (~w7922 & w40541);
assign w7924 = (~w44344 & w47215) | (~w44344 & w47216) | (w47215 & w47216);
assign w7925 = w7350 & ~w7369;
assign w7926 = ~w7350 & w7369;
assign w7927 = ~w7925 & ~w7926;
assign w7928 = ~w7527 & ~w7780;
assign w7929 = (w1320 & w7780) | (w1320 & w40542) | (w7780 & w40542);
assign w7930 = (w7009 & ~w7315) | (w7009 & w51897) | (~w7315 & w51897);
assign w7931 = w7315 & w51898;
assign w7932 = ~w7930 & ~w7931;
assign w7933 = ~w7462 & w51899;
assign w7934 = (~w7933 & w7519) | (~w7933 & w40543) | (w7519 & w40543);
assign w7935 = ~w7780 & ~w7934;
assign w7936 = (~w7932 & w7780) | (~w7932 & w40544) | (w7780 & w40544);
assign w7937 = ~w7929 & ~w7936;
assign w7938 = w1120 & ~w7927;
assign w7939 = w7532 & ~w7938;
assign w7940 = w7937 & ~w7939;
assign w7941 = ~w7937 & w7939;
assign w7942 = ~w7940 & ~w7941;
assign w7943 = (w44344 & w50287) | (w44344 & w50288) | (w50287 & w50288);
assign w7944 = w7924 & w7942;
assign w7945 = ~w7943 & ~w7944;
assign w7946 = w7425 & ~w7539;
assign w7947 = ~w7780 & w40546;
assign w7948 = ~w7367 & w47217;
assign w7949 = (~w7413 & w7948) | (~w7413 & w51900) | (w7948 & w51900);
assign w7950 = ~w7426 & w7947;
assign w7951 = ~w7904 & w40547;
assign w7952 = ~w493 & w7923;
assign w7953 = w7902 & w40548;
assign w7954 = (~w7952 & w7782) | (~w7952 & w40549) | (w7782 & w40549);
assign w7955 = w7393 & ~w7442;
assign w7956 = w400 & w7955;
assign w7957 = w7954 & w7956;
assign w7958 = ~w7951 & w7957;
assign w7959 = w400 & ~w7955;
assign w7960 = ~w7954 & w7959;
assign w7961 = (w7959 & w7950) | (w7959 & w49586) | (w7950 & w49586);
assign w7962 = w7924 & w7961;
assign w7963 = ~w7960 & ~w7962;
assign w7964 = ~w7958 & w7963;
assign w7965 = (w612 & w7947) | (w612 & w44346) | (w7947 & w44346);
assign w7966 = ~w7947 & w44347;
assign w7967 = ~w7965 & ~w7966;
assign w7968 = (w7412 & ~w7924) | (w7412 & w40550) | (~w7924 & w40550);
assign w7969 = w7924 & w40551;
assign w7970 = ~w7968 & ~w7969;
assign w7971 = w493 & w7970;
assign w7972 = ~w400 & w52207;
assign w7973 = ~w7951 & w50289;
assign w7974 = w7972 & ~w7973;
assign w7975 = w7964 & w7971;
assign w7976 = ~w7974 & ~w7975;
assign w7977 = ~w7355 & w7365;
assign w7978 = w7373 & ~w7977;
assign w7979 = w7532 & w7536;
assign w7980 = (w7978 & w7780) | (w7978 & w44348) | (w7780 & w44348);
assign w7981 = ~w945 & w7980;
assign w7982 = w945 & ~w7980;
assign w7983 = ~w7981 & ~w7982;
assign w7984 = ~w7319 & w51901;
assign w7985 = (w7984 & ~w7924) | (w7984 & w40552) | (~w7924 & w40552);
assign w7986 = (w754 & w7319) | (w754 & w51902) | (w7319 & w51902);
assign w7987 = w7924 & w40553;
assign w7988 = ~w7985 & ~w7987;
assign w7989 = ~w7367 & w7539;
assign w7990 = ~w7780 & w40554;
assign w7991 = ~w7539 & ~w7978;
assign w7992 = ~w7923 & ~w7990;
assign w7993 = ~w7446 & ~w7991;
assign w7994 = w7992 & w7993;
assign w7995 = w7902 & w40555;
assign w7996 = w754 & w7923;
assign w7997 = (~w7996 & w7782) | (~w7996 & w40556) | (w7782 & w40556);
assign w7998 = ~w7904 & w7994;
assign w7999 = w7997 & ~w7998;
assign w8000 = w7425 & ~w7449;
assign w8001 = w612 & ~w8000;
assign w8002 = (w8001 & w7998) | (w8001 & w40557) | (w7998 & w40557);
assign w8003 = w612 & w8000;
assign w8004 = ~w7998 & w40558;
assign w8005 = ~w8002 & ~w8004;
assign w8006 = w7988 & w8005;
assign w8007 = ~w7944 & w40559;
assign w8008 = (~w754 & w7319) | (~w754 & w51903) | (w7319 & w51903);
assign w8009 = (w8008 & ~w7924) | (w8008 & w40560) | (~w7924 & w40560);
assign w8010 = ~w7319 & w51904;
assign w8011 = w7924 & w40561;
assign w8012 = ~w8009 & ~w8011;
assign w8013 = ~w8007 & w8012;
assign w8014 = w8006 & ~w8013;
assign w8015 = ~w7923 & ~w7929;
assign w8016 = (~w7932 & w7904) | (~w7932 & w40562) | (w7904 & w40562);
assign w8017 = ~w7904 & w40563;
assign w8018 = ~w8016 & ~w8017;
assign w8019 = ~w1120 & ~w8018;
assign w8020 = (~w945 & w7944) | (~w945 & w40564) | (w7944 & w40564);
assign w8021 = ~w8019 & ~w8020;
assign w8022 = w8006 & w8021;
assign w8023 = ~w612 & ~w8000;
assign w8024 = ~w7998 & w40565;
assign w8025 = ~w612 & w8000;
assign w8026 = (w8025 & w7998) | (w8025 & w40566) | (w7998 & w40566);
assign w8027 = ~w8024 & ~w8026;
assign w8028 = w7964 & w8027;
assign w8029 = ~w493 & w7412;
assign w8030 = (w8029 & ~w7924) | (w8029 & w40567) | (~w7924 & w40567);
assign w8031 = ~w493 & ~w7412;
assign w8032 = w7924 & w40568;
assign w8033 = ~w8030 & ~w8032;
assign w8034 = ~w8014 & ~w8022;
assign w8035 = w8028 & w8033;
assign w8036 = w8034 & w8035;
assign w8037 = (w7976 & ~w8034) | (w7976 & w44349) | (~w8034 & w44349);
assign w8038 = w7451 & ~w7991;
assign w8039 = ~w7928 & w8038;
assign w8040 = (~w7442 & ~w7414) | (~w7442 & w40569) | (~w7414 & w40569);
assign w8041 = (w8040 & ~w7375) | (w8040 & w49587) | (~w7375 & w49587);
assign w8042 = ~w7539 & w8040;
assign w8043 = ~w7527 & w8042;
assign w8044 = ~w8041 & ~w8043;
assign w8045 = ~w8039 & w40570;
assign w8046 = (w400 & w8039) | (w400 & w40571) | (w8039 & w40571);
assign w8047 = ~w8045 & ~w8046;
assign w8048 = w7438 & ~w7923;
assign w8049 = (w8048 & w7782) | (w8048 & w40572) | (w7782 & w40572);
assign w8050 = ~w8047 & w8049;
assign w8051 = (~w40573 & w47219) | (~w40573 & w47220) | (w47219 & w47220);
assign w8052 = ~w7543 & ~w8039;
assign w8053 = w7831 & ~w8052;
assign w8054 = ~w8051 & ~w8053;
assign w8055 = (~w351 & ~w8052) | (~w351 & w8071) | (~w8052 & w8071);
assign w8056 = ~w7439 & w7911;
assign w8057 = w252 & w8056;
assign w8058 = (w8057 & w8052) | (w8057 & w49588) | (w8052 & w49588);
assign w8059 = ~w8050 & ~w8054;
assign w8060 = (~w8058 & ~w8059) | (~w8058 & w44350) | (~w8059 & w44350);
assign w8061 = (w252 & w333) | (w252 & w51905) | (w333 & w51905);
assign w8062 = ~w8061 & ~w7924;
assign w8063 = (~w7438 & w8047) | (~w7438 & w47221) | (w8047 & w47221);
assign w8064 = (w47216 & w49589) | (w47216 & w49590) | (w49589 & w49590);
assign w8065 = (~w8064 & w8063) | (~w8064 & w44351) | (w8063 & w44351);
assign w8066 = (w351 & w8052) | (w351 & w40574) | (w8052 & w40574);
assign w8067 = ~w8052 & w40575;
assign w8068 = ~w8066 & ~w8067;
assign w8069 = (w252 & w8068) | (w252 & w44352) | (w8068 & w44352);
assign w8070 = ~w8039 & w49591;
assign w8071 = w7435 & w51906;
assign w8072 = (w8071 & ~w7924) | (w8071 & w49592) | (~w7924 & w49592);
assign w8073 = ~w8060 & ~w8065;
assign w8074 = (~w7831 & w8069) | (~w7831 & w49593) | (w8069 & w49593);
assign w8075 = ~w8073 & ~w8074;
assign w8076 = ~w7808 & ~w7820;
assign w8077 = w7414 & w51907;
assign w8078 = (~w7911 & w7928) | (~w7911 & w40576) | (w7928 & w40576);
assign w8079 = ~w7542 & w44353;
assign w8080 = ~w8076 & w52208;
assign w8081 = ~w7832 & w8076;
assign w8082 = (w8081 & w8079) | (w8081 & w40578) | (w8079 & w40578);
assign w8083 = w7924 & ~w8082;
assign w8084 = ~w8080 & w8083;
assign w8085 = (w44344 & w50290) | (w44344 & w50291) | (w50290 & w50291);
assign w8086 = (~w8085 & ~w8083) | (~w8085 & w40580) | (~w8083 & w40580);
assign w8087 = ~w57 & ~w8086;
assign w8088 = w57 & w7923;
assign w8089 = w7902 & w40581;
assign w8090 = (~w8088 & w7782) | (~w8088 & w40582) | (w7782 & w40582);
assign w8091 = (~w40541 & w44354) | (~w40541 & w44355) | (w44354 & w44355);
assign w8092 = (w8091 & w7782) | (w8091 & w40583) | (w7782 & w40583);
assign w8093 = ~w8082 & w8092;
assign w8094 = w7818 & w7839;
assign w8095 = w80 & w8094;
assign w8096 = (w8095 & w8093) | (w8095 & w44356) | (w8093 & w44356);
assign w8097 = w80 & ~w8094;
assign w8098 = ~w8093 & w44357;
assign w8099 = ~w8096 & ~w8098;
assign w8100 = ~w8087 & w8099;
assign w8101 = ~w8075 & w8100;
assign w8102 = w7841 & ~w7842;
assign w8103 = (w8102 & w7543) | (w8102 & w40584) | (w7543 & w40584);
assign w8104 = (~w7900 & w7913) | (~w7900 & w7917) | (w7913 & w7917);
assign w8105 = ~w7916 & ~w8104;
assign w8106 = (w8105 & ~w8103) | (w8105 & w44358) | (~w8103 & w44358);
assign w8107 = ~w7854 & ~w7920;
assign w8108 = ~w7919 & ~w7924;
assign w8109 = w40585 & ~w7904;
assign w8110 = w8106 & w8109;
assign w8111 = ~w8108 & ~w8110;
assign w8112 = w40586 & ~w7904;
assign w8113 = ~w8106 & w8112;
assign w8114 = (~w7915 & w7887) | (~w7915 & w51908) | (w7887 & w51908);
assign w8115 = ~w7900 & ~w7916;
assign w8116 = ~w7913 & w51909;
assign w8117 = ~w8114 & w8116;
assign w8118 = ~w8103 & w8117;
assign w8119 = ~w7910 & ~w7921;
assign w8120 = ~w8104 & ~w8119;
assign w8121 = ~w7916 & ~w8114;
assign w8122 = ~w8103 & w49594;
assign w8123 = ~w8114 & w51910;
assign w8124 = (w8103 & w49595) | (w8103 & w49596) | (w49595 & w49596);
assign w8125 = ~w8122 & ~w8124;
assign w8126 = ~w7917 & w51911;
assign w8127 = ~w7914 & w8126;
assign w8128 = ~w7872 & w7886;
assign w8129 = ~w7873 & ~w7905;
assign w8130 = w8129 & w51912;
assign w8131 = (w8103 & w49597) | (w8103 & w49598) | (w49597 & w49598);
assign w8132 = ~w8128 & ~w8129;
assign w8133 = ~w8129 & w51913;
assign w8134 = w8127 & w8132;
assign w8135 = (w8103 & w49599) | (w8103 & w49600) | (w49599 & w49600);
assign w8136 = ~w8131 & w8135;
assign w8137 = w8125 & w8136;
assign w8138 = w42 & ~w8113;
assign w8139 = w8111 & w8138;
assign w8140 = w8137 & ~w8139;
assign w8141 = w57 & ~w8085;
assign w8142 = ~w8084 & w8141;
assign w8143 = ~w80 & w8094;
assign w8144 = w8090 & w8143;
assign w8145 = ~w8093 & w8144;
assign w8146 = ~w80 & ~w8094;
assign w8147 = ~w8090 & w8146;
assign w8148 = w8091 & w8146;
assign w8149 = (~w44344 & w47222) | (~w44344 & w47223) | (w47222 & w47223);
assign w8150 = ~w8082 & w8149;
assign w8151 = ~w8147 & ~w8150;
assign w8152 = ~w8145 & w8151;
assign w8153 = ~w8142 & w8152;
assign w8154 = w8099 & ~w8153;
assign w8155 = w8140 & ~w8154;
assign w8156 = ~w8101 & w8155;
assign w8157 = ~w8037 & w8156;
assign w8158 = ~w8050 & ~w8063;
assign w8159 = (w351 & w8063) | (w351 & w44362) | (w8063 & w44362);
assign w8160 = w351 & ~w7831;
assign w8161 = (w7832 & w8052) | (w7832 & w40587) | (w8052 & w40587);
assign w8162 = ~w8052 & w40588;
assign w8163 = ~w8161 & ~w8162;
assign w8164 = w40589 & ~w7904;
assign w8165 = ~w8068 & w8164;
assign w8166 = (w44344 & w50292) | (w44344 & w50293) | (w50292 & w50293);
assign w8167 = w8163 & ~w8166;
assign w8168 = ~w8165 & w8167;
assign w8169 = w252 & ~w8168;
assign w8170 = ~w252 & w8168;
assign w8171 = ~w8087 & ~w8170;
assign w8172 = w8159 & ~w8169;
assign w8173 = w8171 & ~w8172;
assign w8174 = (w8103 & w51914) | (w8103 & w51915) | (w51914 & w51915);
assign w8175 = ~w7872 & w51916;
assign w8176 = w8175 & w52209;
assign w8177 = ~w8174 & ~w8176;
assign w8178 = w8111 & ~w8113;
assign w8179 = ~w8178 & w49603;
assign w8180 = (w8103 & w51917) | (w8103 & w51918) | (w51917 & w51918);
assign w8181 = ~w8118 & ~w8180;
assign w8182 = ~w8180 & w49604;
assign w8183 = w8099 & ~w8182;
assign w8184 = w8140 & ~w8183;
assign w8185 = ~w8179 & ~w8184;
assign w8186 = w8140 & w8153;
assign w8187 = ~w8173 & w8186;
assign w8188 = w8185 & ~w8187;
assign w8189 = ~w8157 & w8188;
assign w8190 = ~a[70] & w7315;
assign w8191 = ~a[71] & ~w8190;
assign w8192 = a[71] & w8190;
assign w8193 = ~w8191 & ~w8192;
assign w8194 = w6264 & ~w8193;
assign w8195 = a[71] & ~w7315;
assign w8196 = w7577 & ~w6769;
assign w8197 = w7568 & ~w6769;
assign w8198 = ~w7579 & ~w8197;
assign w8199 = ~w7314 & w52210;
assign w8200 = ~w8198 & ~w7315;
assign w8201 = ~w8199 & ~w8200;
assign w8202 = (~w8196 & ~w8201) | (~w8196 & w51920) | (~w8201 & w51920);
assign w8203 = (w6264 & w8202) | (w6264 & w51921) | (w8202 & w51921);
assign w8204 = w7887 & ~w8127;
assign w8205 = w6769 & ~w7315;
assign w8206 = (w8199 & w7872) | (w8199 & w51922) | (w7872 & w51922);
assign w8207 = ~w7568 & w8205;
assign w8208 = ~w8206 & ~w8207;
assign w8209 = (w7564 & w8206) | (w7564 & w51923) | (w8206 & w51923);
assign w8210 = w8195 & ~w8198;
assign w8211 = ~w8210 & w52211;
assign w8212 = w7902 & w40591;
assign w8213 = (~w8211 & w7782) | (~w8211 & w51925) | (w7782 & w51925);
assign w8214 = w40592 & ~w7904;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = ~w8194 & ~w7924;
assign w8217 = w8215 & ~w8216;
assign w8218 = ~a[66] & ~a[67];
assign w8219 = ~w7314 & w52212;
assign w8220 = ~a[68] & w8218;
assign w8221 = ~w8220 & ~w7315;
assign w8222 = w7566 & ~w8219;
assign w8223 = a[69] & w8221;
assign w8224 = ~w8222 & ~w8223;
assign w8225 = ~w7314 & w52213;
assign w8226 = a[69] & ~w8225;
assign w8227 = ~w8221 & ~w8226;
assign w8228 = ~w8227 & w7923;
assign w8229 = w7902 & w40593;
assign w8230 = (~w8228 & w7782) | (~w8228 & w40594) | (w7782 & w40594);
assign w8231 = ~w8224 & ~w7923;
assign w8232 = (w8231 & w7782) | (w8231 & w40595) | (w7782 & w40595);
assign w8233 = w8230 & ~w8232;
assign w8234 = a[70] & ~w7315;
assign w8235 = ~w8190 & ~w8234;
assign w8236 = ~w8235 & w7923;
assign w8237 = w7902 & w40596;
assign w8238 = (~w8236 & w7782) | (~w8236 & w40597) | (w7782 & w40597);
assign w8239 = a[70] & ~w7566;
assign w8240 = ~w7568 & ~w8239;
assign w8241 = ~w8240 & ~w7923;
assign w8242 = (w8241 & w7782) | (w8241 & w40598) | (w7782 & w40598);
assign w8243 = w8238 & ~w8242;
assign w8244 = w8233 & w8243;
assign w8245 = ~w6264 & w7568;
assign w8246 = w8195 & w8245;
assign w8247 = (w44344 & w50294) | (w44344 & w50295) | (w50294 & w50295);
assign w8248 = ~w6769 & ~w8247;
assign w8249 = ~w8244 & ~w8248;
assign w8250 = w8196 & ~w7923;
assign w8251 = ~w8192 & w52214;
assign w8252 = ~w8204 & ~w8208;
assign w8253 = ~w7904 & w8252;
assign w8254 = ~w8251 & ~w8253;
assign w8255 = w8202 & ~w7923;
assign w8256 = (w8255 & w7782) | (w8255 & w40601) | (w7782 & w40601);
assign w8257 = ~w8213 & w8256;
assign w8258 = ~w7314 & w52215;
assign w8259 = ~w8200 & ~w8258;
assign w8260 = w8259 & ~w7923;
assign w8261 = w8191 & w52216;
assign w8262 = ~w8257 & ~w8261;
assign w8263 = ~w8254 & w8262;
assign w8264 = ~a[69] & ~w8221;
assign w8265 = ~w8238 & ~w8264;
assign w8266 = (w6737 & w51929) | (w6737 & w51930) | (w51929 & w51930);
assign w8267 = a[69] & a[70];
assign w8268 = (w8267 & w8221) | (w8267 & w51931) | (w8221 & w51931);
assign w8269 = ~w7568 & ~w8268;
assign w8270 = ~w8269 & ~w7923;
assign w8271 = w6264 & w52217;
assign w8272 = w7544 & w8225;
assign w8273 = (~w8272 & w8265) | (~w8272 & w51932) | (w8265 & w51932);
assign w8274 = ~w8217 & w8249;
assign w8275 = w8263 & w8273;
assign w8276 = ~w8274 & ~w8275;
assign w8277 = ~w8233 & ~w8243;
assign w8278 = ~w6264 & w8277;
assign w8279 = ~a[71] & w8190;
assign w8280 = ~a[71] & w7315;
assign w8281 = w7579 & ~w8280;
assign w8282 = ~w8279 & ~w8281;
assign w8283 = (~w8197 & ~w8282) | (~w8197 & w51933) | (~w8282 & w51933);
assign w8284 = w6264 & ~w8283;
assign w8285 = ~w6264 & w8283;
assign w8286 = ~w8284 & ~w8285;
assign w8287 = w8286 & ~w7923;
assign w8288 = ~w6769 & ~w7315;
assign w8289 = (a[72] & w8279) | (a[72] & w51934) | (w8279 & w51934);
assign w8290 = ~w8279 & w51935;
assign w8291 = ~w8289 & ~w8290;
assign w8292 = (~w44364 & w47224) | (~w44364 & w47225) | (w47224 & w47225);
assign w8293 = (w7782 & w49605) | (w7782 & w49606) | (w49605 & w49606);
assign w8294 = w8292 & ~w8293;
assign w8295 = (~w8294 & ~w8277) | (~w8294 & w49607) | (~w8277 & w49607);
assign w8296 = ~w7590 & w7600;
assign w8297 = (~w40541 & w44365) | (~w40541 & w44366) | (w44365 & w44366);
assign w8298 = ~w5330 & w7562;
assign w8299 = w8298 & w52218;
assign w8300 = ~w5330 & ~w7562;
assign w8301 = (w7782 & w44367) | (w7782 & w44368) | (w44367 & w44368);
assign w8302 = ~w8299 & ~w8301;
assign w8303 = ~w8278 & w44369;
assign w8304 = ~w8275 & w44370;
assign w8305 = ~w7648 & ~w7668;
assign w8306 = w7902 & w40606;
assign w8307 = w4056 & w7923;
assign w8308 = (~w8307 & w7782) | (~w8307 & w40607) | (w7782 & w40607);
assign w8309 = w8305 & ~w7923;
assign w8310 = (w8309 & w7782) | (w8309 & w40608) | (w7782 & w40608);
assign w8311 = w8308 & ~w8310;
assign w8312 = w7694 & ~w7724;
assign w8313 = w8311 & ~w8312;
assign w8314 = ~w8311 & w8312;
assign w8315 = ~w8313 & ~w8314;
assign w8316 = ~w3646 & w8315;
assign w8317 = ~w7648 & w51936;
assign w8318 = ~w7724 & ~w8317;
assign w8319 = (w44344 & w50296) | (w44344 & w50297) | (w50296 & w50297);
assign w8320 = w40610 & ~w7904;
assign w8321 = ~w8319 & ~w8320;
assign w8322 = w7682 & w7733;
assign w8323 = ~w3242 & ~w8322;
assign w8324 = w8321 & w8323;
assign w8325 = ~w3242 & w8322;
assign w8326 = ~w8321 & w8325;
assign w8327 = ~w8324 & ~w8326;
assign w8328 = ~w8316 & w8327;
assign w8329 = w7562 & w52218;
assign w8330 = (w7782 & w44371) | (w7782 & w44372) | (w44371 & w44372);
assign w8331 = ~w8329 & ~w8330;
assign w8332 = w5330 & w8331;
assign w8333 = ~w5745 & ~w8291;
assign w8334 = (~w7782 & w44373) | (~w7782 & w44374) | (w44373 & w44374);
assign w8335 = ~w5745 & w8291;
assign w8336 = (w7782 & w44375) | (w7782 & w44376) | (w44375 & w44376);
assign w8337 = ~w8334 & ~w8336;
assign w8338 = w8302 & ~w8337;
assign w8339 = ~w8332 & ~w8338;
assign w8340 = (w7657 & w7613) | (w7657 & w51937) | (w7613 & w51937);
assign w8341 = w4430 & ~w8340;
assign w8342 = ~w4430 & w8340;
assign w8343 = ~w8341 & ~w8342;
assign w8344 = ~w8343 & ~w7923;
assign w8345 = (w6873 & w7305) | (w6873 & w51938) | (w7305 & w51938);
assign w8346 = ~w7305 & w51939;
assign w8347 = ~w8345 & ~w8346;
assign w8348 = w4056 & w8347;
assign w8349 = (~w7782 & w51940) | (~w7782 & w51941) | (w51940 & w51941);
assign w8350 = w4056 & ~w8347;
assign w8351 = (w7782 & w51942) | (w7782 & w51943) | (w51942 & w51943);
assign w8352 = ~w8349 & ~w8351;
assign w8353 = ~w7613 & w51944;
assign w8354 = (w4838 & w7613) | (w4838 & w51945) | (w7613 & w51945);
assign w8355 = ~w8353 & ~w8354;
assign w8356 = ~w8355 & ~w7923;
assign w8357 = (w6895 & w7305) | (w6895 & w51946) | (w7305 & w51946);
assign w8358 = ~w7305 & w51947;
assign w8359 = ~w8357 & ~w8358;
assign w8360 = w4430 & ~w8359;
assign w8361 = (~w7782 & w44377) | (~w7782 & w44378) | (w44377 & w44378);
assign w8362 = w4430 & w8359;
assign w8363 = (w7782 & w44379) | (w7782 & w44380) | (w44379 & w44380);
assign w8364 = ~w8361 & ~w8363;
assign w8365 = w8352 & w8364;
assign w8366 = ~w7591 & w7600;
assign w8367 = w7611 & w7622;
assign w8368 = w8366 & ~w8367;
assign w8369 = ~w8366 & w8367;
assign w8370 = ~w8368 & ~w8369;
assign w8371 = (w6845 & w7305) | (w6845 & w51948) | (w7305 & w51948);
assign w8372 = ~w7305 & w51949;
assign w8373 = ~w8371 & ~w8372;
assign w8374 = ~w8373 & w7923;
assign w8375 = w7902 & w40613;
assign w8376 = (~w8374 & w7782) | (~w8374 & w40614) | (w7782 & w40614);
assign w8377 = w8370 & ~w7923;
assign w8378 = (w8377 & w7782) | (w8377 & w40615) | (w7782 & w40615);
assign w8379 = w8376 & ~w8378;
assign w8380 = ~w4838 & w8379;
assign w8381 = ~w4430 & ~w8359;
assign w8382 = (w7782 & w44381) | (w7782 & w44382) | (w44381 & w44382);
assign w8383 = ~w4430 & w8359;
assign w8384 = (~w7782 & w44383) | (~w7782 & w44384) | (w44383 & w44384);
assign w8385 = ~w8382 & ~w8384;
assign w8386 = w8380 & w8385;
assign w8387 = w8365 & ~w8386;
assign w8388 = w8339 & w8387;
assign w8389 = w8328 & w8388;
assign w8390 = ~w8304 & w8389;
assign w8391 = w4838 & ~w8379;
assign w8392 = w8385 & ~w8391;
assign w8393 = w8365 & ~w8392;
assign w8394 = w3646 & ~w8312;
assign w8395 = w8311 & w8394;
assign w8396 = w3646 & w8312;
assign w8397 = ~w8311 & w8396;
assign w8398 = ~w8395 & ~w8397;
assign w8399 = (~w4056 & w44385) | (~w4056 & w52219) | (w44385 & w52219);
assign w8400 = w8347 & w52219;
assign w8401 = w8399 & ~w8400;
assign w8402 = w8398 & ~w8401;
assign w8403 = ~w8393 & w8402;
assign w8404 = w8328 & ~w8403;
assign w8405 = (~w8404 & w8304) | (~w8404 & w40616) | (w8304 & w40616);
assign w8406 = ~w7695 & w7733;
assign w8407 = ~w7763 & ~w8406;
assign w8408 = w7749 & ~w8407;
assign w8409 = w7734 & w7749;
assign w8410 = (w8409 & w7648) | (w8409 & w40617) | (w7648 & w40617);
assign w8411 = ~w8408 & ~w8410;
assign w8412 = w2896 & w8411;
assign w8413 = (w7713 & ~w8411) | (w7713 & w51950) | (~w8411 & w51950);
assign w8414 = ~w2896 & ~w8411;
assign w8415 = ~w7923 & w51951;
assign w8416 = ~w7904 & w8415;
assign w8417 = (~w2558 & w7894) | (~w2558 & w51952) | (w7894 & w51952);
assign w8418 = (w8417 & w7887) | (w8417 & w51953) | (w7887 & w51953);
assign w8419 = ~w7842 & w51954;
assign w8420 = ~w2558 & w7923;
assign w8421 = (~w8420 & w7782) | (~w8420 & w40618) | (w7782 & w40618);
assign w8422 = ~w8416 & w8421;
assign w8423 = ~w7708 & w7769;
assign w8424 = (~w2285 & ~w7769) | (~w2285 & w51955) | (~w7769 & w51955);
assign w8425 = ~w8416 & w40619;
assign w8426 = w7769 & w51956;
assign w8427 = (w8426 & w8416) | (w8426 & w40620) | (w8416 & w40620);
assign w8428 = ~w8425 & ~w8427;
assign w8429 = ~w7765 & w7769;
assign w8430 = ~w7759 & w8429;
assign w8431 = ~w2285 & w7923;
assign w8432 = w7902 & w40621;
assign w8433 = (~w8431 & w7782) | (~w8431 & w40622) | (w7782 & w40622);
assign w8434 = ~w7923 & ~w8430;
assign w8435 = (w8434 & w7782) | (w8434 & w40623) | (w7782 & w40623);
assign w8436 = w8433 & ~w8435;
assign w8437 = w7482 & w7774;
assign w8438 = ~w2006 & ~w8437;
assign w8439 = ~w8436 & w8438;
assign w8440 = ~w2006 & w8437;
assign w8441 = w8436 & w8440;
assign w8442 = ~w8439 & ~w8441;
assign w8443 = w8428 & w8442;
assign w8444 = (w2285 & ~w7769) | (w2285 & w51957) | (~w7769 & w51957);
assign w8445 = (w8444 & w8416) | (w8444 & w40624) | (w8416 & w40624);
assign w8446 = w7769 & w51958;
assign w8447 = ~w8416 & w40625;
assign w8448 = ~w8445 & ~w8447;
assign w8449 = (w7734 & w7648) | (w7734 & w40626) | (w7648 & w40626);
assign w8450 = ~w8449 & w51959;
assign w8451 = (w3242 & w8449) | (w3242 & w51960) | (w8449 & w51960);
assign w8452 = ~w8450 & ~w8451;
assign w8453 = w7902 & w40627;
assign w8454 = ~w7923 & w51961;
assign w8455 = ~w7904 & w8454;
assign w8456 = (~w7762 & w7923) | (~w7762 & w51962) | (w7923 & w51962);
assign w8457 = (~w8456 & w7782) | (~w8456 & w52084) | (w7782 & w52084);
assign w8458 = ~w8455 & w8457;
assign w8459 = ~w8412 & ~w8414;
assign w8460 = ~w7923 & w8459;
assign w8461 = w2558 & ~w7713;
assign w8462 = w8460 & w8461;
assign w8463 = ~w7904 & w8462;
assign w8464 = w2558 & w7713;
assign w8465 = ~w8460 & w8464;
assign w8466 = w7902 & w40628;
assign w8467 = ~w7782 & w8466;
assign w8468 = ~w8465 & ~w8467;
assign w8469 = ~w8463 & w8468;
assign w8470 = w8458 & w8469;
assign w8471 = ~w2558 & w7713;
assign w8472 = w8460 & w8471;
assign w8473 = ~w7904 & w8472;
assign w8474 = ~w2558 & ~w7713;
assign w8475 = ~w8460 & w8474;
assign w8476 = w7902 & w40629;
assign w8477 = ~w7782 & w8476;
assign w8478 = ~w8475 & ~w8477;
assign w8479 = ~w8473 & w8478;
assign w8480 = (~w7713 & ~w8411) | (~w7713 & w51963) | (~w8411 & w51963);
assign w8481 = ~w2558 & ~w8411;
assign w8482 = w8480 & ~w8481;
assign w8483 = w2558 & w8411;
assign w8484 = ~w8414 & ~w8483;
assign w8485 = ~w7923 & w8484;
assign w8486 = (~w3277 & w7713) | (~w3277 & w51964) | (w7713 & w51964);
assign w8487 = ~w8485 & w8486;
assign w8488 = w7902 & w40630;
assign w8489 = ~w7782 & w8488;
assign w8490 = ~w8487 & ~w8489;
assign w8491 = ~w7923 & w8482;
assign w8492 = ~w7904 & w8491;
assign w8493 = w8490 & ~w8492;
assign w8494 = w8479 & ~w8493;
assign w8495 = ~w8470 & w8494;
assign w8496 = w8448 & w8495;
assign w8497 = w8443 & ~w8496;
assign w8498 = w7496 & w7502;
assign w8499 = (w7482 & w7759) | (w7482 & w40631) | (w7759 & w40631);
assign w8500 = w8498 & ~w8499;
assign w8501 = ~w8498 & w8499;
assign w8502 = ~w8500 & ~w8501;
assign w8503 = w7490 & ~w7491;
assign w8504 = ~w7490 & w7491;
assign w8505 = ~w8503 & ~w8504;
assign w8506 = w7902 & w40632;
assign w8507 = w8505 & w7923;
assign w8508 = (~w8507 & w7782) | (~w8507 & w40633) | (w7782 & w40633);
assign w8509 = ~w7923 & w8502;
assign w8510 = ~w7904 & w8509;
assign w8511 = w8508 & ~w8510;
assign w8512 = (w1738 & w8510) | (w1738 & w40634) | (w8510 & w40634);
assign w8513 = w2006 & w8437;
assign w8514 = ~w8436 & w8513;
assign w8515 = w2006 & ~w8437;
assign w8516 = w8436 & w8515;
assign w8517 = ~w8514 & ~w8516;
assign w8518 = ~w8512 & w8517;
assign w8519 = (w8518 & w8496) | (w8518 & w40648) | (w8496 & w40648);
assign w8520 = ~w8510 & w40635;
assign w8521 = w8437 & w8498;
assign w8522 = w7517 & ~w7523;
assign w8523 = w8521 & w8522;
assign w8524 = w7519 & ~w7523;
assign w8525 = (~w8524 & ~w8430) | (~w8524 & w40636) | (~w8430 & w40636);
assign w8526 = ~w7923 & w8525;
assign w8527 = (~w8522 & w7497) | (~w8522 & w51965) | (w7497 & w51965);
assign w8528 = (w8527 & ~w40637) | (w8527 & w49608) | (~w40637 & w49608);
assign w8529 = w7887 & w51966;
assign w8530 = ~w7910 & w52220;
assign w8531 = ~w1541 & ~w8530;
assign w8532 = (w8531 & ~w8103) | (w8531 & w51968) | (~w8103 & w51968);
assign w8533 = w8526 & ~w8528;
assign w8534 = ~w7904 & w8533;
assign w8535 = w8532 & ~w8534;
assign w8536 = ~w8520 & ~w8535;
assign w8537 = (w3242 & ~w8321) | (w3242 & w51969) | (~w8321 & w51969);
assign w8538 = ~w8321 & w8322;
assign w8539 = w8537 & ~w8538;
assign w8540 = w8536 & ~w8539;
assign w8541 = ~w8519 & w8540;
assign w8542 = w8405 & w8541;
assign w8543 = ~w8479 & w8493;
assign w8544 = w8478 & w44386;
assign w8545 = w8470 & ~w8544;
assign w8546 = w8448 & ~w8545;
assign w8547 = ~w7519 & ~w7523;
assign w8548 = (w8547 & ~w8430) | (w8547 & w40638) | (~w8430 & w40638);
assign w8549 = ~w7468 & ~w7525;
assign w8550 = ~w8548 & ~w8549;
assign w8551 = ~w7780 & w40639;
assign w8552 = ~w7923 & ~w8551;
assign w8553 = ~w8550 & w8552;
assign w8554 = ~w7904 & w8553;
assign w8555 = w7902 & w40640;
assign w8556 = w7524 & w7923;
assign w8557 = w1320 & ~w8556;
assign w8558 = (w8557 & w7782) | (w8557 & w49609) | (w7782 & w49609);
assign w8559 = ~w8554 & w8558;
assign w8560 = w1541 & ~w8528;
assign w8561 = w8526 & w8560;
assign w8562 = ~w7904 & w8561;
assign w8563 = w7887 & w51970;
assign w8564 = ~w7842 & w51971;
assign w8565 = (w8564 & w7543) | (w8564 & w51972) | (w7543 & w51972);
assign w8566 = w1541 & w8530;
assign w8567 = ~w8565 & ~w8566;
assign w8568 = ~w8562 & w8567;
assign w8569 = ~w8559 & w8568;
assign w8570 = ~w8536 & w8569;
assign w8571 = w8443 & ~w8570;
assign w8572 = ~w8545 & w40641;
assign w8573 = w8571 & ~w8572;
assign w8574 = ~w8512 & w8569;
assign w8575 = w8517 & w8574;
assign w8576 = ~w8570 & ~w8575;
assign w8577 = ~w8573 & ~w8576;
assign w8578 = ~w945 & w8018;
assign w8579 = ~w1344 & ~w8018;
assign w8580 = ~w8578 & ~w8579;
assign w8581 = ~w8573 & w51973;
assign w8582 = (w8581 & ~w8405) | (w8581 & w51974) | (~w8405 & w51974);
assign w8583 = (~w8556 & w7782) | (~w8556 & w40642) | (w7782 & w40642);
assign w8584 = ~w8554 & w8583;
assign w8585 = (~w1320 & w8554) | (~w1320 & w40643) | (w8554 & w40643);
assign w8586 = w1120 & w7932;
assign w8587 = (w8586 & w7904) | (w8586 & w40644) | (w7904 & w40644);
assign w8588 = w1120 & ~w7932;
assign w8589 = ~w7904 & w40645;
assign w8590 = ~w8587 & ~w8589;
assign w8591 = ~w8585 & w8590;
assign w8592 = w8033 & w8591;
assign w8593 = w8028 & w8592;
assign w8594 = ~w8014 & w8593;
assign w8595 = w8155 & w8594;
assign w8596 = ~w8101 & w8595;
assign w8597 = w8188 & ~w8596;
assign w8598 = ~w8157 & w8597;
assign w8599 = ~w8573 & w51975;
assign w8600 = ~w8585 & w51976;
assign w8601 = ~w8580 & ~w8591;
assign w8602 = ~w8600 & ~w8601;
assign w8603 = ~w8599 & ~w8602;
assign w8604 = ~w8519 & w51977;
assign w8605 = w8405 & w8604;
assign w8606 = ~w8603 & ~w8605;
assign w8607 = w8598 & ~w8606;
assign w8608 = (w7945 & w8607) | (w7945 & w40646) | (w8607 & w40646);
assign w8609 = ~w8607 & w40647;
assign w8610 = ~w8608 & ~w8609;
assign w8611 = w754 & w8610;
assign w8612 = ~w8559 & ~w8585;
assign w8613 = ~w8443 & w8517;
assign w8614 = w8517 & ~w8543;
assign w8615 = w8546 & w8614;
assign w8616 = ~w8613 & ~w8615;
assign w8617 = w8536 & w52221;
assign w8618 = ~w1320 & w52222;
assign w8619 = ~w8018 & ~w8618;
assign w8620 = (~w8619 & w8542) | (~w8619 & w51979) | (w8542 & w51979);
assign w8621 = (w8577 & ~w8405) | (w8577 & w44388) | (~w8405 & w44388);
assign w8622 = w8189 & w8621;
assign w8623 = ~w1120 & ~w8585;
assign w8624 = w8597 & w40649;
assign w8625 = ~w8622 & ~w8624;
assign w8626 = ~w8620 & ~w8625;
assign w8627 = (w8018 & ~w47226) | (w8018 & w49610) | (~w47226 & w49610);
assign w8628 = ~w8019 & w8590;
assign w8629 = w8621 & w8628;
assign w8630 = w8018 & ~w8189;
assign w8631 = w8629 & ~w8630;
assign w8632 = (~w8631 & w8626) | (~w8631 & w47227) | (w8626 & w47227);
assign w8633 = ~w945 & ~w8632;
assign w8634 = (~w8584 & ~w8189) | (~w8584 & w47228) | (~w8189 & w47228);
assign w8635 = ~w8189 & ~w8584;
assign w8636 = ~w8542 & w44389;
assign w8637 = (w8612 & w8542) | (w8612 & w44390) | (w8542 & w44390);
assign w8638 = ~w8636 & ~w8637;
assign w8639 = ~w8635 & w8638;
assign w8640 = (~w8585 & ~w8597) | (~w8585 & w49611) | (~w8597 & w49611);
assign w8641 = ~w8634 & w8640;
assign w8642 = ~w8639 & ~w8641;
assign w8643 = ~w1120 & ~w8642;
assign w8644 = w8596 & ~w8621;
assign w8645 = ~w8404 & ~w8539;
assign w8646 = ~w8520 & w52221;
assign w8647 = ~w8496 & w44391;
assign w8648 = (~w8646 & ~w40650) | (~w8646 & w51980) | (~w40650 & w51980);
assign w8649 = (~w1541 & ~w8597) | (~w1541 & w40651) | (~w8597 & w40651);
assign w8650 = ~w8622 & w8649;
assign w8651 = w8189 & w8648;
assign w8652 = ~w8644 & w8651;
assign w8653 = ~w8650 & ~w8652;
assign w8654 = ~w8535 & w8568;
assign w8655 = w1320 & w8654;
assign w8656 = (w8655 & w8652) | (w8655 & w44392) | (w8652 & w44392);
assign w8657 = w1320 & ~w8654;
assign w8658 = ~w8652 & w44393;
assign w8659 = ~w8656 & ~w8658;
assign w8660 = ~w8643 & w8659;
assign w8661 = ~w1320 & ~w8654;
assign w8662 = (w8661 & w8652) | (w8661 & w44394) | (w8652 & w44394);
assign w8663 = ~w1320 & w8654;
assign w8664 = ~w8652 & w44395;
assign w8665 = ~w8662 & ~w8664;
assign w8666 = w8189 & ~w8644;
assign w8667 = ~w8512 & ~w8520;
assign w8668 = (~w8616 & ~w40652) | (~w8616 & w44396) | (~w40652 & w44396);
assign w8669 = w8667 & ~w8668;
assign w8670 = ~w8667 & w8668;
assign w8671 = ~w8669 & ~w8670;
assign w8672 = (w8511 & w8644) | (w8511 & w49612) | (w8644 & w49612);
assign w8673 = w8666 & ~w8671;
assign w8674 = ~w8672 & ~w8673;
assign w8675 = (~w1541 & w8673) | (~w1541 & w49613) | (w8673 & w49613);
assign w8676 = w8665 & ~w8675;
assign w8677 = w8660 & ~w8676;
assign w8678 = w1120 & w8642;
assign w8679 = w945 & w8632;
assign w8680 = ~w8678 & ~w8679;
assign w8681 = ~w8677 & w8680;
assign w8682 = ~w8545 & w44397;
assign w8683 = (w8428 & ~w8495) | (w8428 & w44398) | (~w8495 & w44398);
assign w8684 = w8683 & w50184;
assign w8685 = w8189 & w8684;
assign w8686 = (~w2896 & w8390) | (~w2896 & w40654) | (w8390 & w40654);
assign w8687 = w2896 & ~w8539;
assign w8688 = ~w8404 & w8687;
assign w8689 = ~w8390 & w8688;
assign w8690 = (~w8458 & w8390) | (~w8458 & w40655) | (w8390 & w40655);
assign w8691 = ~w8686 & ~w8690;
assign w8692 = (w8479 & ~w8691) | (w8479 & w51981) | (~w8691 & w51981);
assign w8693 = (w8428 & ~w8685) | (w8428 & w47229) | (~w8685 & w47229);
assign w8694 = w8692 & ~w8693;
assign w8695 = w8685 & w47230;
assign w8696 = w8422 & ~w8423;
assign w8697 = ~w8422 & w8423;
assign w8698 = ~w8696 & ~w8697;
assign w8699 = (~w8698 & ~w8597) | (~w8698 & w40656) | (~w8597 & w40656);
assign w8700 = ~w8622 & w8699;
assign w8701 = w2006 & ~w8700;
assign w8702 = ~w8695 & w8701;
assign w8703 = ~w8694 & w8702;
assign w8704 = w8436 & ~w8437;
assign w8705 = ~w8436 & w8437;
assign w8706 = ~w8704 & ~w8705;
assign w8707 = ~w8470 & ~w8493;
assign w8708 = (w8428 & ~w8707) | (w8428 & w44398) | (~w8707 & w44398);
assign w8709 = w8682 & w8708;
assign w8710 = w8442 & w8517;
assign w8711 = w8708 & ~w8710;
assign w8712 = ~w8708 & w8710;
assign w8713 = ~w8711 & ~w8712;
assign w8714 = (w40657 & w44399) | (w40657 & w44400) | (w44399 & w44400);
assign w8715 = (~w40657 & w44401) | (~w40657 & w44402) | (w44401 & w44402);
assign w8716 = ~w8714 & ~w8715;
assign w8717 = w1738 & ~w8716;
assign w8718 = w8666 & w8717;
assign w8719 = w1738 & ~w8706;
assign w8720 = (w8719 & w8644) | (w8719 & w49614) | (w8644 & w49614);
assign w8721 = ~w8718 & ~w8720;
assign w8722 = (w8721 & ~w8702) | (w8721 & w47231) | (~w8702 & w47231);
assign w8723 = (w47216 & w51982) | (w47216 & w51983) | (w51982 & w51983);
assign w8724 = w7713 & ~w8723;
assign w8725 = ~w7713 & w8723;
assign w8726 = ~w8724 & ~w8725;
assign w8727 = (w8726 & ~w8597) | (w8726 & w40658) | (~w8597 & w40658);
assign w8728 = ~w8622 & w8727;
assign w8729 = w8469 & w8479;
assign w8730 = ~w8690 & w44403;
assign w8731 = (w8729 & w8690) | (w8729 & w44404) | (w8690 & w44404);
assign w8732 = ~w8730 & ~w8731;
assign w8733 = w8666 & ~w8732;
assign w8734 = ~w8728 & ~w8733;
assign w8735 = (w2285 & w8733) | (w2285 & w49615) | (w8733 & w49615);
assign w8736 = ~w2285 & ~w8728;
assign w8737 = ~w8733 & w8736;
assign w8738 = ~w8686 & ~w8689;
assign w8739 = w8189 & w8738;
assign w8740 = ~w8644 & w8739;
assign w8741 = (w2558 & ~w8457) | (w2558 & w51984) | (~w8457 & w51984);
assign w8742 = (w8741 & ~w8739) | (w8741 & w47232) | (~w8739 & w47232);
assign w8743 = w8457 & w51985;
assign w8744 = w8739 & w47233;
assign w8745 = ~w8742 & ~w8744;
assign w8746 = ~w8737 & w8745;
assign w8747 = ~w8735 & ~w8746;
assign w8748 = (w8706 & w8644) | (w8706 & w51986) | (w8644 & w51986);
assign w8749 = w8666 & w8716;
assign w8750 = ~w8748 & ~w8749;
assign w8751 = (~w1738 & w8749) | (~w1738 & w51987) | (w8749 & w51987);
assign w8752 = ~w8695 & ~w8700;
assign w8753 = ~w8694 & w8752;
assign w8754 = ~w8718 & w49616;
assign w8755 = ~w8753 & w8754;
assign w8756 = ~w8751 & ~w8755;
assign w8757 = w8722 & w8747;
assign w8758 = w8756 & ~w8757;
assign w8759 = ~w8673 & w49617;
assign w8760 = w8665 & w8759;
assign w8761 = w8660 & ~w8760;
assign w8762 = (~w8633 & w8677) | (~w8633 & w51988) | (w8677 & w51988);
assign w8763 = ~w8633 & w8761;
assign w8764 = ~w8758 & w8763;
assign w8765 = ~w8762 & ~w8764;
assign w8766 = w8302 & ~w8332;
assign w8767 = ~w8275 & w40659;
assign w8768 = (w8337 & ~w40659) | (w8337 & w51989) | (~w40659 & w51989);
assign w8769 = w8766 & ~w8768;
assign w8770 = ~w8766 & w8768;
assign w8771 = ~w8769 & ~w8770;
assign w8772 = (~w8331 & w8644) | (~w8331 & w49618) | (w8644 & w49618);
assign w8773 = ~w8644 & w49619;
assign w8774 = ~w8772 & ~w8773;
assign w8775 = ~w4838 & w8774;
assign w8776 = w4838 & ~w8774;
assign w8777 = w8276 & ~w8278;
assign w8778 = ~w8157 & w47234;
assign w8779 = (w5745 & w8157) | (w5745 & w47235) | (w8157 & w47235);
assign w8780 = w8595 & w49620;
assign w8781 = ~w8621 & w8780;
assign w8782 = ~w8779 & ~w8781;
assign w8783 = ~w8644 & w8778;
assign w8784 = w8782 & ~w8783;
assign w8785 = ~w8294 & w8337;
assign w8786 = w5330 & w8785;
assign w8787 = ~w8784 & w8786;
assign w8788 = w5330 & ~w8785;
assign w8789 = w8784 & w8788;
assign w8790 = ~w8787 & ~w8789;
assign w8791 = (~w8775 & w8790) | (~w8775 & w49621) | (w8790 & w49621);
assign w8792 = w8339 & ~w8380;
assign w8793 = w8364 & w8385;
assign w8794 = (w44406 & w47236) | (w44406 & w47237) | (w47236 & w47237);
assign w8795 = (~w44406 & w47238) | (~w44406 & w47239) | (w47238 & w47239);
assign w8796 = ~w8794 & ~w8795;
assign w8797 = (w7782 & w51990) | (w7782 & w51991) | (w51990 & w51991);
assign w8798 = w8359 & w52223;
assign w8799 = ~w8797 & ~w8798;
assign w8800 = (w8799 & ~w8597) | (w8799 & w40660) | (~w8597 & w40660);
assign w8801 = ~w8622 & w8800;
assign w8802 = w8189 & ~w8796;
assign w8803 = ~w8644 & w8802;
assign w8804 = ~w8801 & ~w8803;
assign w8805 = w4056 & ~w8804;
assign w8806 = (w8339 & ~w44370) | (w8339 & w51992) | (~w44370 & w51992);
assign w8807 = ~w4838 & w8806;
assign w8808 = w4838 & ~w8806;
assign w8809 = ~w8807 & ~w8808;
assign w8810 = w8189 & ~w8809;
assign w8811 = (w8379 & ~w8810) | (w8379 & w47240) | (~w8810 & w47240);
assign w8812 = w8810 & w47241;
assign w8813 = ~w8811 & ~w8812;
assign w8814 = w4430 & ~w8813;
assign w8815 = ~w4056 & w8804;
assign w8816 = (w44406 & w47242) | (w44406 & w47243) | (w47242 & w47243);
assign w8817 = w8364 & ~w8816;
assign w8818 = (w4056 & w8157) | (w4056 & w47244) | (w8157 & w47244);
assign w8819 = w8595 & w51993;
assign w8820 = ~w8621 & w8819;
assign w8821 = w8189 & ~w8817;
assign w8822 = ~w8644 & w8821;
assign w8823 = w8352 & ~w8401;
assign w8824 = w3646 & ~w8823;
assign w8825 = ~w8822 & w47245;
assign w8826 = w3646 & w8823;
assign w8827 = (w8826 & w8822) | (w8826 & w47246) | (w8822 & w47246);
assign w8828 = ~w8825 & ~w8827;
assign w8829 = ~w8815 & w8828;
assign w8830 = ~w8805 & ~w8814;
assign w8831 = w8829 & ~w8830;
assign w8832 = (w8315 & w8644) | (w8315 & w49622) | (w8644 & w49622);
assign w8833 = ~w8386 & w51994;
assign w8834 = (~w8833 & w8767) | (~w8833 & w44407) | (w8767 & w44407);
assign w8835 = w8403 & w8834;
assign w8836 = w8352 & ~w8385;
assign w8837 = w8806 & w8836;
assign w8838 = w8835 & ~w8837;
assign w8839 = w8189 & ~w8838;
assign w8840 = (~w8316 & ~w8839) | (~w8316 & w47247) | (~w8839 & w47247);
assign w8841 = (~w8401 & w8392) | (~w8401 & w51995) | (w8392 & w51995);
assign w8842 = ~w8316 & w8398;
assign w8843 = (~w8842 & ~w8834) | (~w8842 & w51996) | (~w8834 & w51996);
assign w8844 = ~w3242 & w8832;
assign w8845 = (w8834 & w51997) | (w8834 & w51998) | (w51997 & w51998);
assign w8846 = ~w8840 & w8845;
assign w8847 = ~w8844 & ~w8846;
assign w8848 = ~w3646 & ~w8823;
assign w8849 = (w8848 & w8822) | (w8848 & w47248) | (w8822 & w47248);
assign w8850 = ~w3646 & w8823;
assign w8851 = ~w8822 & w47249;
assign w8852 = ~w8849 & ~w8851;
assign w8853 = w8847 & w8852;
assign w8854 = w8791 & ~w8831;
assign w8855 = w8853 & w8854;
assign w8856 = ~w4430 & ~w8379;
assign w8857 = (w8856 & ~w8810) | (w8856 & w47250) | (~w8810 & w47250);
assign w8858 = ~w4430 & w8379;
assign w8859 = w8810 & w47251;
assign w8860 = ~w8857 & ~w8859;
assign w8861 = ~w8815 & w8860;
assign w8862 = w8828 & w8861;
assign w8863 = w8853 & ~w8862;
assign w8864 = ~w8831 & w8863;
assign w8865 = ~w8840 & ~w8843;
assign w8866 = w3242 & ~w8832;
assign w8867 = ~w8865 & w8866;
assign w8868 = (~w3242 & ~w8597) | (~w3242 & w40661) | (~w8597 & w40661);
assign w8869 = ~w8622 & w8868;
assign w8870 = (~w8316 & ~w8834) | (~w8316 & w49623) | (~w8834 & w49623);
assign w8871 = w8189 & ~w8870;
assign w8872 = ~w8644 & w8871;
assign w8873 = ~w8869 & ~w8872;
assign w8874 = w8327 & ~w8539;
assign w8875 = ~w2896 & ~w8874;
assign w8876 = w8873 & w8875;
assign w8877 = ~w2896 & w8874;
assign w8878 = ~w8873 & w8877;
assign w8879 = ~w8876 & ~w8878;
assign w8880 = ~w8867 & w8879;
assign w8881 = (w8880 & ~w8863) | (w8880 & w47252) | (~w8863 & w47252);
assign w8882 = ~w8855 & w8881;
assign w8883 = ~a[64] & ~a[65];
assign w8884 = ~a[66] & w8883;
assign w8885 = ~w8884 & ~w7924;
assign w8886 = (~w8218 & ~w8885) | (~w8218 & w51999) | (~w8885 & w51999);
assign w8887 = ~w8157 & w47253;
assign w8888 = ~w8644 & w8887;
assign w8889 = ~a[67] & ~w8885;
assign w8890 = (w47216 & w52000) | (w47216 & w52001) | (w52000 & w52001);
assign w8891 = ~w8889 & ~w8890;
assign w8892 = (~w8891 & w8157) | (~w8891 & w47254) | (w8157 & w47254);
assign w8893 = w8595 & w49624;
assign w8894 = ~w8621 & w8893;
assign w8895 = ~w8892 & ~w8894;
assign w8896 = ~w8888 & w8895;
assign w8897 = w7315 & ~w8896;
assign w8898 = a[68] & ~w8218;
assign w8899 = a[68] & ~w7924;
assign w8900 = (w47216 & w52002) | (w47216 & w52003) | (w52002 & w52003);
assign w8901 = ~w8899 & ~w8900;
assign w8902 = (w8901 & w8644) | (w8901 & w49625) | (w8644 & w49625);
assign w8903 = ~w8220 & ~w8898;
assign w8904 = ~w8644 & w49626;
assign w8905 = ~w8902 & ~w8904;
assign w8906 = ~w8897 & w8905;
assign w8907 = ~w7315 & w8896;
assign w8908 = (~w6769 & ~w8896) | (~w6769 & w8258) | (~w8896 & w8258);
assign w8909 = ~w8906 & w8908;
assign w8910 = (w8900 & w8644) | (w8900 & w49627) | (w8644 & w49627);
assign w8911 = ~w8221 & ~w8225;
assign w8912 = (w47216 & w52004) | (w47216 & w52005) | (w52004 & w52005);
assign w8913 = w8911 & ~w7924;
assign w8914 = ~w8912 & ~w8913;
assign w8915 = ~w8644 & w49628;
assign w8916 = a[69] & w8900;
assign w8917 = ~w8644 & w49629;
assign w8918 = w8916 & ~w8917;
assign w8919 = w8226 & w8915;
assign w8920 = ~w8918 & ~w8919;
assign w8921 = ~w8910 & ~w8915;
assign w8922 = ~a[69] & w8921;
assign w8923 = w8920 & ~w8922;
assign w8924 = ~w8909 & w8923;
assign w8925 = ~w6769 & w8233;
assign w8926 = w6769 & ~w8233;
assign w8927 = ~w8925 & ~w8926;
assign w8928 = ~w8644 & w49630;
assign w8929 = w8243 & ~w8928;
assign w8930 = ~w8243 & w8928;
assign w8931 = ~w8929 & ~w8930;
assign w8932 = ~w6264 & w8931;
assign w8933 = (w6769 & w8896) | (w6769 & w8205) | (w8896 & w8205);
assign w8934 = ~w8905 & ~w8907;
assign w8935 = w8933 & ~w8934;
assign w8936 = ~w8932 & ~w8935;
assign w8937 = ~w8924 & w8936;
assign w8938 = w6769 & ~w8244;
assign w8939 = ~w8273 & ~w8938;
assign w8940 = ~w8244 & w52006;
assign w8941 = ~w8939 & w52007;
assign w8942 = ~w8644 & w49631;
assign w8943 = w8263 & ~w8942;
assign w8944 = ~w8263 & w8942;
assign w8945 = ~w8943 & ~w8944;
assign w8946 = ~w5745 & w8945;
assign w8947 = w6264 & ~w8931;
assign w8948 = ~w8946 & ~w8947;
assign w8949 = ~w8937 & w8948;
assign w8950 = ~w5330 & ~w8785;
assign w8951 = ~w8784 & w8950;
assign w8952 = ~w5330 & w8785;
assign w8953 = w8784 & w8952;
assign w8954 = ~w8951 & ~w8953;
assign w8955 = ~w8776 & w8954;
assign w8956 = (~w8775 & ~w8954) | (~w8775 & w49621) | (~w8954 & w49621);
assign w8957 = w5745 & ~w8945;
assign w8958 = w8880 & ~w8957;
assign w8959 = ~w8956 & w8958;
assign w8960 = ~w8864 & w8959;
assign w8961 = ~w8949 & w8960;
assign w8962 = ~w8882 & ~w8961;
assign w8963 = w8873 & ~w8874;
assign w8964 = ~w8873 & w8874;
assign w8965 = ~w8963 & ~w8964;
assign w8966 = w2896 & w8965;
assign w8967 = w8458 & ~w8740;
assign w8968 = ~w8458 & w8740;
assign w8969 = ~w8967 & ~w8968;
assign w8970 = ~w2558 & ~w8969;
assign w8971 = ~w8966 & ~w8970;
assign w8972 = ~w8966 & w47255;
assign w8973 = w8722 & w8972;
assign w8974 = w8763 & w8973;
assign w8975 = ~w8961 & w47256;
assign w8976 = (~w8611 & w8975) | (~w8611 & w52008) | (w8975 & w52008);
assign w8977 = ~w754 & ~w7945;
assign w8978 = (w8977 & w8607) | (w8977 & w40662) | (w8607 & w40662);
assign w8979 = ~w7944 & w52009;
assign w8980 = ~w8607 & w40663;
assign w8981 = ~w8978 & ~w8980;
assign w8982 = w7988 & w8012;
assign w8983 = w8021 & ~w8591;
assign w8984 = (w8021 & w8575) | (w8021 & w40664) | (w8575 & w40664);
assign w8985 = ~w8573 & w8984;
assign w8986 = w8536 & w8591;
assign w8987 = ~w8539 & w8986;
assign w8988 = ~w8519 & w8987;
assign w8989 = ~w8519 & w44410;
assign w8990 = w8405 & w8989;
assign w8991 = (w8982 & w8990) | (w8982 & w44411) | (w8990 & w44411);
assign w8992 = ~w8990 & w44412;
assign w8993 = ~w8991 & ~w8992;
assign w8994 = w8666 & ~w8993;
assign w8995 = (w7445 & ~w7924) | (w7445 & w52010) | (~w7924 & w52010);
assign w8996 = w7924 & w52011;
assign w8997 = ~w8995 & ~w8996;
assign w8998 = (w8997 & ~w8597) | (w8997 & w40665) | (~w8597 & w40665);
assign w8999 = ~w8622 & w8998;
assign w9000 = w612 & ~w8999;
assign w9001 = ~w8994 & w9000;
assign w9002 = w754 & ~w8610;
assign w9003 = (~w9001 & w8610) | (~w9001 & w44413) | (w8610 & w44413);
assign w9004 = ~w8633 & w9003;
assign w9005 = w8761 & w9004;
assign w9006 = w8973 & w9005;
assign w9007 = w8541 & w8594;
assign w9008 = w8405 & w9007;
assign w9009 = ~w8577 & w8594;
assign w9010 = w7976 & w8173;
assign w9011 = ~w8036 & w9010;
assign w9012 = ~w9009 & w9011;
assign w9013 = ~w9008 & w9012;
assign w9014 = ~w8075 & w8173;
assign w9015 = (w8153 & ~w8173) | (w8153 & w52012) | (~w8173 & w52012);
assign w9016 = w8125 & ~w8182;
assign w9017 = (w9013 & w49632) | (w9013 & w49633) | (w49632 & w49633);
assign w9018 = w9016 & w52224;
assign w9019 = ~w9017 & ~w9018;
assign w9020 = (w8181 & w8644) | (w8181 & w52013) | (w8644 & w52013);
assign w9021 = w8666 & w9019;
assign w9022 = (~w9020 & ~w9019) | (~w9020 & w52014) | (~w9019 & w52014);
assign w9023 = w8178 & w52225;
assign w9024 = (~w8177 & ~w8111) | (~w8177 & w52015) | (~w8111 & w52015);
assign w9025 = (w9013 & w52016) | (w9013 & w52017) | (w52016 & w52017);
assign w9026 = ~w9023 & ~w9025;
assign w9027 = ~w42 & w9026;
assign w9028 = ~w9022 & w9027;
assign w9029 = w8013 & w8027;
assign w9030 = ~w8519 & w44417;
assign w9031 = w8405 & w9030;
assign w9032 = ~w8006 & w8027;
assign w9033 = (~w7971 & w8006) | (~w7971 & w52018) | (w8006 & w52018);
assign w9034 = (w8033 & w9031) | (w8033 & w49634) | (w9031 & w49634);
assign w9035 = (w400 & w8644) | (w400 & w50002) | (w8644 & w50002);
assign w9036 = w8666 & ~w9034;
assign w9037 = w7964 & ~w7974;
assign w9038 = w351 & w9037;
assign w9039 = (w9038 & w9036) | (w9038 & w50003) | (w9036 & w50003);
assign w9040 = w351 & ~w9037;
assign w9041 = ~w9036 & w50004;
assign w9042 = ~w9039 & ~w9041;
assign w9043 = ~w9008 & ~w9009;
assign w9044 = w8037 & ~w8159;
assign w9045 = ~w9008 & w44419;
assign w9046 = ~w351 & w8158;
assign w9047 = ~w9045 & ~w9046;
assign w9048 = w8666 & w9047;
assign w9049 = (~w252 & ~w8597) | (~w252 & w40666) | (~w8597 & w40666);
assign w9050 = ~w8622 & w9049;
assign w9051 = ~w8169 & ~w8170;
assign w9052 = ~w57 & w9051;
assign w9053 = ~w9050 & w9052;
assign w9054 = ~w9048 & w9053;
assign w9055 = ~w57 & ~w9051;
assign w9056 = w9050 & w9055;
assign w9057 = ~w9051 & w52019;
assign w9058 = ~w9045 & w9057;
assign w9059 = w8666 & w9058;
assign w9060 = ~w9056 & ~w9059;
assign w9061 = ~w9054 & w9060;
assign w9062 = w351 & ~w8037;
assign w9063 = ~w351 & w8037;
assign w9064 = ~w9062 & ~w9063;
assign w9065 = (~w351 & w8101) | (~w351 & w47257) | (w8101 & w47257);
assign w9066 = (~w9065 & w9008) | (~w9065 & w44420) | (w9008 & w44420);
assign w9067 = w8189 & ~w9066;
assign w9068 = w9043 & ~w9064;
assign w9069 = w9067 & ~w9068;
assign w9070 = ~w252 & ~w8158;
assign w9071 = ~w9069 & w9070;
assign w9072 = ~w252 & w8158;
assign w9073 = w9069 & w9072;
assign w9074 = ~w9071 & ~w9073;
assign w9075 = w9061 & w9074;
assign w9076 = w8405 & w8988;
assign w9077 = ~w7971 & w8033;
assign w9078 = w9032 & ~w9077;
assign w9079 = ~w8014 & w52020;
assign w9080 = (w9079 & w9076) | (w9079 & w44422) | (w9076 & w44422);
assign w9081 = ~w9032 & w9077;
assign w9082 = ~w9031 & w44423;
assign w9083 = ~w9080 & ~w9082;
assign w9084 = w8666 & w9083;
assign w9085 = (~w7970 & ~w8597) | (~w7970 & w40667) | (~w8597 & w40667);
assign w9086 = ~w8622 & w9085;
assign w9087 = ~w400 & ~w9086;
assign w9088 = ~w9084 & w9087;
assign w9089 = w8005 & w8027;
assign w9090 = ~w7988 & ~w9089;
assign w9091 = w7988 & ~w8013;
assign w9092 = ~w9089 & ~w9091;
assign w9093 = (w9092 & w9076) | (w9092 & w40669) | (w9076 & w40669);
assign w9094 = w8006 & w8027;
assign w9095 = w8006 & w52021;
assign w9096 = (~w9095 & w9076) | (~w9095 & w40671) | (w9076 & w40671);
assign w9097 = ~w9093 & w9096;
assign w9098 = w8666 & w9097;
assign w9099 = w7999 & ~w8000;
assign w9100 = ~w7999 & w8000;
assign w9101 = ~w9099 & ~w9100;
assign w9102 = w493 & w9101;
assign w9103 = (~w9102 & w8644) | (~w9102 & w40673) | (w8644 & w40673);
assign w9104 = ~w9098 & ~w9103;
assign w9105 = ~w9088 & ~w9104;
assign w9106 = w9075 & w47258;
assign w9107 = (w8086 & w8157) | (w8086 & w40674) | (w8157 & w40674);
assign w9108 = w8595 & w40675;
assign w9109 = ~w8621 & w9108;
assign w9110 = ~w9107 & ~w9109;
assign w9111 = ~w9013 & w40676;
assign w9112 = w8666 & w9111;
assign w9113 = (w8142 & w9013) | (w8142 & w40677) | (w9013 & w40677);
assign w9114 = w9110 & ~w9113;
assign w9115 = ~w9112 & w9114;
assign w9116 = ~w8073 & w52022;
assign w9117 = (w9116 & ~w9043) | (w9116 & w52023) | (~w9043 & w52023);
assign w9118 = (w80 & w9115) | (w80 & w40679) | (w9115 & w40679);
assign w9119 = (w80 & w8644) | (w80 & w49635) | (w8644 & w49635);
assign w9120 = w8099 & w8152;
assign w9121 = ~w3 & ~w9120;
assign w9122 = (w9121 & w9112) | (w9121 & w49636) | (w9112 & w49636);
assign w9123 = ~w3 & w9120;
assign w9124 = ~w9112 & w49637;
assign w9125 = ~w9122 & ~w9124;
assign w9126 = ~w9118 & w9125;
assign w9127 = w9004 & w9126;
assign w9128 = w9106 & w9127;
assign w9129 = w9127 & w47259;
assign w9130 = w9006 & w9129;
assign w9131 = w8962 & w9130;
assign w9132 = ~w8681 & w9004;
assign w9133 = ~w8758 & w9005;
assign w9134 = ~w9132 & ~w9133;
assign w9135 = w9129 & ~w9134;
assign w9136 = ~w8994 & ~w8999;
assign w9137 = (~w612 & w8994) | (~w612 & w40680) | (w8994 & w40680);
assign w9138 = (~w9137 & w8981) | (~w9137 & w44424) | (w8981 & w44424);
assign w9139 = (w400 & w9084) | (w400 & w40681) | (w9084 & w40681);
assign w9140 = (~w9101 & w8644) | (~w9101 & w44425) | (w8644 & w44425);
assign w9141 = ~w9098 & ~w9140;
assign w9142 = (~w493 & w9098) | (~w493 & w44426) | (w9098 & w44426);
assign w9143 = ~w9139 & ~w9142;
assign w9144 = w9138 & w9143;
assign w9145 = ~w9105 & ~w9139;
assign w9146 = ~w351 & ~w9037;
assign w9147 = (w9146 & w9036) | (w9146 & w50005) | (w9036 & w50005);
assign w9148 = ~w351 & w9037;
assign w9149 = ~w9036 & w50006;
assign w9150 = ~w9147 & ~w9149;
assign w9151 = (w8158 & ~w9067) | (w8158 & w40682) | (~w9067 & w40682);
assign w9152 = w9067 & w40683;
assign w9153 = ~w9151 & ~w9152;
assign w9154 = w252 & ~w9153;
assign w9155 = w57 & ~w9051;
assign w9156 = ~w9050 & w9155;
assign w9157 = ~w9048 & w9156;
assign w9158 = w57 & w9051;
assign w9159 = w9050 & w9158;
assign w9160 = w9051 & w52024;
assign w9161 = (w9160 & ~w9043) | (w9160 & w40684) | (~w9043 & w40684);
assign w9162 = w8666 & w9161;
assign w9163 = ~w9159 & ~w9162;
assign w9164 = ~w9157 & w9163;
assign w9165 = (w9043 & w52025) | (w9043 & w52026) | (w52025 & w52026);
assign w9166 = ~w9115 & w9165;
assign w9167 = w9164 & ~w9166;
assign w9168 = w9150 & ~w9154;
assign w9169 = w9167 & w9168;
assign w9170 = w9042 & ~w9145;
assign w9171 = ~w9144 & w9170;
assign w9172 = w9169 & ~w9171;
assign w9173 = ~w9075 & w9167;
assign w9174 = w9126 & ~w9173;
assign w9175 = ~w9173 & w47260;
assign w9176 = (w3 & w40685) | (w3 & w52226) | (w40685 & w52226);
assign w9177 = ~w9112 & w52027;
assign w9178 = w9176 & ~w9177;
assign w9179 = ~w9021 & w40686;
assign w9180 = ~w42 & ~w9026;
assign w9181 = w7872 & w52209;
assign w9182 = ~w7872 & ~w7886;
assign w9183 = (w8103 & w52028) | (w8103 & w52029) | (w52028 & w52029);
assign w9184 = ~w9181 & ~w9183;
assign w9185 = w40687 & w52227;
assign w9186 = ~w8178 & ~w9185;
assign w9187 = (w9013 & w52030) | (w9013 & w52031) | (w52030 & w52031);
assign w9188 = ~w9186 & w9187;
assign w9189 = ~w9180 & ~w9188;
assign w9190 = ~w9179 & w9189;
assign w9191 = ~w9028 & w9178;
assign w9192 = w9190 & ~w9191;
assign w9193 = (w9192 & w9172) | (w9192 & w47261) | (w9172 & w47261);
assign w9194 = ~w9135 & w9193;
assign w9195 = ~w9131 & w9194;
assign w9196 = ~w8764 & w52032;
assign w9197 = ~w8975 & w9196;
assign w9198 = ~w754 & ~w8610;
assign w9199 = (~w9198 & w8764) | (~w9198 & w52033) | (w8764 & w52033);
assign w9200 = w8973 & w40689;
assign w9201 = (~w9199 & ~w8962) | (~w9199 & w52034) | (~w8962 & w52034);
assign w9202 = w8765 & ~w9002;
assign w9203 = ~w8975 & w9202;
assign w9204 = w9201 & ~w9203;
assign w9205 = ~w8610 & w9195;
assign w9206 = ~w9204 & ~w9205;
assign w9207 = ~w9195 & w52035;
assign w9208 = w9206 & ~w9207;
assign w9209 = (w612 & ~w9206) | (w612 & w52036) | (~w9206 & w52036);
assign w9210 = w8761 & w8973;
assign w9211 = ~w8961 & w47262;
assign w9212 = ~w8758 & w8761;
assign w9213 = ~w8677 & ~w8678;
assign w9214 = ~w9212 & w9213;
assign w9215 = (w9214 & ~w8962) | (w9214 & w40690) | (~w8962 & w40690);
assign w9216 = ~w945 & w9195;
assign w9217 = ~w9195 & w9215;
assign w9218 = ~w9216 & ~w9217;
assign w9219 = ~w8633 & ~w8679;
assign w9220 = ~w754 & ~w9219;
assign w9221 = w9218 & w9220;
assign w9222 = ~w754 & w9219;
assign w9223 = ~w9218 & w9222;
assign w9224 = ~w9221 & ~w9223;
assign w9225 = w8659 & w8665;
assign w9226 = ~w8759 & w9225;
assign w9227 = w8973 & w9226;
assign w9228 = ~w8961 & w47263;
assign w9229 = ~w8757 & w52037;
assign w9230 = w9226 & ~w9229;
assign w9231 = (w8665 & w9229) | (w8665 & w52038) | (w9229 & w52038);
assign w9232 = ~w9228 & w9231;
assign w9233 = ~w1120 & w9195;
assign w9234 = ~w9195 & w9232;
assign w9235 = ~w9233 & ~w9234;
assign w9236 = ~w8643 & ~w8678;
assign w9237 = w945 & ~w9236;
assign w9238 = w9235 & w9237;
assign w9239 = w945 & w9236;
assign w9240 = ~w9235 & w9239;
assign w9241 = ~w9238 & ~w9240;
assign w9242 = w9224 & w9241;
assign w9243 = w754 & ~w9219;
assign w9244 = ~w9218 & w9243;
assign w9245 = w754 & w9219;
assign w9246 = w9218 & w9245;
assign w9247 = ~w9244 & ~w9246;
assign w9248 = ~w9242 & w9247;
assign w9249 = ~w2006 & ~w8753;
assign w9250 = ~w8703 & ~w8735;
assign w9251 = ~w9249 & ~w9250;
assign w9252 = w8746 & ~w9249;
assign w9253 = (w8961 & w52039) | (w8961 & w52040) | (w52039 & w52040);
assign w9254 = ~w9251 & ~w9253;
assign w9255 = w8721 & ~w8751;
assign w9256 = ~w9195 & w52041;
assign w9257 = ~w9251 & w9255;
assign w9258 = ~w9251 & w52042;
assign w9259 = w8971 & w9257;
assign w9260 = (~w9258 & ~w8962) | (~w9258 & w40692) | (~w8962 & w40692);
assign w9261 = ~w9195 & ~w9260;
assign w9262 = w8750 & w9192;
assign w9263 = (w9262 & w9172) | (w9262 & w52043) | (w9172 & w52043);
assign w9264 = ~w9135 & w9263;
assign w9265 = ~w9131 & w9264;
assign w9266 = ~w9261 & ~w9265;
assign w9267 = ~w9256 & w9266;
assign w9268 = (w1541 & ~w9266) | (w1541 & w52044) | (~w9266 & w52044);
assign w9269 = ~w8961 & w52045;
assign w9270 = (w8961 & w52046) | (w8961 & w52047) | (w52046 & w52047);
assign w9271 = ~w8759 & ~w9270;
assign w9272 = ~w9195 & w52048;
assign w9273 = (~w9230 & ~w8962) | (~w9230 & w40694) | (~w8962 & w40694);
assign w9274 = ~w9195 & ~w9273;
assign w9275 = w8653 & ~w8654;
assign w9276 = ~w8653 & w8654;
assign w9277 = ~w9275 & ~w9276;
assign w9278 = w9192 & ~w9277;
assign w9279 = (w9278 & w9172) | (w9278 & w52049) | (w9172 & w52049);
assign w9280 = ~w9135 & w9279;
assign w9281 = ~w9131 & w9280;
assign w9282 = w1120 & ~w9281;
assign w9283 = ~w9274 & w9282;
assign w9284 = ~w9272 & w9283;
assign w9285 = w8758 & w8973;
assign w9286 = ~w8675 & ~w8759;
assign w9287 = ~w8757 & w52050;
assign w9288 = (w9286 & w8757) | (w9286 & w52051) | (w8757 & w52051);
assign w9289 = ~w9287 & ~w9288;
assign w9290 = w8962 & w40695;
assign w9291 = (~w9289 & ~w8962) | (~w9289 & w40696) | (~w8962 & w40696);
assign w9292 = ~w9290 & ~w9291;
assign w9293 = (~w1320 & ~w9195) | (~w1320 & w40697) | (~w9195 & w40697);
assign w9294 = ~w9195 & ~w9292;
assign w9295 = w9293 & ~w9294;
assign w9296 = ~w9284 & ~w9295;
assign w9297 = ~w9274 & ~w9281;
assign w9298 = ~w9272 & w9297;
assign w9299 = (~w1120 & ~w9297) | (~w1120 & w52052) | (~w9297 & w52052);
assign w9300 = (w1320 & ~w9195) | (w1320 & w40698) | (~w9195 & w40698);
assign w9301 = ~w9195 & w9292;
assign w9302 = w9300 & ~w9301;
assign w9303 = ~w9284 & w9302;
assign w9304 = ~w9299 & ~w9303;
assign w9305 = w9268 & w9296;
assign w9306 = w9304 & ~w9305;
assign w9307 = ~w945 & ~w9236;
assign w9308 = ~w9235 & w9307;
assign w9309 = ~w945 & w9236;
assign w9310 = w9235 & w9309;
assign w9311 = ~w9308 & ~w9310;
assign w9312 = w9247 & w9311;
assign w9313 = w9306 & w9312;
assign w9314 = ~w9248 & ~w9313;
assign w9315 = ~w1541 & ~w9265;
assign w9316 = ~w9261 & w9315;
assign w9317 = ~w9256 & w9316;
assign w9318 = ~w9302 & w9317;
assign w9319 = w9296 & ~w9318;
assign w9320 = w9311 & ~w9319;
assign w9321 = w9306 & w9320;
assign w9322 = ~w8703 & ~w9249;
assign w9323 = (w8961 & w52053) | (w8961 & w52054) | (w52053 & w52054);
assign w9324 = w2006 & w9195;
assign w9325 = ~w9195 & w9323;
assign w9326 = ~w9324 & ~w9325;
assign w9327 = w9322 & ~w9326;
assign w9328 = ~w9322 & w9326;
assign w9329 = ~w9327 & ~w9328;
assign w9330 = ~w1738 & ~w9329;
assign w9331 = w1738 & ~w9322;
assign w9332 = ~w9326 & w9331;
assign w9333 = w1738 & w9322;
assign w9334 = w9326 & w9333;
assign w9335 = ~w9332 & ~w9334;
assign w9336 = ~w8735 & ~w8737;
assign w9337 = (w8961 & w52055) | (w8961 & w52056) | (w52055 & w52056);
assign w9338 = w9336 & ~w9337;
assign w9339 = w8745 & ~w9336;
assign w9340 = (w8961 & w52057) | (w8961 & w52058) | (w52057 & w52058);
assign w9341 = ~w9195 & w52059;
assign w9342 = w8734 & w9195;
assign w9343 = ~w9341 & ~w9342;
assign w9344 = (~w2006 & w9341) | (~w2006 & w40702) | (w9341 & w40702);
assign w9345 = w9335 & w9344;
assign w9346 = ~w9330 & ~w9345;
assign w9347 = w9242 & w9346;
assign w9348 = ~w9321 & w9347;
assign w9349 = ~w9314 & ~w9348;
assign w9350 = ~a[62] & ~a[63];
assign w9351 = ~a[64] & w9350;
assign w9352 = ~w8644 & w52060;
assign w9353 = (~w9351 & w8644) | (~w9351 & w52061) | (w8644 & w52061);
assign w9354 = a[65] & w9353;
assign w9355 = ~a[65] & ~w9353;
assign w9356 = ~w9352 & ~w9355;
assign w9357 = w9192 & w9356;
assign w9358 = (w9357 & w9172) | (w9357 & w52062) | (w9172 & w52062);
assign w9359 = ~w9135 & w9358;
assign w9360 = ~w9131 & w9359;
assign w9361 = ~w9354 & ~w9360;
assign w9362 = w8883 & ~w9352;
assign w9363 = ~w9195 & w9362;
assign w9364 = w9361 & ~w9363;
assign w9365 = ~w7924 & ~w9364;
assign w9366 = (a[66] & w8644) | (a[66] & w52063) | (w8644 & w52063);
assign w9367 = ~w8644 & w52064;
assign w9368 = ~w9366 & ~w9367;
assign w9369 = a[66] & ~w8883;
assign w9370 = w9195 & w9368;
assign w9371 = ~w8884 & ~w9369;
assign w9372 = ~w9195 & w9371;
assign w9373 = ~w9370 & ~w9372;
assign w9374 = w7924 & w9364;
assign w9375 = (~w7315 & ~w9364) | (~w7315 & w40703) | (~w9364 & w40703);
assign w9376 = ~w9365 & ~w9373;
assign w9377 = w9375 & ~w9376;
assign w9378 = (w7924 & w8644) | (w7924 & w52065) | (w8644 & w52065);
assign w9379 = ~w8644 & w52066;
assign w9380 = ~w9378 & ~w9379;
assign w9381 = ~w8884 & ~w9380;
assign w9382 = (a[67] & w9195) | (a[67] & w40704) | (w9195 & w40704);
assign w9383 = ~w9195 & w40705;
assign w9384 = ~w9382 & ~w9383;
assign w9385 = w8883 & w9380;
assign w9386 = ~w9195 & ~w9385;
assign w9387 = ~w8666 & w9195;
assign w9388 = ~a[66] & ~w9378;
assign w9389 = ~w9386 & ~w9387;
assign w9390 = w9388 & w9389;
assign w9391 = w9384 & ~w9390;
assign w9392 = ~w9384 & w9390;
assign w9393 = ~w9391 & ~w9392;
assign w9394 = ~w9377 & ~w9393;
assign w9395 = (w7315 & w9364) | (w7315 & w40706) | (w9364 & w40706);
assign w9396 = w9373 & ~w9374;
assign w9397 = w9395 & ~w9396;
assign w9398 = ~w8932 & ~w8947;
assign w9399 = (w9398 & w8924) | (w9398 & w52067) | (w8924 & w52067);
assign w9400 = ~w8924 & w52068;
assign w9401 = ~w9399 & ~w9400;
assign w9402 = ~w8931 & w9195;
assign w9403 = ~w9195 & ~w9401;
assign w9404 = ~w9402 & ~w9403;
assign w9405 = ~w5745 & ~w9404;
assign w9406 = ~w8909 & ~w8935;
assign w9407 = ~w9195 & w9406;
assign w9408 = w6264 & ~w8923;
assign w9409 = (w9408 & w9195) | (w9408 & w40707) | (w9195 & w40707);
assign w9410 = w6264 & w8923;
assign w9411 = ~w9195 & w40708;
assign w9412 = ~w9409 & ~w9411;
assign w9413 = ~w9405 & w9412;
assign w9414 = ~w6264 & w8923;
assign w9415 = (w9414 & w9195) | (w9414 & w40709) | (w9195 & w40709);
assign w9416 = ~w6264 & ~w8923;
assign w9417 = ~w9195 & w40710;
assign w9418 = ~w9415 & ~w9417;
assign w9419 = ~w9172 & w9174;
assign w9420 = (~w9178 & w9172) | (~w9178 & w40711) | (w9172 & w40711);
assign w9421 = ~w8897 & ~w8907;
assign w9422 = (w9421 & w9420) | (w9421 & w52069) | (w9420 & w52069);
assign w9423 = ~w9195 & w9422;
assign w9424 = ~w6769 & ~w8905;
assign w9425 = (w9424 & w9195) | (w9424 & w40712) | (w9195 & w40712);
assign w9426 = ~w6769 & w8905;
assign w9427 = ~w9195 & w40713;
assign w9428 = ~w9425 & ~w9427;
assign w9429 = w9418 & ~w9428;
assign w9430 = w9413 & ~w9429;
assign w9431 = ~w9397 & w9430;
assign w9432 = ~w9394 & w9431;
assign w9433 = w6769 & w8905;
assign w9434 = (w9433 & w9195) | (w9433 & w40714) | (w9195 & w40714);
assign w9435 = w6769 & ~w8905;
assign w9436 = ~w9195 & w40715;
assign w9437 = ~w9434 & ~w9436;
assign w9438 = w9418 & w9437;
assign w9439 = w9413 & ~w9438;
assign w9440 = w8784 & ~w8785;
assign w9441 = ~w8784 & w8785;
assign w9442 = ~w9440 & ~w9441;
assign w9443 = w8790 & w8954;
assign w9444 = w9443 & w52228;
assign w9445 = (w8937 & w52071) | (w8937 & w52072) | (w52071 & w52072);
assign w9446 = ~w9444 & ~w9445;
assign w9447 = w9195 & w9442;
assign w9448 = ~w9195 & w9446;
assign w9449 = ~w9447 & ~w9448;
assign w9450 = w4838 & ~w9449;
assign w9451 = ~w8775 & ~w8776;
assign w9452 = w8954 & ~w8957;
assign w9453 = w8790 & w52229;
assign w9454 = w9451 & ~w9453;
assign w9455 = ~w9451 & w9453;
assign w9456 = ~w9454 & ~w9455;
assign w9457 = w8774 & w9195;
assign w9458 = ~w9195 & w9456;
assign w9459 = ~w9457 & ~w9458;
assign w9460 = ~w4430 & w9459;
assign w9461 = ~w9450 & ~w9460;
assign w9462 = w5745 & w9404;
assign w9463 = ~w8946 & ~w8957;
assign w9464 = (w9463 & w8937) | (w9463 & w52073) | (w8937 & w52073);
assign w9465 = ~w8937 & w52074;
assign w9466 = ~w9464 & ~w9465;
assign w9467 = ~w8945 & w9195;
assign w9468 = ~w9195 & ~w9466;
assign w9469 = ~w9467 & ~w9468;
assign w9470 = ~w5330 & ~w9469;
assign w9471 = ~w9462 & ~w9470;
assign w9472 = w9461 & w9471;
assign w9473 = ~w9439 & w9472;
assign w9474 = ~w9432 & w9473;
assign w9475 = w5330 & w9469;
assign w9476 = ~w4838 & w9449;
assign w9477 = ~w9450 & ~w9476;
assign w9478 = ~w9475 & w9477;
assign w9479 = w9461 & ~w9478;
assign w9480 = ~w8814 & w8860;
assign w9481 = w8955 & ~w8957;
assign w9482 = (w9481 & w8937) | (w9481 & w40717) | (w8937 & w40717);
assign w9483 = w8791 & ~w9482;
assign w9484 = (w8906 & w8924) | (w8906 & w40718) | (w8924 & w40718);
assign w9485 = ~w8946 & w8956;
assign w9486 = (w9485 & w9484) | (w9485 & w52075) | (w9484 & w52075);
assign w9487 = ~w9483 & w52076;
assign w9488 = (~w9480 & w9483) | (~w9480 & w52077) | (w9483 & w52077);
assign w9489 = ~w8813 & w9195;
assign w9490 = ~w9195 & w40719;
assign w9491 = ~w9489 & ~w9490;
assign w9492 = w4056 & ~w9491;
assign w9493 = w4430 & ~w9459;
assign w9494 = ~w9492 & ~w9493;
assign w9495 = (w9494 & w9478) | (w9494 & w40720) | (w9478 & w40720);
assign w9496 = w8879 & ~w8966;
assign w9497 = w8955 & w52078;
assign w9498 = ~w8864 & w9497;
assign w9499 = ~w8949 & w9498;
assign w9500 = (~w8867 & ~w8863) | (~w8867 & w47264) | (~w8863 & w47264);
assign w9501 = (w9496 & w9499) | (w9496 & w47265) | (w9499 & w47265);
assign w9502 = ~w9499 & w47266;
assign w9503 = ~w9501 & ~w9502;
assign w9504 = w8965 & w9195;
assign w9505 = ~w9195 & w9503;
assign w9506 = ~w9504 & ~w9505;
assign w9507 = ~w2558 & ~w9506;
assign w9508 = w8847 & ~w8867;
assign w9509 = (w8852 & ~w8861) | (w8852 & w52079) | (~w8861 & w52079);
assign w9510 = ~w8831 & w9509;
assign w9511 = w9481 & ~w9510;
assign w9512 = ~w8831 & w8852;
assign w9513 = ~w8791 & w8862;
assign w9514 = w9512 & ~w9513;
assign w9515 = ~w8949 & w9511;
assign w9516 = (w9508 & w9515) | (w9508 & w40721) | (w9515 & w40721);
assign w9517 = ~w9515 & w40722;
assign w9518 = ~w9516 & ~w9517;
assign w9519 = ~w9195 & ~w9518;
assign w9520 = ~w8832 & ~w8865;
assign w9521 = w9195 & w9520;
assign w9522 = ~w9519 & ~w9521;
assign w9523 = w2896 & w9522;
assign w9524 = ~w9507 & ~w9523;
assign w9525 = (w8860 & ~w8791) | (w8860 & w52080) | (~w8791 & w52080);
assign w9526 = w8860 & w9481;
assign w9527 = ~w8949 & w9526;
assign w9528 = ~w8805 & ~w8815;
assign w9529 = (w40723 & w8949) | (w40723 & w52081) | (w8949 & w52081);
assign w9530 = ~w8815 & ~w9529;
assign w9531 = ~w9195 & w9530;
assign w9532 = ~w3646 & w9192;
assign w9533 = (w9532 & w9172) | (w9532 & w52082) | (w9172 & w52082);
assign w9534 = ~w9135 & w9533;
assign w9535 = ~w9131 & w9534;
assign w9536 = w8828 & w8852;
assign w9537 = ~w3242 & ~w9536;
assign w9538 = (w9537 & w9531) | (w9537 & w40724) | (w9531 & w40724);
assign w9539 = ~w3242 & w9536;
assign w9540 = ~w9535 & w9539;
assign w9541 = ~w9531 & w9540;
assign w9542 = ~w9527 & w40725;
assign w9543 = (w9528 & w9527) | (w9528 & w40726) | (w9527 & w40726);
assign w9544 = ~w9542 & ~w9543;
assign w9545 = ~w9195 & ~w9544;
assign w9546 = w8804 & w9192;
assign w9547 = (w9546 & w9172) | (w9546 & w52085) | (w9172 & w52085);
assign w9548 = ~w9135 & w9547;
assign w9549 = ~w9131 & w9548;
assign w9550 = ~w3646 & ~w9549;
assign w9551 = ~w9545 & w9550;
assign w9552 = ~w9541 & ~w9551;
assign w9553 = ~w9538 & w9552;
assign w9554 = w9524 & w9553;
assign w9555 = ~w2896 & ~w9522;
assign w9556 = ~w9523 & ~w9555;
assign w9557 = w3242 & ~w9536;
assign w9558 = ~w9531 & w40727;
assign w9559 = w3242 & w9536;
assign w9560 = (w9559 & w9531) | (w9559 & w40728) | (w9531 & w40728);
assign w9561 = ~w9558 & ~w9560;
assign w9562 = w9556 & w9561;
assign w9563 = w9524 & ~w9562;
assign w9564 = ~w9554 & ~w9563;
assign w9565 = w9495 & ~w9564;
assign w9566 = ~w9474 & w9565;
assign w9567 = ~w4056 & w9491;
assign w9568 = ~w9545 & ~w9549;
assign w9569 = w3646 & ~w9568;
assign w9570 = ~w9567 & ~w9569;
assign w9571 = w9554 & ~w9570;
assign w9572 = ~w9563 & ~w9571;
assign w9573 = ~w8969 & w9195;
assign w9574 = w8745 & ~w8970;
assign w9575 = (w9574 & ~w8962) | (w9574 & w40729) | (~w8962 & w40729);
assign w9576 = ~w9195 & ~w9575;
assign w9577 = w8962 & w40730;
assign w9578 = w9576 & ~w9577;
assign w9579 = ~w9573 & ~w9578;
assign w9580 = ~w9578 & w40731;
assign w9581 = w2558 & w9506;
assign w9582 = ~w9580 & ~w9581;
assign w9583 = w9572 & w9582;
assign w9584 = w8973 & w40732;
assign w9585 = w8962 & w9584;
assign w9586 = ~w9134 & ~w9145;
assign w9587 = ~w9144 & ~w9145;
assign w9588 = w9150 & ~w9587;
assign w9589 = (w9588 & w9134) | (w9588 & w40733) | (w9134 & w40733);
assign w9590 = (w9042 & w9585) | (w9042 & w40734) | (w9585 & w40734);
assign w9591 = w9074 & ~w9154;
assign w9592 = ~w9153 & w9195;
assign w9593 = ~w9195 & ~w9591;
assign w9594 = w9590 & w9593;
assign w9595 = ~w9195 & w9591;
assign w9596 = ~w9590 & w9595;
assign w9597 = ~w9594 & ~w9596;
assign w9598 = (w57 & ~w9597) | (w57 & w40735) | (~w9597 & w40735);
assign w9599 = w9042 & w9150;
assign w9600 = (~w9587 & w9134) | (~w9587 & w40736) | (w9134 & w40736);
assign w9601 = ~w9585 & w9600;
assign w9602 = w351 & w9195;
assign w9603 = ~w9195 & w9601;
assign w9604 = ~w9602 & ~w9603;
assign w9605 = w9599 & w9604;
assign w9606 = ~w9599 & ~w9604;
assign w9607 = ~w9605 & ~w9606;
assign w9608 = w252 & w9607;
assign w9609 = ~w9598 & ~w9608;
assign w9610 = ~w9131 & ~w9135;
assign w9611 = w9074 & ~w9193;
assign w9612 = w9610 & ~w9611;
assign w9613 = ~w9154 & w9588;
assign w9614 = ~w9586 & w9613;
assign w9615 = ~w9585 & w9614;
assign w9616 = ~w9042 & ~w9154;
assign w9617 = ~w9615 & ~w9616;
assign w9618 = ~w9612 & w9617;
assign w9619 = w57 & w9195;
assign w9620 = w9061 & w9164;
assign w9621 = ~w9618 & w40737;
assign w9622 = (w9620 & w9618) | (w9620 & w40738) | (w9618 & w40738);
assign w9623 = ~w9621 & ~w9622;
assign w9624 = ~w80 & w9623;
assign w9625 = w9609 & ~w9624;
assign w9626 = ~w9118 & ~w9195;
assign w9627 = w3 & w9192;
assign w9628 = (w9627 & w9172) | (w9627 & w52086) | (w9172 & w52086);
assign w9629 = ~w9135 & w9628;
assign w9630 = ~w9131 & w9629;
assign w9631 = w9075 & ~w9616;
assign w9632 = ~w9615 & w9631;
assign w9633 = ~w9626 & ~w9630;
assign w9634 = w9167 & ~w9630;
assign w9635 = ~w9632 & w9634;
assign w9636 = ~w9633 & ~w9635;
assign w9637 = w9125 & ~w9178;
assign w9638 = w42 & ~w9637;
assign w9639 = w9636 & w9638;
assign w9640 = w42 & w9637;
assign w9641 = ~w9636 & w9640;
assign w9642 = ~w9639 & ~w9641;
assign w9643 = w80 & w9195;
assign w9644 = w9164 & ~w9195;
assign w9645 = ~w9632 & w9644;
assign w9646 = ~w9643 & ~w9645;
assign w9647 = ~w9118 & ~w9166;
assign w9648 = w3 & w9647;
assign w9649 = (w9648 & w9645) | (w9648 & w40739) | (w9645 & w40739);
assign w9650 = w3 & ~w9647;
assign w9651 = (w9650 & ~w9195) | (w9650 & w40740) | (~w9195 & w40740);
assign w9652 = ~w9645 & w9651;
assign w9653 = ~w8677 & w47267;
assign w9654 = ~w9212 & w9653;
assign w9655 = ~w9419 & w9654;
assign w9656 = ~w9211 & w9655;
assign w9657 = ~w9128 & w9420;
assign w9658 = ~w9022 & w9180;
assign w9659 = ~w9657 & ~w9658;
assign w9660 = ~w42 & w9022;
assign w9661 = w9657 & ~w9660;
assign w9662 = w9655 & ~w9660;
assign w9663 = ~w9211 & w9662;
assign w9664 = ~w9661 & ~w9663;
assign w9665 = ~w9656 & w9659;
assign w9666 = w9664 & ~w9665;
assign w9667 = ~w9022 & w9188;
assign w9668 = w9657 & ~w9667;
assign w9669 = w9655 & ~w9667;
assign w9670 = ~w9211 & w9669;
assign w9671 = ~w9668 & ~w9670;
assign w9672 = ~w9179 & ~w9657;
assign w9673 = ~w9656 & w9672;
assign w9674 = w9671 & ~w9673;
assign w9675 = ~w9666 & ~w9674;
assign w9676 = ~w9652 & w9675;
assign w9677 = ~w9649 & w9676;
assign w9678 = w9642 & w9677;
assign w9679 = w9138 & ~w9142;
assign w9680 = (~w9104 & ~w9134) | (~w9104 & w40741) | (~w9134 & w40741);
assign w9681 = w8973 & w44428;
assign w9682 = w8962 & w9681;
assign w9683 = ~w9680 & ~w9682;
assign w9684 = ~w400 & w9195;
assign w9685 = ~w9195 & w9683;
assign w9686 = ~w9684 & ~w9685;
assign w9687 = ~w9088 & ~w9139;
assign w9688 = ~w351 & ~w9687;
assign w9689 = w9686 & w9688;
assign w9690 = ~w351 & w9687;
assign w9691 = ~w9686 & w9690;
assign w9692 = ~w9689 & ~w9691;
assign w9693 = ~w9104 & ~w9142;
assign w9694 = w9134 & w9138;
assign w9695 = w8962 & w9006;
assign w9696 = (w9693 & w9695) | (w9693 & w40742) | (w9695 & w40742);
assign w9697 = ~w9195 & ~w9696;
assign w9698 = ~w9695 & w40743;
assign w9699 = ~w9141 & w9195;
assign w9700 = w400 & w9699;
assign w9701 = w400 & ~w9698;
assign w9702 = w9697 & w9701;
assign w9703 = ~w9700 & ~w9702;
assign w9704 = w9692 & w9703;
assign w9705 = w9206 & w52087;
assign w9706 = ~w8611 & ~w9198;
assign w9707 = w8765 & ~w9706;
assign w9708 = ~w9001 & ~w9137;
assign w9709 = ~w9002 & ~w9708;
assign w9710 = w9002 & w9708;
assign w9711 = ~w9709 & ~w9710;
assign w9712 = (w9711 & w8975) | (w9711 & w40744) | (w8975 & w40744);
assign w9713 = w9707 & ~w9708;
assign w9714 = ~w8975 & w9713;
assign w9715 = ~w9136 & w9195;
assign w9716 = ~w9195 & ~w9714;
assign w9717 = ~w9712 & w9716;
assign w9718 = ~w9715 & ~w9717;
assign w9719 = (~w493 & w9717) | (~w493 & w40745) | (w9717 & w40745);
assign w9720 = ~w9705 & ~w9719;
assign w9721 = w9704 & w9720;
assign w9722 = w9678 & w9721;
assign w9723 = w9625 & w9722;
assign w9724 = w9583 & w9723;
assign w9725 = ~w9566 & w9724;
assign w9726 = ~w9209 & w9349;
assign w9727 = w9725 & ~w9726;
assign w9728 = w9636 & ~w9637;
assign w9729 = ~w9636 & w9637;
assign w9730 = ~w9728 & ~w9729;
assign w9731 = ~w42 & ~w9666;
assign w9732 = w9730 & w9731;
assign w9733 = ~w9678 & ~w9732;
assign w9734 = ~w252 & ~w9607;
assign w9735 = (w351 & ~w9686) | (w351 & w40746) | (~w9686 & w40746);
assign w9736 = ~w9686 & w9687;
assign w9737 = w9735 & ~w9736;
assign w9738 = ~w9734 & ~w9737;
assign w9739 = ~w400 & ~w9699;
assign w9740 = w9697 & ~w9698;
assign w9741 = w9739 & ~w9740;
assign w9742 = ~w9717 & w40747;
assign w9743 = ~w9741 & ~w9742;
assign w9744 = w9704 & ~w9743;
assign w9745 = w9738 & ~w9744;
assign w9746 = w9597 & w40748;
assign w9747 = w80 & w9620;
assign w9748 = (w9747 & w9618) | (w9747 & w40749) | (w9618 & w40749);
assign w9749 = w80 & ~w9620;
assign w9750 = ~w9618 & w40750;
assign w9751 = ~w9748 & ~w9750;
assign w9752 = ~w9746 & w9751;
assign w9753 = ~w9624 & ~w9752;
assign w9754 = ~w9645 & w40751;
assign w9755 = ~w3 & ~w9754;
assign w9756 = ~w9646 & w9647;
assign w9757 = w9755 & ~w9756;
assign w9758 = ~w9732 & ~w9757;
assign w9759 = ~w9753 & w9758;
assign w9760 = w9625 & ~w9745;
assign w9761 = w9759 & ~w9760;
assign w9762 = w9195 & w40752;
assign w9763 = w2285 & ~w9577;
assign w9764 = w9576 & w9763;
assign w9765 = ~w9762 & ~w9764;
assign w9766 = (w2006 & ~w9195) | (w2006 & w40753) | (~w9195 & w40753);
assign w9767 = ~w9341 & w9766;
assign w9768 = w9765 & ~w9767;
assign w9769 = w9335 & w9768;
assign w9770 = w9242 & ~w9769;
assign w9771 = w9346 & w9770;
assign w9772 = ~w9321 & w9771;
assign w9773 = ~w9242 & w40754;
assign w9774 = ~w9209 & w9312;
assign w9775 = w9306 & w9774;
assign w9776 = ~w9773 & ~w9775;
assign w9777 = ~w9772 & ~w9776;
assign w9778 = ~w9733 & ~w9761;
assign w9779 = w9723 & ~w9777;
assign w9780 = ~w9778 & ~w9779;
assign w9781 = ~w9727 & w9780;
assign w9782 = w9346 & w9582;
assign w9783 = w9572 & w9782;
assign w9784 = w9769 & w9783;
assign w9785 = ~w9566 & w9784;
assign w9786 = w9346 & ~w9769;
assign w9787 = ~w9268 & ~w9317;
assign w9788 = w9786 & ~w9787;
assign w9789 = ~w9786 & w9787;
assign w9790 = ~w9788 & ~w9789;
assign w9791 = w9785 & ~w9790;
assign w9792 = ~w9785 & w9790;
assign w9793 = ~w9791 & ~w9792;
assign w9794 = w9267 & ~w9781;
assign w9795 = w9781 & ~w9793;
assign w9796 = ~w9794 & ~w9795;
assign w9797 = w1320 & w9796;
assign w9798 = ~w9344 & w9768;
assign w9799 = w9572 & w40755;
assign w9800 = ~w9566 & w9799;
assign w9801 = ~w9344 & ~w9768;
assign w9802 = ~w9330 & w9335;
assign w9803 = w9801 & ~w9802;
assign w9804 = ~w9801 & w9802;
assign w9805 = ~w9803 & ~w9804;
assign w9806 = ~w9566 & w40756;
assign w9807 = (w9805 & w9566) | (w9805 & w40757) | (w9566 & w40757);
assign w9808 = ~w9806 & ~w9807;
assign w9809 = w9329 & ~w9781;
assign w9810 = w9781 & w9808;
assign w9811 = ~w9809 & ~w9810;
assign w9812 = w1541 & ~w9811;
assign w9813 = ~w9797 & ~w9812;
assign w9814 = w9572 & ~w9581;
assign w9815 = ~w9580 & w9765;
assign w9816 = (~w9815 & w9566) | (~w9815 & w40758) | (w9566 & w40758);
assign w9817 = w9572 & w44429;
assign w9818 = ~w9566 & w9817;
assign w9819 = ~w9579 & ~w9781;
assign w9820 = ~w9816 & ~w9818;
assign w9821 = w9781 & w9820;
assign w9822 = ~w9819 & ~w9821;
assign w9823 = w2006 & ~w9822;
assign w9824 = w2006 & ~w9765;
assign w9825 = ~w2006 & w9765;
assign w9826 = ~w9824 & ~w9825;
assign w9827 = ~w9566 & w44430;
assign w9828 = (~w9826 & w9566) | (~w9826 & w44431) | (w9566 & w44431);
assign w9829 = ~w9827 & ~w9828;
assign w9830 = w9781 & w9829;
assign w9831 = w1738 & w9343;
assign w9832 = (w9831 & ~w9781) | (w9831 & w44432) | (~w9781 & w44432);
assign w9833 = w1738 & ~w9343;
assign w9834 = w9781 & w44433;
assign w9835 = ~w9832 & ~w9834;
assign w9836 = ~w9823 & w9835;
assign w9837 = w9813 & w9836;
assign w9838 = ~w9495 & w9570;
assign w9839 = w9473 & w9570;
assign w9840 = ~w9432 & w9839;
assign w9841 = ~w9840 & w40759;
assign w9842 = w9562 & ~w9841;
assign w9843 = ~w9556 & ~w9561;
assign w9844 = w9553 & ~w9556;
assign w9845 = ~w9840 & w40760;
assign w9846 = ~w9843 & ~w9845;
assign w9847 = w9522 & ~w9781;
assign w9848 = ~w9842 & w9846;
assign w9849 = w9781 & w9848;
assign w9850 = ~w9847 & ~w9849;
assign w9851 = ~w2558 & ~w9850;
assign w9852 = w2558 & ~w9781;
assign w9853 = ~w9523 & ~w9842;
assign w9854 = w9781 & w9853;
assign w9855 = ~w9852 & ~w9854;
assign w9856 = ~w9507 & ~w9581;
assign w9857 = w2285 & ~w9856;
assign w9858 = w9855 & w9857;
assign w9859 = w2285 & w9856;
assign w9860 = ~w9855 & w9859;
assign w9861 = ~w9858 & ~w9860;
assign w9862 = ~w9851 & w9861;
assign w9863 = w9837 & w9862;
assign w9864 = ~a[60] & ~a[61];
assign w9865 = ~a[62] & w9864;
assign w9866 = ~w9195 & w9865;
assign w9867 = w9195 & ~w9865;
assign w9868 = ~w9866 & ~w9867;
assign w9869 = a[63] & ~w9868;
assign w9870 = ~w9350 & ~w9869;
assign w9871 = ~a[63] & w9868;
assign w9872 = ~w9866 & ~w9871;
assign w9873 = ~w9781 & w9872;
assign w9874 = ~w9866 & ~w9870;
assign w9875 = w9781 & w9874;
assign w9876 = ~w9873 & ~w9875;
assign w9877 = a[64] & ~w9350;
assign w9878 = ~w9351 & ~w9877;
assign w9879 = ~a[64] & ~w9195;
assign w9880 = a[64] & w9195;
assign w9881 = ~w9879 & ~w9880;
assign w9882 = w8666 & w9878;
assign w9883 = w9781 & w9882;
assign w9884 = w8666 & w9881;
assign w9885 = ~w9781 & w9884;
assign w9886 = ~w9883 & ~w9885;
assign w9887 = ~w9876 & w9886;
assign w9888 = ~w8666 & ~w9881;
assign w9889 = ~w9781 & w9888;
assign w9890 = ~w8666 & ~w9878;
assign w9891 = w9781 & w9890;
assign w9892 = ~w9889 & ~w9891;
assign w9893 = w7924 & w9892;
assign w9894 = ~w9887 & w9893;
assign w9895 = ~w9365 & ~w9374;
assign w9896 = (w9373 & ~w9781) | (w9373 & w40761) | (~w9781 & w40761);
assign w9897 = w9781 & w40762;
assign w9898 = ~w9896 & ~w9897;
assign w9899 = w7315 & w9898;
assign w9900 = ~w9894 & ~w9899;
assign w9901 = ~w9377 & ~w9397;
assign w9902 = w9781 & w9901;
assign w9903 = w6769 & w9393;
assign w9904 = (w9903 & ~w9781) | (w9903 & w40763) | (~w9781 & w40763);
assign w9905 = w6769 & ~w9393;
assign w9906 = w9781 & w40764;
assign w9907 = ~w9904 & ~w9906;
assign w9908 = ~w7315 & w9373;
assign w9909 = (w9908 & ~w9781) | (w9908 & w40765) | (~w9781 & w40765);
assign w9910 = ~w7315 & ~w9373;
assign w9911 = w9781 & w40766;
assign w9912 = ~w9909 & ~w9911;
assign w9913 = w9907 & w9912;
assign w9914 = ~w7924 & ~w9892;
assign w9915 = a[65] & ~w9879;
assign w9916 = ~w9195 & w9781;
assign w9917 = (w9915 & ~w9781) | (w9915 & w40767) | (~w9781 & w40767);
assign w9918 = ~w9352 & w9781;
assign w9919 = w8883 & ~w9195;
assign w9920 = ~w9354 & ~w9355;
assign w9921 = ~w9195 & w9920;
assign w9922 = w9195 & ~w9920;
assign w9923 = ~w9921 & ~w9922;
assign w9924 = (~w9919 & ~w9781) | (~w9919 & w40768) | (~w9781 & w40768);
assign w9925 = ~w9917 & w9924;
assign w9926 = w9918 & w9923;
assign w9927 = ~w9925 & ~w9926;
assign w9928 = ~w9914 & ~w9927;
assign w9929 = ~w7924 & w9887;
assign w9930 = (w9913 & w9894) | (w9913 & w40769) | (w9894 & w40769);
assign w9931 = w9913 & ~w9929;
assign w9932 = w9928 & w9931;
assign w9933 = ~w9930 & ~w9932;
assign w9934 = (w9428 & w9396) | (w9428 & w40770) | (w9396 & w40770);
assign w9935 = (w9437 & w9394) | (w9437 & w40771) | (w9394 & w40771);
assign w9936 = ~w9405 & ~w9462;
assign w9937 = w9418 & ~w9936;
assign w9938 = w9412 & ~w9935;
assign w9939 = w9937 & ~w9938;
assign w9940 = ~w9439 & ~w9462;
assign w9941 = ~w9432 & w9940;
assign w9942 = ~w9462 & ~w9941;
assign w9943 = ~w9939 & ~w9942;
assign w9944 = w5330 & ~w9404;
assign w9945 = ~w9781 & w9944;
assign w9946 = w5330 & ~w9943;
assign w9947 = w9781 & w9946;
assign w9948 = ~w9945 & ~w9947;
assign w9949 = w6264 & w9948;
assign w9950 = ~w5330 & w9404;
assign w9951 = ~w9781 & w9950;
assign w9952 = ~w5330 & w9943;
assign w9953 = w9781 & w9952;
assign w9954 = ~w9951 & ~w9953;
assign w9955 = ~w9394 & ~w9397;
assign w9956 = ~w6769 & ~w9955;
assign w9957 = w9781 & ~w9956;
assign w9958 = w8905 & ~w9423;
assign w9959 = ~w8905 & w9423;
assign w9960 = ~w9958 & ~w9959;
assign w9961 = w8923 & ~w9407;
assign w9962 = ~w8923 & w9407;
assign w9963 = ~w9961 & ~w9962;
assign w9964 = (~w9963 & ~w9781) | (~w9963 & w40772) | (~w9781 & w40772);
assign w9965 = ~w5745 & w9960;
assign w9966 = (w9965 & ~w9781) | (w9965 & w40773) | (~w9781 & w40773);
assign w9967 = w9964 & ~w9966;
assign w9968 = w6769 & w9955;
assign w9969 = ~w9960 & w9963;
assign w9970 = w9968 & w9969;
assign w9971 = w9781 & w9970;
assign w9972 = ~w9949 & w9954;
assign w9973 = w9954 & ~w9971;
assign w9974 = ~w9967 & w9973;
assign w9975 = ~w9972 & ~w9974;
assign w9976 = ~w9956 & ~w9968;
assign w9977 = w6264 & w9960;
assign w9978 = (w9977 & ~w9781) | (w9977 & w40774) | (~w9781 & w40774);
assign w9979 = w6264 & ~w9960;
assign w9980 = w9781 & w40775;
assign w9981 = ~w9978 & ~w9980;
assign w9982 = w9957 & w9963;
assign w9983 = ~w9981 & ~w9982;
assign w9984 = w9412 & w9418;
assign w9985 = w9935 & ~w9984;
assign w9986 = ~w9935 & w9984;
assign w9987 = ~w9985 & ~w9986;
assign w9988 = ~w9781 & ~w9963;
assign w9989 = w9781 & w9987;
assign w9990 = ~w9988 & ~w9989;
assign w9991 = ~w5745 & w9990;
assign w9992 = ~w5745 & w6264;
assign w9993 = w9948 & ~w9992;
assign w9994 = ~w9991 & w9993;
assign w9995 = ~w9983 & w9994;
assign w9996 = ~w9975 & ~w9995;
assign w9997 = ~w9393 & ~w9902;
assign w9998 = w9393 & w9902;
assign w9999 = ~w9997 & ~w9998;
assign w10000 = ~w6769 & ~w9999;
assign w10001 = ~w9470 & ~w9475;
assign w10002 = w9745 & ~w9753;
assign w10003 = w9723 & ~w10002;
assign w10004 = w5330 & ~w9781;
assign w10005 = w9781 & w9941;
assign w10006 = ~w10004 & ~w10005;
assign w10007 = ~w5330 & w10003;
assign w10008 = ~w10006 & ~w10007;
assign w10009 = (~w4838 & w10006) | (~w4838 & w40776) | (w10006 & w40776);
assign w10010 = (~w10001 & w10006) | (~w10001 & w44434) | (w10006 & w44434);
assign w10011 = w10009 & ~w10010;
assign w10012 = ~w10000 & ~w10011;
assign w10013 = ~w9996 & w10012;
assign w10014 = w9933 & w10013;
assign w10015 = ~w6264 & ~w9960;
assign w10016 = (w10015 & ~w9781) | (w10015 & w40777) | (~w9781 & w40777);
assign w10017 = ~w6264 & w9960;
assign w10018 = w9781 & w40778;
assign w10019 = ~w10016 & ~w10018;
assign w10020 = w5745 & ~w9990;
assign w10021 = w9954 & ~w10020;
assign w10022 = ~w9991 & ~w10019;
assign w10023 = w10021 & ~w10022;
assign w10024 = ~w10011 & ~w10023;
assign w10025 = ~w9996 & w10024;
assign w10026 = (w9495 & w9432) | (w9495 & w40779) | (w9432 & w40779);
assign w10027 = ~w9567 & ~w10026;
assign w10028 = w3646 & w10027;
assign w10029 = ~w3646 & ~w9492;
assign w10030 = ~w10027 & w10029;
assign w10031 = ~w10028 & ~w10030;
assign w10032 = w3242 & ~w9568;
assign w10033 = (w10032 & ~w9781) | (w10032 & w40780) | (~w9781 & w40780);
assign w10034 = w3242 & w9568;
assign w10035 = w9781 & w40781;
assign w10036 = ~w10033 & ~w10035;
assign w10037 = (~w9479 & w9432) | (~w9479 & w40782) | (w9432 & w40782);
assign w10038 = ~w9493 & w10037;
assign w10039 = ~w9432 & w40783;
assign w10040 = w9478 & ~w10039;
assign w10041 = ~w9450 & w10037;
assign w10042 = ~w10040 & w10041;
assign w10043 = ~w9460 & w10038;
assign w10044 = ~w10042 & ~w10043;
assign w10045 = w9781 & ~w10044;
assign w10046 = w4430 & ~w9450;
assign w10047 = ~w10040 & w10046;
assign w10048 = (~w9459 & ~w9781) | (~w9459 & w40784) | (~w9781 & w40784);
assign w10049 = ~w10045 & ~w10048;
assign w10050 = ~w4056 & w10049;
assign w10051 = ~w9492 & ~w9567;
assign w10052 = w10038 & ~w10051;
assign w10053 = ~w10038 & w10051;
assign w10054 = ~w10052 & ~w10053;
assign w10055 = w9491 & ~w9781;
assign w10056 = w9781 & ~w10054;
assign w10057 = ~w10055 & ~w10056;
assign w10058 = w3646 & ~w10057;
assign w10059 = w10036 & ~w10058;
assign w10060 = ~w10050 & w10059;
assign w10061 = (w4838 & ~w10006) | (w4838 & w40785) | (~w10006 & w40785);
assign w10062 = ~w10001 & w10008;
assign w10063 = w10061 & ~w10062;
assign w10064 = ~w9475 & ~w10039;
assign w10065 = ~w9477 & ~w10064;
assign w10066 = ~w9449 & ~w9781;
assign w10067 = ~w10040 & ~w10065;
assign w10068 = w9781 & w10067;
assign w10069 = ~w10066 & ~w10068;
assign w10070 = ~w4430 & ~w10069;
assign w10071 = (~w10070 & w10062) | (~w10070 & w40786) | (w10062 & w40786);
assign w10072 = w10060 & w10071;
assign w10073 = ~w10025 & w10072;
assign w10074 = ~w10014 & w10073;
assign w10075 = ~w9538 & ~w9541;
assign w10076 = ~w3242 & w10075;
assign w10077 = w9561 & ~w10076;
assign w10078 = w9561 & w10075;
assign w10079 = ~w9840 & w40787;
assign w10080 = w10078 & ~w10079;
assign w10081 = ~w10078 & w10079;
assign w10082 = ~w10080 & ~w10081;
assign w10083 = ~w9781 & w10077;
assign w10084 = w9781 & w10082;
assign w10085 = ~w10083 & ~w10084;
assign w10086 = w2896 & ~w10085;
assign w10087 = ~w3242 & w9568;
assign w10088 = (w10087 & ~w9781) | (w10087 & w40788) | (~w9781 & w40788);
assign w10089 = ~w3242 & ~w9568;
assign w10090 = w9781 & w40789;
assign w10091 = ~w10088 & ~w10090;
assign w10092 = ~w10086 & w10091;
assign w10093 = ~w3646 & w10057;
assign w10094 = w10036 & w10093;
assign w10095 = w4430 & w10069;
assign w10096 = w9781 & w40790;
assign w10097 = w4056 & ~w9459;
assign w10098 = (w10097 & ~w9781) | (w10097 & w40791) | (~w9781 & w40791);
assign w10099 = ~w10096 & ~w10098;
assign w10100 = ~w10095 & w10099;
assign w10101 = (~w10094 & ~w10060) | (~w10094 & w40792) | (~w10060 & w40792);
assign w10102 = w10092 & w10101;
assign w10103 = w9863 & w10102;
assign w10104 = ~w10074 & w10103;
assign w10105 = ~w9566 & w9583;
assign w10106 = (w9769 & w9313) | (w9769 & w40793) | (w9313 & w40793);
assign w10107 = ~w9209 & w9743;
assign w10108 = w10106 & w10107;
assign w10109 = ~w10105 & w10108;
assign w10110 = ~w9720 & w9743;
assign w10111 = w9704 & ~w10110;
assign w10112 = w9609 & w10111;
assign w10113 = w10111 & w50185;
assign w10114 = w9609 & ~w9738;
assign w10115 = (~w10114 & w10109) | (~w10114 & w40795) | (w10109 & w40795);
assign w10116 = ~w9746 & w9781;
assign w10117 = w10115 & w10116;
assign w10118 = ~w9624 & w9751;
assign w10119 = ~w3 & ~w10118;
assign w10120 = (w10119 & w9781) | (w10119 & w40796) | (w9781 & w40796);
assign w10121 = ~w10117 & w10120;
assign w10122 = ~w3 & w10118;
assign w10123 = ~w9781 & w40797;
assign w10124 = ~w9746 & w10122;
assign w10125 = w9781 & w10124;
assign w10126 = w10115 & w10125;
assign w10127 = ~w10123 & ~w10126;
assign w10128 = ~w10121 & w10127;
assign w10129 = w9752 & ~w10114;
assign w10130 = (w10129 & w10109) | (w10129 & w40798) | (w10109 & w40798);
assign w10131 = ~w9624 & w9781;
assign w10132 = ~w10130 & w10131;
assign w10133 = ~w3 & ~w9781;
assign w10134 = ~w9649 & ~w9652;
assign w10135 = ~w9757 & w10134;
assign w10136 = ~w42 & w10135;
assign w10137 = (w10136 & w9781) | (w10136 & w40799) | (w9781 & w40799);
assign w10138 = ~w10132 & w10137;
assign w10139 = ~w42 & ~w10135;
assign w10140 = ~w9781 & w40800;
assign w10141 = ~w9624 & w10139;
assign w10142 = w9781 & w10141;
assign w10143 = ~w10130 & w10142;
assign w10144 = ~w10140 & ~w10143;
assign w10145 = ~w10138 & w10144;
assign w10146 = w10128 & w10145;
assign w10147 = (w10111 & ~w9349) | (w10111 & w40801) | (~w9349 & w40801);
assign w10148 = ~w10109 & w10147;
assign w10149 = (w9738 & w10109) | (w9738 & w40802) | (w10109 & w40802);
assign w10150 = ~w9608 & w9781;
assign w10151 = ~w10149 & w10150;
assign w10152 = ~w9598 & ~w9746;
assign w10153 = w80 & w10152;
assign w10154 = (w10153 & w9781) | (w10153 & w40803) | (w9781 & w40803);
assign w10155 = ~w10151 & w10154;
assign w10156 = w80 & ~w10152;
assign w10157 = ~w9781 & w40804;
assign w10158 = ~w9608 & w10156;
assign w10159 = w9781 & w10158;
assign w10160 = ~w10149 & w10159;
assign w10161 = ~w10157 & ~w10160;
assign w10162 = ~w10155 & w10161;
assign w10163 = ~w9737 & w9781;
assign w10164 = ~w10148 & w10163;
assign w10165 = ~w9608 & ~w9734;
assign w10166 = w57 & w10165;
assign w10167 = (w10166 & w9781) | (w10166 & w40805) | (w9781 & w40805);
assign w10168 = ~w10164 & w10167;
assign w10169 = w57 & ~w10165;
assign w10170 = (w10169 & w10109) | (w10169 & w40806) | (w10109 & w40806);
assign w10171 = w10163 & w10170;
assign w10172 = ~w9781 & w40807;
assign w10173 = ~w10171 & ~w10172;
assign w10174 = ~w10168 & w10173;
assign w10175 = w10162 & ~w10174;
assign w10176 = ~w80 & ~w10152;
assign w10177 = (w10176 & w9781) | (w10176 & w40808) | (w9781 & w40808);
assign w10178 = ~w10151 & w10177;
assign w10179 = ~w80 & w10152;
assign w10180 = ~w9781 & w40809;
assign w10181 = ~w9608 & w10179;
assign w10182 = w9781 & w10181;
assign w10183 = ~w10149 & w10182;
assign w10184 = ~w10180 & ~w10183;
assign w10185 = ~w10178 & w10184;
assign w10186 = w3 & w10118;
assign w10187 = (w10186 & w9781) | (w10186 & w40810) | (w9781 & w40810);
assign w10188 = ~w10117 & w10187;
assign w10189 = w3 & ~w10118;
assign w10190 = ~w9781 & w40811;
assign w10191 = ~w9746 & w10189;
assign w10192 = w9781 & w10191;
assign w10193 = w10115 & w10192;
assign w10194 = ~w10190 & ~w10193;
assign w10195 = ~w10188 & w10194;
assign w10196 = w10185 & w10195;
assign w10197 = ~w10175 & w10196;
assign w10198 = w9666 & w9730;
assign w10199 = w9642 & ~w10198;
assign w10200 = ~w9624 & ~w10130;
assign w10201 = ~w10134 & ~w10199;
assign w10202 = ~w9757 & ~w10199;
assign w10203 = ~w10200 & w10202;
assign w10204 = ~w10201 & ~w10203;
assign w10205 = ~w9757 & ~w10200;
assign w10206 = ~w9674 & w9730;
assign w10207 = w9642 & w10134;
assign w10208 = ~w10206 & w10207;
assign w10209 = ~w10205 & w10208;
assign w10210 = ~w10132 & ~w10133;
assign w10211 = w42 & w10135;
assign w10212 = (w10211 & w10132) | (w10211 & w40812) | (w10132 & w40812);
assign w10213 = w42 & ~w10135;
assign w10214 = ~w10132 & w40813;
assign w10215 = ~w10212 & ~w10214;
assign w10216 = w10204 & ~w10209;
assign w10217 = w10215 & w10216;
assign w10218 = (w10217 & w10197) | (w10217 & w40814) | (w10197 & w40814);
assign w10219 = w9703 & ~w10110;
assign w10220 = (w10219 & ~w9349) | (w10219 & w40815) | (~w9349 & w40815);
assign w10221 = ~w10109 & w10220;
assign w10222 = w351 & ~w9781;
assign w10223 = w9781 & w10221;
assign w10224 = ~w10222 & ~w10223;
assign w10225 = w9692 & ~w9737;
assign w10226 = w252 & ~w10225;
assign w10227 = w10224 & w10226;
assign w10228 = w252 & w10225;
assign w10229 = ~w10224 & w10228;
assign w10230 = ~w10227 & ~w10229;
assign w10231 = w9348 & w9583;
assign w10232 = ~w9566 & w10231;
assign w10233 = ~w9720 & ~w9742;
assign w10234 = ~w9742 & w9777;
assign w10235 = ~w10232 & w10234;
assign w10236 = ~w10233 & ~w10235;
assign w10237 = w400 & ~w9781;
assign w10238 = w9781 & ~w10236;
assign w10239 = ~w10237 & ~w10238;
assign w10240 = w9703 & ~w9741;
assign w10241 = ~w351 & ~w10240;
assign w10242 = ~w10239 & w10241;
assign w10243 = ~w351 & w10240;
assign w10244 = w10239 & w10243;
assign w10245 = ~w10242 & ~w10244;
assign w10246 = w10230 & w10245;
assign w10247 = ~w9719 & ~w9742;
assign w10248 = w9705 & w10247;
assign w10249 = w9777 & w10247;
assign w10250 = ~w10232 & w10249;
assign w10251 = ~w10248 & ~w10250;
assign w10252 = w9781 & ~w10251;
assign w10253 = ~w9705 & ~w10247;
assign w10254 = (w10253 & w10232) | (w10253 & w40816) | (w10232 & w40816);
assign w10255 = w9718 & ~w9781;
assign w10256 = w9781 & w10254;
assign w10257 = ~w10255 & ~w10256;
assign w10258 = (~w400 & ~w10257) | (~w400 & w40817) | (~w10257 & w40817);
assign w10259 = w351 & w10240;
assign w10260 = ~w10239 & w10259;
assign w10261 = w351 & ~w10240;
assign w10262 = w10239 & w10261;
assign w10263 = ~w10260 & ~w10262;
assign w10264 = ~w10258 & w10263;
assign w10265 = ~w9209 & ~w9705;
assign w10266 = ~w9349 & ~w10265;
assign w10267 = (w10106 & w9566) | (w10106 & w40818) | (w9566 & w40818);
assign w10268 = w10266 & ~w10267;
assign w10269 = ~w10232 & w40819;
assign w10270 = ~w10268 & ~w10269;
assign w10271 = (w493 & w9781) | (w493 & w40820) | (w9781 & w40820);
assign w10272 = w9781 & w10270;
assign w10273 = w10271 & ~w10272;
assign w10274 = w9319 & ~w9769;
assign w10275 = w9346 & w10274;
assign w10276 = w9306 & ~w10275;
assign w10277 = ~w10275 & w40821;
assign w10278 = w9319 & w9582;
assign w10279 = w9346 & w10278;
assign w10280 = w9572 & w10279;
assign w10281 = w9241 & ~w10277;
assign w10282 = w9241 & w10280;
assign w10283 = ~w9566 & w10282;
assign w10284 = w9224 & w9247;
assign w10285 = ~w10283 & w40822;
assign w10286 = (w10284 & w10283) | (w10284 & w40823) | (w10283 & w40823);
assign w10287 = ~w10285 & ~w10286;
assign w10288 = w9218 & ~w9219;
assign w10289 = ~w9218 & w9219;
assign w10290 = ~w10288 & ~w10289;
assign w10291 = (w612 & w9781) | (w612 & w40824) | (w9781 & w40824);
assign w10292 = w9781 & ~w10287;
assign w10293 = w10291 & ~w10292;
assign w10294 = ~w10273 & ~w10293;
assign w10295 = (~w493 & w9781) | (~w493 & w40825) | (w9781 & w40825);
assign w10296 = w9781 & ~w10270;
assign w10297 = w10295 & ~w10296;
assign w10298 = w400 & ~w10252;
assign w10299 = w10257 & w10298;
assign w10300 = ~w10297 & ~w10299;
assign w10301 = ~w10294 & w10300;
assign w10302 = w10264 & ~w10301;
assign w10303 = w10246 & ~w10302;
assign w10304 = w10276 & w10280;
assign w10305 = ~w9566 & w10304;
assign w10306 = w9241 & w9311;
assign w10307 = ~w10275 & w40826;
assign w10308 = (w10306 & w10275) | (w10306 & w40827) | (w10275 & w40827);
assign w10309 = ~w10307 & ~w10308;
assign w10310 = w10305 & w10306;
assign w10311 = ~w10305 & ~w10309;
assign w10312 = ~w10310 & ~w10311;
assign w10313 = w9235 & ~w9236;
assign w10314 = ~w9235 & w9236;
assign w10315 = ~w10313 & ~w10314;
assign w10316 = w9781 & ~w10312;
assign w10317 = ~w9781 & ~w10315;
assign w10318 = ~w10316 & ~w10317;
assign w10319 = ~w754 & ~w10318;
assign w10320 = w9781 & w10287;
assign w10321 = ~w9781 & w10290;
assign w10322 = (~w612 & w9781) | (~w612 & w40828) | (w9781 & w40828);
assign w10323 = ~w10320 & w10322;
assign w10324 = ~w10319 & ~w10323;
assign w10325 = w10300 & w10324;
assign w10326 = w10246 & w10325;
assign w10327 = w1541 & w9195;
assign w10328 = w8758 & ~w9269;
assign w10329 = ~w9195 & w10328;
assign w10330 = ~w10327 & ~w10329;
assign w10331 = w9286 & w10330;
assign w10332 = ~w9286 & ~w10330;
assign w10333 = ~w10331 & ~w10332;
assign w10334 = ~w9295 & w9318;
assign w10335 = w9783 & ~w10334;
assign w10336 = ~w9295 & ~w9302;
assign w10337 = (~w9268 & ~w9346) | (~w9268 & w40829) | (~w9346 & w40829);
assign w10338 = ~w9317 & ~w10337;
assign w10339 = w10336 & ~w10338;
assign w10340 = ~w9566 & w10335;
assign w10341 = w10339 & ~w10340;
assign w10342 = ~w9317 & ~w10336;
assign w10343 = ~w10337 & w10342;
assign w10344 = w9783 & w10342;
assign w10345 = ~w9566 & w10344;
assign w10346 = ~w10343 & ~w10345;
assign w10347 = ~w9781 & w10333;
assign w10348 = ~w10341 & w10346;
assign w10349 = w9781 & w10348;
assign w10350 = ~w10347 & ~w10349;
assign w10351 = w1120 & ~w10350;
assign w10352 = (~w945 & w10350) | (~w945 & w40830) | (w10350 & w40830);
assign w10353 = ~w9284 & ~w9299;
assign w10354 = w1120 & ~w9298;
assign w10355 = (~w10354 & ~w9781) | (~w10354 & w40831) | (~w9781 & w40831);
assign w10356 = w9781 & w40832;
assign w10357 = ~w10355 & ~w10356;
assign w10358 = ~w9295 & ~w10353;
assign w10359 = w9781 & w40833;
assign w10360 = w9299 & ~w9781;
assign w10361 = ~w10359 & ~w10360;
assign w10362 = ~w10357 & w10361;
assign w10363 = ~w10350 & w40834;
assign w10364 = ~w10362 & ~w10363;
assign w10365 = w754 & w10318;
assign w10366 = ~w10352 & ~w10365;
assign w10367 = ~w10364 & w10366;
assign w10368 = w10326 & ~w10367;
assign w10369 = ~w10303 & ~w10368;
assign w10370 = ~w2006 & w9822;
assign w10371 = ~w2285 & ~w9856;
assign w10372 = ~w9855 & w10371;
assign w10373 = ~w2285 & w9856;
assign w10374 = w9855 & w10373;
assign w10375 = ~w10372 & ~w10374;
assign w10376 = ~w10370 & w10375;
assign w10377 = ~w1320 & ~w9796;
assign w10378 = ~w1541 & w9811;
assign w10379 = ~w1738 & ~w9343;
assign w10380 = (w10379 & ~w9781) | (w10379 & w44435) | (~w9781 & w44435);
assign w10381 = ~w1738 & w9343;
assign w10382 = w9781 & w44436;
assign w10383 = ~w10380 & ~w10382;
assign w10384 = ~w10378 & w10383;
assign w10385 = w9813 & ~w10384;
assign w10386 = ~w10377 & ~w10385;
assign w10387 = w9837 & ~w10376;
assign w10388 = w10386 & ~w10387;
assign w10389 = ~w2896 & w10085;
assign w10390 = w2558 & w9850;
assign w10391 = ~w10389 & ~w10390;
assign w10392 = w9863 & ~w10391;
assign w10393 = w10388 & ~w10392;
assign w10394 = ~w10369 & w10393;
assign w10395 = w10218 & w10394;
assign w10396 = ~w10104 & w10395;
assign w10397 = ~w1120 & w10350;
assign w10398 = w10350 & w40830;
assign w10399 = (w945 & ~w10350) | (w945 & w40834) | (~w10350 & w40834);
assign w10400 = ~w10362 & ~w10399;
assign w10401 = ~w10365 & ~w10398;
assign w10402 = ~w10400 & w10401;
assign w10403 = w10326 & ~w10402;
assign w10404 = ~w10303 & ~w10403;
assign w10405 = ~w57 & w10165;
assign w10406 = (w10405 & w10164) | (w10405 & w40835) | (w10164 & w40835);
assign w10407 = ~w57 & ~w10165;
assign w10408 = ~w10164 & w40836;
assign w10409 = ~w10406 & ~w10408;
assign w10410 = w10162 & w10409;
assign w10411 = ~w10224 & ~w10225;
assign w10412 = w10224 & w10225;
assign w10413 = ~w10411 & ~w10412;
assign w10414 = ~w252 & ~w10413;
assign w10415 = w10410 & ~w10414;
assign w10416 = w10146 & w10415;
assign w10417 = w10404 & w10416;
assign w10418 = (w10218 & ~w10404) | (w10218 & w40837) | (~w10404 & w40837);
assign w10419 = ~w10396 & ~w10418;
assign w10420 = ~w10025 & ~w10063;
assign w10421 = ~w10014 & w10420;
assign w10422 = w10092 & ~w10094;
assign w10423 = w10100 & w10422;
assign w10424 = (w10423 & ~w10388) | (w10423 & w40838) | (~w10388 & w40838);
assign w10425 = ~w10421 & w10424;
assign w10426 = w10391 & ~w10422;
assign w10427 = ~w10100 & w10391;
assign w10428 = w10060 & w10427;
assign w10429 = ~w10426 & ~w10428;
assign w10430 = ~w10070 & w10391;
assign w10431 = w10060 & w10430;
assign w10432 = w9863 & ~w10431;
assign w10433 = w10429 & w10432;
assign w10434 = w10388 & ~w10433;
assign w10435 = ~w10425 & w10434;
assign w10436 = w10404 & ~w10418;
assign w10437 = ~w10396 & w10436;
assign w10438 = ~w10425 & w40839;
assign w10439 = w10437 & ~w10438;
assign w10440 = ~w10104 & w10394;
assign w10441 = (w10417 & w10104) | (w10417 & w40840) | (w10104 & w40840);
assign w10442 = w252 & ~w10218;
assign w10443 = ~w10413 & ~w10442;
assign w10444 = ~w10441 & w10443;
assign w10445 = ~w10439 & ~w10444;
assign w10446 = w10324 & ~w10367;
assign w10447 = w10300 & w10446;
assign w10448 = w10302 & ~w10447;
assign w10449 = w10245 & ~w10448;
assign w10450 = (w10230 & w10218) | (w10230 & w44437) | (w10218 & w44437);
assign w10451 = (w10393 & w10074) | (w10393 & w40841) | (w10074 & w40841);
assign w10452 = w10324 & ~w10402;
assign w10453 = (w10294 & w10402) | (w10294 & w44438) | (w10402 & w44438);
assign w10454 = w10300 & ~w10453;
assign w10455 = w10264 & ~w10454;
assign w10456 = ~w10449 & ~w10450;
assign w10457 = ~w10450 & w10455;
assign w10458 = ~w10451 & w10457;
assign w10459 = ~w10456 & ~w10458;
assign w10460 = ~w57 & w10459;
assign w10461 = ~w10445 & w10460;
assign w10462 = (w10459 & w10439) | (w10459 & w40842) | (w10439 & w40842);
assign w10463 = w57 & ~w10462;
assign w10464 = ~w10461 & ~w10463;
assign w10465 = ~w10398 & ~w10418;
assign w10466 = ~w10396 & w10465;
assign w10467 = ~w10425 & w40843;
assign w10468 = w10466 & ~w10467;
assign w10469 = ~w10351 & ~w10362;
assign w10470 = ~w10433 & w40844;
assign w10471 = (~w10400 & w10425) | (~w10400 & w40845) | (w10425 & w40845);
assign w10472 = w10466 & w44439;
assign w10473 = (~w754 & w10396) | (~w754 & w40846) | (w10396 & w40846);
assign w10474 = ~w10319 & ~w10365;
assign w10475 = w612 & ~w10474;
assign w10476 = ~w10473 & w10475;
assign w10477 = ~w10472 & w10476;
assign w10478 = w612 & w10474;
assign w10479 = w10471 & w10478;
assign w10480 = w10468 & w10479;
assign w10481 = w10473 & w10478;
assign w10482 = ~w10480 & ~w10481;
assign w10483 = ~w10477 & w10482;
assign w10484 = w10393 & w10446;
assign w10485 = (~w10452 & w10104) | (~w10452 & w40847) | (w10104 & w40847);
assign w10486 = ~w612 & ~w10418;
assign w10487 = ~w10320 & ~w10321;
assign w10488 = (~w10487 & w10396) | (~w10487 & w40848) | (w10396 & w40848);
assign w10489 = w10419 & w10485;
assign w10490 = ~w10488 & ~w10489;
assign w10491 = ~w10319 & ~w10402;
assign w10492 = w10323 & ~w10491;
assign w10493 = w10293 & ~w10491;
assign w10494 = ~w10418 & w10493;
assign w10495 = ~w10319 & ~w10367;
assign w10496 = w10435 & w10495;
assign w10497 = (~w10492 & w10396) | (~w10492 & w40849) | (w10396 & w40849);
assign w10498 = ~w10496 & ~w10497;
assign w10499 = ~w10490 & w40850;
assign w10500 = w10483 & ~w10499;
assign w10501 = ~w612 & w10474;
assign w10502 = ~w10473 & w10501;
assign w10503 = ~w10472 & w10502;
assign w10504 = ~w612 & ~w10474;
assign w10505 = w10471 & w10504;
assign w10506 = w10468 & w10505;
assign w10507 = w10473 & w10504;
assign w10508 = ~w10506 & ~w10507;
assign w10509 = ~w10503 & w10508;
assign w10510 = (w10399 & w10425) | (w10399 & w44440) | (w10425 & w44440);
assign w10511 = w10466 & w47268;
assign w10512 = ~w754 & w10362;
assign w10513 = (w10512 & ~w10468) | (w10512 & w40852) | (~w10468 & w40852);
assign w10514 = ~w754 & ~w10362;
assign w10515 = w10468 & w40853;
assign w10516 = ~w10513 & ~w10515;
assign w10517 = w10509 & w10516;
assign w10518 = w10500 & ~w10517;
assign w10519 = ~w10433 & w40854;
assign w10520 = ~w10297 & ~w10418;
assign w10521 = ~w10396 & w10520;
assign w10522 = (w10453 & w10425) | (w10453 & w40855) | (w10425 & w40855);
assign w10523 = w10521 & ~w10522;
assign w10524 = (~w400 & w10396) | (~w400 & w40856) | (w10396 & w40856);
assign w10525 = ~w10258 & ~w10299;
assign w10526 = ~w351 & ~w10525;
assign w10527 = ~w10523 & w40857;
assign w10528 = ~w351 & w10525;
assign w10529 = (w10528 & w10523) | (w10528 & w40858) | (w10523 & w40858);
assign w10530 = ~w10527 & ~w10529;
assign w10531 = w10245 & w10263;
assign w10532 = w10393 & w10447;
assign w10533 = ~w10258 & ~w10454;
assign w10534 = (w10533 & w10104) | (w10533 & w40859) | (w10104 & w40859);
assign w10535 = w10531 & ~w10534;
assign w10536 = ~w10531 & w10534;
assign w10537 = ~w10535 & ~w10536;
assign w10538 = w10239 & ~w10240;
assign w10539 = ~w10239 & w10240;
assign w10540 = ~w10538 & ~w10539;
assign w10541 = ~w10419 & ~w10540;
assign w10542 = w252 & ~w10541;
assign w10543 = w10419 & w10537;
assign w10544 = w10542 & ~w10543;
assign w10545 = w10530 & ~w10544;
assign w10546 = (~w493 & w10490) | (~w493 & w40860) | (w10490 & w40860);
assign w10547 = ~w10293 & ~w10452;
assign w10548 = (w10547 & w10425) | (w10547 & w40861) | (w10425 & w40861);
assign w10549 = (w493 & w10396) | (w493 & w44441) | (w10396 & w44441);
assign w10550 = w10419 & ~w10548;
assign w10551 = ~w10273 & ~w10297;
assign w10552 = w400 & ~w10551;
assign w10553 = ~w10550 & w44442;
assign w10554 = w400 & w10551;
assign w10555 = (w10554 & w10550) | (w10554 & w44443) | (w10550 & w44443);
assign w10556 = ~w10553 & ~w10555;
assign w10557 = ~w10546 & w10556;
assign w10558 = w10545 & w10557;
assign w10559 = ~w10518 & w10558;
assign w10560 = w351 & ~w10525;
assign w10561 = (w10560 & w10523) | (w10560 & w40862) | (w10523 & w40862);
assign w10562 = w351 & w10525;
assign w10563 = ~w10523 & w40863;
assign w10564 = ~w10561 & ~w10563;
assign w10565 = ~w400 & ~w10551;
assign w10566 = (w10565 & w10550) | (w10565 & w44444) | (w10550 & w44444);
assign w10567 = ~w400 & w10551;
assign w10568 = ~w10550 & w44445;
assign w10569 = ~w10566 & ~w10568;
assign w10570 = w10564 & w10569;
assign w10571 = w10545 & ~w10570;
assign w10572 = (w57 & w10396) | (w57 & w40864) | (w10396 & w40864);
assign w10573 = (~w10414 & w10302) | (~w10414 & w40865) | (w10302 & w40865);
assign w10574 = w10326 & w40866;
assign w10575 = w10573 & ~w10574;
assign w10576 = ~w10418 & w10575;
assign w10577 = ~w10440 & w10576;
assign w10578 = w10174 & w10409;
assign w10579 = w80 & ~w10578;
assign w10580 = (w10579 & w10440) | (w10579 & w40867) | (w10440 & w40867);
assign w10581 = ~w10572 & w10580;
assign w10582 = w80 & w10578;
assign w10583 = w57 & w10582;
assign w10584 = (w10583 & w10396) | (w10583 & w40868) | (w10396 & w40868);
assign w10585 = ~w10440 & w40869;
assign w10586 = ~w10584 & ~w10585;
assign w10587 = ~w10581 & w10586;
assign w10588 = ~w10461 & w10587;
assign w10589 = ~w10419 & w10540;
assign w10590 = ~w252 & ~w10589;
assign w10591 = w10419 & ~w10537;
assign w10592 = w10590 & ~w10591;
assign w10593 = w10588 & ~w10592;
assign w10594 = ~w10175 & w10185;
assign w10595 = ~w10418 & w10594;
assign w10596 = ~w10396 & w10595;
assign w10597 = w10404 & w10415;
assign w10598 = (w10597 & w10104) | (w10597 & w40870) | (w10104 & w40870);
assign w10599 = w10596 & ~w10598;
assign w10600 = ~w10128 & ~w10418;
assign w10601 = (w10195 & w10396) | (w10195 & w40871) | (w10396 & w40871);
assign w10602 = w10128 & w10195;
assign w10603 = ~w3 & w10602;
assign w10604 = (w10603 & w10396) | (w10603 & w40872) | (w10396 & w40872);
assign w10605 = ~w10597 & w10602;
assign w10606 = w10394 & w10602;
assign w10607 = ~w10104 & w10606;
assign w10608 = ~w10605 & ~w10607;
assign w10609 = w10596 & ~w10608;
assign w10610 = ~w10604 & ~w10609;
assign w10611 = ~w10599 & ~w10601;
assign w10612 = w10610 & ~w10611;
assign w10613 = w10128 & w10410;
assign w10614 = w10575 & w10613;
assign w10615 = (w10614 & w10104) | (w10614 & w40873) | (w10104 & w40873);
assign w10616 = w10128 & ~w10197;
assign w10617 = ~w10615 & ~w10616;
assign w10618 = w10135 & ~w10210;
assign w10619 = ~w10135 & w10210;
assign w10620 = ~w10618 & ~w10619;
assign w10621 = ~w42 & ~w10620;
assign w10622 = ~w9730 & w10134;
assign w10623 = ~w10205 & w10622;
assign w10624 = w10204 & ~w10623;
assign w10625 = ~w42 & w10624;
assign w10626 = ~w10621 & ~w10625;
assign w10627 = ~w10617 & w10626;
assign w10628 = w10145 & w10617;
assign w10629 = ~w10627 & ~w10628;
assign w10630 = w10612 & w10629;
assign w10631 = w10174 & ~w10418;
assign w10632 = ~w10396 & w10631;
assign w10633 = w10409 & w10575;
assign w10634 = (w10633 & w10104) | (w10633 & w40874) | (w10104 & w40874);
assign w10635 = w10632 & ~w10634;
assign w10636 = (w80 & w10396) | (w80 & w40875) | (w10396 & w40875);
assign w10637 = ~w10635 & ~w10636;
assign w10638 = w10162 & w10185;
assign w10639 = ~w3 & ~w10638;
assign w10640 = (w10639 & w10635) | (w10639 & w40876) | (w10635 & w40876);
assign w10641 = ~w3 & w10638;
assign w10642 = ~w10635 & w40877;
assign w10643 = ~w10640 & ~w10642;
assign w10644 = ~w10630 & w10643;
assign w10645 = w10593 & w10644;
assign w10646 = ~w10571 & w10645;
assign w10647 = ~w10559 & w10646;
assign w10648 = ~w10572 & ~w10577;
assign w10649 = w10578 & ~w10648;
assign w10650 = (~w10578 & w10440) | (~w10578 & w40878) | (w10440 & w40878);
assign w10651 = ~w10572 & w10650;
assign w10652 = ~w80 & ~w10651;
assign w10653 = ~w10649 & w10652;
assign w10654 = w3 & ~w10638;
assign w10655 = ~w10635 & w40879;
assign w10656 = w3 & w10638;
assign w10657 = (w10656 & w10635) | (w10656 & w40880) | (w10635 & w40880);
assign w10658 = ~w10655 & ~w10657;
assign w10659 = ~w10653 & w10658;
assign w10660 = w10463 & w10587;
assign w10661 = w10659 & ~w10660;
assign w10662 = w10644 & ~w10661;
assign w10663 = w42 & w10620;
assign w10664 = (w10627 & ~w10612) | (w10627 & w44446) | (~w10612 & w44446);
assign w10665 = w9642 & ~w10209;
assign w10666 = ~w10623 & ~w10665;
assign w10667 = w10663 & w10666;
assign w10668 = ~w10621 & ~w10667;
assign w10669 = w10617 & ~w10668;
assign w10670 = (~w10669 & w10612) | (~w10669 & w44447) | (w10612 & w44447);
assign w10671 = ~w10664 & w10670;
assign w10672 = ~w10662 & w10671;
assign w10673 = ~w10647 & w10672;
assign w10674 = ~w10351 & ~w10397;
assign w10675 = w10419 & ~w10435;
assign w10676 = (w10674 & w10675) | (w10674 & w40882) | (w10675 & w40882);
assign w10677 = ~w10675 & w40883;
assign w10678 = ~w10676 & ~w10677;
assign w10679 = ~w945 & ~w10678;
assign w10680 = (w10468 & w44448) | (w10468 & w44449) | (w44448 & w44449);
assign w10681 = ~w10362 & w10511;
assign w10682 = w10680 & ~w10681;
assign w10683 = ~w10679 & ~w10682;
assign w10684 = w10500 & w10683;
assign w10685 = w10570 & w10684;
assign w10686 = w10645 & w10685;
assign w10687 = w9835 & w10383;
assign w10688 = ~w9851 & w10429;
assign w10689 = w10429 & w9862;
assign w10690 = w10429 & ~w10431;
assign w10691 = (w10376 & ~w10429) | (w10376 & w40885) | (~w10429 & w40885);
assign w10692 = w10421 & w10691;
assign w10693 = ~w10692 & w40886;
assign w10694 = (~w10687 & w10692) | (~w10687 & w44450) | (w10692 & w44450);
assign w10695 = w10419 & ~w10694;
assign w10696 = w10687 & w10693;
assign w10697 = w10695 & ~w10696;
assign w10698 = w9343 & ~w9830;
assign w10699 = ~w9343 & w9830;
assign w10700 = ~w10698 & ~w10699;
assign w10701 = (w10700 & w10396) | (w10700 & w44451) | (w10396 & w44451);
assign w10702 = (~w10701 & ~w10695) | (~w10701 & w44452) | (~w10695 & w44452);
assign w10703 = ~w1541 & ~w10702;
assign w10704 = ~w9812 & w10384;
assign w10705 = (w10704 & w10692) | (w10704 & w44453) | (w10692 & w44453);
assign w10706 = w10419 & ~w10705;
assign w10707 = ~w9812 & ~w10378;
assign w10708 = (w10383 & w10692) | (w10383 & w44454) | (w10692 & w44454);
assign w10709 = ~w10707 & ~w10708;
assign w10710 = w10706 & ~w10709;
assign w10711 = ~w1738 & ~w9781;
assign w10712 = ~w9800 & ~w9801;
assign w10713 = w9781 & w10712;
assign w10714 = ~w10711 & ~w10713;
assign w10715 = w9802 & w10714;
assign w10716 = ~w9802 & ~w10714;
assign w10717 = ~w10715 & ~w10716;
assign w10718 = (w10717 & w10396) | (w10717 & w44455) | (w10396 & w44455);
assign w10719 = ~w1320 & ~w10718;
assign w10720 = ~w10710 & w10719;
assign w10721 = (w9822 & w10396) | (w9822 & w44456) | (w10396 & w44456);
assign w10722 = ~w9823 & ~w10370;
assign w10723 = w10421 & ~w10690;
assign w10724 = w10429 & w52230;
assign w10725 = (w10722 & w10724) | (w10722 & w44457) | (w10724 & w44457);
assign w10726 = w10419 & ~w10725;
assign w10727 = ~w10724 & w44458;
assign w10728 = ~w1738 & w10721;
assign w10729 = ~w1738 & ~w10727;
assign w10730 = w10726 & w10729;
assign w10731 = ~w10728 & ~w10730;
assign w10732 = ~w10720 & w10731;
assign w10733 = ~w10703 & w10732;
assign w10734 = w9861 & w10375;
assign w10735 = (w10734 & ~w10429) | (w10734 & w40888) | (~w10429 & w40888);
assign w10736 = w10421 & w10735;
assign w10737 = w10688 & ~w10734;
assign w10738 = ~w10723 & w10737;
assign w10739 = ~w10688 & w10734;
assign w10740 = ~w10736 & ~w10739;
assign w10741 = ~w10738 & w10740;
assign w10742 = ~w9855 & ~w9856;
assign w10743 = w9855 & w9856;
assign w10744 = ~w10742 & ~w10743;
assign w10745 = w10419 & w10741;
assign w10746 = (w10744 & w10396) | (w10744 & w40889) | (w10396 & w40889);
assign w10747 = ~w10745 & ~w10746;
assign w10748 = ~w10745 & w40890;
assign w10749 = ~w10058 & ~w10093;
assign w10750 = ~w10025 & w10071;
assign w10751 = ~w10014 & w10750;
assign w10752 = w10050 & w10749;
assign w10753 = w10100 & w10749;
assign w10754 = (~w10752 & w10751) | (~w10752 & w40891) | (w10751 & w40891);
assign w10755 = (~w3242 & w10396) | (~w3242 & w44459) | (w10396 & w44459);
assign w10756 = ~w10058 & w10754;
assign w10757 = w10419 & w10756;
assign w10758 = ~w10755 & ~w10757;
assign w10759 = w10036 & w10091;
assign w10760 = ~w2896 & ~w10759;
assign w10761 = ~w10757 & w44460;
assign w10762 = ~w2896 & w10759;
assign w10763 = (w10762 & w10757) | (w10762 & w44461) | (w10757 & w44461);
assign w10764 = ~w10761 & ~w10763;
assign w10765 = ~w9851 & ~w10390;
assign w10766 = w10765 & w52231;
assign w10767 = (w10074 & w44462) | (w10074 & w44463) | (w44462 & w44463);
assign w10768 = ~w10766 & ~w10767;
assign w10769 = ~w2285 & w52232;
assign w10770 = w10419 & ~w10768;
assign w10771 = w10769 & ~w10770;
assign w10772 = ~w10086 & ~w10389;
assign w10773 = w10091 & w10101;
assign w10774 = (w10772 & w10074) | (w10772 & w40894) | (w10074 & w40894);
assign w10775 = ~w10074 & w40895;
assign w10776 = ~w10774 & ~w10775;
assign w10777 = (w10085 & w10396) | (w10085 & w40896) | (w10396 & w40896);
assign w10778 = w10419 & ~w10776;
assign w10779 = ~w10777 & ~w10778;
assign w10780 = (w2558 & w10778) | (w2558 & w40897) | (w10778 & w40897);
assign w10781 = ~w10771 & ~w10780;
assign w10782 = w10764 & w10781;
assign w10783 = w10764 & w40898;
assign w10784 = w10733 & w10783;
assign w10785 = ~w10050 & ~w10749;
assign w10786 = (w10785 & w10751) | (w10785 & w40899) | (w10751 & w40899);
assign w10787 = w10754 & ~w10786;
assign w10788 = (~w10057 & w10396) | (~w10057 & w40900) | (w10396 & w40900);
assign w10789 = w10419 & w10787;
assign w10790 = ~w10788 & ~w10789;
assign w10791 = w3242 & ~w10790;
assign w10792 = (w4056 & w10751) | (w4056 & w40901) | (w10751 & w40901);
assign w10793 = ~w10751 & w40902;
assign w10794 = ~w10792 & ~w10793;
assign w10795 = w3646 & w10049;
assign w10796 = (w10795 & ~w10419) | (w10795 & w40903) | (~w10419 & w40903);
assign w10797 = w3646 & ~w10049;
assign w10798 = w10419 & w40904;
assign w10799 = ~w10796 & ~w10798;
assign w10800 = w4430 & ~w10421;
assign w10801 = ~w4430 & w10421;
assign w10802 = ~w10800 & ~w10801;
assign w10803 = w10419 & ~w10802;
assign w10804 = w4056 & w10069;
assign w10805 = (w10804 & ~w10419) | (w10804 & w40905) | (~w10419 & w40905);
assign w10806 = w4056 & ~w10069;
assign w10807 = w10419 & w40906;
assign w10808 = ~w10805 & ~w10807;
assign w10809 = w10799 & ~w10808;
assign w10810 = ~w10789 & w40907;
assign w10811 = ~w3646 & ~w10049;
assign w10812 = (w10811 & ~w10419) | (w10811 & w40908) | (~w10419 & w40908);
assign w10813 = ~w3646 & w10049;
assign w10814 = w10419 & w40909;
assign w10815 = ~w10812 & ~w10814;
assign w10816 = ~w10810 & w10815;
assign w10817 = ~w10809 & w10816;
assign w10818 = ~w10791 & ~w10817;
assign w10819 = ~w10757 & w44464;
assign w10820 = w2896 & ~w10819;
assign w10821 = ~w10758 & w10759;
assign w10822 = w10820 & ~w10821;
assign w10823 = ~w10818 & ~w10822;
assign w10824 = ~w10778 & w40910;
assign w10825 = w10419 & w10768;
assign w10826 = (w9850 & w10396) | (w9850 & w40911) | (w10396 & w40911);
assign w10827 = w2285 & ~w10826;
assign w10828 = ~w10825 & w10827;
assign w10829 = ~w10824 & ~w10828;
assign w10830 = ~w10748 & ~w10771;
assign w10831 = ~w10829 & w10830;
assign w10832 = w10419 & w44465;
assign w10833 = w1738 & ~w10721;
assign w10834 = ~w10832 & w10833;
assign w10835 = (w2006 & w10745) | (w2006 & w44466) | (w10745 & w44466);
assign w10836 = ~w10834 & ~w10835;
assign w10837 = ~w10831 & w10836;
assign w10838 = w1320 & w10383;
assign w10839 = (w10838 & w10692) | (w10838 & w44467) | (w10692 & w44467);
assign w10840 = w1320 & w10707;
assign w10841 = ~w10839 & ~w10840;
assign w10842 = w1320 & w10718;
assign w10843 = w10706 & ~w10841;
assign w10844 = ~w10842 & ~w10843;
assign w10845 = w1541 & ~w10701;
assign w10846 = ~w10697 & w10845;
assign w10847 = w10844 & ~w10846;
assign w10848 = ~w10720 & ~w10847;
assign w10849 = ~w1320 & ~w10419;
assign w10850 = w10419 & w44468;
assign w10851 = ~w10849 & ~w10850;
assign w10852 = ~w9797 & ~w10377;
assign w10853 = ~w1120 & w10852;
assign w10854 = ~w10851 & w10853;
assign w10855 = ~w1120 & ~w10852;
assign w10856 = w10851 & w10855;
assign w10857 = ~w10854 & ~w10856;
assign w10858 = ~w10848 & w10857;
assign w10859 = w10733 & ~w10837;
assign w10860 = w10858 & ~w10859;
assign w10861 = w10784 & ~w10823;
assign w10862 = w10860 & ~w10861;
assign w10863 = w945 & w10678;
assign w10864 = w10851 & ~w10852;
assign w10865 = ~w10851 & w10852;
assign w10866 = ~w10864 & ~w10865;
assign w10867 = w1120 & w10866;
assign w10868 = ~w10863 & ~w10867;
assign w10869 = ~w10862 & w10868;
assign w10870 = w10686 & ~w10869;
assign w10871 = ~w9932 & w40912;
assign w10872 = (~w9996 & w10871) | (~w9996 & w44469) | (w10871 & w44469);
assign w10873 = ~w10218 & ~w10872;
assign w10874 = w10417 & ~w10872;
assign w10875 = (~w10873 & w10440) | (~w10873 & w40913) | (w10440 & w40913);
assign w10876 = ~w4838 & w10218;
assign w10877 = ~w10441 & w10876;
assign w10878 = w10875 & ~w10877;
assign w10879 = ~w10011 & ~w10063;
assign w10880 = w4430 & ~w10879;
assign w10881 = ~w10878 & w10880;
assign w10882 = w4430 & w10879;
assign w10883 = w10878 & w10882;
assign w10884 = ~w10881 & ~w10883;
assign w10885 = ~w9404 & ~w9781;
assign w10886 = w9781 & ~w9943;
assign w10887 = ~w10885 & ~w10886;
assign w10888 = w9981 & ~w10000;
assign w10889 = ~w9932 & w40914;
assign w10890 = w10019 & ~w10020;
assign w10891 = ~w10889 & w10890;
assign w10892 = w9948 & w9954;
assign w10893 = w10890 & w10892;
assign w10894 = ~w10889 & w10893;
assign w10895 = ~w9991 & ~w10892;
assign w10896 = ~w10891 & w10895;
assign w10897 = w9991 & w10892;
assign w10898 = ~w10894 & ~w10897;
assign w10899 = ~w10896 & w10898;
assign w10900 = ~w10396 & w40915;
assign w10901 = ~w4838 & ~w10900;
assign w10902 = ~w10419 & w10887;
assign w10903 = w10901 & ~w10902;
assign w10904 = w4838 & w10887;
assign w10905 = (w10904 & w10396) | (w10904 & w40916) | (w10396 & w40916);
assign w10906 = w4838 & ~w10899;
assign w10907 = w10419 & w10906;
assign w10908 = ~w10905 & ~w10907;
assign w10909 = ~w9991 & ~w10020;
assign w10910 = w10019 & ~w10889;
assign w10911 = w10909 & ~w10910;
assign w10912 = ~w10909 & w10910;
assign w10913 = ~w10911 & ~w10912;
assign w10914 = w5330 & w9990;
assign w10915 = (w10914 & w10396) | (w10914 & w40917) | (w10396 & w40917);
assign w10916 = w5330 & ~w10913;
assign w10917 = w10419 & w10916;
assign w10918 = ~w10915 & ~w10917;
assign w10919 = w10908 & ~w10918;
assign w10920 = ~w10903 & ~w10919;
assign w10921 = w10884 & w10920;
assign w10922 = ~w4056 & ~w10069;
assign w10923 = (w10922 & ~w10419) | (w10922 & w40918) | (~w10419 & w40918);
assign w10924 = ~w4056 & w10069;
assign w10925 = w10419 & w40919;
assign w10926 = ~w10923 & ~w10925;
assign w10927 = w10799 & w10926;
assign w10928 = ~w4430 & ~w10879;
assign w10929 = w10878 & w10928;
assign w10930 = ~w4430 & w10879;
assign w10931 = ~w10878 & w10930;
assign w10932 = ~w10929 & ~w10931;
assign w10933 = w10927 & w10932;
assign w10934 = ~w10791 & w10933;
assign w10935 = ~w10921 & w10934;
assign w10936 = a[62] & ~a[63];
assign w10937 = w10218 & w10936;
assign w10938 = ~w10104 & w40920;
assign w10939 = ~w9781 & w9868;
assign w10940 = w10146 & w10939;
assign w10941 = ~w10217 & w10939;
assign w10942 = ~w10197 & w10940;
assign w10943 = ~w10941 & ~w10942;
assign w10944 = ~a[63] & ~w9781;
assign w10945 = ~w10942 & w40921;
assign w10946 = ~w10417 & w10937;
assign w10947 = a[63] & ~w10943;
assign w10948 = ~w10946 & ~w10947;
assign w10949 = w10394 & w10945;
assign w10950 = ~w10104 & w10949;
assign w10951 = w10948 & ~w10950;
assign w10952 = w10196 & ~w10410;
assign w10953 = w10146 & ~w10952;
assign w10954 = w10217 & ~w10953;
assign w10955 = w10575 & ~w10954;
assign w10956 = w9868 & w10955;
assign w10957 = a[63] & w10940;
assign w10958 = w10597 & w10957;
assign w10959 = ~w10440 & w10958;
assign w10960 = w10945 & ~w10956;
assign w10961 = ~w10959 & ~w10960;
assign w10962 = ~w9869 & ~w9871;
assign w10963 = w9781 & ~w10962;
assign w10964 = ~a[63] & w10003;
assign w10965 = w10963 & ~w10964;
assign w10966 = w10218 & ~w10369;
assign w10967 = w10434 & w10966;
assign w10968 = ~w10425 & w10967;
assign w10969 = ~w10418 & ~w10968;
assign w10970 = ~a[62] & a[63];
assign w10971 = w9781 & w10970;
assign w10972 = (w10971 & w10968) | (w10971 & w40922) | (w10968 & w40922);
assign w10973 = ~w10396 & w40923;
assign w10974 = ~w10972 & ~w10973;
assign w10975 = ~w10938 & w10951;
assign w10976 = w10961 & w10975;
assign w10977 = w10974 & w10976;
assign w10978 = a[62] & ~w9864;
assign w10979 = ~w9865 & ~w10978;
assign w10980 = ~w10218 & w10979;
assign w10981 = w10394 & ~w10980;
assign w10982 = ~w10104 & w10981;
assign w10983 = a[62] & ~w9781;
assign w10984 = ~a[62] & w9781;
assign w10985 = ~w10983 & ~w10984;
assign w10986 = w10218 & w10985;
assign w10987 = ~w10955 & w10986;
assign w10988 = w10394 & w10986;
assign w10989 = ~w10104 & w10988;
assign w10990 = ~w10987 & ~w10989;
assign w10991 = ~w10418 & w10979;
assign w10992 = ~w10982 & w10991;
assign w10993 = w10990 & ~w10992;
assign w10994 = ~a[58] & ~a[59];
assign w10995 = ~a[60] & w10994;
assign w10996 = ~w9781 & ~w10995;
assign w10997 = a[61] & ~w10996;
assign w10998 = w9781 & w10995;
assign w10999 = a[60] & ~a[61];
assign w11000 = ~w10998 & ~w10999;
assign w11001 = ~a[61] & ~w10996;
assign w11002 = ~w10998 & ~w11001;
assign w11003 = (w11002 & w10968) | (w11002 & w40924) | (w10968 & w40924);
assign w11004 = ~w10997 & w11000;
assign w11005 = ~w10968 & w40925;
assign w11006 = ~w11003 & ~w11005;
assign w11007 = w9195 & w10993;
assign w11008 = w11006 & ~w11007;
assign w11009 = ~w9195 & ~w10993;
assign w11010 = ~w11008 & ~w11009;
assign w11011 = (w8666 & ~w10976) | (w8666 & w40926) | (~w10976 & w40926);
assign w11012 = w11010 & ~w11011;
assign w11013 = ~w10936 & ~w10970;
assign w11014 = ~w8666 & w11013;
assign w11015 = ~w10944 & w11014;
assign w11016 = ~w9781 & ~w9871;
assign w11017 = ~w10963 & ~w11016;
assign w11018 = ~w8666 & w11017;
assign w11019 = ~w10396 & w40927;
assign w11020 = a[63] & ~w8666;
assign w11021 = ~w9781 & w11020;
assign w11022 = w10943 & w11021;
assign w11023 = (w11022 & w10440) | (w11022 & w40928) | (w10440 & w40928);
assign w11024 = ~w11019 & ~w11023;
assign w11025 = ~w10419 & w11015;
assign w11026 = w11024 & ~w11025;
assign w11027 = ~w9894 & ~w9929;
assign w11028 = ~w9914 & w11027;
assign w11029 = ~w10218 & w11028;
assign w11030 = w10394 & ~w11029;
assign w11031 = ~w10418 & w11028;
assign w11032 = ~w10104 & w11030;
assign w11033 = ~w7315 & w9927;
assign w11034 = (w11033 & w11032) | (w11033 & w40929) | (w11032 & w40929);
assign w11035 = ~w7315 & ~w9927;
assign w11036 = ~w11032 & w40930;
assign w11037 = ~w11034 & ~w11036;
assign w11038 = w9928 & w11027;
assign w11039 = ~w9894 & ~w11038;
assign w11040 = w7315 & ~w11039;
assign w11041 = ~w7315 & w11039;
assign w11042 = ~w11040 & ~w11041;
assign w11043 = ~w10418 & w11042;
assign w11044 = ~w10396 & w11043;
assign w11045 = w6769 & ~w9898;
assign w11046 = (w11045 & w10396) | (w11045 & w40931) | (w10396 & w40931);
assign w11047 = w6769 & w9898;
assign w11048 = ~w10396 & w40932;
assign w11049 = ~w11046 & ~w11048;
assign w11050 = w11037 & w11049;
assign w11051 = w8666 & w9876;
assign w11052 = ~w8666 & ~w9876;
assign w11053 = ~w11051 & ~w11052;
assign w11054 = ~w10418 & w11053;
assign w11055 = ~w10396 & w11054;
assign w11056 = w9781 & w9878;
assign w11057 = ~w9781 & w9881;
assign w11058 = ~w11056 & ~w11057;
assign w11059 = w11055 & w11058;
assign w11060 = ~w11055 & ~w11058;
assign w11061 = ~w11059 & ~w11060;
assign w11062 = ~w7924 & w11061;
assign w11063 = w11026 & w11050;
assign w11064 = ~w11062 & w11063;
assign w11065 = ~w11012 & w11064;
assign w11066 = w7315 & ~w9927;
assign w11067 = (w11066 & w11032) | (w11066 & w40933) | (w11032 & w40933);
assign w11068 = w7315 & w9927;
assign w11069 = ~w11032 & w40934;
assign w11070 = ~w11067 & ~w11069;
assign w11071 = w7924 & ~w11058;
assign w11072 = (w11071 & w10396) | (w11071 & w40935) | (w10396 & w40935);
assign w11073 = w7924 & w11058;
assign w11074 = ~w10396 & w40936;
assign w11075 = ~w11072 & ~w11074;
assign w11076 = w11070 & w11075;
assign w11077 = w11050 & ~w11076;
assign w11078 = ~w6264 & w10218;
assign w11079 = w10394 & w11078;
assign w11080 = ~w10104 & w11079;
assign w11081 = ~w6264 & w10418;
assign w11082 = ~w11080 & ~w11081;
assign w11083 = ~w10418 & w10871;
assign w11084 = ~w10396 & w11083;
assign w11085 = w11082 & ~w11084;
assign w11086 = w9981 & w10019;
assign w11087 = ~w5745 & w11086;
assign w11088 = ~w11085 & w11087;
assign w11089 = ~w5745 & ~w11086;
assign w11090 = w11085 & w11089;
assign w11091 = ~w11088 & ~w11090;
assign w11092 = (w9912 & w11038) | (w9912 & w40937) | (w11038 & w40937);
assign w11093 = w9907 & ~w10000;
assign w11094 = w11092 & ~w11093;
assign w11095 = ~w11092 & w11093;
assign w11096 = ~w11094 & ~w11095;
assign w11097 = w9999 & w10218;
assign w11098 = w10394 & w11097;
assign w11099 = ~w10104 & w11098;
assign w11100 = w9999 & w10418;
assign w11101 = ~w11099 & ~w11100;
assign w11102 = ~w10418 & w11096;
assign w11103 = ~w10396 & w11102;
assign w11104 = w11101 & ~w11103;
assign w11105 = w6264 & w11104;
assign w11106 = ~w6769 & w9898;
assign w11107 = (w11106 & w10396) | (w11106 & w40938) | (w10396 & w40938);
assign w11108 = ~w6769 & ~w9898;
assign w11109 = ~w10396 & w40939;
assign w11110 = ~w11107 & ~w11109;
assign w11111 = ~w11105 & w11110;
assign w11112 = w11091 & w11111;
assign w11113 = ~w11077 & w11112;
assign w11114 = ~w11065 & w11113;
assign w11115 = w11085 & ~w11086;
assign w11116 = ~w11085 & w11086;
assign w11117 = ~w11115 & ~w11116;
assign w11118 = w5745 & w11117;
assign w11119 = ~w6264 & ~w11104;
assign w11120 = w11091 & w11119;
assign w11121 = ~w11118 & ~w11120;
assign w11122 = ~w5330 & ~w9990;
assign w11123 = (w11122 & w10396) | (w11122 & w40940) | (w10396 & w40940);
assign w11124 = ~w5330 & w10913;
assign w11125 = w10419 & w11124;
assign w11126 = ~w11123 & ~w11125;
assign w11127 = w10908 & w11126;
assign w11128 = ~w10903 & ~w11127;
assign w11129 = w10884 & w11128;
assign w11130 = w11121 & ~w11129;
assign w11131 = w10934 & w11130;
assign w11132 = ~w11114 & w11131;
assign w11133 = ~w10935 & ~w11132;
assign w11134 = w10784 & ~w10867;
assign w11135 = ~w10863 & w11134;
assign w11136 = ~w11133 & w11135;
assign w11137 = w10870 & ~w11136;
assign w11138 = w10673 & ~w11137;
assign w11139 = ~w10869 & ~w11136;
assign w11140 = w10684 & w44470;
assign w11141 = ~w10559 & ~w10571;
assign w11142 = ~w10559 & w40942;
assign w11143 = (~w11142 & w11136) | (~w11142 & w48733) | (w11136 & w48733);
assign w11144 = ~w11138 & w11143;
assign w11145 = (w10464 & w11144) | (w10464 & w44472) | (w11144 & w44472);
assign w11146 = ~w11144 & w44473;
assign w11147 = ~w11145 & ~w11146;
assign w11148 = w80 & w11147;
assign w11149 = ~w80 & ~w11147;
assign w11150 = w10530 & w10564;
assign w11151 = ~w10500 & w10557;
assign w11152 = w10517 & w10557;
assign w11153 = ~w11151 & w50186;
assign w11154 = ~w11137 & w48734;
assign w11155 = (w10569 & w11137) | (w10569 & w44475) | (w11137 & w44475);
assign w11156 = w11153 & w11155;
assign w11157 = (w11150 & w11156) | (w11150 & w48735) | (w11156 & w48735);
assign w11158 = ~w11156 & w48736;
assign w11159 = ~w11157 & ~w11158;
assign w11160 = w252 & w11159;
assign w11161 = ~w10518 & ~w10546;
assign w11162 = (w11161 & w11136) | (w11161 & w44476) | (w11136 & w44476);
assign w11163 = ~w11137 & w47269;
assign w11164 = ~w11138 & w11162;
assign w11165 = ~w11163 & ~w11164;
assign w11166 = w10556 & w10569;
assign w11167 = (~w11166 & w11164) | (~w11166 & w47270) | (w11164 & w47270);
assign w11168 = ~w351 & ~w11167;
assign w11169 = w11165 & w11166;
assign w11170 = w11168 & ~w11169;
assign w11171 = ~w11160 & ~w11170;
assign w11172 = w10483 & ~w10673;
assign w11173 = ~w11137 & ~w11172;
assign w11174 = (w10517 & w11136) | (w10517 & w44477) | (w11136 & w44477);
assign w11175 = ~w11173 & ~w11174;
assign w11176 = ~w11137 & w44478;
assign w11177 = ~w11175 & ~w11176;
assign w11178 = ~w10499 & ~w10546;
assign w11179 = ~w400 & w11178;
assign w11180 = (w11179 & w11175) | (w11179 & w44479) | (w11175 & w44479);
assign w11181 = ~w400 & ~w11178;
assign w11182 = ~w11175 & w44480;
assign w11183 = ~w11180 & ~w11182;
assign w11184 = w351 & ~w11166;
assign w11185 = (w11184 & w11164) | (w11184 & w47271) | (w11164 & w47271);
assign w11186 = w351 & w11166;
assign w11187 = ~w11164 & w47272;
assign w11188 = ~w11185 & ~w11187;
assign w11189 = w11183 & w11188;
assign w11190 = w400 & ~w11178;
assign w11191 = (w11190 & w11175) | (w11190 & w44481) | (w11175 & w44481);
assign w11192 = w400 & w11178;
assign w11193 = ~w11175 & w44482;
assign w11194 = ~w11191 & ~w11193;
assign w11195 = w10483 & w10509;
assign w11196 = (w10516 & w11136) | (w10516 & w44483) | (w11136 & w44483);
assign w11197 = ~w11195 & ~w11196;
assign w11198 = w10516 & w11195;
assign w11199 = (w11198 & w11136) | (w11198 & w44484) | (w11136 & w44484);
assign w11200 = ~w10472 & ~w10473;
assign w11201 = w10474 & ~w11200;
assign w11202 = ~w10474 & w11200;
assign w11203 = ~w11201 & ~w11202;
assign w11204 = w11138 & ~w11203;
assign w11205 = ~w11138 & ~w11199;
assign w11206 = ~w11197 & w11205;
assign w11207 = ~w11206 & w47273;
assign w11208 = w11194 & ~w11207;
assign w11209 = w11189 & ~w11208;
assign w11210 = w11171 & ~w11209;
assign w11211 = ~w252 & ~w11159;
assign w11212 = w57 & ~w11211;
assign w11213 = ~w11210 & w11212;
assign w11214 = ~w10069 & ~w10803;
assign w11215 = w10069 & w10803;
assign w11216 = ~w11214 & ~w11215;
assign w11217 = w10808 & w10926;
assign w11218 = w10921 & w11113;
assign w11219 = ~w11065 & w11218;
assign w11220 = w10921 & w11120;
assign w11221 = ~w11219 & ~w11220;
assign w11222 = ~w11118 & w11127;
assign w11223 = w10921 & ~w11222;
assign w11224 = w10932 & ~w11223;
assign w11225 = w11221 & w11224;
assign w11226 = w11217 & ~w11225;
assign w11227 = ~w11217 & w11225;
assign w11228 = ~w11226 & ~w11227;
assign w11229 = w11138 & ~w11216;
assign w11230 = ~w11138 & w11228;
assign w11231 = ~w11229 & ~w11230;
assign w11232 = w3646 & ~w11231;
assign w11233 = w11112 & w40945;
assign w11234 = ~w11065 & w11233;
assign w11235 = ~w5330 & ~w11121;
assign w11236 = w9990 & ~w10419;
assign w11237 = w10419 & ~w10913;
assign w11238 = ~w11236 & ~w11237;
assign w11239 = (~w11238 & w11121) | (~w11238 & w40946) | (w11121 & w40946);
assign w11240 = ~w11234 & w11239;
assign w11241 = w5330 & w11121;
assign w11242 = (~w10903 & ~w11121) | (~w10903 & w40947) | (~w11121 & w40947);
assign w11243 = w11112 & w40948;
assign w11244 = ~w11065 & w11243;
assign w11245 = ~w11242 & ~w11244;
assign w11246 = ~w11240 & ~w11245;
assign w11247 = w10884 & w10932;
assign w11248 = w10908 & ~w11247;
assign w11249 = ~w11246 & w11248;
assign w11250 = ~w10673 & ~w11249;
assign w11251 = ~w11136 & ~w11249;
assign w11252 = w10870 & w11251;
assign w11253 = ~w11250 & ~w11252;
assign w11254 = w10908 & ~w11246;
assign w11255 = w11247 & ~w11254;
assign w11256 = w10878 & ~w10879;
assign w11257 = ~w10878 & w10879;
assign w11258 = ~w11256 & ~w11257;
assign w11259 = ~w4056 & ~w11258;
assign w11260 = w11138 & w11259;
assign w11261 = ~w4056 & ~w11255;
assign w11262 = ~w11253 & w11261;
assign w11263 = ~w11260 & ~w11262;
assign w11264 = ~w11114 & w11241;
assign w11265 = ~w11240 & ~w11264;
assign w11266 = ~w10903 & w10908;
assign w11267 = w11265 & ~w11266;
assign w11268 = ~w11265 & w11266;
assign w11269 = ~w11267 & ~w11268;
assign w11270 = ~w11138 & w11269;
assign w11271 = ~w5330 & ~w10419;
assign w11272 = ~w9991 & ~w10891;
assign w11273 = w10419 & w11272;
assign w11274 = ~w11271 & ~w11273;
assign w11275 = w10892 & w11274;
assign w11276 = ~w10892 & ~w11274;
assign w11277 = ~w11275 & ~w11276;
assign w11278 = w11246 & w11277;
assign w11279 = ~w11136 & ~w11278;
assign w11280 = ~w10673 & ~w11246;
assign w11281 = w11277 & ~w11280;
assign w11282 = w10870 & w11279;
assign w11283 = w11281 & ~w11282;
assign w11284 = (~w4430 & w11282) | (~w4430 & w40949) | (w11282 & w40949);
assign w11285 = ~w11270 & w11284;
assign w11286 = w11263 & ~w11285;
assign w11287 = ~w11282 & w40950;
assign w11288 = w4430 & w11269;
assign w11289 = ~w11138 & w11288;
assign w11290 = ~w11287 & ~w11289;
assign w11291 = ~w11234 & ~w11235;
assign w11292 = ~w11264 & w11291;
assign w11293 = w10673 & w11292;
assign w11294 = ~w11137 & w11293;
assign w11295 = w11238 & ~w11292;
assign w11296 = w11240 & ~w11264;
assign w11297 = ~w11295 & ~w11296;
assign w11298 = w4838 & w11238;
assign w11299 = ~w11137 & w50300;
assign w11300 = (w4838 & w11295) | (w4838 & w50301) | (w11295 & w50301);
assign w11301 = ~w11294 & w11300;
assign w11302 = ~w11299 & ~w11301;
assign w11303 = w11290 & ~w11302;
assign w11304 = ~w11077 & w11110;
assign w11305 = (w11304 & w11012) | (w11304 & w50510) | (w11012 & w50510);
assign w11306 = w11091 & ~w11118;
assign w11307 = ~w11119 & ~w11306;
assign w11308 = ~w11105 & w11305;
assign w11309 = w11307 & ~w11308;
assign w11310 = w5745 & ~w11309;
assign w11311 = ~w11114 & ~w11120;
assign w11312 = ~w11309 & w11311;
assign w11313 = (w11312 & w11137) | (w11312 & w50511) | (w11137 & w50511);
assign w11314 = w11117 & w52233;
assign w11315 = ~w11313 & ~w11314;
assign w11316 = w5330 & w11315;
assign w11317 = ~w4838 & w11297;
assign w11318 = ~w11294 & w11317;
assign w11319 = ~w4838 & ~w11238;
assign w11320 = w11294 & w11319;
assign w11321 = ~w11318 & ~w11320;
assign w11322 = w11290 & w11321;
assign w11323 = w11286 & ~w11322;
assign w11324 = (~w11255 & w11252) | (~w11255 & w40951) | (w11252 & w40951);
assign w11325 = w11138 & ~w11258;
assign w11326 = ~w11324 & ~w11325;
assign w11327 = w4056 & w11326;
assign w11328 = ~w3646 & w11231;
assign w11329 = ~w11327 & ~w11328;
assign w11330 = ~w11323 & w11329;
assign w11331 = w11286 & w50303;
assign w11332 = w11330 & ~w11331;
assign w11333 = w10799 & w10815;
assign w11334 = (w10808 & ~w11221) | (w10808 & w40953) | (~w11221 & w40953);
assign w11335 = ~w10673 & ~w11334;
assign w11336 = ~w11136 & ~w11334;
assign w11337 = (~w11335 & ~w11336) | (~w11335 & w40954) | (~w11336 & w40954);
assign w11338 = ~w3646 & w10673;
assign w11339 = ~w11137 & w11338;
assign w11340 = w11337 & ~w11339;
assign w11341 = (~w3242 & ~w11340) | (~w3242 & w48737) | (~w11340 & w48737);
assign w11342 = w11333 & ~w11340;
assign w11343 = w11341 & ~w11342;
assign w11344 = (w11330 & w50304) | (w11330 & w50305) | (w50304 & w50305);
assign w11345 = ~w10791 & ~w10810;
assign w11346 = ~w10809 & w10815;
assign w11347 = (w11221 & w44485) | (w11221 & w44486) | (w44485 & w44486);
assign w11348 = ~w11345 & w52234;
assign w11349 = ~w11347 & ~w11348;
assign w11350 = ~w11137 & w44487;
assign w11351 = (~w11349 & w11137) | (~w11349 & w44488) | (w11137 & w44488);
assign w11352 = ~w11350 & ~w11351;
assign w11353 = ~w2896 & ~w11352;
assign w11354 = w3242 & w11333;
assign w11355 = ~w11340 & w11354;
assign w11356 = w3242 & ~w11333;
assign w11357 = w11340 & w11356;
assign w11358 = ~w11355 & ~w11357;
assign w11359 = ~w11353 & w11358;
assign w11360 = w10823 & ~w10935;
assign w11361 = (w10764 & w11132) | (w10764 & w40957) | (w11132 & w40957);
assign w11362 = ~w10771 & ~w10828;
assign w11363 = ~w10780 & w11362;
assign w11364 = (w11363 & w11361) | (w11363 & w44489) | (w11361 & w44489);
assign w11365 = ~w10824 & ~w11362;
assign w11366 = (w11365 & ~w11361) | (w11365 & w44490) | (~w11361 & w44490);
assign w11367 = ~w11364 & ~w11366;
assign w11368 = ~w11138 & w11367;
assign w11369 = ~w10825 & ~w10826;
assign w11370 = w10673 & w11369;
assign w11371 = ~w11137 & w11370;
assign w11372 = (~w2006 & w11137) | (~w2006 & w44491) | (w11137 & w44491);
assign w11373 = ~w11368 & w11372;
assign w11374 = ~w10748 & ~w10835;
assign w11375 = ~w10771 & ~w10829;
assign w11376 = (w10782 & w11132) | (w10782 & w40958) | (w11132 & w40958);
assign w11377 = (w11374 & w11376) | (w11374 & w44492) | (w11376 & w44492);
assign w11378 = ~w11376 & w44493;
assign w11379 = ~w11377 & ~w11378;
assign w11380 = ~w11138 & w11379;
assign w11381 = w10673 & ~w10747;
assign w11382 = ~w11137 & w11381;
assign w11383 = (~w1738 & w11137) | (~w1738 & w44494) | (w11137 & w44494);
assign w11384 = ~w11380 & w11383;
assign w11385 = ~w11373 & ~w11384;
assign w11386 = ~w10647 & w44495;
assign w11387 = ~w11137 & w11386;
assign w11388 = ~w10818 & ~w10935;
assign w11389 = ~w11132 & w11388;
assign w11390 = ~w10673 & w11389;
assign w11391 = w10686 & w11389;
assign w11392 = ~w10869 & w11391;
assign w11393 = w10764 & ~w10822;
assign w11394 = w2558 & w11393;
assign w11395 = ~w11392 & w40959;
assign w11396 = ~w11387 & w11395;
assign w11397 = w2558 & ~w11393;
assign w11398 = (w11397 & w11392) | (w11397 & w40960) | (w11392 & w40960);
assign w11399 = w11386 & w11397;
assign w11400 = ~w11137 & w11399;
assign w11401 = ~w11398 & ~w11400;
assign w11402 = ~w11396 & w11401;
assign w11403 = ~w10780 & ~w10824;
assign w11404 = w11361 & ~w11403;
assign w11405 = ~w11361 & w11403;
assign w11406 = ~w11404 & ~w11405;
assign w11407 = ~w2285 & ~w10779;
assign w11408 = ~w11137 & w44496;
assign w11409 = ~w2285 & w11406;
assign w11410 = ~w11138 & w11409;
assign w11411 = ~w11408 & ~w11410;
assign w11412 = w11402 & w11411;
assign w11413 = w11385 & w11412;
assign w11414 = w11359 & w11413;
assign w11415 = (w10783 & w11132) | (w10783 & w40961) | (w11132 & w40961);
assign w11416 = w10731 & w10837;
assign w11417 = ~w11415 & w11416;
assign w11418 = ~w10831 & ~w10835;
assign w11419 = w10731 & ~w10834;
assign w11420 = (~w11419 & w11415) | (~w11419 & w44497) | (w11415 & w44497);
assign w11421 = ~w10721 & ~w10832;
assign w11422 = ~w11417 & ~w11420;
assign w11423 = ~w11138 & w11422;
assign w11424 = (~w1541 & w11423) | (~w1541 & w44499) | (w11423 & w44499);
assign w11425 = ~w10703 & ~w10846;
assign w11426 = w10731 & ~w11425;
assign w11427 = ~w10731 & w11425;
assign w11428 = ~w11426 & ~w11427;
assign w11429 = ~w11415 & w44500;
assign w11430 = (~w11428 & w11415) | (~w11428 & w44501) | (w11415 & w44501);
assign w11431 = ~w11429 & ~w11430;
assign w11432 = ~w11137 & w44502;
assign w11433 = ~w11138 & w11431;
assign w11434 = (~w1320 & w11433) | (~w1320 & w44503) | (w11433 & w44503);
assign w11435 = ~w11424 & ~w11434;
assign w11436 = w11414 & w11435;
assign w11437 = ~w10862 & ~w10867;
assign w11438 = (w11134 & w11132) | (w11134 & w40962) | (w11132 & w40962);
assign w11439 = ~w11437 & ~w11438;
assign w11440 = ~w945 & w11439;
assign w11441 = w945 & ~w11439;
assign w11442 = ~w11440 & ~w11441;
assign w11443 = ~w11138 & ~w11442;
assign w11444 = ~w10678 & ~w11443;
assign w11445 = (~w10679 & ~w10673) | (~w10679 & w44504) | (~w10673 & w44504);
assign w11446 = w11139 & w11445;
assign w11447 = w945 & w11439;
assign w11448 = w11446 & ~w11447;
assign w11449 = (~w754 & ~w11446) | (~w754 & w44505) | (~w11446 & w44505);
assign w11450 = ~w11444 & w11449;
assign w11451 = ~w754 & w10673;
assign w11452 = ~w11137 & w11451;
assign w11453 = ~w11446 & ~w11452;
assign w11454 = w10516 & ~w10682;
assign w11455 = ~w612 & ~w11454;
assign w11456 = ~w11453 & w11455;
assign w11457 = ~w612 & w11454;
assign w11458 = w11453 & w11457;
assign w11459 = ~w11456 & ~w11458;
assign w11460 = ~w11450 & w11459;
assign w11461 = ~w10710 & ~w10718;
assign w11462 = ~w11137 & w44506;
assign w11463 = ~w10720 & w10844;
assign w11464 = ~w10703 & w10731;
assign w11465 = w10846 & ~w11463;
assign w11466 = ~w11463 & w11464;
assign w11467 = (w11466 & w11415) | (w11466 & w44507) | (w11415 & w44507);
assign w11468 = ~w11465 & ~w11467;
assign w11469 = ~w11138 & w11468;
assign w11470 = ~w10846 & w11463;
assign w11471 = (w11464 & w11415) | (w11464 & w44508) | (w11415 & w44508);
assign w11472 = w11470 & ~w11471;
assign w11473 = w1120 & w11462;
assign w11474 = w1120 & ~w11472;
assign w11475 = w11469 & w11474;
assign w11476 = ~w11473 & ~w11475;
assign w11477 = ~w10733 & ~w10848;
assign w11478 = ~w10848 & w11416;
assign w11479 = (~w11477 & w11415) | (~w11477 & w44509) | (w11415 & w44509);
assign w11480 = w10857 & ~w10867;
assign w11481 = w10686 & w10863;
assign w11482 = w10673 & ~w10866;
assign w11483 = ~w11481 & w11482;
assign w11484 = (~w11480 & ~w10673) | (~w11480 & w44510) | (~w10673 & w44510);
assign w11485 = w11479 & w11484;
assign w11486 = (w11480 & ~w10673) | (w11480 & w44511) | (~w10673 & w44511);
assign w11487 = ~w11479 & w11486;
assign w11488 = ~w11485 & ~w11487;
assign w11489 = ~w11483 & w11488;
assign w11490 = w945 & w11489;
assign w11491 = w11476 & ~w11490;
assign w11492 = w11460 & w11491;
assign w11493 = w11436 & w11492;
assign w11494 = w10673 & w40963;
assign w11495 = w11305 & ~w11494;
assign w11496 = w10673 & ~w11494;
assign w11497 = ~w11137 & w11496;
assign w11498 = ~w11495 & ~w11497;
assign w11499 = (w10784 & w11132) | (w10784 & w40964) | (w11132 & w40964);
assign w11500 = w10862 & ~w11499;
assign w11501 = (w11305 & w11500) | (w11305 & w44512) | (w11500 & w44512);
assign w11502 = w6264 & ~w10867;
assign w11503 = ~w11481 & w11502;
assign w11504 = ~w11501 & w11503;
assign w11505 = ~w11498 & ~w11504;
assign w11506 = ~w11105 & ~w11119;
assign w11507 = ~w5745 & ~w11506;
assign w11508 = (w11507 & w11498) | (w11507 & w44513) | (w11498 & w44513);
assign w11509 = ~w5745 & w11506;
assign w11510 = ~w11498 & w44514;
assign w11511 = ~w11508 & ~w11510;
assign w11512 = ~w9898 & ~w11044;
assign w11513 = w9898 & w11044;
assign w11514 = ~w11512 & ~w11513;
assign w11515 = ~w11062 & w11075;
assign w11516 = (w11026 & ~w11010) | (w11026 & w40965) | (~w11010 & w40965);
assign w11517 = w11515 & w11516;
assign w11518 = w11037 & w11076;
assign w11519 = (w11518 & ~w11516) | (w11518 & w44515) | (~w11516 & w44515);
assign w11520 = w11049 & w11110;
assign w11521 = w11037 & ~w11520;
assign w11522 = ~w11037 & w11520;
assign w11523 = ~w11521 & ~w11522;
assign w11524 = w11519 & w11520;
assign w11525 = ~w11519 & ~w11523;
assign w11526 = ~w11524 & ~w11525;
assign w11527 = ~w10673 & ~w11526;
assign w11528 = w10686 & ~w11526;
assign w11529 = (~w11527 & ~w11139) | (~w11527 & w40966) | (~w11139 & w40966);
assign w11530 = w10673 & w11514;
assign w11531 = ~w11137 & w11530;
assign w11532 = w11529 & ~w11531;
assign w11533 = ~w6264 & w11532;
assign w11534 = w11075 & ~w11517;
assign w11535 = ~w10673 & w11534;
assign w11536 = w10686 & w11534;
assign w11537 = ~w11136 & w40967;
assign w11538 = ~w11535 & ~w11537;
assign w11539 = ~w7315 & w10673;
assign w11540 = ~w11137 & w11539;
assign w11541 = w11538 & ~w11540;
assign w11542 = w11037 & w11070;
assign w11543 = w11541 & ~w11542;
assign w11544 = ~w11541 & w11542;
assign w11545 = ~w11543 & ~w11544;
assign w11546 = w6264 & ~w11532;
assign w11547 = (w6769 & w11532) | (w6769 & w7545) | (w11532 & w7545);
assign w11548 = (~w11533 & ~w11545) | (~w11533 & w44516) | (~w11545 & w44516);
assign w11549 = ~w6769 & w11542;
assign w11550 = ~w11541 & w11549;
assign w11551 = ~w6769 & ~w11542;
assign w11552 = w11541 & w11551;
assign w11553 = ~w11546 & ~w11552;
assign w11554 = ~w11550 & w11553;
assign w11555 = w11511 & w11554;
assign w11556 = ~w11515 & ~w11516;
assign w11557 = ~w11137 & w44517;
assign w11558 = ~w11517 & ~w11556;
assign w11559 = (w11558 & w11137) | (w11558 & w44518) | (w11137 & w44518);
assign w11560 = ~w11557 & ~w11559;
assign w11561 = w7315 & ~w11560;
assign w11562 = ~w7315 & w11560;
assign w11563 = w8666 & ~w11010;
assign w11564 = ~w8666 & w11010;
assign w11565 = ~w11563 & ~w11564;
assign w11566 = (w11565 & w11137) | (w11565 & w44519) | (w11137 & w44519);
assign w11567 = ~w7924 & w10977;
assign w11568 = ~w11566 & w11567;
assign w11569 = ~w7924 & ~w10977;
assign w11570 = w11566 & w11569;
assign w11571 = ~w11568 & ~w11570;
assign w11572 = ~w11562 & w11571;
assign w11573 = ~w11561 & ~w11572;
assign w11574 = w11511 & ~w11548;
assign w11575 = w11555 & w11573;
assign w11576 = ~w11574 & ~w11575;
assign w11577 = ~w5330 & ~w11315;
assign w11578 = w11286 & w50306;
assign w11579 = (w5745 & w11505) | (w5745 & w50307) | (w11505 & w50307);
assign w11580 = w11505 & w11506;
assign w11581 = w11579 & ~w11580;
assign w11582 = w11578 & w40968;
assign w11583 = w11576 & w11582;
assign w11584 = w10419 & w10997;
assign w11585 = ~w10969 & ~w11002;
assign w11586 = ~w11584 & ~w11585;
assign w11587 = w10969 & ~w11000;
assign w11588 = w11586 & ~w11587;
assign w11589 = ~w9195 & w11588;
assign w11590 = w9195 & ~w11588;
assign w11591 = ~w11589 & ~w11590;
assign w11592 = ~w10673 & ~w11591;
assign w11593 = (~w11591 & w11133) | (~w11591 & w40969) | (w11133 & w40969);
assign w11594 = w10870 & w11593;
assign w11595 = (w10993 & w11594) | (w10993 & w44520) | (w11594 & w44520);
assign w11596 = ~w11594 & w44521;
assign w11597 = ~w11595 & ~w11596;
assign w11598 = ~w8666 & w11597;
assign w11599 = w10685 & w44522;
assign w11600 = ~w11136 & w40970;
assign w11601 = (~a[59] & w10647) | (~a[59] & w40971) | (w10647 & w40971);
assign w11602 = ~a[56] & ~a[57];
assign w11603 = ~a[58] & w11602;
assign w11604 = ~w10419 & ~w11603;
assign w11605 = ~w9781 & w11604;
assign w11606 = ~w11601 & w11605;
assign w11607 = ~w11600 & w11606;
assign w11608 = w10419 & w11602;
assign w11609 = ~a[58] & w11608;
assign w11610 = ~w9781 & ~w11609;
assign w11611 = w10994 & w11610;
assign w11612 = ~w10673 & w11611;
assign w11613 = (w11611 & w11133) | (w11611 & w40972) | (w11133 & w40972);
assign w11614 = w10870 & w11613;
assign w11615 = ~w11612 & ~w11614;
assign w11616 = ~w11607 & w11615;
assign w11617 = ~a[60] & w10419;
assign w11618 = a[60] & ~w10419;
assign w11619 = ~w11617 & ~w11618;
assign w11620 = a[59] & w11610;
assign w11621 = w11619 & ~w11620;
assign w11622 = a[60] & ~w10994;
assign w11623 = ~w10995 & ~w11622;
assign w11624 = a[58] & ~a[59];
assign w11625 = w9781 & w11624;
assign w11626 = ~w11623 & ~w11625;
assign w11627 = ~w10673 & ~w11626;
assign w11628 = (~w11626 & w11133) | (~w11626 & w40973) | (w11133 & w40973);
assign w11629 = w10870 & w11628;
assign w11630 = ~w11627 & ~w11629;
assign w11631 = w10673 & w11621;
assign w11632 = ~w11137 & w11631;
assign w11633 = w11630 & ~w11632;
assign w11634 = w11616 & ~w11633;
assign w11635 = a[59] & w10673;
assign w11636 = ~w11137 & w11635;
assign w11637 = ~w11601 & ~w11604;
assign w11638 = ~w11601 & w44523;
assign w11639 = ~w11600 & w11638;
assign w11640 = ~w11636 & w11639;
assign w11641 = w9781 & w10419;
assign w11642 = ~w11603 & ~w11624;
assign w11643 = w11641 & ~w11642;
assign w11644 = ~w11640 & ~w11643;
assign w11645 = ~w11634 & w11644;
assign w11646 = ~w9195 & ~w11645;
assign w11647 = (w10661 & w10559) | (w10661 & w40974) | (w10559 & w40974);
assign w11648 = ~w9781 & ~w10419;
assign w11649 = ~w11641 & ~w11648;
assign w11650 = ~w10593 & w10661;
assign w11651 = w10644 & ~w11650;
assign w11652 = w10994 & ~w11649;
assign w11653 = w11651 & ~w11652;
assign w11654 = ~w11647 & w11653;
assign w11655 = w10685 & w11653;
assign w11656 = ~w11136 & w40975;
assign w11657 = ~w11654 & ~w11656;
assign w11658 = w10995 & ~w11649;
assign w11659 = w11651 & w11658;
assign w11660 = w10671 & w11617;
assign w11661 = ~w10671 & w11658;
assign w11662 = ~w11660 & ~w11661;
assign w11663 = ~w11659 & w11662;
assign w11664 = w10419 & ~w10671;
assign w11665 = ~w10419 & w10671;
assign w11666 = ~w11664 & ~w11665;
assign w11667 = ~w9781 & ~w10662;
assign w11668 = ~w11141 & ~w11666;
assign w11669 = w11667 & w11668;
assign w11670 = ~w11663 & ~w11669;
assign w11671 = w10685 & ~w11663;
assign w11672 = w11139 & w11671;
assign w11673 = ~w11670 & ~w11672;
assign w11674 = ~w10995 & w11649;
assign w11675 = ~w9781 & ~w10994;
assign w11676 = w11617 & w11675;
assign w11677 = a[61] & ~w11676;
assign w11678 = ~w11674 & w11677;
assign w11679 = w10673 & w11677;
assign w11680 = ~w11137 & w11679;
assign w11681 = ~w11678 & ~w11680;
assign w11682 = w11657 & ~w11673;
assign w11683 = ~w11681 & ~w11682;
assign w11684 = ~w11658 & ~w11674;
assign w11685 = ~a[61] & ~w11684;
assign w11686 = ~w11138 & w11685;
assign w11687 = ~a[61] & w11617;
assign w11688 = w11138 & w11687;
assign w11689 = ~w11686 & ~w11688;
assign w11690 = ~w11683 & w11689;
assign w11691 = w9195 & ~w11643;
assign w11692 = ~w11640 & w11691;
assign w11693 = ~w11634 & w11692;
assign w11694 = ~w11645 & w44524;
assign w11695 = w11690 & w40976;
assign w11696 = ~w11694 & ~w11695;
assign w11697 = w10977 & ~w11566;
assign w11698 = ~w10977 & w11566;
assign w11699 = ~w11697 & ~w11698;
assign w11700 = w7924 & w11699;
assign w11701 = w8666 & ~w11597;
assign w11702 = ~w11561 & ~w11701;
assign w11703 = ~w11700 & w11702;
assign w11704 = w11555 & w11703;
assign w11705 = w11696 & w11704;
assign w11706 = ~w11344 & w11493;
assign w11707 = w11493 & ~w11705;
assign w11708 = w11583 & w11707;
assign w11709 = ~w11706 & ~w11708;
assign w11710 = w11453 & ~w11454;
assign w11711 = ~w11453 & w11454;
assign w11712 = ~w11710 & ~w11711;
assign w11713 = w612 & ~w11712;
assign w11714 = ~w11423 & w44525;
assign w11715 = ~w11380 & ~w11382;
assign w11716 = (w1738 & w11380) | (w1738 & w44526) | (w11380 & w44526);
assign w11717 = ~w11714 & ~w11716;
assign w11718 = ~w2558 & ~w11393;
assign w11719 = ~w11392 & w40977;
assign w11720 = ~w11387 & w11719;
assign w11721 = ~w2558 & w11393;
assign w11722 = (w11721 & w11392) | (w11721 & w40978) | (w11392 & w40978);
assign w11723 = w11386 & w11721;
assign w11724 = ~w11137 & w11723;
assign w11725 = ~w11722 & ~w11724;
assign w11726 = ~w11720 & w11725;
assign w11727 = w2896 & w10790;
assign w11728 = ~w11137 & w44527;
assign w11729 = w2896 & w11349;
assign w11730 = ~w11138 & w11729;
assign w11731 = ~w11728 & ~w11730;
assign w11732 = w11726 & w11731;
assign w11733 = w11412 & ~w11732;
assign w11734 = ~w11368 & ~w11371;
assign w11735 = (w2006 & w11368) | (w2006 & w44528) | (w11368 & w44528);
assign w11736 = ~w11137 & w44529;
assign w11737 = ~w11138 & w11406;
assign w11738 = ~w11736 & ~w11737;
assign w11739 = ~w11737 & w44530;
assign w11740 = ~w11735 & ~w11739;
assign w11741 = ~w11733 & w11740;
assign w11742 = w11435 & ~w11717;
assign w11743 = w11385 & w11435;
assign w11744 = ~w11741 & w11743;
assign w11745 = (~w11742 & w11741) | (~w11742 & w44531) | (w11741 & w44531);
assign w11746 = ~w11460 & ~w11713;
assign w11747 = w11491 & ~w11746;
assign w11748 = ~w11745 & w11747;
assign w11749 = w11446 & w44532;
assign w11750 = w754 & ~w10678;
assign w11751 = ~w11443 & w11750;
assign w11752 = ~w11749 & ~w11751;
assign w11753 = ~w945 & ~w11489;
assign w11754 = w11752 & ~w11753;
assign w11755 = ~w11138 & w44533;
assign w11756 = ~w1120 & ~w11462;
assign w11757 = ~w11755 & w11756;
assign w11758 = ~w11433 & w44534;
assign w11759 = ~w11757 & ~w11758;
assign w11760 = w11754 & w11759;
assign w11761 = ~w11491 & w11754;
assign w11762 = w11460 & ~w11761;
assign w11763 = ~w11760 & w11762;
assign w11764 = (w493 & w11206) | (w493 & w44535) | (w11206 & w44535);
assign w11765 = w11194 & w11764;
assign w11766 = w11189 & ~w11765;
assign w11767 = w11189 & w44536;
assign w11768 = ~w11763 & w11767;
assign w11769 = ~w11748 & w11768;
assign w11770 = w11768 & w44537;
assign w11771 = (~w11213 & ~w11709) | (~w11213 & w44538) | (~w11709 & w44538);
assign w11772 = ~w10544 & ~w10592;
assign w11773 = w50186 & w50308;
assign w11774 = ~w252 & w11138;
assign w11775 = (w10530 & w11137) | (w10530 & w47274) | (w11137 & w47274);
assign w11776 = ~w11773 & w11775;
assign w11777 = ~w11774 & ~w11776;
assign w11778 = w11772 & ~w11777;
assign w11779 = ~w11772 & w11777;
assign w11780 = ~w11778 & ~w11779;
assign w11781 = ~w57 & w11210;
assign w11782 = (w11781 & w11708) | (w11781 & w50309) | (w11708 & w50309);
assign w11783 = (w11781 & ~w11768) | (w11781 & w50512) | (~w11768 & w50512);
assign w11784 = ~w57 & w11211;
assign w11785 = ~w11780 & ~w11784;
assign w11786 = (w11785 & w11769) | (w11785 & w44539) | (w11769 & w44539);
assign w11787 = ~w11782 & w11786;
assign w11788 = w11771 & ~w11787;
assign w11789 = ~w11149 & w52235;
assign w11790 = w10653 & w11138;
assign w11791 = (~w10463 & w10559) | (~w10463 & w44541) | (w10559 & w44541);
assign w11792 = ~w10461 & ~w10673;
assign w11793 = ~w11137 & ~w11792;
assign w11794 = (w11791 & w11136) | (w11791 & w48738) | (w11136 & w48738);
assign w11795 = ~w11793 & ~w11794;
assign w11796 = w10587 & ~w10653;
assign w11797 = ~w80 & w10673;
assign w11798 = ~w11793 & w48739;
assign w11799 = (w11796 & w11137) | (w11796 & w44542) | (w11137 & w44542);
assign w11800 = ~w11795 & w11799;
assign w11801 = ~w11798 & ~w11800;
assign w11802 = ~w11790 & w11801;
assign w11803 = (w3 & ~w11801) | (w3 & w44543) | (~w11801 & w44543);
assign w11804 = ~w3 & ~w11790;
assign w11805 = w11801 & w11804;
assign w11806 = (~w11713 & ~w11762) | (~w11713 & w44544) | (~w11762 & w44544);
assign w11807 = ~w11748 & w11806;
assign w11808 = ~w11148 & ~w11211;
assign w11809 = ~w57 & w11780;
assign w11810 = w11808 & ~w11809;
assign w11811 = w11171 & ~w11766;
assign w11812 = w11810 & ~w11811;
assign w11813 = w11807 & w11812;
assign w11814 = w11709 & w11813;
assign w11815 = ~w11210 & w11810;
assign w11816 = w10643 & ~w11650;
assign w11817 = ~w11647 & w11816;
assign w11818 = w10612 & ~w11817;
assign w11819 = ~w10612 & w11817;
assign w11820 = ~w11818 & ~w11819;
assign w11821 = w10685 & w11816;
assign w11822 = w11647 & w11821;
assign w11823 = ~w11136 & w40979;
assign w11824 = w11820 & ~w11823;
assign w11825 = ~w11820 & w11823;
assign w11826 = ~w11824 & ~w11825;
assign w11827 = ~w10630 & ~w11826;
assign w11828 = ~w42 & ~w11827;
assign w11829 = ~w10588 & ~w10653;
assign w11830 = ~w10653 & w11791;
assign w11831 = ~w11829 & ~w11830;
assign w11832 = w11140 & ~w11829;
assign w11833 = ~w11136 & w40980;
assign w11834 = ~w11831 & ~w11833;
assign w11835 = w10643 & w10658;
assign w11836 = ~w10673 & w11835;
assign w11837 = (w11835 & w11133) | (w11835 & w40981) | (w11133 & w40981);
assign w11838 = w10870 & w11837;
assign w11839 = ~w11836 & ~w11838;
assign w11840 = w10637 & ~w10638;
assign w11841 = ~w10637 & w10638;
assign w11842 = ~w11840 & ~w11841;
assign w11843 = w10673 & w11842;
assign w11844 = ~w11137 & w11843;
assign w11845 = w10673 & ~w11842;
assign w11846 = ~w11137 & w11845;
assign w11847 = w11839 & ~w11846;
assign w11848 = w11834 & ~w11847;
assign w11849 = ~w11834 & w11839;
assign w11850 = ~w11844 & w11849;
assign w11851 = ~w11848 & ~w11850;
assign w11852 = ~w11138 & w11826;
assign w11853 = (w42 & ~w11826) | (w42 & w40982) | (~w11826 & w40982);
assign w11854 = w11851 & w11853;
assign w11855 = ~w11828 & ~w11854;
assign w11856 = ~w11138 & w48740;
assign w11857 = w80 & ~w11856;
assign w11858 = ~w10464 & ~w11144;
assign w11859 = w11857 & ~w11858;
assign w11860 = w57 & ~w11859;
assign w11861 = ~w11780 & w11860;
assign w11862 = ~w11149 & ~w11803;
assign w11863 = ~w11861 & w11862;
assign w11864 = ~w11861 & w40983;
assign w11865 = ~w11815 & w11864;
assign w11866 = (w11865 & ~w11709) | (w11865 & w44545) | (~w11709 & w44545);
assign w11867 = ~w42 & w11851;
assign w11868 = ~w11805 & ~w11867;
assign w11869 = ~w11855 & ~w11868;
assign w11870 = (w11709 & w44546) | (w11709 & w44547) | (w44546 & w44547);
assign w11871 = ~w11803 & ~w11805;
assign w11872 = w11870 & w11871;
assign w11873 = w11805 & w11855;
assign w11874 = ~w11803 & ~w11873;
assign w11875 = ~w11802 & ~w11870;
assign w11876 = (w44540 & w50513) | (w44540 & w50514) | (w50513 & w50514);
assign w11877 = ~w11875 & ~w11876;
assign w11878 = w11789 & w11872;
assign w11879 = w11877 & ~w11878;
assign w11880 = ~w11815 & w11863;
assign w11881 = (w11880 & ~w11709) | (w11880 & w50515) | (~w11709 & w50515);
assign w11882 = ~w11805 & ~w11881;
assign w11883 = ~w11851 & ~w11882;
assign w11884 = w11827 & w11851;
assign w11885 = w11882 & w11884;
assign w11886 = ~w11883 & ~w11885;
assign w11887 = ~w42 & w11886;
assign w11888 = w11879 & w11887;
assign w11889 = ~w11695 & w44548;
assign w11890 = w11571 & ~w11700;
assign w11891 = w11889 & w11890;
assign w11892 = ~w11869 & ~w11891;
assign w11893 = ~w11815 & w40986;
assign w11894 = w7315 & w11869;
assign w11895 = (~w11894 & w11814) | (~w11894 & w40987) | (w11814 & w40987);
assign w11896 = w11571 & w11892;
assign w11897 = (w11896 & w11814) | (w11896 & w40988) | (w11814 & w40988);
assign w11898 = w11895 & ~w11897;
assign w11899 = ~w11561 & ~w11562;
assign w11900 = w11898 & ~w11899;
assign w11901 = ~w11898 & w11899;
assign w11902 = ~w11900 & ~w11901;
assign w11903 = ~w6769 & w11902;
assign w11904 = ~w11646 & ~w11693;
assign w11905 = ~w11869 & w11904;
assign w11906 = (w11709 & w44549) | (w11709 & w44550) | (w44549 & w44550);
assign w11907 = w11690 & ~w11906;
assign w11908 = ~w11690 & w11906;
assign w11909 = ~w11907 & ~w11908;
assign w11910 = w8666 & ~w11909;
assign w11911 = w11690 & ~w11693;
assign w11912 = ~w11646 & ~w11911;
assign w11913 = (w8666 & w11911) | (w8666 & w44551) | (w11911 & w44551);
assign w11914 = ~w11869 & ~w11913;
assign w11915 = ~w8666 & w11912;
assign w11916 = w11914 & ~w11915;
assign w11917 = ~w11815 & w40990;
assign w11918 = ~w11597 & w11916;
assign w11919 = (w11918 & w11814) | (w11918 & w40991) | (w11814 & w40991);
assign w11920 = w11597 & ~w11916;
assign w11921 = (~w11920 & w11814) | (~w11920 & w40992) | (w11814 & w40992);
assign w11922 = ~w11919 & w11921;
assign w11923 = ~w11889 & ~w11890;
assign w11924 = w11892 & ~w11923;
assign w11925 = ~w11815 & w40993;
assign w11926 = ~w11699 & w11869;
assign w11927 = (~w11926 & w11814) | (~w11926 & w40994) | (w11814 & w40994);
assign w11928 = ~w11866 & w11924;
assign w11929 = w11927 & ~w11928;
assign w11930 = (~w7315 & w11928) | (~w7315 & w40995) | (w11928 & w40995);
assign w11931 = ~w7924 & ~w11922;
assign w11932 = ~w11930 & ~w11931;
assign w11933 = ~w11928 & w40996;
assign w11934 = w7924 & w11922;
assign w11935 = ~w11930 & w11934;
assign w11936 = ~w11933 & ~w11935;
assign w11937 = w11910 & w11932;
assign w11938 = w11936 & ~w11937;
assign w11939 = (w6264 & w11902) | (w6264 & w7544) | (w11902 & w7544);
assign w11940 = ~a[54] & ~a[55];
assign w11941 = ~a[56] & w11940;
assign w11942 = w11138 & ~w11941;
assign w11943 = ~w11815 & w40997;
assign w11944 = a[57] & w11869;
assign w11945 = (~w11944 & w11814) | (~w11944 & w40998) | (w11814 & w40998);
assign w11946 = ~a[57] & ~w11869;
assign w11947 = (w11709 & w44552) | (w11709 & w44553) | (w44552 & w44553);
assign w11948 = w11945 & ~w11947;
assign w11949 = w11602 & ~w11869;
assign w11950 = (w11709 & w44554) | (w11709 & w44555) | (w44554 & w44555);
assign w11951 = w11945 & ~w11950;
assign w11952 = ~w11138 & w11940;
assign w11953 = ~a[56] & w11952;
assign w11954 = ~w11869 & w11952;
assign w11955 = (w11709 & w44556) | (w11709 & w44557) | (w44556 & w44557);
assign w11956 = ~w11953 & ~w11955;
assign w11957 = w11945 & w44558;
assign w11958 = ~w11951 & w11956;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = a[58] & ~w11602;
assign w11961 = ~w11603 & ~w11960;
assign w11962 = ~w11869 & w11961;
assign w11963 = (w11709 & w44559) | (w11709 & w44560) | (w44559 & w44560);
assign w11964 = a[58] & w11138;
assign w11965 = ~a[58] & ~w11138;
assign w11966 = w11869 & ~w11965;
assign w11967 = (~w11965 & w11854) | (~w11965 & w44561) | (w11854 & w44561);
assign w11968 = ~w11861 & w41003;
assign w11969 = ~w11964 & w11966;
assign w11970 = ~w11815 & w41004;
assign w11971 = (~w11969 & w11814) | (~w11969 & w41005) | (w11814 & w41005);
assign w11972 = ~w11963 & w11971;
assign w11973 = w10419 & ~w11972;
assign w11974 = ~w11959 & ~w11973;
assign w11975 = ~w10419 & w11138;
assign w11976 = w10419 & ~w11138;
assign w11977 = ~w11975 & ~w11976;
assign w11978 = w11603 & ~w11977;
assign w11979 = ~w11603 & w11977;
assign w11980 = ~w11978 & ~w11979;
assign w11981 = ~w11869 & w11980;
assign w11982 = (w11709 & w44562) | (w11709 & w44563) | (w44562 & w44563);
assign w11983 = ~a[59] & ~w11966;
assign w11984 = (w11983 & w11814) | (w11983 & w41007) | (w11814 & w41007);
assign w11985 = ~w11982 & w11984;
assign w11986 = ~w11965 & w11979;
assign w11987 = ~w11869 & ~w11986;
assign w11988 = (w11709 & w44564) | (w11709 & w44565) | (w44564 & w44565);
assign w11989 = ~w11866 & w11987;
assign w11990 = w11988 & ~w11989;
assign w11991 = w11868 & w11978;
assign w11992 = w42 & w11842;
assign w11993 = ~w11828 & ~w11992;
assign w11994 = w11138 & ~w11993;
assign w11995 = w11978 & ~w11994;
assign w11996 = ~w10419 & ~w11602;
assign w11997 = w11965 & w11996;
assign w11998 = a[59] & ~w11997;
assign w11999 = ~w11995 & w11998;
assign w12000 = ~w11991 & w11999;
assign w12001 = ~w11815 & w41009;
assign w12002 = (~w12000 & w11814) | (~w12000 & w41010) | (w11814 & w41010);
assign w12003 = w11984 & w44566;
assign w12004 = ~w9781 & ~w12002;
assign w12005 = ~w11990 & w12004;
assign w12006 = ~w12003 & ~w12005;
assign w12007 = w11971 & w44567;
assign w12008 = ~w12005 & w41011;
assign w12009 = ~w11974 & w12008;
assign w12010 = w11138 & w11619;
assign w12011 = ~w11138 & w11623;
assign w12012 = ~w12010 & ~w12011;
assign w12013 = ~w11600 & w11637;
assign w12014 = ~w11608 & ~w12013;
assign w12015 = ~w11138 & w11624;
assign w12016 = w12014 & ~w12015;
assign w12017 = ~w11609 & w11636;
assign w12018 = w9781 & ~w12017;
assign w12019 = ~w12016 & w12018;
assign w12020 = ~w9781 & w12017;
assign w12021 = w11616 & ~w12020;
assign w12022 = ~w12019 & w12021;
assign w12023 = ~w11869 & w12022;
assign w12024 = (w11709 & w44568) | (w11709 & w44569) | (w44568 & w44569);
assign w12025 = w12012 & ~w12024;
assign w12026 = ~w12012 & w12024;
assign w12027 = ~w12025 & ~w12026;
assign w12028 = ~w9195 & w12027;
assign w12029 = (~w12002 & w11989) | (~w12002 & w41013) | (w11989 & w41013);
assign w12030 = ~w11985 & ~w12029;
assign w12031 = ~w12029 & w44570;
assign w12032 = ~w12028 & ~w12031;
assign w12033 = ~w12009 & w12032;
assign w12034 = ~w8666 & w11909;
assign w12035 = w9195 & w12012;
assign w12036 = ~w12024 & w12035;
assign w12037 = w9195 & ~w12012;
assign w12038 = w12024 & w12037;
assign w12039 = ~w12036 & ~w12038;
assign w12040 = ~w11931 & w47275;
assign w12041 = ~w11934 & w12034;
assign w12042 = w12040 & ~w12041;
assign w12043 = (w11939 & ~w11938) | (w11939 & w44571) | (~w11938 & w44571);
assign w12044 = w11939 & w12042;
assign w12045 = ~w12033 & w12044;
assign w12046 = ~w12043 & ~w12045;
assign w12047 = ~w12007 & w12039;
assign w12048 = w12006 & w12047;
assign w12049 = ~w11974 & w12048;
assign w12050 = w9781 & w12039;
assign w12051 = w12030 & w12050;
assign w12052 = ~w11910 & ~w12028;
assign w12053 = ~w12051 & w12052;
assign w12054 = ~w12049 & w12053;
assign w12055 = w7545 & ~w11902;
assign w12056 = w6769 & w11545;
assign w12057 = ~w6769 & ~w11545;
assign w12058 = ~w12056 & ~w12057;
assign w12059 = (~w11573 & ~w11696) | (~w11573 & w41014) | (~w11696 & w41014);
assign w12060 = w6769 & ~w11870;
assign w12061 = w11870 & ~w12059;
assign w12062 = ~w12060 & ~w12061;
assign w12063 = w12058 & ~w12062;
assign w12064 = ~w12058 & w12062;
assign w12065 = ~w12063 & ~w12064;
assign w12066 = ~w12055 & ~w12065;
assign w12067 = w11932 & ~w12034;
assign w12068 = w12066 & w12067;
assign w12069 = ~w12054 & w12068;
assign w12070 = (~w6264 & ~w40996) | (~w6264 & w44572) | (~w40996 & w44572);
assign w12071 = ~w11935 & w12070;
assign w12072 = ~w11903 & w12071;
assign w12073 = w12066 & ~w12072;
assign w12074 = (~w12073 & w12054) | (~w12073 & w41015) | (w12054 & w41015);
assign w12075 = w12046 & w12074;
assign w12076 = ~w11575 & w44573;
assign w12077 = ~w5330 & ~w11869;
assign w12078 = w12076 & w41016;
assign w12079 = w5330 & ~w11869;
assign w12080 = (w12079 & ~w12076) | (w12079 & w41017) | (~w12076 & w41017);
assign w12081 = ~w12078 & ~w12080;
assign w12082 = ~w4838 & ~w11315;
assign w12083 = ~w12081 & w12082;
assign w12084 = ~w11866 & w12083;
assign w12085 = ~w4838 & w11315;
assign w12086 = ~w11815 & w41018;
assign w12087 = (w12086 & ~w11709) | (w12086 & w44574) | (~w11709 & w44574);
assign w12088 = w12081 & w12085;
assign w12089 = ~w12087 & ~w12088;
assign w12090 = ~w12084 & w12089;
assign w12091 = ~w4838 & ~w11577;
assign w12092 = ~w11705 & w12091;
assign w12093 = w4838 & w11315;
assign w12094 = ~w6027 & ~w11316;
assign w12095 = ~w12093 & ~w12094;
assign w12096 = ~w11869 & ~w12095;
assign w12097 = (w12096 & ~w12092) | (w12096 & w48741) | (~w12092 & w48741);
assign w12098 = w4838 & ~w11316;
assign w12099 = (w12098 & ~w12076) | (w12098 & w41019) | (~w12076 & w41019);
assign w12100 = w12097 & ~w12099;
assign w12101 = ~w11238 & w11294;
assign w12102 = ~w11294 & w11297;
assign w12103 = ~w12101 & ~w12102;
assign w12104 = w4430 & w12103;
assign w12105 = w12097 & w41020;
assign w12106 = ~w11866 & w12105;
assign w12107 = w4430 & ~w12103;
assign w12108 = (w12107 & ~w12097) | (w12107 & w41021) | (~w12097 & w41021);
assign w12109 = ~w11815 & w41022;
assign w12110 = (w12109 & ~w11709) | (w12109 & w44575) | (~w11709 & w44575);
assign w12111 = ~w12108 & ~w12110;
assign w12112 = ~w12106 & w12111;
assign w12113 = w12090 & w12112;
assign w12114 = (w11302 & w11315) | (w11302 & w41023) | (w11315 & w41023);
assign w12115 = w11321 & ~w12114;
assign w12116 = w4430 & ~w12115;
assign w12117 = ~w11316 & w11321;
assign w12118 = w12116 & ~w12117;
assign w12119 = ~w11705 & w12116;
assign w12120 = (~w12118 & ~w12119) | (~w12118 & w44576) | (~w12119 & w44576);
assign w12121 = ~w4430 & w11321;
assign w12122 = ~w12114 & w12121;
assign w12123 = ~w11270 & ~w11283;
assign w12124 = (~w12123 & w12114) | (~w12123 & w50310) | (w12114 & w50310);
assign w12125 = ~w11316 & w12121;
assign w12126 = w12124 & ~w12125;
assign w12127 = ~w11705 & w12124;
assign w12128 = (~w12126 & ~w12127) | (~w12126 & w44577) | (~w12127 & w44577);
assign w12129 = w12120 & ~w12128;
assign w12130 = ~w4056 & ~w11869;
assign w12131 = w12129 & w12130;
assign w12132 = ~w11866 & w12131;
assign w12133 = ~w11869 & ~w12122;
assign w12134 = ~w12125 & w12133;
assign w12135 = ~w11705 & w12133;
assign w12136 = w12076 & w12135;
assign w12137 = ~w12134 & ~w12136;
assign w12138 = ~w4056 & w12123;
assign w12139 = (w12138 & w12137) | (w12138 & w44578) | (w12137 & w44578);
assign w12140 = ~w11815 & w41024;
assign w12141 = (w12140 & ~w11709) | (w12140 & w44579) | (~w11709 & w44579);
assign w12142 = ~w12139 & ~w12141;
assign w12143 = ~w12132 & w12142;
assign w12144 = ~w4430 & ~w12103;
assign w12145 = w12097 & w41025;
assign w12146 = ~w11866 & w12145;
assign w12147 = ~w4430 & w12103;
assign w12148 = (w12147 & ~w12097) | (w12147 & w41026) | (~w12097 & w41026);
assign w12149 = ~w11815 & w41027;
assign w12150 = (w12149 & ~w11709) | (w12149 & w44580) | (~w11709 & w44580);
assign w12151 = ~w12148 & ~w12150;
assign w12152 = ~w12146 & w12151;
assign w12153 = w12143 & w12152;
assign w12154 = ~w12113 & w12153;
assign w12155 = (w12123 & w11866) | (w12123 & w41028) | (w11866 & w41028);
assign w12156 = w11870 & w12129;
assign w12157 = ~w12155 & ~w12156;
assign w12158 = w4056 & w12157;
assign w12159 = ~w12154 & ~w12158;
assign w12160 = w12120 & w12128;
assign w12161 = w4056 & ~w11870;
assign w12162 = w11870 & ~w12160;
assign w12163 = ~w12161 & ~w12162;
assign w12164 = w11263 & ~w11327;
assign w12165 = ~w3646 & w12164;
assign w12166 = w12163 & w12165;
assign w12167 = ~w3646 & ~w12164;
assign w12168 = ~w12163 & w12167;
assign w12169 = ~w12166 & ~w12168;
assign w12170 = w12159 & w12169;
assign w12171 = ~w12057 & ~w12059;
assign w12172 = ~w12056 & ~w12171;
assign w12173 = ~w11546 & ~w11869;
assign w12174 = ~w11533 & w12172;
assign w12175 = w12173 & ~w12174;
assign w12176 = w5745 & w11869;
assign w12177 = ~w11815 & w41029;
assign w12178 = ~w11866 & w12175;
assign w12179 = w11511 & ~w11581;
assign w12180 = ~w5330 & ~w12179;
assign w12181 = (w12180 & w12178) | (w12180 & w41031) | (w12178 & w41031);
assign w12182 = ~w5330 & w12179;
assign w12183 = ~w12178 & w41032;
assign w12184 = ~w12181 & ~w12183;
assign w12185 = w4838 & ~w11315;
assign w12186 = ~w11815 & w41033;
assign w12187 = (w12186 & ~w11709) | (w12186 & w44581) | (~w11709 & w44581);
assign w12188 = w12081 & w12185;
assign w12189 = ~w12187 & ~w12188;
assign w12190 = ~w12081 & w12093;
assign w12191 = ~w11866 & w12190;
assign w12192 = w12189 & ~w12191;
assign w12193 = w12152 & w12192;
assign w12194 = w12143 & w12193;
assign w12195 = w12184 & w12194;
assign w12196 = ~w11533 & ~w11546;
assign w12197 = w6264 & ~w11870;
assign w12198 = w11870 & w12172;
assign w12199 = ~w12197 & ~w12198;
assign w12200 = w12196 & ~w12199;
assign w12201 = ~w12196 & w12199;
assign w12202 = ~w12200 & ~w12201;
assign w12203 = w5745 & ~w12202;
assign w12204 = ~w4056 & w11869;
assign w12205 = (w11709 & w48742) | (w11709 & w48743) | (w48742 & w48743);
assign w12206 = ~w11869 & w12160;
assign w12207 = w12160 & w41035;
assign w12208 = w12164 & ~w12206;
assign w12209 = w11326 & ~w12205;
assign w12210 = w12205 & ~w12207;
assign w12211 = ~w12208 & w12210;
assign w12212 = ~w12209 & ~w12211;
assign w12213 = w3646 & w12212;
assign w12214 = ~w12203 & ~w12213;
assign w12215 = w12170 & ~w12195;
assign w12216 = w12214 & ~w12215;
assign w12217 = ~w12075 & w12216;
assign w12218 = (~w11332 & w41036) | (~w11332 & w41037) | (w41036 & w41037);
assign w12219 = w11436 & ~w11705;
assign w12220 = w11583 & w12219;
assign w12221 = ~w11744 & w41038;
assign w12222 = ~w12220 & w41039;
assign w12223 = w11476 & ~w11757;
assign w12224 = w12222 & ~w12223;
assign w12225 = ~w12222 & w12223;
assign w12226 = ~w12224 & ~w12225;
assign w12227 = ~w11462 & ~w11755;
assign w12228 = ~w11870 & w12227;
assign w12229 = w11870 & w12226;
assign w12230 = ~w12228 & ~w12229;
assign w12231 = (~w945 & w12229) | (~w945 & w44582) | (w12229 & w44582);
assign w12232 = ~w11744 & w44583;
assign w12233 = ~w12220 & w41040;
assign w12234 = ~w11490 & ~w11753;
assign w12235 = w11476 & ~w12234;
assign w12236 = ~w12233 & w12235;
assign w12237 = ~w11476 & w12234;
assign w12238 = (w12220 & w44584) | (w12220 & w44585) | (w44584 & w44585);
assign w12239 = ~w12236 & w12238;
assign w12240 = w11489 & ~w11870;
assign w12241 = w11870 & w12239;
assign w12242 = ~w12241 & w44586;
assign w12243 = ~w12231 & ~w12242;
assign w12244 = w11385 & ~w11741;
assign w12245 = ~w11716 & ~w12244;
assign w12246 = w11583 & ~w11705;
assign w12247 = (w11344 & ~w11583) | (w11344 & w50516) | (~w11583 & w50516);
assign w12248 = ~w11869 & ~w12245;
assign w12249 = w11414 & ~w11869;
assign w12250 = ~w12248 & w52236;
assign w12251 = ~w11815 & w41043;
assign w12252 = w1541 & w11869;
assign w12253 = ~w11866 & ~w12250;
assign w12254 = ~w11424 & ~w11714;
assign w12255 = w1320 & ~w12254;
assign w12256 = (w12255 & w12253) | (w12255 & w41045) | (w12253 & w41045);
assign w12257 = w1320 & w12254;
assign w12258 = ~w12253 & w41046;
assign w12259 = ~w12256 & ~w12258;
assign w12260 = ~w11424 & ~w11869;
assign w12261 = w11717 & ~w12244;
assign w12262 = w12260 & ~w12261;
assign w12263 = ~w11869 & w48744;
assign w12264 = ~w12262 & w52237;
assign w12265 = ~w11815 & w41048;
assign w12266 = w1320 & w11869;
assign w12267 = ~w11866 & ~w12264;
assign w12268 = ~w11434 & ~w11758;
assign w12269 = ~w1120 & ~w12268;
assign w12270 = (w12269 & w12267) | (w12269 & w41050) | (w12267 & w41050);
assign w12271 = ~w1120 & w12268;
assign w12272 = ~w12267 & w41051;
assign w12273 = ~w12270 & ~w12272;
assign w12274 = w12259 & w12273;
assign w12275 = w12243 & w12274;
assign w12276 = ~w11412 & ~w11739;
assign w12277 = w11359 & ~w12276;
assign w12278 = ~w11705 & w12277;
assign w12279 = w11583 & w12278;
assign w12280 = ~w11733 & ~w11739;
assign w12281 = ~w11373 & ~w11735;
assign w12282 = ~w12279 & w44587;
assign w12283 = (w12281 & w12279) | (w12281 & w44588) | (w12279 & w44588);
assign w12284 = ~w12282 & ~w12283;
assign w12285 = w11734 & ~w11870;
assign w12286 = w11870 & ~w12284;
assign w12287 = ~w12285 & ~w12286;
assign w12288 = w1738 & w12287;
assign w12289 = w1738 & ~w11735;
assign w12290 = ~w1738 & w11735;
assign w12291 = ~w12289 & ~w12290;
assign w12292 = ~w12281 & w12291;
assign w12293 = w12280 & w12291;
assign w12294 = (~w12292 & w12279) | (~w12292 & w44589) | (w12279 & w44589);
assign w12295 = w1738 & w12281;
assign w12296 = (w12295 & w12279) | (w12295 & w44590) | (w12279 & w44590);
assign w12297 = w12294 & ~w12296;
assign w12298 = w11870 & w12297;
assign w12299 = w11715 & ~w12298;
assign w12300 = ~w11715 & w12298;
assign w12301 = ~w12299 & ~w12300;
assign w12302 = w1541 & w12301;
assign w12303 = ~w12288 & ~w12302;
assign w12304 = w12275 & w12303;
assign w12305 = ~w1738 & ~w12287;
assign w12306 = w11402 & ~w11732;
assign w12307 = (w11402 & w11359) | (w11402 & w12306) | (w11359 & w12306);
assign w12308 = (~w12246 & w44591) | (~w12246 & w44592) | (w44591 & w44592);
assign w12309 = (w12246 & w44593) | (w12246 & w44594) | (w44593 & w44594);
assign w12310 = ~w12308 & ~w12309;
assign w12311 = w11870 & ~w12310;
assign w12312 = ~w2006 & ~w11738;
assign w12313 = ~w12311 & w12312;
assign w12314 = ~w2006 & w11738;
assign w12315 = w12311 & w12314;
assign w12316 = ~w12313 & ~w12315;
assign w12317 = ~w12305 & w12316;
assign w12318 = w11402 & w11726;
assign w12319 = ~w11731 & ~w11869;
assign w12320 = w11359 & ~w11869;
assign w12321 = (w12320 & w12246) | (w12320 & w41058) | (w12246 & w41058);
assign w12322 = ~w12319 & ~w12321;
assign w12323 = ~w11815 & w41059;
assign w12324 = ~w2558 & w11869;
assign w12325 = (~w12324 & w11814) | (~w12324 & w41060) | (w11814 & w41060);
assign w12326 = ~w11866 & ~w12322;
assign w12327 = w12325 & ~w12326;
assign w12328 = (w12318 & w12326) | (w12318 & w41061) | (w12326 & w41061);
assign w12329 = ~w12326 & w41062;
assign w12330 = ~w12328 & ~w12329;
assign w12331 = ~w12328 & w50311;
assign w12332 = (w2006 & w12311) | (w2006 & w48745) | (w12311 & w48745);
assign w12333 = w11738 & w12311;
assign w12334 = w12332 & ~w12333;
assign w12335 = ~w12331 & ~w12334;
assign w12336 = (w12317 & w12331) | (w12317 & w44595) | (w12331 & w44595);
assign w12337 = ~w11353 & w11731;
assign w12338 = w2558 & ~w12337;
assign w12339 = w12338 & w52238;
assign w12340 = w2558 & w12337;
assign w12341 = (w12246 & w44596) | (w12246 & w44597) | (w44596 & w44597);
assign w12342 = ~w12339 & ~w12341;
assign w12343 = w2558 & ~w11352;
assign w12344 = ~w11870 & w12343;
assign w12345 = w11870 & ~w12342;
assign w12346 = ~w12344 & ~w12345;
assign w12347 = ~w2285 & ~w12318;
assign w12348 = w12327 & w12347;
assign w12349 = ~w2285 & w12318;
assign w12350 = (w12349 & w12326) | (w12349 & w41064) | (w12326 & w41064);
assign w12351 = w12346 & ~w12350;
assign w12352 = ~w12348 & w12351;
assign w12353 = w12317 & w12352;
assign w12354 = (~w11869 & w11332) | (~w11869 & w44598) | (w11332 & w44598);
assign w12355 = ~w12246 & w12354;
assign w12356 = (w12355 & w11814) | (w12355 & w41065) | (w11814 & w41065);
assign w12357 = w3242 & w11869;
assign w12358 = ~w11815 & w41066;
assign w12359 = (~w12357 & w11814) | (~w12357 & w41067) | (w11814 & w41067);
assign w12360 = ~w12356 & w12359;
assign w12361 = ~w11343 & w11358;
assign w12362 = ~w2558 & w12337;
assign w12363 = w12362 & w52238;
assign w12364 = ~w2558 & ~w12337;
assign w12365 = (w12246 & w44599) | (w12246 & w44600) | (w44599 & w44600);
assign w12366 = ~w12363 & ~w12365;
assign w12367 = ~w2558 & w11352;
assign w12368 = ~w11870 & w12367;
assign w12369 = w11870 & ~w12366;
assign w12370 = ~w12368 & ~w12369;
assign w12371 = w2896 & w12361;
assign w12372 = ~w12360 & w12371;
assign w12373 = w2896 & ~w12361;
assign w12374 = w12360 & w12373;
assign w12375 = w12370 & ~w12374;
assign w12376 = ~w12372 & w12375;
assign w12377 = ~w2896 & ~w12361;
assign w12378 = ~w12360 & w12377;
assign w12379 = ~w2896 & w12361;
assign w12380 = w12360 & w12379;
assign w12381 = ~w12378 & ~w12380;
assign w12382 = ~w11232 & ~w11328;
assign w12383 = (~w11327 & ~w11286) | (~w11327 & w44601) | (~w11286 & w44601);
assign w12384 = ~w11578 & w12383;
assign w12385 = ~w11316 & w12383;
assign w12386 = ~w12384 & w52239;
assign w12387 = w12382 & ~w12386;
assign w12388 = ~w12382 & w12386;
assign w12389 = ~w12387 & ~w12388;
assign w12390 = w11231 & ~w11870;
assign w12391 = w11870 & ~w12389;
assign w12392 = ~w12390 & ~w12391;
assign w12393 = ~w3242 & ~w12392;
assign w12394 = w12381 & w12393;
assign w12395 = w12376 & ~w12394;
assign w12396 = w12353 & ~w12395;
assign w12397 = ~w12336 & ~w12396;
assign w12398 = ~w12396 & w47276;
assign w12399 = ~w12178 & w41069;
assign w12400 = (w12179 & w12178) | (w12179 & w41070) | (w12178 & w41070);
assign w12401 = ~w12399 & ~w12400;
assign w12402 = (w5330 & w12400) | (w5330 & w50312) | (w12400 & w50312);
assign w12403 = ~w5745 & ~w12196;
assign w12404 = ~w12199 & w12403;
assign w12405 = ~w5745 & w12196;
assign w12406 = w12199 & w12405;
assign w12407 = ~w12404 & ~w12406;
assign w12408 = ~w12402 & w12407;
assign w12409 = (~w12213 & ~w12159) | (~w12213 & w41071) | (~w12159 & w41071);
assign w12410 = w12195 & ~w12213;
assign w12411 = ~w12408 & w12410;
assign w12412 = ~w12409 & ~w12411;
assign w12413 = w12398 & w12412;
assign w12414 = w42 & ~w11879;
assign w12415 = ~w42 & ~w11886;
assign w12416 = w11852 & ~w11882;
assign w12417 = w11851 & ~w12416;
assign w12418 = w42 & ~w11883;
assign w12419 = ~w12417 & w12418;
assign w12420 = ~w12415 & ~w12419;
assign w12421 = ~w12414 & w12420;
assign w12422 = w11459 & ~w11713;
assign w12423 = ~w11869 & ~w12422;
assign w12424 = ~w11815 & w41072;
assign w12425 = w11712 & w11869;
assign w12426 = (~w12425 & w11814) | (~w12425 & w41073) | (w11814 & w41073);
assign w12427 = ~w11866 & w12423;
assign w12428 = w12426 & ~w12427;
assign w12429 = ~w11450 & w11760;
assign w12430 = w11745 & w12429;
assign w12431 = ~w12220 & w41074;
assign w12432 = ~w11450 & w11761;
assign w12433 = ~w11869 & ~w12432;
assign w12434 = ~w11450 & w12433;
assign w12435 = ~w12431 & w12434;
assign w12436 = ~w11866 & w12435;
assign w12437 = (~w493 & w11866) | (~w493 & w41075) | (w11866 & w41075);
assign w12438 = ~w12428 & w12437;
assign w12439 = ~w11866 & w41076;
assign w12440 = w12428 & w12439;
assign w12441 = ~w12438 & ~w12440;
assign w12442 = (~w11869 & ~w11709) | (~w11869 & w41077) | (~w11709 & w41077);
assign w12443 = w493 & w11865;
assign w12444 = w493 & w11869;
assign w12445 = (~w12444 & w11814) | (~w12444 & w44602) | (w11814 & w44602);
assign w12446 = ~w11866 & w12442;
assign w12447 = w12445 & ~w12446;
assign w12448 = ~w11207 & ~w11764;
assign w12449 = w400 & ~w12448;
assign w12450 = w12447 & w12449;
assign w12451 = w400 & w12448;
assign w12452 = ~w12447 & w12451;
assign w12453 = ~w12450 & ~w12452;
assign w12454 = w12441 & w12453;
assign w12455 = ~w11450 & w11752;
assign w12456 = w11491 & ~w12455;
assign w12457 = ~w12233 & w12456;
assign w12458 = w11753 & ~w12455;
assign w12459 = w12433 & ~w12458;
assign w12460 = ~w12431 & w12459;
assign w12461 = ~w11866 & w41078;
assign w12462 = ~w11444 & ~w11448;
assign w12463 = ~w11870 & w12462;
assign w12464 = ~w12461 & ~w12463;
assign w12465 = ~w12461 & w50517;
assign w12466 = ~w11866 & w41079;
assign w12467 = ~w12428 & w12466;
assign w12468 = (w493 & w11866) | (w493 & w41080) | (w11866 & w41080);
assign w12469 = w12428 & w12468;
assign w12470 = ~w12467 & ~w12469;
assign w12471 = ~w12465 & w12470;
assign w12472 = w12454 & ~w12471;
assign w12473 = ~w11207 & w11492;
assign w12474 = w11436 & w12473;
assign w12475 = ~w11344 & w12474;
assign w12476 = ~w11705 & w12474;
assign w12477 = w11583 & w12476;
assign w12478 = ~w12475 & ~w12477;
assign w12479 = ~w11207 & w11713;
assign w12480 = ~w11207 & ~w11760;
assign w12481 = w11762 & w12480;
assign w12482 = ~w12479 & ~w12481;
assign w12483 = ~w11746 & w41081;
assign w12484 = ~w11745 & w12483;
assign w12485 = w11183 & ~w11764;
assign w12486 = w12482 & w44603;
assign w12487 = w11194 & ~w11869;
assign w12488 = (w12487 & ~w12478) | (w12487 & w44604) | (~w12478 & w44604);
assign w12489 = ~w11866 & w12488;
assign w12490 = ~w11815 & w41082;
assign w12491 = w351 & w11869;
assign w12492 = (~w12491 & w11814) | (~w12491 & w41083) | (w11814 & w41083);
assign w12493 = ~w12489 & w12492;
assign w12494 = ~w11170 & w11188;
assign w12495 = ~w252 & ~w12494;
assign w12496 = (w12495 & w12489) | (w12495 & w41084) | (w12489 & w41084);
assign w12497 = ~w252 & w12494;
assign w12498 = ~w12489 & w41085;
assign w12499 = ~w12496 & ~w12498;
assign w12500 = ~w11170 & ~w11209;
assign w12501 = w11493 & w12500;
assign w12502 = ~w11160 & ~w11211;
assign w12503 = (~w12502 & w11769) | (~w12502 & w41086) | (w11769 & w41086);
assign w12504 = (w12501 & w12246) | (w12501 & w41087) | (w12246 & w41087);
assign w12505 = w12503 & ~w12504;
assign w12506 = w12501 & w12502;
assign w12507 = ~w12247 & w12506;
assign w12508 = ~w11769 & w41088;
assign w12509 = ~w12507 & ~w12508;
assign w12510 = ~w11159 & ~w11870;
assign w12511 = ~w12505 & w12509;
assign w12512 = w11870 & w12511;
assign w12513 = ~w12510 & ~w12512;
assign w12514 = (~w57 & w12512) | (~w57 & w41089) | (w12512 & w41089);
assign w12515 = w12499 & ~w12514;
assign w12516 = w12482 & w44605;
assign w12517 = w11183 & w11194;
assign w12518 = w12478 & w44606;
assign w12519 = (w12517 & ~w12478) | (w12517 & w44607) | (~w12478 & w44607);
assign w12520 = ~w12518 & ~w12519;
assign w12521 = w11177 & ~w11178;
assign w12522 = ~w11177 & w11178;
assign w12523 = ~w12521 & ~w12522;
assign w12524 = w11870 & w12520;
assign w12525 = ~w11870 & ~w12523;
assign w12526 = ~w12524 & ~w12525;
assign w12527 = (w351 & w12524) | (w351 & w41090) | (w12524 & w41090);
assign w12528 = ~w400 & ~w12448;
assign w12529 = ~w12447 & w12528;
assign w12530 = ~w400 & w12448;
assign w12531 = w12447 & w12530;
assign w12532 = ~w12529 & ~w12531;
assign w12533 = ~w12527 & w12532;
assign w12534 = ~w12512 & w41091;
assign w12535 = ~w11783 & ~w11784;
assign w12536 = ~w11782 & w12535;
assign w12537 = w11771 & w12536;
assign w12538 = (w11780 & ~w12537) | (w11780 & w41092) | (~w12537 & w41092);
assign w12539 = w11771 & w11787;
assign w12540 = w11870 & w12539;
assign w12541 = (~w80 & ~w12539) | (~w80 & w41093) | (~w12539 & w41093);
assign w12542 = ~w12538 & w12541;
assign w12543 = ~w12534 & ~w12542;
assign w12544 = w80 & ~w11869;
assign w12545 = (w11709 & w50518) | (w11709 & w50519) | (w50518 & w50519);
assign w12546 = ~w11788 & w12545;
assign w12547 = ~w80 & ~w11869;
assign w12548 = ~w11213 & w12547;
assign w12549 = (w12548 & ~w11709) | (w12548 & w50520) | (~w11709 & w50520);
assign w12550 = ~w11787 & ~w11866;
assign w12551 = w12549 & w12550;
assign w12552 = ~w12546 & ~w12551;
assign w12553 = w3 & w11147;
assign w12554 = ~w12552 & w12553;
assign w12555 = w3 & ~w11147;
assign w12556 = w12552 & w12555;
assign w12557 = ~w12554 & ~w12556;
assign w12558 = w12543 & w12557;
assign w12559 = ~w12524 & w41095;
assign w12560 = w252 & ~w12494;
assign w12561 = ~w12489 & w41096;
assign w12562 = w252 & w12494;
assign w12563 = (w12562 & w12489) | (w12562 & w41097) | (w12489 & w41097);
assign w12564 = ~w12561 & ~w12563;
assign w12565 = ~w12559 & w12564;
assign w12566 = w12515 & ~w12565;
assign w12567 = w12558 & ~w12566;
assign w12568 = w12515 & w12533;
assign w12569 = ~w12472 & w12568;
assign w12570 = w12567 & ~w12569;
assign w12571 = w11147 & ~w12552;
assign w12572 = ~w11147 & w12552;
assign w12573 = ~w12571 & ~w12572;
assign w12574 = ~w12538 & ~w12540;
assign w12575 = w80 & ~w12574;
assign w12576 = ~w3 & w12573;
assign w12577 = w12557 & w12575;
assign w12578 = ~w12576 & ~w12577;
assign w12579 = ~w11888 & w12578;
assign w12580 = ~w12570 & w12579;
assign w12581 = w12421 & ~w12580;
assign w12582 = (w12413 & w12580) | (w12413 & w47277) | (w12580 & w47277);
assign w12583 = ~w12217 & w12582;
assign w12584 = w3242 & w12392;
assign w12585 = w12381 & ~w12584;
assign w12586 = w12376 & ~w12585;
assign w12587 = w12353 & ~w12586;
assign w12588 = ~w12336 & ~w12587;
assign w12589 = ~w12587 & w47276;
assign w12590 = (~w612 & w12461) | (~w612 & w44608) | (w12461 & w44608);
assign w12591 = (~w754 & w12241) | (~w754 & w44609) | (w12241 & w44609);
assign w12592 = ~w12590 & ~w12591;
assign w12593 = w12454 & w12592;
assign w12594 = w12454 & w41098;
assign w12595 = ~w1541 & ~w12301;
assign w12596 = ~w12253 & w41099;
assign w12597 = (w12254 & w12253) | (w12254 & w41100) | (w12253 & w41100);
assign w12598 = ~w12596 & ~w12597;
assign w12599 = ~w1320 & ~w12598;
assign w12600 = ~w12595 & ~w12599;
assign w12601 = w12275 & ~w12600;
assign w12602 = ~w12229 & w50313;
assign w12603 = ~w12267 & w41101;
assign w12604 = (w12268 & w12267) | (w12268 & w41102) | (w12267 & w41102);
assign w12605 = ~w12603 & ~w12604;
assign w12606 = w1120 & ~w12605;
assign w12607 = ~w12602 & ~w12606;
assign w12608 = (w12243 & w12606) | (w12243 & w44610) | (w12606 & w44610);
assign w12609 = ~w12601 & ~w12608;
assign w12610 = w12594 & w12609;
assign w12611 = ~w12589 & w12610;
assign w12612 = w12558 & w12594;
assign w12613 = w12421 & w12612;
assign w12614 = w12611 & w12613;
assign w12615 = ~w12581 & ~w12614;
assign w12616 = ~w12583 & ~w12615;
assign w12617 = ~a[52] & ~a[53];
assign w12618 = ~a[54] & w12617;
assign w12619 = w11870 & w12618;
assign w12620 = ~w11870 & ~w12618;
assign w12621 = ~w12589 & w12609;
assign w12622 = ~w12580 & w41104;
assign w12623 = w12612 & w41104;
assign w12624 = a[55] & w12620;
assign w12625 = (~w12624 & w12583) | (~w12624 & w41105) | (w12583 & w41105);
assign w12626 = w11940 & ~w12619;
assign w12627 = (w12626 & w12583) | (w12626 & w41106) | (w12583 & w41106);
assign w12628 = w12625 & ~w12627;
assign w12629 = a[55] & ~w12619;
assign w12630 = w12629 & w50187;
assign w12631 = w12628 & ~w12630;
assign w12632 = w12398 & w12588;
assign w12633 = w12612 & w47278;
assign w12634 = ~w12632 & w12633;
assign w12635 = ~w12581 & ~w12634;
assign w12636 = (w12412 & w12075) | (w12412 & w12724) | (w12075 & w12724);
assign w12637 = ~w12635 & ~w12636;
assign w12638 = ~w12398 & w12613;
assign w12639 = w12621 & w12638;
assign w12640 = ~w12581 & ~w12639;
assign w12641 = a[56] & ~w11940;
assign w12642 = ~w11941 & ~w12641;
assign w12643 = ~w11138 & w12642;
assign w12644 = w12640 & w12643;
assign w12645 = ~w12637 & w12644;
assign w12646 = ~a[56] & ~w11870;
assign w12647 = a[56] & w11870;
assign w12648 = ~w12646 & ~w12647;
assign w12649 = ~w11138 & ~w12648;
assign w12650 = ~w12580 & w41107;
assign w12651 = w12612 & w41107;
assign w12652 = w12621 & w12651;
assign w12653 = ~w12650 & ~w12652;
assign w12654 = w11888 & w12649;
assign w12655 = (~w12654 & w12583) | (~w12654 & w41108) | (w12583 & w41108);
assign w12656 = ~w12645 & w12655;
assign w12657 = ~w12648 & w50187;
assign w12658 = w12640 & w12642;
assign w12659 = ~w12637 & w12658;
assign w12660 = w11138 & ~w12659;
assign w12661 = ~w12657 & w12660;
assign w12662 = w12660 & w47279;
assign w12663 = ~w10419 & w12656;
assign w12664 = ~w12631 & w12663;
assign w12665 = ~w12662 & ~w12664;
assign w12666 = ~w12637 & w12640;
assign w12667 = w10419 & ~w11959;
assign w12668 = ~w10419 & w11959;
assign w12669 = ~w12667 & ~w12668;
assign w12670 = ~w12637 & w44611;
assign w12671 = w9781 & ~w11972;
assign w12672 = ~w12670 & w12671;
assign w12673 = w9781 & w11972;
assign w12674 = w12670 & w12673;
assign w12675 = ~w12672 & ~w12674;
assign w12676 = (w10419 & ~w12660) | (w10419 & w47280) | (~w12660 & w47280);
assign w12677 = ~w12631 & w12656;
assign w12678 = w12676 & ~w12677;
assign w12679 = a[56] & a[57];
assign w12680 = w11951 & ~w12679;
assign w12681 = w11956 & ~w11957;
assign w12682 = ~w11942 & ~w11948;
assign w12683 = w12681 & ~w12682;
assign w12684 = ~w11138 & ~w12680;
assign w12685 = ~w11941 & ~w12647;
assign w12686 = w12684 & ~w12685;
assign w12687 = w11942 & ~w11945;
assign w12688 = ~w12686 & ~w12687;
assign w12689 = (w12683 & w12583) | (w12683 & w44612) | (w12583 & w44612);
assign w12690 = w12688 & ~w12689;
assign w12691 = w12616 & ~w12680;
assign w12692 = w12690 & ~w12691;
assign w12693 = (w12675 & w12664) | (w12675 & w47281) | (w12664 & w47281);
assign w12694 = w12675 & ~w12692;
assign w12695 = ~w12678 & w12694;
assign w12696 = ~w12693 & ~w12695;
assign w12697 = w11972 & ~w12670;
assign w12698 = ~w11972 & w12670;
assign w12699 = ~w12697 & ~w12698;
assign w12700 = ~w9781 & ~w12699;
assign w12701 = ~w12028 & w12039;
assign w12702 = ~w12009 & ~w12031;
assign w12703 = w12701 & ~w12702;
assign w12704 = ~w12701 & w12702;
assign w12705 = ~w12703 & ~w12704;
assign w12706 = ~w12583 & w41109;
assign w12707 = (w12705 & w12583) | (w12705 & w41110) | (w12583 & w41110);
assign w12708 = ~w12706 & ~w12707;
assign w12709 = ~w8666 & w12708;
assign w12710 = (~w12028 & ~w12030) | (~w12028 & w50521) | (~w12030 & w50521);
assign w12711 = (w8666 & w12049) | (w8666 & w50522) | (w12049 & w50522);
assign w12712 = ~w12049 & w50523;
assign w12713 = ~w12711 & ~w12712;
assign w12714 = w11909 & w12713;
assign w12715 = w12640 & w12714;
assign w12716 = ~w12637 & w12715;
assign w12717 = ~w12580 & w41111;
assign w12718 = w12612 & w41111;
assign w12719 = w12621 & w12718;
assign w12720 = ~w11909 & ~w12713;
assign w12721 = (~w12720 & w12583) | (~w12720 & w41112) | (w12583 & w41112);
assign w12722 = ~w12716 & w12721;
assign w12723 = w12075 & w12412;
assign w12724 = ~w12216 & w12412;
assign w12725 = w12713 & ~w12724;
assign w12726 = ~w12723 & w12725;
assign w12727 = ~w12635 & w12726;
assign w12728 = ~w12616 & w12727;
assign w12729 = (~w7924 & w12616) | (~w7924 & w41113) | (w12616 & w41113);
assign w12730 = w12722 & w12729;
assign w12731 = ~w12709 & ~w12730;
assign w12732 = w8666 & ~w12708;
assign w12733 = ~w11974 & ~w12007;
assign w12734 = w9781 & ~w12733;
assign w12735 = ~w9781 & w12733;
assign w12736 = ~w12734 & ~w12735;
assign w12737 = (~w12736 & w12583) | (~w12736 & w41114) | (w12583 & w41114);
assign w12738 = w9195 & ~w12030;
assign w12739 = ~w12737 & w12738;
assign w12740 = w9195 & w12030;
assign w12741 = w12737 & w12740;
assign w12742 = ~w12739 & ~w12741;
assign w12743 = ~w12732 & ~w12742;
assign w12744 = w12731 & w50524;
assign w12745 = w12696 & w12744;
assign w12746 = (~w41115 & w50314) | (~w41115 & w50315) | (w50314 & w50315);
assign w12747 = w7924 & ~w12034;
assign w12748 = (w12747 & w12049) | (w12747 & w41116) | (w12049 & w41116);
assign w12749 = (~w41116 & w50316) | (~w41116 & w50317) | (w50316 & w50317);
assign w12750 = ~w12746 & ~w12749;
assign w12751 = w7315 & ~w12750;
assign w12752 = ~w7315 & w12750;
assign w12753 = ~w12751 & ~w12752;
assign w12754 = ~w7315 & w11929;
assign w12755 = w11933 & ~w12750;
assign w12756 = w12750 & w12754;
assign w12757 = ~w12755 & ~w12756;
assign w12758 = w12640 & ~w12757;
assign w12759 = (~w6769 & ~w12758) | (~w6769 & w50318) | (~w12758 & w50318);
assign w12760 = ~w11929 & w50188;
assign w12761 = w12759 & ~w12760;
assign w12762 = (w12042 & w12009) | (w12042 & w50525) | (w12009 & w50525);
assign w12763 = w11938 & ~w12762;
assign w12764 = ~w6769 & w12763;
assign w12765 = w6769 & ~w12763;
assign w12766 = ~w12764 & ~w12765;
assign w12767 = w12640 & ~w12766;
assign w12768 = (~w11902 & ~w12767) | (~w11902 & w50319) | (~w12767 & w50319);
assign w12769 = w12216 & w12609;
assign w12770 = ~w12589 & w12769;
assign w12771 = ~w12075 & w12770;
assign w12772 = ~w12413 & w12621;
assign w12773 = ~w12771 & ~w12772;
assign w12774 = (w11902 & w12580) | (w11902 & w44613) | (w12580 & w44613);
assign w12775 = ~w12766 & w12774;
assign w12776 = (w12613 & w12771) | (w12613 & w41118) | (w12771 & w41118);
assign w12777 = w12775 & ~w12776;
assign w12778 = (w6264 & w12776) | (w6264 & w44614) | (w12776 & w44614);
assign w12779 = ~w12768 & w12778;
assign w12780 = ~w12761 & ~w12779;
assign w12781 = w12758 & w50320;
assign w12782 = w6769 & ~w11929;
assign w12783 = w12782 & w50188;
assign w12784 = ~w12781 & ~w12783;
assign w12785 = ~w12746 & ~w12748;
assign w12786 = w11922 & w50189;
assign w12787 = ~w12746 & w12749;
assign w12788 = ~w12639 & w50321;
assign w12789 = ~w12637 & w12788;
assign w12790 = ~w7315 & ~w12789;
assign w12791 = ~w12786 & w12790;
assign w12792 = w12784 & ~w12791;
assign w12793 = ~w12768 & ~w12777;
assign w12794 = (~w6264 & w12768) | (~w6264 & w44615) | (w12768 & w44615);
assign w12795 = w12072 & w12763;
assign w12796 = w12046 & ~w12055;
assign w12797 = ~w12795 & w12796;
assign w12798 = (~w41120 & w47282) | (~w41120 & w47283) | (w47282 & w47283);
assign w12799 = (w41120 & w47284) | (w41120 & w47285) | (w47284 & w47285);
assign w12800 = ~w12798 & ~w12799;
assign w12801 = w5745 & ~w12800;
assign w12802 = ~w12794 & ~w12801;
assign w12803 = w12780 & ~w12792;
assign w12804 = w12802 & ~w12803;
assign w12805 = ~w12786 & ~w12789;
assign w12806 = w7315 & ~w12805;
assign w12807 = w12780 & ~w12806;
assign w12808 = w12804 & ~w12807;
assign w12809 = (w7924 & w12716) | (w7924 & w48746) | (w12716 & w48746);
assign w12810 = w12030 & ~w12737;
assign w12811 = (w12583 & w50526) | (w12583 & w50527) | (w50526 & w50527);
assign w12812 = ~w12810 & ~w12811;
assign w12813 = ~w9195 & ~w12812;
assign w12814 = (~w12809 & w12730) | (~w12809 & w48747) | (w12730 & w48747);
assign w12815 = ~w12732 & ~w12809;
assign w12816 = ~w12813 & w12815;
assign w12817 = ~w12814 & ~w12816;
assign w12818 = ~w12203 & w12407;
assign w12819 = w12075 & ~w12818;
assign w12820 = ~w12075 & w12818;
assign w12821 = ~w12819 & ~w12820;
assign w12822 = (w12202 & w12637) | (w12202 & w44616) | (w12637 & w44616);
assign w12823 = ~w12637 & w44617;
assign w12824 = ~w12822 & ~w12823;
assign w12825 = (w5330 & w12823) | (w5330 & w50528) | (w12823 & w50528);
assign w12826 = ~w5745 & w12800;
assign w12827 = ~w12825 & ~w12826;
assign w12828 = ~w12817 & w12827;
assign w12829 = ~w12808 & w12828;
assign w12830 = ~w12745 & w12829;
assign w12831 = ~w12073 & w12408;
assign w12832 = ~w12069 & w12831;
assign w12833 = w12046 & w12832;
assign w12834 = (w12184 & w12202) | (w12184 & w50529) | (w12202 & w50529);
assign w12835 = ~w12402 & ~w12834;
assign w12836 = w12193 & ~w12835;
assign w12837 = (w12833 & w50530) | (w12833 & w50531) | (w50530 & w50531);
assign w12838 = w3646 & w52240;
assign w12839 = ~w12837 & ~w12838;
assign w12840 = (w12212 & w12583) | (w12212 & w41122) | (w12583 & w41122);
assign w12841 = ~w12839 & w12840;
assign w12842 = w12840 & w44618;
assign w12843 = ~w3242 & ~w12212;
assign w12844 = (w12843 & ~w12666) | (w12843 & w44619) | (~w12666 & w44619);
assign w12845 = ~w12842 & ~w12844;
assign w12846 = ~w12584 & ~w12724;
assign w12847 = ~w12723 & w12846;
assign w12848 = (~w12393 & w12723) | (~w12393 & w44620) | (w12723 & w44620);
assign w12849 = ~w3242 & ~w12636;
assign w12850 = ~w12848 & ~w12849;
assign w12851 = (w12392 & w12847) | (w12392 & w50532) | (w12847 & w50532);
assign w12852 = (w12584 & ~w12635) | (w12584 & w44621) | (~w12635 & w44621);
assign w12853 = ~w12851 & ~w12852;
assign w12854 = w12666 & w12850;
assign w12855 = w12853 & ~w12854;
assign w12856 = w12853 & w50322;
assign w12857 = w12845 & ~w12856;
assign w12858 = ~w12113 & w12152;
assign w12859 = w12408 & ~w12858;
assign w12860 = ~w12073 & w12859;
assign w12861 = ~w12069 & w12860;
assign w12862 = ~w12836 & ~w12858;
assign w12863 = w12046 & w12861;
assign w12864 = ~w12862 & ~w12863;
assign w12865 = (w4056 & w12863) | (w4056 & w41123) | (w12863 & w41123);
assign w12866 = ~w12863 & w41124;
assign w12867 = ~w12865 & ~w12866;
assign w12868 = (w12157 & w12616) | (w12157 & w41125) | (w12616 & w41125);
assign w12869 = ~w12157 & ~w12867;
assign w12870 = w12666 & w12869;
assign w12871 = ~w12868 & ~w12870;
assign w12872 = ~w12870 & w47287;
assign w12873 = (~w12212 & ~w12666) | (~w12212 & w44622) | (~w12666 & w44622);
assign w12874 = (w3242 & ~w12840) | (w3242 & w47288) | (~w12840 & w47288);
assign w12875 = ~w12873 & w12874;
assign w12876 = ~w12872 & ~w12875;
assign w12877 = ~w2896 & ~w12855;
assign w12878 = w12360 & ~w12361;
assign w12879 = ~w12360 & w12361;
assign w12880 = ~w12878 & ~w12879;
assign w12881 = ~w2896 & ~w12880;
assign w12882 = ~w12848 & ~w12881;
assign w12883 = w2896 & ~w12880;
assign w12884 = w12848 & ~w12883;
assign w12885 = ~w12616 & ~w12884;
assign w12886 = ~w12381 & w12848;
assign w12887 = ~w12583 & w41126;
assign w12888 = w2896 & w12880;
assign w12889 = ~w12848 & w12888;
assign w12890 = ~w12882 & w12885;
assign w12891 = (w2558 & w12890) | (w2558 & w44624) | (w12890 & w44624);
assign w12892 = ~w12877 & ~w12891;
assign w12893 = w12857 & ~w12876;
assign w12894 = w12892 & ~w12893;
assign w12895 = (w12827 & w12803) | (w12827 & w47289) | (w12803 & w47289);
assign w12896 = w12184 & ~w12402;
assign w12897 = w12407 & ~w12896;
assign w12898 = (w12897 & w12075) | (w12897 & w48748) | (w12075 & w48748);
assign w12899 = w12640 & ~w12898;
assign w12900 = w5330 & w11888;
assign w12901 = w12897 & ~w12900;
assign w12902 = (w12901 & w12075) | (w12901 & w48749) | (w12075 & w48749);
assign w12903 = ~w12401 & ~w12902;
assign w12904 = ~w12580 & w41127;
assign w12905 = w12612 & w41127;
assign w12906 = w12621 & w12905;
assign w12907 = ~w12904 & ~w12906;
assign w12908 = ~w12583 & ~w12907;
assign w12909 = ~w12903 & ~w12908;
assign w12910 = ~w12637 & w12899;
assign w12911 = w12909 & ~w12910;
assign w12912 = (w12407 & w12075) | (w12407 & w48750) | (w12075 & w48750);
assign w12913 = w12896 & ~w12912;
assign w12914 = ~w4838 & ~w12913;
assign w12915 = ~w4838 & ~w12401;
assign w12916 = ~w12583 & w41128;
assign w12917 = ~w12914 & ~w12916;
assign w12918 = ~w12911 & ~w12917;
assign w12919 = (~w12835 & ~w12832) | (~w12835 & w41129) | (~w12832 & w41129);
assign w12920 = w12090 & ~w12919;
assign w12921 = w12640 & ~w12920;
assign w12922 = ~w12637 & w12921;
assign w12923 = ~w11866 & ~w12081;
assign w12924 = w11315 & ~w12923;
assign w12925 = ~w11315 & w12923;
assign w12926 = ~w12924 & ~w12925;
assign w12927 = ~w12580 & w41130;
assign w12928 = w12612 & w41130;
assign w12929 = w12621 & w12928;
assign w12930 = ~w12927 & ~w12929;
assign w12931 = ~w12583 & ~w12930;
assign w12932 = w12919 & w12926;
assign w12933 = w4430 & w12192;
assign w12934 = ~w12932 & w12933;
assign w12935 = ~w12931 & w12934;
assign w12936 = ~w12090 & w12919;
assign w12937 = (~w12613 & w12580) | (~w12613 & ~w12421) | (w12580 & ~w12421);
assign w12938 = ~w12570 & w12578;
assign w12939 = w11888 & ~w12938;
assign w12940 = w12937 & ~w12939;
assign w12941 = ~w12773 & ~w12940;
assign w12942 = (~w12192 & w12580) | (~w12192 & w41131) | (w12580 & w41131);
assign w12943 = w12919 & w12942;
assign w12944 = w4430 & w12936;
assign w12945 = w12942 & w48751;
assign w12946 = (~w12944 & w12941) | (~w12944 & w41132) | (w12941 & w41132);
assign w12947 = ~w12922 & w12935;
assign w12948 = w12946 & ~w12947;
assign w12949 = ~w12918 & w12948;
assign w12950 = ~w12823 & w50533;
assign w12951 = ~w12583 & w41133;
assign w12952 = w12913 & ~w12951;
assign w12953 = ~w12911 & ~w12952;
assign w12954 = (w4838 & w12911) | (w4838 & w41134) | (w12911 & w41134);
assign w12955 = ~w12950 & ~w12954;
assign w12956 = w12949 & ~w12955;
assign w12957 = (w12580 & w47290) | (w12580 & w47291) | (w47290 & w47291);
assign w12958 = w12152 & ~w12957;
assign w12959 = ~w12581 & w12864;
assign w12960 = w12773 & w12959;
assign w12961 = (w12192 & w12919) | (w12192 & w50534) | (w12919 & w50534);
assign w12962 = (~w12961 & w12960) | (~w12961 & w41135) | (w12960 & w41135);
assign w12963 = (~w4430 & w44625) | (~w4430 & ~w12937) | (w44625 & ~w12937);
assign w12964 = ~w12771 & w41136;
assign w12965 = ~w12863 & w47292;
assign w12966 = (w12965 & w12964) | (w12965 & w44626) | (w12964 & w44626);
assign w12967 = ~w11866 & w12100;
assign w12968 = ~w12103 & ~w12967;
assign w12969 = w12103 & w12967;
assign w12970 = ~w12968 & ~w12969;
assign w12971 = (w12970 & w12637) | (w12970 & w44627) | (w12637 & w44627);
assign w12972 = ~w12966 & ~w12971;
assign w12973 = ~w12962 & w12972;
assign w12974 = (~w4056 & ~w12972) | (~w4056 & w47293) | (~w12972 & w47293);
assign w12975 = w12192 & ~w12932;
assign w12976 = ~w12931 & w12975;
assign w12977 = ~w12922 & w12976;
assign w12978 = (w12943 & w12773) | (w12943 & w41137) | (w12773 & w41137);
assign w12979 = ~w12936 & ~w12978;
assign w12980 = ~w12977 & w12979;
assign w12981 = ~w12977 & w41138;
assign w12982 = ~w12974 & ~w12981;
assign w12983 = ~w12956 & w12982;
assign w12984 = ~w12895 & w12983;
assign w12985 = w12894 & w12984;
assign w12986 = ~w12830 & w12985;
assign w12987 = ~w12949 & ~w12981;
assign w12988 = ~w12949 & w12982;
assign w12989 = (~w3646 & w12870) | (~w3646 & w47294) | (w12870 & w47294);
assign w12990 = w4056 & ~w12962;
assign w12991 = w12972 & w12990;
assign w12992 = ~w12989 & ~w12991;
assign w12993 = w12857 & w12992;
assign w12994 = ~w12988 & w12993;
assign w12995 = w12894 & ~w12994;
assign w12996 = (~w12995 & w12830) | (~w12995 & w47295) | (w12830 & w47295);
assign w12997 = ~w12230 & w50190;
assign w12998 = ~w12302 & w50323;
assign w12999 = (w12335 & w12395) | (w12335 & w50324) | (w12395 & w50324);
assign w13000 = w12412 & w12999;
assign w13001 = ~w12587 & w44628;
assign w13002 = (w12998 & w12215) | (w12998 & w41140) | (w12215 & w41140);
assign w13003 = (~w13001 & ~w13000) | (~w13001 & w41141) | (~w13000 & w41141);
assign w13004 = w12412 & w50325;
assign w13005 = w12075 & w13004;
assign w13006 = w12259 & ~w12600;
assign w13007 = ~w12606 & ~w13006;
assign w13008 = ~w13005 & w41142;
assign w13009 = w12273 & ~w13008;
assign w13010 = ~w945 & w12230;
assign w13011 = ~w12639 & w50326;
assign w13012 = ~w12637 & w13011;
assign w13013 = w13009 & ~w13012;
assign w13014 = ~w12997 & w13013;
assign w13015 = ~w12230 & w50191;
assign w13016 = ~w12639 & w50327;
assign w13017 = ~w12637 & w13016;
assign w13018 = ~w13009 & ~w13017;
assign w13019 = ~w13015 & w13018;
assign w13020 = ~w13014 & ~w13019;
assign w13021 = ~w754 & ~w13020;
assign w13022 = ~w12242 & ~w12591;
assign w13023 = w12607 & ~w13006;
assign w13024 = ~w13005 & w41144;
assign w13025 = ~w12273 & w12607;
assign w13026 = ~w12231 & ~w13025;
assign w13027 = ~w13024 & w13026;
assign w13028 = (w754 & w12637) | (w754 & w44629) | (w12637 & w44629);
assign w13029 = w12666 & ~w13027;
assign w13030 = (w13022 & w13029) | (w13022 & w44630) | (w13029 & w44630);
assign w13031 = ~w13029 & w44631;
assign w13032 = ~w13030 & ~w13031;
assign w13033 = ~w612 & ~w13032;
assign w13034 = ~w13021 & ~w13033;
assign w13035 = ~w13005 & w41145;
assign w13036 = w1120 & ~w13035;
assign w13037 = ~w1120 & ~w13006;
assign w13038 = ~w13005 & w41146;
assign w13039 = (~w13038 & w12583) | (~w13038 & w44632) | (w12583 & w44632);
assign w13040 = ~w13036 & ~w13038;
assign w13041 = (~w12605 & ~w13039) | (~w12605 & w41147) | (~w13039 & w41147);
assign w13042 = ~w12637 & w44633;
assign w13043 = w13040 & w13042;
assign w13044 = ~w13041 & ~w13043;
assign w13045 = ~w945 & w13044;
assign w13046 = w754 & w13020;
assign w13047 = ~w13045 & ~w13046;
assign w13048 = w945 & w12605;
assign w13049 = ~w12637 & w44634;
assign w13050 = w13040 & w13049;
assign w13051 = w945 & ~w12605;
assign w13052 = (w13051 & ~w13039) | (w13051 & w41148) | (~w13039 & w41148);
assign w13053 = ~w13050 & ~w13052;
assign w13054 = (~w12595 & w12587) | (~w12595 & w44635) | (w12587 & w44635);
assign w13055 = (w13054 & ~w12724) | (w13054 & w41149) | (~w12724 & w41149);
assign w13056 = w12075 & w13000;
assign w13057 = ~w12303 & ~w12595;
assign w13058 = (~w13057 & w13056) | (~w13057 & w44636) | (w13056 & w44636);
assign w13059 = w12259 & ~w12599;
assign w13060 = w13058 & ~w13059;
assign w13061 = ~w13058 & w13059;
assign w13062 = ~w13060 & ~w13061;
assign w13063 = w1120 & w52241;
assign w13064 = w12666 & w13062;
assign w13065 = w13063 & ~w13064;
assign w13066 = w13053 & ~w13065;
assign w13067 = ~w12302 & w13055;
assign w13068 = (w12412 & w12075) | (w12412 & w44638) | (w12075 & w44638);
assign w13069 = w13067 & ~w13068;
assign w13070 = ~w12302 & ~w12595;
assign w13071 = ~w12288 & ~w13070;
assign w13072 = w13000 & w13071;
assign w13073 = ~w12217 & w13072;
assign w13074 = ~w12288 & w12397;
assign w13075 = w13070 & ~w13074;
assign w13076 = w12588 & w13071;
assign w13077 = ~w13075 & ~w13076;
assign w13078 = ~w13073 & w13077;
assign w13079 = ~w13069 & w13078;
assign w13080 = (w12301 & w12637) | (w12301 & w44639) | (w12637 & w44639);
assign w13081 = w12666 & w13079;
assign w13082 = ~w13080 & ~w13081;
assign w13083 = (w1320 & w13081) | (w1320 & w44640) | (w13081 & w44640);
assign w13084 = (~w12598 & w12637) | (~w12598 & w44641) | (w12637 & w44641);
assign w13085 = ~w1120 & ~w13084;
assign w13086 = w12666 & ~w13062;
assign w13087 = w13085 & ~w13086;
assign w13088 = ~w13083 & ~w13087;
assign w13089 = w13066 & ~w13088;
assign w13090 = w13047 & ~w13089;
assign w13091 = w13034 & ~w13090;
assign w13092 = ~w12601 & w44642;
assign w13093 = w12770 & w41150;
assign w13094 = ~w12589 & w13092;
assign w13095 = ~w12413 & w13094;
assign w13096 = ~w612 & ~w13095;
assign w13097 = ~w13093 & w13096;
assign w13098 = w612 & ~w12591;
assign w13099 = w12770 & w41151;
assign w13100 = ~w12601 & w44643;
assign w13101 = ~w12589 & w13100;
assign w13102 = ~w12413 & w13101;
assign w13103 = (~w13102 & ~w41151) | (~w13102 & w47296) | (~w41151 & w47296);
assign w13104 = w12464 & ~w13102;
assign w13105 = ~w13099 & w13104;
assign w13106 = ~w13097 & w13105;
assign w13107 = (w493 & ~w13106) | (w493 & w50535) | (~w13106 & w50535);
assign w13108 = (~w12464 & ~w41152) | (~w12464 & w47297) | (~w41152 & w47297);
assign w13109 = w13107 & ~w13108;
assign w13110 = ~w400 & w13109;
assign w13111 = (w400 & ~w13107) | (w400 & w47298) | (~w13107 & w47298);
assign w13112 = ~w12590 & w13095;
assign w13113 = w12770 & w41153;
assign w13114 = ~w13112 & ~w13113;
assign w13115 = ~w13113 & w50328;
assign w13116 = w12428 & ~w12436;
assign w13117 = ~w12428 & w12436;
assign w13118 = ~w13116 & ~w13117;
assign w13119 = (w13118 & w12637) | (w13118 & w44644) | (w12637 & w44644);
assign w13120 = ~w13115 & ~w13119;
assign w13121 = w12441 & w12470;
assign w13122 = w12666 & w13121;
assign w13123 = w13120 & ~w13122;
assign w13124 = ~w13113 & w50329;
assign w13125 = ~w12583 & w44646;
assign w13126 = w13124 & ~w13125;
assign w13127 = ~w12470 & w12666;
assign w13128 = w13126 & ~w13127;
assign w13129 = ~w13123 & ~w13128;
assign w13130 = ~w13111 & ~w13129;
assign w13131 = ~w13110 & ~w13130;
assign w13132 = w12453 & w12532;
assign w13133 = ~w12637 & w44647;
assign w13134 = w12447 & ~w12448;
assign w13135 = ~w12447 & w12448;
assign w13136 = ~w13134 & ~w13135;
assign w13137 = (w400 & w12583) | (w400 & w41154) | (w12583 & w41154);
assign w13138 = w13136 & ~w13137;
assign w13139 = ~w13113 & w50330;
assign w13140 = w12441 & ~w13139;
assign w13141 = (~w13136 & w12637) | (~w13136 & w44648) | (w12637 & w44648);
assign w13142 = ~w13133 & ~w13141;
assign w13143 = ~w13140 & ~w13142;
assign w13144 = ~w13133 & ~w13138;
assign w13145 = w13140 & w13144;
assign w13146 = ~w13145 & w44649;
assign w13147 = w612 & w13032;
assign w13148 = ~w13146 & ~w13147;
assign w13149 = w13131 & w13148;
assign w13150 = ~w13091 & w13149;
assign w13151 = w11879 & ~w12419;
assign w13152 = ~w12414 & ~w13151;
assign w13153 = (w12612 & w12771) | (w12612 & w50536) | (w12771 & w50536);
assign w13154 = w12938 & ~w13153;
assign w13155 = w11879 & w12415;
assign w13156 = ~w13152 & ~w13154;
assign w13157 = ~w12414 & ~w13155;
assign w13158 = w13154 & w13157;
assign w13159 = ~w13156 & ~w13158;
assign w13160 = w12770 & w41155;
assign w13161 = ~w12413 & w12611;
assign w13162 = ~w12472 & w12533;
assign w13163 = (w12565 & w12472) | (w12565 & w50537) | (w12472 & w50537);
assign w13164 = w12499 & ~w13163;
assign w13165 = ~w12514 & w13164;
assign w13166 = ~w13161 & w13165;
assign w13167 = (w12543 & w13160) | (w12543 & w48752) | (w13160 & w48752);
assign w13168 = (~w12575 & w44650) | (~w12575 & w52242) | (w44650 & w52242);
assign w13169 = (w3 & w12583) | (w3 & w44651) | (w12583 & w44651);
assign w13170 = ~w13168 & w13169;
assign w13171 = ~w3 & ~w12575;
assign w13172 = (w13171 & w12583) | (w13171 & w41156) | (w12583 & w41156);
assign w13173 = ~w13167 & w13172;
assign w13174 = w12573 & ~w13173;
assign w13175 = ~w13170 & w13174;
assign w13176 = ~w3 & ~w12573;
assign w13177 = w12640 & w13176;
assign w13178 = ~w12637 & w13177;
assign w13179 = ~w12557 & ~w12581;
assign w13180 = w42 & ~w13179;
assign w13181 = ~w13168 & w13180;
assign w13182 = w42 & ~w13178;
assign w13183 = w13168 & w13182;
assign w13184 = ~w13181 & ~w13183;
assign w13185 = (~w13159 & w13184) | (~w13159 & w48753) | (w13184 & w48753);
assign w13186 = (~w12534 & w13160) | (~w12534 & w50538) | (w13160 & w50538);
assign w13187 = (w12542 & w12583) | (w12542 & w41157) | (w12583 & w41157);
assign w13188 = ~w12575 & ~w13187;
assign w13189 = w13186 & ~w13188;
assign w13190 = (~w12575 & w44652) | (~w12575 & w52242) | (w44652 & w52242);
assign w13191 = w12666 & ~w13190;
assign w13192 = w80 & w12640;
assign w13193 = ~w12637 & w13192;
assign w13194 = w12574 & ~w13193;
assign w13195 = ~w13188 & w44653;
assign w13196 = (~w3 & w13193) | (~w3 & w44654) | (w13193 & w44654);
assign w13197 = ~w13191 & w13196;
assign w13198 = ~w13195 & ~w13197;
assign w13199 = ~w42 & w12573;
assign w13200 = ~w13173 & w13199;
assign w13201 = ~w13170 & w13200;
assign w13202 = ~w12639 & w50331;
assign w13203 = ~w12637 & w50539;
assign w13204 = ~w13168 & w13203;
assign w13205 = ~w12637 & w50540;
assign w13206 = w13168 & w13205;
assign w13207 = ~w13204 & ~w13206;
assign w13208 = ~w13201 & w13207;
assign w13209 = w13198 & w13208;
assign w13210 = w13185 & ~w13209;
assign w13211 = ~w13161 & w13164;
assign w13212 = ~w13160 & w50541;
assign w13213 = (w57 & w13160) | (w57 & w50542) | (w13160 & w50542);
assign w13214 = ~w13212 & ~w13213;
assign w13215 = w12513 & w12666;
assign w13216 = ~w13214 & w13215;
assign w13217 = (~w12513 & w13214) | (~w12513 & w44655) | (w13214 & w44655);
assign w13218 = ~w13216 & ~w13217;
assign w13219 = w80 & ~w13218;
assign w13220 = w12471 & w12532;
assign w13221 = (w12075 & w50332) | (w12075 & w50333) | (w50332 & w50333);
assign w13222 = w12593 & w12609;
assign w13223 = ~w12632 & w13222;
assign w13224 = ~w12472 & w12532;
assign w13225 = ~w13223 & w13224;
assign w13226 = (~w13225 & ~w13114) | (~w13225 & w44656) | (~w13114 & w44656);
assign w13227 = ~w12559 & w52243;
assign w13228 = w12526 & ~w12666;
assign w13229 = ~w13226 & ~w13227;
assign w13230 = ~w13228 & ~w13229;
assign w13231 = ~w12527 & ~w12559;
assign w13232 = ~w12637 & w44657;
assign w13233 = w13226 & w13232;
assign w13234 = (~w252 & ~w13226) | (~w252 & w50543) | (~w13226 & w50543);
assign w13235 = w13230 & w13234;
assign w13236 = w12493 & ~w12494;
assign w13237 = ~w12493 & w12494;
assign w13238 = ~w13236 & ~w13237;
assign w13239 = (~w13238 & w12637) | (~w13238 & w44658) | (w12637 & w44658);
assign w13240 = w12499 & w12564;
assign w13241 = (w13240 & ~w41159) | (w13240 & w47299) | (~w41159 & w47299);
assign w13242 = ~w13239 & ~w13241;
assign w13243 = ~w13025 & w13162;
assign w13244 = w12243 & w13243;
assign w13245 = ~w12593 & w13162;
assign w13246 = ~w12559 & ~w13245;
assign w13247 = (w13246 & w13024) | (w13246 & w50334) | (w13024 & w50334);
assign w13248 = (~w13240 & ~w41159) | (~w13240 & w47300) | (~w41159 & w47300);
assign w13249 = ~w13239 & ~w13248;
assign w13250 = ~w57 & w13247;
assign w13251 = w13242 & w13250;
assign w13252 = ~w57 & ~w13247;
assign w13253 = w13249 & w13252;
assign w13254 = ~w13251 & ~w13253;
assign w13255 = ~w13235 & w13254;
assign w13256 = ~w13219 & w13255;
assign w13257 = ~w13210 & w13256;
assign w13258 = w12316 & ~w12334;
assign w13259 = w12352 & ~w12586;
assign w13260 = ~w12724 & w13259;
assign w13261 = ~w12395 & w13259;
assign w13262 = ~w12331 & ~w13261;
assign w13263 = (w13262 & w12723) | (w13262 & w50335) | (w12723 & w50335);
assign w13264 = ~w12616 & w13263;
assign w13265 = (w13258 & w13264) | (w13258 & w41161) | (w13264 & w41161);
assign w13266 = ~w13264 & w41162;
assign w13267 = ~w13265 & ~w13266;
assign w13268 = w1738 & ~w13267;
assign w13269 = w12335 & ~w13261;
assign w13270 = (w13269 & w12723) | (w13269 & w44659) | (w12723 & w44659);
assign w13271 = w12316 & ~w13270;
assign w13272 = (w1738 & w12637) | (w1738 & w44660) | (w12637 & w44660);
assign w13273 = w12666 & w13271;
assign w13274 = ~w12288 & ~w12305;
assign w13275 = w1541 & ~w13274;
assign w13276 = (w13275 & w13273) | (w13275 & w44661) | (w13273 & w44661);
assign w13277 = w1541 & w13274;
assign w13278 = ~w13273 & w44662;
assign w13279 = ~w13276 & ~w13278;
assign w13280 = ~w13268 & w13279;
assign w13281 = w12346 & ~w12586;
assign w13282 = ~w12724 & w13281;
assign w13283 = ~w12395 & w13281;
assign w13284 = w2285 & ~w12330;
assign w13285 = ~w13283 & w13284;
assign w13286 = (w13285 & w12723) | (w13285 & w44663) | (w12723 & w44663);
assign w13287 = ~w2285 & ~w12330;
assign w13288 = ~w12724 & w41163;
assign w13289 = w13283 & w13287;
assign w13290 = (~w13289 & w12723) | (~w13289 & w44664) | (w12723 & w44664);
assign w13291 = ~w13286 & w13290;
assign w13292 = ~w12616 & ~w13291;
assign w13293 = ~w12583 & w41164;
assign w13294 = ~w2285 & w12330;
assign w13295 = ~w13283 & w13294;
assign w13296 = (w13295 & w12723) | (w13295 & w44665) | (w12723 & w44665);
assign w13297 = ~w12724 & w41165;
assign w13298 = w12331 & w13283;
assign w13299 = (~w13298 & w12723) | (~w13298 & w44666) | (w12723 & w44666);
assign w13300 = ~w13296 & w13299;
assign w13301 = ~w13293 & w13300;
assign w13302 = ~w13292 & w13301;
assign w13303 = (w2006 & ~w13301) | (w2006 & w47301) | (~w13301 & w47301);
assign w13304 = ~w12585 & ~w12883;
assign w13305 = ~w12724 & ~w13304;
assign w13306 = ~w12394 & ~w12883;
assign w13307 = (w13306 & w12723) | (w13306 & w50336) | (w12723 & w50336);
assign w13308 = ~w12583 & w41166;
assign w13309 = ~w12616 & w13307;
assign w13310 = ~w13308 & ~w13309;
assign w13311 = w12346 & w12370;
assign w13312 = ~w2285 & ~w13311;
assign w13313 = (w13312 & w13309) | (w13312 & w41167) | (w13309 & w41167);
assign w13314 = ~w2285 & w13311;
assign w13315 = ~w13309 & w41168;
assign w13316 = ~w13313 & ~w13315;
assign w13317 = ~w13303 & ~w13316;
assign w13318 = w13301 & w47302;
assign w13319 = ~w1738 & ~w13258;
assign w13320 = (w13319 & w13264) | (w13319 & w41169) | (w13264 & w41169);
assign w13321 = ~w1738 & w13258;
assign w13322 = ~w13264 & w41170;
assign w13323 = ~w13320 & ~w13322;
assign w13324 = ~w13318 & w13323;
assign w13325 = ~w13317 & w13324;
assign w13326 = ~w12890 & w44667;
assign w13327 = w2285 & w13311;
assign w13328 = (w13327 & w13309) | (w13327 & w41171) | (w13309 & w41171);
assign w13329 = w2285 & ~w13311;
assign w13330 = ~w13309 & w41172;
assign w13331 = ~w13328 & ~w13330;
assign w13332 = ~w13303 & w13331;
assign w13333 = ~w13326 & w13332;
assign w13334 = w13325 & ~w13333;
assign w13335 = w13280 & ~w13334;
assign w13336 = w13257 & w13335;
assign w13337 = w13150 & w13336;
assign w13338 = w13280 & ~w13325;
assign w13339 = ~w1320 & w13082;
assign w13340 = ~w13273 & w44668;
assign w13341 = (w13274 & w13273) | (w13274 & w44669) | (w13273 & w44669);
assign w13342 = ~w13340 & ~w13341;
assign w13343 = ~w1541 & ~w13342;
assign w13344 = ~w13339 & ~w13343;
assign w13345 = ~w13338 & w13344;
assign w13346 = ~w13046 & w44670;
assign w13347 = w13034 & ~w13346;
assign w13348 = w13345 & w13347;
assign w13349 = w13150 & ~w13348;
assign w13350 = w13150 & w48754;
assign w13351 = w3 & ~w13189;
assign w13352 = ~w13191 & ~w13194;
assign w13353 = w13351 & ~w13352;
assign w13354 = w13208 & w13353;
assign w13355 = w13185 & ~w13354;
assign w13356 = w13209 & ~w13219;
assign w13357 = ~w13229 & w44671;
assign w13358 = (w252 & ~w44671) | (w252 & w50337) | (~w44671 & w50337);
assign w13359 = (~w351 & w13145) | (~w351 & w44672) | (w13145 & w44672);
assign w13360 = ~w13358 & ~w13359;
assign w13361 = w13106 & w50338;
assign w13362 = ~w493 & ~w12464;
assign w13363 = (w13362 & ~w41152) | (w13362 & w47303) | (~w41152 & w47303);
assign w13364 = ~w13361 & ~w13363;
assign w13365 = ~w13361 & w47304;
assign w13366 = w13129 & ~w13365;
assign w13367 = w400 & ~w13364;
assign w13368 = ~w13366 & ~w13367;
assign w13369 = w13255 & ~w13360;
assign w13370 = ~w13146 & w13255;
assign w13371 = ~w13368 & w13370;
assign w13372 = ~w13369 & ~w13371;
assign w13373 = ~w80 & w13218;
assign w13374 = w13242 & w13247;
assign w13375 = ~w13247 & w13249;
assign w13376 = ~w13374 & ~w13375;
assign w13377 = w57 & w13376;
assign w13378 = ~w13373 & ~w13377;
assign w13379 = w13355 & ~w13356;
assign w13380 = w13355 & w13378;
assign w13381 = (~w13379 & ~w13372) | (~w13379 & w44673) | (~w13372 & w44673);
assign w13382 = ~w13350 & ~w13381;
assign w13383 = w12996 & w13337;
assign w13384 = w13382 & ~w13383;
assign w13385 = ~w12745 & ~w12817;
assign w13386 = w7315 & ~w13385;
assign w13387 = ~w7315 & w13385;
assign w13388 = ~w13386 & ~w13387;
assign w13389 = (w12805 & w13384) | (w12805 & w44674) | (w13384 & w44674);
assign w13390 = ~w13384 & w44675;
assign w13391 = ~w13389 & ~w13390;
assign w13392 = w6769 & ~w13391;
assign w13393 = w12722 & ~w12728;
assign w13394 = w12696 & ~w12700;
assign w13395 = ~w12695 & w48755;
assign w13396 = ~w12732 & ~w12813;
assign w13397 = (w13396 & ~w48755) | (w13396 & w50544) | (~w48755 & w50544);
assign w13398 = ~w12709 & ~w13397;
assign w13399 = w7924 & ~w13398;
assign w13400 = ~w7924 & w13398;
assign w13401 = ~w13399 & ~w13400;
assign w13402 = (w13393 & w13384) | (w13393 & w44677) | (w13384 & w44677);
assign w13403 = ~w13384 & w44678;
assign w13404 = ~w13402 & ~w13403;
assign w13405 = ~w7315 & ~w13404;
assign w13406 = ~w13392 & ~w13405;
assign w13407 = ~w12806 & ~w12817;
assign w13408 = w13382 & w47305;
assign w13409 = ~w12791 & w52244;
assign w13410 = (w13409 & ~w13382) | (w13409 & w47306) | (~w13382 & w47306);
assign w13411 = ~w13408 & ~w13410;
assign w13412 = ~w12761 & w12784;
assign w13413 = ~w6264 & ~w13412;
assign w13414 = w13411 & w13413;
assign w13415 = ~w6264 & w13412;
assign w13416 = ~w13411 & w13415;
assign w13417 = ~w13414 & ~w13416;
assign w13418 = ~w12779 & ~w12794;
assign w13419 = w12792 & w52244;
assign w13420 = ~w12761 & ~w13419;
assign w13421 = w13418 & ~w13420;
assign w13422 = ~w13418 & w13420;
assign w13423 = ~w13421 & ~w13422;
assign w13424 = w12793 & w13384;
assign w13425 = ~w13384 & w13423;
assign w13426 = ~w13424 & ~w13425;
assign w13427 = w5745 & w13426;
assign w13428 = w13417 & ~w13427;
assign w13429 = w13406 & w13428;
assign w13430 = ~w9195 & w13394;
assign w13431 = w9195 & ~w13394;
assign w13432 = ~w13430 & ~w13431;
assign w13433 = ~w13384 & w13432;
assign w13434 = ~w8666 & w12812;
assign w13435 = (w13434 & w13384) | (w13434 & w44679) | (w13384 & w44679);
assign w13436 = ~w8666 & ~w12812;
assign w13437 = ~w13384 & w44680;
assign w13438 = ~w13435 & ~w13437;
assign w13439 = ~w12813 & ~w13395;
assign w13440 = w8666 & ~w13439;
assign w13441 = ~w8666 & w13439;
assign w13442 = ~w13440 & ~w13441;
assign w13443 = ~w7924 & w12708;
assign w13444 = (w13443 & w13384) | (w13443 & w44681) | (w13384 & w44681);
assign w13445 = ~w7924 & ~w12708;
assign w13446 = ~w13384 & w44682;
assign w13447 = ~w13444 & ~w13446;
assign w13448 = w13438 & w13447;
assign w13449 = ~w12678 & ~w12692;
assign w13450 = w12675 & ~w12700;
assign w13451 = ~w13449 & w50545;
assign w13452 = (w13450 & w13449) | (w13450 & w50546) | (w13449 & w50546);
assign w13453 = ~w13451 & ~w13452;
assign w13454 = ~w9195 & w12699;
assign w13455 = w13382 & w47307;
assign w13456 = ~w9195 & ~w13453;
assign w13457 = (w13456 & ~w13382) | (w13456 & w47308) | (~w13382 & w47308);
assign w13458 = ~w13455 & ~w13457;
assign w13459 = w8666 & w12812;
assign w13460 = ~w13384 & w50547;
assign w13461 = w8666 & ~w12812;
assign w13462 = (w13461 & w13384) | (w13461 & w44683) | (w13384 & w44683);
assign w13463 = w13458 & ~w13462;
assign w13464 = ~w13460 & w13463;
assign w13465 = w13448 & ~w13464;
assign w13466 = w7315 & w13404;
assign w13467 = (w12708 & w13384) | (w12708 & w44684) | (w13384 & w44684);
assign w13468 = ~w13384 & w44685;
assign w13469 = ~w13467 & ~w13468;
assign w13470 = w13372 & w13378;
assign w13471 = ~w13219 & ~w13470;
assign w13472 = ~w12995 & w13335;
assign w13473 = w13150 & w13472;
assign w13474 = ~w12986 & w13473;
assign w13475 = (~w41173 & w44686) | (~w41173 & w44687) | (w44686 & w44687);
assign w13476 = w12708 & w13210;
assign w13477 = ~w13475 & w48757;
assign w13478 = w7924 & ~w13477;
assign w13479 = w13469 & w13478;
assign w13480 = ~w13466 & ~w13479;
assign w13481 = ~w13465 & w13480;
assign w13482 = w13429 & ~w13481;
assign w13483 = ~w6769 & w13391;
assign w13484 = w6264 & ~w13412;
assign w13485 = ~w13415 & ~w13484;
assign w13486 = w13411 & ~w13485;
assign w13487 = ~w13411 & w13485;
assign w13488 = ~w13486 & ~w13487;
assign w13489 = ~w13483 & ~w13488;
assign w13490 = w13428 & ~w13489;
assign w13491 = ~w12918 & ~w12954;
assign w13492 = (~w12950 & w12804) | (~w12950 & w44688) | (w12804 & w44688);
assign w13493 = w13491 & w13492;
assign w13494 = ~w12830 & w13493;
assign w13495 = ~w12830 & w13492;
assign w13496 = ~w13491 & ~w13495;
assign w13497 = w13382 & w47309;
assign w13498 = ~w13494 & ~w13496;
assign w13499 = ~w13384 & w13498;
assign w13500 = ~w13497 & ~w13499;
assign w13501 = (w4430 & w13499) | (w4430 & w47310) | (w13499 & w47310);
assign w13502 = ~w12825 & ~w12950;
assign w13503 = w12792 & ~w12794;
assign w13504 = (w13503 & w12817) | (w13503 & w44689) | (w12817 & w44689);
assign w13505 = w12744 & w13503;
assign w13506 = w12696 & w13505;
assign w13507 = ~w12780 & ~w12794;
assign w13508 = ~w12826 & ~w13507;
assign w13509 = ~w13506 & w44690;
assign w13510 = ~w12801 & ~w13509;
assign w13511 = w13502 & ~w13510;
assign w13512 = ~w13502 & w13510;
assign w13513 = ~w13511 & ~w13512;
assign w13514 = w13382 & w47311;
assign w13515 = ~w13384 & ~w13513;
assign w13516 = ~w13514 & ~w13515;
assign w13517 = (~w4838 & w13515) | (~w4838 & w47312) | (w13515 & w47312);
assign w13518 = ~w13501 & ~w13517;
assign w13519 = ~w5745 & ~w13426;
assign w13520 = ~w13506 & w48758;
assign w13521 = ~w5745 & w13520;
assign w13522 = w5745 & ~w13520;
assign w13523 = ~w13521 & ~w13522;
assign w13524 = (~w12800 & w13384) | (~w12800 & w44691) | (w13384 & w44691);
assign w13525 = ~w13384 & w44692;
assign w13526 = ~w13524 & ~w13525;
assign w13527 = w5330 & w13526;
assign w13528 = ~w13519 & ~w13527;
assign w13529 = w13518 & w13528;
assign w13530 = ~w13490 & w13529;
assign w13531 = ~w13482 & w13530;
assign w13532 = ~w12891 & ~w13326;
assign w13533 = w12876 & w12984;
assign w13534 = ~w12830 & w13533;
assign w13535 = (~w12991 & ~w12987) | (~w12991 & w41174) | (~w12987 & w41174);
assign w13536 = ~w12989 & w13535;
assign w13537 = w12876 & ~w13536;
assign w13538 = w12857 & ~w13537;
assign w13539 = (~w12877 & w13534) | (~w12877 & w44693) | (w13534 & w44693);
assign w13540 = w13382 & w47313;
assign w13541 = (w13539 & ~w13382) | (w13539 & w47314) | (~w13382 & w47314);
assign w13542 = (w13532 & w13541) | (w13532 & w50615) | (w13541 & w50615);
assign w13543 = ~w13541 & w50616;
assign w13544 = ~w13542 & ~w13543;
assign w13545 = ~w2285 & ~w13544;
assign w13546 = w2285 & ~w13532;
assign w13547 = w13539 & w13546;
assign w13548 = w2285 & w13326;
assign w13549 = w13382 & w47315;
assign w13550 = ~w13384 & w13547;
assign w13551 = ~w13549 & ~w13550;
assign w13552 = w2285 & w13532;
assign w13553 = ~w13539 & w13552;
assign w13554 = ~w13384 & w13553;
assign w13555 = w2558 & w13552;
assign w13556 = w13382 & w47316;
assign w13557 = ~w13554 & ~w13556;
assign w13558 = w13551 & w13557;
assign w13559 = ~w12856 & ~w12877;
assign w13560 = w12845 & ~w13537;
assign w13561 = ~w13534 & w13560;
assign w13562 = (w13559 & w13534) | (w13559 & w44694) | (w13534 & w44694);
assign w13563 = ~w13534 & w44695;
assign w13564 = ~w13562 & ~w13563;
assign w13565 = w13382 & w47317;
assign w13566 = ~w13384 & ~w13564;
assign w13567 = ~w13566 & w47318;
assign w13568 = w13558 & ~w13567;
assign w13569 = w12845 & ~w12875;
assign w13570 = ~w12872 & ~w13536;
assign w13571 = ~w12872 & w12984;
assign w13572 = ~w12830 & w13571;
assign w13573 = (w13569 & w13572) | (w13569 & w44696) | (w13572 & w44696);
assign w13574 = ~w13572 & w44697;
assign w13575 = ~w13573 & ~w13574;
assign w13576 = ~w13384 & ~w13575;
assign w13577 = ~w12841 & ~w12873;
assign w13578 = w13382 & w47319;
assign w13579 = ~w13576 & ~w13578;
assign w13580 = (~w2896 & w13576) | (~w2896 & w47320) | (w13576 & w47320);
assign w13581 = (w2558 & w13566) | (w2558 & w47321) | (w13566 & w47321);
assign w13582 = ~w13580 & ~w13581;
assign w13583 = w13568 & ~w13582;
assign w13584 = ~w13545 & ~w13583;
assign w13585 = ~w13515 & w47322;
assign w13586 = ~w5330 & ~w12800;
assign w13587 = (w13586 & w13384) | (w13586 & w44698) | (w13384 & w44698);
assign w13588 = ~w5330 & w12800;
assign w13589 = ~w13384 & w44699;
assign w13590 = ~w13587 & ~w13589;
assign w13591 = ~w13585 & w13590;
assign w13592 = w13518 & ~w13591;
assign w13593 = w12948 & ~w12981;
assign w13594 = w4056 & ~w12987;
assign w13595 = ~w4056 & w12987;
assign w13596 = ~w13594 & ~w13595;
assign w13597 = ~w12830 & w48759;
assign w13598 = (w13596 & w12830) | (w13596 & w48760) | (w12830 & w48760);
assign w13599 = ~w13597 & ~w13598;
assign w13600 = ~w13384 & w13599;
assign w13601 = w3646 & ~w12973;
assign w13602 = (w13601 & w13384) | (w13601 & w44701) | (w13384 & w44701);
assign w13603 = w3646 & w12973;
assign w13604 = ~w13384 & w44702;
assign w13605 = ~w13602 & ~w13604;
assign w13606 = (~w12918 & w12830) | (~w12918 & w44703) | (w12830 & w44703);
assign w13607 = w13593 & ~w13606;
assign w13608 = ~w13593 & w13606;
assign w13609 = ~w13607 & ~w13608;
assign w13610 = w13382 & w47323;
assign w13611 = ~w13384 & w13609;
assign w13612 = ~w13610 & ~w13611;
assign w13613 = ~w13611 & w47324;
assign w13614 = w13605 & ~w13613;
assign w13615 = ~w12872 & ~w12989;
assign w13616 = (w13535 & w12830) | (w13535 & w44704) | (w12830 & w44704);
assign w13617 = w13615 & ~w13616;
assign w13618 = ~w13615 & w13616;
assign w13619 = ~w13617 & ~w13618;
assign w13620 = w13382 & w47325;
assign w13621 = ~w13384 & w13619;
assign w13622 = ~w13620 & ~w13621;
assign w13623 = ~w13621 & w47326;
assign w13624 = ~w13499 & w47327;
assign w13625 = ~w13623 & ~w13624;
assign w13626 = w13614 & w13625;
assign w13627 = ~w13592 & w13626;
assign w13628 = w13584 & w13627;
assign w13629 = ~a[52] & ~w13384;
assign w13630 = ~a[50] & ~a[51];
assign w13631 = ~a[52] & w13630;
assign w13632 = ~w12666 & ~w13631;
assign w13633 = ~a[53] & ~w13632;
assign w13634 = (w13633 & w13384) | (w13633 & w44705) | (w13384 & w44705);
assign w13635 = a[53] & w13632;
assign w13636 = ~w12617 & ~w13635;
assign w13637 = w12666 & w13631;
assign w13638 = w13349 & w44706;
assign w13639 = w13337 & w13636;
assign w13640 = w12996 & w13639;
assign w13641 = w13381 & w13636;
assign w13642 = ~w13640 & ~w13641;
assign w13643 = w13642 & w44707;
assign w13644 = ~w13634 & w13643;
assign w13645 = a[54] & ~w12666;
assign w13646 = ~a[54] & w12666;
assign w13647 = a[54] & ~w12617;
assign w13648 = ~w12618 & ~w13647;
assign w13649 = ~w13645 & ~w13646;
assign w13650 = w13382 & w47328;
assign w13651 = (w13648 & ~w13382) | (w13648 & w47329) | (~w13382 & w47329);
assign w13652 = ~w13650 & ~w13651;
assign w13653 = (w11870 & ~w13642) | (w11870 & w44708) | (~w13642 & w44708);
assign w13654 = w11870 & w13633;
assign w13655 = (w13654 & w13384) | (w13654 & w44709) | (w13384 & w44709);
assign w13656 = ~w13653 & ~w13655;
assign w13657 = ~w13653 & w48761;
assign w13658 = ~w13644 & ~w13652;
assign w13659 = w13657 & ~w13658;
assign w13660 = w12656 & ~w12661;
assign w13661 = w12631 & ~w13660;
assign w13662 = ~w12631 & w13660;
assign w13663 = ~w13661 & ~w13662;
assign w13664 = ~w12657 & ~w12659;
assign w13665 = w13382 & w47330;
assign w13666 = (w13663 & ~w13382) | (w13663 & w47331) | (~w13382 & w47331);
assign w13667 = ~w13665 & ~w13666;
assign w13668 = w10419 & w13667;
assign w13669 = ~w10419 & ~w13667;
assign w13670 = ~w13668 & ~w13669;
assign w13671 = ~w13659 & w13670;
assign w13672 = w12665 & ~w12678;
assign w13673 = w9781 & ~w12692;
assign w13674 = ~w13384 & w44710;
assign w13675 = w9781 & w12692;
assign w13676 = (w13675 & w13384) | (w13675 & w44711) | (w13384 & w44711);
assign w13677 = ~w13674 & ~w13676;
assign w13678 = ~w13668 & w13677;
assign w13679 = (w13678 & w13659) | (w13678 & w48762) | (w13659 & w48762);
assign w13680 = (~w11138 & w13653) | (~w11138 & w48763) | (w13653 & w48763);
assign w13681 = ~w11138 & ~w13652;
assign w13682 = ~w13644 & w13681;
assign w13683 = ~w13680 & ~w13682;
assign w13684 = ~w11870 & ~w12666;
assign w13685 = ~w13209 & w13684;
assign w13686 = ~w13353 & ~w13684;
assign w13687 = w13185 & w13686;
assign w13688 = ~w13685 & ~w13687;
assign w13689 = ~w13475 & w48764;
assign w13690 = ~w12619 & ~w12620;
assign w13691 = ~w12666 & ~w13690;
assign w13692 = w12666 & w13690;
assign w13693 = ~w13691 & ~w13692;
assign w13694 = a[55] & ~w13693;
assign w13695 = a[55] & ~w13646;
assign w13696 = ~a[55] & w13646;
assign w13697 = ~w13695 & ~w13696;
assign w13698 = (~w13697 & w13384) | (~w13697 & w44712) | (w13384 & w44712);
assign w13699 = ~a[55] & ~w13692;
assign w13700 = ~w13384 & w44713;
assign w13701 = ~w13698 & ~w13700;
assign w13702 = ~w13210 & w13694;
assign w13703 = ~w13689 & w13702;
assign w13704 = w13701 & ~w13703;
assign w13705 = w13678 & ~w13704;
assign w13706 = w13683 & w13705;
assign w13707 = (w12692 & w13384) | (w12692 & w44714) | (w13384 & w44714);
assign w13708 = ~w13384 & w44715;
assign w13709 = ~w13707 & ~w13708;
assign w13710 = ~w9781 & w13709;
assign w13711 = ~w12699 & w13384;
assign w13712 = ~w13384 & w13453;
assign w13713 = ~w13711 & ~w13712;
assign w13714 = w9195 & ~w13713;
assign w13715 = w13448 & ~w13710;
assign w13716 = ~w13714 & w13715;
assign w13717 = ~w13706 & w13716;
assign w13718 = ~w13679 & w13717;
assign w13719 = ~w13531 & w13628;
assign w13720 = w13584 & w14045;
assign w13721 = w13718 & w13720;
assign w13722 = ~w13719 & ~w13721;
assign w13723 = (w4056 & w13611) | (w4056 & w47332) | (w13611 & w47332);
assign w13724 = ~w3646 & w12973;
assign w13725 = (w13724 & w13384) | (w13724 & w44716) | (w13384 & w44716);
assign w13726 = ~w3646 & ~w12973;
assign w13727 = ~w13384 & w44717;
assign w13728 = ~w13725 & ~w13727;
assign w13729 = ~w13723 & w13728;
assign w13730 = w13605 & ~w13623;
assign w13731 = ~w13729 & w13730;
assign w13732 = ~w3242 & ~w13622;
assign w13733 = w2896 & w13579;
assign w13734 = ~w13732 & ~w13733;
assign w13735 = ~w13731 & w13734;
assign w13736 = ~w13545 & ~w13568;
assign w13737 = w13735 & ~w13736;
assign w13738 = w13584 & ~w13737;
assign w13739 = w13722 & ~w13738;
assign w13740 = ~w13065 & ~w13088;
assign w13741 = ~w12995 & w41175;
assign w13742 = (w13088 & w13338) | (w13088 & w44718) | (w13338 & w44718);
assign w13743 = ~w13065 & ~w13742;
assign w13744 = (w13743 & w12986) | (w13743 & w44719) | (w12986 & w44719);
assign w13745 = (w13044 & w13384) | (w13044 & w44720) | (w13384 & w44720);
assign w13746 = ~w12995 & w41176;
assign w13747 = ~w12986 & w13746;
assign w13748 = w13066 & ~w13742;
assign w13749 = (w13748 & w12986) | (w13748 & w44721) | (w12986 & w44721);
assign w13750 = ~w13045 & ~w13749;
assign w13751 = ~w13384 & w13750;
assign w13752 = (~w13045 & w13384) | (~w13045 & w44722) | (w13384 & w44722);
assign w13753 = ~w13745 & w13752;
assign w13754 = ~w13053 & ~w13744;
assign w13755 = w13045 & ~w13744;
assign w13756 = (~w13754 & w13384) | (~w13754 & w44723) | (w13384 & w44723);
assign w13757 = (w48765 & w50339) | (w48765 & w44723) | (w50339 & w44723);
assign w13758 = ~w13753 & w13757;
assign w13759 = ~w13021 & ~w13046;
assign w13760 = w612 & w13759;
assign w13761 = (w13760 & w13751) | (w13760 & w47334) | (w13751 & w47334);
assign w13762 = w612 & ~w13759;
assign w13763 = ~w13751 & w47335;
assign w13764 = ~w13761 & ~w13763;
assign w13765 = ~w13758 & w13764;
assign w13766 = ~w13751 & w47336;
assign w13767 = (w13759 & w13751) | (w13759 & w47337) | (w13751 & w47337);
assign w13768 = ~w13766 & ~w13767;
assign w13769 = ~w612 & w13768;
assign w13770 = ~w13765 & ~w13769;
assign w13771 = (~w13147 & w13090) | (~w13147 & w44724) | (w13090 & w44724);
assign w13772 = w13472 & w13771;
assign w13773 = ~w12986 & w13772;
assign w13774 = ~w13348 & w13771;
assign w13775 = (~w13774 & ~w13772) | (~w13774 & w41177) | (~w13772 & w41177);
assign w13776 = ~w13384 & ~w13775;
assign w13777 = ~w13110 & ~w13111;
assign w13778 = ~w13384 & w44725;
assign w13779 = ~w400 & ~w13364;
assign w13780 = (w48766 & w50340) | (w48766 & w44673) | (w50340 & w44673);
assign w13781 = w400 & w13364;
assign w13782 = (w48767 & w50341) | (w48767 & w44673) | (w50341 & w44673);
assign w13783 = (~w13780 & ~w13775) | (~w13780 & w44726) | (~w13775 & w44726);
assign w13784 = w351 & ~w13129;
assign w13785 = w13784 & w13783;
assign w13786 = ~w13778 & w13785;
assign w13787 = w351 & w13129;
assign w13788 = w13777 & w13787;
assign w13789 = ~w13384 & w44727;
assign w13790 = (w13775 & w48768) | (w13775 & w48769) | (w48768 & w48769);
assign w13791 = ~w13789 & ~w13790;
assign w13792 = ~w13786 & w13791;
assign w13793 = ~w13109 & w13364;
assign w13794 = ~w400 & w13793;
assign w13795 = (w13794 & w13776) | (w13794 & w47339) | (w13776 & w47339);
assign w13796 = ~w400 & ~w13793;
assign w13797 = ~w13776 & w47340;
assign w13798 = ~w13795 & ~w13797;
assign w13799 = w13792 & w13798;
assign w13800 = w400 & ~w13793;
assign w13801 = (w13800 & w13776) | (w13800 & w47341) | (w13776 & w47341);
assign w13802 = w400 & w13793;
assign w13803 = ~w13776 & w47342;
assign w13804 = ~w13801 & ~w13803;
assign w13805 = ~w13021 & ~w13047;
assign w13806 = ~w13021 & w13748;
assign w13807 = (~w13805 & w13747) | (~w13805 & w44728) | (w13747 & w44728);
assign w13808 = w13382 & w47343;
assign w13809 = ~w13384 & w13807;
assign w13810 = ~w13033 & ~w13147;
assign w13811 = w493 & w13810;
assign w13812 = (w13811 & w13809) | (w13811 & w47344) | (w13809 & w47344);
assign w13813 = w493 & ~w13810;
assign w13814 = ~w13809 & w47345;
assign w13815 = ~w13812 & ~w13814;
assign w13816 = w13804 & ~w13815;
assign w13817 = w13799 & ~w13816;
assign w13818 = ~w13770 & w13817;
assign w13819 = (w13333 & w12994) | (w13333 & w41178) | (w12994 & w41178);
assign w13820 = ~w13338 & ~w13343;
assign w13821 = (w13820 & w12986) | (w13820 & w48770) | (w12986 & w48770);
assign w13822 = ~w13083 & ~w13339;
assign w13823 = ~w13821 & w13822;
assign w13824 = ~w13339 & ~w13823;
assign w13825 = ~w13065 & ~w13087;
assign w13826 = w1320 & ~w12666;
assign w13827 = w12666 & ~w13058;
assign w13828 = ~w13826 & ~w13827;
assign w13829 = w13059 & ~w13828;
assign w13830 = ~w13059 & w13828;
assign w13831 = ~w13829 & ~w13830;
assign w13832 = w13384 & w13831;
assign w13833 = ~w13384 & w13825;
assign w13834 = ~w13824 & w13833;
assign w13835 = ~w13832 & ~w13834;
assign w13836 = ~w13384 & ~w13823;
assign w13837 = ~w13339 & ~w13825;
assign w13838 = ~w13384 & w50548;
assign w13839 = w945 & ~w13838;
assign w13840 = w13835 & w13839;
assign w13841 = ~w13753 & w13756;
assign w13842 = (~w754 & w13753) | (~w754 & w50549) | (w13753 & w50549);
assign w13843 = ~w13769 & ~w13842;
assign w13844 = w13765 & w13840;
assign w13845 = w13843 & ~w13844;
assign w13846 = (w13129 & w13778) | (w13129 & w50550) | (w13778 & w50550);
assign w13847 = ~w13778 & w50551;
assign w13848 = ~w13846 & ~w13847;
assign w13849 = ~w351 & w13848;
assign w13850 = (w13809 & w50617) | (w13809 & w50618) | (w50617 & w50618);
assign w13851 = (w13810 & w13809) | (w13810 & w50619) | (w13809 & w50619);
assign w13852 = w13850 & ~w13851;
assign w13853 = w13804 & ~w13852;
assign w13854 = w13799 & ~w13853;
assign w13855 = (~w13849 & w13853) | (~w13849 & w50552) | (w13853 & w50552);
assign w13856 = w13818 & ~w13845;
assign w13857 = w13855 & ~w13856;
assign w13858 = (~w13146 & w13366) | (~w13146 & w50553) | (w13366 & w50553);
assign w13859 = ~w13359 & ~w13858;
assign w13860 = ~w13349 & w13859;
assign w13861 = ~w13474 & w13860;
assign w13862 = ~w13474 & w41179;
assign w13863 = w13254 & ~w13377;
assign w13864 = (w13863 & ~w13382) | (w13863 & w47346) | (~w13382 & w47346);
assign w13865 = ~w13235 & ~w13862;
assign w13866 = w13864 & ~w13865;
assign w13867 = ~w13235 & w13377;
assign w13868 = ~w13235 & ~w13254;
assign w13869 = ~w13379 & w50192;
assign w13870 = ~w13867 & ~w13869;
assign w13871 = w13382 & w47347;
assign w13872 = ~w13862 & ~w13870;
assign w13873 = ~w13871 & ~w13872;
assign w13874 = ~w13866 & w13873;
assign w13875 = ~w80 & ~w13874;
assign w13876 = ~w13235 & ~w13358;
assign w13877 = (~w13876 & w13474) | (~w13876 & w41180) | (w13474 & w41180);
assign w13878 = ~w13384 & ~w13877;
assign w13879 = w13357 & ~w13381;
assign w13880 = (~w13879 & ~w13878) | (~w13879 & w44730) | (~w13878 & w44730);
assign w13881 = ~w57 & ~w13880;
assign w13882 = w80 & w13874;
assign w13883 = ~w13881 & ~w13882;
assign w13884 = w57 & w13880;
assign w13885 = w13364 & ~w13366;
assign w13886 = (w13131 & w13773) | (w13131 & w41181) | (w13773 & w41181);
assign w13887 = ~w13384 & w13886;
assign w13888 = ~w13146 & ~w13359;
assign w13889 = w252 & ~w13888;
assign w13890 = (w13889 & w13887) | (w13889 & w47349) | (w13887 & w47349);
assign w13891 = w252 & w13888;
assign w13892 = ~w13887 & w47350;
assign w13893 = ~w13890 & ~w13892;
assign w13894 = ~w13884 & w13893;
assign w13895 = (~w13875 & ~w13883) | (~w13875 & w49638) | (~w13883 & w49638);
assign w13896 = ~w13219 & ~w13373;
assign w13897 = w13255 & ~w13862;
assign w13898 = (~w13377 & ~w13382) | (~w13377 & w47351) | (~w13382 & w47351);
assign w13899 = ~w13897 & w13898;
assign w13900 = (w13896 & w13899) | (w13896 & w44731) | (w13899 & w44731);
assign w13901 = ~w13899 & w44732;
assign w13902 = ~w13900 & ~w13901;
assign w13903 = w3 & ~w13902;
assign w13904 = (w13198 & w13475) | (w13198 & w47352) | (w13475 & w47352);
assign w13905 = w13168 & w13178;
assign w13906 = ~w13168 & w13179;
assign w13907 = ~w13905 & ~w13906;
assign w13908 = ~w13175 & w13907;
assign w13909 = w11879 & ~w13154;
assign w13910 = w13154 & ~w13155;
assign w13911 = ~w13909 & ~w13910;
assign w13912 = w13908 & ~w13904;
assign w13913 = ~w13908 & w13911;
assign w13914 = (w13475 & w48771) | (w13475 & w48772) | (w48771 & w48772);
assign w13915 = ~w13912 & ~w13914;
assign w13916 = ~w42 & w13915;
assign w13917 = w13198 & ~w13353;
assign w13918 = w13382 & w47353;
assign w13919 = (w13917 & w13918) | (w13917 & w44733) | (w13918 & w44733);
assign w13920 = ~w13918 & w44734;
assign w13921 = ~w13919 & ~w13920;
assign w13922 = w13159 & ~w13908;
assign w13923 = w42 & ~w13922;
assign w13924 = ~w13904 & w13923;
assign w13925 = w42 & ~w13908;
assign w13926 = w13904 & w13925;
assign w13927 = ~w13924 & ~w13926;
assign w13928 = w13921 & ~w13927;
assign w13929 = ~w13916 & ~w13928;
assign w13930 = ~w13903 & ~w13929;
assign w13931 = w13895 & w13930;
assign w13932 = ~w3 & w13902;
assign w13933 = ~w13929 & w13932;
assign w13934 = (~w13933 & ~w13895) | (~w13933 & w44735) | (~w13895 & w44735);
assign w13935 = w13857 & ~w13934;
assign w13936 = ~w13834 & w50554;
assign w13937 = ~w945 & ~w13936;
assign w13938 = w13082 & w13384;
assign w13939 = w13821 & ~w13822;
assign w13940 = w1120 & w13938;
assign w13941 = w1120 & ~w13939;
assign w13942 = w13836 & w13941;
assign w13943 = ~w13940 & ~w13942;
assign w13944 = ~w13268 & w13323;
assign w13945 = ~w13317 & ~w13318;
assign w13946 = ~w13944 & ~w13945;
assign w13947 = (w41178 & w44736) | (w41178 & w44737) | (w44736 & w44737);
assign w13948 = (~w13946 & w12986) | (~w13946 & w44738) | (w12986 & w44738);
assign w13949 = ~w13268 & w13325;
assign w13950 = (w13949 & w12986) | (w13949 & w44739) | (w12986 & w44739);
assign w13951 = w13948 & ~w13950;
assign w13952 = w13382 & w47354;
assign w13953 = ~w13384 & w13951;
assign w13954 = ~w13952 & ~w13953;
assign w13955 = (w1541 & w13953) | (w1541 & w47355) | (w13953 & w47355);
assign w13956 = w13316 & w13331;
assign w13957 = (~w13326 & w12994) | (~w13326 & w41182) | (w12994 & w41182);
assign w13958 = w13956 & w13957;
assign w13959 = ~w12986 & w13958;
assign w13960 = ~w13303 & ~w13318;
assign w13961 = ~w12986 & w44740;
assign w13962 = w13316 & ~w13960;
assign w13963 = ~w13316 & w13960;
assign w13964 = ~w13962 & ~w13963;
assign w13965 = (w13964 & w12986) | (w13964 & w44741) | (w12986 & w44741);
assign w13966 = w13382 & w47356;
assign w13967 = ~w13961 & ~w13965;
assign w13968 = ~w13384 & w13967;
assign w13969 = ~w13966 & ~w13968;
assign w13970 = (w1738 & w13968) | (w1738 & w47357) | (w13968 & w47357);
assign w13971 = ~w13955 & ~w13970;
assign w13972 = w13310 & ~w13311;
assign w13973 = ~w13310 & w13311;
assign w13974 = ~w13972 & ~w13973;
assign w13975 = (~w13956 & w12986) | (~w13956 & w41183) | (w12986 & w41183);
assign w13976 = w13382 & w47358;
assign w13977 = ~w13959 & ~w13975;
assign w13978 = ~w13384 & w13977;
assign w13979 = ~w13976 & ~w13978;
assign w13980 = w2006 & w13979;
assign w13981 = w13971 & ~w13980;
assign w13982 = ~w13953 & w47359;
assign w13983 = ~w1320 & ~w13342;
assign w13984 = w13384 & ~w13983;
assign w13985 = ~w13268 & w13316;
assign w13986 = w13819 & w13985;
assign w13987 = ~w12986 & w13986;
assign w13988 = ~w13268 & ~w13325;
assign w13989 = ~w13987 & ~w13988;
assign w13990 = w13279 & ~w13343;
assign w13991 = ~w1320 & w13990;
assign w13992 = (w41184 & w12986) | (w41184 & w48773) | (w12986 & w48773);
assign w13993 = ~w1320 & ~w13990;
assign w13994 = (w13993 & w41185) | (w13993 & w13987) | (w41185 & w13987);
assign w13995 = ~w13992 & ~w13994;
assign w13996 = ~w13384 & w13995;
assign w13997 = ~w13984 & ~w13996;
assign w13998 = ~w13982 & ~w13997;
assign w13999 = ~w13968 & w47360;
assign w14000 = (~w2006 & w13978) | (~w2006 & w47361) | (w13978 & w47361);
assign w14001 = ~w13999 & ~w14000;
assign w14002 = w13971 & ~w14001;
assign w14003 = w13998 & ~w14002;
assign w14004 = ~w13981 & w14003;
assign w14005 = w1541 & w13384;
assign w14006 = ~w13384 & w13989;
assign w14007 = ~w14005 & ~w14006;
assign w14008 = w13990 & w14007;
assign w14009 = ~w13990 & ~w14007;
assign w14010 = ~w14008 & ~w14009;
assign w14011 = w1320 & ~w14010;
assign w14012 = (~w1120 & ~w13384) | (~w1120 & w50555) | (~w13384 & w50555);
assign w14013 = ~w13384 & w50556;
assign w14014 = w14012 & ~w14013;
assign w14015 = (~w14014 & w14010) | (~w14014 & w44742) | (w14010 & w44742);
assign w14016 = ~w13937 & ~w13943;
assign w14017 = ~w13937 & w14015;
assign w14018 = ~w14004 & w14017;
assign w14019 = (~w14016 & w14004) | (~w14016 & w44743) | (w14004 & w44743);
assign w14020 = w13943 & w13998;
assign w14021 = ~w14002 & w14020;
assign w14022 = w13818 & ~w14021;
assign w14023 = ~w14019 & w14022;
assign w14024 = w13935 & ~w14023;
assign w14025 = ~w13739 & w14024;
assign w14026 = (w13818 & w14018) | (w13818 & w41186) | (w14018 & w41186);
assign w14027 = w13935 & ~w14026;
assign w14028 = ~w13887 & w47362;
assign w14029 = (w13888 & w13887) | (w13888 & w47363) | (w13887 & w47363);
assign w14030 = ~w14028 & ~w14029;
assign w14031 = ~w252 & ~w14030;
assign w14032 = ~w14030 & w48774;
assign w14033 = w13883 & ~w14032;
assign w14034 = w13916 & w13921;
assign w14035 = (~w14034 & w13929) | (~w14034 & w47364) | (w13929 & w47364);
assign w14036 = w13931 & ~w14033;
assign w14037 = (w14035 & ~w13931) | (w14035 & w44744) | (~w13931 & w44744);
assign w14038 = (w14037 & ~w13935) | (w14037 & w44745) | (~w13935 & w44745);
assign w14039 = ~w14025 & w14038;
assign w14040 = (w13737 & w13856) | (w13737 & w44746) | (w13856 & w44746);
assign w14041 = w13737 & w13818;
assign w14042 = ~w14019 & w14041;
assign w14043 = ~w14040 & ~w14042;
assign w14044 = ~w13531 & w13627;
assign w14045 = w13429 & w13627;
assign w14046 = w13718 & w14045;
assign w14047 = ~w14044 & ~w14046;
assign w14048 = ~w14031 & w14047;
assign w14049 = ~w14043 & w14048;
assign w14050 = w13584 & w14021;
assign w14051 = w13818 & ~w14050;
assign w14052 = (~w14031 & w13856) | (~w14031 & w44747) | (w13856 & w44747);
assign w14053 = ~w14050 & w47365;
assign w14054 = ~w14019 & w14053;
assign w14055 = ~w14052 & ~w14054;
assign w14056 = ~w14054 & w44748;
assign w14057 = (w14056 & ~w14048) | (w14056 & w49639) | (~w14048 & w49639);
assign w14058 = ~w14036 & w41187;
assign w14059 = ~w14027 & w14058;
assign w14060 = ~w14025 & w14059;
assign w14061 = (~w80 & w14025) | (~w80 & w44749) | (w14025 & w44749);
assign w14062 = ~w14057 & w14060;
assign w14063 = ~w14061 & ~w14062;
assign w14064 = ~w13875 & ~w13882;
assign w14065 = ~w3 & w14064;
assign w14066 = (w14065 & w14062) | (w14065 & w44750) | (w14062 & w44750);
assign w14067 = ~w3 & ~w14064;
assign w14068 = ~w14062 & w44751;
assign w14069 = ~w14066 & ~w14068;
assign w14070 = w3 & ~w14064;
assign w14071 = (w14070 & w14062) | (w14070 & w44752) | (w14062 & w44752);
assign w14072 = w3 & w14064;
assign w14073 = ~w14062 & w44753;
assign w14074 = ~w14071 & ~w14073;
assign w14075 = w13458 & ~w13714;
assign w14076 = ~w13706 & ~w13710;
assign w14077 = ~w13679 & w14076;
assign w14078 = w14075 & w14077;
assign w14079 = (w13458 & ~w14077) | (w13458 & w47366) | (~w14077 & w47366);
assign w14080 = w8666 & ~w14079;
assign w14081 = ~w8666 & w14079;
assign w14082 = ~w14080 & ~w14081;
assign w14083 = w14039 & w14082;
assign w14084 = w12812 & ~w13433;
assign w14085 = ~w12812 & w13433;
assign w14086 = ~w14084 & ~w14085;
assign w14087 = w7924 & w14086;
assign w14088 = (w14087 & ~w14039) | (w14087 & w41188) | (~w14039 & w41188);
assign w14089 = w7924 & ~w14086;
assign w14090 = w14039 & w41189;
assign w14091 = ~w14088 & ~w14090;
assign w14092 = ~w14075 & ~w14077;
assign w14093 = (w13713 & w14025) | (w13713 & w44754) | (w14025 & w44754);
assign w14094 = ~w14078 & ~w14092;
assign w14095 = ~w14025 & w44755;
assign w14096 = ~w14093 & ~w14095;
assign w14097 = ~w8666 & w14096;
assign w14098 = ~w7924 & w14086;
assign w14099 = w14039 & w41190;
assign w14100 = ~w7924 & ~w14086;
assign w14101 = (w14100 & ~w14039) | (w14100 & w41191) | (~w14039 & w41191);
assign w14102 = ~w14099 & ~w14101;
assign w14103 = (w14091 & w14097) | (w14091 & w41192) | (w14097 & w41192);
assign w14104 = ~w13392 & ~w13483;
assign w14105 = w13481 & ~w13718;
assign w14106 = ~w13405 & ~w14105;
assign w14107 = w14104 & ~w14106;
assign w14108 = ~w14104 & w14106;
assign w14109 = ~w14107 & ~w14108;
assign w14110 = (w13391 & w14025) | (w13391 & w44756) | (w14025 & w44756);
assign w14111 = w14039 & ~w14109;
assign w14112 = ~w14110 & ~w14111;
assign w14113 = ~w14111 & w47367;
assign w14114 = w13438 & w13464;
assign w14115 = w7924 & w13469;
assign w14116 = w13447 & ~w14115;
assign w14117 = (w13438 & w14115) | (w13438 & w50557) | (w14115 & w50557);
assign w14118 = ~w14115 & w50558;
assign w14119 = ~w14117 & ~w14118;
assign w14120 = (~w14077 & w47368) | (~w14077 & w47369) | (w47368 & w47369);
assign w14121 = (w14077 & w47370) | (w14077 & w47371) | (w47370 & w47371);
assign w14122 = ~w14120 & ~w14121;
assign w14123 = (w13469 & w14025) | (w13469 & w44757) | (w14025 & w44757);
assign w14124 = ~w14025 & w44758;
assign w14125 = ~w14123 & ~w14124;
assign w14126 = ~w7315 & w14125;
assign w14127 = ~w13405 & ~w13466;
assign w14128 = ~w13465 & ~w13479;
assign w14129 = (w14128 & ~w13717) | (w14128 & w48775) | (~w13717 & w48775);
assign w14130 = w14127 & ~w14129;
assign w14131 = ~w14127 & w14129;
assign w14132 = ~w14130 & ~w14131;
assign w14133 = (~w14025 & w47372) | (~w14025 & w47373) | (w47372 & w47373);
assign w14134 = ~w14025 & w47374;
assign w14135 = w14133 & ~w14134;
assign w14136 = ~w14126 & ~w14135;
assign w14137 = w13429 & w13718;
assign w14138 = ~w13490 & ~w13519;
assign w14139 = ~w13482 & w14138;
assign w14140 = ~w14137 & w14139;
assign w14141 = ~w14137 & w47375;
assign w14142 = (~w5330 & w14137) | (~w5330 & w47376) | (w14137 & w47376);
assign w14143 = ~w14141 & ~w14142;
assign w14144 = ~w4838 & w13526;
assign w14145 = (w14144 & ~w14039) | (w14144 & w41195) | (~w14039 & w41195);
assign w14146 = ~w4838 & ~w13526;
assign w14147 = w14039 & w41196;
assign w14148 = ~w14145 & ~w14147;
assign w14149 = ~w13406 & w13489;
assign w14150 = w13481 & w13489;
assign w14151 = (~w14149 & w13718) | (~w14149 & w41197) | (w13718 & w41197);
assign w14152 = w14151 & w47377;
assign w14153 = (w5745 & ~w14151) | (w5745 & w47378) | (~w14151 & w47378);
assign w14154 = ~w14152 & ~w14153;
assign w14155 = w14039 & w14154;
assign w14156 = w5330 & ~w13426;
assign w14157 = (w14156 & ~w14039) | (w14156 & w41198) | (~w14039 & w41198);
assign w14158 = w14039 & w41199;
assign w14159 = ~w14157 & ~w14158;
assign w14160 = w14148 & w14159;
assign w14161 = (w13406 & w13718) | (w13406 & w41200) | (w13718 & w41200);
assign w14162 = ~w13483 & ~w14161;
assign w14163 = w13488 & ~w14162;
assign w14164 = w14151 & ~w14163;
assign w14165 = w13411 & ~w13412;
assign w14166 = ~w13411 & w13412;
assign w14167 = ~w14165 & ~w14166;
assign w14168 = w14039 & w14164;
assign w14169 = ~w14168 & w44760;
assign w14170 = (w6264 & w14111) | (w6264 & w44761) | (w14111 & w44761);
assign w14171 = ~w14169 & ~w14170;
assign w14172 = w14160 & w14171;
assign w14173 = w7315 & w13469;
assign w14174 = (w14173 & w14025) | (w14173 & w44762) | (w14025 & w44762);
assign w14175 = w7315 & ~w14122;
assign w14176 = ~w14025 & w47379;
assign w14177 = ~w14174 & ~w14176;
assign w14178 = ~w6769 & w13404;
assign w14179 = (w14178 & w14025) | (w14178 & w44763) | (w14025 & w44763);
assign w14180 = ~w6769 & w14132;
assign w14181 = ~w14025 & w48776;
assign w14182 = ~w14179 & ~w14181;
assign w14183 = w14177 & w14182;
assign w14184 = (~w14135 & ~w14182) | (~w14135 & w47380) | (~w14182 & w47380);
assign w14185 = ~w14113 & w14184;
assign w14186 = w14172 & ~w14185;
assign w14187 = ~w14113 & w14136;
assign w14188 = ~w14103 & w14187;
assign w14189 = w14186 & ~w14188;
assign w14190 = ~w13517 & ~w13585;
assign w14191 = ~w13490 & w13528;
assign w14192 = ~w13482 & w14191;
assign w14193 = (w13590 & w14137) | (w13590 & w41201) | (w14137 & w41201);
assign w14194 = w14190 & ~w14193;
assign w14195 = ~w14190 & w14193;
assign w14196 = ~w14194 & ~w14195;
assign w14197 = (w13516 & w14025) | (w13516 & w44764) | (w14025 & w44764);
assign w14198 = w14039 & w14196;
assign w14199 = ~w14197 & ~w14198;
assign w14200 = (~w4430 & w14198) | (~w4430 & w47381) | (w14198 & w47381);
assign w14201 = (~w13526 & ~w14039) | (~w13526 & w44765) | (~w14039 & w44765);
assign w14202 = w14039 & w44766;
assign w14203 = ~w14201 & ~w14202;
assign w14204 = w4838 & ~w14203;
assign w14205 = (w5745 & w14168) | (w5745 & w44767) | (w14168 & w44767);
assign w14206 = ~w5330 & w13426;
assign w14207 = (w14206 & ~w14039) | (w14206 & w41202) | (~w14039 & w41202);
assign w14208 = w14039 & w41203;
assign w14209 = ~w14207 & ~w14208;
assign w14210 = ~w14205 & w14209;
assign w14211 = w14160 & ~w14210;
assign w14212 = ~w14204 & ~w14211;
assign w14213 = ~w14211 & w41204;
assign w14214 = (w14213 & ~w14186) | (w14213 & w44768) | (~w14186 & w44768);
assign w14215 = ~w13580 & ~w13733;
assign w14216 = ~w13731 & ~w13732;
assign w14217 = (~w14215 & ~w14047) | (~w14215 & w41205) | (~w14047 & w41205);
assign w14218 = w14215 & w14216;
assign w14219 = w14047 & w14218;
assign w14220 = ~w14217 & ~w14219;
assign w14221 = (~w13579 & w14025) | (~w13579 & w44769) | (w14025 & w44769);
assign w14222 = w14039 & w14220;
assign w14223 = ~w14221 & ~w14222;
assign w14224 = ~w14222 & w44770;
assign w14225 = ~w13567 & ~w13581;
assign w14226 = w14218 & w14225;
assign w14227 = w14047 & w14226;
assign w14228 = ~w13580 & w14225;
assign w14229 = w13580 & ~w14225;
assign w14230 = ~w14228 & ~w14229;
assign w14231 = (w14230 & ~w14047) | (w14230 & w41206) | (~w14047 & w41206);
assign w14232 = ~w2896 & w13384;
assign w14233 = ~w13384 & w13561;
assign w14234 = ~w14232 & ~w14233;
assign w14235 = w13559 & ~w14234;
assign w14236 = ~w13559 & w14234;
assign w14237 = ~w14235 & ~w14236;
assign w14238 = (w14237 & w14025) | (w14237 & w44771) | (w14025 & w44771);
assign w14239 = ~w14227 & ~w14231;
assign w14240 = w14039 & w14239;
assign w14241 = ~w14238 & ~w14240;
assign w14242 = ~w14240 & w44772;
assign w14243 = ~w14224 & ~w14242;
assign w14244 = ~w13592 & ~w13624;
assign w14245 = ~w13531 & w14244;
assign w14246 = w13429 & w14244;
assign w14247 = w13718 & w14246;
assign w14248 = ~w14245 & ~w14247;
assign w14249 = w13605 & w13728;
assign w14250 = ~w13723 & ~w14249;
assign w14251 = w13613 & ~w14249;
assign w14252 = w13723 & w14249;
assign w14253 = ~w14251 & ~w14252;
assign w14254 = (w14253 & ~w14248) | (w14253 & w41207) | (~w14248 & w41207);
assign w14255 = ~w14248 & w44773;
assign w14256 = w14254 & ~w14255;
assign w14257 = w12973 & ~w13600;
assign w14258 = ~w12973 & w13600;
assign w14259 = ~w14257 & ~w14258;
assign w14260 = w14039 & w14256;
assign w14261 = (~w14259 & w14025) | (~w14259 & w44774) | (w14025 & w44774);
assign w14262 = ~w14260 & ~w14261;
assign w14263 = (~w3242 & w14260) | (~w3242 & w44775) | (w14260 & w44775);
assign w14264 = (~w13622 & w14025) | (~w13622 & w44776) | (w14025 & w44776);
assign w14265 = ~w13623 & ~w13732;
assign w14266 = w13605 & ~w13729;
assign w14267 = (~w14248 & w44777) | (~w14248 & w44778) | (w44777 & w44778);
assign w14268 = ~w14025 & w44779;
assign w14269 = (w14248 & w44780) | (w14248 & w44781) | (w44780 & w44781);
assign w14270 = (w41209 & w14025) | (w41209 & w47382) | (w14025 & w47382);
assign w14271 = w2896 & ~w14269;
assign w14272 = w14268 & w14271;
assign w14273 = ~w14270 & ~w14272;
assign w14274 = ~w14263 & w14273;
assign w14275 = w14243 & w14274;
assign w14276 = ~w13613 & ~w13723;
assign w14277 = w14248 & ~w14276;
assign w14278 = ~w14248 & w14276;
assign w14279 = ~w14277 & ~w14278;
assign w14280 = (w13612 & w14025) | (w13612 & w44782) | (w14025 & w44782);
assign w14281 = w14039 & ~w14279;
assign w14282 = ~w14280 & ~w14281;
assign w14283 = (w3646 & w14281) | (w3646 & w44783) | (w14281 & w44783);
assign w14284 = ~w13501 & ~w13624;
assign w14285 = ~w13517 & ~w13591;
assign w14286 = ~w13517 & w14192;
assign w14287 = ~w14137 & w14286;
assign w14288 = (w14284 & w14287) | (w14284 & w41210) | (w14287 & w41210);
assign w14289 = ~w14287 & w41211;
assign w14290 = ~w14288 & ~w14289;
assign w14291 = (~w13500 & w14025) | (~w13500 & w44784) | (w14025 & w44784);
assign w14292 = w14039 & ~w14290;
assign w14293 = ~w14291 & ~w14292;
assign w14294 = (w4056 & w14292) | (w4056 & w44785) | (w14292 & w44785);
assign w14295 = ~w14283 & w14294;
assign w14296 = ~w14281 & w44786;
assign w14297 = ~w14198 & w44787;
assign w14298 = ~w14296 & ~w14297;
assign w14299 = ~w14295 & w14298;
assign w14300 = w14275 & w14299;
assign w14301 = ~w12666 & w13384;
assign w14302 = w12666 & ~w13384;
assign w14303 = ~w14301 & ~w14302;
assign w14304 = ~w13631 & w14303;
assign w14305 = ~w13384 & w13636;
assign w14306 = ~w13634 & ~w14305;
assign w14307 = w14304 & ~w14306;
assign w14308 = ~a[53] & ~w14307;
assign w14309 = ~w14036 & w41212;
assign w14310 = ~w14027 & w14309;
assign w14311 = a[53] & ~w13629;
assign w14312 = (~w14311 & w14025) | (~w14311 & w49640) | (w14025 & w49640);
assign w14313 = ~w14019 & w14051;
assign w14314 = (~w14304 & w41213) | (~w14304 & w13933) | (w41213 & w13933);
assign w14315 = ~w13856 & w44788;
assign w14316 = ~w14313 & w14315;
assign w14317 = w13631 & ~w14303;
assign w14318 = w14304 & w14306;
assign w14319 = ~w14317 & ~w14318;
assign w14320 = ~w14316 & ~w14319;
assign w14321 = w14047 & ~w14319;
assign w14322 = ~w14043 & w14321;
assign w14323 = ~w14320 & ~w14322;
assign w14324 = w14039 & ~w14323;
assign w14325 = ~w14312 & ~w14324;
assign w14326 = ~w12666 & ~w13630;
assign w14327 = ~w14036 & w41214;
assign w14328 = ~a[53] & w13629;
assign w14329 = (w14328 & w14025) | (w14328 & w49641) | (w14025 & w49641);
assign w14330 = ~a[53] & w14317;
assign w14331 = ~w13384 & w14330;
assign w14332 = ~w14036 & w41215;
assign w14333 = ~w14027 & w14332;
assign w14334 = (~w14331 & w14025) | (~w14331 & w49642) | (w14025 & w49642);
assign w14335 = ~w14329 & w14334;
assign w14336 = ~w14325 & w14335;
assign w14337 = ~a[48] & ~a[49];
assign w14338 = ~a[50] & w14337;
assign w14339 = ~w13384 & w14338;
assign w14340 = w13384 & ~w14338;
assign w14341 = a[51] & w14340;
assign w14342 = ~w13630 & ~w14341;
assign w14343 = ~a[51] & ~w14340;
assign w14344 = ~w14339 & ~w14343;
assign w14345 = (w14344 & w14025) | (w14344 & w44789) | (w14025 & w44789);
assign w14346 = ~w14339 & ~w14342;
assign w14347 = ~w14025 & w44790;
assign w14348 = ~w14345 & ~w14347;
assign w14349 = a[52] & ~w13630;
assign w14350 = ~w13631 & ~w14349;
assign w14351 = a[52] & w13384;
assign w14352 = ~w13629 & ~w14351;
assign w14353 = ~w12666 & ~w14352;
assign w14354 = (w14353 & w14025) | (w14353 & w44791) | (w14025 & w44791);
assign w14355 = ~w12666 & ~w14350;
assign w14356 = ~w14025 & w44792;
assign w14357 = ~w14354 & ~w14356;
assign w14358 = w14348 & w14357;
assign w14359 = ~w13644 & w13656;
assign w14360 = ~w14036 & w41216;
assign w14361 = ~w14027 & w14360;
assign w14362 = ~w14025 & w14361;
assign w14363 = (w13681 & w14025) | (w13681 & w49643) | (w14025 & w49643);
assign w14364 = ~w11138 & w13652;
assign w14365 = ~w14025 & w49644;
assign w14366 = ~w14363 & ~w14365;
assign w14367 = w12666 & w14350;
assign w14368 = ~w14025 & w44793;
assign w14369 = w12666 & w14352;
assign w14370 = (w14369 & w14025) | (w14369 & w44794) | (w14025 & w44794);
assign w14371 = ~w14368 & ~w14370;
assign w14372 = w14366 & w14371;
assign w14373 = ~w14358 & w14372;
assign w14374 = ~w14325 & w49645;
assign w14375 = w14373 & ~w14374;
assign w14376 = w13652 & ~w14362;
assign w14377 = ~w13652 & w14362;
assign w14378 = ~w14376 & ~w14377;
assign w14379 = w11138 & ~w14378;
assign w14380 = ~w11870 & w14366;
assign w14381 = ~w14336 & w14380;
assign w14382 = ~w14379 & ~w14381;
assign w14383 = ~w14375 & w14382;
assign w14384 = ~w13659 & w13683;
assign w14385 = ~w14025 & w44795;
assign w14386 = ~w13704 & ~w14385;
assign w14387 = w10419 & ~w14386;
assign w14388 = w13704 & w14385;
assign w14389 = w14387 & ~w14388;
assign w14390 = (~w14389 & ~w14382) | (~w14389 & w49646) | (~w14382 & w49646);
assign w14391 = ~w10419 & ~w13704;
assign w14392 = (w14391 & ~w14039) | (w14391 & w41217) | (~w14039 & w41217);
assign w14393 = ~w10419 & w13704;
assign w14394 = w14039 & w41218;
assign w14395 = ~w14392 & ~w14394;
assign w14396 = w13683 & ~w13704;
assign w14397 = w13671 & ~w14396;
assign w14398 = (w9781 & w14397) | (w9781 & w41219) | (w14397 & w41219);
assign w14399 = ~w14397 & w41220;
assign w14400 = ~w14398 & ~w14399;
assign w14401 = w14037 & w14400;
assign w14402 = w9195 & w13709;
assign w14403 = (w14402 & w14025) | (w14402 & w49647) | (w14025 & w49647);
assign w14404 = w9195 & ~w13709;
assign w14405 = ~w14025 & w49648;
assign w14406 = ~w14403 & ~w14405;
assign w14407 = ~w13659 & ~w14396;
assign w14408 = ~w13670 & ~w14407;
assign w14409 = ~w14397 & ~w14408;
assign w14410 = ~w9781 & ~w13667;
assign w14411 = (w14410 & w14025) | (w14410 & w44796) | (w14025 & w44796);
assign w14412 = ~w9781 & ~w14409;
assign w14413 = ~w14025 & w44797;
assign w14414 = ~w14411 & ~w14413;
assign w14415 = w14406 & w14414;
assign w14416 = w14395 & w14415;
assign w14417 = (w14382 & w49649) | (w14382 & w49650) | (w49649 & w49650);
assign w14418 = w8666 & ~w14096;
assign w14419 = w14091 & ~w14418;
assign w14420 = ~w14126 & ~w14419;
assign w14421 = ~w14103 & w14420;
assign w14422 = (~w13709 & w14025) | (~w13709 & w49651) | (w14025 & w49651);
assign w14423 = ~w14025 & w49652;
assign w14424 = ~w14422 & ~w14423;
assign w14425 = ~w9195 & ~w14424;
assign w14426 = w9781 & w13667;
assign w14427 = (w14426 & w14025) | (w14426 & w44798) | (w14025 & w44798);
assign w14428 = w9781 & w14409;
assign w14429 = ~w14025 & w44799;
assign w14430 = ~w14427 & ~w14429;
assign w14431 = w14406 & ~w14430;
assign w14432 = ~w14425 & ~w14431;
assign w14433 = w14183 & w14432;
assign w14434 = w14172 & w14433;
assign w14435 = ~w14421 & w14434;
assign w14436 = (w14300 & w14189) | (w14300 & w41222) | (w14189 & w41222);
assign w14437 = w14434 & w44800;
assign w14438 = ~w14417 & w14437;
assign w14439 = ~w14436 & ~w14438;
assign w14440 = ~w13738 & w13981;
assign w14441 = ~w13982 & ~w14002;
assign w14442 = (w14441 & ~w13722) | (w14441 & w41223) | (~w13722 & w41223);
assign w14443 = ~w14036 & w41224;
assign w14444 = ~w14027 & w14443;
assign w14445 = ~w14025 & w44801;
assign w14446 = (~w13954 & w14025) | (~w13954 & w49653) | (w14025 & w49653);
assign w14447 = ~w14445 & ~w14446;
assign w14448 = ~w14036 & w41225;
assign w14449 = w13722 & w41226;
assign w14450 = w14001 & ~w14449;
assign w14451 = ~w13970 & ~w14450;
assign w14452 = (~w13982 & w14025) | (~w13982 & w49654) | (w14025 & w49654);
assign w14453 = w14451 & ~w14452;
assign w14454 = ~w14447 & ~w14453;
assign w14455 = (~w1320 & w14447) | (~w1320 & w50559) | (w14447 & w50559);
assign w14456 = w1320 & w14010;
assign w14457 = (w13722 & w48777) | (w13722 & w48778) | (w48777 & w48778);
assign w14458 = (w14003 & ~w13722) | (w14003 & w41227) | (~w13722 & w41227);
assign w14459 = ~w1320 & ~w14010;
assign w14460 = w14011 & w14442;
assign w14461 = ~w14442 & w14459;
assign w14462 = ~w14460 & ~w14461;
assign w14463 = (~w14010 & w14025) | (~w14010 & w48779) | (w14025 & w48779);
assign w14464 = w14462 & ~w14463;
assign w14465 = w14464 & w41228;
assign w14466 = ~w14455 & ~w14465;
assign w14467 = (~w1120 & ~w14464) | (~w1120 & w41229) | (~w14464 & w41229);
assign w14468 = (w1120 & w14025) | (w1120 & w44802) | (w14025 & w44802);
assign w14469 = ~w14011 & ~w14458;
assign w14470 = w14039 & w14469;
assign w14471 = w13943 & ~w14014;
assign w14472 = ~w945 & w14471;
assign w14473 = (w14472 & w14470) | (w14472 & w44803) | (w14470 & w44803);
assign w14474 = ~w945 & ~w14471;
assign w14475 = ~w14470 & w44804;
assign w14476 = ~w14473 & ~w14475;
assign w14477 = ~w14467 & w14476;
assign w14478 = ~w14466 & w14477;
assign w14479 = w945 & ~w14471;
assign w14480 = (w14479 & w14470) | (w14479 & w44805) | (w14470 & w44805);
assign w14481 = w945 & w14471;
assign w14482 = ~w14470 & w44806;
assign w14483 = ~w14480 & ~w14482;
assign w14484 = ~w13738 & ~w14019;
assign w14485 = w13722 & w14484;
assign w14486 = (~w14021 & w14018) | (~w14021 & w41230) | (w14018 & w41230);
assign w14487 = ~w13840 & ~w13842;
assign w14488 = w14487 & ~w14486;
assign w14489 = (w14488 & ~w13722) | (w14488 & w49655) | (~w13722 & w49655);
assign w14490 = ~w13840 & ~w14486;
assign w14491 = w754 & ~w13841;
assign w14492 = (w13722 & w49656) | (w13722 & w49657) | (w49656 & w49657);
assign w14493 = ~w14485 & w41232;
assign w14494 = ~w754 & w13841;
assign w14495 = (w14494 & w14485) | (w14494 & w41233) | (w14485 & w41233);
assign w14496 = ~w14493 & ~w14495;
assign w14497 = (w13841 & w14025) | (w13841 & w44807) | (w14025 & w44807);
assign w14498 = w14496 & ~w14497;
assign w14499 = w14039 & w41234;
assign w14500 = w14498 & ~w14499;
assign w14501 = w14498 & w41235;
assign w14502 = (~w13937 & ~w14039) | (~w13937 & w41236) | (~w14039 & w41236);
assign w14503 = ~w13840 & ~w13937;
assign w14504 = ~w13970 & ~w14001;
assign w14505 = w13998 & ~w14504;
assign w14506 = ~w14004 & w14015;
assign w14507 = ~w13943 & ~w14503;
assign w14508 = ~w14503 & w14506;
assign w14509 = ~w14507 & w52245;
assign w14510 = (w14039 & w44810) | (w14039 & w44811) | (w44810 & w44811);
assign w14511 = (~w13936 & w14025) | (~w13936 & w44812) | (w14025 & w44812);
assign w14512 = ~w754 & ~w14511;
assign w14513 = ~w14510 & w14512;
assign w14514 = w14483 & w41238;
assign w14515 = ~w14478 & w14514;
assign w14516 = ~w14447 & w50560;
assign w14517 = ~w14467 & ~w14516;
assign w14518 = (~w14465 & w14516) | (~w14465 & w41239) | (w14516 & w41239);
assign w14519 = w14476 & ~w14518;
assign w14520 = w14515 & ~w14519;
assign w14521 = w612 & ~w14500;
assign w14522 = w754 & w14509;
assign w14523 = ~w14502 & w14522;
assign w14524 = w754 & w14511;
assign w14525 = ~w14523 & ~w14524;
assign w14526 = ~w14501 & ~w14525;
assign w14527 = ~w14521 & ~w14526;
assign w14528 = (w13969 & w14025) | (w13969 & w48780) | (w14025 & w48780);
assign w14529 = ~w13980 & ~w14000;
assign w14530 = (w14529 & ~w13722) | (w14529 & w41240) | (~w13722 & w41240);
assign w14531 = ~w13970 & ~w13999;
assign w14532 = ~w13980 & w14531;
assign w14533 = (w13722 & w48781) | (w13722 & w48782) | (w48781 & w48782);
assign w14534 = ~w14025 & w48783;
assign w14535 = ~w14000 & ~w14531;
assign w14536 = (w14535 & ~w13722) | (w14535 & w48784) | (~w13722 & w48784);
assign w14537 = ~w14039 & w41241;
assign w14538 = ~w1541 & ~w14536;
assign w14539 = w14534 & w14538;
assign w14540 = ~w14537 & ~w14539;
assign w14541 = w13722 & w41242;
assign w14542 = (w13979 & w14025) | (w13979 & w44813) | (w14025 & w44813);
assign w14543 = ~w14530 & ~w14541;
assign w14544 = w14039 & w14543;
assign w14545 = ~w14542 & ~w14544;
assign w14546 = ~w14544 & w44814;
assign w14547 = w14540 & ~w14546;
assign w14548 = w14039 & w47383;
assign w14549 = ~w14528 & ~w14548;
assign w14550 = ~w14548 & w48785;
assign w14551 = (w1738 & w14544) | (w1738 & w44815) | (w14544 & w44815);
assign w14552 = ~w13545 & w13558;
assign w14553 = ~w13567 & ~w13582;
assign w14554 = w14552 & ~w14553;
assign w14555 = ~w14552 & w14553;
assign w14556 = ~w14554 & ~w14555;
assign w14557 = w14047 & w41243;
assign w14558 = (~w14556 & ~w14047) | (~w14556 & w41244) | (~w14047 & w41244);
assign w14559 = ~w14557 & ~w14558;
assign w14560 = (~w13544 & w14025) | (~w13544 & w44816) | (w14025 & w44816);
assign w14561 = w14039 & ~w14559;
assign w14562 = ~w14560 & ~w14561;
assign w14563 = ~w14561 & w44817;
assign w14564 = ~w14551 & ~w14563;
assign w14565 = (~w14550 & ~w14547) | (~w14550 & w47384) | (~w14547 & w47384);
assign w14566 = w14527 & w14565;
assign w14567 = (w14566 & ~w14515) | (w14566 & w47385) | (~w14515 & w47385);
assign w14568 = ~w14439 & w14567;
assign w14569 = w14039 & w41245;
assign w14570 = ~w14264 & ~w14569;
assign w14571 = ~w14569 & w44818;
assign w14572 = (w2558 & w14222) | (w2558 & w44819) | (w14222 & w44819);
assign w14573 = ~w14571 & ~w14572;
assign w14574 = w14243 & ~w14573;
assign w14575 = ~w14292 & w44820;
assign w14576 = ~w14260 & w44821;
assign w14577 = ~w14283 & ~w14576;
assign w14578 = ~w14296 & w14575;
assign w14579 = w14577 & ~w14578;
assign w14580 = w14275 & ~w14579;
assign w14581 = ~w14574 & ~w14580;
assign w14582 = w14566 & ~w14581;
assign w14583 = ~w14520 & w14582;
assign w14584 = (w14527 & w14478) | (w14527 & w41246) | (w14478 & w41246);
assign w14585 = (~w2285 & w14240) | (~w2285 & w44822) | (w14240 & w44822);
assign w14586 = (~w2006 & w14561) | (~w2006 & w44823) | (w14561 & w44823);
assign w14587 = ~w14585 & ~w14586;
assign w14588 = w14547 & w14587;
assign w14589 = w14565 & w41247;
assign w14590 = ~w14520 & w14589;
assign w14591 = (~w14584 & w14520) | (~w14584 & w41248) | (w14520 & w41248);
assign w14592 = (~w13880 & w14025) | (~w13880 & w49658) | (w14025 & w49658);
assign w14593 = w14039 & ~w14057;
assign w14594 = ~w14592 & ~w14593;
assign w14595 = w13881 & w14037;
assign w14596 = ~w13884 & ~w14595;
assign w14597 = w13893 & w14055;
assign w14598 = ~w14049 & w14597;
assign w14599 = ~w14596 & ~w14598;
assign w14600 = ~w14594 & ~w14599;
assign w14601 = (~w80 & w14594) | (~w80 & w41249) | (w14594 & w41249);
assign w14602 = (w80 & w14598) | (w80 & w41250) | (w14598 & w41250);
assign w14603 = ~w14594 & w14602;
assign w14604 = (w14037 & w14313) | (w14037 & w47386) | (w14313 & w47386);
assign w14605 = w14037 & w14047;
assign w14606 = ~w14043 & w14605;
assign w14607 = w252 & ~w14034;
assign w14608 = ~w13933 & w50193;
assign w14609 = ~w14030 & ~w14608;
assign w14610 = w14030 & w14608;
assign w14611 = ~w14609 & ~w14610;
assign w14612 = w13893 & ~w14031;
assign w14613 = (w14612 & w14606) | (w14612 & w44824) | (w14606 & w44824);
assign w14614 = ~w14606 & w44825;
assign w14615 = ~w14613 & ~w14614;
assign w14616 = ~w57 & ~w14615;
assign w14617 = ~w14603 & ~w14616;
assign w14618 = w13798 & w13804;
assign w14619 = ~w13770 & w13815;
assign w14620 = ~w13770 & w41251;
assign w14621 = (w14620 & w13737) | (w14620 & w49659) | (w13737 & w49659);
assign w14622 = ~w14019 & w14621;
assign w14623 = ~w13845 & w14619;
assign w14624 = ~w13852 & ~w14623;
assign w14625 = w13815 & ~w14021;
assign w14626 = w13770 & ~w13852;
assign w14627 = w14625 & ~w14626;
assign w14628 = (w14618 & w14623) | (w14618 & w41252) | (w14623 & w41252);
assign w14629 = w14618 & w14627;
assign w14630 = ~w14019 & w14629;
assign w14631 = ~w14628 & ~w14630;
assign w14632 = w13722 & w14622;
assign w14633 = w14631 & ~w14632;
assign w14634 = ~w14632 & w49660;
assign w14635 = w13792 & ~w13849;
assign w14636 = ~w14036 & w41253;
assign w14637 = ~w14027 & w14636;
assign w14638 = ~w14025 & w14637;
assign w14639 = ~w14036 & w41254;
assign w14640 = ~w14027 & w14639;
assign w14641 = ~w14025 & w14640;
assign w14642 = (~w13848 & w14025) | (~w13848 & w44826) | (w14025 & w44826);
assign w14643 = ~w14634 & w14641;
assign w14644 = ~w14642 & ~w14643;
assign w14645 = (~w252 & ~w14644) | (~w252 & w41255) | (~w14644 & w41255);
assign w14646 = ~w14618 & w14624;
assign w14647 = ~w14019 & w14627;
assign w14648 = w14646 & ~w14647;
assign w14649 = w13722 & w48786;
assign w14650 = w14648 & ~w14649;
assign w14651 = w400 & w13804;
assign w14652 = w13798 & ~w14651;
assign w14653 = ~w14039 & w14652;
assign w14654 = w14039 & w48787;
assign w14655 = ~w14653 & ~w14654;
assign w14656 = ~w14654 & w41256;
assign w14657 = ~w14645 & ~w14656;
assign w14658 = w14617 & w14657;
assign w14659 = (~w351 & w14654) | (~w351 & w41257) | (w14654 & w41257);
assign w14660 = w13845 & ~w14486;
assign w14661 = (~w13770 & w14485) | (~w13770 & w41258) | (w14485 & w41258);
assign w14662 = (w493 & w14025) | (w493 & w44827) | (w14025 & w44827);
assign w14663 = w14039 & ~w14661;
assign w14664 = ~w14662 & ~w14663;
assign w14665 = w13815 & ~w13852;
assign w14666 = w400 & ~w14665;
assign w14667 = ~w14663 & w44828;
assign w14668 = w400 & w14665;
assign w14669 = (w14668 & w14663) | (w14668 & w44829) | (w14663 & w44829);
assign w14670 = ~w14667 & ~w14669;
assign w14671 = ~w14659 & w14670;
assign w14672 = ~w400 & w14665;
assign w14673 = ~w14663 & w44830;
assign w14674 = ~w400 & ~w14665;
assign w14675 = (w14674 & w14663) | (w14674 & w44831) | (w14663 & w44831);
assign w14676 = ~w14673 & ~w14675;
assign w14677 = (~w612 & w14025) | (~w612 & w44832) | (w14025 & w44832);
assign w14678 = (~w13758 & w14485) | (~w13758 & w41259) | (w14485 & w41259);
assign w14679 = w14039 & w14678;
assign w14680 = ~w14677 & ~w14679;
assign w14681 = w13764 & ~w13769;
assign w14682 = ~w493 & ~w14681;
assign w14683 = (w14682 & w14679) | (w14682 & w44833) | (w14679 & w44833);
assign w14684 = ~w493 & w14681;
assign w14685 = ~w14679 & w44834;
assign w14686 = ~w14683 & ~w14685;
assign w14687 = w14676 & ~w14686;
assign w14688 = w14671 & ~w14687;
assign w14689 = w14658 & ~w14688;
assign w14690 = (w252 & ~w14638) | (w252 & w49661) | (~w14638 & w49661);
assign w14691 = w14644 & w14690;
assign w14692 = w57 & w14615;
assign w14693 = ~w14691 & ~w14692;
assign w14694 = w14617 & ~w14693;
assign w14695 = (~w14694 & w14688) | (~w14694 & w41260) | (w14688 & w41260);
assign w14696 = ~w14601 & w14695;
assign w14697 = ~w14583 & w14696;
assign w14698 = w14591 & w14697;
assign w14699 = ~w14568 & w14698;
assign w14700 = w493 & w14681;
assign w14701 = (w14700 & w14679) | (w14700 & w44835) | (w14679 & w44835);
assign w14702 = w493 & ~w14681;
assign w14703 = ~w14679 & w44836;
assign w14704 = ~w14701 & ~w14703;
assign w14705 = w14676 & w14704;
assign w14706 = w14671 & ~w14705;
assign w14707 = w14658 & ~w14706;
assign w14708 = (w14698 & w47387) | (w14698 & w47388) | (w47387 & w47388);
assign w14709 = (w14033 & w14313) | (w14033 & w47389) | (w14313 & w47389);
assign w14710 = w14033 & w14047;
assign w14711 = ~w14043 & w14710;
assign w14712 = (~w14709 & ~w14710) | (~w14709 & w49662) | (~w14710 & w49662);
assign w14713 = w13895 & ~w13903;
assign w14714 = (w14711 & w47390) | (w14711 & w47391) | (w47390 & w47391);
assign w14715 = ~w13916 & w13921;
assign w14716 = w14714 & ~w14715;
assign w14717 = ~w14036 & w41263;
assign w14718 = ~w14027 & w14717;
assign w14719 = ~w14025 & w14718;
assign w14720 = (~w3 & w14025) | (~w3 & w44837) | (w14025 & w44837);
assign w14721 = w14712 & w14719;
assign w14722 = ~w14720 & ~w14721;
assign w14723 = ~w13903 & ~w13932;
assign w14724 = ~w42 & ~w14723;
assign w14725 = (w14724 & w14721) | (w14724 & w44838) | (w14721 & w44838);
assign w14726 = ~w42 & w14723;
assign w14727 = ~w14721 & w44839;
assign w14728 = ~w14725 & ~w14727;
assign w14729 = (w14699 & w47392) | (w14699 & w47393) | (w47392 & w47393);
assign w14730 = w13921 & ~w14714;
assign w14731 = w14722 & ~w14723;
assign w14732 = ~w14722 & w14723;
assign w14733 = ~w14731 & ~w14732;
assign w14734 = ~w14730 & w14733;
assign w14735 = ~w42 & ~w14734;
assign w14736 = ~w14708 & w14735;
assign w14737 = ~w14729 & ~w14736;
assign w14738 = w42 & ~w14723;
assign w14739 = (~w14738 & w14721) | (~w14738 & w44842) | (w14721 & w44842);
assign w14740 = ~w14025 & w47394;
assign w14741 = w14714 & w14740;
assign w14742 = ~w14739 & ~w14741;
assign w14743 = w42 & w14723;
assign w14744 = ~w14721 & w44843;
assign w14745 = ~w14025 & w47395;
assign w14746 = ~w14714 & w14745;
assign w14747 = ~w14744 & ~w14746;
assign w14748 = ~w14716 & ~w14730;
assign w14749 = w14742 & w14747;
assign w14750 = ~w42 & ~w14748;
assign w14751 = ~w14749 & ~w14750;
assign w14752 = w14069 & w14728;
assign w14753 = ~w14751 & ~w14752;
assign w14754 = w14074 & ~w14601;
assign w14755 = ~w14694 & w14754;
assign w14756 = ~w14751 & w14755;
assign w14757 = ~w14689 & w14756;
assign w14758 = (~w14753 & ~w14756) | (~w14753 & w44844) | (~w14756 & w44844);
assign w14759 = w14707 & ~w14753;
assign w14760 = w14584 & w14759;
assign w14761 = ~w14758 & ~w14760;
assign w14762 = ~w14580 & w41264;
assign w14763 = ~w14438 & w41265;
assign w14764 = ~w14520 & w44845;
assign w14765 = ~w14763 & w14764;
assign w14766 = (w14761 & w14763) | (w14761 & w44846) | (w14763 & w44846);
assign w14767 = w14069 & w14074;
assign w14768 = (w41266 & ~w14698) | (w41266 & w44847) | (~w14698 & w44847);
assign w14769 = (w14698 & w44848) | (w14698 & w44849) | (w44848 & w44849);
assign w14770 = ~w14768 & ~w14769;
assign w14771 = ~w14766 & ~w14770;
assign w14772 = w14063 & ~w14064;
assign w14773 = ~w14063 & w14064;
assign w14774 = ~w14772 & ~w14773;
assign w14775 = w14766 & w14774;
assign w14776 = (~w14775 & w14770) | (~w14775 & w47396) | (w14770 & w47396);
assign w14777 = ~w14737 & w14776;
assign w14778 = (~w14691 & w14688) | (~w14691 & w48788) | (w14688 & w48788);
assign w14779 = w14657 & ~w14706;
assign w14780 = w14778 & ~w14779;
assign w14781 = (w14778 & w14520) | (w14778 & w47397) | (w14520 & w47397);
assign w14782 = w14591 & w14781;
assign w14783 = ~w14568 & w14782;
assign w14784 = (w14782 & w44850) | (w14782 & w44851) | (w44850 & w44851);
assign w14785 = ~w14766 & ~w14784;
assign w14786 = w57 & ~w14780;
assign w14787 = ~w14783 & w14786;
assign w14788 = (w14782 & w44852) | (w14782 & w44853) | (w44852 & w44853);
assign w14789 = ~w14784 & w48789;
assign w14790 = ~w80 & w14761;
assign w14791 = ~w14765 & w14790;
assign w14792 = ~w14601 & ~w14603;
assign w14793 = (~w14792 & w14765) | (~w14792 & w44854) | (w14765 & w44854);
assign w14794 = ~w3 & w14792;
assign w14795 = w14791 & w14794;
assign w14796 = w14794 & ~w14788;
assign w14797 = (~w14795 & ~w14785) | (~w14795 & w47398) | (~w14785 & w47398);
assign w14798 = ~w3 & w14793;
assign w14799 = (w14798 & ~w14785) | (w14798 & w47399) | (~w14785 & w47399);
assign w14800 = w14797 & ~w14799;
assign w14801 = w14785 & ~w14787;
assign w14802 = w80 & ~w14615;
assign w14803 = (w14802 & ~w14785) | (w14802 & w47400) | (~w14785 & w47400);
assign w14804 = w80 & w14615;
assign w14805 = w14785 & w47401;
assign w14806 = ~w14803 & ~w14805;
assign w14807 = w14800 & w14806;
assign w14808 = (w14686 & w14520) | (w14686 & w47402) | (w14520 & w47402);
assign w14809 = w14591 & w14808;
assign w14810 = (w14705 & ~w14809) | (w14705 & w44855) | (~w14809 & w44855);
assign w14811 = ~w14766 & ~w14810;
assign w14812 = ~w14810 & w41270;
assign w14813 = (w14809 & w44856) | (w14809 & w44857) | (w44856 & w44857);
assign w14814 = ~w14656 & ~w14659;
assign w14815 = ~w14655 & w14766;
assign w14816 = ~w14814 & ~w14766;
assign w14817 = ~w14813 & w14816;
assign w14818 = ~w14815 & ~w14817;
assign w14819 = ~w14810 & w47403;
assign w14820 = w14818 & w47404;
assign w14821 = ~w252 & w14766;
assign w14822 = w14656 & ~w14766;
assign w14823 = ~w14821 & ~w14822;
assign w14824 = ~w14812 & w14823;
assign w14825 = ~w14645 & ~w14691;
assign w14826 = ~w57 & ~w14825;
assign w14827 = (w14826 & w14812) | (w14826 & w47405) | (w14812 & w47405);
assign w14828 = ~w57 & w14825;
assign w14829 = ~w14812 & w47406;
assign w14830 = ~w14827 & ~w14829;
assign w14831 = ~w14820 & w14830;
assign w14832 = w14807 & w14831;
assign w14833 = ~w14583 & w14591;
assign w14834 = w14686 & w14704;
assign w14835 = (~w14834 & w14568) | (~w14834 & w41272) | (w14568 & w41272);
assign w14836 = w14809 & w44858;
assign w14837 = w14680 & ~w14681;
assign w14838 = ~w14680 & w14681;
assign w14839 = ~w14837 & ~w14838;
assign w14840 = ~w14839 & w14766;
assign w14841 = ~w14766 & ~w14835;
assign w14842 = (w14841 & w48790) | (w14841 & w48791) | (w48790 & w48791);
assign w14843 = w14670 & w14676;
assign w14844 = (w14809 & w44860) | (w14809 & w44861) | (w44860 & w44861);
assign w14845 = w14676 & w14766;
assign w14846 = w14844 & ~w14845;
assign w14847 = ~w14664 & ~w14665;
assign w14848 = w14664 & w14665;
assign w14849 = ~w14847 & ~w14848;
assign w14850 = w14761 & w14849;
assign w14851 = ~w14765 & w14850;
assign w14852 = w14670 & ~w14851;
assign w14853 = ~w14811 & w14852;
assign w14854 = ~w14846 & ~w14853;
assign w14855 = (w351 & w14853) | (w351 & w41274) | (w14853 & w41274);
assign w14856 = ~w14842 & ~w14855;
assign w14857 = ~w14510 & ~w14511;
assign w14858 = ~w14857 & w14766;
assign w14859 = ~w14520 & w44862;
assign w14860 = ~w14758 & ~w14859;
assign w14861 = w14483 & ~w14519;
assign w14862 = ~w14513 & w14861;
assign w14863 = w14565 & ~w14862;
assign w14864 = ~w14763 & w14863;
assign w14865 = ~w14478 & w14483;
assign w14866 = ~w14513 & w14865;
assign w14867 = ~w14761 & ~w14866;
assign w14868 = w14525 & ~w14867;
assign w14869 = ~w14860 & w14864;
assign w14870 = w14868 & ~w14869;
assign w14871 = w14300 & w14565;
assign w14872 = ~w14214 & w14871;
assign w14873 = w14435 & w14871;
assign w14874 = ~w14417 & w14873;
assign w14875 = ~w14872 & ~w14874;
assign w14876 = (w14565 & ~w41264) | (w14565 & w47407) | (~w41264 & w47407);
assign w14877 = ~w14874 & w44863;
assign w14878 = ~w14513 & w14525;
assign w14879 = ~w14861 & ~w14878;
assign w14880 = (w14879 & ~w14877) | (w14879 & w47408) | (~w14877 & w47408);
assign w14881 = (~w14858 & w14870) | (~w14858 & w44864) | (w14870 & w44864);
assign w14882 = w612 & ~w14881;
assign w14883 = (~w14526 & w14478) | (~w14526 & w44865) | (w14478 & w44865);
assign w14884 = ~w14876 & ~w14883;
assign w14885 = (~w14526 & ~w14515) | (~w14526 & w44866) | (~w14515 & w44866);
assign w14886 = (w14885 & ~w14875) | (w14885 & w41275) | (~w14875 & w41275);
assign w14887 = ~w14766 & w14886;
assign w14888 = w14500 & ~w14887;
assign w14889 = (w14866 & w14763) | (w14866 & w44867) | (w14763 & w44867);
assign w14890 = w14521 & w14758;
assign w14891 = ~w14501 & ~w14890;
assign w14892 = (w14875 & w47409) | (w14875 & w47410) | (w47409 & w47410);
assign w14893 = ~w14766 & w14892;
assign w14894 = w14525 & ~w14891;
assign w14895 = ~w14889 & w14894;
assign w14896 = ~w14893 & ~w14895;
assign w14897 = ~w14888 & w14896;
assign w14898 = w14896 & w44868;
assign w14899 = ~w14882 & ~w14898;
assign w14900 = w14856 & w14899;
assign w14901 = ~w14874 & w47411;
assign w14902 = (~w14516 & ~w14875) | (~w14516 & w44869) | (~w14875 & w44869);
assign w14903 = ~w14766 & w14902;
assign w14904 = ~w14465 & ~w14467;
assign w14905 = w945 & w14904;
assign w14906 = (w14905 & w14765) | (w14905 & w44870) | (w14765 & w44870);
assign w14907 = ~w14903 & w14906;
assign w14908 = w945 & ~w14904;
assign w14909 = ~w14765 & w44871;
assign w14910 = ~w14516 & w14908;
assign w14911 = (w14910 & ~w14875) | (w14910 & w44872) | (~w14875 & w44872);
assign w14912 = ~w14766 & w14911;
assign w14913 = ~w14909 & ~w14912;
assign w14914 = ~w14907 & w14913;
assign w14915 = (w14516 & w14859) | (w14516 & w41277) | (w14859 & w41277);
assign w14916 = ~w14455 & ~w14915;
assign w14917 = ~w14877 & ~w14916;
assign w14918 = ~w14766 & ~w14901;
assign w14919 = ~w1320 & ~w14761;
assign w14920 = w14877 & w14919;
assign w14921 = w14454 & ~w14920;
assign w14922 = ~w14916 & w48792;
assign w14923 = (w1120 & w14920) | (w1120 & w41278) | (w14920 & w41278);
assign w14924 = ~w14918 & w14923;
assign w14925 = ~w14922 & ~w14924;
assign w14926 = w14914 & w14925;
assign w14927 = ~w945 & ~w14904;
assign w14928 = (w14927 & w14765) | (w14927 & w44873) | (w14765 & w44873);
assign w14929 = ~w14903 & w14928;
assign w14930 = ~w945 & w14904;
assign w14931 = ~w14765 & w44874;
assign w14932 = ~w14516 & w14930;
assign w14933 = (w14932 & ~w14875) | (w14932 & w44875) | (~w14875 & w44875);
assign w14934 = ~w14766 & w14933;
assign w14935 = ~w14931 & ~w14934;
assign w14936 = ~w14929 & w14935;
assign w14937 = (w14874 & w48793) | (w14874 & w48794) | (w48793 & w48794);
assign w14938 = ~w14466 & ~w14467;
assign w14939 = ~w14761 & ~w14938;
assign w14940 = w14567 & w41280;
assign w14941 = ~w14763 & w14940;
assign w14942 = ~w14939 & ~w14941;
assign w14943 = ~w14937 & ~w14942;
assign w14944 = ~w945 & w14761;
assign w14945 = ~w14765 & w14944;
assign w14946 = w14476 & w14483;
assign w14947 = w754 & w14946;
assign w14948 = (w14947 & w14765) | (w14947 & w44876) | (w14765 & w44876);
assign w14949 = ~w14943 & w14948;
assign w14950 = w754 & ~w14946;
assign w14951 = (w14875 & w44877) | (w14875 & w44878) | (w44877 & w44878);
assign w14952 = ~w14942 & w14951;
assign w14953 = ~w14765 & w44879;
assign w14954 = ~w14952 & ~w14953;
assign w14955 = ~w14949 & w14954;
assign w14956 = w14936 & w14955;
assign w14957 = ~w14926 & w14956;
assign w14958 = ~w612 & w14881;
assign w14959 = ~w14943 & ~w14945;
assign w14960 = ~w754 & w14946;
assign w14961 = (w14960 & w14943) | (w14960 & w44880) | (w14943 & w44880);
assign w14962 = ~w754 & ~w14946;
assign w14963 = ~w14943 & w44881;
assign w14964 = ~w14961 & ~w14963;
assign w14965 = ~w14958 & w14964;
assign w14966 = ~w14957 & w14965;
assign w14967 = ~w14918 & ~w14921;
assign w14968 = ~w14917 & ~w14967;
assign w14969 = ~w14967 & w47412;
assign w14970 = w14914 & w14969;
assign w14971 = w14956 & ~w14970;
assign w14972 = w14966 & ~w14971;
assign w14973 = (w14900 & ~w14966) | (w14900 & w44882) | (~w14966 & w44882);
assign w14974 = (w44882 & w47413) | (w44882 & w47414) | (w47413 & w47414);
assign w14975 = (~w14841 & w48795) | (~w14841 & w48796) | (w48795 & w48796);
assign w14976 = (~w493 & ~w14896) | (~w493 & w44883) | (~w14896 & w44883);
assign w14977 = ~w14975 & ~w14976;
assign w14978 = (w252 & ~w14818) | (w252 & w47415) | (~w14818 & w47415);
assign w14979 = ~w351 & w14854;
assign w14980 = ~w14978 & ~w14979;
assign w14981 = w14856 & ~w14977;
assign w14982 = w14980 & ~w14981;
assign w14983 = w14832 & ~w14982;
assign w14984 = w14785 & w14788;
assign w14985 = ~w80 & w14615;
assign w14986 = (w14985 & ~w14785) | (w14985 & w47416) | (~w14785 & w47416);
assign w14987 = w14785 & w47417;
assign w14988 = ~w14986 & ~w14987;
assign w14989 = w57 & ~w14825;
assign w14990 = ~w14812 & w47418;
assign w14991 = w57 & w14825;
assign w14992 = (w14991 & w14812) | (w14991 & w47419) | (w14812 & w47419);
assign w14993 = ~w14990 & ~w14992;
assign w14994 = w14988 & w14993;
assign w14995 = w14807 & ~w14994;
assign w14996 = ~w14733 & ~w14766;
assign w14997 = ~w14708 & w14996;
assign w14998 = w14733 & ~w14766;
assign w14999 = w14708 & w14998;
assign w15000 = ~w14997 & ~w14999;
assign w15001 = w42 & ~w14775;
assign w15002 = (w14737 & ~w44884) | (w14737 & w47420) | (~w44884 & w47420);
assign w15003 = ~w14765 & w44885;
assign w15004 = ~w14793 & ~w15003;
assign w15005 = w3 & ~w15004;
assign w15006 = w14789 & w15005;
assign w15007 = w3 & w15004;
assign w15008 = ~w14789 & w15007;
assign w15009 = ~w15006 & ~w15008;
assign w15010 = ~w14777 & ~w15009;
assign w15011 = ~w15002 & ~w15010;
assign w15012 = ~w14995 & w15011;
assign w15013 = ~w14983 & w15012;
assign w15014 = ~w14974 & w15013;
assign w15015 = (~w14777 & ~w15013) | (~w14777 & w47421) | (~w15013 & w47421);
assign w15016 = ~w14546 & ~w14564;
assign w15017 = w14540 & ~w14550;
assign w15018 = w15016 & ~w15017;
assign w15019 = ~w15016 & w15017;
assign w15020 = ~w15018 & ~w15019;
assign w15021 = w14581 & ~w14585;
assign w15022 = ~w14563 & ~w14586;
assign w15023 = ~w14546 & ~w14551;
assign w15024 = w15022 & w15023;
assign w15025 = (w15020 & ~w14439) | (w15020 & w41281) | (~w14439 & w41281);
assign w15026 = w14439 & w41282;
assign w15027 = ~w15025 & ~w15026;
assign w15028 = w14761 & w50194;
assign w15029 = ~w14766 & ~w15027;
assign w15030 = ~w15028 & ~w15029;
assign w15031 = (~w1320 & w15029) | (~w1320 & w47423) | (w15029 & w47423);
assign w15032 = w1320 & w15030;
assign w15033 = ~w14438 & w41283;
assign w15034 = ~w14546 & w14564;
assign w15035 = (w15034 & ~w44886) | (w15034 & w47424) | (~w44886 & w47424);
assign w15036 = ~w14766 & w15035;
assign w15037 = (w15022 & ~w41283) | (w15022 & w44887) | (~w41283 & w44887);
assign w15038 = ~w14586 & ~w15023;
assign w15039 = w15038 & ~w15037;
assign w15040 = w14761 & w50195;
assign w15041 = ~w14766 & w15039;
assign w15042 = ~w15040 & ~w15041;
assign w15043 = ~w15036 & w15042;
assign w15044 = (w1541 & ~w15042) | (w1541 & w47426) | (~w15042 & w47426);
assign w15045 = ~w15032 & ~w15044;
assign w15046 = ~w15031 & ~w15045;
assign w15047 = (~w1541 & w14766) | (~w1541 & w47427) | (w14766 & w47427);
assign w15048 = w15042 & w15047;
assign w15049 = ~w15031 & ~w15048;
assign w15050 = ~w14562 & w14761;
assign w15051 = ~w14765 & w15050;
assign w15052 = w41283 & w44888;
assign w15053 = ~w15037 & ~w15052;
assign w15054 = ~w14766 & w15053;
assign w15055 = (w1738 & w14765) | (w1738 & w44889) | (w14765 & w44889);
assign w15056 = ~w15054 & w15055;
assign w15057 = w15049 & w15056;
assign w15058 = ~w15046 & ~w15057;
assign w15059 = w14274 & w14299;
assign w15060 = (w15059 & w14189) | (w15059 & w41284) | (w14189 & w41284);
assign w15061 = w14434 & w44890;
assign w15062 = ~w14417 & w15061;
assign w15063 = w14274 & ~w14579;
assign w15064 = ~w14571 & ~w15063;
assign w15065 = ~w14224 & ~w14572;
assign w15066 = w15064 & w15065;
assign w15067 = ~w15062 & w41285;
assign w15068 = (~w15065 & ~w41286) | (~w15065 & w44891) | (~w41286 & w44891);
assign w15069 = ~w15067 & ~w15068;
assign w15070 = ~w14766 & ~w15069;
assign w15071 = ~w14223 & w14761;
assign w15072 = ~w14765 & w15071;
assign w15073 = (w2285 & w14765) | (w2285 & w44892) | (w14765 & w44892);
assign w15074 = ~w15070 & w15073;
assign w15075 = w41285 & w44893;
assign w15076 = w2285 & ~w14223;
assign w15077 = w3096 & w14223;
assign w15078 = ~w15076 & ~w15077;
assign w15079 = (~w15078 & ~w41285) | (~w15078 & w44894) | (~w41285 & w44894);
assign w15080 = ~w15075 & ~w15079;
assign w15081 = ~w14766 & ~w15080;
assign w15082 = w2006 & w14241;
assign w15083 = ~w15081 & w15082;
assign w15084 = w2006 & ~w14241;
assign w15085 = w15081 & w15084;
assign w15086 = ~w15083 & ~w15085;
assign w15087 = ~w15074 & w15086;
assign w15088 = (~w14297 & w14189) | (~w14297 & w41287) | (w14189 & w41287);
assign w15089 = w14434 & w44895;
assign w15090 = ~w14417 & w15089;
assign w15091 = ~w14294 & ~w14296;
assign w15092 = (w15091 & w15090) | (w15091 & w41288) | (w15090 & w41288);
assign w15093 = w14273 & ~w14571;
assign w15094 = ~w14761 & ~w15093;
assign w15095 = w14567 & w41289;
assign w15096 = ~w14763 & w15095;
assign w15097 = ~w15094 & ~w15096;
assign w15098 = ~w14570 & w14761;
assign w15099 = ~w14765 & w15098;
assign w15100 = w15097 & ~w15099;
assign w15101 = ~w14263 & w52246;
assign w15102 = ~w14766 & w15101;
assign w15103 = w15100 & ~w15102;
assign w15104 = ~w14263 & ~w15093;
assign w15105 = w15104 & w52246;
assign w15106 = ~w14766 & w15105;
assign w15107 = (~w2558 & w14766) | (~w2558 & w48797) | (w14766 & w48797);
assign w15108 = ~w15103 & w15107;
assign w15109 = ~w14262 & w14766;
assign w15110 = w14262 & w14761;
assign w15111 = ~w14765 & w15110;
assign w15112 = (w44897 & w48798) | (w44897 & w48799) | (w48798 & w48799);
assign w15113 = ~w15111 & ~w15112;
assign w15114 = ~w14295 & ~w14296;
assign w15115 = ~w14263 & ~w14576;
assign w15116 = w15114 & ~w15115;
assign w15117 = ~w14283 & ~w14575;
assign w15118 = ~w15090 & w48800;
assign w15119 = w15116 & ~w15118;
assign w15120 = w2896 & w15109;
assign w15121 = w2896 & ~w15119;
assign w15122 = w15113 & w15121;
assign w15123 = ~w15120 & ~w15122;
assign w15124 = ~w15108 & w15123;
assign w15125 = w15087 & w15124;
assign w15126 = ~w15111 & w44898;
assign w15127 = ~w2896 & ~w15109;
assign w15128 = ~w15126 & w15127;
assign w15129 = ~w14283 & ~w14296;
assign w15130 = ~w14575 & ~w15129;
assign w15131 = w14294 & ~w15129;
assign w15132 = w14575 & w15129;
assign w15133 = ~w15131 & ~w15132;
assign w15134 = (w15133 & ~w41290) | (w15133 & w44899) | (~w41290 & w44899);
assign w15135 = ~w14283 & w15092;
assign w15136 = w15134 & ~w15135;
assign w15137 = ~w14282 & w14766;
assign w15138 = ~w14766 & w15136;
assign w15139 = ~w15137 & ~w15138;
assign w15140 = (w3242 & w15138) | (w3242 & w44900) | (w15138 & w44900);
assign w15141 = ~w15128 & ~w15140;
assign w15142 = ~w15138 & w44901;
assign w15143 = (w4056 & w15090) | (w4056 & w41291) | (w15090 & w41291);
assign w15144 = ~w15090 & w41292;
assign w15145 = ~w15143 & ~w15144;
assign w15146 = w14293 & w14761;
assign w15147 = ~w14765 & w15146;
assign w15148 = ~w14293 & ~w15145;
assign w15149 = ~w14766 & w15148;
assign w15150 = w14293 & w15145;
assign w15151 = ~w15147 & ~w15150;
assign w15152 = ~w15149 & w15151;
assign w15153 = ~w3646 & w15152;
assign w15154 = ~w15142 & ~w15153;
assign w15155 = w15141 & ~w15154;
assign w15156 = w15125 & ~w15155;
assign w15157 = w14148 & ~w14204;
assign w15158 = (~w14184 & w14103) | (~w14184 & w47428) | (w14103 & w47428);
assign w15159 = ~w14421 & w14433;
assign w15160 = ~w15158 & ~w15159;
assign w15161 = w14136 & w14416;
assign w15162 = ~w14103 & w15161;
assign w15163 = w14184 & w14416;
assign w15164 = ~w15162 & ~w15163;
assign w15165 = ~w14390 & ~w15164;
assign w15166 = ~w14113 & w14210;
assign w15167 = ~w14171 & w14210;
assign w15168 = w14159 & ~w15167;
assign w15169 = ~w15157 & ~w15166;
assign w15170 = w15168 & w15169;
assign w15171 = w15157 & ~w15168;
assign w15172 = ~w15170 & ~w15171;
assign w15173 = w15157 & w15166;
assign w15174 = (w15173 & w15165) | (w15173 & w44902) | (w15165 & w44902);
assign w15175 = ~w15157 & w15168;
assign w15176 = ~w15165 & w44903;
assign w15177 = ~w15176 & w49663;
assign w15178 = ~w14766 & w15177;
assign w15179 = w14203 & w14761;
assign w15180 = ~w14765 & w15179;
assign w15181 = (~w4430 & w14765) | (~w4430 & w44904) | (w14765 & w44904);
assign w15182 = ~w15178 & w15181;
assign w15183 = (w4056 & w15178) | (w4056 & w47429) | (w15178 & w47429);
assign w15184 = ~w4056 & ~w4430;
assign w15185 = (w15184 & w14765) | (w15184 & w44905) | (w14765 & w44905);
assign w15186 = ~w15178 & w15185;
assign w15187 = ~w14200 & ~w14297;
assign w15188 = ~w14189 & w14212;
assign w15189 = ~w14417 & w14435;
assign w15190 = (w15187 & w15189) | (w15187 & w47430) | (w15189 & w47430);
assign w15191 = ~w15189 & w47431;
assign w15192 = ~w15190 & ~w15191;
assign w15193 = ~w14199 & w14766;
assign w15194 = ~w14766 & w15192;
assign w15195 = ~w15193 & ~w15194;
assign w15196 = ~w15186 & w15195;
assign w15197 = ~w15183 & ~w15196;
assign w15198 = ~w14140 & w14155;
assign w15199 = w13426 & ~w14155;
assign w15200 = ~w15198 & ~w15199;
assign w15201 = w14159 & w14209;
assign w15202 = ~w14171 & ~w14205;
assign w15203 = ~w14113 & ~w14205;
assign w15204 = w15201 & ~w15202;
assign w15205 = ~w15165 & w44906;
assign w15206 = ~w15201 & w15203;
assign w15207 = (w15206 & w15165) | (w15206 & w44907) | (w15165 & w44907);
assign w15208 = ~w15205 & ~w15207;
assign w15209 = ~w15201 & w15202;
assign w15210 = w15201 & ~w15203;
assign w15211 = ~w15202 & w15210;
assign w15212 = ~w15209 & ~w15211;
assign w15213 = w15208 & w15212;
assign w15214 = w15200 & w14766;
assign w15215 = ~w14766 & ~w15213;
assign w15216 = ~w15214 & ~w15215;
assign w15217 = ~w15215 & w47432;
assign w15218 = (~w14113 & w15165) | (~w14113 & w44908) | (w15165 & w44908);
assign w15219 = ~w14170 & ~w15218;
assign w15220 = ~w15219 & ~w14766;
assign w15221 = ~w5745 & w14761;
assign w15222 = ~w14765 & w15221;
assign w15223 = ~w14169 & ~w14205;
assign w15224 = ~w5330 & ~w15223;
assign w15225 = (w15224 & w14765) | (w15224 & w44909) | (w14765 & w44909);
assign w15226 = ~w15220 & w15225;
assign w15227 = ~w5330 & w15223;
assign w15228 = ~w14765 & w44910;
assign w15229 = (w15227 & w15218) | (w15227 & w47433) | (w15218 & w47433);
assign w15230 = w15229 & ~w14766;
assign w15231 = ~w15228 & ~w15230;
assign w15232 = ~w15226 & w15231;
assign w15233 = ~w15217 & w15232;
assign w15234 = ~w15197 & w15233;
assign w15235 = ~w14416 & w14432;
assign w15236 = ~w14389 & w14432;
assign w15237 = (~w15235 & w14383) | (~w15235 & w41293) | (w14383 & w41293);
assign w15238 = (~w14103 & w15237) | (~w14103 & w44911) | (w15237 & w44911);
assign w15239 = (w15237 & w47434) | (w15237 & w47435) | (w47434 & w47435);
assign w15240 = w14761 & ~w15239;
assign w15241 = ~w14126 & w14177;
assign w15242 = w15238 & ~w15241;
assign w15243 = (w15242 & w14765) | (w15242 & w44912) | (w14765 & w44912);
assign w15244 = (~w14126 & w14765) | (~w14126 & w44913) | (w14765 & w44913);
assign w15245 = w14177 & w14419;
assign w15246 = w14103 & w14177;
assign w15247 = (~w15246 & w15237) | (~w15246 & w47436) | (w15237 & w47436);
assign w15248 = ~w14761 & w15247;
assign w15249 = w14764 & w15247;
assign w15250 = ~w14763 & w15249;
assign w15251 = ~w15248 & ~w15250;
assign w15252 = w15242 & w50196;
assign w15253 = ~w15250 & w41294;
assign w15254 = w15244 & w15253;
assign w15255 = ~w15252 & ~w15254;
assign w15256 = ~w14126 & ~w15246;
assign w15257 = (w15256 & w15237) | (w15256 & w48802) | (w15237 & w48802);
assign w15258 = ~w14761 & ~w15257;
assign w15259 = w14764 & ~w15257;
assign w15260 = ~w14763 & w15259;
assign w15261 = ~w15258 & ~w15260;
assign w15262 = w6769 & w14761;
assign w15263 = ~w14765 & w15262;
assign w15264 = w15261 & ~w15263;
assign w15265 = ~w14135 & w14182;
assign w15266 = w6264 & w15265;
assign w15267 = (w15266 & ~w15261) | (w15266 & w41295) | (~w15261 & w41295);
assign w15268 = w6264 & ~w15265;
assign w15269 = w15261 & w41296;
assign w15270 = ~w15267 & ~w15269;
assign w15271 = w15255 & w15270;
assign w15272 = w14083 & w14086;
assign w15273 = ~w14083 & ~w14086;
assign w15274 = ~w15272 & ~w15273;
assign w15275 = w14102 & w14419;
assign w15276 = (w15275 & ~w15237) | (w15275 & w47437) | (~w15237 & w47437);
assign w15277 = ~w14761 & ~w15276;
assign w15278 = w14764 & ~w15276;
assign w15279 = ~w14763 & w15278;
assign w15280 = ~w15277 & ~w15279;
assign w15281 = w14761 & ~w15274;
assign w15282 = ~w14765 & w15281;
assign w15283 = w15280 & ~w15282;
assign w15284 = (~w14418 & ~w15237) | (~w14418 & w47438) | (~w15237 & w47438);
assign w15285 = ~w14091 & ~w15284;
assign w15286 = w14761 & ~w15285;
assign w15287 = w14091 & w14102;
assign w15288 = ~w15284 & ~w15287;
assign w15289 = ~w14765 & w15286;
assign w15290 = w15288 & ~w15289;
assign w15291 = ~w15283 & ~w15290;
assign w15292 = ~w15283 & w41297;
assign w15293 = w15244 & w15251;
assign w15294 = w6769 & ~w15243;
assign w15295 = ~w15293 & w15294;
assign w15296 = ~w15292 & ~w15295;
assign w15297 = (w7315 & w15283) | (w7315 & w41298) | (w15283 & w41298);
assign w15298 = ~w14415 & ~w14425;
assign w15299 = w15298 & w50197;
assign w15300 = ~w8666 & w15299;
assign w15301 = ~w15284 & ~w15300;
assign w15302 = w14418 & w15237;
assign w15303 = ~w15299 & w15302;
assign w15304 = w15301 & ~w15303;
assign w15305 = w14097 & ~w15237;
assign w15306 = (~w15305 & w14765) | (~w15305 & w44914) | (w14765 & w44914);
assign w15307 = ~w14766 & w15304;
assign w15308 = w15306 & ~w15307;
assign w15309 = (~w7924 & w15307) | (~w7924 & w48803) | (w15307 & w48803);
assign w15310 = ~w15297 & w15309;
assign w15311 = w15296 & ~w15310;
assign w15312 = w9781 & w50197;
assign w15313 = (w14383 & w47439) | (w14383 & w47440) | (w47439 & w47440);
assign w15314 = ~w15312 & ~w15313;
assign w15315 = w14764 & ~w15314;
assign w15316 = ~w14763 & w15315;
assign w15317 = w13667 & ~w14039;
assign w15318 = w14039 & w14409;
assign w15319 = ~w15317 & ~w15318;
assign w15320 = ~w15316 & w41300;
assign w15321 = (w15319 & w15316) | (w15319 & w41301) | (w15316 & w41301);
assign w15322 = ~w15320 & ~w15321;
assign w15323 = ~w9195 & ~w15322;
assign w15324 = w14406 & ~w14425;
assign w15325 = w14430 & w50197;
assign w15326 = w14414 & ~w15325;
assign w15327 = w15324 & w15326;
assign w15328 = w14430 & ~w15324;
assign w15329 = ~w15326 & w15328;
assign w15330 = ~w15327 & ~w15329;
assign w15331 = w14424 & w14766;
assign w15332 = ~w14766 & ~w15330;
assign w15333 = ~w15331 & ~w15332;
assign w15334 = ~w15332 & w47441;
assign w15335 = ~w15323 & ~w15334;
assign w15336 = w9195 & ~w15319;
assign w15337 = (w15336 & w15316) | (w15336 & w41302) | (w15316 & w41302);
assign w15338 = w9195 & w15319;
assign w15339 = ~w15316 & w41303;
assign w15340 = ~w15337 & ~w15339;
assign w15341 = w14383 & ~w14761;
assign w15342 = w14567 & w41304;
assign w15343 = ~w14763 & w15342;
assign w15344 = ~w15341 & ~w15343;
assign w15345 = w10419 & w14761;
assign w15346 = ~w14765 & w15345;
assign w15347 = w15344 & ~w15346;
assign w15348 = ~w14389 & w14395;
assign w15349 = ~w9781 & ~w15348;
assign w15350 = w15347 & w15349;
assign w15351 = ~w9781 & w15348;
assign w15352 = ~w15347 & w15351;
assign w15353 = ~w15350 & ~w15352;
assign w15354 = w15340 & w15353;
assign w15355 = w15335 & ~w15354;
assign w15356 = ~w6264 & ~w15265;
assign w15357 = (w15356 & ~w15261) | (w15356 & w41305) | (~w15261 & w41305);
assign w15358 = ~w6264 & w15265;
assign w15359 = w15261 & w41306;
assign w15360 = ~w15357 & ~w15359;
assign w15361 = w14112 & w14761;
assign w15362 = ~w14765 & w15361;
assign w15363 = ~w14113 & ~w14170;
assign w15364 = ~w15165 & w44915;
assign w15365 = w14761 & ~w15364;
assign w15366 = ~w14765 & w15365;
assign w15367 = (~w15363 & w15165) | (~w15363 & w48804) | (w15165 & w48804);
assign w15368 = ~w15165 & w48805;
assign w15369 = ~w15367 & ~w15368;
assign w15370 = ~w15366 & w15369;
assign w15371 = ~w15362 & ~w15370;
assign w15372 = (w5745 & w15370) | (w5745 & w44916) | (w15370 & w44916);
assign w15373 = w15360 & ~w15372;
assign w15374 = (~w8666 & w15332) | (~w8666 & w47442) | (w15332 & w47442);
assign w15375 = w15360 & w44917;
assign w15376 = ~w15355 & w15375;
assign w15377 = w15271 & ~w15311;
assign w15378 = w15376 & ~w15377;
assign w15379 = ~w14358 & w14371;
assign w15380 = ~w11870 & w15379;
assign w15381 = w11870 & ~w15379;
assign w15382 = ~w15380 & ~w15381;
assign w15383 = w15382 & ~w14766;
assign w15384 = w11138 & ~w14336;
assign w15385 = ~w15383 & w15384;
assign w15386 = w11138 & w14336;
assign w15387 = w15383 & w15386;
assign w15388 = ~w15385 & ~w15387;
assign w15389 = w14039 & w14350;
assign w15390 = ~w14039 & w14352;
assign w15391 = ~w15389 & ~w15390;
assign w15392 = ~w12666 & w14348;
assign w15393 = w14761 & w15391;
assign w15394 = ~w14765 & w15393;
assign w15395 = ~w15391 & w15392;
assign w15396 = ~w14763 & w44918;
assign w15397 = ~w15394 & ~w15396;
assign w15398 = ~w14584 & w14757;
assign w15399 = ~w14590 & w15398;
assign w15400 = w15398 & w50342;
assign w15401 = ~w14568 & w15400;
assign w15402 = ~w14758 & ~w14759;
assign w15403 = ~w14348 & ~w14371;
assign w15404 = (w15403 & w14758) | (w15403 & w47443) | (w14758 & w47443);
assign w15405 = (w15404 & ~w15400) | (w15404 & w44919) | (~w15400 & w44919);
assign w15406 = w12666 & ~w14348;
assign w15407 = ~w15392 & ~w15406;
assign w15408 = w15391 & w15407;
assign w15409 = (~w15408 & w14761) | (~w15408 & w41307) | (w14761 & w41307);
assign w15410 = w11870 & w15409;
assign w15411 = ~w15405 & w15410;
assign w15412 = w15397 & w15411;
assign w15413 = ~a[50] & w14039;
assign w15414 = ~a[50] & a[51];
assign w15415 = ~w12666 & ~w15414;
assign w15416 = ~a[51] & ~w15413;
assign w15417 = w15415 & ~w15416;
assign w15418 = ~w14339 & ~w14340;
assign w15419 = w14039 & w15418;
assign w15420 = a[51] & ~w15419;
assign w15421 = ~a[51] & w15419;
assign w15422 = ~w15420 & ~w15421;
assign w15423 = ~w14039 & ~w15418;
assign w15424 = ~w12666 & ~w15423;
assign w15425 = w15422 & w15424;
assign w15426 = ~w14761 & ~w15425;
assign w15427 = w14567 & w41308;
assign w15428 = ~w14763 & w15427;
assign w15429 = ~w15426 & ~w15428;
assign w15430 = w14761 & ~w15417;
assign w15431 = ~w14765 & w15430;
assign w15432 = w15429 & ~w15431;
assign w15433 = ~w14039 & ~w14752;
assign w15434 = ~w14751 & w15433;
assign w15435 = ~w15423 & ~w15434;
assign w15436 = ~w15434 & w41309;
assign w15437 = w14695 & w14754;
assign w15438 = w15436 & ~w15437;
assign w15439 = w14707 & w15435;
assign w15440 = w14567 & w15439;
assign w15441 = ~w15438 & ~w15440;
assign w15442 = (~w14039 & w14761) | (~w14039 & w15423) | (w14761 & w15423);
assign w15443 = ~w14763 & ~w15441;
assign w15444 = a[51] & ~w12666;
assign w15445 = ~w15443 & w41310;
assign w15446 = ~w15432 & ~w15445;
assign w15447 = (w15409 & w15401) | (w15409 & w41311) | (w15401 & w41311);
assign w15448 = w15397 & w15447;
assign w15449 = ~w15412 & ~w15446;
assign w15450 = (~w11870 & ~w15447) | (~w11870 & w47444) | (~w15447 & w47444);
assign w15451 = ~w15449 & ~w15450;
assign w15452 = a[50] & ~w14039;
assign w15453 = ~w15413 & ~w15452;
assign w15454 = (~w15453 & w14520) | (~w15453 & w47445) | (w14520 & w47445);
assign w15455 = w15399 & w15454;
assign w15456 = ~w14568 & w15455;
assign w15457 = a[50] & ~w14337;
assign w15458 = ~w14338 & ~w15457;
assign w15459 = w14565 & ~w15458;
assign w15460 = ~w14860 & w41312;
assign w15461 = ~w14759 & ~w15453;
assign w15462 = ~w14758 & w15461;
assign w15463 = ~w14761 & ~w15458;
assign w15464 = ~w13384 & ~w15462;
assign w15465 = ~w15463 & w15464;
assign w15466 = ~a[46] & ~a[47];
assign w15467 = ~a[48] & w15466;
assign w15468 = ~w14039 & ~w15467;
assign w15469 = a[48] & ~a[49];
assign w15470 = w14039 & w15467;
assign w15471 = ~w15469 & ~w15470;
assign w15472 = a[49] & ~w15468;
assign w15473 = w15471 & ~w15472;
assign w15474 = ~w14761 & w15473;
assign w15475 = w14567 & w41313;
assign w15476 = ~w14763 & w15475;
assign w15477 = ~w15474 & ~w15476;
assign w15478 = ~a[49] & ~w15468;
assign w15479 = ~w15470 & ~w15478;
assign w15480 = w14761 & w15479;
assign w15481 = ~w14765 & w15480;
assign w15482 = w15477 & ~w15481;
assign w15483 = ~w15456 & w47446;
assign w15484 = ~w15482 & ~w15483;
assign w15485 = ~w15462 & ~w15463;
assign w15486 = ~w15456 & w15485;
assign w15487 = ~w15460 & w15486;
assign w15488 = (w13384 & ~w15486) | (w13384 & w41314) | (~w15486 & w41314);
assign w15489 = ~w15484 & ~w15488;
assign w15490 = a[51] & ~w15413;
assign w15491 = ~w13630 & ~w15490;
assign w15492 = ~w15422 & ~w15423;
assign w15493 = ~w14761 & ~w15492;
assign w15494 = w14567 & w41315;
assign w15495 = ~w14763 & w15494;
assign w15496 = ~w15493 & ~w15495;
assign w15497 = w14761 & ~w15491;
assign w15498 = ~w14765 & w15497;
assign w15499 = w15496 & ~w15498;
assign w15500 = (w41316 & w15441) | (w41316 & w44920) | (w15441 & w44920);
assign w15501 = ~w15499 & ~w15500;
assign w15502 = (w12666 & w15499) | (w12666 & w44921) | (w15499 & w44921);
assign w15503 = ~w15489 & ~w15502;
assign w15504 = ~w15489 & w41317;
assign w15505 = ~w15449 & w41318;
assign w15506 = ~w15504 & w15505;
assign w15507 = w14336 & ~w15383;
assign w15508 = ~w14336 & w15383;
assign w15509 = ~w15507 & ~w15508;
assign w15510 = ~w11138 & ~w15509;
assign w15511 = ~w10419 & ~w15510;
assign w15512 = w15347 & ~w15348;
assign w15513 = ~w15347 & w15348;
assign w15514 = ~w15512 & ~w15513;
assign w15515 = w9781 & w15340;
assign w15516 = w15514 & w15515;
assign w15517 = w15335 & ~w15516;
assign w15518 = w10419 & w15388;
assign w15519 = ~w15449 & w47447;
assign w15520 = ~w15504 & w15519;
assign w15521 = w14366 & ~w14379;
assign w15522 = ~w14336 & ~w15381;
assign w15523 = ~w15380 & ~w15522;
assign w15524 = w15521 & ~w15523;
assign w15525 = ~w15521 & w15523;
assign w15526 = ~w15524 & ~w15525;
assign w15527 = ~w14378 & w14766;
assign w15528 = ~w14766 & w15526;
assign w15529 = ~w15527 & ~w15528;
assign w15530 = w11976 & ~w15509;
assign w15531 = ~w15529 & ~w15530;
assign w15532 = w15517 & w15531;
assign w15533 = ~w15520 & w15532;
assign w15534 = w15511 & w15517;
assign w15535 = ~w15506 & w15534;
assign w15536 = ~w15533 & ~w15535;
assign w15537 = w15376 & w44922;
assign w15538 = w15536 & w15537;
assign w15539 = ~w15194 & w47448;
assign w15540 = ~w4838 & w15200;
assign w15541 = w15540 & w14766;
assign w15542 = (~w4838 & ~w15208) | (~w4838 & w41319) | (~w15208 & w41319);
assign w15543 = ~w14766 & w15542;
assign w15544 = ~w15541 & ~w15543;
assign w15545 = ~w14765 & w44923;
assign w15546 = ~w15176 & w49664;
assign w15547 = ~w14766 & w15546;
assign w15548 = ~w15545 & ~w15547;
assign w15549 = w15544 & w15548;
assign w15550 = ~w15539 & w15549;
assign w15551 = ~w15197 & ~w15550;
assign w15552 = ~w15220 & ~w15222;
assign w15553 = w5330 & w15223;
assign w15554 = w15552 & w15553;
assign w15555 = (~w5745 & w14765) | (~w5745 & w44924) | (w14765 & w44924);
assign w15556 = ~w15370 & w15555;
assign w15557 = w5330 & ~w15223;
assign w15558 = ~w14765 & w44925;
assign w15559 = ~w15219 & w15557;
assign w15560 = ~w14766 & w15559;
assign w15561 = ~w15558 & ~w15560;
assign w15562 = ~w15556 & w15561;
assign w15563 = ~w15554 & w15562;
assign w15564 = ~w15373 & w15563;
assign w15565 = ~w15307 & w48806;
assign w15566 = ~w15297 & ~w15565;
assign w15567 = w15296 & ~w15566;
assign w15568 = w15271 & w15563;
assign w15569 = ~w15567 & w15568;
assign w15570 = w15234 & ~w15564;
assign w15571 = ~w15569 & w15570;
assign w15572 = ~w15551 & ~w15571;
assign w15573 = w15058 & w15156;
assign w15574 = w15572 & w15573;
assign w15575 = ~w15538 & w15574;
assign w15576 = ~w15070 & ~w15072;
assign w15577 = ~w2285 & ~w15576;
assign w15578 = (~w15106 & ~w15100) | (~w15106 & w44926) | (~w15100 & w44926);
assign w15579 = w2558 & ~w15578;
assign w15580 = ~w15577 & ~w15579;
assign w15581 = w15087 & ~w15580;
assign w15582 = w3646 & ~w15152;
assign w15583 = ~w15142 & w15582;
assign w15584 = w15141 & ~w15583;
assign w15585 = w15125 & ~w15584;
assign w15586 = ~w15581 & ~w15585;
assign w15587 = ~w1738 & ~w15033;
assign w15588 = ~w15399 & ~w15402;
assign w15589 = w15033 & w15588;
assign w15590 = w14586 & ~w15589;
assign w15591 = w14241 & ~w15587;
assign w15592 = ~w15081 & w15591;
assign w15593 = ~w14241 & ~w15587;
assign w15594 = w15081 & w15593;
assign w15595 = ~w15592 & ~w15594;
assign w15596 = w15590 & w15595;
assign w15597 = ~w15033 & ~w14766;
assign w15598 = w14562 & ~w15597;
assign w15599 = w2006 & ~w15037;
assign w15600 = (~w1738 & w14766) | (~w1738 & w48807) | (w14766 & w48807);
assign w15601 = ~w15598 & w15600;
assign w15602 = w14562 & w15021;
assign w15603 = ~w1738 & ~w14241;
assign w15604 = w1738 & w14241;
assign w15605 = ~w2006 & ~w15604;
assign w15606 = ~w1738 & w14241;
assign w15607 = w1738 & ~w14241;
assign w15608 = ~w2006 & ~w15607;
assign w15609 = (w15588 & w44927) | (w15588 & w44928) | (w44927 & w44928);
assign w15610 = w15081 & w15609;
assign w15611 = (w15588 & w44929) | (w15588 & w44930) | (w44929 & w44930);
assign w15612 = ~w15081 & w15611;
assign w15613 = ~w15610 & ~w15612;
assign w15614 = w15049 & ~w15596;
assign w15615 = ~w15601 & w15613;
assign w15616 = w15614 & w15615;
assign w15617 = ~w15046 & ~w15616;
assign w15618 = ~w15058 & ~w15617;
assign w15619 = w15586 & ~w15617;
assign w15620 = ~w15618 & ~w15619;
assign w15621 = w14900 & ~w14966;
assign w15622 = w14982 & ~w15621;
assign w15623 = ~w15002 & w15009;
assign w15624 = ~w14995 & w15623;
assign w15625 = (~w14983 & w47449) | (~w14983 & w47450) | (w47449 & w47450);
assign w15626 = ~w15620 & w50198;
assign w15627 = w15015 & ~w15626;
assign w15628 = a[49] & ~w14766;
assign w15629 = ~a[49] & w14766;
assign w15630 = ~w15628 & ~w15629;
assign w15631 = ~w15468 & ~w15470;
assign w15632 = ~w15630 & ~w15631;
assign w15633 = w15630 & w15631;
assign w15634 = ~w15632 & ~w15633;
assign w15635 = ~a[48] & ~w15630;
assign w15636 = ~w15469 & ~w15635;
assign w15637 = ~w15626 & w48808;
assign w15638 = (w15636 & w15626) | (w15636 & w48809) | (w15626 & w48809);
assign w15639 = ~w15637 & ~w15638;
assign w15640 = ~w13384 & w15639;
assign w15641 = ~a[44] & ~a[45];
assign w15642 = ~a[46] & w15641;
assign w15643 = w14766 & ~w15642;
assign w15644 = ~w14777 & w50199;
assign w15645 = ~w14766 & w15642;
assign w15646 = ~a[47] & ~w15643;
assign w15647 = ~w15645 & ~w15646;
assign w15648 = ~w15234 & ~w15551;
assign w15649 = ~w15585 & w44932;
assign w15650 = w15388 & ~w15510;
assign w15651 = w15451 & ~w15504;
assign w15652 = (w15650 & w15504) | (w15650 & w44933) | (w15504 & w44933);
assign w15653 = w15518 & ~w15652;
assign w15654 = ~w15506 & w15511;
assign w15655 = (w15529 & w15506) | (w15529 & w44934) | (w15506 & w44934);
assign w15656 = ~w15653 & ~w15655;
assign w15657 = w15378 & w15649;
assign w15658 = ~w15656 & w15657;
assign w15659 = ~w15564 & ~w15569;
assign w15660 = (~w15551 & w15569) | (~w15551 & w44935) | (w15569 & w44935);
assign w15661 = w15311 & w15375;
assign w15662 = (w15233 & w15516) | (w15233 & w44936) | (w15516 & w44936);
assign w15663 = w15661 & w15662;
assign w15664 = w15660 & ~w15663;
assign w15665 = w15649 & ~w15664;
assign w15666 = ~w15658 & ~w15665;
assign w15667 = ~w15617 & w47451;
assign w15668 = ~w15156 & ~w15581;
assign w15669 = (~w14777 & w15156) | (~w14777 & w44937) | (w15156 & w44937);
assign w15670 = ~w15667 & w15669;
assign w15671 = ~w15014 & w15670;
assign w15672 = w15666 & w15671;
assign w15673 = w15058 & ~w15616;
assign w15674 = w15622 & ~w15673;
assign w15675 = ~w14777 & w14832;
assign w15676 = w14973 & w15675;
assign w15677 = ~w15674 & w15676;
assign w15678 = ~w14983 & w15624;
assign w15679 = (~w14777 & w14983) | (~w14777 & w47452) | (w14983 & w47452);
assign w15680 = ~w15677 & ~w15679;
assign w15681 = ~w15672 & w15680;
assign w15682 = ~a[47] & ~w15645;
assign w15683 = (w15682 & w15672) | (w15682 & w47453) | (w15672 & w47453);
assign w15684 = (w15647 & w15626) | (w15647 & w48811) | (w15626 & w48811);
assign w15685 = ~w15683 & ~w15684;
assign w15686 = ~w15683 & w48812;
assign w15687 = a[46] & ~a[47];
assign w15688 = (w15672 & w48813) | (w15672 & w48814) | (w48813 & w48814);
assign w15689 = a[48] & ~w14766;
assign w15690 = ~a[48] & w14766;
assign w15691 = ~w15689 & ~w15690;
assign w15692 = a[48] & ~w15466;
assign w15693 = ~w15672 & w47455;
assign w15694 = ~w15467 & ~w15692;
assign w15695 = (w15694 & w15672) | (w15694 & w47456) | (w15672 & w47456);
assign w15696 = ~w15693 & ~w15695;
assign w15697 = ~w15688 & w15696;
assign w15698 = ~w15686 & w15697;
assign w15699 = ~w14039 & w50200;
assign w15700 = ~w15685 & w15699;
assign w15701 = w13384 & ~w15639;
assign w15702 = ~w15700 & ~w15701;
assign w15703 = ~w15698 & w15702;
assign w15704 = ~w15640 & ~w15703;
assign w15705 = ~w13384 & w15482;
assign w15706 = w13384 & ~w15482;
assign w15707 = ~w15705 & ~w15706;
assign w15708 = ~w15672 & w48815;
assign w15709 = w15487 & w15707;
assign w15710 = ~w15487 & ~w15707;
assign w15711 = ~w15709 & ~w15710;
assign w15712 = w15487 & w15708;
assign w15713 = ~w15708 & w15711;
assign w15714 = ~w15712 & ~w15713;
assign w15715 = ~w12666 & w15714;
assign w15716 = w12666 & ~w15489;
assign w15717 = ~w12666 & w15489;
assign w15718 = ~w15716 & ~w15717;
assign w15719 = ~w15501 & ~w15718;
assign w15720 = w15501 & w15718;
assign w15721 = ~w15719 & ~w15720;
assign w15722 = ~w15677 & w44938;
assign w15723 = (w15721 & w15672) | (w15721 & w47457) | (w15672 & w47457);
assign w15724 = ~w15677 & w44939;
assign w15725 = (~w11870 & w15672) | (~w11870 & w47458) | (w15672 & w47458);
assign w15726 = ~w15723 & w15725;
assign w15727 = ~w15715 & ~w15726;
assign w15728 = ~w15704 & w15727;
assign w15729 = w12666 & w15711;
assign w15730 = ~w15677 & w44940;
assign w15731 = (w15729 & w15672) | (w15729 & w47459) | (w15672 & w47459);
assign w15732 = w12666 & w15709;
assign w15733 = ~w15672 & w47460;
assign w15734 = ~w15731 & ~w15733;
assign w15735 = ~w15672 & w47461;
assign w15736 = ~w15723 & ~w15735;
assign w15737 = ~w15726 & ~w15734;
assign w15738 = w11870 & ~w15736;
assign w15739 = ~w15737 & ~w15738;
assign w15740 = ~w15653 & ~w15654;
assign w15741 = w9781 & ~w15529;
assign w15742 = w15740 & w15741;
assign w15743 = (w15742 & w15672) | (w15742 & w47462) | (w15672 & w47462);
assign w15744 = w9781 & w15529;
assign w15745 = ~w15740 & w15744;
assign w15746 = ~w15677 & w44941;
assign w15747 = (~w15745 & w15672) | (~w15745 & w47463) | (w15672 & w47463);
assign w15748 = ~w15650 & w15651;
assign w15749 = ~w15652 & ~w15748;
assign w15750 = w10419 & ~w15509;
assign w15751 = ~w15672 & w47464;
assign w15752 = w10419 & ~w15749;
assign w15753 = (w15752 & w15672) | (w15752 & w47465) | (w15672 & w47465);
assign w15754 = ~w15751 & ~w15753;
assign w15755 = ~w15743 & w15747;
assign w15756 = w15754 & w15755;
assign w15757 = w15446 & ~w15503;
assign w15758 = w11870 & ~w15757;
assign w15759 = ~w11870 & w15757;
assign w15760 = ~w15758 & ~w15759;
assign w15761 = ~w15677 & w44942;
assign w15762 = ~w15448 & ~w15760;
assign w15763 = w15448 & w15760;
assign w15764 = ~w15762 & ~w15763;
assign w15765 = (w15764 & w15672) | (w15764 & w47466) | (w15672 & w47466);
assign w15766 = ~w15677 & w44943;
assign w15767 = ~w15672 & w15766;
assign w15768 = (~w11138 & w15672) | (~w11138 & w47467) | (w15672 & w47467);
assign w15769 = ~w15765 & w15768;
assign w15770 = ~w10419 & w15509;
assign w15771 = ~w15672 & w47468;
assign w15772 = ~w10419 & w15749;
assign w15773 = (w15772 & w15672) | (w15772 & w47469) | (w15672 & w47469);
assign w15774 = ~w15771 & ~w15773;
assign w15775 = w15769 & w15774;
assign w15776 = w15756 & ~w15775;
assign w15777 = w15739 & w15776;
assign w15778 = ~w15672 & w47470;
assign w15779 = w11138 & w15764;
assign w15780 = (w15779 & w15672) | (w15779 & w47471) | (w15672 & w47471);
assign w15781 = ~w15778 & ~w15780;
assign w15782 = w15774 & w15781;
assign w15783 = w15756 & ~w15782;
assign w15784 = w9781 & ~w15656;
assign w15785 = ~w9781 & w15656;
assign w15786 = ~w15784 & ~w15785;
assign w15787 = ~w15514 & ~w15786;
assign w15788 = ~w15677 & w44944;
assign w15789 = (~w15787 & w15672) | (~w15787 & w47472) | (w15672 & w47472);
assign w15790 = w14974 & ~w15674;
assign w15791 = (w15678 & w15674) | (w15678 & w44945) | (w15674 & w44945);
assign w15792 = ~w15649 & ~w15668;
assign w15793 = w15378 & ~w15656;
assign w15794 = ~w15663 & ~w15668;
assign w15795 = w15660 & w15794;
assign w15796 = ~w15793 & w15795;
assign w15797 = ~w15792 & ~w15796;
assign w15798 = (~w14995 & w14982) | (~w14995 & w47473) | (w14982 & w47473);
assign w15799 = ~w14974 & w15798;
assign w15800 = ~w15618 & ~w15799;
assign w15801 = ~w14777 & w15514;
assign w15802 = w15786 & w15801;
assign w15803 = w15625 & ~w15800;
assign w15804 = w15802 & ~w15803;
assign w15805 = w15791 & w15797;
assign w15806 = w15804 & ~w15805;
assign w15807 = w15789 & ~w15806;
assign w15808 = w9195 & ~w15807;
assign w15809 = (w15740 & w15672) | (w15740 & w47474) | (w15672 & w47474);
assign w15810 = ~w9781 & ~w15529;
assign w15811 = ~w15809 & w15810;
assign w15812 = ~w9781 & w15529;
assign w15813 = w15809 & w15812;
assign w15814 = ~w15811 & ~w15813;
assign w15815 = ~w15808 & w15814;
assign w15816 = ~w15783 & w15815;
assign w15817 = (~w15374 & w15354) | (~w15374 & w44946) | (w15354 & w44946);
assign w15818 = (w7924 & ~w15536) | (w7924 & w48816) | (~w15536 & w48816);
assign w15819 = w15536 & w48817;
assign w15820 = ~w15818 & ~w15819;
assign w15821 = (~w15820 & w15672) | (~w15820 & w47475) | (w15672 & w47475);
assign w15822 = w15308 & ~w15821;
assign w15823 = ~w15308 & w15821;
assign w15824 = ~w15822 & ~w15823;
assign w15825 = w7315 & ~w15824;
assign w15826 = ~w15309 & w15817;
assign w15827 = (~w15565 & ~w41324) | (~w15565 & w48818) | (~w41324 & w48818);
assign w15828 = w15292 & ~w15827;
assign w15829 = (w15828 & w15672) | (w15828 & w47476) | (w15672 & w47476);
assign w15830 = ~w15672 & w47477;
assign w15831 = w15233 & ~w15564;
assign w15832 = ~w15569 & w15831;
assign w15833 = w44947 & w47478;
assign w15834 = ~w15658 & w15833;
assign w15835 = ~w15197 & w15586;
assign w15836 = ~w15673 & w15835;
assign w15837 = w15668 & ~w15673;
assign w15838 = (w15566 & ~w41324) | (w15566 & w48819) | (~w41324 & w48819);
assign w15839 = w7315 & ~w14777;
assign w15840 = w15291 & ~w15839;
assign w15841 = w15838 & ~w15840;
assign w15842 = w15058 & ~w15837;
assign w15843 = ~w15799 & w15842;
assign w15844 = w15841 & w15843;
assign w15845 = (w15836 & w15658) | (w15836 & w48820) | (w15658 & w48820);
assign w15846 = w15844 & ~w15845;
assign w15847 = w7315 & w15625;
assign w15848 = w15841 & ~w15847;
assign w15849 = w15297 & ~w15827;
assign w15850 = ~w15848 & ~w15849;
assign w15851 = ~w15829 & ~w15830;
assign w15852 = ~w15846 & w15850;
assign w15853 = w15851 & w15852;
assign w15854 = (~w6769 & ~w15851) | (~w6769 & w48821) | (~w15851 & w48821);
assign w15855 = ~w15825 & ~w15854;
assign w15856 = w9781 & w15514;
assign w15857 = (w15353 & ~w15656) | (w15353 & w48822) | (~w15656 & w48822);
assign w15858 = ~w15334 & ~w15374;
assign w15859 = w15340 & ~w15858;
assign w15860 = ~w15340 & w15858;
assign w15861 = ~w15859 & ~w15860;
assign w15862 = w15323 & ~w15858;
assign w15863 = ~w15323 & w15858;
assign w15864 = ~w15862 & ~w15863;
assign w15865 = w15857 & ~w15861;
assign w15866 = ~w15857 & ~w15864;
assign w15867 = ~w15865 & ~w15866;
assign w15868 = ~w15672 & w47479;
assign w15869 = (~w15867 & w15672) | (~w15867 & w48823) | (w15672 & w48823);
assign w15870 = ~w15868 & ~w15869;
assign w15871 = (w7924 & w15869) | (w7924 & w47480) | (w15869 & w47480);
assign w15872 = ~w9195 & w15857;
assign w15873 = w9195 & ~w15857;
assign w15874 = ~w15872 & ~w15873;
assign w15875 = ~w15681 & w15874;
assign w15876 = ~w8666 & w15322;
assign w15877 = (w15876 & w15681) | (w15876 & w47481) | (w15681 & w47481);
assign w15878 = ~w8666 & ~w15322;
assign w15879 = ~w15681 & w47482;
assign w15880 = ~w15877 & ~w15879;
assign w15881 = ~w7315 & ~w15308;
assign w15882 = ~w15821 & w15881;
assign w15883 = ~w7315 & w15308;
assign w15884 = w15821 & w15883;
assign w15885 = ~w15882 & ~w15884;
assign w15886 = ~w15869 & w47483;
assign w15887 = w15885 & ~w15886;
assign w15888 = ~w15871 & ~w15880;
assign w15889 = w15887 & ~w15888;
assign w15890 = w15855 & ~w15889;
assign w15891 = w6769 & w15853;
assign w15892 = w15255 & ~w15295;
assign w15893 = ~w15292 & ~w15838;
assign w15894 = w15892 & ~w15893;
assign w15895 = ~w15892 & w15893;
assign w15896 = ~w15894 & ~w15895;
assign w15897 = ~w15243 & ~w15293;
assign w15898 = w15681 & w15897;
assign w15899 = ~w15681 & w15896;
assign w15900 = ~w15898 & ~w15899;
assign w15901 = ~w6264 & ~w15900;
assign w15902 = ~w15891 & ~w15901;
assign w15903 = ~w15890 & w15902;
assign w15904 = ~w15890 & w48824;
assign w15905 = (w15777 & w15704) | (w15777 & w48825) | (w15704 & w48825);
assign w15906 = w15904 & ~w15905;
assign w15907 = ~w9195 & w15807;
assign w15908 = w8666 & ~w15322;
assign w15909 = (w15908 & w15681) | (w15908 & w47484) | (w15681 & w47484);
assign w15910 = w8666 & w15322;
assign w15911 = ~w15681 & w47485;
assign w15912 = ~w15909 & ~w15911;
assign w15913 = ~w15907 & w15912;
assign w15914 = ~w15825 & w48826;
assign w15915 = w15913 & w15914;
assign w15916 = w15903 & ~w15915;
assign w15917 = ~w15360 & ~w15681;
assign w15918 = w15270 & ~w15917;
assign w15919 = w15296 & ~w15838;
assign w15920 = w15255 & ~w15919;
assign w15921 = w15271 & ~w15567;
assign w15922 = w41324 & w44948;
assign w15923 = w15921 & ~w15922;
assign w15924 = ~w15681 & ~w15923;
assign w15925 = w15264 & w15265;
assign w15926 = ~w15264 & ~w15265;
assign w15927 = ~w15925 & ~w15926;
assign w15928 = ~w15924 & w15927;
assign w15929 = w6264 & w15923;
assign w15930 = w15627 & w15929;
assign w15931 = ~w15928 & ~w15930;
assign w15932 = ~w15918 & ~w15920;
assign w15933 = w15931 & ~w15932;
assign w15934 = ~w5745 & ~w15933;
assign w15935 = w6264 & w15900;
assign w15936 = ~w15934 & ~w15935;
assign w15937 = ~w15916 & w15936;
assign w15938 = ~w15906 & w15937;
assign w15939 = w5745 & w15933;
assign w15940 = ~w15625 & ~w15799;
assign w15941 = ~w14777 & w15940;
assign w15942 = w15046 & w15623;
assign w15943 = ~w15941 & w15942;
assign w15944 = (w15539 & ~w15666) | (w15539 & w48827) | (~w15666 & w48827);
assign w15945 = w15943 & w15944;
assign w15946 = w15376 & w44949;
assign w15947 = (w15183 & ~w44947) | (w15183 & w47486) | (~w44947 & w47486);
assign w15948 = w15183 & w15946;
assign w15949 = ~w15656 & w15948;
assign w15950 = ~w15947 & ~w15949;
assign w15951 = ~w4056 & w15549;
assign w15952 = (~w15186 & ~w44950) | (~w15186 & w47487) | (~w44950 & w47487);
assign w15953 = ~w15186 & w15946;
assign w15954 = ~w15656 & w15953;
assign w15955 = ~w15952 & ~w15954;
assign w15956 = w15950 & ~w15955;
assign w15957 = ~w15195 & ~w15956;
assign w15958 = ~w15677 & w44951;
assign w15959 = ~w15672 & w15958;
assign w15960 = ~w15957 & ~w15959;
assign w15961 = (w15196 & ~w44950) | (w15196 & w47488) | (~w44950 & w47488);
assign w15962 = w15196 & w15946;
assign w15963 = ~w15656 & w15962;
assign w15964 = ~w15961 & ~w15963;
assign w15965 = w15950 & ~w15964;
assign w15966 = ~w3646 & ~w15965;
assign w15967 = ~w15677 & w44952;
assign w15968 = ~w15672 & w15967;
assign w15969 = ~w15966 & ~w15968;
assign w15970 = w15944 & w47489;
assign w15971 = w15960 & ~w15969;
assign w15972 = ~w15970 & ~w15971;
assign w15973 = ~w15178 & ~w15180;
assign w15974 = w4056 & ~w15973;
assign w15975 = w15681 & ~w15974;
assign w15976 = w41325 & w44953;
assign w15977 = w15232 & w15659;
assign w15978 = w15544 & ~w15977;
assign w15979 = ~w15976 & w15978;
assign w15980 = ~w15217 & ~w15979;
assign w15981 = ~w15182 & w15548;
assign w15982 = w15183 & w15548;
assign w15983 = ~w15980 & w15982;
assign w15984 = w4056 & ~w15981;
assign w15985 = w15980 & w15984;
assign w15986 = ~w15681 & w47490;
assign w15987 = ~w15975 & ~w15986;
assign w15988 = w15972 & ~w15987;
assign w15989 = ~w15217 & w15544;
assign w15990 = ~w15976 & ~w15977;
assign w15991 = w15989 & ~w15990;
assign w15992 = ~w15989 & w15990;
assign w15993 = ~w15991 & ~w15992;
assign w15994 = ~w15216 & w15681;
assign w15995 = ~w15681 & w15993;
assign w15996 = ~w15994 & ~w15995;
assign w15997 = ~w4430 & w15996;
assign w15998 = ~w15672 & w47491;
assign w15999 = (w15980 & w15672) | (w15980 & w47492) | (w15672 & w47492);
assign w16000 = ~w15998 & ~w15999;
assign w16001 = ~w4056 & ~w15981;
assign w16002 = w16000 & w16001;
assign w16003 = ~w4056 & w15981;
assign w16004 = ~w16000 & w16003;
assign w16005 = ~w16002 & ~w16004;
assign w16006 = ~w15997 & w16005;
assign w16007 = w4430 & ~w15996;
assign w16008 = (w15373 & w15567) | (w15373 & w47493) | (w15567 & w47493);
assign w16009 = ~w15556 & ~w16008;
assign w16010 = (w16009 & ~w41325) | (w16009 & w44954) | (~w41325 & w44954);
assign w16011 = w5330 & ~w16010;
assign w16012 = ~w5330 & w16010;
assign w16013 = ~w16011 & ~w16012;
assign w16014 = w15223 & ~w15552;
assign w16015 = ~w15223 & w15552;
assign w16016 = ~w16014 & ~w16015;
assign w16017 = w16013 & ~w16016;
assign w16018 = ~w15681 & w16017;
assign w16019 = (~w5330 & ~w15666) | (~w5330 & w48828) | (~w15666 & w48828);
assign w16020 = w15943 & w16019;
assign w16021 = w16018 & ~w16020;
assign w16022 = ~w16013 & w16016;
assign w16023 = ~w15677 & w44955;
assign w16024 = ~w15672 & w16023;
assign w16025 = ~w16022 & ~w16024;
assign w16026 = ~w16021 & w16025;
assign w16027 = (~w4838 & w16021) | (~w4838 & w47494) | (w16021 & w47494);
assign w16028 = ~w16007 & ~w16027;
assign w16029 = ~w15672 & w47495;
assign w16030 = ~w15372 & ~w15556;
assign w16031 = w15360 & ~w15923;
assign w16032 = ~w16030 & w16031;
assign w16033 = ~w15681 & ~w16032;
assign w16034 = w16030 & ~w16031;
assign w16035 = ~w5330 & w16029;
assign w16036 = ~w5330 & ~w16034;
assign w16037 = w16033 & w16036;
assign w16038 = ~w16035 & ~w16037;
assign w16039 = ~w16024 & w47496;
assign w16040 = ~w16021 & w16039;
assign w16041 = w16038 & ~w16040;
assign w16042 = w15988 & ~w16006;
assign w16043 = w15988 & ~w16041;
assign w16044 = w16028 & w16043;
assign w16045 = ~w16042 & ~w16044;
assign w16046 = w15123 & ~w15584;
assign w16047 = ~w15108 & ~w15579;
assign w16048 = w16046 & ~w16047;
assign w16049 = ~w16046 & w16047;
assign w16050 = ~w16048 & ~w16049;
assign w16051 = ~w15140 & ~w15142;
assign w16052 = ~w15582 & w16051;
assign w16053 = w15123 & ~w15128;
assign w16054 = ~w15140 & ~w15154;
assign w16055 = w16052 & ~w16054;
assign w16056 = w16053 & w16055;
assign w16057 = w15572 & w50201;
assign w16058 = w16050 & ~w16057;
assign w16059 = ~w16050 & w16057;
assign w16060 = ~w16058 & ~w16059;
assign w16061 = ~w15672 & w48829;
assign w16062 = ~w15681 & ~w16060;
assign w16063 = ~w16061 & ~w16062;
assign w16064 = (w2285 & w16062) | (w2285 & w48830) | (w16062 & w48830);
assign w16065 = ~w15109 & ~w15126;
assign w16066 = ~w15677 & w44957;
assign w16067 = ~w15672 & w16066;
assign w16068 = ~w15153 & w16052;
assign w16069 = ~w15648 & w16068;
assign w16070 = ~w15664 & w16069;
assign w16071 = w15378 & w16069;
assign w16072 = ~w15656 & w16071;
assign w16073 = ~w16070 & ~w16072;
assign w16074 = w16053 & ~w16054;
assign w16075 = ~w16053 & w16054;
assign w16076 = ~w16074 & ~w16075;
assign w16077 = w16073 & ~w16076;
assign w16078 = ~w16073 & w16076;
assign w16079 = ~w16077 & ~w16078;
assign w16080 = ~w15681 & ~w16079;
assign w16081 = ~w16067 & ~w16080;
assign w16082 = (~w2558 & w16080) | (~w2558 & w48831) | (w16080 & w48831);
assign w16083 = ~w16064 & ~w16082;
assign w16084 = w15582 & ~w16051;
assign w16085 = ~w16052 & ~w16084;
assign w16086 = ~w15153 & ~w15582;
assign w16087 = w15572 & w16086;
assign w16088 = ~w15538 & w16087;
assign w16089 = (w16085 & w15538) | (w16085 & w41327) | (w15538 & w41327);
assign w16090 = ~w15538 & w41328;
assign w16091 = ~w16089 & ~w16090;
assign w16092 = ~w2896 & ~w15139;
assign w16093 = ~w15672 & w48832;
assign w16094 = ~w2896 & w16091;
assign w16095 = ~w15681 & w16094;
assign w16096 = ~w16093 & ~w16095;
assign w16097 = (w2558 & w15672) | (w2558 & w48833) | (w15672 & w48833);
assign w16098 = ~w16080 & w16097;
assign w16099 = w16096 & ~w16098;
assign w16100 = (w15965 & w15672) | (w15965 & w48834) | (w15672 & w48834);
assign w16101 = w15960 & ~w16100;
assign w16102 = w3646 & ~w15945;
assign w16103 = ~w16101 & w16102;
assign w16104 = (~w41326 & w44958) | (~w41326 & w44959) | (w44958 & w44959);
assign w16105 = ~w16088 & ~w16104;
assign w16106 = ~w15672 & w48835;
assign w16107 = (w16105 & w15672) | (w16105 & w48836) | (w15672 & w48836);
assign w16108 = ~w16106 & ~w16107;
assign w16109 = w3242 & ~w16108;
assign w16110 = ~w2285 & w16063;
assign w16111 = ~w16103 & ~w16109;
assign w16112 = ~w16110 & w16111;
assign w16113 = w16083 & ~w16099;
assign w16114 = w16112 & ~w16113;
assign w16115 = w16045 & w16114;
assign w16116 = w16045 & w47497;
assign w16117 = ~w15938 & w16116;
assign w16118 = ~w15044 & ~w15048;
assign w16119 = ~w15596 & w15615;
assign w16120 = ~w2006 & ~w14241;
assign w16121 = ~w15081 & w16120;
assign w16122 = ~w2006 & w14241;
assign w16123 = w15081 & w16122;
assign w16124 = ~w16121 & ~w16123;
assign w16125 = ~w15056 & ~w16124;
assign w16126 = ~w15056 & ~w15074;
assign w16127 = w15086 & w16126;
assign w16128 = ~w16125 & ~w16127;
assign w16129 = w16119 & w16128;
assign w16130 = w15124 & w15154;
assign w16131 = w15124 & ~w15584;
assign w16132 = (w15580 & w15584) | (w15580 & w44960) | (w15584 & w44960);
assign w16133 = w16119 & w16132;
assign w16134 = w15648 & w16130;
assign w16135 = w16133 & ~w16134;
assign w16136 = ~w16129 & ~w16135;
assign w16137 = ~w16129 & w16130;
assign w16138 = ~w15663 & w16137;
assign w16139 = w15660 & w16138;
assign w16140 = ~w15793 & w16139;
assign w16141 = ~w16118 & ~w16136;
assign w16142 = ~w16140 & w16141;
assign w16143 = w16118 & w16136;
assign w16144 = w16138 & w48837;
assign w16145 = ~w15793 & w16144;
assign w16146 = ~w16143 & ~w16145;
assign w16147 = ~w15672 & w48838;
assign w16148 = ~w16142 & w16146;
assign w16149 = ~w15681 & w16148;
assign w16150 = ~w16147 & ~w16149;
assign w16151 = ~w16149 & w48839;
assign w16152 = ~w15051 & ~w15054;
assign w16153 = (~w16152 & w15672) | (~w16152 & w48840) | (w15672 & w48840);
assign w16154 = ~w15156 & w44961;
assign w16155 = ~w15648 & w16124;
assign w16156 = w15586 & w16155;
assign w16157 = ~w16154 & ~w16156;
assign w16158 = w1738 & w16157;
assign w16159 = w15794 & w44962;
assign w16160 = ~w15793 & w16159;
assign w16161 = ~w16158 & ~w16160;
assign w16162 = (~w1738 & w16156) | (~w1738 & w44963) | (w16156 & w44963);
assign w16163 = w15793 & w16162;
assign w16164 = ~w15795 & ~w16157;
assign w16165 = ~w1738 & w16164;
assign w16166 = ~w16163 & ~w16165;
assign w16167 = w16161 & w16166;
assign w16168 = w16153 & ~w16167;
assign w16169 = ~w1738 & w16152;
assign w16170 = w16157 & ~w16169;
assign w16171 = w15794 & w44964;
assign w16172 = ~w15793 & w16171;
assign w16173 = ~w16170 & ~w16172;
assign w16174 = ~w15056 & ~w16157;
assign w16175 = ~w15796 & w16174;
assign w16176 = w16173 & ~w16175;
assign w16177 = ~w15677 & w44965;
assign w16178 = ~w15672 & w16177;
assign w16179 = ~w16176 & ~w16178;
assign w16180 = ~w16178 & w48841;
assign w16181 = ~w16168 & w16180;
assign w16182 = (~w16142 & w15672) | (~w16142 & w48842) | (w15672 & w48842);
assign w16183 = ~w1320 & w16147;
assign w16184 = ~w1320 & w16146;
assign w16185 = w16182 & w16184;
assign w16186 = ~w16183 & ~w16185;
assign w16187 = ~w16181 & w16186;
assign w16188 = ~w16151 & ~w16187;
assign w16189 = (w41323 & w44966) | (w41323 & w44967) | (w44966 & w44967);
assign w16190 = (~w41323 & w44968) | (~w41323 & w44969) | (w44968 & w44969);
assign w16191 = ~w16189 & ~w16190;
assign w16192 = (w14968 & w15672) | (w14968 & w48843) | (w15672 & w48843);
assign w16193 = (~w41323 & w44970) | (~w41323 & w44971) | (w44970 & w44971);
assign w16194 = ~w1120 & ~w14968;
assign w16195 = (w41323 & w44972) | (w41323 & w44973) | (w44972 & w44973);
assign w16196 = ~w16193 & ~w16195;
assign w16197 = ~w15677 & w44974;
assign w16198 = ~w15672 & w16197;
assign w16199 = w16196 & ~w16198;
assign w16200 = (w945 & w16198) | (w945 & w48844) | (w16198 & w48844);
assign w16201 = w945 & w16191;
assign w16202 = w16192 & w16201;
assign w16203 = ~w16200 & ~w16202;
assign w16204 = ~w15663 & w16130;
assign w16205 = w15660 & w16204;
assign w16206 = ~w15048 & w16135;
assign w16207 = ~w15048 & w16129;
assign w16208 = ~w15044 & ~w16207;
assign w16209 = ~w16206 & w16208;
assign w16210 = w16205 & w16208;
assign w16211 = ~w15793 & w16210;
assign w16212 = ~w16209 & ~w16211;
assign w16213 = ~w15031 & ~w15032;
assign w16214 = w1120 & ~w16213;
assign w16215 = ~w1320 & w16214;
assign w16216 = ~w15672 & w48845;
assign w16217 = (w16214 & w16211) | (w16214 & w48846) | (w16211 & w48846);
assign w16218 = ~w15681 & w16217;
assign w16219 = ~w16216 & ~w16218;
assign w16220 = w1120 & w16213;
assign w16221 = ~w16211 & w48847;
assign w16222 = ~w15681 & w16221;
assign w16223 = w1320 & w16220;
assign w16224 = ~w15672 & w48848;
assign w16225 = ~w16222 & ~w16224;
assign w16226 = w16219 & w16225;
assign w16227 = w16203 & w16226;
assign w16228 = (w1541 & w16178) | (w1541 & w48849) | (w16178 & w48849);
assign w16229 = (w1541 & ~w16166) | (w1541 & w44975) | (~w16166 & w44975);
assign w16230 = w16153 & w16229;
assign w16231 = ~w16228 & ~w16230;
assign w16232 = ~w16151 & w16231;
assign w16233 = w16191 & w16192;
assign w16234 = w16199 & ~w16233;
assign w16235 = ~w15672 & w48850;
assign w16236 = ~w15681 & ~w16212;
assign w16237 = ~w16235 & ~w16236;
assign w16238 = ~w1120 & w16213;
assign w16239 = (w16238 & w16236) | (w16238 & w48851) | (w16236 & w48851);
assign w16240 = ~w1120 & ~w16213;
assign w16241 = ~w16236 & w48852;
assign w16242 = ~w16239 & ~w16241;
assign w16243 = ~w945 & w16234;
assign w16244 = w16242 & ~w16243;
assign w16245 = w16203 & ~w16244;
assign w16246 = w16227 & ~w16232;
assign w16247 = ~w16188 & w16246;
assign w16248 = ~w16245 & ~w16247;
assign w16249 = w5330 & ~w16029;
assign w16250 = ~w15681 & w48853;
assign w16251 = w16249 & ~w16250;
assign w16252 = ~w16040 & w16251;
assign w16253 = w15988 & ~w16252;
assign w16254 = w16028 & w16253;
assign w16255 = w16114 & ~w16254;
assign w16256 = w16045 & w16255;
assign w16257 = ~w14241 & ~w15081;
assign w16258 = w14241 & w15081;
assign w16259 = ~w16257 & ~w16258;
assign w16260 = ~w15672 & w48854;
assign w16261 = ~w15571 & w44976;
assign w16262 = ~w15074 & w16132;
assign w16263 = (w16262 & w15538) | (w16262 & w41329) | (w15538 & w41329);
assign w16264 = ~w15074 & ~w16263;
assign w16265 = w15086 & w16124;
assign w16266 = ~w16264 & ~w16265;
assign w16267 = w16264 & w16265;
assign w16268 = ~w15681 & w48855;
assign w16269 = ~w16260 & ~w16268;
assign w16270 = ~w1738 & ~w16269;
assign w16271 = w1738 & ~w16260;
assign w16272 = ~w16268 & w16271;
assign w16273 = ~w15579 & ~w16131;
assign w16274 = ~w15074 & ~w15577;
assign w16275 = (w16273 & w15538) | (w16273 & w41330) | (w15538 & w41330);
assign w16276 = ~w16274 & ~w16275;
assign w16277 = ~w15672 & w48856;
assign w16278 = ~w16263 & ~w16276;
assign w16279 = ~w15681 & w16278;
assign w16280 = ~w16277 & ~w16279;
assign w16281 = w2006 & ~w16280;
assign w16282 = ~w16272 & ~w16281;
assign w16283 = ~w16270 & ~w16282;
assign w16284 = ~w3242 & w15152;
assign w16285 = ~w15672 & w48857;
assign w16286 = ~w3242 & ~w16105;
assign w16287 = ~w15681 & w16286;
assign w16288 = ~w16285 & ~w16287;
assign w16289 = w2896 & w15139;
assign w16290 = ~w15672 & w48858;
assign w16291 = w2896 & ~w16091;
assign w16292 = ~w15681 & w16291;
assign w16293 = ~w16290 & ~w16292;
assign w16294 = w16288 & w16293;
assign w16295 = w16099 & ~w16294;
assign w16296 = (~w16110 & w16295) | (~w16110 & w48859) | (w16295 & w48859);
assign w16297 = ~w16283 & ~w16296;
assign w16298 = w16248 & w16297;
assign w16299 = ~w16256 & w16298;
assign w16300 = ~w16117 & w16299;
assign w16301 = ~w15672 & w47498;
assign w16302 = (w14966 & w15619) | (w14966 & w44977) | (w15619 & w44977);
assign w16303 = ~w14882 & ~w14972;
assign w16304 = (w16303 & w15575) | (w16303 & w41331) | (w15575 & w41331);
assign w16305 = ~w14882 & ~w16304;
assign w16306 = ~w15681 & ~w16305;
assign w16307 = ~w14957 & w14964;
assign w16308 = ~w14882 & ~w14958;
assign w16309 = ~w16307 & ~w16308;
assign w16310 = w14971 & ~w16308;
assign w16311 = (~w41323 & w44978) | (~w41323 & w44979) | (w44978 & w44979);
assign w16312 = ~w16309 & ~w16311;
assign w16313 = w493 & w16301;
assign w16314 = w493 & w16312;
assign w16315 = w16306 & w16314;
assign w16316 = ~w16313 & ~w16315;
assign w16317 = w14936 & ~w14970;
assign w16318 = w754 & w16317;
assign w16319 = (w16318 & w15617) | (w16318 & w47499) | (w15617 & w47499);
assign w16320 = w15792 & w16319;
assign w16321 = w15795 & w16319;
assign w16322 = (~w16320 & ~w16321) | (~w16320 & w44980) | (~w16321 & w44980);
assign w16323 = ~w14926 & w14936;
assign w16324 = ~w754 & ~w16323;
assign w16325 = w15836 & w16324;
assign w16326 = ~w15834 & w16325;
assign w16327 = (w16317 & w15617) | (w16317 & w47500) | (w15617 & w47500);
assign w16328 = ~w15837 & w16327;
assign w16329 = w16324 & ~w16328;
assign w16330 = w14926 & ~w15617;
assign w16331 = w16318 & ~w16330;
assign w16332 = ~w16329 & ~w16331;
assign w16333 = ~w16326 & w16332;
assign w16334 = w16322 & w16333;
assign w16335 = w14946 & ~w14959;
assign w16336 = ~w14946 & w14959;
assign w16337 = ~w16335 & ~w16336;
assign w16338 = w612 & ~w16337;
assign w16339 = (w16338 & w15672) | (w16338 & w47501) | (w15672 & w47501);
assign w16340 = ~w16334 & w16339;
assign w16341 = w612 & w16337;
assign w16342 = ~w15672 & w47502;
assign w16343 = w16341 & w16322;
assign w16344 = w16333 & w16343;
assign w16345 = ~w16342 & ~w16344;
assign w16346 = ~w16340 & w16345;
assign w16347 = w16316 & w16346;
assign w16348 = ~w612 & w16337;
assign w16349 = (w16348 & w15672) | (w16348 & w47503) | (w15672 & w47503);
assign w16350 = ~w16334 & w16349;
assign w16351 = ~w612 & ~w16337;
assign w16352 = ~w15672 & w47504;
assign w16353 = w16351 & w16322;
assign w16354 = w16333 & w16353;
assign w16355 = ~w16352 & ~w16354;
assign w16356 = ~w16350 & w16355;
assign w16357 = w14914 & w14936;
assign w16358 = (~w14969 & w15575) | (~w14969 & w41332) | (w15575 & w41332);
assign w16359 = w16357 & ~w16358;
assign w16360 = ~w16357 & w16358;
assign w16361 = ~w15681 & w47505;
assign w16362 = ~w945 & w14936;
assign w16363 = w14914 & ~w16362;
assign w16364 = ~w15672 & w47506;
assign w16365 = ~w754 & ~w16364;
assign w16366 = ~w16361 & w16365;
assign w16367 = w16356 & ~w16366;
assign w16368 = w16347 & ~w16367;
assign w16369 = ~w15681 & w47507;
assign w16370 = ~w16301 & ~w16369;
assign w16371 = ~w493 & w16370;
assign w16372 = ~w14898 & ~w14976;
assign w16373 = w16304 & ~w16372;
assign w16374 = ~w16304 & w16372;
assign w16375 = w14897 & w15681;
assign w16376 = ~w15681 & w47508;
assign w16377 = ~w16375 & ~w16376;
assign w16378 = w400 & w16377;
assign w16379 = ~w16371 & ~w16378;
assign w16380 = ~w16368 & w16379;
assign w16381 = w351 & w14842;
assign w16382 = ~w14777 & ~w16381;
assign w16383 = w16382 & ~w15791;
assign w16384 = w15669 & ~w16381;
assign w16385 = ~w15667 & w16384;
assign w16386 = ~w15014 & w16385;
assign w16387 = w15666 & w16386;
assign w16388 = ~w16383 & ~w16387;
assign w16389 = w14899 & ~w14972;
assign w16390 = w351 & w14977;
assign w16391 = (~w41333 & w47509) | (~w41333 & w47510) | (w47509 & w47510);
assign w16392 = ~w16388 & ~w16391;
assign w16393 = ~w351 & ~w14842;
assign w16394 = w16389 & w16393;
assign w16395 = (w16394 & w15575) | (w16394 & w41334) | (w15575 & w41334);
assign w16396 = ~w14977 & w16393;
assign w16397 = ~w14854 & ~w16396;
assign w16398 = (~w41334 & w47511) | (~w41334 & w47512) | (w47511 & w47512);
assign w16399 = ~w16388 & w47513;
assign w16400 = ~w15672 & w47514;
assign w16401 = ~w14820 & ~w14978;
assign w16402 = ~w57 & ~w16401;
assign w16403 = ~w16400 & w16402;
assign w16404 = ~w16399 & w16403;
assign w16405 = ~w57 & w16401;
assign w16406 = w16400 & w16405;
assign w16407 = ~w16398 & w16405;
assign w16408 = w16392 & w16407;
assign w16409 = ~w16406 & ~w16408;
assign w16410 = ~w16404 & w16409;
assign w16411 = ~w16395 & ~w16396;
assign w16412 = w16392 & w16411;
assign w16413 = ~w252 & ~w14854;
assign w16414 = (w16413 & ~w16392) | (w16413 & w47515) | (~w16392 & w47515);
assign w16415 = ~w252 & w14854;
assign w16416 = w16392 & w47516;
assign w16417 = ~w16414 & ~w16416;
assign w16418 = w16410 & w16417;
assign w16419 = ~w15677 & w44981;
assign w16420 = ~w15672 & w16419;
assign w16421 = w14966 & ~w14976;
assign w16422 = (w16421 & w15619) | (w16421 & w44982) | (w15619 & w44982);
assign w16423 = ~w14976 & ~w16389;
assign w16424 = (~w16423 & w15575) | (~w16423 & w41335) | (w15575 & w41335);
assign w16425 = ~w15681 & w16424;
assign w16426 = ~w16420 & ~w16425;
assign w16427 = ~w14842 & ~w14975;
assign w16428 = w351 & w16427;
assign w16429 = (w16428 & w16425) | (w16428 & w47517) | (w16425 & w47517);
assign w16430 = w351 & ~w16427;
assign w16431 = ~w16425 & w47518;
assign w16432 = ~w16429 & ~w16431;
assign w16433 = ~w400 & ~w16377;
assign w16434 = w16432 & ~w16433;
assign w16435 = ~w14975 & w16393;
assign w16436 = (~w16435 & w15672) | (~w16435 & w47519) | (w15672 & w47519);
assign w16437 = ~w351 & ~w16427;
assign w16438 = ~w15672 & w47520;
assign w16439 = (w41335 & w47521) | (w41335 & w47522) | (w47521 & w47522);
assign w16440 = ~w15681 & w16439;
assign w16441 = ~w16438 & ~w16440;
assign w16442 = ~w16425 & w16436;
assign w16443 = w16441 & ~w16442;
assign w16444 = w252 & ~w14854;
assign w16445 = w16412 & w16444;
assign w16446 = w252 & w14854;
assign w16447 = (w16446 & ~w16392) | (w16446 & w47523) | (~w16392 & w47523);
assign w16448 = ~w16443 & ~w16447;
assign w16449 = ~w16445 & w16448;
assign w16450 = w14824 & ~w14825;
assign w16451 = ~w14824 & w14825;
assign w16452 = ~w16450 & ~w16451;
assign w16453 = ~w15575 & w41336;
assign w16454 = ~w14973 & w14982;
assign w16455 = ~w14820 & ~w16454;
assign w16456 = w14830 & w14993;
assign w16457 = (~w16456 & w16453) | (~w16456 & w41337) | (w16453 & w41337);
assign w16458 = ~w16453 & w41338;
assign w16459 = w15681 & ~w16452;
assign w16460 = ~w16457 & ~w16458;
assign w16461 = ~w15681 & w16460;
assign w16462 = ~w16459 & ~w16461;
assign w16463 = ~w80 & ~w16462;
assign w16464 = w57 & ~w16401;
assign w16465 = (w16464 & w16399) | (w16464 & w41339) | (w16399 & w41339);
assign w16466 = w57 & w16401;
assign w16467 = ~w16399 & w41340;
assign w16468 = ~w16465 & ~w16467;
assign w16469 = ~w16463 & w16468;
assign w16470 = w16418 & ~w16449;
assign w16471 = w16469 & ~w16470;
assign w16472 = w16418 & w16434;
assign w16473 = ~w16380 & w16472;
assign w16474 = w16471 & ~w16473;
assign w16475 = (w14806 & w15672) | (w14806 & w41341) | (w15672 & w41341);
assign w16476 = w14831 & ~w16454;
assign w16477 = (w14994 & w16453) | (w14994 & w41342) | (w16453 & w41342);
assign w16478 = w16475 & ~w16477;
assign w16479 = w14789 & ~w15004;
assign w16480 = ~w14789 & w15004;
assign w16481 = ~w16479 & ~w16480;
assign w16482 = w14800 & ~w15010;
assign w16483 = (w16482 & ~w41343) | (w16482 & w44983) | (~w41343 & w44983);
assign w16484 = w16478 & ~w16483;
assign w16485 = ~w16478 & w16483;
assign w16486 = ~w16484 & ~w16485;
assign w16487 = w15009 & w15798;
assign w16488 = ~w15790 & w16487;
assign w16489 = (w16488 & w15797) | (w16488 & w41344) | (w15797 & w41344);
assign w16490 = w14770 & ~w15000;
assign w16491 = (w41344 & w44984) | (w41344 & w44985) | (w44984 & w44985);
assign w16492 = w42 & ~w16491;
assign w16493 = ~w14776 & ~w16489;
assign w16494 = w16492 & ~w16493;
assign w16495 = w14708 & ~w14733;
assign w16496 = w14733 & w14748;
assign w16497 = ~w14708 & w16496;
assign w16498 = ~w16495 & ~w16497;
assign w16499 = (w41344 & w44986) | (w41344 & w44987) | (w44986 & w44987);
assign w16500 = w14776 & ~w16498;
assign w16501 = (~w41344 & w44988) | (~w41344 & w44989) | (w44988 & w44989);
assign w16502 = ~w16499 & ~w16501;
assign w16503 = ~w42 & w16502;
assign w16504 = (~w16503 & ~w16486) | (~w16503 & w44990) | (~w16486 & w44990);
assign w16505 = w16486 & w16503;
assign w16506 = w14615 & ~w14801;
assign w16507 = ~w14984 & ~w16506;
assign w16508 = w16507 & ~w16475;
assign w16509 = ~w16478 & ~w16508;
assign w16510 = w14806 & w14988;
assign w16511 = (w14993 & w16453) | (w14993 & w41345) | (w16453 & w41345);
assign w16512 = ~w15681 & ~w16511;
assign w16513 = (w3 & w16509) | (w3 & w44991) | (w16509 & w44991);
assign w16514 = ~w16505 & w16513;
assign w16515 = ~w16504 & ~w16514;
assign w16516 = ~w16279 & w48860;
assign w16517 = ~w16272 & w16516;
assign w16518 = ~w16270 & ~w16517;
assign w16519 = w16232 & ~w16518;
assign w16520 = ~w16188 & w16227;
assign w16521 = ~w16519 & w16520;
assign w16522 = ~w16245 & ~w16521;
assign w16523 = (w16515 & w16521) | (w16515 & w41346) | (w16521 & w41346);
assign w16524 = w16474 & w16523;
assign w16525 = (w16524 & w16117) | (w16524 & w41347) | (w16117 & w41347);
assign w16526 = w80 & w16462;
assign w16527 = ~w16509 & w44992;
assign w16528 = ~w16505 & ~w16527;
assign w16529 = ~w16504 & ~w16528;
assign w16530 = ~w16526 & ~w16529;
assign w16531 = ~w16474 & w16530;
assign w16532 = w15681 & w41348;
assign w16533 = (w754 & ~w16358) | (w754 & w41349) | (~w16358 & w41349);
assign w16534 = ~w15681 & w48861;
assign w16535 = ~w16532 & ~w16534;
assign w16536 = w16356 & ~w16535;
assign w16537 = w16347 & ~w16536;
assign w16538 = w16434 & w16537;
assign w16539 = w16410 & w48862;
assign w16540 = w16538 & w16539;
assign w16541 = (~w16529 & w16540) | (~w16529 & w41350) | (w16540 & w41350);
assign w16542 = ~w16531 & ~w16541;
assign w16543 = (~w15715 & w15703) | (~w15715 & w41351) | (w15703 & w41351);
assign w16544 = w15734 & ~w16543;
assign w16545 = w11870 & ~w16544;
assign w16546 = ~w11870 & w16544;
assign w16547 = ~w16545 & ~w16546;
assign w16548 = ~w16542 & w41352;
assign w16549 = (w15736 & w16542) | (w15736 & w41353) | (w16542 & w41353);
assign w16550 = w16523 & ~w16531;
assign w16551 = ~w16531 & w41354;
assign w16552 = (w16551 & w16117) | (w16551 & w41355) | (w16117 & w41355);
assign w16553 = ~w16549 & ~w16552;
assign w16554 = ~w16525 & w16548;
assign w16555 = w16553 & ~w16554;
assign w16556 = ~w16542 & ~w16550;
assign w16557 = w16299 & ~w16542;
assign w16558 = ~w16117 & w16557;
assign w16559 = ~w16556 & ~w16558;
assign w16560 = w16346 & w16356;
assign w16561 = ~w16299 & ~w16522;
assign w16562 = w16116 & ~w16522;
assign w16563 = ~w15938 & w16562;
assign w16564 = ~w16561 & ~w16563;
assign w16565 = ~w16366 & w16535;
assign w16566 = ~w16563 & w41356;
assign w16567 = ~w16366 & ~w16566;
assign w16568 = ~w16566 & w48863;
assign w16569 = w16346 & ~w16568;
assign w16570 = ~w16559 & ~w16569;
assign w16571 = w16316 & ~w16371;
assign w16572 = (w16571 & w16558) | (w16571 & w48864) | (w16558 & w48864);
assign w16573 = ~w16558 & w48865;
assign w16574 = ~w16572 & ~w16573;
assign w16575 = ~w16570 & w16574;
assign w16576 = ~w16569 & w16572;
assign w16577 = ~w400 & ~w16576;
assign w16578 = ~w16575 & w16577;
assign w16579 = ~w16525 & ~w16542;
assign w16580 = ~w16525 & w48866;
assign w16581 = ~w16378 & ~w16580;
assign w16582 = ~w16563 & w41357;
assign w16583 = ~w16368 & ~w16371;
assign w16584 = ~w16582 & w16583;
assign w16585 = ~w16581 & ~w16584;
assign w16586 = w16380 & ~w16582;
assign w16587 = (w400 & w16558) | (w400 & w47524) | (w16558 & w47524);
assign w16588 = ~w16377 & ~w16587;
assign w16589 = ~w16559 & ~w16586;
assign w16590 = ~w16588 & ~w16589;
assign w16591 = ~w16590 & w48867;
assign w16592 = ~w16578 & ~w16591;
assign w16593 = ~w612 & ~w16579;
assign w16594 = w16568 & ~w16593;
assign w16595 = ~w15681 & ~w16334;
assign w16596 = w16337 & ~w16595;
assign w16597 = ~w16337 & w16595;
assign w16598 = ~w16596 & ~w16597;
assign w16599 = w16559 & w16598;
assign w16600 = ~w16594 & ~w16599;
assign w16601 = (~w16560 & w16558) | (~w16560 & w48868) | (w16558 & w48868);
assign w16602 = ~w16567 & w16601;
assign w16603 = w16600 & ~w16602;
assign w16604 = ~w493 & ~w16603;
assign w16605 = w400 & w16576;
assign w16606 = w400 & w16574;
assign w16607 = ~w16570 & w16606;
assign w16608 = ~w16605 & ~w16607;
assign w16609 = ~w16604 & w16608;
assign w16610 = ~w16361 & ~w16364;
assign w16611 = ~w16564 & ~w16565;
assign w16612 = w16559 & w16610;
assign w16613 = (~w16566 & w16558) | (~w16566 & w48869) | (w16558 & w48869);
assign w16614 = ~w16611 & w16613;
assign w16615 = ~w16612 & ~w16614;
assign w16616 = (~w612 & w16614) | (~w612 & w41358) | (w16614 & w41358);
assign w16617 = w16045 & w48870;
assign w16618 = ~w15938 & w16617;
assign w16619 = (w16518 & w16256) | (w16518 & w41360) | (w16256 & w41360);
assign w16620 = w16232 & w16242;
assign w16621 = w16188 & w16242;
assign w16622 = (~w16621 & w16618) | (~w16621 & w41361) | (w16618 & w41361);
assign w16623 = w16226 & w16622;
assign w16624 = (w16550 & w16117) | (w16550 & w41362) | (w16117 & w41362);
assign w16625 = (w945 & w16531) | (w945 & w41363) | (w16531 & w41363);
assign w16626 = (~w41363 & w44993) | (~w41363 & w44994) | (w44993 & w44994);
assign w16627 = ~w16550 & w16625;
assign w16628 = (~w16626 & w16564) | (~w16626 & w41364) | (w16564 & w41364);
assign w16629 = ~w16234 & w16624;
assign w16630 = (~w945 & w16531) | (~w945 & w41365) | (w16531 & w41365);
assign w16631 = (w16234 & ~w16630) | (w16234 & w44995) | (~w16630 & w44995);
assign w16632 = ~w16563 & w41366;
assign w16633 = ~w16631 & ~w16632;
assign w16634 = (~w754 & w16633) | (~w754 & w44996) | (w16633 & w44996);
assign w16635 = w16628 & w48871;
assign w16636 = w16634 & ~w16635;
assign w16637 = ~w16616 & ~w16636;
assign w16638 = (~w16619 & w15938) | (~w16619 & w41367) | (w15938 & w41367);
assign w16639 = w16242 & w50202;
assign w16640 = ~w16188 & ~w16639;
assign w16641 = w16232 & w16638;
assign w16642 = w16640 & ~w16641;
assign w16643 = w16242 & w16525;
assign w16644 = w16642 & ~w16643;
assign w16645 = (w16622 & w16558) | (w16622 & w48872) | (w16558 & w48872);
assign w16646 = ~w16213 & w16237;
assign w16647 = w16213 & ~w16237;
assign w16648 = ~w16646 & ~w16647;
assign w16649 = ~w1120 & ~w16542;
assign w16650 = w16648 & ~w16649;
assign w16651 = w16550 & w16648;
assign w16652 = ~w16300 & w16651;
assign w16653 = ~w16650 & ~w16652;
assign w16654 = ~w16645 & w16653;
assign w16655 = ~w16644 & ~w16654;
assign w16656 = (~w945 & w16654) | (~w945 & w41369) | (w16654 & w41369);
assign w16657 = (w16623 & ~w16628) | (w16623 & w44997) | (~w16628 & w44997);
assign w16658 = ~w16623 & w16633;
assign w16659 = (w754 & ~w16633) | (w754 & w44998) | (~w16633 & w44998);
assign w16660 = ~w16657 & w16659;
assign w16661 = ~w16656 & ~w16660;
assign w16662 = w16637 & ~w16661;
assign w16663 = w612 & w16615;
assign w16664 = w493 & ~w16602;
assign w16665 = w16600 & w16664;
assign w16666 = ~w16663 & ~w16665;
assign w16667 = ~w16662 & w16666;
assign w16668 = ~w16181 & ~w16638;
assign w16669 = w16231 & ~w16668;
assign w16670 = ~w16559 & ~w16669;
assign w16671 = ~w16151 & w16186;
assign w16672 = w1120 & ~w16671;
assign w16673 = w1120 & ~w16150;
assign w16674 = ~w16558 & w48873;
assign w16675 = (w16672 & w16558) | (w16672 & w41370) | (w16558 & w41370);
assign w16676 = w16669 & w16675;
assign w16677 = ~w16674 & ~w16676;
assign w16678 = w1120 & w16671;
assign w16679 = ~w16559 & w48874;
assign w16680 = w16677 & ~w16679;
assign w16681 = ~w16654 & w41371;
assign w16682 = w16680 & ~w16681;
assign w16683 = w16637 & w16682;
assign w16684 = ~w1120 & w16671;
assign w16685 = ~w1120 & w16150;
assign w16686 = ~w16558 & w48875;
assign w16687 = (w16684 & w16558) | (w16684 & w41372) | (w16558 & w41372);
assign w16688 = w16669 & w16687;
assign w16689 = ~w16686 & ~w16688;
assign w16690 = ~w1120 & ~w16671;
assign w16691 = ~w16559 & w48876;
assign w16692 = w16689 & ~w16691;
assign w16693 = ~w16168 & w16179;
assign w16694 = ~w1541 & w16638;
assign w16695 = w1541 & ~w16638;
assign w16696 = ~w16559 & w41373;
assign w16697 = w1320 & ~w16693;
assign w16698 = (w16697 & w16559) | (w16697 & w48877) | (w16559 & w48877);
assign w16699 = w1320 & w16693;
assign w16700 = ~w16559 & w48878;
assign w16701 = ~w16698 & ~w16700;
assign w16702 = w16692 & w16701;
assign w16703 = ~w16270 & ~w16272;
assign w16704 = ~w16256 & ~w16296;
assign w16705 = (~w16516 & w16117) | (~w16516 & w41374) | (w16117 & w41374);
assign w16706 = w16703 & ~w16705;
assign w16707 = ~w16703 & w16705;
assign w16708 = ~w16706 & ~w16707;
assign w16709 = ~w16559 & ~w16708;
assign w16710 = ~w16558 & w48879;
assign w16711 = ~w1541 & ~w16710;
assign w16712 = ~w16709 & w16711;
assign w16713 = ~w1320 & w16693;
assign w16714 = (w16713 & w16559) | (w16713 & w48880) | (w16559 & w48880);
assign w16715 = ~w1320 & ~w16693;
assign w16716 = ~w16559 & w48881;
assign w16717 = ~w16714 & ~w16716;
assign w16718 = ~w16712 & w16717;
assign w16719 = w16702 & ~w16718;
assign w16720 = w16683 & ~w16719;
assign w16721 = w16667 & ~w16720;
assign w16722 = (w16609 & w16720) | (w16609 & w48882) | (w16720 & w48882);
assign w16723 = (w16592 & w16721) | (w16592 & w44999) | (w16721 & w44999);
assign w16724 = ~w16380 & w16434;
assign w16725 = w16449 & ~w16724;
assign w16726 = (w16725 & w16563) | (w16725 & w41376) | (w16563 & w41376);
assign w16727 = ~w16558 & w47525;
assign w16728 = ~w16559 & w41377;
assign w16729 = ~w16727 & ~w16728;
assign w16730 = w16410 & w16468;
assign w16731 = ~w80 & ~w16730;
assign w16732 = (w16731 & w16728) | (w16731 & w47526) | (w16728 & w47526);
assign w16733 = ~w80 & w16730;
assign w16734 = ~w16728 & w47527;
assign w16735 = ~w16732 & ~w16734;
assign w16736 = w16418 & ~w16725;
assign w16737 = w16418 & w16538;
assign w16738 = ~w16563 & w41378;
assign w16739 = ~w16736 & ~w16738;
assign w16740 = (w16526 & w16558) | (w16526 & w41379) | (w16558 & w41379);
assign w16741 = ~w16739 & ~w16740;
assign w16742 = ~w16468 & ~w16526;
assign w16743 = ~w16558 & w41380;
assign w16744 = ~w16742 & ~w16743;
assign w16745 = w80 & w16579;
assign w16746 = ~w16462 & ~w16745;
assign w16747 = ~w16741 & w16744;
assign w16748 = ~w16746 & ~w16747;
assign w16749 = (w16463 & w16558) | (w16463 & w41381) | (w16558 & w41381);
assign w16750 = ~w16526 & ~w16749;
assign w16751 = w16468 & w16739;
assign w16752 = ~w16750 & w16751;
assign w16753 = (w3 & w16750) | (w3 & w47528) | (w16750 & w47528);
assign w16754 = ~w16748 & w16753;
assign w16755 = w16735 & ~w16754;
assign w16756 = ~w16443 & ~w16724;
assign w16757 = ~w16563 & w41382;
assign w16758 = w16756 & ~w16757;
assign w16759 = w14854 & ~w16412;
assign w16760 = ~w14854 & w16412;
assign w16761 = ~w16759 & ~w16760;
assign w16762 = w252 & w16761;
assign w16763 = ~w252 & ~w16761;
assign w16764 = ~w16542 & w16763;
assign w16765 = ~w16525 & w16764;
assign w16766 = ~w16762 & ~w16765;
assign w16767 = ~w16559 & ~w16758;
assign w16768 = ~w16558 & w41383;
assign w16769 = ~w16762 & ~w16763;
assign w16770 = (w16769 & w16558) | (w16769 & w41384) | (w16558 & w41384);
assign w16771 = ~w16768 & ~w16770;
assign w16772 = ~w16758 & ~w16766;
assign w16773 = ~w16767 & ~w16771;
assign w16774 = ~w16772 & ~w16773;
assign w16775 = ~w16773 & w47529;
assign w16776 = w80 & w16730;
assign w16777 = (w16776 & w16728) | (w16776 & w47530) | (w16728 & w47530);
assign w16778 = w80 & ~w16730;
assign w16779 = ~w16728 & w47531;
assign w16780 = ~w16777 & ~w16779;
assign w16781 = w16775 & w16780;
assign w16782 = ~w16748 & ~w16752;
assign w16783 = (~w3 & w16748) | (~w3 & w47532) | (w16748 & w47532);
assign w16784 = ~w80 & w15681;
assign w16785 = ~w16512 & ~w16784;
assign w16786 = w16510 & ~w16785;
assign w16787 = ~w16510 & w16785;
assign w16788 = ~w16786 & ~w16787;
assign w16789 = ~w16474 & ~w16526;
assign w16790 = ~w16563 & w41385;
assign w16791 = ~w16789 & ~w16790;
assign w16792 = ~w3 & ~w16529;
assign w16793 = (w3 & w16558) | (w3 & w41386) | (w16558 & w41386);
assign w16794 = w16791 & w16793;
assign w16795 = ~w16794 & w47533;
assign w16796 = (~w16788 & w16794) | (~w16788 & w47534) | (w16794 & w47534);
assign w16797 = ~w16795 & ~w16796;
assign w16798 = ~w42 & w16797;
assign w16799 = ~w16783 & ~w16798;
assign w16800 = w16755 & ~w16781;
assign w16801 = w16799 & ~w16800;
assign w16802 = ~w16527 & ~w16791;
assign w16803 = ~w16513 & ~w16802;
assign w16804 = ~w42 & w16486;
assign w16805 = w42 & ~w16486;
assign w16806 = ~w16804 & ~w16805;
assign w16807 = ~w16503 & ~w16806;
assign w16808 = ~w16803 & w16807;
assign w16809 = ~w16494 & w16806;
assign w16810 = w16803 & w16809;
assign w16811 = ~w16808 & ~w16810;
assign w16812 = w42 & ~w16797;
assign w16813 = w16811 & ~w16812;
assign w16814 = (~w16432 & w16558) | (~w16432 & w41387) | (w16558 & w41387);
assign w16815 = ~w16443 & ~w16814;
assign w16816 = ~w16433 & ~w16586;
assign w16817 = ~w16815 & w16816;
assign w16818 = w16426 & ~w16427;
assign w16819 = ~w16426 & w16427;
assign w16820 = ~w16818 & ~w16819;
assign w16821 = (w16820 & w16559) | (w16820 & w47535) | (w16559 & w47535);
assign w16822 = w16579 & w16758;
assign w16823 = ~w351 & w16822;
assign w16824 = ~w16817 & w47536;
assign w16825 = w252 & ~w16824;
assign w16826 = (~w351 & w16590) | (~w351 & w48883) | (w16590 & w48883);
assign w16827 = ~w16825 & ~w16826;
assign w16828 = w16813 & w16827;
assign w16829 = ~w16801 & w16828;
assign w16830 = ~w16723 & w16829;
assign w16831 = w16038 & ~w16251;
assign w16832 = ~w15938 & ~w15939;
assign w16833 = ~w16558 & w41388;
assign w16834 = (w16832 & w16558) | (w16832 & w41389) | (w16558 & w41389);
assign w16835 = ~w16833 & ~w16834;
assign w16836 = w16831 & w16835;
assign w16837 = ~w16831 & ~w16835;
assign w16838 = ~w16836 & ~w16837;
assign w16839 = w4838 & w16838;
assign w16840 = w15880 & ~w15913;
assign w16841 = w15777 & ~w16840;
assign w16842 = (w15880 & w15816) | (w15880 & w16840) | (w15816 & w16840);
assign w16843 = (w16842 & w15728) | (w16842 & w41390) | (w15728 & w41390);
assign w16844 = w15914 & ~w16843;
assign w16845 = ~w15890 & ~w15891;
assign w16846 = w6264 & w16845;
assign w16847 = ~w16844 & w16846;
assign w16848 = ~w16542 & ~w16847;
assign w16849 = ~w16558 & w41391;
assign w16850 = ~w16624 & w16848;
assign w16851 = ~w16849 & ~w16850;
assign w16852 = ~w16844 & w16845;
assign w16853 = ~w6264 & ~w16852;
assign w16854 = w16848 & ~w16853;
assign w16855 = ~w16624 & w16854;
assign w16856 = w15900 & w16855;
assign w16857 = ~w16851 & ~w16856;
assign w16858 = ~w15934 & ~w15939;
assign w16859 = ~w5330 & ~w16858;
assign w16860 = w16857 & w16859;
assign w16861 = ~w5330 & w16858;
assign w16862 = ~w16857 & w16861;
assign w16863 = ~w16860 & ~w16862;
assign w16864 = ~w16839 & w16863;
assign w16865 = (~w4838 & w16558) | (~w4838 & w41392) | (w16558 & w41392);
assign w16866 = w16026 & ~w16865;
assign w16867 = (w41393 & ~w15937) | (w41393 & w50343) | (~w15937 & w50343);
assign w16868 = ~w16027 & ~w16251;
assign w16869 = ~w16867 & w16868;
assign w16870 = (~w16869 & w16558) | (~w16869 & w47537) | (w16558 & w47537);
assign w16871 = ~w16251 & ~w16867;
assign w16872 = w16027 & ~w16871;
assign w16873 = w16040 & ~w16871;
assign w16874 = w16579 & w16873;
assign w16875 = ~w16872 & ~w16874;
assign w16876 = ~w16866 & ~w16870;
assign w16877 = w16875 & ~w16876;
assign w16878 = (w4430 & w16876) | (w4430 & w47538) | (w16876 & w47538);
assign w16879 = ~w4838 & ~w16838;
assign w16880 = ~w16878 & ~w16879;
assign w16881 = ~w16864 & w16880;
assign w16882 = ~w4430 & w16877;
assign w16883 = ~w15997 & ~w16007;
assign w16884 = (w41394 & w16558) | (w41394 & w47539) | (w16558 & w47539);
assign w16885 = ~w16558 & w47540;
assign w16886 = ~w16884 & ~w16885;
assign w16887 = w16883 & ~w16886;
assign w16888 = ~w16883 & w16886;
assign w16889 = ~w16887 & ~w16888;
assign w16890 = ~w4056 & ~w16889;
assign w16891 = ~w16882 & ~w16890;
assign w16892 = ~w16881 & w16891;
assign w16893 = w2006 & w52247;
assign w16894 = ~w2006 & ~w52247;
assign w16895 = ~w16559 & w41396;
assign w16896 = ~w1738 & w16280;
assign w16897 = (w16896 & w16559) | (w16896 & w48884) | (w16559 & w48884);
assign w16898 = ~w1738 & ~w16280;
assign w16899 = ~w16559 & w48885;
assign w16900 = ~w16897 & ~w16899;
assign w16901 = ~w16115 & w16298;
assign w16902 = (w16901 & w15938) | (w16901 & w41397) | (w15938 & w41397);
assign w16903 = ~w16110 & w16524;
assign w16904 = ~w16902 & w16903;
assign w16905 = w16064 & ~w16542;
assign w16906 = ~w16110 & ~w16905;
assign w16907 = ~w15939 & ~w16103;
assign w16908 = w16045 & w16907;
assign w16909 = w16045 & w41398;
assign w16910 = ~w15938 & w16909;
assign w16911 = w16111 & ~w16254;
assign w16912 = w16045 & w16911;
assign w16913 = w16096 & w16293;
assign w16914 = w16288 & w16913;
assign w16915 = ~w16912 & w16914;
assign w16916 = ~w16082 & ~w16099;
assign w16917 = (~w16916 & w16910) | (~w16916 & w41399) | (w16910 & w41399);
assign w16918 = ~w16904 & ~w16917;
assign w16919 = ~w16906 & w16918;
assign w16920 = (~w2285 & w16531) | (~w2285 & w48886) | (w16531 & w48886);
assign w16921 = ~w16063 & ~w16920;
assign w16922 = ~w16531 & w48887;
assign w16923 = ~w16300 & w16922;
assign w16924 = ~w16921 & ~w16923;
assign w16925 = (w16110 & w16558) | (w16110 & w41400) | (w16558 & w41400);
assign w16926 = w16924 & ~w16925;
assign w16927 = ~w16559 & ~w16917;
assign w16928 = w16918 & w48888;
assign w16929 = (~w2006 & w16559) | (~w2006 & w41401) | (w16559 & w41401);
assign w16930 = w16926 & w16929;
assign w16931 = ~w16928 & ~w16930;
assign w16932 = w16081 & ~w16556;
assign w16933 = ~w16558 & w16932;
assign w16934 = w2558 & w16081;
assign w16935 = ~w16082 & ~w16934;
assign w16936 = (w16096 & w16912) | (w16096 & w41402) | (w16912 & w41402);
assign w16937 = ~w16935 & ~w16936;
assign w16938 = w16096 & w16909;
assign w16939 = ~w15938 & w16938;
assign w16940 = w16937 & ~w16939;
assign w16941 = w16096 & w16935;
assign w16942 = ~w16915 & w16941;
assign w16943 = w16909 & w16941;
assign w16944 = ~w15938 & w16943;
assign w16945 = ~w16942 & ~w16944;
assign w16946 = ~w16940 & w16945;
assign w16947 = ~w16559 & ~w16946;
assign w16948 = ~w16933 & ~w16947;
assign w16949 = (~w2285 & w16947) | (~w2285 & w41403) | (w16947 & w41403);
assign w16950 = w2285 & ~w16933;
assign w16951 = ~w16947 & w16950;
assign w16952 = (w16915 & w15938) | (w16915 & w41404) | (w15938 & w41404);
assign w16953 = w16288 & ~w16912;
assign w16954 = ~w16913 & ~w16953;
assign w16955 = w16909 & ~w16913;
assign w16956 = ~w15938 & w16955;
assign w16957 = ~w16954 & ~w16956;
assign w16958 = ~w16952 & w16957;
assign w16959 = ~w16559 & w16958;
assign w16960 = w15139 & w15681;
assign w16961 = ~w15681 & ~w16091;
assign w16962 = ~w16960 & ~w16961;
assign w16963 = ~w16556 & w16962;
assign w16964 = ~w16558 & w16963;
assign w16965 = ~w2558 & ~w16964;
assign w16966 = ~w16959 & w16965;
assign w16967 = ~w16951 & ~w16966;
assign w16968 = ~w16949 & ~w16967;
assign w16969 = w16931 & w16968;
assign w16970 = w16926 & ~w16927;
assign w16971 = w2006 & ~w16919;
assign w16972 = ~w16970 & w16971;
assign w16973 = w1738 & ~w16280;
assign w16974 = ~w16895 & w16973;
assign w16975 = w1738 & w16280;
assign w16976 = w16895 & w16975;
assign w16977 = ~w16974 & ~w16976;
assign w16978 = ~w16972 & w16977;
assign w16979 = (w16900 & w16969) | (w16900 & w47541) | (w16969 & w47541);
assign w16980 = w16028 & ~w16252;
assign w16981 = ~w15997 & w16041;
assign w16982 = ~w15939 & w16981;
assign w16983 = w16980 & w16982;
assign w16984 = ~w15997 & ~w16980;
assign w16985 = ~w15987 & w16005;
assign w16986 = ~w16984 & w16985;
assign w16987 = w16984 & ~w16985;
assign w16988 = ~w16986 & ~w16987;
assign w16989 = ~w15938 & w41405;
assign w16990 = (w16988 & w15938) | (w16988 & w41406) | (w15938 & w41406);
assign w16991 = ~w16989 & ~w16990;
assign w16992 = w15981 & w16000;
assign w16993 = ~w15981 & ~w16000;
assign w16994 = ~w16992 & ~w16993;
assign w16995 = (w16991 & w16558) | (w16991 & w48889) | (w16558 & w48889);
assign w16996 = ~w16558 & w41407;
assign w16997 = ~w16995 & ~w16996;
assign w16998 = ~w16995 & w41408;
assign w16999 = w16005 & ~w16986;
assign w17000 = w16005 & w16982;
assign w17001 = (~w16999 & w15938) | (~w16999 & w41409) | (w15938 & w41409);
assign w17002 = (~w17001 & w16558) | (~w17001 & w47542) | (w16558 & w47542);
assign w17003 = ~w3646 & ~w16556;
assign w17004 = ~w16558 & w17003;
assign w17005 = w15972 & ~w16103;
assign w17006 = ~w3242 & w17005;
assign w17007 = ~w17004 & w17006;
assign w17008 = ~w17002 & w17007;
assign w17009 = ~w3242 & ~w17005;
assign w17010 = w17004 & w17009;
assign w17011 = ~w17001 & w17009;
assign w17012 = (w17011 & w16558) | (w17011 & w47543) | (w16558 & w47543);
assign w17013 = ~w17010 & ~w17012;
assign w17014 = ~w17008 & w17013;
assign w17015 = w16254 & w16908;
assign w17016 = ~w15938 & w17015;
assign w17017 = ~w16103 & ~w16254;
assign w17018 = w16045 & w17017;
assign w17019 = ~w16109 & w16288;
assign w17020 = w17018 & ~w17019;
assign w17021 = ~w17018 & w17019;
assign w17022 = ~w17020 & ~w17021;
assign w17023 = w17016 & w17022;
assign w17024 = ~w17016 & ~w17022;
assign w17025 = ~w17023 & ~w17024;
assign w17026 = ~w16558 & w41410;
assign w17027 = ~w16559 & w17025;
assign w17028 = ~w17026 & ~w17027;
assign w17029 = (~w2896 & w17027) | (~w2896 & w41411) | (w17027 & w41411);
assign w17030 = w3242 & ~w17005;
assign w17031 = ~w17004 & w17030;
assign w17032 = ~w17002 & w17031;
assign w17033 = w3242 & w17005;
assign w17034 = w17004 & w17033;
assign w17035 = ~w17001 & w17033;
assign w17036 = (w17035 & w16558) | (w17035 & w47544) | (w16558 & w47544);
assign w17037 = ~w17034 & ~w17036;
assign w17038 = ~w17032 & w17037;
assign w17039 = ~w17029 & w17038;
assign w17040 = w16998 & w17014;
assign w17041 = w17039 & ~w17040;
assign w17042 = ~w17027 & w48890;
assign w17043 = ~w17041 & ~w17042;
assign w17044 = ~w16959 & ~w16964;
assign w17045 = (w2558 & w16959) | (w2558 & w48891) | (w16959 & w48891);
assign w17046 = ~w16949 & ~w17045;
assign w17047 = w16900 & w16931;
assign w17048 = w17046 & w17047;
assign w17049 = ~w17043 & w17048;
assign w17050 = ~w16979 & ~w17049;
assign w17051 = w16892 & ~w17050;
assign w17052 = ~w3646 & ~w16997;
assign w17053 = w4056 & ~w16883;
assign w17054 = ~w16886 & w17053;
assign w17055 = w4056 & w16883;
assign w17056 = w16886 & w17055;
assign w17057 = ~w17054 & ~w17056;
assign w17058 = ~w17052 & w17057;
assign w17059 = w17014 & ~w17042;
assign w17060 = w17058 & w17059;
assign w17061 = ~w17043 & w47545;
assign w17062 = ~w16979 & ~w17061;
assign w17063 = ~w15871 & ~w16842;
assign w17064 = ~w15871 & w16841;
assign w17065 = ~w15728 & w17064;
assign w17066 = ~w17063 & ~w17065;
assign w17067 = (w41413 & w16531) | (w41413 & w47546) | (w16531 & w47546);
assign w17068 = (w41414 & w16531) | (w41414 & w47547) | (w16531 & w47547);
assign w17069 = ~w17067 & ~w17068;
assign w17070 = w15824 & w17068;
assign w17071 = ~w16624 & w17070;
assign w17072 = w15824 & w17067;
assign w17073 = ~w16525 & w17072;
assign w17074 = ~w17071 & ~w17073;
assign w17075 = (~w15824 & w16624) | (~w15824 & w47548) | (w16624 & w47548);
assign w17076 = w17074 & ~w17075;
assign w17077 = ~w6769 & ~w17076;
assign w17078 = w17074 & w47549;
assign w17079 = w7924 & ~w16843;
assign w17080 = ~w7924 & w16843;
assign w17081 = ~w17079 & ~w17080;
assign w17082 = (~w17081 & w16558) | (~w17081 & w41415) | (w16558 & w41415);
assign w17083 = ~w15870 & ~w17082;
assign w17084 = w15870 & ~w17081;
assign w17085 = w16579 & w17084;
assign w17086 = ~w17083 & ~w17085;
assign w17087 = ~w17083 & w47550;
assign w17088 = ~w17078 & ~w17087;
assign w17089 = ~w17077 & ~w17088;
assign w17090 = w15900 & ~w16855;
assign w17091 = ~w15900 & w16855;
assign w17092 = ~w17090 & ~w17091;
assign w17093 = w5745 & w17092;
assign w17094 = ~w15854 & ~w15891;
assign w17095 = w15887 & w17066;
assign w17096 = ~w15825 & ~w17095;
assign w17097 = ~w17094 & w17096;
assign w17098 = w17094 & ~w17096;
assign w17099 = ~w16558 & w47551;
assign w17100 = ~w17097 & ~w17098;
assign w17101 = ~w16559 & w17100;
assign w17102 = ~w17099 & ~w17101;
assign w17103 = ~w6264 & w17102;
assign w17104 = ~w17093 & ~w17103;
assign w17105 = ~w17089 & w17104;
assign w17106 = ~w5745 & ~w17092;
assign w17107 = (w6264 & w17101) | (w6264 & w47552) | (w17101 & w47552);
assign w17108 = ~w17106 & ~w17107;
assign w17109 = ~w17093 & ~w17108;
assign w17110 = w15322 & ~w15875;
assign w17111 = ~w15322 & w15875;
assign w17112 = ~w17110 & ~w17111;
assign w17113 = ~w15816 & ~w15907;
assign w17114 = w15777 & ~w15907;
assign w17115 = (~w17113 & w15728) | (~w17113 & w41416) | (w15728 & w41416);
assign w17116 = ~w8666 & ~w17115;
assign w17117 = w8666 & w17115;
assign w17118 = ~w16542 & w41417;
assign w17119 = (~w17112 & w16624) | (~w17112 & w47553) | (w16624 & w47553);
assign w17120 = ~w16542 & w47554;
assign w17121 = ~w16525 & w17120;
assign w17122 = w7924 & ~w17121;
assign w17123 = ~w17119 & w17122;
assign w17124 = (w15739 & w15704) | (w15739 & w41418) | (w15704 & w41418);
assign w17125 = w15781 & ~w17124;
assign w17126 = ~w15769 & ~w17125;
assign w17127 = w15754 & w17126;
assign w17128 = w15509 & w15681;
assign w17129 = ~w15681 & w15749;
assign w17130 = ~w17128 & ~w17129;
assign w17131 = (w10419 & w16558) | (w10419 & w41419) | (w16558 & w41419);
assign w17132 = ~w17130 & ~w17131;
assign w17133 = (~w17127 & w16558) | (~w17127 & w47555) | (w16558 & w47555);
assign w17134 = ~w17132 & ~w17133;
assign w17135 = ~w15754 & ~w17126;
assign w17136 = ~w15774 & ~w17126;
assign w17137 = w16579 & w17136;
assign w17138 = ~w17135 & ~w17137;
assign w17139 = ~w17134 & w17138;
assign w17140 = (w9781 & w17134) | (w9781 & w47556) | (w17134 & w47556);
assign w17141 = w15774 & w15814;
assign w17142 = ~w17127 & w17141;
assign w17143 = (~w17142 & w16558) | (~w17142 & w41420) | (w16558 & w41420);
assign w17144 = w15529 & ~w15809;
assign w17145 = ~w15529 & w15809;
assign w17146 = ~w17144 & ~w17145;
assign w17147 = w16550 & ~w17146;
assign w17148 = ~w16300 & w17147;
assign w17149 = ~w9781 & ~w16542;
assign w17150 = ~w17146 & ~w17149;
assign w17151 = w15774 & ~w17127;
assign w17152 = ~w15755 & ~w16542;
assign w17153 = ~w15814 & ~w17151;
assign w17154 = ~w17151 & w17152;
assign w17155 = ~w16525 & w17154;
assign w17156 = ~w17153 & ~w17155;
assign w17157 = ~w17148 & ~w17150;
assign w17158 = ~w17143 & w17157;
assign w17159 = w17156 & ~w17158;
assign w17160 = ~w17158 & w41421;
assign w17161 = ~w15808 & ~w15907;
assign w17162 = w15755 & ~w17141;
assign w17163 = w15756 & ~w15769;
assign w17164 = ~w17125 & w17163;
assign w17165 = ~w17162 & ~w17164;
assign w17166 = w17161 & ~w17165;
assign w17167 = ~w17161 & w17165;
assign w17168 = ~w17166 & ~w17167;
assign w17169 = (w17168 & w16558) | (w17168 & w48892) | (w16558 & w48892);
assign w17170 = ~w16558 & w41422;
assign w17171 = ~w17169 & ~w17170;
assign w17172 = ~w17169 & w41423;
assign w17173 = ~w17123 & ~w17172;
assign w17174 = ~w17160 & w17173;
assign w17175 = ~w17140 & w17174;
assign w17176 = ~w16558 & w41424;
assign w17177 = ~w9387 & ~w17176;
assign w17178 = ~w16559 & w41425;
assign w17179 = w17177 & ~w17178;
assign w17180 = ~w7924 & ~w17112;
assign w17181 = (w17180 & w16624) | (w17180 & w47557) | (w16624 & w47557);
assign w17182 = ~w7924 & w17121;
assign w17183 = ~w17181 & ~w17182;
assign w17184 = (~w8666 & w17169) | (~w8666 & w41426) | (w17169 & w41426);
assign w17185 = w17183 & ~w17184;
assign w17186 = ~w17159 & ~w17179;
assign w17187 = w17185 & ~w17186;
assign w17188 = (~w17123 & w17186) | (~w17123 & w41427) | (w17186 & w41427);
assign w17189 = ~w17175 & ~w17188;
assign w17190 = w7315 & ~w17086;
assign w17191 = ~w17077 & ~w17190;
assign w17192 = ~w17105 & ~w17109;
assign w17193 = ~w17109 & w17191;
assign w17194 = ~w17189 & w17193;
assign w17195 = ~w17192 & ~w17194;
assign w17196 = ~a[42] & ~a[43];
assign w17197 = ~a[44] & w17196;
assign w17198 = ~w15681 & w17197;
assign w17199 = w15681 & ~w17197;
assign w17200 = a[45] & w17199;
assign w17201 = ~w15641 & ~w17200;
assign w17202 = ~w17198 & ~w17201;
assign w17203 = a[45] & ~w17198;
assign w17204 = ~w17199 & ~w17203;
assign w17205 = w14766 & w17202;
assign w17206 = (w17205 & w16558) | (w17205 & w41428) | (w16558 & w41428);
assign w17207 = w14766 & ~w17204;
assign w17208 = ~w16558 & w41429;
assign w17209 = ~w17206 & ~w17208;
assign w17210 = ~a[46] & ~w15681;
assign w17211 = a[46] & w15681;
assign w17212 = a[46] & ~w15641;
assign w17213 = ~w15642 & ~w17212;
assign w17214 = ~w17210 & ~w17211;
assign w17215 = ~w16558 & w41430;
assign w17216 = (w17213 & w16558) | (w17213 & w41431) | (w16558 & w41431);
assign w17217 = ~w17215 & ~w17216;
assign w17218 = w17209 & ~w17217;
assign w17219 = ~w14766 & ~w17202;
assign w17220 = (w17219 & w16558) | (w17219 & w41432) | (w16558 & w41432);
assign w17221 = ~w14766 & w17204;
assign w17222 = ~w16558 & w41433;
assign w17223 = ~w17220 & ~w17222;
assign w17224 = (w14039 & w17218) | (w14039 & w47558) | (w17218 & w47558);
assign w17225 = ~w14766 & ~w15641;
assign w17226 = w15681 & w17225;
assign w17227 = ~w16529 & w17226;
assign w17228 = a[46] & ~w17227;
assign w17229 = ~w14766 & ~w15681;
assign w17230 = w14766 & w15681;
assign w17231 = ~w17229 & ~w17230;
assign w17232 = w15642 & ~w17231;
assign w17233 = ~w15642 & w17231;
assign w17234 = ~w17232 & ~w17233;
assign w17235 = (~w17234 & w16531) | (~w17234 & w48893) | (w16531 & w48893);
assign w17236 = ~a[47] & ~w17228;
assign w17237 = ~a[47] & w17235;
assign w17238 = (~w17236 & w16624) | (~w17236 & w48894) | (w16624 & w48894);
assign w17239 = w14766 & w15641;
assign w17240 = ~w17225 & ~w17239;
assign w17241 = w15681 & ~w17240;
assign w17242 = ~w16542 & w17241;
assign w17243 = ~w16525 & w17242;
assign w17244 = ~w17212 & w17240;
assign w17245 = (~w17244 & w16531) | (~w17244 & w48895) | (w16531 & w48895);
assign w17246 = ~w16531 & w48896;
assign w17247 = ~w16300 & w17246;
assign w17248 = ~w15681 & ~w17245;
assign w17249 = ~w17247 & ~w17248;
assign w17250 = ~w17243 & w17249;
assign w17251 = ~w17238 & ~w17250;
assign w17252 = w15687 & w17231;
assign w17253 = w16579 & w17252;
assign w17254 = ~w16531 & w48897;
assign w17255 = ~w16300 & w17254;
assign w17256 = a[47] & ~w17235;
assign w17257 = ~w17255 & ~w17256;
assign w17258 = w16542 & w17210;
assign w17259 = w16524 & w17210;
assign w17260 = (w17259 & w16117) | (w17259 & w41434) | (w16117 & w41434);
assign w17261 = ~w17258 & ~w17260;
assign w17262 = ~w17257 & w17261;
assign w17263 = ~w17253 & ~w17262;
assign w17264 = ~w17251 & w17263;
assign w17265 = ~w14039 & w17223;
assign w17266 = ~w17218 & w17265;
assign w17267 = w17264 & ~w17266;
assign w17268 = ~w17224 & ~w17267;
assign w17269 = ~w15686 & ~w15700;
assign w17270 = ~w15688 & w17269;
assign w17271 = (w17270 & w16558) | (w17270 & w41435) | (w16558 & w41435);
assign w17272 = w15696 & ~w17271;
assign w17273 = ~w15696 & w17271;
assign w17274 = ~w17272 & ~w17273;
assign w17275 = ~w13384 & w17274;
assign w17276 = w16553 & w48898;
assign w17277 = w11138 & w17125;
assign w17278 = ~w16542 & w17277;
assign w17279 = ~w16525 & w17278;
assign w17280 = w15769 & w17124;
assign w17281 = (w17280 & w16558) | (w17280 & w41436) | (w16558 & w41436);
assign w17282 = ~w17279 & ~w17281;
assign w17283 = w11138 & w17124;
assign w17284 = ~w17125 & ~w17283;
assign w17285 = ~w15765 & ~w15767;
assign w17286 = ~w17284 & ~w17285;
assign w17287 = ~w16556 & ~w17285;
assign w17288 = ~w16558 & w17287;
assign w17289 = ~w17286 & ~w17288;
assign w17290 = ~w17288 & w41437;
assign w17291 = w17282 & w17290;
assign w17292 = ~w17276 & ~w17291;
assign w17293 = (w16542 & w48899) | (w16542 & w48900) | (w48899 & w48900);
assign w17294 = ~w16531 & w49665;
assign w17295 = ~w16300 & w17294;
assign w17296 = ~w17293 & ~w17295;
assign w17297 = ~w16542 & w48901;
assign w17298 = ~w16525 & w17297;
assign w17299 = w17296 & ~w17298;
assign w17300 = w12666 & ~w15704;
assign w17301 = ~w12666 & w15704;
assign w17302 = ~w17300 & ~w17301;
assign w17303 = (w17302 & w16531) | (w17302 & w41438) | (w16531 & w41438);
assign w17304 = w15714 & ~w17303;
assign w17305 = w15714 & w16524;
assign w17306 = (w17305 & w16117) | (w17305 & w41439) | (w16117 & w41439);
assign w17307 = ~w17304 & ~w17306;
assign w17308 = ~w15714 & w17303;
assign w17309 = ~w16531 & w48902;
assign w17310 = ~w16300 & w17309;
assign w17311 = (w11870 & ~w17303) | (w11870 & w48903) | (~w17303 & w48903);
assign w17312 = ~w17310 & ~w17311;
assign w17313 = w17307 & ~w17312;
assign w17314 = ~w15698 & ~w15700;
assign w17315 = ~w15640 & ~w15701;
assign w17316 = w17314 & ~w17315;
assign w17317 = ~w17314 & w17315;
assign w17318 = ~w17316 & ~w17317;
assign w17319 = ~w16558 & w41440;
assign w17320 = (w17318 & w16558) | (w17318 & w41441) | (w16558 & w41441);
assign w17321 = ~w17319 & ~w17320;
assign w17322 = w12666 & w17321;
assign w17323 = w17299 & w17313;
assign w17324 = ~w17322 & ~w17323;
assign w17325 = w17292 & w17324;
assign w17326 = w17324 & w41442;
assign w17327 = w17268 & w17326;
assign w17328 = w13384 & ~w17274;
assign w17329 = ~w12666 & ~w17321;
assign w17330 = ~w17328 & ~w17329;
assign w17331 = w17325 & ~w17330;
assign w17332 = w17282 & w17289;
assign w17333 = ~w10419 & ~w17332;
assign w17334 = ~w16624 & w17308;
assign w17335 = w17307 & ~w17334;
assign w17336 = ~w11870 & ~w17335;
assign w17337 = w17299 & ~w17336;
assign w17338 = w17292 & ~w17337;
assign w17339 = ~w17333 & ~w17338;
assign w17340 = ~w17331 & w17339;
assign w17341 = ~w17327 & w17340;
assign w17342 = ~w9781 & w17139;
assign w17343 = w17187 & ~w17342;
assign w17344 = w17105 & w17343;
assign w17345 = w17341 & w17344;
assign w17346 = ~w17195 & ~w17345;
assign w17347 = w16857 & ~w16858;
assign w17348 = ~w16857 & w16858;
assign w17349 = ~w17347 & ~w17348;
assign w17350 = w5330 & w17349;
assign w17351 = w16880 & ~w17350;
assign w17352 = ~w17051 & w17062;
assign w17353 = ~w17061 & w41443;
assign w17354 = w17346 & w17353;
assign w17355 = ~w17352 & ~w17354;
assign w17356 = ~w17354 & w41444;
assign w17357 = (w16813 & w16800) | (w16813 & w47559) | (w16800 & w47559);
assign w17358 = ~w16558 & w48904;
assign w17359 = w1541 & ~w17358;
assign w17360 = ~w16559 & w16708;
assign w17361 = w17359 & ~w17360;
assign w17362 = w16717 & w17361;
assign w17363 = w16702 & ~w17362;
assign w17364 = w16683 & ~w17363;
assign w17365 = w16667 & ~w17364;
assign w17366 = w16609 & w16827;
assign w17367 = ~w17365 & w17366;
assign w17368 = (~w57 & w16773) | (~w57 & w47560) | (w16773 & w47560);
assign w17369 = w16780 & ~w17368;
assign w17370 = ~w252 & w16824;
assign w17371 = w17369 & ~w17370;
assign w17372 = w16799 & w17371;
assign w17373 = ~w16592 & w16827;
assign w17374 = w17372 & ~w17373;
assign w17375 = ~w17367 & w17374;
assign w17376 = (w17357 & w17367) | (w17357 & w45000) | (w17367 & w45000);
assign w17377 = w16592 & w17372;
assign w17378 = ~w16722 & w17377;
assign w17379 = w17376 & ~w17378;
assign w17380 = (~w17379 & ~w41444) | (~w17379 & w47561) | (~w41444 & w47561);
assign w17381 = ~w17322 & ~w17329;
assign w17382 = (~w17328 & w17267) | (~w17328 & w41445) | (w17267 & w41445);
assign w17383 = ~w17275 & ~w17382;
assign w17384 = (w17381 & w17382) | (w17381 & w48905) | (w17382 & w48905);
assign w17385 = ~w17322 & ~w17384;
assign w17386 = ~w17313 & w17385;
assign w17387 = ~w17276 & w17337;
assign w17388 = ~w17386 & w17387;
assign w17389 = ~w17276 & w17299;
assign w17390 = ~w17336 & ~w17386;
assign w17391 = ~w17389 & ~w17390;
assign w17392 = w16555 & ~w17380;
assign w17393 = ~w17388 & ~w17391;
assign w17394 = w17380 & w17393;
assign w17395 = ~w17392 & ~w17394;
assign w17396 = ~w17140 & ~w17342;
assign w17397 = w17341 & w17396;
assign w17398 = (~w17140 & ~w17341) | (~w17140 & w41446) | (~w17341 & w41446);
assign w17399 = ~w9195 & w17398;
assign w17400 = w9195 & ~w17398;
assign w17401 = ~w17399 & ~w17400;
assign w17402 = ~w17379 & ~w17401;
assign w17403 = (w17159 & w17356) | (w17159 & w48906) | (w17356 & w48906);
assign w17404 = ~w17356 & w48907;
assign w17405 = ~w17403 & ~w17404;
assign w17406 = ~w8666 & w17405;
assign w17407 = ~w17341 & ~w17396;
assign w17408 = ~w17397 & ~w17407;
assign w17409 = w17139 & w17379;
assign w17410 = w16830 & w17139;
assign w17411 = w17355 & w17410;
assign w17412 = ~w17409 & ~w17411;
assign w17413 = ~w17379 & ~w17408;
assign w17414 = ~w17356 & w17413;
assign w17415 = w17412 & ~w17414;
assign w17416 = w17412 & w41447;
assign w17417 = w8666 & w17159;
assign w17418 = (w17417 & w17356) | (w17417 & w48908) | (w17356 & w48908);
assign w17419 = w8666 & ~w17159;
assign w17420 = ~w17356 & w48909;
assign w17421 = ~w17418 & ~w17420;
assign w17422 = ~w17416 & w17421;
assign w17423 = ~w17406 & ~w17422;
assign w17424 = ~w17119 & ~w17121;
assign w17425 = ~w17123 & w17183;
assign w17426 = ~w17140 & ~w17160;
assign w17427 = w9195 & ~w17159;
assign w17428 = ~w17184 & ~w17427;
assign w17429 = ~w17172 & ~w17428;
assign w17430 = ~w17172 & w17426;
assign w17431 = (w17430 & ~w17341) | (w17430 & w41448) | (~w17341 & w41448);
assign w17432 = ~w17429 & ~w17431;
assign w17433 = w17425 & w17432;
assign w17434 = ~w17425 & ~w17432;
assign w17435 = ~w17433 & ~w17434;
assign w17436 = w7315 & w17424;
assign w17437 = ~w17380 & w17436;
assign w17438 = w7315 & w17435;
assign w17439 = w17380 & w17438;
assign w17440 = ~w17437 & ~w17439;
assign w17441 = (~w17189 & ~w17341) | (~w17189 & w41449) | (~w17341 & w41449);
assign w17442 = ~w17087 & ~w17190;
assign w17443 = ~w17441 & w17442;
assign w17444 = ~w17345 & w41450;
assign w17445 = w17051 & w16830;
assign w17446 = ~w17444 & w17445;
assign w17447 = w16829 & ~w17062;
assign w17448 = ~w16723 & w17447;
assign w17449 = ~w17376 & ~w17448;
assign w17450 = ~w17446 & w17449;
assign w17451 = w17443 & w17450;
assign w17452 = w17441 & ~w17442;
assign w17453 = ~w17448 & w17452;
assign w17454 = ~w17379 & w17453;
assign w17455 = w17086 & w17443;
assign w17456 = w17086 & ~w17378;
assign w17457 = w17376 & w17456;
assign w17458 = ~w17455 & ~w17457;
assign w17459 = w16830 & w17086;
assign w17460 = w17355 & w17459;
assign w17461 = w17458 & ~w17460;
assign w17462 = ~w17446 & w17454;
assign w17463 = w17461 & ~w17462;
assign w17464 = (~w6769 & ~w17450) | (~w6769 & w41451) | (~w17450 & w41451);
assign w17465 = w17463 & w17464;
assign w17466 = w17440 & ~w17465;
assign w17467 = ~w17172 & ~w17184;
assign w17468 = (w17426 & ~w17341) | (w17426 & w48910) | (~w17341 & w48910);
assign w17469 = ~w17427 & ~w17468;
assign w17470 = w17467 & ~w17469;
assign w17471 = ~w17467 & w17469;
assign w17472 = ~w17470 & ~w17471;
assign w17473 = w17171 & ~w17380;
assign w17474 = w17380 & ~w17472;
assign w17475 = ~w17473 & ~w17474;
assign w17476 = w7924 & ~w17475;
assign w17477 = w17466 & ~w17476;
assign w17478 = ~w17423 & w17477;
assign w17479 = ~w17077 & ~w17078;
assign w17480 = (~w17190 & w17441) | (~w17190 & w48911) | (w17441 & w48911);
assign w17481 = w17479 & ~w17480;
assign w17482 = ~w17479 & w17480;
assign w17483 = ~w17481 & ~w17482;
assign w17484 = w17076 & ~w17380;
assign w17485 = w17380 & ~w17483;
assign w17486 = ~w17484 & ~w17485;
assign w17487 = ~w6264 & ~w17486;
assign w17488 = (~w17089 & ~w17441) | (~w17089 & w48912) | (~w17441 & w48912);
assign w17489 = w6264 & ~w17488;
assign w17490 = ~w6264 & w17488;
assign w17491 = ~w17489 & ~w17490;
assign w17492 = w17380 & ~w17491;
assign w17493 = ~w5745 & ~w17102;
assign w17494 = (w17493 & ~w17380) | (w17493 & w48913) | (~w17380 & w48913);
assign w17495 = ~w5745 & w17102;
assign w17496 = w17380 & w48914;
assign w17497 = ~w17494 & ~w17496;
assign w17498 = ~w17451 & w17463;
assign w17499 = (w6769 & ~w17463) | (w6769 & w41452) | (~w17463 & w41452);
assign w17500 = w5745 & w17102;
assign w17501 = (w17500 & ~w17380) | (w17500 & w48915) | (~w17380 & w48915);
assign w17502 = w5745 & ~w17102;
assign w17503 = w17380 & w48916;
assign w17504 = ~w17501 & ~w17503;
assign w17505 = ~w17499 & w17504;
assign w17506 = w17487 & w17497;
assign w17507 = w17505 & ~w17506;
assign w17508 = ~w17380 & w17424;
assign w17509 = w17380 & w17435;
assign w17510 = ~w17508 & ~w17509;
assign w17511 = ~w7315 & w17510;
assign w17512 = ~w7924 & w17475;
assign w17513 = ~w17511 & ~w17512;
assign w17514 = w17466 & ~w17513;
assign w17515 = ~w17478 & w41453;
assign w17516 = ~w16839 & ~w16879;
assign w17517 = (w16863 & ~w41454) | (w16863 & w47562) | (~w41454 & w47562);
assign w17518 = w17516 & ~w17517;
assign w17519 = ~w17516 & w17517;
assign w17520 = ~w17518 & ~w17519;
assign w17521 = w16838 & ~w17380;
assign w17522 = w17380 & w17520;
assign w17523 = ~w17521 & ~w17522;
assign w17524 = w4430 & w17523;
assign w17525 = ~w4430 & ~w17523;
assign w17526 = ~w17524 & ~w17525;
assign w17527 = w17349 & w17379;
assign w17528 = w16830 & w17349;
assign w17529 = w17355 & w17528;
assign w17530 = ~w17527 & ~w17529;
assign w17531 = w16863 & ~w17350;
assign w17532 = ~w17345 & w41455;
assign w17533 = (w17531 & w17345) | (w17531 & w41456) | (w17345 & w41456);
assign w17534 = ~w17532 & ~w17533;
assign w17535 = ~w17379 & w17534;
assign w17536 = ~w17356 & w17535;
assign w17537 = w17530 & ~w17536;
assign w17538 = (~w4838 & ~w17530) | (~w4838 & w41457) | (~w17530 & w41457);
assign w17539 = ~w17103 & ~w17107;
assign w17540 = ~w17089 & w17539;
assign w17541 = (w17191 & w17175) | (w17191 & w50344) | (w17175 & w50344);
assign w17542 = w17540 & w50203;
assign w17543 = ~w17093 & ~w17106;
assign w17544 = w17107 & ~w17543;
assign w17545 = ~w17107 & w17543;
assign w17546 = ~w17544 & ~w17545;
assign w17547 = w17542 & ~w17543;
assign w17548 = ~w17542 & ~w17546;
assign w17549 = ~w17547 & ~w17548;
assign w17550 = w5330 & ~w17092;
assign w17551 = ~w17380 & w17550;
assign w17552 = w5330 & ~w17549;
assign w17553 = w17380 & w17552;
assign w17554 = ~w17551 & ~w17553;
assign w17555 = w4838 & w17537;
assign w17556 = ~w17538 & w17554;
assign w17557 = ~w17555 & ~w17556;
assign w17558 = w17526 & w17557;
assign w17559 = ~w16890 & w17057;
assign w17560 = ~w16881 & ~w16882;
assign w17561 = (~w47563 & w48917) | (~w47563 & w48918) | (w48917 & w48918);
assign w17562 = (w47563 & w48919) | (w47563 & w48920) | (w48919 & w48920);
assign w17563 = ~w17561 & ~w17562;
assign w17564 = ~w16889 & ~w17380;
assign w17565 = w17380 & w17563;
assign w17566 = ~w17564 & ~w17565;
assign w17567 = ~w3646 & w17566;
assign w17568 = ~w16878 & ~w16882;
assign w17569 = ~w16864 & ~w16879;
assign w17570 = ~w16879 & ~w17350;
assign w17571 = (~w17569 & ~w41459) | (~w17569 & w47564) | (~w41459 & w47564);
assign w17572 = w17568 & ~w17571;
assign w17573 = ~w17568 & w17571;
assign w17574 = ~w17572 & ~w17573;
assign w17575 = w16877 & ~w17380;
assign w17576 = w17380 & w17574;
assign w17577 = ~w17575 & ~w17576;
assign w17578 = w4056 & w17577;
assign w17579 = ~w17524 & ~w17567;
assign w17580 = ~w17578 & w17579;
assign w17581 = w6264 & w17486;
assign w17582 = (w17497 & ~w17581) | (w17497 & w48921) | (~w17581 & w48921);
assign w17583 = ~w17558 & w47565;
assign w17584 = ~w17515 & w17583;
assign w17585 = a[44] & w16559;
assign w17586 = ~a[44] & ~w16559;
assign w17587 = ~w17585 & ~w17586;
assign w17588 = ~w17380 & w17587;
assign w17589 = a[44] & ~w17196;
assign w17590 = ~w17197 & ~w17589;
assign w17591 = ~w17379 & w17590;
assign w17592 = ~w17356 & w17591;
assign w17593 = (w15681 & w17356) | (w15681 & w47566) | (w17356 & w47566);
assign w17594 = ~w17588 & w17593;
assign w17595 = ~a[42] & w17380;
assign w17596 = ~a[40] & ~a[41];
assign w17597 = ~a[42] & w17596;
assign w17598 = w16559 & ~w17597;
assign w17599 = a[42] & w16559;
assign w17600 = ~w17378 & ~w17599;
assign w17601 = ~a[42] & w17598;
assign w17602 = ~a[43] & ~w17601;
assign w17603 = w17376 & ~w17600;
assign w17604 = w17602 & ~w17603;
assign w17605 = w41444 & w47567;
assign w17606 = w17604 & ~w17605;
assign w17607 = ~w16559 & w17597;
assign w17608 = ~w17196 & ~w17598;
assign w17609 = ~w15681 & w17590;
assign w17610 = ~w17608 & ~w17609;
assign w17611 = (~w17607 & w17356) | (~w17607 & w47568) | (w17356 & w47568);
assign w17612 = ~w15681 & w17587;
assign w17613 = ~w17380 & w17612;
assign w17614 = w17611 & ~w17613;
assign w17615 = ~w17595 & w17606;
assign w17616 = w17614 & ~w17615;
assign w17617 = (w14766 & w17616) | (w14766 & w48922) | (w17616 & w48922);
assign w17618 = ~w14766 & ~w17594;
assign w17619 = ~w17616 & w17618;
assign w17620 = a[45] & w17586;
assign w17621 = ~w17198 & ~w17199;
assign w17622 = ~w16559 & w17621;
assign w17623 = w16559 & ~w17621;
assign w17624 = ~w17622 & ~w17623;
assign w17625 = w15681 & ~w17196;
assign w17626 = ~a[44] & w17625;
assign w17627 = w17620 & w17625;
assign w17628 = ~a[45] & ~w17624;
assign w17629 = a[45] & ~w17626;
assign w17630 = w17624 & w17629;
assign w17631 = ~w17627 & ~w17630;
assign w17632 = ~w17628 & w17631;
assign w17633 = ~a[45] & ~w17586;
assign w17634 = w17380 & w17632;
assign w17635 = ~w17620 & ~w17633;
assign w17636 = ~w17380 & w17635;
assign w17637 = ~w17634 & ~w17636;
assign w17638 = ~w17619 & ~w17637;
assign w17639 = ~w17617 & ~w17638;
assign w17640 = ~w17381 & w17383;
assign w17641 = ~w17384 & ~w17640;
assign w17642 = w17051 & ~w17444;
assign w17643 = (w16609 & w17364) | (w16609 & w48882) | (w17364 & w48882);
assign w17644 = w17062 & w48923;
assign w17645 = ~w17642 & w17644;
assign w17646 = (w16830 & w17642) | (w16830 & w47569) | (w17642 & w47569);
assign w17647 = w17357 & ~w17372;
assign w17648 = w17641 & ~w17647;
assign w17649 = w11870 & w17648;
assign w17650 = ~w17646 & w17649;
assign w17651 = w11870 & w17321;
assign w17652 = (w17651 & w17356) | (w17651 & w47570) | (w17356 & w47570);
assign w17653 = ~w17650 & ~w17652;
assign w17654 = ~w13384 & w17268;
assign w17655 = w13384 & ~w17268;
assign w17656 = ~w17654 & ~w17655;
assign w17657 = ~w17379 & ~w17656;
assign w17658 = ~w17356 & w17657;
assign w17659 = w12666 & w17274;
assign w17660 = (w17659 & w17356) | (w17659 & w47571) | (w17356 & w47571);
assign w17661 = w12666 & ~w17274;
assign w17662 = ~w17356 & w47572;
assign w17663 = ~w17660 & ~w17662;
assign w17664 = w17653 & w17663;
assign w17665 = ~w17224 & ~w17266;
assign w17666 = (w17665 & ~w17376) | (w17665 & w48924) | (~w17376 & w48924);
assign w17667 = w13384 & ~w17264;
assign w17668 = (w17667 & w17356) | (w17667 & w47573) | (w17356 & w47573);
assign w17669 = w13384 & w17264;
assign w17670 = ~w17356 & w47574;
assign w17671 = ~w17668 & ~w17670;
assign w17672 = ~w12666 & ~w17274;
assign w17673 = (w17672 & w17356) | (w17672 & w47575) | (w17356 & w47575);
assign w17674 = ~w12666 & w17274;
assign w17675 = ~w17356 & w47576;
assign w17676 = ~w17673 & ~w17675;
assign w17677 = w17671 & w17676;
assign w17678 = (w17321 & w17356) | (w17321 & w47577) | (w17356 & w47577);
assign w17679 = ~w17646 & w17648;
assign w17680 = ~w17678 & ~w17679;
assign w17681 = ~w17678 & w48925;
assign w17682 = ~w17313 & ~w17336;
assign w17683 = w17385 & ~w17682;
assign w17684 = ~w17385 & w17682;
assign w17685 = ~w17683 & ~w17684;
assign w17686 = w17335 & ~w17380;
assign w17687 = w17380 & w17685;
assign w17688 = ~w17686 & ~w17687;
assign w17689 = w11138 & w17688;
assign w17690 = ~w17681 & ~w17689;
assign w17691 = w17664 & ~w17677;
assign w17692 = w17690 & ~w17691;
assign w17693 = w17209 & w17223;
assign w17694 = (w17217 & ~w17380) | (w17217 & w48926) | (~w17380 & w48926);
assign w17695 = w17380 & w48927;
assign w17696 = ~w17694 & ~w17695;
assign w17697 = ~w14039 & ~w17696;
assign w17698 = w17692 & ~w17697;
assign w17699 = w17639 & w17698;
assign w17700 = w14039 & w17696;
assign w17701 = (w17264 & w17356) | (w17264 & w47578) | (w17356 & w47578);
assign w17702 = ~w17356 & w47579;
assign w17703 = ~w17701 & ~w17702;
assign w17704 = ~w13384 & ~w17703;
assign w17705 = w17664 & ~w17704;
assign w17706 = ~w17700 & w17705;
assign w17707 = w17692 & ~w17706;
assign w17708 = ~w11138 & ~w17688;
assign w17709 = ~w17291 & ~w17333;
assign w17710 = w17276 & ~w17709;
assign w17711 = ~w17276 & w17709;
assign w17712 = ~w17710 & ~w17711;
assign w17713 = w17388 & ~w17709;
assign w17714 = ~w17388 & ~w17712;
assign w17715 = ~w17713 & ~w17714;
assign w17716 = w17332 & ~w17380;
assign w17717 = w17380 & ~w17715;
assign w17718 = ~w17716 & ~w17717;
assign w17719 = w9781 & ~w17718;
assign w17720 = w10419 & ~w17395;
assign w17721 = ~w17708 & ~w17719;
assign w17722 = ~w17720 & w17721;
assign w17723 = ~w17707 & w17722;
assign w17724 = ~w17699 & w17723;
assign w17725 = ~w9781 & w17718;
assign w17726 = ~w10419 & w17395;
assign w17727 = ~w17725 & ~w17726;
assign w17728 = ~w17719 & ~w17727;
assign w17729 = w9195 & ~w17415;
assign w17730 = ~w17406 & ~w17729;
assign w17731 = ~w17728 & w17730;
assign w17732 = w17507 & w17513;
assign w17733 = w17731 & w17732;
assign w17734 = ~w17724 & w17733;
assign w17735 = w17584 & ~w17734;
assign w17736 = ~w17043 & ~w17060;
assign w17737 = w17351 & ~w17736;
assign w17738 = ~w17345 & w41460;
assign w17739 = ~w16881 & w47580;
assign w17740 = ~w17736 & ~w17739;
assign w17741 = w17046 & ~w17740;
assign w17742 = ~w17738 & w17741;
assign w17743 = (~w16968 & w17738) | (~w16968 & w47581) | (w17738 & w47581);
assign w17744 = ~w16966 & ~w17736;
assign w17745 = w17351 & w17744;
assign w17746 = w17346 & w17745;
assign w17747 = ~w17739 & w17744;
assign w17748 = (w16949 & w17746) | (w16949 & w41461) | (w17746 & w41461);
assign w17749 = w17743 & ~w17748;
assign w17750 = w17380 & w17749;
assign w17751 = w41444 & w47582;
assign w17752 = w17062 & w17378;
assign w17753 = w17376 & ~w17752;
assign w17754 = ~w17746 & w41462;
assign w17755 = w50243 & w50345;
assign w17756 = ~w17754 & ~w17755;
assign w17757 = ~w17751 & w17756;
assign w17758 = ~w17750 & w17757;
assign w17759 = ~w2006 & w17758;
assign w17760 = (~w2558 & w17752) | (~w2558 & w45001) | (w17752 & w45001);
assign w17761 = (~w17044 & w17356) | (~w17044 & w47583) | (w17356 & w47583);
assign w17762 = (~w17747 & ~w17346) | (~w17747 & w41463) | (~w17346 & w41463);
assign w17763 = ~w17753 & w17762;
assign w17764 = ~w17356 & w17763;
assign w17765 = w17045 & ~w17740;
assign w17766 = ~w17738 & w17765;
assign w17767 = ~w17379 & w17766;
assign w17768 = w16966 & ~w17740;
assign w17769 = ~w17738 & w17768;
assign w17770 = ~w17356 & w17767;
assign w17771 = ~w17769 & ~w17770;
assign w17772 = ~w17761 & ~w17764;
assign w17773 = w17771 & ~w17772;
assign w17774 = ~w2285 & w17773;
assign w17775 = ~w17759 & ~w17774;
assign w17776 = (w17042 & w17752) | (w17042 & w45002) | (w17752 & w45002);
assign w17777 = (~w17029 & w17356) | (~w17029 & w47584) | (w17356 & w47584);
assign w17778 = ~w16998 & ~w17058;
assign w17779 = ~w16881 & w48928;
assign w17780 = (~w47585 & w48929) | (~w47585 & w48930) | (w48929 & w48930);
assign w17781 = w17038 & ~w17780;
assign w17782 = w17014 & ~w17781;
assign w17783 = ~w17777 & w17782;
assign w17784 = ~w17042 & ~w17740;
assign w17785 = ~w17738 & w17784;
assign w17786 = ~w17379 & w17785;
assign w17787 = ~w17028 & w17379;
assign w17788 = w16830 & ~w17028;
assign w17789 = w17355 & w17788;
assign w17790 = ~w17787 & ~w17789;
assign w17791 = ~w17356 & w17786;
assign w17792 = w17790 & ~w17791;
assign w17793 = w17790 & w41464;
assign w17794 = ~w17783 & w17793;
assign w17795 = (w2285 & w17770) | (w2285 & w47586) | (w17770 & w47586);
assign w17796 = (w2285 & ~w17763) | (w2285 & w45003) | (~w17763 & w45003);
assign w17797 = ~w17761 & w17796;
assign w17798 = ~w17795 & ~w17797;
assign w17799 = ~w17794 & w17798;
assign w17800 = ~w17379 & ~w17446;
assign w17801 = ~w17002 & ~w17004;
assign w17802 = w17005 & ~w17801;
assign w17803 = ~w17005 & w17801;
assign w17804 = ~w17802 & ~w17803;
assign w17805 = w17380 & ~w17781;
assign w17806 = (w17804 & ~w17800) | (w17804 & w41465) | (~w17800 & w41465);
assign w17807 = ~w17805 & ~w17806;
assign w17808 = (~w17753 & ~w41444) | (~w17753 & w48931) | (~w41444 & w48931);
assign w17809 = ~w17038 & w17780;
assign w17810 = (~w47585 & w48932) | (~w47585 & w48933) | (w48932 & w48933);
assign w17811 = (~w17809 & w17356) | (~w17809 & w48934) | (w17356 & w48934);
assign w17812 = ~w17807 & w17811;
assign w17813 = (~w2896 & w17807) | (~w2896 & w48935) | (w17807 & w48935);
assign w17814 = ~w17783 & w17792;
assign w17815 = w2558 & ~w17814;
assign w17816 = ~w17813 & ~w17815;
assign w17817 = w17799 & ~w17816;
assign w17818 = w17775 & ~w17817;
assign w17819 = ~w16712 & ~w17361;
assign w17820 = (w17819 & w17354) | (w17819 & w41466) | (w17354 & w41466);
assign w17821 = ~w17354 & w45005;
assign w17822 = ~w17820 & ~w17821;
assign w17823 = ~w16709 & ~w16710;
assign w17824 = ~w17380 & w17823;
assign w17825 = w17380 & w17822;
assign w17826 = ~w17824 & ~w17825;
assign w17827 = w1320 & w17826;
assign w17828 = ~w17062 & w17376;
assign w17829 = ~w16969 & ~w16972;
assign w17830 = (w17829 & ~w17376) | (w17829 & w45006) | (~w17376 & w45006);
assign w17831 = ~w17738 & w47588;
assign w17832 = w17830 & ~w17831;
assign w17833 = (~w1738 & w17356) | (~w1738 & w47589) | (w17356 & w47589);
assign w17834 = w17380 & w17832;
assign w17835 = ~w17833 & ~w17834;
assign w17836 = w16900 & w16977;
assign w17837 = w1541 & w17836;
assign w17838 = ~w17835 & w17837;
assign w17839 = w1541 & ~w17836;
assign w17840 = w17835 & w17839;
assign w17841 = ~w17838 & ~w17840;
assign w17842 = ~w17827 & w17841;
assign w17843 = ~w1320 & ~w17826;
assign w17844 = w16693 & ~w16696;
assign w17845 = ~w16693 & w16696;
assign w17846 = ~w17844 & ~w17845;
assign w17847 = w1320 & ~w16712;
assign w17848 = ~w1320 & w16712;
assign w17849 = ~w17847 & ~w17848;
assign w17850 = (w41466 & w47590) | (w41466 & w47591) | (w47590 & w47591);
assign w17851 = (~w41466 & w47592) | (~w41466 & w47593) | (w47592 & w47593);
assign w17852 = ~w17850 & ~w17851;
assign w17853 = ~w17356 & w47594;
assign w17854 = ~w17852 & w17853;
assign w17855 = w17853 & w48936;
assign w17856 = w1120 & ~w17846;
assign w17857 = (w17856 & w17852) | (w17856 & w45007) | (w17852 & w45007);
assign w17858 = ~w17855 & ~w17857;
assign w17859 = ~w17843 & w17858;
assign w17860 = ~w17842 & w17859;
assign w17861 = w2006 & ~w17758;
assign w17862 = w16931 & ~w16972;
assign w17863 = ~w17742 & w45008;
assign w17864 = w17808 & ~w17863;
assign w17865 = ~w16919 & ~w16970;
assign w17866 = (w17865 & w17356) | (w17865 & w47595) | (w17356 & w47595);
assign w17867 = ~w17864 & ~w17866;
assign w17868 = (~w2006 & w17448) | (~w2006 & w41467) | (w17448 & w41467);
assign w17869 = ~w16723 & w45009;
assign w17870 = w17642 & w17869;
assign w17871 = ~w17868 & ~w17870;
assign w17872 = (w17862 & w17742) | (w17862 & w45010) | (w17742 & w45010);
assign w17873 = w17871 & w17872;
assign w17874 = (w1738 & ~w17871) | (w1738 & w45011) | (~w17871 & w45011);
assign w17875 = ~w17867 & w17874;
assign w17876 = ~w17861 & ~w17875;
assign w17877 = (w17876 & w17842) | (w17876 & w48937) | (w17842 & w48937);
assign w17878 = ~w17818 & w17877;
assign w17879 = ~w17867 & ~w17873;
assign w17880 = (~w1738 & w17867) | (~w1738 & w45012) | (w17867 & w45012);
assign w17881 = ~w1541 & ~w17836;
assign w17882 = ~w17835 & w17881;
assign w17883 = ~w1541 & w17836;
assign w17884 = w17835 & w17883;
assign w17885 = ~w17882 & ~w17884;
assign w17886 = ~w17880 & w17885;
assign w17887 = w17859 & w17886;
assign w17888 = ~w17860 & ~w17887;
assign w17889 = (~w17092 & w17356) | (~w17092 & w45013) | (w17356 & w45013);
assign w17890 = w17380 & ~w17549;
assign w17891 = ~w17889 & ~w17890;
assign w17892 = ~w17890 & w45014;
assign w17893 = ~w17538 & w17892;
assign w17894 = ~w17525 & ~w17555;
assign w17895 = ~w17893 & w17894;
assign w17896 = w17580 & ~w17895;
assign w17897 = ~w16998 & ~w17052;
assign w17898 = w16892 & ~w17444;
assign w17899 = w17057 & ~w17898;
assign w17900 = ~w17897 & w17899;
assign w17901 = w17897 & ~w17899;
assign w17902 = ~w16997 & ~w17380;
assign w17903 = w17380 & ~w17900;
assign w17904 = ~w17901 & w17903;
assign w17905 = ~w17902 & ~w17904;
assign w17906 = w3646 & ~w17566;
assign w17907 = ~w4056 & ~w17577;
assign w17908 = ~w17567 & w17907;
assign w17909 = ~w17906 & ~w17908;
assign w17910 = w3242 & w17905;
assign w17911 = w17909 & ~w17910;
assign w17912 = ~w17896 & w17911;
assign w17913 = ~w17888 & w17912;
assign w17914 = ~w17878 & w17913;
assign w17915 = ~w17735 & w17914;
assign w17916 = ~w16797 & w17380;
assign w17917 = w42 & ~w16782;
assign w17918 = ~w17370 & w17645;
assign w17919 = ~w16723 & w16827;
assign w17920 = ~w17370 & ~w17919;
assign w17921 = ~w16775 & ~w17920;
assign w17922 = (w17369 & w17918) | (w17369 & w45015) | (w17918 & w45015);
assign w17923 = w16735 & ~w17922;
assign w17924 = ~w17916 & w17917;
assign w17925 = ~w3 & w17917;
assign w17926 = w17923 & w17925;
assign w17927 = ~w17924 & ~w17926;
assign w17928 = w3 & ~w17923;
assign w17929 = w16797 & w17380;
assign w17930 = ~w17928 & w17929;
assign w17931 = ~w17927 & ~w17930;
assign w17932 = w42 & w16782;
assign w17933 = w17808 & w17932;
assign w17934 = ~w3 & w16797;
assign w17935 = w17933 & w17934;
assign w17936 = ~w17923 & w17935;
assign w17937 = w3 & w16797;
assign w17938 = w17933 & w17937;
assign w17939 = w17923 & w17938;
assign w17940 = ~w17936 & ~w17939;
assign w17941 = ~w16755 & ~w16783;
assign w17942 = ~w16783 & w17369;
assign w17943 = (w17942 & w17918) | (w17942 & w45016) | (w17918 & w45016);
assign w17944 = ~w17941 & ~w17943;
assign w17945 = ~w16486 & w16803;
assign w17946 = w16486 & ~w16503;
assign w17947 = ~w16803 & w17946;
assign w17948 = ~w17945 & ~w17947;
assign w17949 = ~w42 & w17948;
assign w17950 = w16797 & ~w17949;
assign w17951 = w16798 & w17944;
assign w17952 = ~w42 & ~w17950;
assign w17953 = ~w17944 & w17952;
assign w17954 = ~w17951 & ~w17953;
assign w17955 = w17940 & w17954;
assign w17956 = ~w17931 & w17955;
assign w17957 = ~w3 & w17380;
assign w17958 = ~w17923 & w17957;
assign w17959 = w3 & w17380;
assign w17960 = w17923 & w17959;
assign w17961 = ~w17958 & ~w17960;
assign w17962 = (~w17368 & w17918) | (~w17368 & w45017) | (w17918 & w45017);
assign w17963 = w16735 & w16780;
assign w17964 = w16729 & ~w16730;
assign w17965 = ~w16729 & w16730;
assign w17966 = ~w17964 & ~w17965;
assign w17967 = ~w17808 & ~w17966;
assign w17968 = w17380 & ~w17963;
assign w17969 = ~w17962 & w17968;
assign w17970 = w17380 & w17963;
assign w17971 = w17962 & w17970;
assign w17972 = ~w17969 & ~w17971;
assign w17973 = ~w17967 & w17972;
assign w17974 = ~w3 & ~w17973;
assign w17975 = ~w42 & ~w16782;
assign w17976 = w17961 & w17975;
assign w17977 = ~w42 & w16782;
assign w17978 = ~w17961 & w17977;
assign w17979 = ~w17974 & ~w17978;
assign w17980 = ~w17976 & w17979;
assign w17981 = (~w16825 & ~w17450) | (~w16825 & w45018) | (~w17450 & w45018);
assign w17982 = ~w16723 & ~w16826;
assign w17983 = ~w17645 & w17982;
assign w17984 = ~w17981 & ~w17983;
assign w17985 = ~w17367 & ~w17919;
assign w17986 = ~w17645 & ~w17985;
assign w17987 = w17808 & ~w17986;
assign w17988 = ~w16824 & ~w17987;
assign w17989 = w17380 & w17986;
assign w17990 = w252 & w17989;
assign w17991 = ~w17988 & ~w17990;
assign w17992 = ~w17984 & w17991;
assign w17993 = ~w17356 & w45019;
assign w17994 = (w17365 & w17354) | (w17365 & w41468) | (w17354 & w41468);
assign w17995 = w16722 & ~w17994;
assign w17996 = (~w17643 & w17994) | (~w17643 & w45020) | (w17994 & w45020);
assign w17997 = w17993 & w17996;
assign w17998 = ~w351 & ~w17380;
assign w17999 = ~w16591 & ~w16826;
assign w18000 = w252 & ~w17999;
assign w18001 = (w18000 & w17997) | (w18000 & w48938) | (w17997 & w48938);
assign w18002 = w252 & w17999;
assign w18003 = ~w17997 & w48939;
assign w18004 = ~w18001 & ~w18003;
assign w18005 = (w57 & ~w17991) | (w57 & w45021) | (~w17991 & w45021);
assign w18006 = w18004 & ~w18005;
assign w18007 = ~w252 & w17999;
assign w18008 = (w18007 & w17997) | (w18007 & w48940) | (w17997 & w48940);
assign w18009 = ~w252 & ~w17999;
assign w18010 = ~w17997 & w48941;
assign w18011 = ~w18008 & ~w18010;
assign w18012 = w17993 & w17995;
assign w18013 = ~w16604 & ~w16721;
assign w18014 = ~w17994 & w18013;
assign w18015 = w17808 & ~w18014;
assign w18016 = w16578 & w18015;
assign w18017 = ~w16575 & ~w16576;
assign w18018 = ~w17380 & ~w18017;
assign w18019 = ~w16608 & ~w18014;
assign w18020 = ~w18018 & ~w18019;
assign w18021 = ~w18012 & ~w18016;
assign w18022 = w18020 & w18021;
assign w18023 = w18021 & w45022;
assign w18024 = w18011 & ~w18023;
assign w18025 = (~w17920 & ~w17645) | (~w17920 & w45023) | (~w17645 & w45023);
assign w18026 = ~w57 & w18025;
assign w18027 = w17808 & ~w18026;
assign w18028 = w57 & ~w18025;
assign w18029 = w16774 & ~w18028;
assign w18030 = w18027 & w18029;
assign w18031 = ~w17367 & w18028;
assign w18032 = w18027 & ~w18031;
assign w18033 = w80 & w18030;
assign w18034 = w80 & ~w16774;
assign w18035 = ~w18032 & w18034;
assign w18036 = ~w18033 & ~w18035;
assign w18037 = ~w57 & w17992;
assign w18038 = w18036 & ~w18037;
assign w18039 = w18006 & ~w18024;
assign w18040 = w18038 & ~w18039;
assign w18041 = w3 & w17973;
assign w18042 = ~w80 & ~w18030;
assign w18043 = ~w16774 & ~w18032;
assign w18044 = w18042 & ~w18043;
assign w18045 = ~w18041 & ~w18044;
assign w18046 = ~w17956 & w18045;
assign w18047 = ~w17956 & ~w17980;
assign w18048 = ~w18040 & w18046;
assign w18049 = ~w18047 & ~w18048;
assign w18050 = w17799 & w17876;
assign w18051 = ~w3242 & ~w17905;
assign w18052 = w2896 & w17812;
assign w18053 = ~w18051 & ~w18052;
assign w18054 = w18050 & w48942;
assign w18055 = ~w17888 & ~w18054;
assign w18056 = ~w17878 & w18055;
assign w18057 = ~w17061 & w41469;
assign w18058 = w16680 & ~w16719;
assign w18059 = w18057 & w18058;
assign w18060 = ~w945 & w18058;
assign w18061 = w945 & ~w18058;
assign w18062 = ~w18060 & ~w18061;
assign w18063 = ~w18059 & w18062;
assign w18064 = w17051 & w18062;
assign w18065 = ~w17444 & w18064;
assign w18066 = ~w18063 & ~w18065;
assign w18067 = ~w945 & w18059;
assign w18068 = ~w17642 & w18067;
assign w18069 = w18066 & ~w18068;
assign w18070 = (w16655 & w18069) | (w16655 & w48943) | (w18069 & w48943);
assign w18071 = ~w16681 & w18058;
assign w18072 = ~w16656 & ~w18071;
assign w18073 = ~w16656 & w18057;
assign w18074 = ~w17642 & w18073;
assign w18075 = ~w18072 & ~w18074;
assign w18076 = ~w18069 & w18084;
assign w18077 = ~w18070 & ~w18076;
assign w18078 = w754 & w18077;
assign w18079 = w16660 & ~w17448;
assign w18080 = (~w16636 & ~w17800) | (~w16636 & w41470) | (~w17800 & w41470);
assign w18081 = ~w16657 & ~w16658;
assign w18082 = ~w754 & w18081;
assign w18083 = ~w18075 & ~w18080;
assign w18084 = w17808 & w18075;
assign w18085 = w18082 & w18084;
assign w18086 = ~w18083 & ~w18085;
assign w18087 = ~w16636 & ~w17379;
assign w18088 = ~w17356 & w18087;
assign w18089 = w16661 & w18057;
assign w18090 = ~w17642 & w18089;
assign w18091 = ~w18072 & ~w18081;
assign w18092 = ~w18090 & w18091;
assign w18093 = w18088 & w18092;
assign w18094 = ~w17808 & ~w18081;
assign w18095 = ~w18093 & ~w18094;
assign w18096 = ~w18093 & w48944;
assign w18097 = w18086 & w18096;
assign w18098 = ~w18078 & ~w18097;
assign w18099 = w18086 & w18095;
assign w18100 = ~w612 & ~w18099;
assign w18101 = ~w18098 & ~w18100;
assign w18102 = (~w16680 & w17752) | (~w16680 & w45024) | (w17752 & w45024);
assign w18103 = (w16692 & w17356) | (w16692 & w48945) | (w17356 & w48945);
assign w18104 = (~w17361 & w17354) | (~w17361 & w41471) | (w17354 & w41471);
assign w18105 = w16718 & ~w18104;
assign w18106 = w16701 & ~w18105;
assign w18107 = ~w18103 & ~w18106;
assign w18108 = w16680 & w16702;
assign w18109 = (w18108 & ~w17447) | (w18108 & w41472) | (~w17447 & w41472);
assign w18110 = ~w17379 & w18109;
assign w18111 = ~w17446 & w18110;
assign w18112 = w1320 & w16559;
assign w18113 = ~w16670 & ~w18112;
assign w18114 = w16671 & ~w18113;
assign w18115 = ~w16671 & w18113;
assign w18116 = ~w18114 & ~w18115;
assign w18117 = ~w18105 & w18111;
assign w18118 = (w18116 & w17356) | (w18116 & w41473) | (w17356 & w41473);
assign w18119 = ~w18117 & ~w18118;
assign w18120 = ~w18107 & w18119;
assign w18121 = ~w945 & ~w18120;
assign w18122 = (~w17846 & w17852) | (~w17846 & w41474) | (w17852 & w41474);
assign w18123 = ~w1120 & ~w17854;
assign w18124 = ~w18122 & w18123;
assign w18125 = ~w18121 & ~w18124;
assign w18126 = ~w16660 & w18072;
assign w18127 = (~w18126 & w17642) | (~w18126 & w41475) | (w17642 & w41475);
assign w18128 = (w612 & w17356) | (w612 & w41476) | (w17356 & w41476);
assign w18129 = w18088 & w18127;
assign w18130 = ~w18128 & ~w18129;
assign w18131 = ~w16616 & ~w16663;
assign w18132 = w493 & ~w18131;
assign w18133 = (w18132 & w18129) | (w18132 & w41477) | (w18129 & w41477);
assign w18134 = w493 & w18131;
assign w18135 = ~w18129 & w41478;
assign w18136 = ~w18133 & ~w18135;
assign w18137 = ~w16662 & ~w16663;
assign w18138 = ~w16720 & w18137;
assign w18139 = w18057 & w18137;
assign w18140 = (~w18138 & w17642) | (~w18138 & w41479) | (w17642 & w41479);
assign w18141 = ~w493 & ~w18140;
assign w18142 = w493 & ~w18138;
assign w18143 = (w18142 & w17642) | (w18142 & w41480) | (w17642 & w41480);
assign w18144 = w17380 & ~w18143;
assign w18145 = ~w18141 & w18144;
assign w18146 = w493 & w17828;
assign w18147 = w16603 & ~w18146;
assign w18148 = ~w400 & w16603;
assign w18149 = (w18148 & ~w18144) | (w18148 & w41481) | (~w18144 & w41481);
assign w18150 = ~w400 & ~w18147;
assign w18151 = w18145 & w18150;
assign w18152 = ~w18149 & ~w18151;
assign w18153 = w18136 & w18152;
assign w18154 = w18125 & w18153;
assign w18155 = ~w18101 & w18154;
assign w18156 = (w18155 & ~w18055) | (w18155 & w47596) | (~w18055 & w47596);
assign w18157 = w18049 & w18156;
assign w18158 = ~w17915 & w18157;
assign w18159 = w400 & ~w16603;
assign w18160 = (w18159 & ~w18144) | (w18159 & w41482) | (~w18144 & w41482);
assign w18161 = w400 & w18147;
assign w18162 = w18145 & w18161;
assign w18163 = ~w18160 & ~w18162;
assign w18164 = ~w18153 & w18163;
assign w18165 = (~w351 & ~w18021) | (~w351 & w41483) | (~w18021 & w41483);
assign w18166 = ~w18153 & w41484;
assign w18167 = ~w493 & ~w18131;
assign w18168 = ~w18129 & w41485;
assign w18169 = ~w493 & w18131;
assign w18170 = (w18169 & w18129) | (w18169 & w41486) | (w18129 & w41486);
assign w18171 = ~w18168 & ~w18170;
assign w18172 = w18163 & w18171;
assign w18173 = ~w18165 & w18172;
assign w18174 = w945 & w18120;
assign w18175 = ~w754 & ~w18077;
assign w18176 = ~w18174 & ~w18175;
assign w18177 = ~w18100 & w18176;
assign w18178 = ~w18101 & ~w18177;
assign w18179 = (~w18166 & w18178) | (~w18166 & w41487) | (w18178 & w41487);
assign w18180 = w18006 & w18046;
assign w18181 = ~w18179 & w18180;
assign w18182 = w18049 & ~w18181;
assign w18183 = ~w18158 & ~w18182;
assign w18184 = ~w17720 & ~w17726;
assign w18185 = ~w17707 & ~w17708;
assign w18186 = ~w17699 & w18185;
assign w18187 = w18184 & ~w18186;
assign w18188 = ~w18184 & w18186;
assign w18189 = ~w18187 & ~w18188;
assign w18190 = ~w18158 & w41488;
assign w18191 = (w18189 & w18158) | (w18189 & w41489) | (w18158 & w41489);
assign w18192 = ~w18190 & ~w18191;
assign w18193 = ~w17689 & ~w17708;
assign w18194 = ~w17697 & ~w17700;
assign w18195 = ~w17639 & w18194;
assign w18196 = (~w17697 & w17639) | (~w17697 & w41490) | (w17639 & w41490);
assign w18197 = ~w17704 & ~w18196;
assign w18198 = w17677 & ~w18197;
assign w18199 = w17664 & ~w17681;
assign w18200 = ~w18198 & w18199;
assign w18201 = w17681 & ~w18193;
assign w18202 = ~w17681 & w18193;
assign w18203 = ~w18201 & ~w18202;
assign w18204 = ~w18193 & w18200;
assign w18205 = ~w18200 & ~w18203;
assign w18206 = ~w18204 & ~w18205;
assign w18207 = ~w18158 & w41491;
assign w18208 = ~w18183 & w18206;
assign w18209 = ~w18207 & ~w18208;
assign w18210 = (w10419 & w18208) | (w10419 & w41492) | (w18208 & w41492);
assign w18211 = w9781 & ~w18192;
assign w18212 = ~w18210 & ~w18211;
assign w18213 = w17653 & ~w17681;
assign w18214 = w17663 & ~w18198;
assign w18215 = ~w18213 & ~w18214;
assign w18216 = ~w18158 & w41493;
assign w18217 = ~w18200 & ~w18215;
assign w18218 = ~w18183 & w18217;
assign w18219 = ~w18216 & ~w18218;
assign w18220 = (w11138 & w18218) | (w11138 & w41494) | (w18218 & w41494);
assign w18221 = ~w18208 & w41495;
assign w18222 = ~w18220 & ~w18221;
assign w18223 = w18212 & ~w18222;
assign w18224 = ~w9781 & w18192;
assign w18225 = ~w18223 & ~w18224;
assign w18226 = ~w17724 & ~w17728;
assign w18227 = ~w17416 & ~w17729;
assign w18228 = w18226 & ~w18227;
assign w18229 = ~w18226 & w18227;
assign w18230 = ~w18228 & ~w18229;
assign w18231 = w8666 & w17415;
assign w18232 = ~w18158 & w41496;
assign w18233 = w8666 & ~w18230;
assign w18234 = ~w18183 & w18233;
assign w18235 = ~w18232 & ~w18234;
assign w18236 = w8666 & ~w17405;
assign w18237 = ~w17406 & ~w18236;
assign w18238 = ~w17728 & ~w17729;
assign w18239 = (~w17416 & w17724) | (~w17416 & w41497) | (w17724 & w41497);
assign w18240 = w18237 & ~w18239;
assign w18241 = ~w18237 & w18239;
assign w18242 = ~w18240 & ~w18241;
assign w18243 = w7924 & ~w17405;
assign w18244 = ~w18158 & w41498;
assign w18245 = w7924 & w18242;
assign w18246 = ~w18183 & w18245;
assign w18247 = ~w18244 & ~w18246;
assign w18248 = w18235 & w18247;
assign w18249 = ~w17719 & ~w17725;
assign w18250 = (~w17720 & w18186) | (~w17720 & w41499) | (w18186 & w41499);
assign w18251 = w18249 & ~w18250;
assign w18252 = ~w18249 & w18250;
assign w18253 = ~w18251 & ~w18252;
assign w18254 = w9195 & w17718;
assign w18255 = ~w18158 & w41500;
assign w18256 = w9195 & ~w18253;
assign w18257 = ~w18183 & w18256;
assign w18258 = ~w18255 & ~w18257;
assign w18259 = ~w8666 & ~w17415;
assign w18260 = ~w18158 & w41501;
assign w18261 = ~w8666 & w18230;
assign w18262 = ~w18183 & w18261;
assign w18263 = ~w18260 & ~w18262;
assign w18264 = w18258 & w18263;
assign w18265 = (~w7924 & w18158) | (~w7924 & w45025) | (w18158 & w45025);
assign w18266 = ~w18183 & w18242;
assign w18267 = w18265 & ~w18266;
assign w18268 = ~w17476 & ~w17512;
assign w18269 = (~w17423 & w17724) | (~w17423 & w41503) | (w17724 & w41503);
assign w18270 = w18268 & ~w18269;
assign w18271 = ~w18268 & w18269;
assign w18272 = ~w18270 & ~w18271;
assign w18273 = (~w7315 & w18158) | (~w7315 & w45026) | (w18158 & w45026);
assign w18274 = ~w18183 & w18272;
assign w18275 = w18273 & ~w18274;
assign w18276 = ~w18267 & ~w18275;
assign w18277 = w18248 & ~w18264;
assign w18278 = w18276 & ~w18277;
assign w18279 = ~w18158 & w41505;
assign w18280 = (w18269 & w18158) | (w18269 & w41506) | (w18158 & w41506);
assign w18281 = ~w18279 & ~w18280;
assign w18282 = w7315 & ~w18268;
assign w18283 = w18281 & w18282;
assign w18284 = w7315 & w18268;
assign w18285 = ~w18281 & w18284;
assign w18286 = ~w18283 & ~w18285;
assign w18287 = (w18286 & w18277) | (w18286 & w41507) | (w18277 & w41507);
assign w18288 = w18225 & ~w18287;
assign w18289 = w17718 & w18183;
assign w18290 = ~w18183 & ~w18253;
assign w18291 = ~w18289 & ~w18290;
assign w18292 = ~w9195 & w18291;
assign w18293 = w18248 & ~w18292;
assign w18294 = w18278 & ~w18293;
assign w18295 = ~w17526 & ~w17557;
assign w18296 = ~w17558 & ~w18295;
assign w18297 = ~w17515 & w17582;
assign w18298 = w17554 & ~w17892;
assign w18299 = ~w17538 & ~w17555;
assign w18300 = w18298 & w18299;
assign w18301 = (w18300 & w17734) | (w18300 & w41508) | (w17734 & w41508);
assign w18302 = w18296 & ~w18301;
assign w18303 = ~w18296 & w18301;
assign w18304 = ~w18302 & ~w18303;
assign w18305 = ~w18158 & w41509;
assign w18306 = ~w18183 & ~w18304;
assign w18307 = ~w18305 & ~w18306;
assign w18308 = (w4056 & w18306) | (w4056 & w41510) | (w18306 & w41510);
assign w18309 = (w18298 & w17515) | (w18298 & w41511) | (w17515 & w41511);
assign w18310 = w17733 & w18298;
assign w18311 = ~w17724 & w18310;
assign w18312 = ~w18309 & ~w18311;
assign w18313 = w18297 & ~w18298;
assign w18314 = ~w17734 & w18313;
assign w18315 = w18312 & ~w18314;
assign w18316 = ~w4838 & ~w17891;
assign w18317 = ~w18158 & w41512;
assign w18318 = ~w4838 & w18315;
assign w18319 = ~w18183 & w18318;
assign w18320 = ~w18317 & ~w18319;
assign w18321 = ~w17554 & ~w18299;
assign w18322 = w17554 & w18299;
assign w18323 = ~w18321 & ~w18322;
assign w18324 = ~w18311 & w41513;
assign w18325 = ~w18301 & ~w18324;
assign w18326 = w4430 & ~w17537;
assign w18327 = ~w18158 & w41514;
assign w18328 = w4430 & w18325;
assign w18329 = ~w18183 & w18328;
assign w18330 = ~w18327 & ~w18329;
assign w18331 = w18320 & w18330;
assign w18332 = ~w18308 & w18331;
assign w18333 = ~w17487 & ~w17581;
assign w18334 = ~w17499 & ~w17514;
assign w18335 = ~w17478 & w18334;
assign w18336 = w17731 & w18334;
assign w18337 = w18333 & w18335;
assign w18338 = w18333 & w18336;
assign w18339 = ~w17724 & w18338;
assign w18340 = ~w18337 & ~w18339;
assign w18341 = ~w18339 & w41515;
assign w18342 = w17497 & w17504;
assign w18343 = w18341 & ~w18342;
assign w18344 = ~w18341 & w18342;
assign w18345 = ~w18343 & ~w18344;
assign w18346 = w17102 & ~w17492;
assign w18347 = ~w17102 & w17492;
assign w18348 = ~w18346 & ~w18347;
assign w18349 = (~w5330 & w18158) | (~w5330 & w45027) | (w18158 & w45027);
assign w18350 = ~w18183 & w18345;
assign w18351 = w18349 & ~w18350;
assign w18352 = ~w17724 & w18336;
assign w18353 = ~w18333 & ~w18335;
assign w18354 = ~w18352 & w18353;
assign w18355 = w18340 & ~w18354;
assign w18356 = ~w5745 & w17486;
assign w18357 = ~w18158 & w41516;
assign w18358 = ~w5745 & w18355;
assign w18359 = ~w18183 & w18358;
assign w18360 = ~w18357 & ~w18359;
assign w18361 = ~w18351 & ~w18360;
assign w18362 = ~w18182 & ~w18348;
assign w18363 = (w5330 & w18158) | (w5330 & w45028) | (w18158 & w45028);
assign w18364 = ~w18183 & ~w18345;
assign w18365 = w18363 & ~w18364;
assign w18366 = w17440 & ~w17511;
assign w18367 = ~w17423 & w18268;
assign w18368 = w18366 & w18367;
assign w18369 = (w18368 & w17724) | (w18368 & w41517) | (w17724 & w41517);
assign w18370 = ~w6769 & w17498;
assign w18371 = ~w17499 & ~w18370;
assign w18372 = w17440 & ~w17513;
assign w18373 = w18371 & ~w18372;
assign w18374 = ~w18371 & w18372;
assign w18375 = ~w18373 & ~w18374;
assign w18376 = w18369 & w18371;
assign w18377 = ~w18369 & w18375;
assign w18378 = ~w18376 & ~w18377;
assign w18379 = w6264 & w17498;
assign w18380 = ~w18158 & w41518;
assign w18381 = w6264 & ~w18378;
assign w18382 = ~w18183 & w18381;
assign w18383 = ~w18380 & ~w18382;
assign w18384 = ~w18365 & w18383;
assign w18385 = ~w18361 & w18384;
assign w18386 = w18332 & w18385;
assign w18387 = ~w17476 & ~w18270;
assign w18388 = w18366 & ~w18387;
assign w18389 = ~w18366 & w18387;
assign w18390 = ~w18388 & ~w18389;
assign w18391 = ~w18158 & w45029;
assign w18392 = ~w18183 & ~w18390;
assign w18393 = ~w18391 & ~w18392;
assign w18394 = ~w18392 & w45030;
assign w18395 = w18286 & ~w18394;
assign w18396 = w18386 & w18395;
assign w18397 = ~w18294 & w18396;
assign w18398 = ~a[38] & ~a[39];
assign w18399 = ~a[40] & w18398;
assign w18400 = ~w17380 & ~w18399;
assign w18401 = a[41] & w18400;
assign w18402 = ~w17596 & ~w18401;
assign w18403 = (w18402 & w18158) | (w18402 & w41519) | (w18158 & w41519);
assign w18404 = ~a[41] & ~w18400;
assign w18405 = ~w18182 & w18404;
assign w18406 = w17380 & w18399;
assign w18407 = (~w18406 & w18158) | (~w18406 & w45031) | (w18158 & w45031);
assign w18408 = (~w16559 & ~w18407) | (~w16559 & w41520) | (~w18407 & w41520);
assign w18409 = w16559 & ~w18406;
assign w18410 = (w18409 & w18158) | (w18409 & w45032) | (w18158 & w45032);
assign w18411 = ~w18403 & w18410;
assign w18412 = a[42] & ~w17380;
assign w18413 = a[42] & ~w17596;
assign w18414 = ~w17597 & ~w18413;
assign w18415 = ~w17595 & ~w18412;
assign w18416 = ~w18158 & w41521;
assign w18417 = (w18414 & w18158) | (w18414 & w41522) | (w18158 & w41522);
assign w18418 = ~w18416 & ~w18417;
assign w18419 = ~w18411 & ~w18418;
assign w18420 = ~w18408 & ~w18419;
assign w18421 = ~w18419 & w41523;
assign w18422 = ~a[43] & ~w17598;
assign w18423 = ~w17380 & ~w18422;
assign w18424 = ~a[43] & ~w17595;
assign w18425 = ~w17608 & ~w18424;
assign w18426 = ~w18423 & ~w18425;
assign w18427 = ~w17607 & ~w18426;
assign w18428 = ~w15681 & w18427;
assign w18429 = w15681 & ~w18427;
assign w18430 = ~w18428 & ~w18429;
assign w18431 = (~w18430 & w18158) | (~w18430 & w41524) | (w18158 & w41524);
assign w18432 = ~w17588 & ~w17592;
assign w18433 = w14766 & ~w18432;
assign w18434 = w18431 & w18433;
assign w18435 = w14766 & w18432;
assign w18436 = ~w18431 & w18435;
assign w18437 = ~w18434 & ~w18436;
assign w18438 = ~w17598 & ~w17607;
assign w18439 = w17380 & ~w18438;
assign w18440 = ~w17380 & w18438;
assign w18441 = ~w18439 & ~w18440;
assign w18442 = (a[43] & w18158) | (a[43] & w45033) | (w18158 & w45033);
assign w18443 = ~w18183 & w18441;
assign w18444 = w18442 & ~w18443;
assign w18445 = ~w17584 & w17912;
assign w18446 = w17733 & w17912;
assign w18447 = ~w17724 & w18446;
assign w18448 = ~w18445 & ~w18447;
assign w18449 = w18054 & w18155;
assign w18450 = w18448 & w18449;
assign w18451 = (~w18164 & w18178) | (~w18164 & w47597) | (w18178 & w47597);
assign w18452 = ~w17816 & w18050;
assign w18453 = ~w17775 & w17876;
assign w18454 = ~w18452 & ~w18453;
assign w18455 = ~w17860 & w18155;
assign w18456 = ~w18452 & w47598;
assign w18457 = w18455 & ~w18456;
assign w18458 = ~w18451 & ~w18457;
assign w18459 = ~w18450 & w18458;
assign w18460 = ~w17595 & ~w17597;
assign w18461 = ~w18182 & ~w18460;
assign w18462 = ~a[43] & w18441;
assign w18463 = w18049 & w18462;
assign w18464 = (w18463 & ~w18459) | (w18463 & w45034) | (~w18459 & w45034);
assign w18465 = w18183 & w18424;
assign w18466 = ~w18464 & ~w18465;
assign w18467 = ~w18444 & w18466;
assign w18468 = ~w15681 & w18437;
assign w18469 = ~w18420 & w18468;
assign w18470 = ~w17617 & ~w17619;
assign w18471 = w17637 & w50204;
assign w18472 = (w18158 & w45035) | (w18158 & w45036) | (w45035 & w45036);
assign w18473 = ~w18471 & ~w18472;
assign w18474 = w14039 & ~w18473;
assign w18475 = w18431 & ~w18432;
assign w18476 = ~w18431 & w18432;
assign w18477 = ~w18475 & ~w18476;
assign w18478 = ~w14766 & w18477;
assign w18479 = ~w18474 & ~w18478;
assign w18480 = ~w18469 & w18479;
assign w18481 = w18437 & ~w18467;
assign w18482 = ~w18421 & w18481;
assign w18483 = w18480 & ~w18482;
assign w18484 = w17671 & ~w18197;
assign w18485 = w12666 & ~w18484;
assign w18486 = ~w12666 & w18484;
assign w18487 = ~w18485 & ~w18486;
assign w18488 = (~w18487 & w18158) | (~w18487 & w41527) | (w18158 & w41527);
assign w18489 = ~w17274 & ~w17658;
assign w18490 = w17274 & w17658;
assign w18491 = ~w18489 & ~w18490;
assign w18492 = ~w11870 & ~w18491;
assign w18493 = ~w18488 & w18492;
assign w18494 = ~w11870 & w18491;
assign w18495 = w18488 & w18494;
assign w18496 = ~w18493 & ~w18495;
assign w18497 = ~w13384 & w18196;
assign w18498 = w13384 & ~w18196;
assign w18499 = ~w18497 & ~w18498;
assign w18500 = (w18499 & w18158) | (w18499 & w41528) | (w18158 & w41528);
assign w18501 = ~w12666 & w17703;
assign w18502 = ~w18500 & w18501;
assign w18503 = ~w12666 & ~w17703;
assign w18504 = w18500 & w18503;
assign w18505 = ~w18502 & ~w18504;
assign w18506 = w18496 & w18505;
assign w18507 = w17639 & ~w18194;
assign w18508 = ~w18195 & ~w18507;
assign w18509 = ~w18158 & w41529;
assign w18510 = (w18508 & w18158) | (w18508 & w41530) | (w18158 & w41530);
assign w18511 = ~w18509 & ~w18510;
assign w18512 = w13384 & ~w18511;
assign w18513 = ~w14039 & w18473;
assign w18514 = ~w18512 & ~w18513;
assign w18515 = w18506 & w18514;
assign w18516 = (w18515 & ~w18480) | (w18515 & w41531) | (~w18480 & w41531);
assign w18517 = ~w13384 & w18511;
assign w18518 = w12666 & ~w17703;
assign w18519 = ~w18500 & w18518;
assign w18520 = w12666 & w17703;
assign w18521 = w18500 & w18520;
assign w18522 = ~w18519 & ~w18521;
assign w18523 = ~w18517 & w18522;
assign w18524 = w18506 & ~w18523;
assign w18525 = ~w18218 & w41532;
assign w18526 = w11870 & w18491;
assign w18527 = ~w18488 & w18526;
assign w18528 = w11870 & ~w18491;
assign w18529 = w18488 & w18528;
assign w18530 = ~w18527 & ~w18529;
assign w18531 = ~w18525 & w18530;
assign w18532 = w18212 & w18531;
assign w18533 = ~w18524 & w18532;
assign w18534 = ~w18288 & w18397;
assign w18535 = w18397 & w18533;
assign w18536 = ~w18516 & w18535;
assign w18537 = ~w18534 & ~w18536;
assign w18538 = ~w2285 & ~w17813;
assign w18539 = (w18538 & ~w18448) | (w18538 & w41533) | (~w18448 & w41533);
assign w18540 = ~w17813 & ~w18053;
assign w18541 = w2558 & ~w18540;
assign w18542 = ~w17813 & w17912;
assign w18543 = w18541 & ~w18542;
assign w18544 = w17584 & w18541;
assign w18545 = ~w17734 & w18544;
assign w18546 = ~w18545 & w41534;
assign w18547 = ~w18539 & w18546;
assign w18548 = ~w18183 & w18547;
assign w18549 = w17794 & w17812;
assign w18550 = ~w18182 & w18549;
assign w18551 = ~w18158 & w18550;
assign w18552 = ~w2558 & ~w17813;
assign w18553 = w17814 & w18552;
assign w18554 = (w18553 & ~w18448) | (w18553 & w41535) | (~w18448 & w41535);
assign w18555 = ~w3095 & ~w18554;
assign w18556 = ~w17813 & ~w18052;
assign w18557 = w18448 & w41536;
assign w18558 = (w18556 & ~w18448) | (w18556 & w41537) | (~w18448 & w41537);
assign w18559 = ~w18557 & ~w18558;
assign w18560 = ~w18158 & w41538;
assign w18561 = ~w18183 & w18559;
assign w18562 = ~w18560 & ~w18561;
assign w18563 = ~w18551 & w18555;
assign w18564 = ~w18548 & w18563;
assign w18565 = ~w18562 & ~w18564;
assign w18566 = w2285 & w17814;
assign w18567 = ~w2558 & w18540;
assign w18568 = ~w18545 & w41539;
assign w18569 = ~w18448 & w18552;
assign w18570 = w18568 & ~w18569;
assign w18571 = w2285 & ~w17814;
assign w18572 = (w18566 & w18183) | (w18566 & w41540) | (w18183 & w41540);
assign w18573 = ~w18183 & w41541;
assign w18574 = ~w18572 & ~w18573;
assign w18575 = w2285 & w17816;
assign w18576 = (w18575 & ~w18448) | (w18575 & w41542) | (~w18448 & w41542);
assign w18577 = ~w2285 & ~w17794;
assign w18578 = w18053 & w18577;
assign w18579 = ~w17816 & w18577;
assign w18580 = ~w2558 & w18566;
assign w18581 = ~w18579 & ~w18580;
assign w18582 = (w18581 & ~w18448) | (w18581 & w41543) | (~w18448 & w41543);
assign w18583 = ~w18576 & w18582;
assign w18584 = w2006 & ~w17773;
assign w18585 = (w18584 & w18183) | (w18584 & w41544) | (w18183 & w41544);
assign w18586 = w2006 & w17773;
assign w18587 = ~w18183 & w41545;
assign w18588 = ~w18585 & ~w18587;
assign w18589 = w18574 & w18588;
assign w18590 = ~w18565 & w18589;
assign w18591 = w2558 & w18562;
assign w18592 = (w17814 & w18183) | (w17814 & w41546) | (w18183 & w41546);
assign w18593 = ~w18183 & w41547;
assign w18594 = ~w18592 & ~w18593;
assign w18595 = ~w2285 & w18594;
assign w18596 = ~w18591 & ~w18595;
assign w18597 = w18590 & ~w18596;
assign w18598 = w17841 & w17885;
assign w18599 = w1320 & ~w1541;
assign w18600 = w18598 & w18599;
assign w18601 = w1320 & w1541;
assign w18602 = ~w18598 & w18601;
assign w18603 = ~w18600 & ~w18602;
assign w18604 = w18183 & w18603;
assign w18605 = ~w18452 & w47599;
assign w18606 = w17912 & w18605;
assign w18607 = ~w17735 & w18606;
assign w18608 = ~w18051 & w47600;
assign w18609 = w17775 & ~w17799;
assign w18610 = w18608 & ~w18609;
assign w18611 = ~w17875 & w18610;
assign w18612 = w18605 & ~w18611;
assign w18613 = (~w18612 & w17735) | (~w18612 & w41548) | (w17735 & w41548);
assign w18614 = w1320 & ~w18598;
assign w18615 = ~w18613 & w18614;
assign w18616 = w1320 & w18598;
assign w18617 = w18613 & w18616;
assign w18618 = ~w18615 & ~w18617;
assign w18619 = ~w18183 & w18618;
assign w18620 = ~w18604 & ~w18619;
assign w18621 = w17818 & w18610;
assign w18622 = w18448 & w18621;
assign w18623 = ~w17875 & ~w17880;
assign w18624 = ~w17818 & ~w17861;
assign w18625 = w18623 & ~w18624;
assign w18626 = ~w18623 & w18624;
assign w18627 = ~w18625 & ~w18626;
assign w18628 = w18448 & w41549;
assign w18629 = ~w18622 & ~w18627;
assign w18630 = ~w18628 & ~w18629;
assign w18631 = ~w18183 & w18630;
assign w18632 = w17879 & ~w18182;
assign w18633 = ~w18158 & w18632;
assign w18634 = (~w1541 & w18158) | (~w1541 & w45037) | (w18158 & w45037);
assign w18635 = ~w18631 & w18634;
assign w18636 = w1541 & w17841;
assign w18637 = w17885 & ~w18636;
assign w18638 = ~w1320 & ~w18598;
assign w18639 = ~w18612 & w18638;
assign w18640 = ~w18607 & w18639;
assign w18641 = ~w1320 & w18598;
assign w18642 = w18605 & w41550;
assign w18643 = ~w17735 & w18642;
assign w18644 = w18612 & w18641;
assign w18645 = ~w18643 & ~w18644;
assign w18646 = ~w18640 & w18645;
assign w18647 = ~w18183 & ~w18646;
assign w18648 = ~w1320 & ~w18637;
assign w18649 = ~w18158 & w41551;
assign w18650 = ~w18647 & ~w18649;
assign w18651 = ~w18635 & w18650;
assign w18652 = ~w18620 & ~w18651;
assign w18653 = w17886 & w18454;
assign w18654 = (w18653 & ~w18448) | (w18653 & w41552) | (~w18448 & w41552);
assign w18655 = ~w18158 & w45038;
assign w18656 = w17841 & ~w18654;
assign w18657 = ~w18183 & w18656;
assign w18658 = ~w18655 & ~w18657;
assign w18659 = ~w17827 & ~w17843;
assign w18660 = w1120 & ~w18659;
assign w18661 = (w18660 & w18657) | (w18660 & w45039) | (w18657 & w45039);
assign w18662 = w1120 & w18659;
assign w18663 = ~w18657 & w45040;
assign w18664 = ~w18661 & ~w18663;
assign w18665 = ~w18652 & w18664;
assign w18666 = (w17773 & w18183) | (w17773 & w41553) | (w18183 & w41553);
assign w18667 = ~w18183 & w41554;
assign w18668 = ~w18666 & ~w18667;
assign w18669 = ~w2006 & ~w18668;
assign w18670 = ~w17774 & ~w17799;
assign w18671 = ~w17774 & w17816;
assign w18672 = (w18671 & ~w18448) | (w18671 & w41555) | (~w18448 & w41555);
assign w18673 = ~w18670 & ~w18672;
assign w18674 = ~w18158 & w41556;
assign w18675 = ~w18183 & w18673;
assign w18676 = ~w17759 & ~w17861;
assign w18677 = ~w1738 & ~w18676;
assign w18678 = (w18677 & w18675) | (w18677 & w41557) | (w18675 & w41557);
assign w18679 = ~w1738 & w18676;
assign w18680 = ~w18675 & w41558;
assign w18681 = ~w18678 & ~w18680;
assign w18682 = ~w18669 & w18681;
assign w18683 = w18665 & w18682;
assign w18684 = ~w18597 & w18683;
assign w18685 = ~w17567 & ~w17906;
assign w18686 = ~w17515 & w41559;
assign w18687 = ~w17524 & ~w17578;
assign w18688 = ~w17907 & ~w18687;
assign w18689 = w17895 & ~w18688;
assign w18690 = ~w17907 & w18689;
assign w18691 = (w18690 & w17734) | (w18690 & w41560) | (w17734 & w41560);
assign w18692 = w18685 & ~w18688;
assign w18693 = ~w18685 & w18688;
assign w18694 = ~w18692 & ~w18693;
assign w18695 = w18685 & w18691;
assign w18696 = ~w18691 & w18694;
assign w18697 = ~w18695 & ~w18696;
assign w18698 = ~w18158 & w41561;
assign w18699 = ~w18183 & w18697;
assign w18700 = ~w18698 & ~w18699;
assign w18701 = ~w18699 & w41562;
assign w18702 = ~w17896 & w17909;
assign w18703 = (w18702 & w17734) | (w18702 & w41563) | (w17734 & w41563);
assign w18704 = ~w3242 & w18703;
assign w18705 = w3242 & ~w18703;
assign w18706 = ~w18704 & ~w18705;
assign w18707 = ~w18183 & w18706;
assign w18708 = ~w2896 & w17905;
assign w18709 = (w18708 & w18183) | (w18708 & w41564) | (w18183 & w41564);
assign w18710 = ~w2896 & ~w17905;
assign w18711 = ~w18183 & w41565;
assign w18712 = ~w18709 & ~w18711;
assign w18713 = ~w18701 & w18712;
assign w18714 = (~w3242 & w18699) | (~w3242 & w41566) | (w18699 & w41566);
assign w18715 = ~w17578 & ~w17907;
assign w18716 = w3646 & w18715;
assign w18717 = (w17895 & w17734) | (w17895 & w41567) | (w17734 & w41567);
assign w18718 = ~w17524 & ~w18717;
assign w18719 = w4056 & w18716;
assign w18720 = ~w18158 & w41568;
assign w18721 = w18716 & ~w18718;
assign w18722 = ~w18183 & w18721;
assign w18723 = ~w18720 & ~w18722;
assign w18724 = w3646 & ~w18715;
assign w18725 = w18718 & w18724;
assign w18726 = w3646 & w17907;
assign w18727 = ~w18158 & w41569;
assign w18728 = ~w18183 & w18725;
assign w18729 = ~w18727 & ~w18728;
assign w18730 = w18723 & w18729;
assign w18731 = ~w18714 & ~w18730;
assign w18732 = w18713 & ~w18731;
assign w18733 = w2896 & ~w17905;
assign w18734 = (w18733 & w18183) | (w18733 & w41570) | (w18183 & w41570);
assign w18735 = w2896 & w17905;
assign w18736 = ~w18183 & w41571;
assign w18737 = ~w18734 & ~w18736;
assign w18738 = ~w18565 & w18737;
assign w18739 = w18589 & w18738;
assign w18740 = ~w18732 & w18739;
assign w18741 = w18684 & ~w18740;
assign w18742 = ~w17854 & ~w18122;
assign w18743 = w17858 & ~w18124;
assign w18744 = w17842 & ~w18654;
assign w18745 = ~w17843 & ~w18744;
assign w18746 = w18183 & w18742;
assign w18747 = (~w18743 & w18158) | (~w18743 & w41572) | (w18158 & w41572);
assign w18748 = w18745 & w18747;
assign w18749 = (w18743 & w18158) | (w18743 & w41573) | (w18158 & w41573);
assign w18750 = ~w18745 & w18749;
assign w18751 = ~w18748 & ~w18750;
assign w18752 = ~w18746 & w18751;
assign w18753 = w945 & w18752;
assign w18754 = (w18125 & ~w18055) | (w18125 & w47601) | (~w18055 & w47601);
assign w18755 = ~w18078 & ~w18175;
assign w18756 = ~w18174 & ~w18755;
assign w18757 = (w18756 & w17915) | (w18756 & w41574) | (w17915 & w41574);
assign w18758 = w18174 & w18755;
assign w18759 = w18125 & w18755;
assign w18760 = (~w18758 & w18056) | (~w18758 & w41575) | (w18056 & w41575);
assign w18761 = w17914 & ~w18758;
assign w18762 = ~w17735 & w18761;
assign w18763 = ~w18760 & ~w18762;
assign w18764 = ~w18183 & w41576;
assign w18765 = ~w18077 & w18183;
assign w18766 = (w612 & ~w18183) | (w612 & w41577) | (~w18183 & w41577);
assign w18767 = ~w18764 & w18766;
assign w18768 = ~w945 & w18120;
assign w18769 = (w41578 & ~w18055) | (w41578 & w47602) | (~w18055 & w47602);
assign w18770 = (w18055 & w47603) | (w18055 & w47604) | (w47603 & w47604);
assign w18771 = w17914 & ~w18174;
assign w18772 = ~w17735 & w18771;
assign w18773 = ~w18770 & ~w18772;
assign w18774 = ~w17915 & w18769;
assign w18775 = w18773 & ~w18774;
assign w18776 = w945 & ~w18120;
assign w18777 = (w41580 & ~w18055) | (w41580 & w47605) | (~w18055 & w47605);
assign w18778 = (w18055 & w47606) | (w18055 & w47607) | (w47606 & w47607);
assign w18779 = w17914 & ~w18121;
assign w18780 = ~w17735 & w18779;
assign w18781 = ~w18778 & ~w18780;
assign w18782 = ~w17915 & w18777;
assign w18783 = w18781 & ~w18782;
assign w18784 = ~w18120 & ~w18182;
assign w18785 = ~w18158 & w18784;
assign w18786 = ~w18783 & ~w18785;
assign w18787 = ~w18183 & w18775;
assign w18788 = w18786 & ~w18787;
assign w18789 = ~w754 & w18788;
assign w18790 = ~w18764 & ~w18765;
assign w18791 = ~w612 & ~w18790;
assign w18792 = ~w18789 & ~w18791;
assign w18793 = ~w18767 & ~w18792;
assign w18794 = ~w18753 & ~w18793;
assign w18795 = ~w17498 & w18183;
assign w18796 = ~w18183 & w18378;
assign w18797 = ~w18795 & ~w18796;
assign w18798 = ~w6264 & ~w18797;
assign w18799 = w6769 & ~w18393;
assign w18800 = ~w18798 & ~w18799;
assign w18801 = w18386 & ~w18800;
assign w18802 = w5745 & ~w17486;
assign w18803 = ~w18158 & w41582;
assign w18804 = w5745 & ~w18355;
assign w18805 = ~w18183 & w18804;
assign w18806 = ~w18803 & ~w18805;
assign w18807 = ~w18365 & ~w18806;
assign w18808 = w4838 & w17891;
assign w18809 = ~w18158 & w41583;
assign w18810 = w4838 & ~w18315;
assign w18811 = ~w18183 & w18810;
assign w18812 = ~w18809 & ~w18811;
assign w18813 = ~w18351 & w18812;
assign w18814 = ~w18807 & w18813;
assign w18815 = w18332 & ~w18814;
assign w18816 = ~w4056 & w18307;
assign w18817 = ~w18158 & w41584;
assign w18818 = ~w4430 & ~w18817;
assign w18819 = ~w18183 & w18325;
assign w18820 = w18818 & ~w18819;
assign w18821 = ~w18308 & w18820;
assign w18822 = ~w18816 & ~w18821;
assign w18823 = ~w18815 & w18822;
assign w18824 = ~w18801 & w18823;
assign w18825 = w18794 & w18824;
assign w18826 = w18741 & w18825;
assign w18827 = w18537 & w18826;
assign w18828 = w754 & ~w18788;
assign w18829 = ~w18767 & ~w18828;
assign w18830 = ~w18791 & ~w18829;
assign w18831 = w18715 & w18718;
assign w18832 = ~w18715 & ~w18718;
assign w18833 = ~w18183 & w41585;
assign w18834 = (~w3646 & ~w18183) | (~w3646 & w41586) | (~w18183 & w41586);
assign w18835 = ~w18833 & w18834;
assign w18836 = ~w18714 & ~w18835;
assign w18837 = w18737 & w18836;
assign w18838 = ~w18713 & w18737;
assign w18839 = ~w18837 & ~w18838;
assign w18840 = w18590 & ~w18839;
assign w18841 = (~w18676 & w18675) | (~w18676 & w41587) | (w18675 & w41587);
assign w18842 = ~w18675 & w41588;
assign w18843 = ~w18841 & ~w18842;
assign w18844 = w1738 & w18843;
assign w18845 = ~w18631 & ~w18633;
assign w18846 = (w1541 & w18631) | (w1541 & w41589) | (w18631 & w41589);
assign w18847 = w18650 & w18846;
assign w18848 = ~w18620 & ~w18847;
assign w18849 = ~w18844 & w18848;
assign w18850 = w18665 & ~w18849;
assign w18851 = ~w945 & ~w18752;
assign w18852 = w18658 & ~w18659;
assign w18853 = ~w18658 & w18659;
assign w18854 = ~w18852 & ~w18853;
assign w18855 = ~w1120 & ~w18854;
assign w18856 = ~w18830 & ~w18851;
assign w18857 = ~w18855 & w18856;
assign w18858 = ~w18850 & w18857;
assign w18859 = w18684 & ~w18840;
assign w18860 = w18858 & ~w18859;
assign w18861 = ~w18794 & ~w18830;
assign w18862 = ~w18860 & ~w18861;
assign w18863 = ~w18457 & w41590;
assign w18864 = ~w18450 & w18863;
assign w18865 = ~w17974 & ~w18045;
assign w18866 = ~w17974 & w18040;
assign w18867 = ~w18865 & w50205;
assign w18868 = w16782 & ~w17961;
assign w18869 = ~w16782 & w17961;
assign w18870 = ~w18868 & ~w18869;
assign w18871 = w18867 & ~w18870;
assign w18872 = ~w18867 & w18870;
assign w18873 = ~w18871 & ~w18872;
assign w18874 = (~w18044 & w18158) | (~w18044 & w41592) | (w18158 & w41592);
assign w18875 = w18040 & ~w18864;
assign w18876 = w18874 & ~w18875;
assign w18877 = ~w3 & ~w18182;
assign w18878 = ~w18158 & w18877;
assign w18879 = ~w17974 & ~w18041;
assign w18880 = ~w18878 & w18879;
assign w18881 = ~w18158 & w41593;
assign w18882 = w18876 & w18880;
assign w18883 = ~w18880 & ~w18881;
assign w18884 = ~w18876 & w18883;
assign w18885 = ~w18882 & ~w18884;
assign w18886 = w42 & ~w18183;
assign w18887 = ~w18873 & w18886;
assign w18888 = w18885 & ~w18887;
assign w18889 = ~w16797 & w17944;
assign w18890 = ~w17944 & w17950;
assign w18891 = ~w18889 & ~w18890;
assign w18892 = ~w18867 & w18891;
assign w18893 = w18873 & ~w18892;
assign w18894 = ~w42 & ~w18893;
assign w18895 = w18885 & w41594;
assign w18896 = ~w18894 & ~w18895;
assign w18897 = w18885 & w18894;
assign w18898 = w18004 & w18166;
assign w18899 = w18004 & w18173;
assign w18900 = ~w18178 & w18899;
assign w18901 = ~w18898 & ~w18900;
assign w18902 = w18004 & ~w18024;
assign w18903 = ~w18457 & ~w18901;
assign w18904 = ~w18902 & ~w18903;
assign w18905 = w18024 & w18449;
assign w18906 = w18448 & w18905;
assign w18907 = ~w18904 & ~w18906;
assign w18908 = (w57 & w18904) | (w57 & w47608) | (w18904 & w47608);
assign w18909 = ~w18183 & ~w18908;
assign w18910 = ~w18904 & w47609;
assign w18911 = (~w17992 & ~w18907) | (~w17992 & w18005) | (~w18907 & w18005);
assign w18912 = w18909 & ~w18911;
assign w18913 = w80 & w18183;
assign w18914 = w18036 & ~w18044;
assign w18915 = ~w18912 & w41595;
assign w18916 = (w18914 & w18912) | (w18914 & w41596) | (w18912 & w41596);
assign w18917 = ~w18915 & ~w18916;
assign w18918 = w3 & ~w18917;
assign w18919 = ~w18897 & w18918;
assign w18920 = ~w18896 & ~w18919;
assign w18921 = w18004 & w18011;
assign w18922 = (~w18023 & w18457) | (~w18023 & w41597) | (w18457 & w41597);
assign w18923 = ~w18023 & w18449;
assign w18924 = w18448 & w18923;
assign w18925 = ~w18922 & ~w18924;
assign w18926 = (~w18921 & w18924) | (~w18921 & w41598) | (w18924 & w41598);
assign w18927 = w18921 & w18925;
assign w18928 = ~w252 & w18011;
assign w18929 = w18004 & ~w18928;
assign w18930 = w18183 & w18929;
assign w18931 = ~w18183 & ~w18926;
assign w18932 = ~w18927 & w18931;
assign w18933 = ~w18930 & ~w18932;
assign w18934 = ~w18932 & w41599;
assign w18935 = w18909 & ~w18910;
assign w18936 = ~w80 & ~w17992;
assign w18937 = (w18936 & ~w18909) | (w18936 & w41600) | (~w18909 & w41600);
assign w18938 = ~w80 & w17992;
assign w18939 = w18909 & w41601;
assign w18940 = ~w18937 & ~w18939;
assign w18941 = ~w18934 & w18940;
assign w18942 = w351 & ~w18022;
assign w18943 = (w18942 & w18450) | (w18942 & w41602) | (w18450 & w41602);
assign w18944 = ~w18183 & w18943;
assign w18945 = ~w351 & w18022;
assign w18946 = ~w18450 & w41603;
assign w18947 = (w18945 & w18450) | (w18945 & w41604) | (w18450 & w41604);
assign w18948 = ~w18946 & ~w18947;
assign w18949 = ~w18158 & w41605;
assign w18950 = ~w18450 & w41606;
assign w18951 = ~w18183 & w18950;
assign w18952 = ~w18949 & ~w18951;
assign w18953 = ~w18944 & w18948;
assign w18954 = w18952 & w18953;
assign w18955 = ~w252 & ~w18954;
assign w18956 = (~w57 & w18932) | (~w57 & w45041) | (w18932 & w45041);
assign w18957 = ~w18955 & ~w18956;
assign w18958 = w252 & w18954;
assign w18959 = w18098 & w18125;
assign w18960 = (~w18178 & w18056) | (~w18178 & w41607) | (w18056 & w41607);
assign w18961 = w17914 & ~w18178;
assign w18962 = ~w17735 & w18961;
assign w18963 = ~w18960 & ~w18962;
assign w18964 = w18136 & w18171;
assign w18965 = ~w18962 & w41608;
assign w18966 = ~w18183 & ~w18965;
assign w18967 = ~w18183 & w41609;
assign w18968 = ~w18158 & w41610;
assign w18969 = w18152 & w18163;
assign w18970 = ~w351 & ~w18969;
assign w18971 = ~w18968 & w18970;
assign w18972 = ~w18967 & w18971;
assign w18973 = ~w351 & w18969;
assign w18974 = w18171 & w18973;
assign w18975 = ~w18183 & w41611;
assign w18976 = w18968 & w18973;
assign w18977 = ~w18975 & ~w18976;
assign w18978 = ~w18972 & w18977;
assign w18979 = ~w18958 & w18978;
assign w18980 = w18941 & w18979;
assign w18981 = ~w18158 & w41612;
assign w18982 = (~w18175 & w18762) | (~w18175 & w41613) | (w18762 & w41613);
assign w18983 = ~w18183 & w18982;
assign w18984 = ~w18097 & ~w18100;
assign w18985 = w400 & ~w18984;
assign w18986 = ~w18983 & w41614;
assign w18987 = w400 & w18984;
assign w18988 = (w18987 & w18983) | (w18987 & w41615) | (w18983 & w41615);
assign w18989 = ~w18986 & ~w18988;
assign w18990 = ~w18963 & ~w18964;
assign w18991 = w18966 & ~w18990;
assign w18992 = w18130 & ~w18131;
assign w18993 = ~w18130 & w18131;
assign w18994 = ~w18992 & ~w18993;
assign w18995 = w18183 & ~w18994;
assign w18996 = ~w18991 & ~w18995;
assign w18997 = w400 & ~w493;
assign w18998 = ~w18991 & w41616;
assign w18999 = w18989 & w18998;
assign w19000 = ~w400 & w493;
assign w19001 = ~w18984 & w19000;
assign w19002 = (w19001 & w18983) | (w19001 & w41617) | (w18983 & w41617);
assign w19003 = w18984 & w19000;
assign w19004 = ~w18983 & w41618;
assign w19005 = ~w19002 & ~w19004;
assign w19006 = w351 & w18969;
assign w19007 = ~w18968 & w19006;
assign w19008 = ~w18967 & w19007;
assign w19009 = w351 & ~w18969;
assign w19010 = w18171 & w19009;
assign w19011 = ~w18183 & w41619;
assign w19012 = w18968 & w19009;
assign w19013 = ~w19011 & ~w19012;
assign w19014 = ~w19008 & w19013;
assign w19015 = w19005 & w19014;
assign w19016 = ~w18999 & w19015;
assign w19017 = w18941 & ~w18957;
assign w19018 = w18980 & ~w19016;
assign w19019 = ~w19017 & ~w19018;
assign w19020 = ~w3 & w18917;
assign w19021 = ~w17992 & ~w18935;
assign w19022 = w80 & ~w19021;
assign w19023 = w17992 & w18935;
assign w19024 = w19022 & ~w19023;
assign w19025 = ~w18897 & ~w19020;
assign w19026 = ~w19024 & w19025;
assign w19027 = w19019 & w19026;
assign w19028 = (w18920 & ~w19019) | (w18920 & w41620) | (~w19019 & w41620);
assign w19029 = ~w18862 & ~w19028;
assign w19030 = ~w18827 & w19029;
assign w19031 = ~w18983 & w41621;
assign w19032 = (w18984 & w18983) | (w18984 & w41622) | (w18983 & w41622);
assign w19033 = ~w19031 & ~w19032;
assign w19034 = ~w493 & ~w19033;
assign w19035 = w400 & ~w18996;
assign w19036 = ~w19034 & ~w19035;
assign w19037 = w18980 & w19036;
assign w19038 = w19019 & w41623;
assign w19039 = w18920 & ~w19038;
assign w19040 = ~w19030 & w19039;
assign w19041 = w18533 & ~w18516;
assign w19042 = w18288 & w50206;
assign w19043 = w18397 & w18840;
assign w19044 = ~w18850 & ~w18855;
assign w19045 = ~w18824 & w18840;
assign w19046 = w18741 & ~w19045;
assign w19047 = w19043 & w19044;
assign w19048 = ~w19042 & w19047;
assign w19049 = w19044 & ~w19046;
assign w19050 = ~w19048 & ~w19049;
assign w19051 = ~w18753 & ~w18851;
assign w19052 = ~w19050 & w19051;
assign w19053 = ~w18789 & ~w18828;
assign w19054 = ~w18753 & ~w19053;
assign w19055 = ~w18828 & ~w18851;
assign w19056 = (w19055 & ~w19050) | (w19055 & w45044) | (~w19050 & w45044);
assign w19057 = ~w19030 & w48946;
assign w19058 = (~w18789 & w19030) | (~w18789 & w41624) | (w19030 & w41624);
assign w19059 = w19056 & w19058;
assign w19060 = ~w19057 & ~w19059;
assign w19061 = ~w19040 & w48947;
assign w19062 = w19060 & ~w19061;
assign w19063 = w18562 & w19039;
assign w19064 = ~w19030 & w19063;
assign w19065 = w18397 & w18837;
assign w19066 = ~w19042 & w19065;
assign w19067 = w18824 & w41625;
assign w19068 = ~w18839 & ~w19067;
assign w19069 = ~w2558 & ~w18562;
assign w19070 = ~w18591 & ~w19069;
assign w19071 = w19065 & w19070;
assign w19072 = ~w19042 & w19071;
assign w19073 = ~w19068 & ~w19070;
assign w19074 = ~w19066 & w19073;
assign w19075 = w19068 & w19070;
assign w19076 = ~w19072 & ~w19075;
assign w19077 = ~w19074 & w19076;
assign w19078 = ~w19040 & w19077;
assign w19079 = ~w19064 & ~w19078;
assign w19080 = ~w2285 & ~w19079;
assign w19081 = (w2285 & w19030) | (w2285 & w41626) | (w19030 & w41626);
assign w19082 = ~w19078 & w19081;
assign w19083 = ~w18701 & ~w18836;
assign w19084 = w18397 & ~w19083;
assign w19085 = ~w19042 & w19084;
assign w19086 = w18712 & w18737;
assign w19087 = w18824 & w41627;
assign w19088 = ~w19083 & ~w19087;
assign w19089 = w19084 & w19086;
assign w19090 = ~w19042 & w19089;
assign w19091 = ~w19086 & ~w19088;
assign w19092 = ~w19085 & w19091;
assign w19093 = w19086 & w19088;
assign w19094 = ~w19090 & ~w19093;
assign w19095 = ~w19092 & w19094;
assign w19096 = ~w19040 & w19095;
assign w19097 = w17905 & ~w18707;
assign w19098 = ~w17905 & w18707;
assign w19099 = ~w19097 & ~w19098;
assign w19100 = w19039 & ~w19099;
assign w19101 = ~w19030 & w19100;
assign w19102 = (~w2558 & w19030) | (~w2558 & w41628) | (w19030 & w41628);
assign w19103 = ~w19096 & w19102;
assign w19104 = ~w19082 & ~w19103;
assign w19105 = w18730 & ~w18835;
assign w19106 = w18824 & w19105;
assign w19107 = (w19106 & w18536) | (w19106 & w41629) | (w18536 & w41629);
assign w19108 = (~w18835 & ~w18824) | (~w18835 & w41630) | (~w18824 & w41630);
assign w19109 = ~w18701 & ~w18714;
assign w19110 = w19108 & ~w19109;
assign w19111 = ~w19108 & w19109;
assign w19112 = ~w19110 & ~w19111;
assign w19113 = w19107 & w19112;
assign w19114 = ~w19107 & ~w19112;
assign w19115 = ~w19113 & ~w19114;
assign w19116 = ~w19030 & w41631;
assign w19117 = ~w19040 & w19115;
assign w19118 = ~w19116 & ~w19117;
assign w19119 = ~w19117 & w41632;
assign w19120 = ~w19096 & ~w19101;
assign w19121 = (w2558 & w19096) | (w2558 & w41633) | (w19096 & w41633);
assign w19122 = ~w19119 & ~w19121;
assign w19123 = w19104 & ~w19122;
assign w19124 = ~w19080 & ~w19123;
assign w19125 = w2285 & w19069;
assign w19126 = w18397 & w45045;
assign w19127 = ~w19042 & w19126;
assign w19128 = ~w18839 & ~w19069;
assign w19129 = ~w18591 & ~w19128;
assign w19130 = ~w18591 & ~w18838;
assign w19131 = w18824 & w41634;
assign w19132 = ~w2285 & ~w19069;
assign w19133 = w18397 & w45046;
assign w19134 = ~w19042 & w19133;
assign w19135 = (w2285 & w19131) | (w2285 & w45047) | (w19131 & w45047);
assign w19136 = ~w19127 & w19135;
assign w19137 = ~w19131 & w45048;
assign w19138 = ~w19134 & ~w19137;
assign w19139 = ~w19136 & w19138;
assign w19140 = w2339 & w18594;
assign w19141 = (w19140 & w19040) | (w19140 & w41635) | (w19040 & w41635);
assign w19142 = w2339 & ~w18594;
assign w19143 = ~w19040 & w41636;
assign w19144 = ~w19141 & ~w19143;
assign w19145 = w2006 & ~w18595;
assign w19146 = w18574 & ~w19069;
assign w19147 = w19145 & ~w19146;
assign w19148 = ~w18591 & w19145;
assign w19149 = ~w19068 & w19148;
assign w19150 = ~w19066 & w19149;
assign w19151 = ~w19147 & ~w19150;
assign w19152 = ~w19040 & w19151;
assign w19153 = w18840 & ~w19067;
assign w19154 = ~w18597 & ~w19153;
assign w19155 = w18590 & w19065;
assign w19156 = ~w19042 & w19155;
assign w19157 = w19154 & ~w19156;
assign w19158 = w18668 & w19157;
assign w19159 = w18669 & ~w19157;
assign w19160 = ~w19158 & ~w19159;
assign w19161 = (w18668 & w19040) | (w18668 & w41637) | (w19040 & w41637);
assign w19162 = w19152 & w19160;
assign w19163 = ~w19161 & ~w19162;
assign w19164 = w19144 & ~w19163;
assign w19165 = ~w2006 & w18594;
assign w19166 = (w19165 & w19040) | (w19165 & w41638) | (w19040 & w41638);
assign w19167 = ~w2006 & ~w18594;
assign w19168 = ~w19040 & w41639;
assign w19169 = ~w19166 & ~w19168;
assign w19170 = w1738 & w19169;
assign w19171 = ~w19164 & ~w19170;
assign w19172 = ~w4056 & w18183;
assign w19173 = ~w18183 & w18718;
assign w19174 = ~w19172 & ~w19173;
assign w19175 = w18715 & ~w19174;
assign w19176 = ~w18715 & w19174;
assign w19177 = ~w19175 & ~w19176;
assign w19178 = w18537 & w18824;
assign w19179 = w19105 & ~w19178;
assign w19180 = ~w19105 & w19178;
assign w19181 = ~w19179 & ~w19180;
assign w19182 = w19040 & w19177;
assign w19183 = ~w19040 & w19181;
assign w19184 = ~w19182 & ~w19183;
assign w19185 = ~w3242 & w19184;
assign w19186 = (w2896 & w19117) | (w2896 & w41640) | (w19117 & w41640);
assign w19187 = w19104 & ~w19186;
assign w19188 = ~w19185 & w19187;
assign w19189 = ~w19171 & ~w19188;
assign w19190 = w18681 & ~w18844;
assign w19191 = ~w18597 & ~w18740;
assign w19192 = ~w18669 & w19191;
assign w19193 = ~w19045 & w19192;
assign w19194 = ~w19042 & w19043;
assign w19195 = w19193 & ~w19194;
assign w19196 = w19190 & ~w19195;
assign w19197 = ~w19190 & w19195;
assign w19198 = ~w19196 & ~w19197;
assign w19199 = w18843 & w19040;
assign w19200 = ~w19040 & ~w19198;
assign w19201 = ~w19199 & ~w19200;
assign w19202 = w1541 & ~w19201;
assign w19203 = w2006 & ~w18594;
assign w19204 = (w19203 & w19040) | (w19203 & w41641) | (w19040 & w41641);
assign w19205 = w2006 & w18594;
assign w19206 = ~w19040 & w41642;
assign w19207 = ~w19204 & ~w19206;
assign w19208 = ~w1738 & w19207;
assign w19209 = ~w19162 & w41643;
assign w19210 = ~w19208 & ~w19209;
assign w19211 = (w18594 & w19040) | (w18594 & w41644) | (w19040 & w41644);
assign w19212 = ~w19040 & w41645;
assign w19213 = ~w19211 & ~w19212;
assign w19214 = w1738 & w19213;
assign w19215 = ~w19164 & ~w19214;
assign w19216 = w19210 & ~w19215;
assign w19217 = (~w19202 & w19215) | (~w19202 & w20063) | (w19215 & w20063);
assign w19218 = w19124 & w19189;
assign w19219 = w19124 & ~w19171;
assign w19220 = ~w19216 & ~w19219;
assign w19221 = ~w18308 & ~w18816;
assign w19222 = ~w18351 & w18806;
assign w19223 = w18395 & ~w18799;
assign w19224 = ~w18294 & w19223;
assign w19225 = (w18800 & w18294) | (w18800 & w41646) | (w18294 & w41646);
assign w19226 = w18383 & ~w19225;
assign w19227 = w18383 & ~w18800;
assign w19228 = w18288 & ~w19227;
assign w19229 = (w19222 & w19225) | (w19222 & w45049) | (w19225 & w45049);
assign w19230 = w18288 & w45050;
assign w19231 = ~w19041 & w19230;
assign w19232 = ~w19229 & ~w19231;
assign w19233 = ~w18361 & ~w18365;
assign w19234 = w18812 & ~w19233;
assign w19235 = w18331 & ~w19234;
assign w19236 = ~w18820 & ~w19235;
assign w19237 = w18812 & ~w18820;
assign w19238 = (w19237 & w19231) | (w19237 & w47610) | (w19231 & w47610);
assign w19239 = w18307 & w19039;
assign w19240 = ~w19030 & w19239;
assign w19241 = (w41647 & w19030) | (w41647 & w45051) | (w19030 & w45051);
assign w19242 = (w41648 & w19030) | (w41648 & w45052) | (w19030 & w45052);
assign w19243 = ~w19241 & ~w19242;
assign w19244 = ~w19240 & w19243;
assign w19245 = ~w3646 & w19244;
assign w19246 = w18330 & ~w18820;
assign w19247 = w18320 & ~w19234;
assign w19248 = (w18812 & w19231) | (w18812 & w47611) | (w19231 & w47611);
assign w19249 = w19247 & ~w19248;
assign w19250 = ~w19030 & w41649;
assign w19251 = (w19249 & w19030) | (w19249 & w45053) | (w19030 & w45053);
assign w19252 = ~w19250 & ~w19251;
assign w19253 = w4056 & w19246;
assign w19254 = (w19253 & w19251) | (w19253 & w41650) | (w19251 & w41650);
assign w19255 = w4056 & ~w19246;
assign w19256 = ~w19251 & w41651;
assign w19257 = ~w19254 & ~w19256;
assign w19258 = w3242 & ~w19184;
assign w19259 = w3646 & ~w19244;
assign w19260 = ~w19258 & ~w19259;
assign w19261 = ~w17891 & w18183;
assign w19262 = ~w18183 & w18315;
assign w19263 = ~w19261 & ~w19262;
assign w19264 = w18320 & w18812;
assign w19265 = w19232 & w19233;
assign w19266 = ~w19264 & w19265;
assign w19267 = w19264 & ~w19265;
assign w19268 = ~w19030 & w45054;
assign w19269 = ~w19040 & w41652;
assign w19270 = ~w19268 & ~w19269;
assign w19271 = ~w19269 & w45055;
assign w19272 = w19257 & w19271;
assign w19273 = ~w19245 & w19272;
assign w19274 = w19260 & ~w19273;
assign w19275 = ~w1541 & w19201;
assign w19276 = w18397 & w48948;
assign w19277 = ~w19042 & w19276;
assign w19278 = ~w18740 & w41653;
assign w19279 = ~w19045 & w19278;
assign w19280 = (~w18844 & w19045) | (~w18844 & w41654) | (w19045 & w41654);
assign w19281 = ~w19277 & ~w19280;
assign w19282 = ~w18635 & ~w18846;
assign w19283 = w19281 & ~w19282;
assign w19284 = ~w19281 & w19282;
assign w19285 = ~w19030 & w48949;
assign w19286 = ~w19040 & w41655;
assign w19287 = ~w19285 & ~w19286;
assign w19288 = ~w1320 & ~w19287;
assign w19289 = ~w19275 & ~w19288;
assign w19290 = (w19289 & w19218) | (w19289 & w41656) | (w19218 & w41656);
assign w19291 = w19274 & w19289;
assign w19292 = ~w19220 & w19291;
assign w19293 = ~w19290 & ~w19292;
assign w19294 = ~w18291 & w19039;
assign w19295 = ~w19030 & w19294;
assign w19296 = w18258 & ~w18292;
assign w19297 = w18225 & ~w18533;
assign w19298 = w19296 & ~w19297;
assign w19299 = w18225 & w18515;
assign w19300 = ~w18483 & w19299;
assign w19301 = w19298 & ~w19300;
assign w19302 = w18225 & w50206;
assign w19303 = ~w19296 & w19302;
assign w19304 = ~w19301 & ~w19303;
assign w19305 = ~w19030 & w41657;
assign w19306 = ~w8666 & w19304;
assign w19307 = (w19306 & w19030) | (w19306 & w45056) | (w19030 & w45056);
assign w19308 = ~w19305 & ~w19307;
assign w19309 = ~w18220 & w18515;
assign w19310 = ~w18483 & w19309;
assign w19311 = ~w18524 & w18531;
assign w19312 = ~w18220 & ~w19311;
assign w19313 = ~w18210 & ~w19312;
assign w19314 = (~w18221 & w19310) | (~w18221 & w41658) | (w19310 & w41658);
assign w19315 = ~w18211 & ~w18224;
assign w19316 = w19314 & ~w19315;
assign w19317 = ~w19314 & w19315;
assign w19318 = ~w19316 & ~w19317;
assign w19319 = w9195 & w18192;
assign w19320 = ~w19030 & w41659;
assign w19321 = w9195 & w19318;
assign w19322 = ~w19040 & w19321;
assign w19323 = ~w19320 & ~w19322;
assign w19324 = w19308 & w19323;
assign w19325 = w18235 & w18263;
assign w19326 = (w18258 & w19300) | (w18258 & w41660) | (w19300 & w41660);
assign w19327 = w19325 & ~w19326;
assign w19328 = ~w19325 & w19326;
assign w19329 = ~w19327 & ~w19328;
assign w19330 = (w19329 & w19030) | (w19329 & w41661) | (w19030 & w41661);
assign w19331 = ~w17415 & w18183;
assign w19332 = ~w18183 & w18230;
assign w19333 = ~w19331 & ~w19332;
assign w19334 = w19039 & ~w19333;
assign w19335 = ~w19030 & w19334;
assign w19336 = (w7924 & w19030) | (w7924 & w41662) | (w19030 & w41662);
assign w19337 = ~w19330 & w19336;
assign w19338 = ~w18291 & ~w19302;
assign w19339 = w8666 & ~w19338;
assign w19340 = (w19339 & w19030) | (w19339 & w41663) | (w19030 & w41663);
assign w19341 = w18291 & w19302;
assign w19342 = (w19341 & w19030) | (w19341 & w41664) | (w19030 & w41664);
assign w19343 = w19340 & ~w19342;
assign w19344 = ~w19337 & ~w19343;
assign w19345 = ~w19324 & w19344;
assign w19346 = w18247 & ~w18267;
assign w19347 = ~w18235 & w19346;
assign w19348 = w18264 & w19346;
assign w19349 = (w19348 & w19300) | (w19348 & w41665) | (w19300 & w41665);
assign w19350 = ~w19347 & ~w19349;
assign w19351 = w18247 & w19350;
assign w19352 = (w19351 & w19030) | (w19351 & w41666) | (w19030 & w41666);
assign w19353 = ~w7315 & w19039;
assign w19354 = ~w19030 & w19353;
assign w19355 = ~w18275 & w18286;
assign w19356 = w6769 & w19355;
assign w19357 = (w19356 & w19030) | (w19356 & w41667) | (w19030 & w41667);
assign w19358 = ~w19352 & w19357;
assign w19359 = w6769 & ~w19355;
assign w19360 = w19351 & w19359;
assign w19361 = ~w19040 & w19360;
assign w19362 = ~w19030 & w41668;
assign w19363 = ~w19361 & ~w19362;
assign w19364 = ~w19358 & w19363;
assign w19365 = ~w19030 & w41669;
assign w19366 = ~w7924 & w19329;
assign w19367 = ~w19040 & w19366;
assign w19368 = ~w19365 & ~w19367;
assign w19369 = (w18264 & w19300) | (w18264 & w41670) | (w19300 & w41670);
assign w19370 = w18235 & ~w19346;
assign w19371 = ~w19369 & w19370;
assign w19372 = w19350 & ~w19371;
assign w19373 = ~w7315 & ~w19372;
assign w19374 = ~w19040 & w19373;
assign w19375 = ~w8666 & w18183;
assign w19376 = ~w18183 & w18239;
assign w19377 = ~w19375 & ~w19376;
assign w19378 = w18237 & ~w19377;
assign w19379 = ~w18237 & w19377;
assign w19380 = ~w19378 & ~w19379;
assign w19381 = ~w19030 & w41671;
assign w19382 = ~w19374 & ~w19381;
assign w19383 = w19368 & w19382;
assign w19384 = w19364 & w19383;
assign w19385 = ~w19040 & w19304;
assign w19386 = w8666 & ~w19295;
assign w19387 = ~w19385 & w19386;
assign w19388 = ~w19337 & ~w19387;
assign w19389 = ~w19310 & ~w19312;
assign w19390 = ~w18210 & ~w18221;
assign w19391 = w19389 & ~w19390;
assign w19392 = ~w19389 & w19390;
assign w19393 = ~w19391 & ~w19392;
assign w19394 = ~w19040 & ~w19393;
assign w19395 = w18209 & w19039;
assign w19396 = ~w19030 & w19395;
assign w19397 = w9781 & ~w19396;
assign w19398 = ~w19394 & w19397;
assign w19399 = ~w9195 & ~w18192;
assign w19400 = w19040 & w19399;
assign w19401 = ~w9195 & ~w19318;
assign w19402 = ~w19040 & w19401;
assign w19403 = ~w19400 & ~w19402;
assign w19404 = ~w19398 & w19403;
assign w19405 = w19388 & w19404;
assign w19406 = ~w19352 & ~w19354;
assign w19407 = w19355 & ~w19406;
assign w19408 = ~w19355 & w19406;
assign w19409 = ~w19407 & ~w19408;
assign w19410 = ~w6769 & ~w19409;
assign w19411 = ~w19040 & w19372;
assign w19412 = w19040 & ~w19380;
assign w19413 = ~w19411 & ~w19412;
assign w19414 = w7315 & ~w19413;
assign w19415 = w19364 & w19414;
assign w19416 = ~w19410 & ~w19415;
assign w19417 = ~w19345 & w19384;
assign w19418 = ~w19405 & w19417;
assign w19419 = w19416 & ~w19418;
assign w19420 = ~w17380 & w18183;
assign w19421 = w17380 & ~w18183;
assign w19422 = ~w19420 & ~w19421;
assign w19423 = ~w18827 & ~w18862;
assign w19424 = ~w17380 & ~w19026;
assign w19425 = w19019 & ~w19037;
assign w19426 = (w18183 & w19425) | (w18183 & w45057) | (w19425 & w45057);
assign w19427 = (w18920 & ~w19425) | (w18920 & w45058) | (~w19425 & w45058);
assign w19428 = ~w19426 & w19427;
assign w19429 = ~w19018 & w41672;
assign w19430 = ~w19020 & w19429;
assign w19431 = ~w17380 & w18920;
assign w19432 = ~w18183 & w18897;
assign w19433 = (~w19432 & w19430) | (~w19432 & w45059) | (w19430 & w45059);
assign w19434 = ~w19422 & ~w19430;
assign w19435 = w19433 & ~w19434;
assign w19436 = ~w19428 & w19435;
assign w19437 = ~w19423 & ~w19436;
assign w19438 = w19428 & ~w19433;
assign w19439 = w18399 & w19422;
assign w19440 = ~w19438 & w19439;
assign w19441 = ~w19437 & w19440;
assign w19442 = ~a[40] & ~w18183;
assign w19443 = ~w19030 & w41673;
assign w19444 = ~w18399 & ~w19422;
assign w19445 = (~w19444 & w19030) | (~w19444 & w41674) | (w19030 & w41674);
assign w19446 = ~w19443 & ~w19445;
assign w19447 = ~a[41] & ~w19446;
assign w19448 = ~w19441 & w19447;
assign w19449 = w18897 & w19420;
assign w19450 = (w19449 & ~w19429) | (w19449 & w45060) | (~w19429 & w45060);
assign w19451 = (w19450 & w18827) | (w19450 & w41675) | (w18827 & w41675);
assign w19452 = ~w18406 & ~w19442;
assign w19453 = ~w19451 & w19452;
assign w19454 = w17380 & ~w18398;
assign w19455 = ~w17380 & w18398;
assign w19456 = ~w19454 & ~w19455;
assign w19457 = w19442 & w19456;
assign w19458 = a[41] & ~w19457;
assign w19459 = (w19458 & w19030) | (w19458 & w45061) | (w19030 & w45061);
assign w19460 = w19445 & w19453;
assign w19461 = w19459 & ~w19460;
assign w19462 = ~a[36] & ~a[37];
assign w19463 = ~a[38] & w19462;
assign w19464 = ~w18183 & w19463;
assign w19465 = w18183 & ~w19463;
assign w19466 = ~w19464 & ~w19465;
assign w19467 = a[39] & ~w19466;
assign w19468 = ~w18398 & ~w19467;
assign w19469 = ~w19464 & ~w19468;
assign w19470 = a[40] & ~w18398;
assign w19471 = ~w18399 & ~w19470;
assign w19472 = w17380 & ~w19469;
assign w19473 = ~w19471 & ~w19472;
assign w19474 = ~w17380 & w19469;
assign w19475 = ~w19473 & ~w19474;
assign w19476 = a[40] & w18183;
assign w19477 = ~w19442 & ~w19476;
assign w19478 = ~a[39] & w19466;
assign w19479 = ~w19464 & ~w19478;
assign w19480 = w17380 & ~w19479;
assign w19481 = ~w19477 & ~w19480;
assign w19482 = ~w17380 & w19479;
assign w19483 = (w19475 & w19030) | (w19475 & w41676) | (w19030 & w41676);
assign w19484 = ~w19481 & ~w19482;
assign w19485 = ~w19030 & w41677;
assign w19486 = ~w19483 & ~w19485;
assign w19487 = w16559 & w19486;
assign w19488 = ~w19461 & ~w19487;
assign w19489 = ~w19448 & w19488;
assign w19490 = w18437 & ~w18478;
assign w19491 = ~w15681 & ~w18420;
assign w19492 = ~w18421 & ~w18467;
assign w19493 = ~w19491 & ~w19492;
assign w19494 = w19490 & ~w19493;
assign w19495 = ~w19490 & w19493;
assign w19496 = ~w19494 & ~w19495;
assign w19497 = ~w19030 & w41678;
assign w19498 = (w19496 & w19030) | (w19496 & w41679) | (w19030 & w41679);
assign w19499 = ~w19497 & ~w19498;
assign w19500 = w14039 & ~w19499;
assign w19501 = ~w18421 & ~w19491;
assign w19502 = (w19501 & w19030) | (w19501 & w41680) | (w19030 & w41680);
assign w19503 = ~w14766 & ~w18467;
assign w19504 = (~w19030 & w45062) | (~w19030 & w45063) | (w45062 & w45063);
assign w19505 = ~w14766 & w18467;
assign w19506 = (w19030 & w45064) | (w19030 & w45065) | (w45064 & w45065);
assign w19507 = ~w19504 & ~w19506;
assign w19508 = ~w19500 & w19507;
assign w19509 = ~w16559 & ~w19486;
assign w19510 = ~w18408 & ~w18411;
assign w19511 = ~w15681 & ~w18418;
assign w19512 = (~w19030 & w45066) | (~w19030 & w45067) | (w45066 & w45067);
assign w19513 = ~w15681 & w18418;
assign w19514 = (w19030 & w45068) | (w19030 & w45069) | (w45068 & w45069);
assign w19515 = ~w19512 & ~w19514;
assign w19516 = ~w19509 & w19515;
assign w19517 = w19508 & w19516;
assign w19518 = ~w19489 & w19517;
assign w19519 = ~w14039 & w19499;
assign w19520 = w15681 & w18418;
assign w19521 = (~w19030 & w45070) | (~w19030 & w45071) | (w45070 & w45071);
assign w19522 = w15681 & ~w18418;
assign w19523 = (w19030 & w45072) | (w19030 & w45073) | (w45072 & w45073);
assign w19524 = ~w19521 & ~w19523;
assign w19525 = w14766 & w18467;
assign w19526 = (~w19030 & w45074) | (~w19030 & w45075) | (w45074 & w45075);
assign w19527 = w14766 & ~w18467;
assign w19528 = (w19030 & w45076) | (w19030 & w45077) | (w45076 & w45077);
assign w19529 = ~w19526 & ~w19528;
assign w19530 = w19524 & w19529;
assign w19531 = (~w19519 & ~w19508) | (~w19519 & w45078) | (~w19508 & w45078);
assign w19532 = ~w19518 & w19531;
assign w19533 = (w18514 & ~w18480) | (w18514 & w41682) | (~w18480 & w41682);
assign w19534 = ~w18517 & ~w19533;
assign w19535 = w18505 & ~w19534;
assign w19536 = w18496 & w18530;
assign w19537 = w18530 & w18920;
assign w19538 = (~w19536 & w19027) | (~w19536 & w41683) | (w19027 & w41683);
assign w19539 = w18522 & ~w19535;
assign w19540 = w19538 & ~w19539;
assign w19541 = w18522 & w18530;
assign w19542 = ~w19535 & w19541;
assign w19543 = ~w19540 & ~w19542;
assign w19544 = w18488 & ~w18491;
assign w19545 = ~w18488 & w18491;
assign w19546 = ~w19544 & ~w19545;
assign w19547 = w19039 & w19546;
assign w19548 = ~w19030 & w19547;
assign w19549 = ~w18496 & ~w19540;
assign w19550 = ~w19548 & ~w19549;
assign w19551 = ~w19040 & w19543;
assign w19552 = w19550 & ~w19551;
assign w19553 = ~w11138 & w19552;
assign w19554 = w18219 & w19039;
assign w19555 = ~w19030 & w19554;
assign w19556 = ~w18220 & ~w18525;
assign w19557 = w18506 & ~w19534;
assign w19558 = w18496 & ~w19541;
assign w19559 = ~w19557 & ~w19558;
assign w19560 = w19556 & ~w19559;
assign w19561 = ~w19556 & w19559;
assign w19562 = ~w19560 & ~w19561;
assign w19563 = ~w19040 & w19562;
assign w19564 = (w10419 & w19563) | (w10419 & w41684) | (w19563 & w41684);
assign w19565 = ~w19553 & ~w19564;
assign w19566 = ~w17703 & ~w18500;
assign w19567 = w17703 & w18500;
assign w19568 = ~w19566 & ~w19567;
assign w19569 = w19039 & ~w19568;
assign w19570 = w18505 & w18522;
assign w19571 = w19534 & ~w19570;
assign w19572 = ~w19534 & w19570;
assign w19573 = ~w19571 & ~w19572;
assign w19574 = ~w19030 & w41685;
assign w19575 = w11870 & w19573;
assign w19576 = (w19575 & w19030) | (w19575 & w41686) | (w19030 & w41686);
assign w19577 = ~w19574 & ~w19576;
assign w19578 = ~w18512 & ~w18517;
assign w19579 = ~w18483 & ~w18513;
assign w19580 = w19578 & ~w19579;
assign w19581 = ~w19578 & w19579;
assign w19582 = ~w19580 & ~w19581;
assign w19583 = w12666 & w18511;
assign w19584 = ~w19030 & w41687;
assign w19585 = w12666 & ~w19582;
assign w19586 = (w19585 & w19030) | (w19585 & w41688) | (w19030 & w41688);
assign w19587 = ~w19584 & ~w19586;
assign w19588 = w19577 & w19587;
assign w19589 = ~w18478 & ~w19494;
assign w19590 = ~w18474 & ~w18513;
assign w19591 = w19589 & ~w19590;
assign w19592 = ~w19589 & w19590;
assign w19593 = ~w19591 & ~w19592;
assign w19594 = ~w19030 & w45079;
assign w19595 = (w19593 & w19030) | (w19593 & w45080) | (w19030 & w45080);
assign w19596 = ~w19594 & ~w19595;
assign w19597 = ~w13384 & ~w19596;
assign w19598 = w13384 & w18473;
assign w19599 = ~w19030 & w41689;
assign w19600 = w13384 & ~w19593;
assign w19601 = (w19600 & w19030) | (w19600 & w41690) | (w19030 & w41690);
assign w19602 = ~w19599 & ~w19601;
assign w19603 = ~w12666 & ~w18511;
assign w19604 = ~w19030 & w41691;
assign w19605 = ~w12666 & w19582;
assign w19606 = (w19605 & w19030) | (w19605 & w41692) | (w19030 & w41692);
assign w19607 = ~w19604 & ~w19606;
assign w19608 = w19602 & w19607;
assign w19609 = w19588 & ~w19608;
assign w19610 = (~w11870 & w19030) | (~w11870 & w41693) | (w19030 & w41693);
assign w19611 = (w19573 & w19030) | (w19573 & w45081) | (w19030 & w45081);
assign w19612 = w19610 & ~w19611;
assign w19613 = w11138 & ~w19552;
assign w19614 = (~w19612 & w19552) | (~w19612 & w45082) | (w19552 & w45082);
assign w19615 = ~w19609 & w19614;
assign w19616 = w19588 & ~w19597;
assign w19617 = (w19565 & ~w19615) | (w19565 & w41694) | (~w19615 & w41694);
assign w19618 = ~w19532 & w19617;
assign w19619 = (~w10419 & w19030) | (~w10419 & w41695) | (w19030 & w41695);
assign w19620 = ~w19563 & w19619;
assign w19621 = ~w19612 & ~w19620;
assign w19622 = ~w19613 & w19621;
assign w19623 = ~w19609 & w19622;
assign w19624 = (~w19620 & w19553) | (~w19620 & w41696) | (w19553 & w41696);
assign w19625 = ~w19623 & ~w19624;
assign w19626 = ~w19394 & ~w19396;
assign w19627 = ~w9781 & ~w19626;
assign w19628 = w19417 & ~w19627;
assign w19629 = ~w19625 & w19628;
assign w19630 = ~w19618 & w19629;
assign w19631 = w19419 & ~w19630;
assign w19632 = w18383 & ~w18798;
assign w19633 = ~w18294 & w41697;
assign w19634 = ~w18516 & w19633;
assign w19635 = ~w18288 & w19224;
assign w19636 = (~w18799 & ~w19224) | (~w18799 & w41698) | (~w19224 & w41698);
assign w19637 = ~w19634 & w19636;
assign w19638 = w19632 & ~w19637;
assign w19639 = ~w19632 & w19637;
assign w19640 = ~w19638 & ~w19639;
assign w19641 = w5745 & ~w18797;
assign w19642 = ~w19030 & w41699;
assign w19643 = w5745 & w19640;
assign w19644 = ~w19040 & w19643;
assign w19645 = ~w19642 & ~w19644;
assign w19646 = ~w18394 & ~w18799;
assign w19647 = w18286 & ~w18294;
assign w19648 = ~w19646 & ~w19647;
assign w19649 = ~w19635 & ~w19648;
assign w19650 = ~w19634 & w19649;
assign w19651 = w19042 & ~w19646;
assign w19652 = w19650 & ~w19651;
assign w19653 = ~w6264 & ~w18393;
assign w19654 = ~w19030 & w41700;
assign w19655 = ~w6264 & w19652;
assign w19656 = ~w19040 & w19655;
assign w19657 = ~w19654 & ~w19656;
assign w19658 = w19645 & w19657;
assign w19659 = w4430 & ~w19270;
assign w19660 = ~w5745 & w19039;
assign w19661 = ~w19030 & w19660;
assign w19662 = ~w19041 & w19228;
assign w19663 = w19226 & ~w19662;
assign w19664 = (~w19663 & w19030) | (~w19663 & w41701) | (w19030 & w41701);
assign w19665 = ~w19661 & ~w19664;
assign w19666 = w18360 & w18806;
assign w19667 = ~w5330 & ~w19666;
assign w19668 = w19665 & w19667;
assign w19669 = ~w5330 & w19666;
assign w19670 = ~w19665 & w19669;
assign w19671 = ~w19668 & ~w19670;
assign w19672 = ~w4838 & w19671;
assign w19673 = ~w19246 & w19252;
assign w19674 = ~w4056 & ~w19673;
assign w19675 = w19246 & ~w19252;
assign w19676 = w19674 & ~w19675;
assign w19677 = ~w19659 & ~w19672;
assign w19678 = ~w19676 & ~w19677;
assign w19679 = ~w19218 & w41702;
assign w19680 = w19658 & ~w19679;
assign w19681 = ~w19245 & w19257;
assign w19682 = w19260 & ~w19681;
assign w19683 = w19188 & ~w19682;
assign w19684 = w19219 & ~w19683;
assign w19685 = w19217 & ~w19684;
assign w19686 = ~w5745 & ~w19640;
assign w19687 = ~w19040 & w19686;
assign w19688 = ~w19030 & w41703;
assign w19689 = ~w19687 & ~w19688;
assign w19690 = w6264 & w18393;
assign w19691 = ~w19030 & w41704;
assign w19692 = w6264 & ~w19652;
assign w19693 = ~w19040 & w19692;
assign w19694 = ~w19691 & ~w19693;
assign w19695 = w19689 & w19694;
assign w19696 = w19645 & ~w19695;
assign w19697 = w5330 & ~w19666;
assign w19698 = ~w19665 & w19697;
assign w19699 = w5330 & w19666;
assign w19700 = w19665 & w19699;
assign w19701 = ~w19698 & ~w19700;
assign w19702 = ~w19696 & w19701;
assign w19703 = w19672 & ~w19702;
assign w19704 = ~w19659 & ~w19703;
assign w19705 = ~w19676 & ~w19704;
assign w19706 = w19685 & ~w19705;
assign w19707 = ~w19631 & w19680;
assign w19708 = w19706 & ~w19707;
assign w19709 = (w19671 & w19696) | (w19671 & w41705) | (w19696 & w41705);
assign w19710 = w4838 & ~w19709;
assign w19711 = w19419 & w19710;
assign w19712 = w4838 & ~w19658;
assign w19713 = w19702 & w19712;
assign w19714 = ~w18351 & ~w18365;
assign w19715 = w18360 & w19663;
assign w19716 = w18806 & ~w19715;
assign w19717 = w5330 & w19040;
assign w19718 = ~w19040 & w19716;
assign w19719 = ~w19717 & ~w19718;
assign w19720 = w19714 & ~w19719;
assign w19721 = ~w19714 & w19719;
assign w19722 = ~w19720 & ~w19721;
assign w19723 = ~w19665 & ~w19666;
assign w19724 = w6027 & ~w19723;
assign w19725 = w19665 & w19666;
assign w19726 = w19724 & ~w19725;
assign w19727 = w19722 & ~w19726;
assign w19728 = ~w19713 & w19727;
assign w19729 = ~w19711 & w19728;
assign w19730 = w19629 & w19728;
assign w19731 = ~w19618 & w19730;
assign w19732 = ~w19729 & ~w19731;
assign w19733 = w19274 & ~w19676;
assign w19734 = ~w19220 & w19733;
assign w19735 = ~w19732 & w19734;
assign w19736 = w19708 & ~w19735;
assign w19737 = ~w19293 & ~w19736;
assign w19738 = w18849 & ~w19279;
assign w19739 = w18849 & w19043;
assign w19740 = ~w19042 & w19739;
assign w19741 = ~w19738 & ~w19740;
assign w19742 = ~w18652 & w19741;
assign w19743 = w18664 & ~w18855;
assign w19744 = ~w945 & ~w18652;
assign w19745 = ~w19743 & w19744;
assign w19746 = w19741 & w19745;
assign w19747 = ~w945 & ~w18854;
assign w19748 = ~w19030 & w41706;
assign w19749 = ~w19040 & w19746;
assign w19750 = ~w19748 & ~w19749;
assign w19751 = ~w945 & w19743;
assign w19752 = ~w19040 & w41707;
assign w19753 = w19750 & ~w19752;
assign w19754 = w19050 & ~w19051;
assign w19755 = ~w19030 & w41708;
assign w19756 = w754 & ~w19755;
assign w19757 = ~w19040 & w41709;
assign w19758 = w19756 & ~w19757;
assign w19759 = w19753 & ~w19758;
assign w19760 = ~w18635 & ~w19280;
assign w19761 = ~w19277 & w19760;
assign w19762 = ~w18846 & ~w19761;
assign w19763 = ~w19040 & w19762;
assign w19764 = ~w1320 & w19039;
assign w19765 = ~w19030 & w19764;
assign w19766 = ~w18620 & w18650;
assign w19767 = w1120 & w19766;
assign w19768 = (w19767 & w19030) | (w19767 & w41710) | (w19030 & w41710);
assign w19769 = ~w19763 & w19768;
assign w19770 = w1120 & ~w19766;
assign w19771 = ~w19030 & w41711;
assign w19772 = ~w18846 & w19770;
assign w19773 = ~w19761 & w19772;
assign w19774 = ~w19040 & w19773;
assign w19775 = ~w19771 & ~w19774;
assign w19776 = ~w19769 & w19775;
assign w19777 = w945 & ~w18652;
assign w19778 = w19743 & w19777;
assign w19779 = w19741 & w19778;
assign w19780 = w945 & w18854;
assign w19781 = ~w19030 & w41712;
assign w19782 = ~w19040 & w19779;
assign w19783 = ~w19781 & ~w19782;
assign w19784 = w945 & ~w19743;
assign w19785 = ~w19040 & w41713;
assign w19786 = w19783 & ~w19785;
assign w19787 = w19776 & w19786;
assign w19788 = w19759 & ~w19787;
assign w19789 = ~w19030 & w41714;
assign w19790 = (w19050 & w19030) | (w19050 & w41715) | (w19030 & w41715);
assign w19791 = ~w19789 & ~w19790;
assign w19792 = w19051 & w19791;
assign w19793 = ~w754 & ~w19792;
assign w19794 = ~w19051 & ~w19791;
assign w19795 = w19793 & ~w19794;
assign w19796 = ~w19788 & ~w19795;
assign w19797 = (~w612 & w19788) | (~w612 & w41716) | (w19788 & w41716);
assign w19798 = ~w19056 & w19058;
assign w19799 = ~w19030 & w45083;
assign w19800 = ~w18767 & ~w18791;
assign w19801 = ~w493 & ~w19800;
assign w19802 = ~w19798 & w45084;
assign w19803 = ~w493 & w19800;
assign w19804 = (w19803 & w19798) | (w19803 & w45085) | (w19798 & w45085);
assign w19805 = ~w19802 & ~w19804;
assign w19806 = ~w19062 & w19805;
assign w19807 = w19806 & ~w19797;
assign w19808 = w612 & w19805;
assign w19809 = ~w19798 & w45086;
assign w19810 = (w19800 & w19798) | (w19800 & w45087) | (w19798 & w45087);
assign w19811 = ~w19809 & ~w19810;
assign w19812 = w493 & w19811;
assign w19813 = (~w19812 & ~w19796) | (~w19812 & w41717) | (~w19796 & w41717);
assign w19814 = ~w19807 & w19813;
assign w19815 = (~w18934 & w19030) | (~w18934 & w41718) | (w19030 & w41718);
assign w19816 = w80 & w19039;
assign w19817 = ~w19030 & w19816;
assign w19818 = w19016 & ~w19036;
assign w19819 = w18979 & ~w19818;
assign w19820 = ~w19815 & ~w19817;
assign w19821 = ~w19817 & w41721;
assign w19822 = ~w19820 & ~w19821;
assign w19823 = w18940 & ~w19024;
assign w19824 = w19822 & ~w19823;
assign w19825 = ~w19822 & w19823;
assign w19826 = ~w19824 & ~w19825;
assign w19827 = ~w3 & ~w19826;
assign w19828 = ~w18918 & ~w19020;
assign w19829 = (~w19024 & ~w18980) | (~w19024 & w41722) | (~w18980 & w41722);
assign w19830 = w19019 & w19829;
assign w19831 = w18826 & ~w19830;
assign w19832 = w18537 & w19831;
assign w19833 = ~w18860 & w41723;
assign w19834 = w19429 & ~w19833;
assign w19835 = ~w19832 & w19834;
assign w19836 = ~w19828 & ~w19835;
assign w19837 = w19828 & ~w19832;
assign w19838 = w19834 & w19837;
assign w19839 = ~w18917 & w19040;
assign w19840 = ~w19040 & ~w19838;
assign w19841 = ~w19836 & w19840;
assign w19842 = ~w19839 & ~w19841;
assign w19843 = ~w19841 & w41724;
assign w19844 = ~w19040 & w41725;
assign w19845 = ~w19030 & w45088;
assign w19846 = ~w18934 & ~w18956;
assign w19847 = (w19846 & w19030) | (w19846 & w41726) | (w19030 & w41726);
assign w19848 = ~w19845 & ~w19847;
assign w19849 = w19844 & w19848;
assign w19850 = ~w19844 & ~w19848;
assign w19851 = ~w19849 & ~w19850;
assign w19852 = w80 & w19851;
assign w19853 = (~w19843 & ~w19851) | (~w19843 & w41727) | (~w19851 & w41727);
assign w19854 = ~w19827 & w19853;
assign w19855 = ~w80 & ~w19851;
assign w19856 = (~w19818 & w18827) | (~w19818 & w41728) | (w18827 & w41728);
assign w19857 = ~w19040 & w41729;
assign w19858 = ~w19030 & w41730;
assign w19859 = ~w18955 & ~w18958;
assign w19860 = w57 & ~w19859;
assign w19861 = ~w19857 & w48950;
assign w19862 = w57 & w19859;
assign w19863 = (w19862 & w19857) | (w19862 & w48951) | (w19857 & w48951);
assign w19864 = ~w19861 & ~w19863;
assign w19865 = ~w19855 & w19864;
assign w19866 = ~w57 & w19859;
assign w19867 = (w19866 & w19030) | (w19866 & w48952) | (w19030 & w48952);
assign w19868 = ~w19857 & w19867;
assign w19869 = ~w57 & ~w19859;
assign w19870 = w18978 & w19869;
assign w19871 = ~w19040 & w41731;
assign w19872 = ~w19030 & w48953;
assign w19873 = ~w19871 & ~w19872;
assign w19874 = ~w19868 & w19873;
assign w19875 = w18978 & w19014;
assign w19876 = ~w18999 & w19005;
assign w19877 = ~w19875 & ~w19876;
assign w19878 = w18978 & w19818;
assign w19879 = ~w19877 & ~w19878;
assign w19880 = (w19879 & w19030) | (w19879 & w41732) | (w19030 & w41732);
assign w19881 = w18978 & w19016;
assign w19882 = (w19881 & w18860) | (w19881 & w41733) | (w18860 & w41733);
assign w19883 = ~w18827 & w19882;
assign w19884 = w19036 & ~w19875;
assign w19885 = w18826 & w19884;
assign w19886 = w18537 & w19885;
assign w19887 = ~w18860 & w41734;
assign w19888 = ~w19886 & ~w19887;
assign w19889 = ~w19883 & w19888;
assign w19890 = ~w18967 & ~w18968;
assign w19891 = w18969 & ~w19890;
assign w19892 = ~w18969 & w19890;
assign w19893 = ~w19891 & ~w19892;
assign w19894 = ~w19030 & w41735;
assign w19895 = w19880 & w19889;
assign w19896 = ~w19894 & ~w19895;
assign w19897 = ~w19895 & w48954;
assign w19898 = w19874 & ~w19897;
assign w19899 = ~w18860 & w41736;
assign w19900 = w18826 & ~w19034;
assign w19901 = w18537 & w19900;
assign w19902 = ~w19899 & ~w19901;
assign w19903 = w18989 & w19005;
assign w19904 = ~w18997 & w19903;
assign w19905 = ~w19028 & w19904;
assign w19906 = w400 & ~w19039;
assign w19907 = ~w19902 & w19906;
assign w19908 = ~w19901 & w41737;
assign w19909 = ~w351 & ~w18996;
assign w19910 = ~w19907 & w41738;
assign w19911 = ~w351 & w18996;
assign w19912 = (w19911 & w19907) | (w19911 & w41739) | (w19907 & w41739);
assign w19913 = ~w19910 & ~w19912;
assign w19914 = w252 & w19894;
assign w19915 = w252 & w19889;
assign w19916 = w19880 & w19915;
assign w19917 = ~w19914 & ~w19916;
assign w19918 = w19913 & w19917;
assign w19919 = w19898 & ~w19918;
assign w19920 = w19865 & ~w19919;
assign w19921 = w19854 & ~w19920;
assign w19922 = (w3 & w19841) | (w3 & w45089) | (w19841 & w45089);
assign w19923 = w19826 & w19922;
assign w19924 = (~w18918 & ~w19837) | (~w18918 & w45090) | (~w19837 & w45090);
assign w19925 = w42 & ~w18885;
assign w19926 = ~w18888 & ~w19925;
assign w19927 = w19924 & w19926;
assign w19928 = w18896 & ~w19926;
assign w19929 = ~w19924 & w19928;
assign w19930 = ~w19927 & ~w19929;
assign w19931 = (w42 & w19841) | (w42 & w41740) | (w19841 & w41740);
assign w19932 = w19930 & ~w19931;
assign w19933 = w493 & w19030;
assign w19934 = ~w493 & ~w19039;
assign w19935 = ~w19423 & w19934;
assign w19936 = ~w19933 & ~w19935;
assign w19937 = w19033 & ~w19936;
assign w19938 = ~w19033 & w19936;
assign w19939 = ~w19937 & ~w19938;
assign w19940 = w400 & ~w19939;
assign w19941 = w19932 & ~w19940;
assign w19942 = ~w19923 & w19941;
assign w19943 = (w19942 & w19920) | (w19942 & w41741) | (w19920 & w41741);
assign w19944 = ~w19814 & w19943;
assign w19945 = w612 & w19796;
assign w19946 = ~w19944 & ~w19945;
assign w19947 = ~w19286 & w48955;
assign w19948 = ~w19763 & ~w19765;
assign w19949 = ~w1120 & ~w19766;
assign w19950 = ~w19763 & w41742;
assign w19951 = ~w1120 & w19766;
assign w19952 = (w19951 & w19763) | (w19951 & w41743) | (w19763 & w41743);
assign w19953 = ~w19950 & ~w19952;
assign w19954 = ~w19947 & w19953;
assign w19955 = w19759 & w19954;
assign w19956 = ~w612 & w19955;
assign w19957 = w19945 & ~w19955;
assign w19958 = ~w19956 & ~w19957;
assign w19959 = w351 & w18996;
assign w19960 = ~w19907 & w41744;
assign w19961 = w351 & ~w18996;
assign w19962 = (w19961 & w19907) | (w19961 & w41745) | (w19907 & w41745);
assign w19963 = ~w19960 & ~w19962;
assign w19964 = ~w400 & ~w19033;
assign w19965 = ~w19936 & w19964;
assign w19966 = ~w400 & w19033;
assign w19967 = w19936 & w19966;
assign w19968 = ~w19965 & ~w19967;
assign w19969 = w19963 & w19968;
assign w19970 = w19918 & ~w19969;
assign w19971 = w19898 & ~w19970;
assign w19972 = w19865 & ~w19971;
assign w19973 = ~w19923 & w19932;
assign w19974 = (w19973 & w19972) | (w19973 & w41746) | (w19972 & w41746);
assign w19975 = (w612 & ~w19060) | (w612 & w48956) | (~w19060 & w48956);
assign w19976 = w493 & ~w19800;
assign w19977 = ~w19803 & ~w19976;
assign w19978 = ~w19798 & w48957;
assign w19979 = (w19977 & w19798) | (w19977 & w48958) | (w19798 & w48958);
assign w19980 = ~w19978 & ~w19979;
assign w19981 = ~w19975 & ~w19980;
assign w19982 = w19955 & w19981;
assign w19983 = w19942 & ~w19982;
assign w19984 = ~w19921 & w19983;
assign w19985 = ~w19814 & w19984;
assign w19986 = (~w19974 & ~w19984) | (~w19974 & w41747) | (~w19984 & w41747);
assign w19987 = ~w19797 & w19986;
assign w19988 = (~w19958 & w19736) | (~w19958 & w45091) | (w19736 & w45091);
assign w19989 = w19987 & ~w19988;
assign w19990 = w19737 & ~w19946;
assign w19991 = w19989 & ~w19990;
assign w19992 = w19062 & ~w19991;
assign w19993 = ~w19062 & w19991;
assign w19994 = ~w19992 & ~w19993;
assign w19995 = ~w493 & ~w19994;
assign w19996 = ~w19735 & w19986;
assign w19997 = w19708 & w19996;
assign w19998 = ~w19293 & w19944;
assign w19999 = w19986 & ~w19998;
assign w20000 = (~w19999 & ~w19996) | (~w19999 & w41748) | (~w19996 & w41748);
assign w20001 = w19776 & ~w19954;
assign w20002 = (~w20001 & w19732) | (~w20001 & w41749) | (w19732 & w41749);
assign w20003 = w19293 & w19954;
assign w20004 = w19776 & ~w20003;
assign w20005 = w19708 & w20002;
assign w20006 = w19753 & w19786;
assign w20007 = ~w20005 & w45092;
assign w20008 = ~w754 & w20000;
assign w20009 = w19753 & ~w20000;
assign w20010 = ~w20007 & w20009;
assign w20011 = ~w19758 & ~w19795;
assign w20012 = ~w20010 & w45093;
assign w20013 = (w20011 & w20010) | (w20011 & w45094) | (w20010 & w45094);
assign w20014 = ~w20012 & ~w20013;
assign w20015 = ~w612 & w20014;
assign w20016 = ~w19995 & ~w20015;
assign w20017 = w493 & w19994;
assign w20018 = w19955 & ~w19975;
assign w20019 = w19062 & ~w19945;
assign w20020 = ~w19797 & ~w20019;
assign w20021 = ~w20018 & w20020;
assign w20022 = ~w19293 & w20020;
assign w20023 = (~w20021 & w19736) | (~w20021 & w45095) | (w19736 & w45095);
assign w20024 = ~w19980 & w20023;
assign w20025 = w19980 & ~w20023;
assign w20026 = ~w20024 & ~w20025;
assign w20027 = ~w19811 & w20000;
assign w20028 = ~w20000 & w20026;
assign w20029 = ~w20027 & ~w20028;
assign w20030 = ~w400 & w20029;
assign w20031 = ~w20017 & ~w20030;
assign w20032 = ~w20016 & w20031;
assign w20033 = ~w19736 & w19998;
assign w20034 = ~w4838 & w19658;
assign w20035 = w19671 & w20034;
assign w20036 = (~w19659 & ~w20034) | (~w19659 & w41750) | (~w20034 & w41750);
assign w20037 = ~w19703 & w20036;
assign w20038 = w19629 & ~w20037;
assign w20039 = (w20035 & w19418) | (w20035 & w41751) | (w19418 & w41751);
assign w20040 = w19704 & ~w20039;
assign w20041 = ~w19618 & w20038;
assign w20042 = w20040 & ~w20041;
assign w20043 = w19732 & w20042;
assign w20044 = w19124 & w19733;
assign w20045 = ~w19216 & ~w19684;
assign w20046 = w19986 & w20045;
assign w20047 = ~w20043 & w41752;
assign w20048 = w20046 & ~w20047;
assign w20049 = ~w1541 & w20000;
assign w20050 = ~w20033 & w20048;
assign w20051 = ~w20049 & ~w20050;
assign w20052 = ~w19202 & ~w19275;
assign w20053 = ~w1320 & ~w20052;
assign w20054 = ~w20051 & w20053;
assign w20055 = ~w1320 & w20052;
assign w20056 = w20051 & w20055;
assign w20057 = ~w20054 & ~w20056;
assign w20058 = w19215 & w19685;
assign w20059 = ~w19275 & ~w20058;
assign w20060 = ~w19275 & w19734;
assign w20061 = (~w20059 & w20043) | (~w20059 & w45096) | (w20043 & w45096);
assign w20062 = w19124 & ~w19683;
assign w20063 = ~w19202 & ~w19210;
assign w20064 = ~w20062 & w20063;
assign w20065 = (w20064 & w20043) | (w20064 & w41753) | (w20043 & w41753);
assign w20066 = ~w20061 & ~w20065;
assign w20067 = ~w20033 & w20066;
assign w20068 = w20066 & w41754;
assign w20069 = w1320 & w20000;
assign w20070 = ~w19288 & ~w19947;
assign w20071 = w1120 & ~w20070;
assign w20072 = (w20071 & ~w20000) | (w20071 & w45097) | (~w20000 & w45097);
assign w20073 = ~w20068 & w20072;
assign w20074 = w1120 & ~w19947;
assign w20075 = w20000 & w45098;
assign w20076 = w19986 & w20070;
assign w20077 = w1120 & w20076;
assign w20078 = w20066 & w41755;
assign w20079 = ~w20075 & ~w20078;
assign w20080 = ~w20073 & w20079;
assign w20081 = w20057 & w20080;
assign w20082 = ~w19944 & ~w19974;
assign w20083 = w1120 & w20082;
assign w20084 = w19766 & ~w19948;
assign w20085 = ~w19766 & w19948;
assign w20086 = ~w20084 & ~w20085;
assign w20087 = w20083 & ~w20086;
assign w20088 = ~w20083 & w20086;
assign w20089 = ~w20087 & ~w20088;
assign w20090 = ~w1120 & w19947;
assign w20091 = ~w20074 & ~w20090;
assign w20092 = w19986 & w20091;
assign w20093 = w20086 & ~w20092;
assign w20094 = ~w20086 & w20092;
assign w20095 = ~w20093 & ~w20094;
assign w20096 = w19737 & ~w20089;
assign w20097 = ~w19737 & ~w20095;
assign w20098 = ~w20096 & ~w20097;
assign w20099 = ~w945 & w20098;
assign w20100 = (~w1120 & ~w20000) | (~w1120 & w45099) | (~w20000 & w45099);
assign w20101 = ~w20066 & w41756;
assign w20102 = w20100 & ~w20101;
assign w20103 = w20067 & w20076;
assign w20104 = w20102 & ~w20103;
assign w20105 = ~w20099 & ~w20104;
assign w20106 = ~w20081 & w20105;
assign w20107 = ~w945 & w20057;
assign w20108 = w20106 & ~w20107;
assign w20109 = (~w20098 & ~w20079) | (~w20098 & w45100) | (~w20079 & w45100);
assign w20110 = w945 & ~w20098;
assign w20111 = (~w20006 & w20005) | (~w20006 & w45101) | (w20005 & w45101);
assign w20112 = ~w945 & w19753;
assign w20113 = w19786 & ~w20112;
assign w20114 = w20000 & w20113;
assign w20115 = ~w20007 & ~w20111;
assign w20116 = ~w20000 & w20115;
assign w20117 = ~w20114 & ~w20116;
assign w20118 = ~w754 & w20117;
assign w20119 = ~w20109 & ~w20118;
assign w20120 = ~w20110 & w20119;
assign w20121 = ~w20108 & w20120;
assign w20122 = w19683 & w20044;
assign w20123 = w2006 & w19213;
assign w20124 = ~w2006 & ~w19213;
assign w20125 = ~w20123 & ~w20124;
assign w20126 = w20062 & ~w20125;
assign w20127 = ~w20062 & w20125;
assign w20128 = ~w20126 & ~w20127;
assign w20129 = ~w20043 & w41757;
assign w20130 = (w20128 & w20043) | (w20128 & w41758) | (w20043 & w41758);
assign w20131 = ~w20129 & ~w20130;
assign w20132 = ~w19213 & w20000;
assign w20133 = ~w20000 & ~w20131;
assign w20134 = ~w20132 & ~w20133;
assign w20135 = ~w1738 & ~w20134;
assign w20136 = w19170 & w20044;
assign w20137 = ~w20062 & ~w20123;
assign w20138 = w19170 & ~w20137;
assign w20139 = w19144 & ~w20138;
assign w20140 = (w20139 & w20043) | (w20139 & w45102) | (w20043 & w45102);
assign w20141 = w19208 & ~w20062;
assign w20142 = (w20141 & w20043) | (w20141 & w41759) | (w20043 & w41759);
assign w20143 = w20140 & ~w20142;
assign w20144 = ~w20000 & w20143;
assign w20145 = ~w1541 & w19163;
assign w20146 = (w20145 & ~w20143) | (w20145 & w41760) | (~w20143 & w41760);
assign w20147 = ~w1541 & ~w19163;
assign w20148 = w20143 & w41761;
assign w20149 = ~w20146 & ~w20148;
assign w20150 = ~w20135 & w20149;
assign w20151 = w1738 & w20134;
assign w20152 = w19122 & w19733;
assign w20153 = ~w20043 & w20152;
assign w20154 = ~w19185 & ~w19682;
assign w20155 = ~w19186 & w20154;
assign w20156 = w19122 & ~w20155;
assign w20157 = ~w19103 & ~w20156;
assign w20158 = w19986 & w20157;
assign w20159 = ~w20153 & w20158;
assign w20160 = ~w20033 & w20159;
assign w20161 = ~w2285 & w20000;
assign w20162 = ~w20160 & ~w20161;
assign w20163 = ~w19080 & ~w19082;
assign w20164 = w2006 & w20163;
assign w20165 = ~w20162 & w20164;
assign w20166 = w2006 & ~w20163;
assign w20167 = w20162 & w20166;
assign w20168 = ~w20165 & ~w20167;
assign w20169 = ~w20151 & w20168;
assign w20170 = w20150 & ~w20169;
assign w20171 = ~w19120 & ~w19999;
assign w20172 = ~w19997 & w20171;
assign w20173 = ~w19119 & ~w19186;
assign w20174 = w19733 & w20154;
assign w20175 = w20173 & w20174;
assign w20176 = ~w19103 & ~w19121;
assign w20177 = ~w19119 & ~w20155;
assign w20178 = w20176 & ~w20177;
assign w20179 = ~w20176 & w20177;
assign w20180 = ~w20178 & ~w20179;
assign w20181 = ~w20043 & w45103;
assign w20182 = (w20180 & w20043) | (w20180 & w45104) | (w20043 & w45104);
assign w20183 = ~w20181 & ~w20182;
assign w20184 = ~w20000 & ~w20183;
assign w20185 = ~w20172 & ~w20184;
assign w20186 = (~w2285 & w20184) | (~w2285 & w41762) | (w20184 & w41762);
assign w20187 = (w2285 & w19997) | (w2285 & w41763) | (w19997 & w41763);
assign w20188 = ~w20184 & w20187;
assign w20189 = ~w20154 & ~w20173;
assign w20190 = w20154 & w20173;
assign w20191 = ~w20189 & ~w20190;
assign w20192 = (w20191 & w20043) | (w20191 & w41764) | (w20043 & w41764);
assign w20193 = (w19986 & w20043) | (w19986 & w45105) | (w20043 & w45105);
assign w20194 = ~w20192 & w20193;
assign w20195 = ~w20033 & w20194;
assign w20196 = ~w19118 & ~w19999;
assign w20197 = ~w19997 & w20196;
assign w20198 = (w2558 & w19997) | (w2558 & w41765) | (w19997 & w41765);
assign w20199 = ~w20195 & w20198;
assign w20200 = ~w20188 & w20199;
assign w20201 = ~w20186 & ~w20200;
assign w20202 = ~w2006 & ~w20163;
assign w20203 = ~w20162 & w20202;
assign w20204 = ~w2006 & w20163;
assign w20205 = w20162 & w20204;
assign w20206 = ~w20203 & ~w20205;
assign w20207 = w20201 & w20206;
assign w20208 = ~w20195 & ~w20197;
assign w20209 = (~w2558 & w20195) | (~w2558 & w41766) | (w20195 & w41766);
assign w20210 = ~w20188 & ~w20209;
assign w20211 = w20150 & ~w20210;
assign w20212 = w20207 & w20211;
assign w20213 = ~w20170 & ~w20212;
assign w20214 = w20051 & ~w20052;
assign w20215 = ~w20051 & w20052;
assign w20216 = ~w20214 & ~w20215;
assign w20217 = w1320 & ~w20216;
assign w20218 = ~w19163 & w20144;
assign w20219 = w1541 & ~w20218;
assign w20220 = w19163 & ~w20144;
assign w20221 = w20219 & ~w20220;
assign w20222 = w20105 & ~w20217;
assign w20223 = ~w20221 & w20222;
assign w20224 = w20213 & w20223;
assign w20225 = w612 & ~w20014;
assign w20226 = w754 & ~w20117;
assign w20227 = ~w20225 & ~w20226;
assign w20228 = w20031 & w20227;
assign w20229 = (w20228 & w20224) | (w20228 & w41767) | (w20224 & w41767);
assign w20230 = ~w19185 & ~w19258;
assign w20231 = ~w19271 & ~w19676;
assign w20232 = ~w19259 & ~w19681;
assign w20233 = ~w19259 & w20231;
assign w20234 = (~w20232 & w20043) | (~w20232 & w41768) | (w20043 & w41768);
assign w20235 = ~w20230 & ~w20234;
assign w20236 = w20230 & w20234;
assign w20237 = ~w19184 & w20000;
assign w20238 = ~w20000 & ~w20235;
assign w20239 = ~w20236 & w20238;
assign w20240 = ~w20237 & ~w20239;
assign w20241 = ~w20239 & w45106;
assign w20242 = w4056 & w20000;
assign w20243 = ~w19271 & ~w20043;
assign w20244 = ~w20000 & w20243;
assign w20245 = ~w20242 & ~w20244;
assign w20246 = w19257 & ~w19676;
assign w20247 = ~w3646 & w20246;
assign w20248 = w20245 & w20247;
assign w20249 = ~w3646 & ~w20246;
assign w20250 = ~w20245 & w20249;
assign w20251 = ~w20248 & ~w20250;
assign w20252 = ~w20241 & w20251;
assign w20253 = (w19257 & w20043) | (w19257 & w45107) | (w20043 & w45107);
assign w20254 = w3646 & w20000;
assign w20255 = ~w20000 & w20253;
assign w20256 = ~w20254 & ~w20255;
assign w20257 = ~w19245 & ~w19259;
assign w20258 = ~w3242 & w20257;
assign w20259 = ~w20256 & w20258;
assign w20260 = ~w3242 & ~w20257;
assign w20261 = w20256 & w20260;
assign w20262 = ~w20259 & ~w20261;
assign w20263 = w20252 & w20262;
assign w20264 = w19364 & ~w19410;
assign w20265 = ~w19618 & ~w19625;
assign w20266 = ~w19618 & w45108;
assign w20267 = ~w19345 & w19383;
assign w20268 = ~w19414 & ~w20267;
assign w20269 = w19405 & ~w19414;
assign w20270 = ~w20266 & w20269;
assign w20271 = ~w20268 & ~w20270;
assign w20272 = w20264 & ~w20271;
assign w20273 = ~w20264 & w20271;
assign w20274 = ~w20272 & ~w20273;
assign w20275 = w19409 & w20000;
assign w20276 = ~w20000 & w20274;
assign w20277 = ~w20275 & ~w20276;
assign w20278 = w6264 & w20277;
assign w20279 = w6264 & ~w19631;
assign w20280 = ~w6264 & w19631;
assign w20281 = ~w20279 & ~w20280;
assign w20282 = ~w18393 & w19040;
assign w20283 = ~w19040 & w19652;
assign w20284 = ~w20282 & ~w20283;
assign w20285 = ~w20000 & w45109;
assign w20286 = (~w20284 & w20000) | (~w20284 & w45110) | (w20000 & w45110);
assign w20287 = ~w20285 & ~w20286;
assign w20288 = ~w5745 & w20287;
assign w20289 = ~w20278 & ~w20288;
assign w20290 = ~w19631 & w20035;
assign w20291 = ~w19703 & ~w19713;
assign w20292 = ~w19726 & w20291;
assign w20293 = w19631 & w19710;
assign w20294 = w20292 & ~w20293;
assign w20295 = ~w20290 & w20294;
assign w20296 = w4430 & w19722;
assign w20297 = (w20296 & w20000) | (w20296 & w45111) | (w20000 & w45111);
assign w20298 = w4430 & ~w19722;
assign w20299 = ~w20000 & w45112;
assign w20300 = ~w20297 & ~w20299;
assign w20301 = ~w19271 & ~w19659;
assign w20302 = ~w19703 & w19732;
assign w20303 = (w20301 & ~w20302) | (w20301 & w41769) | (~w20302 & w41769);
assign w20304 = w20302 & w41770;
assign w20305 = ~w20303 & ~w20304;
assign w20306 = w19270 & w20000;
assign w20307 = ~w20000 & ~w20305;
assign w20308 = ~w20306 & ~w20307;
assign w20309 = w4056 & w20308;
assign w20310 = w20300 & ~w20309;
assign w20311 = ~w19696 & w19986;
assign w20312 = ~w19631 & w19658;
assign w20313 = w20311 & ~w20312;
assign w20314 = (w20313 & w19736) | (w20313 & w45113) | (w19736 & w45113);
assign w20315 = ~w5330 & ~w19999;
assign w20316 = ~w19997 & w20315;
assign w20317 = w19671 & w19701;
assign w20318 = ~w4838 & ~w20317;
assign w20319 = (~w20318 & w19997) | (~w20318 & w41771) | (w19997 & w41771);
assign w20320 = ~w4838 & w20317;
assign w20321 = ~w19997 & w41772;
assign w20322 = w20313 & ~w20320;
assign w20323 = ~w20033 & w20322;
assign w20324 = ~w20321 & ~w20323;
assign w20325 = ~w20314 & w20319;
assign w20326 = w20324 & ~w20325;
assign w20327 = w19694 & w19986;
assign w20328 = ~w19631 & w19657;
assign w20329 = w20327 & ~w20328;
assign w20330 = (w20329 & w19736) | (w20329 & w45114) | (w19736 & w45114);
assign w20331 = w5745 & ~w19999;
assign w20332 = ~w19997 & w20331;
assign w20333 = w19645 & w19689;
assign w20334 = w5330 & ~w20333;
assign w20335 = (w20334 & w19997) | (w20334 & w41773) | (w19997 & w41773);
assign w20336 = ~w20330 & w20335;
assign w20337 = w5330 & w20333;
assign w20338 = w20329 & w20337;
assign w20339 = ~w20033 & w20338;
assign w20340 = ~w19997 & w41774;
assign w20341 = ~w20339 & ~w20340;
assign w20342 = ~w20336 & w20341;
assign w20343 = ~w20326 & w20342;
assign w20344 = w20310 & w20343;
assign w20345 = w20289 & w20344;
assign w20346 = w20263 & w20345;
assign w20347 = w5745 & ~w20287;
assign w20348 = ~w20330 & ~w20332;
assign w20349 = ~w5330 & ~w20333;
assign w20350 = (w20349 & w20332) | (w20349 & w45115) | (w20332 & w45115);
assign w20351 = ~w5330 & w20333;
assign w20352 = ~w20332 & w45116;
assign w20353 = ~w20350 & ~w20352;
assign w20354 = ~w20347 & w20353;
assign w20355 = w20344 & ~w20354;
assign w20356 = ~w4430 & ~w19722;
assign w20357 = (w20356 & w20000) | (w20356 & w45117) | (w20000 & w45117);
assign w20358 = ~w4430 & w19722;
assign w20359 = ~w20000 & w45118;
assign w20360 = ~w20357 & ~w20359;
assign w20361 = w4838 & w20317;
assign w20362 = (w20361 & w19997) | (w20361 & w41775) | (w19997 & w41775);
assign w20363 = ~w20314 & w20362;
assign w20364 = w4838 & ~w20317;
assign w20365 = w20313 & w20364;
assign w20366 = ~w20033 & w20365;
assign w20367 = ~w19997 & w41776;
assign w20368 = ~w20366 & ~w20367;
assign w20369 = ~w20363 & w20368;
assign w20370 = w20360 & w20369;
assign w20371 = w20310 & ~w20370;
assign w20372 = ~w4056 & ~w20308;
assign w20373 = w3646 & ~w20246;
assign w20374 = w20245 & w20373;
assign w20375 = w3646 & w20246;
assign w20376 = ~w20245 & w20375;
assign w20377 = ~w20374 & ~w20376;
assign w20378 = ~w20372 & w20377;
assign w20379 = ~w20371 & w20378;
assign w20380 = ~w20355 & w20379;
assign w20381 = w20263 & ~w20380;
assign w20382 = w20256 & ~w20257;
assign w20383 = ~w20256 & w20257;
assign w20384 = ~w20382 & ~w20383;
assign w20385 = w3242 & w20384;
assign w20386 = (~w2896 & w20239) | (~w2896 & w45119) | (w20239 & w45119);
assign w20387 = ~w20241 & ~w20386;
assign w20388 = ~w20385 & w20387;
assign w20389 = (~w20241 & w20385) | (~w20241 & w45120) | (w20385 & w45120);
assign w20390 = w20201 & w41777;
assign w20391 = ~w20170 & ~w20390;
assign w20392 = ~w20389 & ~w20391;
assign w20393 = w20121 & w20392;
assign w20394 = ~w20346 & ~w20381;
assign w20395 = w20393 & w20394;
assign w20396 = w20229 & ~w20395;
assign w20397 = ~w19467 & ~w19478;
assign w20398 = ~w19040 & w20397;
assign w20399 = w19040 & ~w20397;
assign w20400 = ~w20398 & ~w20399;
assign w20401 = ~a[38] & ~w19040;
assign w20402 = a[39] & ~w20401;
assign w20403 = ~a[39] & w20401;
assign w20404 = ~w20402 & ~w20403;
assign w20405 = ~w20000 & w20400;
assign w20406 = w20000 & w20404;
assign w20407 = ~w20405 & ~w20406;
assign w20408 = a[38] & w18183;
assign w20409 = ~a[34] & ~a[35];
assign w20410 = ~a[36] & w20409;
assign w20411 = ~w20408 & w20410;
assign w20412 = w19040 & ~w20411;
assign w20413 = ~a[35] & ~w19040;
assign w20414 = ~a[34] & w20413;
assign w20415 = ~a[36] & w20414;
assign w20416 = a[37] & ~w20415;
assign w20417 = ~w20412 & ~w20416;
assign w20418 = ~w18183 & w20417;
assign w20419 = w20401 & ~w20418;
assign w20420 = ~a[38] & ~w18183;
assign w20421 = ~w18183 & ~w19040;
assign w20422 = ~w20420 & ~w20421;
assign w20423 = ~w20417 & w20422;
assign w20424 = ~w20419 & ~w20423;
assign w20425 = ~a[36] & ~a[38];
assign w20426 = ~a[37] & ~w20425;
assign w20427 = w20415 & w20426;
assign w20428 = w20408 & ~w20427;
assign w20429 = w19040 & ~w20410;
assign w20430 = ~w20420 & w20429;
assign w20431 = a[37] & ~w20430;
assign w20432 = w20409 & w20421;
assign w20433 = ~w20426 & ~w20432;
assign w20434 = ~w20431 & w20433;
assign w20435 = ~w20428 & ~w20434;
assign w20436 = ~w17380 & ~w20424;
assign w20437 = w20000 & w20436;
assign w20438 = ~w17380 & ~w20435;
assign w20439 = ~w20000 & w20438;
assign w20440 = ~w20437 & ~w20439;
assign w20441 = ~w20407 & w20440;
assign w20442 = ~w19040 & w19471;
assign w20443 = w19040 & w19477;
assign w20444 = ~w20442 & ~w20443;
assign w20445 = w19040 & w19478;
assign w20446 = ~w19464 & ~w20445;
assign w20447 = ~w19040 & w19468;
assign w20448 = w20446 & ~w20447;
assign w20449 = w17380 & ~w20448;
assign w20450 = ~w17380 & w20448;
assign w20451 = ~w20449 & ~w20450;
assign w20452 = ~w19974 & w20451;
assign w20453 = ~w19985 & w20452;
assign w20454 = ~w16559 & w20444;
assign w20455 = w20453 & ~w20454;
assign w20456 = ~w19998 & w20453;
assign w20457 = ~w19735 & w20453;
assign w20458 = w19708 & w20457;
assign w20459 = ~w20456 & ~w20458;
assign w20460 = ~w16559 & ~w20444;
assign w20461 = ~w20458 & w41778;
assign w20462 = (w20455 & w19736) | (w20455 & w48959) | (w19736 & w48959);
assign w20463 = ~w20461 & ~w20462;
assign w20464 = w17380 & w20424;
assign w20465 = w20000 & w20464;
assign w20466 = w17380 & w20435;
assign w20467 = ~w20000 & w20466;
assign w20468 = ~w20465 & ~w20467;
assign w20469 = ~w20463 & w20468;
assign w20470 = ~w20441 & w20469;
assign w20471 = w16559 & ~w20444;
assign w20472 = (w20471 & w20458) | (w20471 & w41779) | (w20458 & w41779);
assign w20473 = w16559 & w20444;
assign w20474 = ~w20458 & w41780;
assign w20475 = ~w20472 & ~w20474;
assign w20476 = ~w19487 & ~w19509;
assign w20477 = ~w19974 & w20476;
assign w20478 = ~w19985 & w20477;
assign w20479 = ~w19998 & w20478;
assign w20480 = ~w19735 & w20478;
assign w20481 = w19708 & w20480;
assign w20482 = ~w19448 & ~w19461;
assign w20483 = w15681 & w20482;
assign w20484 = (w20483 & w20481) | (w20483 & w41781) | (w20481 & w41781);
assign w20485 = w15681 & ~w20482;
assign w20486 = ~w20481 & w41782;
assign w20487 = ~w20484 & ~w20486;
assign w20488 = w20475 & w20487;
assign w20489 = ~w20470 & w20488;
assign w20490 = ~w19489 & ~w19509;
assign w20491 = ~w19974 & w20490;
assign w20492 = ~w19985 & w20491;
assign w20493 = ~w19998 & w20492;
assign w20494 = ~w19735 & w20492;
assign w20495 = (~w20493 & ~w20494) | (~w20493 & w45121) | (~w20494 & w45121);
assign w20496 = w15681 & ~w19999;
assign w20497 = ~w19997 & w20496;
assign w20498 = w20495 & ~w20497;
assign w20499 = w19515 & w19524;
assign w20500 = w14766 & ~w20499;
assign w20501 = w14766 & w20499;
assign w20502 = (w20500 & w20497) | (w20500 & w45122) | (w20497 & w45122);
assign w20503 = ~w20497 & w45123;
assign w20504 = ~w20502 & ~w20503;
assign w20505 = w18467 & ~w19502;
assign w20506 = ~w18467 & w19502;
assign w20507 = ~w20505 & ~w20506;
assign w20508 = w19524 & ~w20490;
assign w20509 = w19515 & ~w20508;
assign w20510 = ~w14766 & ~w20509;
assign w20511 = w14766 & w20509;
assign w20512 = ~w20510 & ~w20511;
assign w20513 = ~w20000 & w20512;
assign w20514 = ~w20507 & ~w20513;
assign w20515 = w20507 & w20513;
assign w20516 = ~w20514 & ~w20515;
assign w20517 = ~w14766 & w20499;
assign w20518 = (w20517 & w20497) | (w20517 & w45124) | (w20497 & w45124);
assign w20519 = ~w14766 & ~w20499;
assign w20520 = ~w20497 & w45125;
assign w20521 = ~w20518 & ~w20520;
assign w20522 = ~w14039 & w20521;
assign w20523 = ~w20481 & w41783;
assign w20524 = (w20482 & w20481) | (w20482 & w41784) | (w20481 & w41784);
assign w20525 = ~w20523 & ~w20524;
assign w20526 = ~w15681 & w20525;
assign w20527 = w20504 & w20526;
assign w20528 = w20522 & ~w20527;
assign w20529 = w20516 & ~w20528;
assign w20530 = w20504 & w20516;
assign w20531 = w20489 & w20530;
assign w20532 = ~w20529 & ~w20531;
assign w20533 = w20521 & ~w20526;
assign w20534 = w14039 & ~w20501;
assign w20535 = ~w20497 & w45126;
assign w20536 = w14039 & ~w20500;
assign w20537 = (w20536 & w20497) | (w20536 & w45127) | (w20497 & w45127);
assign w20538 = ~w20535 & ~w20537;
assign w20539 = ~w20533 & ~w20538;
assign w20540 = w20488 & ~w20538;
assign w20541 = ~w20470 & w20540;
assign w20542 = ~w20539 & ~w20541;
assign w20543 = ~w19500 & ~w19519;
assign w20544 = ~w20507 & ~w20510;
assign w20545 = ~w20511 & ~w20544;
assign w20546 = w20543 & ~w20545;
assign w20547 = ~w20543 & w20545;
assign w20548 = ~w20546 & ~w20547;
assign w20549 = ~w19499 & w20000;
assign w20550 = ~w20000 & ~w20548;
assign w20551 = ~w20549 & ~w20550;
assign w20552 = ~w13384 & ~w20551;
assign w20553 = ~w19597 & w19602;
assign w20554 = w19532 & ~w20553;
assign w20555 = ~w19532 & w20553;
assign w20556 = ~w20554 & ~w20555;
assign w20557 = w19596 & w20000;
assign w20558 = w12666 & ~w20557;
assign w20559 = ~w20000 & w20556;
assign w20560 = w20558 & ~w20559;
assign w20561 = ~w20552 & ~w20560;
assign w20562 = w19577 & ~w19612;
assign w20563 = w19587 & ~w19608;
assign w20564 = w19587 & ~w19597;
assign w20565 = (w20564 & w19518) | (w20564 & w45128) | (w19518 & w45128);
assign w20566 = ~w20563 & ~w20565;
assign w20567 = w20562 & w20566;
assign w20568 = ~w20562 & ~w20566;
assign w20569 = ~w20567 & ~w20568;
assign w20570 = ~w12666 & w19040;
assign w20571 = ~w19040 & w19534;
assign w20572 = ~w20570 & ~w20571;
assign w20573 = w19570 & ~w20572;
assign w20574 = ~w19570 & w20572;
assign w20575 = ~w20573 & ~w20574;
assign w20576 = ~w20000 & w20569;
assign w20577 = w20000 & ~w20575;
assign w20578 = ~w20576 & ~w20577;
assign w20579 = ~w11138 & ~w20578;
assign w20580 = w19587 & w19607;
assign w20581 = w19602 & ~w20555;
assign w20582 = w20580 & ~w20581;
assign w20583 = ~w20580 & w20581;
assign w20584 = ~w20582 & ~w20583;
assign w20585 = w18511 & w19040;
assign w20586 = ~w19040 & ~w19582;
assign w20587 = ~w20585 & ~w20586;
assign w20588 = ~w20000 & w20584;
assign w20589 = w20000 & w20587;
assign w20590 = ~w20588 & ~w20589;
assign w20591 = w11870 & w20590;
assign w20592 = w19577 & ~w20567;
assign w20593 = ~w19553 & ~w19613;
assign w20594 = w20592 & ~w20593;
assign w20595 = ~w20592 & w20593;
assign w20596 = ~w20594 & ~w20595;
assign w20597 = ~w19552 & w20000;
assign w20598 = ~w20000 & ~w20596;
assign w20599 = ~w20597 & ~w20598;
assign w20600 = w10419 & w20599;
assign w20601 = ~w20591 & ~w20600;
assign w20602 = ~w20579 & w20601;
assign w20603 = w20561 & w20602;
assign w20604 = w20542 & w20603;
assign w20605 = w20532 & w20604;
assign w20606 = ~w19532 & ~w19974;
assign w20607 = ~w19985 & w20606;
assign w20608 = ~w19998 & w20607;
assign w20609 = ~w19735 & w20607;
assign w20610 = (~w20608 & ~w20609) | (~w20608 & w45129) | (~w20609 & w45129);
assign w20611 = w13384 & ~w19999;
assign w20612 = ~w19997 & w20611;
assign w20613 = w20610 & ~w20612;
assign w20614 = ~w12666 & ~w20553;
assign w20615 = (w20614 & w20612) | (w20614 & w45130) | (w20612 & w45130);
assign w20616 = ~w12666 & w20553;
assign w20617 = ~w20612 & w45131;
assign w20618 = ~w20615 & ~w20617;
assign w20619 = ~w11870 & ~w20590;
assign w20620 = w20618 & ~w20619;
assign w20621 = w13384 & w20551;
assign w20622 = ~w20560 & w20621;
assign w20623 = w20620 & ~w20622;
assign w20624 = w20602 & ~w20623;
assign w20625 = w19620 & ~w19627;
assign w20626 = ~w19293 & w20625;
assign w20627 = ~w19293 & w19626;
assign w20628 = ~w20082 & w20627;
assign w20629 = ~w20626 & ~w20628;
assign w20630 = w19627 & ~w20265;
assign w20631 = ~w20266 & ~w20630;
assign w20632 = ~w19398 & ~w20631;
assign w20633 = w19626 & ~w19986;
assign w20634 = w20632 & ~w20633;
assign w20635 = ~w19736 & ~w20629;
assign w20636 = w20634 & ~w20635;
assign w20637 = w19626 & w20265;
assign w20638 = (~w20637 & w19997) | (~w20637 & w41785) | (w19997 & w41785);
assign w20639 = w9195 & w19398;
assign w20640 = (~w20639 & w19997) | (~w20639 & w41786) | (w19997 & w41786);
assign w20641 = ~w20635 & w45132;
assign w20642 = w20638 & ~w20640;
assign w20643 = ~w20641 & ~w20642;
assign w20644 = ~w18192 & w19040;
assign w20645 = ~w19040 & ~w19318;
assign w20646 = ~w20644 & ~w20645;
assign w20647 = w19323 & w19403;
assign w20648 = ~w19398 & ~w20266;
assign w20649 = ~w20647 & ~w20648;
assign w20650 = ~w19398 & w20647;
assign w20651 = ~w20266 & w20650;
assign w20652 = w20000 & w20646;
assign w20653 = ~w20649 & ~w20651;
assign w20654 = ~w20000 & w20653;
assign w20655 = ~w20652 & ~w20654;
assign w20656 = ~w8666 & ~w20655;
assign w20657 = w20643 & ~w20656;
assign w20658 = ~w19398 & ~w20000;
assign w20659 = w20638 & ~w20658;
assign w20660 = (~w9195 & w20635) | (~w9195 & w45133) | (w20635 & w45133);
assign w20661 = ~w20659 & w20660;
assign w20662 = ~w19553 & w19577;
assign w20663 = ~w20567 & w20662;
assign w20664 = ~w19613 & ~w20663;
assign w20665 = w19986 & ~w20664;
assign w20666 = (w20665 & w19736) | (w20665 & w45134) | (w19736 & w45134);
assign w20667 = ~w19564 & ~w19620;
assign w20668 = ~w9781 & w20667;
assign w20669 = (w20668 & w19997) | (w20668 & w41787) | (w19997 & w41787);
assign w20670 = ~w20666 & w20669;
assign w20671 = ~w9781 & ~w20667;
assign w20672 = w20665 & w20671;
assign w20673 = ~w20033 & w20672;
assign w20674 = ~w19997 & w41788;
assign w20675 = ~w20673 & ~w20674;
assign w20676 = ~w20670 & w20675;
assign w20677 = ~w20661 & ~w20676;
assign w20678 = w20657 & ~w20677;
assign w20679 = ~w19295 & ~w19385;
assign w20680 = w19308 & ~w19387;
assign w20681 = w19323 & ~w20651;
assign w20682 = ~w20680 & ~w20681;
assign w20683 = w19324 & ~w19387;
assign w20684 = ~w20651 & w20683;
assign w20685 = w20000 & w20679;
assign w20686 = ~w20682 & ~w20684;
assign w20687 = ~w20000 & w20686;
assign w20688 = ~w20685 & ~w20687;
assign w20689 = ~w7924 & w20688;
assign w20690 = ~w19337 & w19368;
assign w20691 = w19387 & ~w20690;
assign w20692 = ~w19387 & w20690;
assign w20693 = ~w20691 & ~w20692;
assign w20694 = w20684 & ~w20690;
assign w20695 = ~w20684 & ~w20693;
assign w20696 = ~w20694 & ~w20695;
assign w20697 = ~w20000 & ~w20696;
assign w20698 = ~w19330 & ~w19335;
assign w20699 = w20000 & w20698;
assign w20700 = ~w20697 & ~w20699;
assign w20701 = ~w7315 & w20700;
assign w20702 = ~w20689 & ~w20701;
assign w20703 = w11138 & ~w20569;
assign w20704 = ~w20000 & w20703;
assign w20705 = w11138 & w20575;
assign w20706 = ~w19999 & w20705;
assign w20707 = ~w19997 & w20706;
assign w20708 = (w10419 & w19997) | (w10419 & w41789) | (w19997 & w41789);
assign w20709 = ~w20704 & w20708;
assign w20710 = ~w20704 & ~w20707;
assign w20711 = ~w10419 & ~w20710;
assign w20712 = ~w20599 & ~w20709;
assign w20713 = ~w20711 & ~w20712;
assign w20714 = w20702 & w20713;
assign w20715 = w20678 & w20714;
assign w20716 = ~w20624 & w20715;
assign w20717 = ~w20605 & w20716;
assign w20718 = w7315 & ~w20700;
assign w20719 = w19368 & ~w19388;
assign w20720 = w20650 & ~w20719;
assign w20721 = ~w19324 & w19388;
assign w20722 = w19368 & ~w20721;
assign w20723 = ~w20266 & w20720;
assign w20724 = w20722 & ~w20723;
assign w20725 = w7315 & ~w20724;
assign w20726 = ~w7315 & w20724;
assign w20727 = ~w20725 & ~w20726;
assign w20728 = ~w20000 & ~w20727;
assign w20729 = ~w6769 & ~w19413;
assign w20730 = (w20729 & w20000) | (w20729 & w45135) | (w20000 & w45135);
assign w20731 = ~w6769 & w19413;
assign w20732 = ~w20000 & w45136;
assign w20733 = ~w20730 & ~w20732;
assign w20734 = ~w20718 & w20733;
assign w20735 = ~w20702 & w20734;
assign w20736 = w9781 & ~w20667;
assign w20737 = (w20736 & w19997) | (w20736 & w41790) | (w19997 & w41790);
assign w20738 = ~w20666 & w20737;
assign w20739 = w9781 & w20667;
assign w20740 = w20665 & w20739;
assign w20741 = ~w20033 & w20740;
assign w20742 = ~w19997 & w41791;
assign w20743 = ~w20741 & ~w20742;
assign w20744 = ~w20738 & w20743;
assign w20745 = ~w20661 & w20744;
assign w20746 = w20657 & ~w20745;
assign w20747 = w8666 & w20655;
assign w20748 = w7924 & ~w20688;
assign w20749 = ~w20747 & ~w20748;
assign w20750 = w20734 & w20749;
assign w20751 = ~w20746 & w20750;
assign w20752 = ~w20735 & ~w20751;
assign w20753 = (~w20752 & w20605) | (~w20752 & w41792) | (w20605 & w41792);
assign w20754 = ~w6264 & ~w20277;
assign w20755 = w6769 & w19413;
assign w20756 = (w20755 & w20000) | (w20755 & w45137) | (w20000 & w45137);
assign w20757 = w6769 & ~w19413;
assign w20758 = ~w20000 & w45138;
assign w20759 = ~w20756 & ~w20758;
assign w20760 = ~w20754 & w20759;
assign w20761 = (w20760 & w20380) | (w20760 & w45139) | (w20380 & w45139);
assign w20762 = w20393 & w20761;
assign w20763 = ~w20753 & w20762;
assign w20764 = w20396 & ~w20763;
assign w20765 = ~w20032 & ~w20764;
assign w20766 = (~w20226 & w20224) | (~w20226 & w41793) | (w20224 & w41793);
assign w20767 = ~w20395 & w20766;
assign w20768 = ~w20763 & w20767;
assign w20769 = ~w20017 & ~w20225;
assign w20770 = w400 & ~w20029;
assign w20771 = ~w20016 & ~w20017;
assign w20772 = ~w20030 & ~w20770;
assign w20773 = ~w20771 & ~w20772;
assign w20774 = (w20773 & ~w20768) | (w20773 & w45140) | (~w20768 & w45140);
assign w20775 = w20346 & ~w20752;
assign w20776 = (w20775 & w20605) | (w20775 & w41794) | (w20605 & w41794);
assign w20777 = w20262 & ~w20760;
assign w20778 = w20252 & w20777;
assign w20779 = w20345 & w20778;
assign w20780 = ~w20389 & ~w20779;
assign w20781 = ~w20381 & w20780;
assign w20782 = ~w20776 & w20781;
assign w20783 = (w19982 & w19732) | (w19982 & w41795) | (w19732 & w41795);
assign w20784 = w19708 & w20783;
assign w20785 = w19293 & w19982;
assign w20786 = ~w19814 & ~w19940;
assign w20787 = ~w20785 & w20786;
assign w20788 = ~w20784 & w20787;
assign w20789 = ~w19852 & ~w19920;
assign w20790 = ~w20784 & w45141;
assign w20791 = ~w19852 & ~w19972;
assign w20792 = ~w20790 & w20791;
assign w20793 = w3 & ~w20000;
assign w20794 = ~w20792 & w20793;
assign w20795 = ~w3 & ~w20000;
assign w20796 = w20792 & w20795;
assign w20797 = ~w20794 & ~w20796;
assign w20798 = w19826 & w20797;
assign w20799 = ~w19827 & w20791;
assign w20800 = ~w20790 & w20799;
assign w20801 = w3 & w19826;
assign w20802 = ~w20800 & ~w20801;
assign w20803 = ~w42 & ~w20000;
assign w20804 = w19842 & ~w20803;
assign w20805 = ~w20000 & ~w20802;
assign w20806 = w19827 & w19931;
assign w20807 = ~w20792 & w20806;
assign w20808 = w42 & ~w19826;
assign w20809 = w20000 & w20808;
assign w20810 = ~w20807 & ~w20809;
assign w20811 = ~w42 & ~w19842;
assign w20812 = ~w20802 & w20811;
assign w20813 = w20810 & ~w20812;
assign w20814 = w19843 & ~w20805;
assign w20815 = w20813 & ~w20814;
assign w20816 = ~w20802 & w20804;
assign w20817 = ~w20798 & w20816;
assign w20818 = w20815 & ~w20817;
assign w20819 = ~w20785 & w45142;
assign w20820 = (~w19970 & w20784) | (~w19970 & w45143) | (w20784 & w45143);
assign w20821 = ~w19897 & w19986;
assign w20822 = (w20821 & w19736) | (w20821 & w45144) | (w19736 & w45144);
assign w20823 = w20820 & w20822;
assign w20824 = w57 & w20000;
assign w20825 = ~w20823 & ~w20824;
assign w20826 = w19864 & w19874;
assign w20827 = w20825 & ~w20826;
assign w20828 = ~w20825 & w20826;
assign w20829 = ~w20827 & ~w20828;
assign w20830 = ~w80 & w20829;
assign w20831 = ~w19852 & ~w19855;
assign w20832 = (w19971 & w20784) | (w19971 & w45145) | (w20784 & w45145);
assign w20833 = w80 & w20000;
assign w20834 = w19864 & ~w20000;
assign w20835 = ~w20832 & w20834;
assign w20836 = (w20831 & w20835) | (w20831 & w45146) | (w20835 & w45146);
assign w20837 = ~w20835 & w45147;
assign w20838 = ~w20836 & ~w20837;
assign w20839 = w3 & ~w20838;
assign w20840 = ~w20830 & ~w20839;
assign w20841 = ~w19940 & w19968;
assign w20842 = ~w19814 & ~w20785;
assign w20843 = ~w20784 & w20842;
assign w20844 = ~w400 & w20000;
assign w20845 = ~w20000 & w20843;
assign w20846 = ~w20844 & ~w20845;
assign w20847 = w20841 & ~w20846;
assign w20848 = ~w20841 & w20846;
assign w20849 = ~w20847 & ~w20848;
assign w20850 = ~w351 & ~w20849;
assign w20851 = ~w20770 & ~w20850;
assign w20852 = ~w351 & w20000;
assign w20853 = ~w20000 & ~w20788;
assign w20854 = w19968 & w20853;
assign w20855 = ~w20852 & ~w20854;
assign w20856 = w19913 & w19963;
assign w20857 = w252 & ~w20856;
assign w20858 = (w20857 & w20854) | (w20857 & w45148) | (w20854 & w45148);
assign w20859 = w252 & w20856;
assign w20860 = ~w20854 & w45149;
assign w20861 = ~w20858 & ~w20860;
assign w20862 = w19897 & w19986;
assign w20863 = w19917 & ~w20862;
assign w20864 = (w19969 & w20784) | (w19969 & w45150) | (w20784 & w45150);
assign w20865 = w19913 & ~w20864;
assign w20866 = ~w19896 & w20000;
assign w20867 = ~w20820 & w20821;
assign w20868 = ~w20866 & ~w20867;
assign w20869 = ~w20863 & ~w20865;
assign w20870 = w20868 & ~w20869;
assign w20871 = w19896 & ~w20082;
assign w20872 = w19737 & w20871;
assign w20873 = w57 & ~w20872;
assign w20874 = ~w20870 & w20873;
assign w20875 = w20861 & ~w20874;
assign w20876 = w20851 & w20875;
assign w20877 = ~w20818 & w20840;
assign w20878 = w20876 & w20877;
assign w20879 = ~w20032 & w20878;
assign w20880 = w20121 & ~w20391;
assign w20881 = w20879 & w20880;
assign w20882 = w20782 & w20881;
assign w20883 = ~w20229 & w20879;
assign w20884 = ~w252 & w20856;
assign w20885 = (w20884 & w20854) | (w20884 & w45151) | (w20854 & w45151);
assign w20886 = ~w252 & ~w20856;
assign w20887 = ~w20854 & w45152;
assign w20888 = ~w20885 & ~w20887;
assign w20889 = w351 & w20849;
assign w20890 = w20888 & ~w20889;
assign w20891 = w20875 & ~w20890;
assign w20892 = ~w20870 & ~w20872;
assign w20893 = ~w57 & ~w20892;
assign w20894 = w80 & ~w20829;
assign w20895 = ~w20893 & ~w20894;
assign w20896 = ~w20891 & w20895;
assign w20897 = ~w19826 & ~w20797;
assign w20898 = ~w20798 & ~w20897;
assign w20899 = ~w3 & w20838;
assign w20900 = ~w42 & w20898;
assign w20901 = ~w20899 & ~w20900;
assign w20902 = w20877 & ~w20896;
assign w20903 = ~w20818 & ~w20901;
assign w20904 = ~w20902 & ~w20903;
assign w20905 = ~w20883 & w20904;
assign w20906 = ~w20882 & w20905;
assign w20907 = ~w400 & ~w20029;
assign w20908 = ~w20906 & ~w20907;
assign w20909 = ~w20908 & w45153;
assign w20910 = ~w20396 & w20879;
assign w20911 = (w20904 & w20396) | (w20904 & w45154) | (w20396 & w45154);
assign w20912 = w20762 & w20879;
assign w20913 = w20762 & w45155;
assign w20914 = w20911 & ~w20913;
assign w20915 = ~w20029 & ~w20914;
assign w20916 = w20770 & w20771;
assign w20917 = w20769 & w20770;
assign w20918 = (~w20916 & ~w20768) | (~w20916 & w45156) | (~w20768 & w45156);
assign w20919 = w351 & w20918;
assign w20920 = ~w20915 & w20919;
assign w20921 = ~w20909 & w20920;
assign w20922 = ~w20915 & w20918;
assign w20923 = ~w20909 & w20922;
assign w20924 = ~w351 & ~w20923;
assign w20925 = w20532 & w20542;
assign w20926 = (~w20621 & ~w20532) | (~w20621 & w41796) | (~w20532 & w41796);
assign w20927 = (w20618 & w20926) | (w20618 & w48960) | (w20926 & w48960);
assign w20928 = w11870 & ~w20927;
assign w20929 = ~w11870 & w20927;
assign w20930 = ~w20928 & ~w20929;
assign w20931 = (w20590 & ~w20906) | (w20590 & w45157) | (~w20906 & w45157);
assign w20932 = w20906 & w45158;
assign w20933 = ~w20931 & ~w20932;
assign w20934 = w11138 & w20933;
assign w20935 = ~w20579 & w20710;
assign w20936 = ~w20561 & w20620;
assign w20937 = ~w20591 & ~w20936;
assign w20938 = w20620 & ~w20621;
assign w20939 = (w20938 & ~w20532) | (w20938 & w41797) | (~w20532 & w41797);
assign w20940 = w20937 & ~w20939;
assign w20941 = ~w20935 & ~w20940;
assign w20942 = w20935 & w20937;
assign w20943 = ~w20939 & w20942;
assign w20944 = w20578 & ~w20906;
assign w20945 = ~w20941 & ~w20943;
assign w20946 = w20906 & w20945;
assign w20947 = ~w20944 & ~w20946;
assign w20948 = ~w10419 & ~w20947;
assign w20949 = ~w20934 & ~w20948;
assign w20950 = ~w20552 & ~w20926;
assign w20951 = w12666 & ~w20950;
assign w20952 = ~w12666 & w20950;
assign w20953 = ~w20951 & ~w20952;
assign w20954 = w20553 & ~w20613;
assign w20955 = ~w20553 & w20613;
assign w20956 = ~w20954 & ~w20955;
assign w20957 = (~w20956 & ~w20906) | (~w20956 & w45159) | (~w20906 & w45159);
assign w20958 = w20953 & w20956;
assign w20959 = w20914 & w20958;
assign w20960 = ~w20957 & ~w20959;
assign w20961 = w11870 & ~w20960;
assign w20962 = ~w11138 & ~w20933;
assign w20963 = ~w20961 & ~w20962;
assign w20964 = ~w20489 & ~w20526;
assign w20965 = w20504 & ~w20964;
assign w20966 = w20522 & ~w20965;
assign w20967 = w20542 & ~w20966;
assign w20968 = w20911 & w48961;
assign w20969 = ~w13384 & w20516;
assign w20970 = ~w20968 & w20969;
assign w20971 = ~w13384 & ~w20516;
assign w20972 = w20968 & w20971;
assign w20973 = ~w20970 & ~w20972;
assign w20974 = ~w13384 & w20925;
assign w20975 = w13384 & ~w20925;
assign w20976 = ~w20974 & ~w20975;
assign w20977 = (w20551 & ~w20906) | (w20551 & w45160) | (~w20906 & w45160);
assign w20978 = ~w20551 & ~w20976;
assign w20979 = w20911 & w48962;
assign w20980 = ~w20977 & ~w20979;
assign w20981 = ~w20977 & w48963;
assign w20982 = w20973 & ~w20981;
assign w20983 = w13384 & ~w20516;
assign w20984 = ~w20968 & w20983;
assign w20985 = w13384 & w20516;
assign w20986 = w20968 & w20985;
assign w20987 = ~w20984 & ~w20986;
assign w20988 = ~w14766 & w20964;
assign w20989 = w14766 & ~w20964;
assign w20990 = ~w20988 & ~w20989;
assign w20991 = w20498 & ~w20499;
assign w20992 = ~w20498 & w20499;
assign w20993 = ~w20991 & ~w20992;
assign w20994 = (w20993 & ~w20906) | (w20993 & w45161) | (~w20906 & w45161);
assign w20995 = ~w20990 & ~w20993;
assign w20996 = w20911 & w48964;
assign w20997 = ~w20994 & ~w20996;
assign w20998 = ~w20994 & w48965;
assign w20999 = w20987 & w20998;
assign w21000 = w20982 & ~w20999;
assign w21001 = ~w11870 & w20960;
assign w21002 = (~w12666 & w20977) | (~w12666 & w48966) | (w20977 & w48966);
assign w21003 = ~w21001 & ~w21002;
assign w21004 = w20949 & w21003;
assign w21005 = w20949 & ~w20963;
assign w21006 = ~w21000 & w21004;
assign w21007 = ~w21005 & ~w21006;
assign w21008 = ~a[36] & ~w20000;
assign w21009 = ~w19040 & ~w20000;
assign w21010 = w19040 & w20000;
assign w21011 = ~w21009 & ~w21010;
assign w21012 = ~w20410 & w21011;
assign w21013 = (w21012 & w20906) | (w21012 & w45162) | (w20906 & w45162);
assign w21014 = ~w20414 & ~w20913;
assign w21015 = w20911 & w21014;
assign w21016 = w20410 & w21010;
assign w21017 = ~w20913 & w21016;
assign w21018 = w20911 & w21017;
assign w21019 = a[37] & ~w21018;
assign w21020 = w21008 & ~w21015;
assign w21021 = w21019 & ~w21020;
assign w21022 = ~w21013 & w21021;
assign w21023 = ~w20000 & ~w20429;
assign w21024 = w21015 & w21023;
assign w21025 = ~w21008 & ~w21016;
assign w21026 = ~w21012 & w21025;
assign w21027 = ~a[37] & ~w21026;
assign w21028 = (w21027 & w20906) | (w21027 & w45163) | (w20906 & w45163);
assign w21029 = ~w21024 & w21028;
assign w21030 = ~w18183 & ~w21029;
assign w21031 = ~w21022 & w21030;
assign w21032 = a[36] & w20000;
assign w21033 = a[36] & ~w20409;
assign w21034 = ~w20410 & ~w21033;
assign w21035 = ~w21008 & ~w21032;
assign w21036 = ~w20906 & w21035;
assign w21037 = w20906 & w21034;
assign w21038 = ~w21036 & ~w21037;
assign w21039 = ~a[32] & ~a[33];
assign w21040 = ~a[34] & w21039;
assign w21041 = w20000 & ~w21040;
assign w21042 = ~a[35] & ~w21041;
assign w21043 = ~w20914 & w21042;
assign w21044 = a[34] & ~a[35];
assign w21045 = ~w20913 & w21044;
assign w21046 = w20911 & w21045;
assign w21047 = ~w20000 & w21040;
assign w21048 = a[35] & ~w21041;
assign w21049 = ~w20902 & w45164;
assign w21050 = ~w20883 & w21049;
assign w21051 = ~w20882 & w21050;
assign w21052 = ~w21047 & ~w21051;
assign w21053 = ~w21046 & w21052;
assign w21054 = ~w21043 & w21053;
assign w21055 = w19040 & w21038;
assign w21056 = ~w21054 & ~w21055;
assign w21057 = ~w19040 & ~w21038;
assign w21058 = ~w21056 & ~w21057;
assign w21059 = ~w21031 & w21058;
assign w21060 = w18183 & w21029;
assign w21061 = w18183 & ~w21013;
assign w21062 = w21021 & w21061;
assign w21063 = ~w21060 & ~w21062;
assign w21064 = ~w19462 & ~w20000;
assign w21065 = ~w21010 & ~w21064;
assign w21066 = a[38] & ~w21065;
assign w21067 = ~a[38] & w21065;
assign w21068 = ~w21066 & ~w21067;
assign w21069 = ~a[37] & ~w20000;
assign w21070 = w20429 & ~w21069;
assign w21071 = ~a[37] & w20000;
assign w21072 = ~w21064 & ~w21071;
assign w21073 = ~w20415 & w21072;
assign w21074 = ~w21070 & ~w21073;
assign w21075 = w18183 & w21074;
assign w21076 = ~w18183 & ~w20415;
assign w21077 = ~w21074 & w21076;
assign w21078 = ~w21075 & ~w21077;
assign w21079 = w20914 & ~w21078;
assign w21080 = w20906 & ~w21078;
assign w21081 = w21068 & ~w21080;
assign w21082 = ~w17380 & ~w21081;
assign w21083 = ~w21068 & w21079;
assign w21084 = w21082 & ~w21083;
assign w21085 = w21063 & ~w21084;
assign w21086 = ~w21059 & w21085;
assign w21087 = ~w20441 & w20468;
assign w21088 = ~w16559 & w21087;
assign w21089 = w16559 & ~w21087;
assign w21090 = ~w21088 & ~w21089;
assign w21091 = w20911 & w48967;
assign w21092 = w20444 & ~w20459;
assign w21093 = ~w20444 & w20459;
assign w21094 = ~w21090 & w21093;
assign w21095 = w20906 & w21094;
assign w21096 = ~w21090 & w21092;
assign w21097 = w20911 & w48968;
assign w21098 = ~w21095 & ~w21097;
assign w21099 = ~w21092 & ~w21093;
assign w21100 = ~w21091 & w21099;
assign w21101 = w21098 & ~w21100;
assign w21102 = ~w20470 & w20475;
assign w21103 = ~w15681 & w21102;
assign w21104 = w15681 & ~w21102;
assign w21105 = ~w21103 & ~w21104;
assign w21106 = w14766 & ~w20525;
assign w21107 = (w21106 & ~w20906) | (w21106 & w45165) | (~w20906 & w45165);
assign w21108 = w14766 & w20525;
assign w21109 = w20906 & w45166;
assign w21110 = ~w21107 & ~w21109;
assign w21111 = ~w15681 & w21110;
assign w21112 = w21101 & w21111;
assign w21113 = (w20525 & ~w20906) | (w20525 & w48969) | (~w20906 & w48969);
assign w21114 = w20906 & w48970;
assign w21115 = ~w21113 & ~w21114;
assign w21116 = ~w14766 & ~w21115;
assign w21117 = ~w21112 & ~w21116;
assign w21118 = w21068 & ~w21079;
assign w21119 = ~w21068 & w21080;
assign w21120 = ~w21118 & ~w21119;
assign w21121 = w17380 & ~w21120;
assign w21122 = w20440 & w20468;
assign w21123 = (w20407 & ~w20906) | (w20407 & w45167) | (~w20906 & w45167);
assign w21124 = w20906 & w45168;
assign w21125 = ~w21123 & ~w21124;
assign w21126 = ~w16559 & w21125;
assign w21127 = ~w21121 & ~w21126;
assign w21128 = w21117 & w21127;
assign w21129 = ~w21086 & w21128;
assign w21130 = (w15681 & ~w21098) | (w15681 & w48971) | (~w21098 & w48971);
assign w21131 = w16559 & ~w21125;
assign w21132 = w21110 & ~w21131;
assign w21133 = ~w21130 & w21132;
assign w21134 = w21117 & ~w21133;
assign w21135 = (~w14039 & w20994) | (~w14039 & w48972) | (w20994 & w48972);
assign w21136 = w20987 & ~w21135;
assign w21137 = w20982 & ~w21136;
assign w21138 = w21004 & ~w21137;
assign w21139 = ~w21134 & w21138;
assign w21140 = ~w21129 & w21139;
assign w21141 = (w21007 & w21129) | (w21007 & w45169) | (w21129 & w45169);
assign w21142 = ~w20746 & ~w20747;
assign w21143 = ~w20624 & w20713;
assign w21144 = ~w20605 & w21143;
assign w21145 = ~w20605 & w41798;
assign w21146 = w21142 & ~w21145;
assign w21147 = ~w20689 & ~w21146;
assign w21148 = ~w20748 & ~w21147;
assign w21149 = w20718 & w20906;
assign w21150 = ~w20701 & ~w21149;
assign w21151 = w7315 & ~w21148;
assign w21152 = w20906 & ~w21151;
assign w21153 = ~w7315 & ~w20700;
assign w21154 = ~w21148 & w21153;
assign w21155 = w20914 & w21154;
assign w21156 = w20700 & ~w21152;
assign w21157 = ~w21155 & ~w21156;
assign w21158 = w21148 & ~w21150;
assign w21159 = w21157 & ~w21158;
assign w21160 = w6769 & ~w21159;
assign w21161 = w7924 & ~w21146;
assign w21162 = ~w7924 & w21146;
assign w21163 = ~w21161 & ~w21162;
assign w21164 = w20914 & w21163;
assign w21165 = ~w20688 & ~w21164;
assign w21166 = w20906 & w21163;
assign w21167 = w20688 & w21166;
assign w21168 = ~w21165 & ~w21167;
assign w21169 = ~w7315 & w21168;
assign w21170 = ~w21160 & ~w21169;
assign w21171 = w20676 & w20744;
assign w21172 = w21144 & ~w21171;
assign w21173 = ~w21144 & w21171;
assign w21174 = ~w21172 & ~w21173;
assign w21175 = ~w9781 & w20676;
assign w21176 = w20744 & ~w21175;
assign w21177 = ~w9195 & ~w21174;
assign w21178 = w20906 & w21177;
assign w21179 = ~w9195 & ~w21176;
assign w21180 = ~w20906 & w21179;
assign w21181 = ~w21178 & ~w21180;
assign w21182 = ~w20605 & w41799;
assign w21183 = w20744 & ~w21182;
assign w21184 = ~w9195 & w21183;
assign w21185 = ~w20636 & ~w20659;
assign w21186 = w9195 & ~w21183;
assign w21187 = (w21185 & ~w20906) | (w21185 & w45170) | (~w20906 & w45170);
assign w21188 = w20914 & w21184;
assign w21189 = w21187 & ~w21188;
assign w21190 = ~w21184 & ~w21186;
assign w21191 = w20906 & w45171;
assign w21192 = ~w8666 & w21181;
assign w21193 = w21181 & ~w21191;
assign w21194 = ~w21189 & w21193;
assign w21195 = ~w21192 & ~w21194;
assign w21196 = ~w8666 & ~w21191;
assign w21197 = ~w21189 & w21196;
assign w21198 = w20745 & ~w21182;
assign w21199 = ~w8666 & w20643;
assign w21200 = ~w21198 & w21199;
assign w21201 = w8666 & ~w20643;
assign w21202 = w8666 & w20745;
assign w21203 = ~w21182 & w21202;
assign w21204 = ~w21201 & ~w21203;
assign w21205 = (w20655 & ~w20906) | (w20655 & w45172) | (~w20906 & w45172);
assign w21206 = w20914 & w21200;
assign w21207 = w21205 & ~w21206;
assign w21208 = ~w21200 & w21204;
assign w21209 = w20906 & w45173;
assign w21210 = ~w7924 & ~w21209;
assign w21211 = ~w21207 & w21210;
assign w21212 = ~w21197 & ~w21211;
assign w21213 = w21195 & w21212;
assign w21214 = ~w21207 & ~w21209;
assign w21215 = w7924 & ~w21214;
assign w21216 = w7315 & ~w21168;
assign w21217 = ~w21215 & ~w21216;
assign w21218 = ~w21213 & w21217;
assign w21219 = w20906 & w21174;
assign w21220 = ~w20906 & w21176;
assign w21221 = ~w21219 & ~w21220;
assign w21222 = ~w20709 & ~w20711;
assign w21223 = w10419 & w20943;
assign w21224 = ~w20943 & w21222;
assign w21225 = ~w21223 & ~w21224;
assign w21226 = (w20599 & ~w20906) | (w20599 & w45174) | (~w20906 & w45174);
assign w21227 = ~w20599 & w21222;
assign w21228 = ~w20943 & w21227;
assign w21229 = w10419 & ~w20599;
assign w21230 = w20943 & w21229;
assign w21231 = ~w21228 & ~w21230;
assign w21232 = ~w20913 & ~w21231;
assign w21233 = w20911 & w21232;
assign w21234 = ~w9781 & ~w21233;
assign w21235 = ~w21226 & w21234;
assign w21236 = w9195 & ~w21221;
assign w21237 = ~w21235 & ~w21236;
assign w21238 = w21212 & w21237;
assign w21239 = ~w21213 & w48973;
assign w21240 = w21170 & ~w21239;
assign w21241 = ~w21141 & w21240;
assign w21242 = ~w6769 & w21159;
assign w21243 = w10419 & w20947;
assign w21244 = w9781 & w20599;
assign w21245 = (w21244 & ~w20906) | (w21244 & w45175) | (~w20906 & w45175);
assign w21246 = w9781 & w21233;
assign w21247 = ~w21245 & ~w21246;
assign w21248 = ~w21243 & w21247;
assign w21249 = w21237 & ~w21248;
assign w21250 = w21212 & w21249;
assign w21251 = ~w21170 & ~w21242;
assign w21252 = ~w21242 & ~w21250;
assign w21253 = w21218 & w21252;
assign w21254 = ~w21251 & ~w21253;
assign w21255 = ~w20624 & w41800;
assign w21256 = ~w20605 & w21255;
assign w21257 = ~w20288 & ~w20347;
assign w21258 = ~w20735 & w20760;
assign w21259 = ~w20751 & w21258;
assign w21260 = ~w20278 & w21257;
assign w21261 = ~w21259 & w21260;
assign w21262 = (w21261 & w20605) | (w21261 & w41801) | (w20605 & w41801);
assign w21263 = ~w5745 & ~w20904;
assign w21264 = w21262 & ~w21263;
assign w21265 = ~w20396 & w45176;
assign w21266 = w21264 & ~w21265;
assign w21267 = ~w20278 & ~w21259;
assign w21268 = ~w21256 & w21267;
assign w21269 = ~w21257 & ~w21268;
assign w21270 = w20906 & w21269;
assign w21271 = ~w21266 & ~w21270;
assign w21272 = w20287 & ~w20906;
assign w21273 = (w5330 & ~w21271) | (w5330 & w45177) | (~w21271 & w45177);
assign w21274 = ~w20278 & ~w20754;
assign w21275 = ~w20753 & w20759;
assign w21276 = ~w21274 & w21275;
assign w21277 = (w20277 & ~w20906) | (w20277 & w45178) | (~w20906 & w45178);
assign w21278 = w21274 & ~w21275;
assign w21279 = w20906 & w21278;
assign w21280 = ~w20912 & w21276;
assign w21281 = w20911 & w21280;
assign w21282 = ~w21279 & ~w21281;
assign w21283 = ~w21277 & w21282;
assign w21284 = (~w5745 & ~w21282) | (~w5745 & w45179) | (~w21282 & w45179);
assign w21285 = ~w20748 & w21142;
assign w21286 = w20702 & ~w21285;
assign w21287 = ~w20718 & ~w21286;
assign w21288 = ~w20717 & w21287;
assign w21289 = ~w6769 & w21288;
assign w21290 = w6769 & ~w21288;
assign w21291 = ~w21289 & ~w21290;
assign w21292 = w19413 & ~w20728;
assign w21293 = ~w19413 & w20728;
assign w21294 = ~w21292 & ~w21293;
assign w21295 = (~w21294 & ~w20906) | (~w21294 & w45180) | (~w20906 & w45180);
assign w21296 = ~w21291 & w21294;
assign w21297 = w20914 & w21296;
assign w21298 = ~w21295 & ~w21297;
assign w21299 = ~w6264 & ~w21298;
assign w21300 = w21271 & w45181;
assign w21301 = w5745 & w21283;
assign w21302 = ~w21300 & ~w21301;
assign w21303 = ~w21284 & w21299;
assign w21304 = (~w21273 & ~w21302) | (~w21273 & w45182) | (~w21302 & w45182);
assign w21305 = ~w20347 & ~w21262;
assign w21306 = w5330 & ~w21305;
assign w21307 = ~w5330 & w21305;
assign w21308 = ~w21306 & ~w21307;
assign w21309 = w20333 & ~w20348;
assign w21310 = ~w20333 & w20348;
assign w21311 = ~w21309 & ~w21310;
assign w21312 = (~w21311 & ~w20906) | (~w21311 & w45183) | (~w20906 & w45183);
assign w21313 = ~w21308 & w21311;
assign w21314 = w20914 & w21313;
assign w21315 = ~w21312 & ~w21314;
assign w21316 = w4838 & w21315;
assign w21317 = ~w20314 & ~w20316;
assign w21318 = w20317 & ~w21317;
assign w21319 = ~w20317 & w21317;
assign w21320 = ~w21318 & ~w21319;
assign w21321 = w20289 & w20342;
assign w21322 = ~w21259 & w21321;
assign w21323 = w20342 & ~w20354;
assign w21324 = ~w20326 & w21323;
assign w21325 = (~w21324 & w21256) | (~w21324 & w41802) | (w21256 & w41802);
assign w21326 = ~w21256 & w21322;
assign w21327 = ~w21323 & ~w21326;
assign w21328 = ~w4838 & w21320;
assign w21329 = ~w21327 & w21328;
assign w21330 = w20914 & w21329;
assign w21331 = (~w21320 & ~w20906) | (~w21320 & w45184) | (~w20906 & w45184);
assign w21332 = ~w21330 & ~w21331;
assign w21333 = w20326 & w21327;
assign w21334 = ~w20369 & w21327;
assign w21335 = (~w21333 & ~w20906) | (~w21333 & w45185) | (~w20906 & w45185);
assign w21336 = ~w4430 & w21335;
assign w21337 = w21332 & w21336;
assign w21338 = ~w21316 & ~w21337;
assign w21339 = w6264 & w21298;
assign w21340 = ~w21273 & ~w21284;
assign w21341 = ~w21339 & w21340;
assign w21342 = w21338 & ~w21341;
assign w21343 = ~w21304 & w21342;
assign w21344 = w20300 & w20360;
assign w21345 = w4430 & ~w20906;
assign w21346 = w20906 & w45186;
assign w21347 = ~w21345 & ~w21346;
assign w21348 = w21344 & ~w21347;
assign w21349 = ~w21344 & w21347;
assign w21350 = ~w21348 & ~w21349;
assign w21351 = w4056 & w21350;
assign w21352 = w21332 & w21335;
assign w21353 = w4430 & ~w21352;
assign w21354 = ~w4838 & ~w21315;
assign w21355 = ~w21337 & w21354;
assign w21356 = ~w21353 & ~w21355;
assign w21357 = ~w21351 & w21356;
assign w21358 = ~w21343 & w21357;
assign w21359 = ~w21254 & w21358;
assign w21360 = w20057 & ~w20217;
assign w21361 = ~w20212 & w41803;
assign w21362 = w41803 & w45187;
assign w21363 = w20390 & w20781;
assign w21364 = ~w20776 & w21363;
assign w21365 = w21362 & ~w21364;
assign w21366 = w20080 & ~w20104;
assign w21367 = w20057 & w21366;
assign w21368 = (w21367 & w21364) | (w21367 & w45188) | (w21364 & w45188);
assign w21369 = w20906 & ~w21368;
assign w21370 = (w20107 & w21364) | (w20107 & w45189) | (w21364 & w45189);
assign w21371 = ~w945 & w21366;
assign w21372 = ~w21370 & ~w21371;
assign w21373 = ~w20068 & ~w20069;
assign w21374 = w20070 & ~w21373;
assign w21375 = ~w20070 & w21373;
assign w21376 = ~w21374 & ~w21375;
assign w21377 = ~w20906 & w21376;
assign w21378 = w21369 & ~w21372;
assign w21379 = ~w20906 & w45190;
assign w21380 = ~w21378 & ~w21379;
assign w21381 = ~w20099 & ~w20110;
assign w21382 = ~w20081 & ~w20104;
assign w21383 = ~w20391 & ~w21382;
assign w21384 = ~w20776 & w45191;
assign w21385 = w20081 & ~w21362;
assign w21386 = ~w20104 & ~w21385;
assign w21387 = ~w21384 & w21386;
assign w21388 = w21381 & ~w21387;
assign w21389 = ~w21381 & w21386;
assign w21390 = ~w21384 & w21389;
assign w21391 = (~w754 & w20906) | (~w754 & w45192) | (w20906 & w45192);
assign w21392 = w20906 & ~w21390;
assign w21393 = ~w21388 & w21392;
assign w21394 = w21391 & ~w21393;
assign w21395 = ~w21380 & ~w21394;
assign w21396 = w612 & ~w20117;
assign w21397 = ~w20106 & ~w20110;
assign w21398 = ~w20224 & w21397;
assign w21399 = w20390 & w21397;
assign w21400 = w20781 & w21399;
assign w21401 = ~w20776 & w21400;
assign w21402 = ~w21398 & ~w21401;
assign w21403 = ~w20118 & ~w20226;
assign w21404 = w612 & ~w21403;
assign w21405 = (w21404 & w21401) | (w21404 & w45193) | (w21401 & w45193);
assign w21406 = w612 & w21403;
assign w21407 = ~w21398 & w21406;
assign w21408 = ~w21401 & w21407;
assign w21409 = ~w20906 & ~w21396;
assign w21410 = w20906 & w45194;
assign w21411 = ~w21409 & ~w21410;
assign w21412 = ~w20902 & w45195;
assign w21413 = ~w20883 & w21412;
assign w21414 = ~w20882 & w21413;
assign w21415 = ~w21390 & w21414;
assign w21416 = ~w21388 & w21415;
assign w21417 = w754 & ~w20906;
assign w21418 = ~w20906 & w45196;
assign w21419 = ~w21416 & ~w21418;
assign w21420 = w20906 & ~w21402;
assign w21421 = ~w21417 & ~w21420;
assign w21422 = w21403 & ~w21421;
assign w21423 = ~w21403 & w21421;
assign w21424 = ~w21422 & ~w21423;
assign w21425 = ~w612 & ~w21424;
assign w21426 = ~w21411 & w21419;
assign w21427 = ~w21395 & w21426;
assign w21428 = ~w21425 & ~w21427;
assign w21429 = w21361 & ~w21364;
assign w21430 = ~w21360 & ~w21429;
assign w21431 = w20216 & ~w20906;
assign w21432 = w20906 & ~w21430;
assign w21433 = ~w21365 & w21432;
assign w21434 = ~w21431 & ~w21433;
assign w21435 = ~w1120 & w21434;
assign w21436 = ~w20902 & w45197;
assign w21437 = ~w20883 & w21436;
assign w21438 = ~w20882 & w21437;
assign w21439 = w20210 & w20775;
assign w21440 = ~w20717 & w21439;
assign w21441 = ~w20135 & ~w20168;
assign w21442 = ~w20135 & w20207;
assign w21443 = ~w21440 & w41804;
assign w21444 = ~w21441 & ~w21443;
assign w21445 = w21438 & w21444;
assign w21446 = ~w1541 & ~w20906;
assign w21447 = ~w21445 & ~w21446;
assign w21448 = w20149 & ~w20221;
assign w21449 = (w1320 & w21447) | (w1320 & w45198) | (w21447 & w45198);
assign w21450 = w21447 & w21448;
assign w21451 = w21449 & ~w21450;
assign w21452 = ~w21435 & ~w21451;
assign w21453 = ~w21428 & w21452;
assign w21454 = w20134 & ~w21438;
assign w21455 = ~w21445 & ~w21454;
assign w21456 = w20151 & ~w20913;
assign w21457 = w20911 & w21456;
assign w21458 = ~w20135 & ~w21457;
assign w21459 = ~w21440 & w41805;
assign w21460 = w20206 & w21459;
assign w21461 = w20168 & ~w21460;
assign w21462 = ~w1541 & w21455;
assign w21463 = ~w1541 & w21461;
assign w21464 = ~w21458 & w21463;
assign w21465 = ~w21462 & ~w21464;
assign w21466 = ~w1320 & ~w21448;
assign w21467 = ~w21447 & w21466;
assign w21468 = ~w1320 & w21448;
assign w21469 = w21447 & w21468;
assign w21470 = ~w21467 & ~w21469;
assign w21471 = w21465 & w21470;
assign w21472 = w20168 & w20206;
assign w21473 = w20201 & ~w21472;
assign w21474 = ~w21440 & w41806;
assign w21475 = w20162 & ~w20163;
assign w21476 = ~w20162 & w20163;
assign w21477 = ~w21475 & ~w21476;
assign w21478 = w2006 & w21474;
assign w21479 = (~w21478 & w20906) | (~w21478 & w45199) | (w20906 & w45199);
assign w21480 = ~w21459 & w21472;
assign w21481 = w20906 & w21480;
assign w21482 = ~w20913 & w21474;
assign w21483 = w20911 & w21482;
assign w21484 = ~w21481 & ~w21483;
assign w21485 = (w1738 & ~w21484) | (w1738 & w45200) | (~w21484 & w45200);
assign w21486 = w1541 & ~w21455;
assign w21487 = ~w21458 & w21461;
assign w21488 = w21486 & ~w21487;
assign w21489 = ~w21485 & ~w21488;
assign w21490 = w21471 & ~w21489;
assign w21491 = w20251 & ~w20380;
assign w21492 = w20251 & w20345;
assign w21493 = w20380 & ~w21259;
assign w21494 = w21492 & w21493;
assign w21495 = ~w21256 & w21494;
assign w21496 = ~w20262 & ~w20385;
assign w21497 = (~w20385 & w20380) | (~w20385 & w45201) | (w20380 & w45201);
assign w21498 = ~w21496 & w52248;
assign w21499 = ~w20387 & w21498;
assign w21500 = w20262 & w52249;
assign w21501 = w20388 & ~w21500;
assign w21502 = w20906 & ~w21501;
assign w21503 = w20240 & ~w20906;
assign w21504 = ~w20906 & w45202;
assign w21505 = ~w2558 & ~w21499;
assign w21506 = w21502 & w21505;
assign w21507 = ~w21504 & ~w21506;
assign w21508 = ~w20371 & ~w20372;
assign w21509 = ~w20355 & w21508;
assign w21510 = ~w20345 & w21509;
assign w21511 = w20760 & w21509;
assign w21512 = ~w20753 & w21511;
assign w21513 = ~w21510 & ~w21512;
assign w21514 = w20251 & w20377;
assign w21515 = ~w3242 & w21514;
assign w21516 = w3646 & w21515;
assign w21517 = ~w20906 & w21516;
assign w21518 = w21513 & w21515;
assign w21519 = w20906 & w21518;
assign w21520 = ~w21517 & ~w21519;
assign w21521 = ~w3242 & ~w21514;
assign w21522 = ~w21513 & w21521;
assign w21523 = w20906 & w21522;
assign w21524 = ~w3646 & w21521;
assign w21525 = ~w20906 & w21524;
assign w21526 = ~w21523 & ~w21525;
assign w21527 = w21520 & w21526;
assign w21528 = w21507 & w21527;
assign w21529 = ~w20902 & w45203;
assign w21530 = ~w20883 & w21529;
assign w21531 = ~w20882 & w21530;
assign w21532 = w20906 & ~w21459;
assign w21533 = w20185 & ~w21531;
assign w21534 = ~w21532 & ~w21533;
assign w21535 = ~w20199 & w20781;
assign w21536 = ~w20776 & w21535;
assign w21537 = w20188 & ~w20209;
assign w21538 = ~w21536 & w21537;
assign w21539 = ~w20913 & w21538;
assign w21540 = w20911 & w21539;
assign w21541 = w20186 & ~w20209;
assign w21542 = ~w21536 & w21541;
assign w21543 = w2006 & ~w21542;
assign w21544 = ~w21540 & w21543;
assign w21545 = ~w21534 & w21544;
assign w21546 = (w20208 & ~w20906) | (w20208 & w45204) | (~w20906 & w45204);
assign w21547 = w2558 & w21536;
assign w21548 = ~w20913 & w21547;
assign w21549 = w20911 & w21548;
assign w21550 = ~w20902 & w45205;
assign w21551 = ~w20883 & w21550;
assign w21552 = w2285 & w20782;
assign w21553 = w2285 & ~w20199;
assign w21554 = (w21553 & w20883) | (w21553 & w45206) | (w20883 & w45206);
assign w21555 = ~w21552 & ~w21554;
assign w21556 = ~w21549 & ~w21555;
assign w21557 = ~w21546 & w21556;
assign w21558 = ~w21545 & ~w21557;
assign w21559 = ~w3242 & w21491;
assign w21560 = w3242 & ~w21491;
assign w21561 = ~w21559 & ~w21560;
assign w21562 = w21495 & ~w21561;
assign w21563 = ~w21495 & w21561;
assign w21564 = ~w21562 & ~w21563;
assign w21565 = ~w20913 & w21564;
assign w21566 = w2896 & ~w20384;
assign w21567 = (w21566 & ~w21565) | (w21566 & w41809) | (~w21565 & w41809);
assign w21568 = w2896 & w20384;
assign w21569 = w21565 & w41810;
assign w21570 = ~w21567 & ~w21569;
assign w21571 = w20300 & w20370;
assign w21572 = w21325 & w21571;
assign w21573 = ~w20309 & ~w20372;
assign w21574 = ~w20300 & w21573;
assign w21575 = w21572 & w21573;
assign w21576 = w20300 & ~w21573;
assign w21577 = ~w21572 & w21576;
assign w21578 = ~w21575 & ~w21577;
assign w21579 = ~w21574 & w21578;
assign w21580 = w20308 & ~w20906;
assign w21581 = ~w3646 & w20906;
assign w21582 = w21579 & w21581;
assign w21583 = ~w3646 & w21580;
assign w21584 = ~w21582 & ~w21583;
assign w21585 = w21570 & w21584;
assign w21586 = w21528 & w21558;
assign w21587 = w21585 & w21586;
assign w21588 = ~w21490 & w21587;
assign w21589 = w20057 & ~w21365;
assign w21590 = ~w21366 & ~w21589;
assign w21591 = w21369 & ~w21590;
assign w21592 = w945 & ~w21377;
assign w21593 = ~w21591 & w21592;
assign w21594 = ~w21394 & ~w21593;
assign w21595 = ~w21425 & w21594;
assign w21596 = ~w21428 & ~w21595;
assign w21597 = w21453 & w21588;
assign w21598 = ~w21596 & ~w21597;
assign w21599 = (~w20830 & w20891) | (~w20830 & w45207) | (w20891 & w45207);
assign w21600 = ~w3 & w21599;
assign w21601 = w3 & ~w21599;
assign w21602 = ~w21600 & ~w21601;
assign w21603 = ~w20838 & ~w21602;
assign w21604 = w20838 & w20904;
assign w21605 = w21602 & w21604;
assign w21606 = ~w21603 & ~w21605;
assign w21607 = ~w20902 & w45208;
assign w21608 = ~w20830 & w20876;
assign w21609 = ~w3 & w21608;
assign w21610 = w21607 & ~w21609;
assign w21611 = w20838 & ~w21610;
assign w21612 = ~w20032 & w20851;
assign w21613 = w20875 & w21612;
assign w21614 = w20840 & w21613;
assign w21615 = w20838 & w21602;
assign w21616 = (~w21615 & w20764) | (~w21615 & w45209) | (w20764 & w45209);
assign w21617 = ~w21602 & ~w21608;
assign w21618 = w20904 & ~w21617;
assign w21619 = ~w20838 & ~w21618;
assign w21620 = w21616 & ~w21619;
assign w21621 = ~w20765 & ~w21606;
assign w21622 = ~w21611 & ~w21620;
assign w21623 = ~w21621 & ~w21622;
assign w21624 = ~w42 & w21623;
assign w21625 = (~w20891 & w20764) | (~w20891 & w45210) | (w20764 & w45210);
assign w21626 = ~w20893 & w20906;
assign w21627 = w21625 & w21626;
assign w21628 = ~w80 & ~w20906;
assign w21629 = ~w21627 & ~w21628;
assign w21630 = ~w20830 & ~w20894;
assign w21631 = ~w3 & w21630;
assign w21632 = (w21631 & w21627) | (w21631 & w45211) | (w21627 & w45211);
assign w21633 = ~w3 & ~w21630;
assign w21634 = ~w21627 & w45212;
assign w21635 = ~w21632 & ~w21634;
assign w21636 = ~w21624 & w21635;
assign w21637 = ~w20764 & w21612;
assign w21638 = w20861 & w20888;
assign w21639 = ~w20889 & w21638;
assign w21640 = (w21639 & w20764) | (w21639 & w45213) | (w20764 & w45213);
assign w21641 = ~w252 & ~w20914;
assign w21642 = w21640 & ~w21641;
assign w21643 = (~w20889 & w20764) | (~w20889 & w45214) | (w20764 & w45214);
assign w21644 = w20855 & ~w20856;
assign w21645 = ~w20855 & w20856;
assign w21646 = ~w21644 & ~w21645;
assign w21647 = ~w20906 & ~w21646;
assign w21648 = w20906 & ~w21638;
assign w21649 = ~w21643 & w21648;
assign w21650 = ~w21647 & ~w21649;
assign w21651 = (~w57 & ~w21650) | (~w57 & w45215) | (~w21650 & w45215);
assign w21652 = ~w20874 & ~w20893;
assign w21653 = (w21652 & w20906) | (w21652 & w45216) | (w20906 & w45216);
assign w21654 = w20861 & w20906;
assign w21655 = ~w21640 & w21654;
assign w21656 = w21653 & ~w21655;
assign w21657 = w20861 & ~w21652;
assign w21658 = w20893 & ~w20906;
assign w21659 = w20906 & w21657;
assign w21660 = ~w21640 & w21659;
assign w21661 = ~w21658 & ~w21660;
assign w21662 = ~w21656 & w21661;
assign w21663 = w80 & ~w21662;
assign w21664 = w20889 & ~w20913;
assign w21665 = w20911 & w21664;
assign w21666 = ~w20850 & ~w21665;
assign w21667 = ~w20764 & w45217;
assign w21668 = ~w351 & ~w21607;
assign w21669 = ~w20889 & ~w21668;
assign w21670 = ~w20849 & ~w20906;
assign w21671 = w21637 & w21669;
assign w21672 = ~w21670 & ~w21671;
assign w21673 = ~w252 & w21672;
assign w21674 = ~w21666 & ~w21667;
assign w21675 = w21673 & ~w21674;
assign w21676 = ~w21663 & w45218;
assign w21677 = ~w20015 & ~w20225;
assign w21678 = ~w20768 & w21677;
assign w21679 = ~w19995 & ~w20017;
assign w21680 = w20906 & ~w21679;
assign w21681 = (~w20225 & w20768) | (~w20225 & w45219) | (w20768 & w45219);
assign w21682 = w21680 & ~w21681;
assign w21683 = ~w19995 & w20769;
assign w21684 = ~w20902 & w45220;
assign w21685 = ~w20883 & w21684;
assign w21686 = ~w20882 & w21685;
assign w21687 = ~w21678 & w21686;
assign w21688 = w19994 & ~w20906;
assign w21689 = ~w21687 & ~w21688;
assign w21690 = ~w21682 & w21689;
assign w21691 = w400 & w21690;
assign w21692 = w20768 & ~w21677;
assign w21693 = ~w20014 & ~w20906;
assign w21694 = w20906 & ~w21678;
assign w21695 = ~w21692 & w21694;
assign w21696 = ~w21693 & ~w21695;
assign w21697 = ~w21695 & w45221;
assign w21698 = ~w21691 & ~w21697;
assign w21699 = ~w400 & ~w21690;
assign w21700 = ~w20921 & ~w21699;
assign w21701 = ~w21698 & w21700;
assign w21702 = w493 & ~w21696;
assign w21703 = w21700 & ~w21702;
assign w21704 = ~w21701 & ~w21703;
assign w21705 = w21676 & ~w21704;
assign w21706 = ~w21704 & w45222;
assign w21707 = ~w21598 & w21706;
assign w21708 = w21359 & w21707;
assign w21709 = ~w21241 & w21708;
assign w21710 = w3 & w21630;
assign w21711 = (w21710 & w20906) | (w21710 & w45223) | (w20906 & w45223);
assign w21712 = ~w21627 & w21711;
assign w21713 = w3 & ~w21630;
assign w21714 = ~w20893 & w21713;
assign w21715 = w20906 & w21714;
assign w21716 = w21625 & w21715;
assign w21717 = ~w20906 & w45224;
assign w21718 = ~w21716 & ~w21717;
assign w21719 = ~w21712 & w21718;
assign w21720 = w252 & ~w21672;
assign w21721 = w252 & ~w21667;
assign w21722 = ~w21666 & w21721;
assign w21723 = ~w21720 & ~w21722;
assign w21724 = w21719 & w21723;
assign w21725 = ~w20924 & w21724;
assign w21726 = ~w21701 & w21725;
assign w21727 = ~w21600 & w21616;
assign w21728 = w42 & ~w20898;
assign w21729 = ~w20900 & ~w21728;
assign w21730 = ~w20818 & w20898;
assign w21731 = ~w21727 & ~w21729;
assign w21732 = w21727 & w21729;
assign w21733 = ~w21731 & ~w21732;
assign w21734 = ~w21730 & w21733;
assign w21735 = w42 & ~w21623;
assign w21736 = ~w21734 & ~w21735;
assign w21737 = ~w21636 & w21736;
assign w21738 = ~w21726 & ~w21737;
assign w21739 = ~w21676 & w21719;
assign w21740 = w21738 & ~w21739;
assign w21741 = ~w80 & w21662;
assign w21742 = w21650 & w45225;
assign w21743 = ~w21663 & w21742;
assign w21744 = ~w21741 & ~w21743;
assign w21745 = (w21636 & w21743) | (w21636 & w45226) | (w21743 & w45226);
assign w21746 = w21736 & ~w21745;
assign w21747 = ~w21740 & w21746;
assign w21748 = ~w21706 & w21747;
assign w21749 = w21302 & w45227;
assign w21750 = w21357 & ~w21749;
assign w21751 = ~w21343 & w21750;
assign w21752 = ~w4056 & ~w21350;
assign w21753 = w20906 & w21579;
assign w21754 = ~w21580 & ~w21753;
assign w21755 = w3646 & w21754;
assign w21756 = ~w21752 & ~w21755;
assign w21757 = ~w21751 & w21756;
assign w21758 = ~w21598 & ~w21757;
assign w21759 = ~w21499 & w21502;
assign w21760 = ~w21503 & ~w21759;
assign w21761 = w2558 & w21760;
assign w21762 = w21513 & ~w21514;
assign w21763 = ~w21513 & w21514;
assign w21764 = w20906 & w45228;
assign w21765 = ~w3646 & w20251;
assign w21766 = w20377 & ~w21765;
assign w21767 = (w3242 & w20906) | (w3242 & w45229) | (w20906 & w45229);
assign w21768 = ~w21764 & w21767;
assign w21769 = (w20384 & ~w21565) | (w20384 & w41811) | (~w21565 & w41811);
assign w21770 = w21565 & w41812;
assign w21771 = ~w21769 & ~w21770;
assign w21772 = ~w2896 & ~w21771;
assign w21773 = w21570 & w21768;
assign w21774 = ~w21772 & ~w21773;
assign w21775 = ~w21761 & w21774;
assign w21776 = w21484 & w45230;
assign w21777 = (~w21542 & ~w21539) | (~w21542 & w47612) | (~w21539 & w47612);
assign w21778 = ~w21534 & w21777;
assign w21779 = (~w2006 & w21534) | (~w2006 & w47613) | (w21534 & w47613);
assign w21780 = ~w21776 & ~w21779;
assign w21781 = w21471 & w21780;
assign w21782 = ~w20199 & ~w21551;
assign w21783 = ~w20782 & ~w21782;
assign w21784 = ~w21549 & ~w21783;
assign w21785 = ~w21546 & w21784;
assign w21786 = ~w2285 & ~w21785;
assign w21787 = ~w21545 & w21786;
assign w21788 = w21781 & ~w21787;
assign w21789 = w21507 & w21558;
assign w21790 = ~w21775 & w21789;
assign w21791 = w21788 & ~w21790;
assign w21792 = w1120 & ~w21434;
assign w21793 = w21595 & ~w21792;
assign w21794 = ~w21428 & ~w21793;
assign w21795 = w21453 & ~w21490;
assign w21796 = ~w21791 & w21795;
assign w21797 = ~w21794 & ~w21796;
assign w21798 = w21747 & w21797;
assign w21799 = ~w21758 & w21798;
assign w21800 = ~w21748 & ~w21799;
assign w21801 = ~w21709 & ~w21800;
assign w21802 = ~w20921 & ~w20924;
assign w21803 = (~w21802 & w21800) | (~w21802 & w41813) | (w21800 & w41813);
assign w21804 = w21359 & ~w21598;
assign w21805 = ~w21241 & w21804;
assign w21806 = ~w21698 & ~w21699;
assign w21807 = ~w21796 & w41814;
assign w21808 = ~w21699 & ~w21702;
assign w21809 = ~w21691 & ~w21808;
assign w21810 = ~w21758 & w21807;
assign w21811 = (~w21809 & w21805) | (~w21809 & w45231) | (w21805 & w45231);
assign w21812 = w21803 & w21811;
assign w21813 = ~w21801 & w21811;
assign w21814 = ~w21803 & ~w21813;
assign w21815 = ~w21800 & w48974;
assign w21816 = ~w21813 & w48975;
assign w21817 = (~w21812 & ~w21814) | (~w21812 & w41815) | (~w21814 & w41815);
assign w21818 = w252 & ~w21817;
assign w21819 = ~w252 & ~w21812;
assign w21820 = ~w21816 & w21819;
assign w21821 = ~w21818 & ~w21820;
assign w21822 = ~w21758 & w21797;
assign w21823 = ~w21805 & w21822;
assign w21824 = ~w20924 & ~w21701;
assign w21825 = w21723 & w21824;
assign w21826 = w21676 & ~w21825;
assign w21827 = w21744 & ~w21826;
assign w21828 = (w21827 & w21823) | (w21827 & w41816) | (w21823 & w41816);
assign w21829 = w21719 & w21828;
assign w21830 = w21635 & w21734;
assign w21831 = w21624 & ~w21830;
assign w21832 = w21624 & w21719;
assign w21833 = w21828 & w21832;
assign w21834 = ~w21831 & ~w21833;
assign w21835 = ~w42 & w21636;
assign w21836 = ~w21829 & w21835;
assign w21837 = w21834 & ~w21836;
assign w21838 = w21635 & w21719;
assign w21839 = w21629 & ~w21630;
assign w21840 = ~w21629 & w21630;
assign w21841 = ~w21839 & ~w21840;
assign w21842 = w21801 & ~w21841;
assign w21843 = (w21838 & w21800) | (w21838 & w41817) | (w21800 & w41817);
assign w21844 = ~w21828 & w21843;
assign w21845 = (~w21838 & w21800) | (~w21838 & w41818) | (w21800 & w41818);
assign w21846 = w21828 & w21845;
assign w21847 = ~w21844 & ~w21846;
assign w21848 = ~w21842 & w21847;
assign w21849 = ~w21837 & ~w21848;
assign w21850 = ~w21805 & w48976;
assign w21851 = ~w21800 & w41819;
assign w21852 = ~w21697 & ~w21702;
assign w21853 = ~w21851 & w48977;
assign w21854 = (w21852 & w21851) | (w21852 & w48978) | (w21851 & w48978);
assign w21855 = ~w21853 & ~w21854;
assign w21856 = ~w400 & w21855;
assign w21857 = (~w21697 & w41820) | (~w21697 & w21823) | (w41820 & w21823);
assign w21858 = ~w21691 & ~w21699;
assign w21859 = ~w21690 & w21801;
assign w21860 = (~w21858 & w21800) | (~w21858 & w41821) | (w21800 & w41821);
assign w21861 = w21857 & w21860;
assign w21862 = (w21858 & w21800) | (w21858 & w41822) | (w21800 & w41822);
assign w21863 = ~w21857 & w21862;
assign w21864 = ~w21861 & ~w21863;
assign w21865 = ~w21859 & w21864;
assign w21866 = (w351 & ~w21864) | (w351 & w48979) | (~w21864 & w48979);
assign w21867 = ~w21856 & ~w21866;
assign w21868 = w400 & ~w21855;
assign w21869 = (w21419 & w21800) | (w21419 & w41823) | (w21800 & w41823);
assign w21870 = (~w612 & ~w21708) | (~w612 & w48980) | (~w21708 & w48980);
assign w21871 = ~w21800 & w21870;
assign w21872 = ~w21451 & ~w21490;
assign w21873 = ~w21490 & w21452;
assign w21874 = w21587 & w21873;
assign w21875 = ~w21254 & w48981;
assign w21876 = ~w21241 & w21875;
assign w21877 = (w21874 & w21751) | (w21874 & w41824) | (w21751 & w41824);
assign w21878 = (~w21792 & w21791) | (~w21792 & w41825) | (w21791 & w41825);
assign w21879 = ~w21593 & w21878;
assign w21880 = (w21380 & w21876) | (w21380 & w41826) | (w21876 & w41826);
assign w21881 = ~w21394 & w21419;
assign w21882 = ~w21869 & ~w21871;
assign w21883 = ~w21871 & w41827;
assign w21884 = ~w21882 & ~w21883;
assign w21885 = ~w21411 & ~w21425;
assign w21886 = ~w493 & ~w21885;
assign w21887 = w21884 & w21886;
assign w21888 = ~w493 & w21885;
assign w21889 = ~w21884 & w21888;
assign w21890 = ~w21887 & ~w21889;
assign w21891 = ~w21868 & w21890;
assign w21892 = w21867 & ~w21891;
assign w21893 = ~w21800 & w41828;
assign w21894 = (w21703 & w21805) | (w21703 & w48982) | (w21805 & w48982);
assign w21895 = (w21824 & w21800) | (w21824 & w41829) | (w21800 & w41829);
assign w21896 = ~w21894 & w21895;
assign w21897 = ~w21893 & ~w21896;
assign w21898 = ~w21675 & w21723;
assign w21899 = w57 & ~w21898;
assign w21900 = ~w21896 & w48983;
assign w21901 = w57 & w21898;
assign w21902 = (w21901 & w21896) | (w21901 & w48984) | (w21896 & w48984);
assign w21903 = ~w21900 & ~w21902;
assign w21904 = ~w21651 & ~w21742;
assign w21905 = ~w21796 & w41830;
assign w21906 = ~w21758 & w21905;
assign w21907 = ~w21805 & w21906;
assign w21908 = ~w21703 & w21825;
assign w21909 = ~w21675 & ~w21908;
assign w21910 = (w21909 & w21805) | (w21909 & w48985) | (w21805 & w48985);
assign w21911 = ~w21800 & w41831;
assign w21912 = ~w21801 & w21910;
assign w21913 = (w21904 & w21912) | (w21904 & w41832) | (w21912 & w41832);
assign w21914 = ~w21912 & w41833;
assign w21915 = ~w21913 & ~w21914;
assign w21916 = ~w80 & w21915;
assign w21917 = w21903 & ~w21916;
assign w21918 = w21864 & w48986;
assign w21919 = ~w21818 & ~w21918;
assign w21920 = w21917 & w21919;
assign w21921 = ~w21892 & w21920;
assign w21922 = ~w57 & w21898;
assign w21923 = ~w21893 & w21922;
assign w21924 = ~w21896 & w21923;
assign w21925 = ~w57 & ~w21898;
assign w21926 = w21893 & w21925;
assign w21927 = (w21925 & w21823) | (w21925 & w41834) | (w21823 & w41834);
assign w21928 = w21895 & w21927;
assign w21929 = ~w21926 & ~w21928;
assign w21930 = ~w21924 & w21929;
assign w21931 = ~w21820 & w21930;
assign w21932 = w21917 & ~w21931;
assign w21933 = ~w21663 & ~w21741;
assign w21934 = ~w21742 & ~w21933;
assign w21935 = ~w21907 & w41835;
assign w21936 = w21934 & ~w21935;
assign w21937 = w21676 & ~w21741;
assign w21938 = ~w21908 & w21937;
assign w21939 = ~w21907 & w21938;
assign w21940 = ~w21741 & w21743;
assign w21941 = (~w21940 & w21800) | (~w21940 & w41836) | (w21800 & w41836);
assign w21942 = ~w21939 & w21941;
assign w21943 = ~w21936 & w21942;
assign w21944 = w21662 & w21801;
assign w21945 = ~w3 & ~w21944;
assign w21946 = ~w21943 & w21945;
assign w21947 = w80 & w21904;
assign w21948 = (w21947 & w21912) | (w21947 & w41837) | (w21912 & w41837);
assign w21949 = w80 & ~w21904;
assign w21950 = ~w21912 & w41838;
assign w21951 = ~w21948 & ~w21950;
assign w21952 = ~w21946 & w21951;
assign w21953 = ~w21849 & w21952;
assign w21954 = ~w21932 & w21953;
assign w21955 = ~w21921 & w21954;
assign w21956 = ~w21943 & ~w21944;
assign w21957 = w3 & ~w21956;
assign w21958 = ~w21828 & ~w21838;
assign w21959 = ~w21829 & ~w21958;
assign w21960 = ~w21734 & ~w21841;
assign w21961 = w21623 & ~w21960;
assign w21962 = ~w21959 & w21961;
assign w21963 = ~w21635 & w21828;
assign w21964 = ~w21623 & ~w21963;
assign w21965 = w42 & ~w21964;
assign w21966 = ~w21962 & w21965;
assign w21967 = w21837 & ~w21966;
assign w21968 = ~w21957 & ~w21967;
assign w21969 = ~w21849 & ~w21968;
assign w21970 = ~w21955 & ~w21969;
assign w21971 = ~w21877 & w21878;
assign w21972 = w21380 & ~w21593;
assign w21973 = (w21972 & w21876) | (w21972 & w41839) | (w21876 & w41839);
assign w21974 = (w21973 & w21800) | (w21973 & w48987) | (w21800 & w48987);
assign w21975 = w945 & w21972;
assign w21976 = ~w21800 & w41840;
assign w21977 = ~w21974 & ~w21976;
assign w21978 = ~w945 & ~w21972;
assign w21979 = ~w21800 & w41841;
assign w21980 = ~w21876 & w41842;
assign w21981 = (w21980 & w21800) | (w21980 & w48988) | (w21800 & w48988);
assign w21982 = ~w21979 & ~w21981;
assign w21983 = w21977 & w21982;
assign w21984 = ~w754 & w21983;
assign w21985 = w21709 & ~w21881;
assign w21986 = (~w21881 & ~w21747) | (~w21881 & w41843) | (~w21747 & w41843);
assign w21987 = ~w21799 & w21986;
assign w21988 = ~w21985 & ~w21987;
assign w21989 = w945 & ~w20906;
assign w21990 = w20906 & w21387;
assign w21991 = ~w21989 & ~w21990;
assign w21992 = w21381 & w21991;
assign w21993 = ~w21381 & ~w21991;
assign w21994 = ~w21992 & ~w21993;
assign w21995 = ~w21880 & ~w21988;
assign w21996 = ~w21800 & w41844;
assign w21997 = ~w21995 & ~w21996;
assign w21998 = ~w21801 & w41845;
assign w21999 = w21997 & ~w21998;
assign w22000 = w21997 & w41846;
assign w22001 = ~w21984 & ~w22000;
assign w22002 = (w1320 & ~w21708) | (w1320 & w47614) | (~w21708 & w47614);
assign w22003 = ~w21800 & w22002;
assign w22004 = ~w21451 & w21470;
assign w22005 = ~w1120 & ~w22004;
assign w22006 = w21489 & ~w21780;
assign w22007 = w21465 & ~w22006;
assign w22008 = (w22007 & w21800) | (w22007 & w41847) | (w21800 & w41847);
assign w22009 = w21528 & w21585;
assign w22010 = w21357 & w22009;
assign w22011 = ~w21343 & w22010;
assign w22012 = ~w21254 & w22011;
assign w22013 = (w21507 & ~w21774) | (w21507 & w41848) | (~w21774 & w41848);
assign w22014 = ~w21786 & ~w22013;
assign w22015 = ~w22009 & w22014;
assign w22016 = w21756 & w22014;
assign w22017 = (~w22015 & w21751) | (~w22015 & w41849) | (w21751 & w41849);
assign w22018 = w21489 & w21558;
assign w22019 = w22017 & w22018;
assign w22020 = ~w21254 & w47615;
assign w22021 = ~w21241 & w22020;
assign w22022 = ~w22019 & ~w22021;
assign w22023 = ~w21800 & w47616;
assign w22024 = w22005 & w22022;
assign w22025 = w22008 & w22024;
assign w22026 = ~w22023 & ~w22025;
assign w22027 = ~w1120 & w22004;
assign w22028 = (w22027 & w21800) | (w22027 & w47617) | (w21800 & w47617);
assign w22029 = (w21800 & w47618) | (w21800 & w47619) | (w47618 & w47619);
assign w22030 = w22028 & ~w22029;
assign w22031 = w22026 & ~w22030;
assign w22032 = ~w21241 & w22012;
assign w22033 = ~w21451 & w22018;
assign w22034 = ~w21781 & w21872;
assign w22035 = ~w22033 & ~w22034;
assign w22036 = ~w22017 & ~w22034;
assign w22037 = (~w22035 & w22032) | (~w22035 & w41850) | (w22032 & w41850);
assign w22038 = ~w21801 & w41851;
assign w22039 = w22026 & w47620;
assign w22040 = ~w945 & ~w22039;
assign w22041 = w754 & ~w21983;
assign w22042 = (w945 & w41852) | (w945 & w22003) | (w41852 & w22003);
assign w22043 = w945 & w22022;
assign w22044 = w22008 & w22043;
assign w22045 = ~w22042 & ~w22044;
assign w22046 = ~w21800 & w41853;
assign w22047 = w1120 & w21434;
assign w22048 = w22037 & w22047;
assign w22049 = ~w22046 & ~w22048;
assign w22050 = ~w1120 & ~w21434;
assign w22051 = (w22050 & w21800) | (w22050 & w41854) | (w21800 & w41854);
assign w22052 = w21435 & ~w22037;
assign w22053 = w22037 & w22051;
assign w22054 = ~w22052 & ~w22053;
assign w22055 = w22026 & ~w22045;
assign w22056 = w22049 & w22054;
assign w22057 = ~w22055 & ~w22056;
assign w22058 = ~w22041 & ~w22057;
assign w22059 = ~w22040 & w22058;
assign w22060 = w22001 & ~w22059;
assign w22061 = ~w21884 & w21885;
assign w22062 = w493 & ~w22061;
assign w22063 = w21884 & ~w21885;
assign w22064 = w22062 & ~w22063;
assign w22065 = w21867 & ~w22064;
assign w22066 = w612 & ~w21999;
assign w22067 = w21931 & ~w22066;
assign w22068 = w21953 & w22067;
assign w22069 = w22065 & w22068;
assign w22070 = ~w22060 & w22069;
assign w22071 = (w22009 & w21751) | (w22009 & w41855) | (w21751 & w41855);
assign w22072 = ~w22013 & ~w22071;
assign w22073 = ~w22032 & w22072;
assign w22074 = ~w22032 & w41856;
assign w22075 = ~w21801 & ~w22074;
assign w22076 = ~w2285 & ~w22073;
assign w22077 = (w21785 & ~w22075) | (w21785 & w41857) | (~w22075 & w41857);
assign w22078 = w22075 & w41858;
assign w22079 = ~w22077 & ~w22078;
assign w22080 = ~w21557 & w21786;
assign w22081 = w21507 & ~w21557;
assign w22082 = (w22081 & ~w21774) | (w22081 & w41859) | (~w21774 & w41859);
assign w22083 = ~w22080 & ~w22082;
assign w22084 = ~w21557 & w21570;
assign w22085 = w21528 & w22084;
assign w22086 = w22083 & ~w22085;
assign w22087 = w21584 & ~w22086;
assign w22088 = w21359 & w22087;
assign w22089 = ~w21241 & w22088;
assign w22090 = w21584 & w22085;
assign w22091 = w22083 & ~w22090;
assign w22092 = w21756 & w22083;
assign w22093 = (~w22091 & w21751) | (~w22091 & w41860) | (w21751 & w41860);
assign w22094 = ~w2006 & w21778;
assign w22095 = ~w22093 & ~w22094;
assign w22096 = ~w22089 & w22095;
assign w22097 = w21558 & w22017;
assign w22098 = ~w21254 & w45232;
assign w22099 = ~w21241 & w22098;
assign w22100 = ~w22097 & ~w22099;
assign w22101 = ~w22096 & w22100;
assign w22102 = ~w21801 & w22101;
assign w22103 = w2006 & ~w22093;
assign w22104 = ~w22089 & w22103;
assign w22105 = ~w22089 & w41861;
assign w22106 = ~w21709 & ~w21778;
assign w22107 = ~w21800 & w22106;
assign w22108 = ~w22105 & ~w22107;
assign w22109 = w21779 & ~w21785;
assign w22110 = ~w21800 & w41862;
assign w22111 = (w21779 & w22089) | (w21779 & w41863) | (w22089 & w41863);
assign w22112 = ~w2339 & ~w22111;
assign w22113 = ~w22110 & w22112;
assign w22114 = (~w1738 & w22107) | (~w1738 & w41864) | (w22107 & w41864);
assign w22115 = w22113 & ~w22114;
assign w22116 = ~w2340 & w22102;
assign w22117 = w22115 & ~w22116;
assign w22118 = w22079 & ~w22117;
assign w22119 = ~w21801 & ~w22104;
assign w22120 = ~w22102 & w22119;
assign w22121 = ~w21800 & w41865;
assign w22122 = ~w21485 & ~w21776;
assign w22123 = ~w1541 & w22122;
assign w22124 = ~w22121 & w22123;
assign w22125 = ~w22120 & w22124;
assign w22126 = ~w1541 & ~w22122;
assign w22127 = (w22126 & w22089) | (w22126 & w41866) | (w22089 & w41866);
assign w22128 = ~w21801 & w22127;
assign w22129 = ~w1541 & w21776;
assign w22130 = w21801 & w22129;
assign w22131 = ~w22102 & w22128;
assign w22132 = ~w22130 & ~w22131;
assign w22133 = ~w22125 & w22132;
assign w22134 = ~w22102 & w22108;
assign w22135 = (~w1738 & ~w22134) | (~w1738 & w41867) | (~w22134 & w41867);
assign w22136 = w22133 & ~w22135;
assign w22137 = ~w22118 & w22136;
assign w22138 = w1541 & w22122;
assign w22139 = (w22138 & w22120) | (w22138 & w41868) | (w22120 & w41868);
assign w22140 = w1541 & ~w22122;
assign w22141 = ~w22120 & w41869;
assign w22142 = ~w22139 & ~w22141;
assign w22143 = (~w1541 & ~w21708) | (~w1541 & w45233) | (~w21708 & w45233);
assign w22144 = ~w21800 & w22143;
assign w22145 = (w21780 & w21800) | (w21780 & w45234) | (w21800 & w45234);
assign w22146 = ~w22144 & w41870;
assign w22147 = ~w21800 & w41871;
assign w22148 = (w21485 & w21800) | (w21485 & w41872) | (w21800 & w41872);
assign w22149 = ~w22147 & ~w22148;
assign w22150 = ~w22146 & w22149;
assign w22151 = w21465 & ~w21488;
assign w22152 = w1320 & ~w22151;
assign w22153 = ~w22150 & w22152;
assign w22154 = w1320 & w22151;
assign w22155 = w22150 & w22154;
assign w22156 = ~w22153 & ~w22155;
assign w22157 = w22142 & w22156;
assign w22158 = ~w22137 & w22157;
assign w22159 = ~w1320 & ~w22151;
assign w22160 = ~w1541 & w22159;
assign w22161 = ~w21800 & w41873;
assign w22162 = ~w21485 & w22159;
assign w22163 = (w22162 & w21800) | (w22162 & w41874) | (w21800 & w41874);
assign w22164 = ~w22161 & ~w22163;
assign w22165 = ~w1320 & w22151;
assign w22166 = w1541 & w22165;
assign w22167 = ~w21800 & w41875;
assign w22168 = w21485 & w22165;
assign w22169 = (w22168 & w21800) | (w22168 & w41876) | (w21800 & w41876);
assign w22170 = ~w22167 & ~w22169;
assign w22171 = w22100 & w22165;
assign w22172 = w22145 & w22171;
assign w22173 = w22170 & ~w22172;
assign w22174 = ~w22146 & ~w22164;
assign w22175 = w22173 & ~w22174;
assign w22176 = ~w22021 & w41877;
assign w22177 = ~w21801 & w22176;
assign w22178 = w1120 & w22004;
assign w22179 = (w22178 & w22177) | (w22178 & w41878) | (w22177 & w41878);
assign w22180 = w1120 & ~w22004;
assign w22181 = ~w22177 & w41879;
assign w22182 = ~w22179 & ~w22181;
assign w22183 = w22175 & w22182;
assign w22184 = w22001 & w22183;
assign w22185 = ~w22038 & w22049;
assign w22186 = w22054 & w22185;
assign w22187 = w945 & w22186;
assign w22188 = ~w22041 & w22187;
assign w22189 = w22184 & ~w22188;
assign w22190 = ~w22158 & w22189;
assign w22191 = w22134 & w41880;
assign w22192 = w2006 & w21785;
assign w22193 = (w22192 & ~w22075) | (w22192 & w41881) | (~w22075 & w41881);
assign w22194 = w2006 & ~w21785;
assign w22195 = w22075 & w41882;
assign w22196 = ~w22193 & ~w22195;
assign w22197 = ~w22191 & w22196;
assign w22198 = w22136 & ~w22197;
assign w22199 = w22157 & ~w22198;
assign w22200 = w22001 & w23685;
assign w22201 = ~w22199 & w22200;
assign w22202 = w22190 & w22201;
assign w22203 = w22070 & ~w22202;
assign w22204 = w21970 & ~w22203;
assign w22205 = ~w22190 & ~w22201;
assign w22206 = w22070 & w22205;
assign w22207 = w21970 & ~w22206;
assign w22208 = ~a[30] & ~a[31];
assign w22209 = ~a[32] & w22208;
assign w22210 = ~w20906 & ~w22209;
assign w22211 = a[33] & w22210;
assign w22212 = ~w21039 & ~w22211;
assign w22213 = w20906 & w22209;
assign w22214 = w20000 & ~w22213;
assign w22215 = ~a[33] & ~w22210;
assign w22216 = w22214 & ~w22215;
assign w22217 = ~w21800 & w41883;
assign w22218 = ~w22212 & w22214;
assign w22219 = (w22218 & w21800) | (w22218 & w41884) | (w21800 & w41884);
assign w22220 = ~w22217 & ~w22219;
assign w22221 = ~a[34] & w20906;
assign w22222 = a[34] & ~w20906;
assign w22223 = a[34] & ~w21039;
assign w22224 = ~w21040 & ~w22223;
assign w22225 = ~w22221 & ~w22222;
assign w22226 = ~w21800 & w41885;
assign w22227 = (w22224 & w21800) | (w22224 & w41886) | (w21800 & w41886);
assign w22228 = ~w22226 & ~w22227;
assign w22229 = ~w22212 & ~w22213;
assign w22230 = ~w20000 & w50207;
assign w22231 = ~w22213 & ~w22215;
assign w22232 = ~w21800 & w45235;
assign w22233 = w22230 & ~w22232;
assign w22234 = w22220 & ~w22228;
assign w22235 = ~w22233 & ~w22234;
assign w22236 = ~w21041 & ~w21047;
assign w22237 = w20906 & ~w22236;
assign w22238 = ~w20906 & w22236;
assign w22239 = ~w22237 & ~w22238;
assign w22240 = ~w21800 & w41888;
assign w22241 = (~w22239 & w21800) | (~w22239 & w41889) | (w21800 & w41889);
assign w22242 = ~w22240 & ~w22241;
assign w22243 = a[35] & ~w19040;
assign w22244 = w20413 & w22242;
assign w22245 = ~w22242 & w22243;
assign w22246 = ~w22244 & ~w22245;
assign w22247 = w22235 & w22246;
assign w22248 = ~a[35] & w19040;
assign w22249 = ~w22242 & w22248;
assign w22250 = a[35] & w19040;
assign w22251 = w22242 & w22250;
assign w22252 = ~w22249 & ~w22251;
assign w22253 = ~w19040 & w21054;
assign w22254 = w19040 & ~w21054;
assign w22255 = ~w22253 & ~w22254;
assign w22256 = w21038 & w50208;
assign w22257 = (w21800 & w48989) | (w21800 & w48990) | (w48989 & w48990);
assign w22258 = ~w22256 & ~w22257;
assign w22259 = w18183 & ~w22258;
assign w22260 = w22252 & ~w22259;
assign w22261 = ~w22247 & w22260;
assign w22262 = ~w21031 & w21063;
assign w22263 = w21058 & ~w22262;
assign w22264 = ~w21058 & w22262;
assign w22265 = ~w22263 & ~w22264;
assign w22266 = ~w21022 & ~w21029;
assign w22267 = ~w21800 & w45236;
assign w22268 = (w22265 & w21800) | (w22265 & w45237) | (w21800 & w45237);
assign w22269 = ~w22267 & ~w22268;
assign w22270 = w17380 & ~w22269;
assign w22271 = ~w18183 & w22258;
assign w22272 = ~w22270 & ~w22271;
assign w22273 = ~w22261 & w22272;
assign w22274 = ~w21800 & w41891;
assign w22275 = ~w21059 & w21063;
assign w22276 = ~w17380 & w21120;
assign w22277 = ~w21121 & ~w22276;
assign w22278 = w22275 & ~w22277;
assign w22279 = ~w22275 & w22277;
assign w22280 = ~w22278 & ~w22279;
assign w22281 = (w22280 & w21800) | (w22280 & w41892) | (w21800 & w41892);
assign w22282 = ~w22274 & ~w22281;
assign w22283 = ~w21086 & ~w21121;
assign w22284 = (w21131 & w22274) | (w21131 & w45238) | (w22274 & w45238);
assign w22285 = w15681 & w22280;
assign w22286 = w21125 & ~w22283;
assign w22287 = ~w22285 & ~w22286;
assign w22288 = w16559 & ~w22287;
assign w22289 = ~w21801 & w22288;
assign w22290 = ~w22284 & ~w22289;
assign w22291 = ~w15681 & w22282;
assign w22292 = ~w22290 & ~w22291;
assign w22293 = ~w17380 & w22269;
assign w22294 = ~w16559 & ~w22283;
assign w22295 = w16559 & w21120;
assign w22296 = w21125 & ~w22295;
assign w22297 = w15681 & w21126;
assign w22298 = (w21800 & w48991) | (w21800 & w48992) | (w48991 & w48992);
assign w22299 = w15681 & ~w22296;
assign w22300 = w22299 & w52250;
assign w22301 = ~w22298 & ~w22300;
assign w22302 = ~w22293 & w22301;
assign w22303 = ~w22292 & w22302;
assign w22304 = (w22303 & w22261) | (w22303 & w45239) | (w22261 & w45239);
assign w22305 = w21141 & ~w21243;
assign w22306 = w9781 & ~w22305;
assign w22307 = ~w9781 & w22305;
assign w22308 = ~w22306 & ~w22307;
assign w22309 = ~w21226 & ~w21233;
assign w22310 = ~w9195 & ~w22309;
assign w22311 = (w22310 & w21801) | (w22310 & w41894) | (w21801 & w41894);
assign w22312 = ~w9195 & w22309;
assign w22313 = ~w21801 & w41895;
assign w22314 = ~w22311 & ~w22313;
assign w22315 = ~w21006 & w41896;
assign w22316 = ~w21140 & w22315;
assign w22317 = ~w21235 & ~w22316;
assign w22318 = ~w9195 & w22317;
assign w22319 = w9195 & ~w22317;
assign w22320 = ~w22318 & ~w22319;
assign w22321 = w8666 & w21221;
assign w22322 = (w22321 & w21801) | (w22321 & w41897) | (w21801 & w41897);
assign w22323 = w8666 & ~w21221;
assign w22324 = ~w21801 & w41898;
assign w22325 = ~w22322 & ~w22324;
assign w22326 = w22314 & w22325;
assign w22327 = ~w20516 & ~w20968;
assign w22328 = w20516 & w20968;
assign w22329 = ~w22327 & ~w22328;
assign w22330 = ~w12666 & ~w22329;
assign w22331 = ~w14303 & w22329;
assign w22332 = ~w22330 & ~w22331;
assign w22333 = ~w21129 & ~w21134;
assign w22334 = (~w20998 & w21129) | (~w20998 & w41899) | (w21129 & w41899);
assign w22335 = w20973 & w21136;
assign w22336 = ~w22334 & w22335;
assign w22337 = w22332 & ~w22336;
assign w22338 = ~w22332 & w22336;
assign w22339 = ~w22337 & ~w22338;
assign w22340 = (~w22339 & w21800) | (~w22339 & w41900) | (w21800 & w41900);
assign w22341 = ~w11870 & ~w20980;
assign w22342 = ~w22340 & w22341;
assign w22343 = ~w11870 & w20980;
assign w22344 = w22340 & w22343;
assign w22345 = ~w22342 & ~w22344;
assign w22346 = w14039 & ~w22333;
assign w22347 = ~w14039 & w22333;
assign w22348 = ~w22346 & ~w22347;
assign w22349 = w13384 & w20997;
assign w22350 = ~w22348 & w22349;
assign w22351 = (w22350 & w21800) | (w22350 & w41901) | (w21800 & w41901);
assign w22352 = w13384 & ~w20997;
assign w22353 = (w22352 & ~w21708) | (w22352 & w45240) | (~w21708 & w45240);
assign w22354 = w22348 & w22352;
assign w22355 = (~w22354 & w21800) | (~w22354 & w45241) | (w21800 & w45241);
assign w22356 = ~w22351 & w22355;
assign w22357 = w20973 & w20987;
assign w22358 = ~w21135 & ~w22334;
assign w22359 = ~w22357 & ~w22358;
assign w22360 = ~w22336 & ~w22359;
assign w22361 = ~w21800 & w41902;
assign w22362 = ~w12666 & ~w22360;
assign w22363 = ~w21801 & w22362;
assign w22364 = ~w22361 & ~w22363;
assign w22365 = w22356 & w22364;
assign w22366 = w22345 & w22365;
assign w22367 = (~w22348 & w21800) | (~w22348 & w41903) | (w21800 & w41903);
assign w22368 = ~w13384 & w20997;
assign w22369 = ~w22367 & w22368;
assign w22370 = ~w13384 & ~w20997;
assign w22371 = w22367 & w22370;
assign w22372 = ~w22369 & ~w22371;
assign w22373 = (~w21131 & w21086) | (~w21131 & w41904) | (w21086 & w41904);
assign w22374 = w15681 & ~w22373;
assign w22375 = ~w15681 & w22373;
assign w22376 = ~w21101 & ~w22375;
assign w22377 = ~w22374 & ~w22376;
assign w22378 = ~w14766 & w22377;
assign w22379 = w14766 & ~w22377;
assign w22380 = ~w22378 & ~w22379;
assign w22381 = ~w21801 & w22380;
assign w22382 = w14039 & ~w21115;
assign w22383 = (w22382 & w21801) | (w22382 & w41905) | (w21801 & w41905);
assign w22384 = w14039 & w21115;
assign w22385 = ~w21801 & w41906;
assign w22386 = ~w22383 & ~w22385;
assign w22387 = w22372 & w22386;
assign w22388 = ~w20961 & ~w21001;
assign w22389 = w21136 & ~w22334;
assign w22390 = w20982 & ~w22389;
assign w22391 = ~w21002 & ~w22390;
assign w22392 = ~w22388 & w22391;
assign w22393 = w22388 & ~w22391;
assign w22394 = ~w21800 & w48993;
assign w22395 = ~w21801 & w41907;
assign w22396 = ~w22394 & ~w22395;
assign w22397 = ~w11138 & w22396;
assign w22398 = w11870 & ~w20980;
assign w22399 = ~w22339 & ~w22398;
assign w22400 = w11870 & w20980;
assign w22401 = w22339 & ~w22400;
assign w22402 = (~w22400 & ~w21708) | (~w22400 & w45242) | (~w21708 & w45242);
assign w22403 = ~w21800 & w22402;
assign w22404 = ~w22401 & ~w22403;
assign w22405 = ~w21801 & w22399;
assign w22406 = w22404 & ~w22405;
assign w22407 = w12666 & w22329;
assign w22408 = ~w21800 & w41908;
assign w22409 = w12666 & w22360;
assign w22410 = ~w21801 & w22409;
assign w22411 = ~w22408 & ~w22410;
assign w22412 = ~w22406 & w22411;
assign w22413 = w22345 & ~w22412;
assign w22414 = ~w22397 & ~w22413;
assign w22415 = w22366 & ~w22387;
assign w22416 = w22414 & ~w22415;
assign w22417 = w21003 & ~w21137;
assign w22418 = ~w21129 & w41909;
assign w22419 = ~w21000 & w21003;
assign w22420 = ~w20934 & w20963;
assign w22421 = ~w22419 & w22420;
assign w22422 = ~w22418 & w22421;
assign w22423 = ~w20948 & ~w21243;
assign w22424 = w20934 & ~w22423;
assign w22425 = ~w20934 & w22423;
assign w22426 = ~w22424 & ~w22425;
assign w22427 = w22422 & ~w22426;
assign w22428 = ~w22422 & w22426;
assign w22429 = ~w22427 & ~w22428;
assign w22430 = ~w21800 & w41910;
assign w22431 = (~w22429 & w21800) | (~w22429 & w41911) | (w21800 & w41911);
assign w22432 = ~w22430 & ~w22431;
assign w22433 = ~w9781 & w22432;
assign w22434 = ~w20961 & ~w22419;
assign w22435 = (w22434 & w21129) | (w22434 & w48994) | (w21129 & w48994);
assign w22436 = ~w11138 & w22435;
assign w22437 = w11138 & ~w22435;
assign w22438 = ~w22436 & ~w22437;
assign w22439 = w10419 & w20933;
assign w22440 = ~w22438 & w22439;
assign w22441 = (w22440 & w21800) | (w22440 & w48995) | (w21800 & w48995);
assign w22442 = w10419 & ~w20933;
assign w22443 = (w22442 & ~w21708) | (w22442 & w45243) | (~w21708 & w45243);
assign w22444 = w22438 & w22442;
assign w22445 = (~w22444 & w21800) | (~w22444 & w48996) | (w21800 & w48996);
assign w22446 = ~w22441 & w22445;
assign w22447 = w9781 & w20947;
assign w22448 = ~w21800 & w41912;
assign w22449 = w9781 & ~w22429;
assign w22450 = ~w21801 & w22449;
assign w22451 = ~w22448 & ~w22450;
assign w22452 = w22446 & w22451;
assign w22453 = ~w22433 & ~w22452;
assign w22454 = ~w16559 & w22282;
assign w22455 = ~w16559 & w22283;
assign w22456 = w16559 & ~w22283;
assign w22457 = ~w22455 & ~w22456;
assign w22458 = (~w22457 & w21800) | (~w22457 & w41913) | (w21800 & w41913);
assign w22459 = ~w15681 & w21125;
assign w22460 = w22459 & ~w22458;
assign w22461 = ~w15681 & ~w21125;
assign w22462 = (w21800 & w48997) | (w21800 & w48998) | (w48997 & w48998);
assign w22463 = ~w22460 & ~w22462;
assign w22464 = ~w22374 & ~w22375;
assign w22465 = (w22464 & w21800) | (w22464 & w41914) | (w21800 & w41914);
assign w22466 = ~w14766 & w21101;
assign w22467 = w22466 & ~w22465;
assign w22468 = ~w14766 & ~w21101;
assign w22469 = (w21800 & w48999) | (w21800 & w49000) | (w48999 & w49000);
assign w22470 = ~w22467 & ~w22469;
assign w22471 = w22463 & w22470;
assign w22472 = w22301 & w22454;
assign w22473 = w22471 & ~w22472;
assign w22474 = ~w22453 & w22473;
assign w22475 = w22416 & w22474;
assign w22476 = w22416 & w41915;
assign w22477 = ~w22304 & w22476;
assign w22478 = w22326 & ~w22453;
assign w22479 = (w11138 & w22395) | (w11138 & w49001) | (w22395 & w49001);
assign w22480 = (~w22438 & w21800) | (~w22438 & w41916) | (w21800 & w41916);
assign w22481 = w20933 & ~w22480;
assign w22482 = ~w20933 & w22480;
assign w22483 = ~w22481 & ~w22482;
assign w22484 = ~w10419 & ~w22483;
assign w22485 = ~w22479 & ~w22484;
assign w22486 = ~w22484 & w49002;
assign w22487 = ~w14039 & w21115;
assign w22488 = (w22487 & w21801) | (w22487 & w41917) | (w21801 & w41917);
assign w22489 = ~w14039 & ~w21115;
assign w22490 = ~w21801 & w41918;
assign w22491 = ~w22488 & ~w22490;
assign w22492 = w14766 & ~w21101;
assign w22493 = ~w22465 & w22492;
assign w22494 = w14766 & w21101;
assign w22495 = w22465 & w22494;
assign w22496 = ~w22493 & ~w22495;
assign w22497 = w22491 & w22496;
assign w22498 = w22366 & w22497;
assign w22499 = w22478 & ~w22486;
assign w22500 = w22478 & ~w22498;
assign w22501 = w22416 & w22500;
assign w22502 = ~w22499 & ~w22501;
assign w22503 = ~w21801 & w41919;
assign w22504 = (w22309 & w21801) | (w22309 & w41920) | (w21801 & w41920);
assign w22505 = ~w22503 & ~w22504;
assign w22506 = w9195 & ~w22505;
assign w22507 = w22325 & w22506;
assign w22508 = ~w21189 & ~w21191;
assign w22509 = w21181 & w52251;
assign w22510 = w8666 & ~w22509;
assign w22511 = ~w8666 & w22509;
assign w22512 = ~w22510 & ~w22511;
assign w22513 = (w22508 & w21801) | (w22508 & w41922) | (w21801 & w41922);
assign w22514 = ~w21801 & w41923;
assign w22515 = ~w22513 & ~w22514;
assign w22516 = (w21221 & w21801) | (w21221 & w41924) | (w21801 & w41924);
assign w22517 = ~w21801 & w41925;
assign w22518 = ~w22516 & ~w22517;
assign w22519 = ~w8666 & w22518;
assign w22520 = ~w7924 & ~w22515;
assign w22521 = ~w22519 & ~w22520;
assign w22522 = ~w22507 & w22521;
assign w22523 = ~w21211 & ~w21215;
assign w22524 = w21195 & ~w21197;
assign w22525 = ~w21197 & w21237;
assign w22526 = (w22525 & w21140) | (w22525 & w41926) | (w21140 & w41926);
assign w22527 = ~w22524 & ~w22526;
assign w22528 = w22523 & ~w22527;
assign w22529 = ~w22523 & w22527;
assign w22530 = ~w22528 & ~w22529;
assign w22531 = ~w21800 & w41927;
assign w22532 = ~w21801 & w22530;
assign w22533 = ~w22531 & ~w22532;
assign w22534 = ~w22532 & w41928;
assign w22535 = ~w21299 & ~w21339;
assign w22536 = ~w21254 & w22535;
assign w22537 = w21254 & ~w22535;
assign w22538 = ~w21239 & w41929;
assign w22539 = ~w21141 & w22538;
assign w22540 = ~w22537 & ~w22539;
assign w22541 = ~w21241 & w22536;
assign w22542 = w22540 & ~w22541;
assign w22543 = ~w21800 & w41930;
assign w22544 = (w22542 & w21800) | (w22542 & w47621) | (w21800 & w47621);
assign w22545 = ~w22543 & ~w22544;
assign w22546 = ~w22544 & w41931;
assign w22547 = ~w21284 & ~w21301;
assign w22548 = (~w21299 & w21254) | (~w21299 & w41932) | (w21254 & w41932);
assign w22549 = ~w21239 & w41933;
assign w22550 = ~w21141 & w22549;
assign w22551 = ~w22550 & w41934;
assign w22552 = (w22547 & w22550) | (w22547 & w41935) | (w22550 & w41935);
assign w22553 = ~w21800 & w45244;
assign w22554 = ~w22551 & ~w22552;
assign w22555 = ~w21801 & w22554;
assign w22556 = (w5330 & w22555) | (w5330 & w45245) | (w22555 & w45245);
assign w22557 = ~w22546 & ~w22556;
assign w22558 = (~w21168 & ~w21708) | (~w21168 & w45246) | (~w21708 & w45246);
assign w22559 = ~w21800 & w22558;
assign w22560 = ~w21169 & ~w21216;
assign w22561 = ~w21213 & ~w21215;
assign w22562 = (w21238 & w21140) | (w21238 & w41936) | (w21140 & w41936);
assign w22563 = w22561 & ~w22562;
assign w22564 = w22560 & ~w22563;
assign w22565 = ~w22560 & w22563;
assign w22566 = ~w22564 & ~w22565;
assign w22567 = ~w21801 & w22566;
assign w22568 = ~w22559 & ~w22567;
assign w22569 = (~w6769 & w22567) | (~w6769 & w41937) | (w22567 & w41937);
assign w22570 = w21238 & w22560;
assign w22571 = w22561 & w22570;
assign w22572 = (w22571 & w21140) | (w22571 & w41938) | (w21140 & w41938);
assign w22573 = ~w21160 & ~w21242;
assign w22574 = ~w21169 & ~w21218;
assign w22575 = w22573 & ~w22574;
assign w22576 = ~w22573 & w22574;
assign w22577 = ~w22575 & ~w22576;
assign w22578 = w22572 & w22573;
assign w22579 = ~w22572 & w22577;
assign w22580 = ~w22578 & ~w22579;
assign w22581 = w6264 & w21159;
assign w22582 = ~w21800 & w41939;
assign w22583 = w6264 & w22580;
assign w22584 = ~w21801 & w22583;
assign w22585 = ~w22582 & ~w22584;
assign w22586 = ~w22569 & w22585;
assign w22587 = w22557 & w22586;
assign w22588 = (w6769 & w21800) | (w6769 & w45247) | (w21800 & w45247);
assign w22589 = ~w22567 & w22588;
assign w22590 = w5745 & ~w21298;
assign w22591 = ~w21800 & w41940;
assign w22592 = w5745 & w22542;
assign w22593 = ~w21801 & w22592;
assign w22594 = ~w22591 & ~w22593;
assign w22595 = ~w6264 & ~w21159;
assign w22596 = ~w21800 & w41941;
assign w22597 = ~w6264 & ~w22580;
assign w22598 = ~w21801 & w22597;
assign w22599 = ~w22596 & ~w22598;
assign w22600 = w22594 & w22599;
assign w22601 = w22585 & w22589;
assign w22602 = w22600 & ~w22601;
assign w22603 = ~w21273 & ~w21300;
assign w22604 = ~w21800 & w41942;
assign w22605 = ~w21284 & ~w22552;
assign w22606 = ~w21801 & w22605;
assign w22607 = ~w22604 & ~w22606;
assign w22608 = ~w22555 & w45248;
assign w22609 = w4838 & w22603;
assign w22610 = w22607 & w22609;
assign w22611 = w4838 & ~w22603;
assign w22612 = (w22611 & w22606) | (w22611 & w41943) | (w22606 & w41943);
assign w22613 = ~w22608 & ~w22612;
assign w22614 = ~w22610 & w22613;
assign w22615 = w22557 & ~w22602;
assign w22616 = w22614 & ~w22615;
assign w22617 = w22557 & w41944;
assign w22618 = w22616 & w41945;
assign w22619 = w22502 & w22618;
assign w22620 = ~w22477 & w22619;
assign w22621 = ~w21254 & w47622;
assign w22622 = ~w21241 & w22621;
assign w22623 = w21584 & ~w21757;
assign w22624 = ~w22622 & w41946;
assign w22625 = ~w2896 & w21527;
assign w22626 = ~w22624 & w22625;
assign w22627 = ~w21801 & ~w22626;
assign w22628 = w21527 & ~w22624;
assign w22629 = w2896 & ~w22628;
assign w22630 = w2896 & ~w21771;
assign w22631 = (w22630 & w21800) | (w22630 & w41947) | (w21800 & w41947);
assign w22632 = w22628 & w22631;
assign w22633 = (w21772 & w21800) | (w21772 & w41948) | (w21800 & w41948);
assign w22634 = ~w22628 & w22633;
assign w22635 = ~w22632 & ~w22634;
assign w22636 = (w21771 & ~w22627) | (w21771 & w47623) | (~w22627 & w47623);
assign w22637 = w22635 & ~w22636;
assign w22638 = w2558 & w22637;
assign w22639 = ~w21800 & w47624;
assign w22640 = ~w22627 & ~w22639;
assign w22641 = w22635 & ~w22640;
assign w22642 = w21507 & ~w21761;
assign w22643 = ~w2285 & ~w22642;
assign w22644 = ~w22641 & w22643;
assign w22645 = ~w2285 & w22642;
assign w22646 = w22641 & w22645;
assign w22647 = ~w22644 & ~w22646;
assign w22648 = ~w22638 & w22647;
assign w22649 = w2285 & w22642;
assign w22650 = ~w22641 & w22649;
assign w22651 = w2285 & ~w22642;
assign w22652 = w22641 & w22651;
assign w22653 = ~w22650 & ~w22652;
assign w22654 = w3646 & ~w20906;
assign w22655 = w20906 & w21513;
assign w22656 = ~w22654 & ~w22655;
assign w22657 = ~w21514 & ~w22656;
assign w22658 = w21514 & w22656;
assign w22659 = ~w22657 & ~w22658;
assign w22660 = ~w21800 & w41949;
assign w22661 = w21527 & ~w21768;
assign w22662 = (w22661 & w22622) | (w22661 & w41950) | (w22622 & w41950);
assign w22663 = (~w22662 & w21800) | (~w22662 & w47625) | (w21800 & w47625);
assign w22664 = ~w22622 & w41951;
assign w22665 = ~w21800 & w49003;
assign w22666 = ~w2896 & ~w22664;
assign w22667 = w22663 & w22666;
assign w22668 = ~w22665 & ~w22667;
assign w22669 = ~w21239 & w41952;
assign w22670 = ~w21141 & w22669;
assign w22671 = ~w21253 & w49004;
assign w22672 = ~w21343 & w41953;
assign w22673 = ~w22671 & w22672;
assign w22674 = ~w22670 & w22673;
assign w22675 = ~w3646 & w21752;
assign w22676 = ~w3646 & w22674;
assign w22677 = w3646 & ~w21752;
assign w22678 = ~w22674 & w22677;
assign w22679 = ~w22676 & ~w22678;
assign w22680 = ~w22675 & w22679;
assign w22681 = ~w3242 & ~w21754;
assign w22682 = (w22681 & w22680) | (w22681 & w41954) | (w22680 & w41954);
assign w22683 = ~w3242 & w21754;
assign w22684 = ~w22680 & w41955;
assign w22685 = ~w22682 & ~w22684;
assign w22686 = w2896 & ~w22660;
assign w22687 = w22663 & ~w22664;
assign w22688 = w22686 & ~w22687;
assign w22689 = w22685 & ~w22688;
assign w22690 = w22668 & ~w22689;
assign w22691 = w3242 & w21754;
assign w22692 = (w22691 & w22680) | (w22691 & w41956) | (w22680 & w41956);
assign w22693 = w3242 & ~w21754;
assign w22694 = ~w22680 & w41957;
assign w22695 = ~w22692 & ~w22694;
assign w22696 = ~w21343 & w21356;
assign w22697 = ~w22671 & w22696;
assign w22698 = ~w22670 & w22697;
assign w22699 = ~w21351 & ~w21752;
assign w22700 = ~w22698 & ~w22699;
assign w22701 = ~w21800 & w41958;
assign w22702 = ~w22674 & ~w22700;
assign w22703 = ~w21801 & w22702;
assign w22704 = ~w22701 & ~w22703;
assign w22705 = (w3646 & w22703) | (w3646 & w41959) | (w22703 & w41959);
assign w22706 = w22668 & ~w22705;
assign w22707 = w22695 & w22706;
assign w22708 = ~w21800 & w49005;
assign w22709 = ~w21337 & ~w21353;
assign w22710 = ~w21254 & w21341;
assign w22711 = ~w21241 & w22710;
assign w22712 = ~w21304 & ~w21316;
assign w22713 = (w22712 & w21241) | (w22712 & w41960) | (w21241 & w41960);
assign w22714 = ~w21354 & ~w22713;
assign w22715 = w22709 & ~w22714;
assign w22716 = ~w21801 & ~w22715;
assign w22717 = ~w22709 & w22714;
assign w22718 = w4056 & w22708;
assign w22719 = w4056 & ~w22717;
assign w22720 = w22716 & w22719;
assign w22721 = ~w22718 & ~w22720;
assign w22722 = ~w22703 & w49006;
assign w22723 = w22721 & ~w22722;
assign w22724 = w22707 & ~w22723;
assign w22725 = ~w22690 & ~w22724;
assign w22726 = ~w2558 & ~w22637;
assign w22727 = ~w22648 & w22653;
assign w22728 = w22653 & ~w22726;
assign w22729 = w22725 & w22728;
assign w22730 = ~w22727 & ~w22729;
assign w22731 = ~w21801 & w45249;
assign w22732 = ~w22708 & ~w22731;
assign w22733 = ~w4056 & w22732;
assign w22734 = ~w21316 & ~w21354;
assign w22735 = ~w21304 & ~w22711;
assign w22736 = (w22735 & w21800) | (w22735 & w45250) | (w21800 & w45250);
assign w22737 = (w22734 & w22736) | (w22734 & w41962) | (w22736 & w41962);
assign w22738 = ~w22736 & w41963;
assign w22739 = ~w22737 & ~w22738;
assign w22740 = ~w4430 & ~w22739;
assign w22741 = ~w22733 & ~w22740;
assign w22742 = w22707 & w22741;
assign w22743 = w22648 & w22742;
assign w22744 = (~w22743 & w22729) | (~w22743 & w41964) | (w22729 & w41964);
assign w22745 = w22620 & ~w22744;
assign w22746 = w7924 & ~w22508;
assign w22747 = (w22746 & w21801) | (w22746 & w41965) | (w21801 & w41965);
assign w22748 = w7924 & w22508;
assign w22749 = ~w21801 & w41966;
assign w22750 = ~w22747 & ~w22749;
assign w22751 = ~w22534 & ~w22750;
assign w22752 = (w7315 & w22532) | (w7315 & w47626) | (w22532 & w47626);
assign w22753 = ~w22751 & ~w22752;
assign w22754 = w22587 & w22753;
assign w22755 = w22616 & ~w22754;
assign w22756 = (w22603 & w22606) | (w22603 & w45251) | (w22606 & w45251);
assign w22757 = ~w22606 & w45252;
assign w22758 = ~w22756 & ~w22757;
assign w22759 = ~w4838 & ~w22758;
assign w22760 = w4430 & w22739;
assign w22761 = ~w22759 & ~w22760;
assign w22762 = (w22761 & ~w22616) | (w22761 & w45253) | (~w22616 & w45253);
assign w22763 = w22743 & ~w22762;
assign w22764 = ~w22730 & ~w22763;
assign w22765 = (w22764 & ~w22620) | (w22764 & w47627) | (~w22620 & w47627);
assign w22766 = w22207 & ~w22765;
assign w22767 = (~w22204 & w22765) | (~w22204 & w41967) | (w22765 & w41967);
assign w22768 = ~w22158 & ~w22199;
assign w22769 = ~w22730 & w45254;
assign w22770 = (~w22066 & w22059) | (~w22066 & w47628) | (w22059 & w47628);
assign w22771 = w22065 & w22770;
assign w22772 = (~w22745 & w45255) | (~w22745 & w45256) | (w45255 & w45256);
assign w22773 = ~w21892 & ~w21918;
assign w22774 = (~w41967 & w47629) | (~w41967 & w47630) | (w47629 & w47630);
assign w22775 = w22767 & w45257;
assign w22776 = ~w22775 & w47631;
assign w22777 = (~w21821 & w22775) | (~w21821 & w47632) | (w22775 & w47632);
assign w22778 = ~w22776 & ~w22777;
assign w22779 = w22758 & ~w22767;
assign w22780 = (w22486 & ~w22416) | (w22486 & w41968) | (~w22416 & w41968);
assign w22781 = ~w22453 & ~w22780;
assign w22782 = w22326 & w22753;
assign w22783 = w22586 & w22782;
assign w22784 = w22475 & w49007;
assign w22785 = w22522 & ~w22534;
assign w22786 = w22753 & ~w22785;
assign w22787 = w22586 & w22786;
assign w22788 = ~w22784 & ~w22787;
assign w22789 = w22781 & w22783;
assign w22790 = ~w22557 & ~w22608;
assign w22791 = w22602 & ~w22608;
assign w22792 = w22788 & w41969;
assign w22793 = ~w22790 & ~w22792;
assign w22794 = w4838 & w22758;
assign w22795 = ~w22759 & ~w22794;
assign w22796 = ~w22793 & ~w22795;
assign w22797 = w22793 & w22795;
assign w22798 = w22767 & w49008;
assign w22799 = ~w22779 & ~w22798;
assign w22800 = w15184 & ~w22799;
assign w22801 = ~w22740 & ~w22760;
assign w22802 = ~w22755 & ~w22759;
assign w22803 = (w22802 & ~w22619) | (w22802 & w50346) | (~w22619 & w50346);
assign w22804 = w4430 & ~w22767;
assign w22805 = ~w22803 & w22767;
assign w22806 = ~w22804 & ~w22805;
assign w22807 = w22801 & ~w22806;
assign w22808 = ~w22801 & w22806;
assign w22809 = ~w22807 & ~w22808;
assign w22810 = ~w22800 & w22809;
assign w22811 = w4056 & w4430;
assign w22812 = w4056 & ~w22779;
assign w22813 = ~w22798 & w22812;
assign w22814 = ~w22811 & ~w22813;
assign w22815 = ~w22810 & w22814;
assign w22816 = ~w22304 & w22475;
assign w22817 = ~w22781 & ~w22816;
assign w22818 = w22782 & w22785;
assign w22819 = ~w22817 & w22818;
assign w22820 = ~w22569 & ~w22589;
assign w22821 = ~w22786 & w22820;
assign w22822 = w22786 & ~w22820;
assign w22823 = ~w22817 & w49009;
assign w22824 = ~w22821 & ~w22822;
assign w22825 = ~w22819 & w22824;
assign w22826 = ~w22823 & ~w22825;
assign w22827 = w22568 & ~w22767;
assign w22828 = w22767 & w22826;
assign w22829 = ~w22827 & ~w22828;
assign w22830 = w6264 & ~w22568;
assign w22831 = w22830 & ~w22767;
assign w22832 = (w6264 & w22825) | (w6264 & w49010) | (w22825 & w49010);
assign w22833 = w22767 & w22832;
assign w22834 = ~w22831 & ~w22833;
assign w22835 = ~w22204 & w22765;
assign w22836 = ~w22477 & w22502;
assign w22837 = w22522 & w22750;
assign w22838 = w22836 & w22837;
assign w22839 = ~w7315 & w22750;
assign w22840 = w7315 & ~w22750;
assign w22841 = ~w22839 & ~w22840;
assign w22842 = ~w22838 & w22841;
assign w22843 = ~w22533 & ~w22842;
assign w22844 = ~w7315 & w22838;
assign w22845 = w22843 & ~w22844;
assign w22846 = w22207 & ~w22533;
assign w22847 = ~w22835 & w22846;
assign w22848 = ~w22845 & ~w22847;
assign w22849 = w22522 & w22836;
assign w22850 = w22839 & ~w22849;
assign w22851 = ~w22786 & ~w22819;
assign w22852 = ~w22850 & ~w22851;
assign w22853 = w6769 & w22207;
assign w22854 = ~w22835 & w22853;
assign w22855 = w6769 & ~w22852;
assign w22856 = ~w22854 & ~w22855;
assign w22857 = w22848 & ~w22856;
assign w22858 = w22834 & w22857;
assign w22859 = ~w6264 & ~w22829;
assign w22860 = ~w22858 & ~w22859;
assign w22861 = (w5745 & w22858) | (w5745 & w41970) | (w22858 & w41970);
assign w22862 = w22585 & w22599;
assign w22863 = ~w22819 & w22821;
assign w22864 = ~w22569 & ~w22863;
assign w22865 = w6264 & ~w22767;
assign w22866 = w22767 & ~w22864;
assign w22867 = ~w22865 & ~w22866;
assign w22868 = w22862 & ~w22867;
assign w22869 = ~w22862 & w22867;
assign w22870 = ~w22868 & ~w22869;
assign w22871 = ~w22861 & w22870;
assign w22872 = ~w21970 & ~w22546;
assign w22873 = ~w22202 & w49011;
assign w22874 = ~w22872 & ~w22873;
assign w22875 = w22788 & w41971;
assign w22876 = ~w22874 & ~w22875;
assign w22877 = ~w22766 & w22876;
assign w22878 = ~w22206 & w49012;
assign w22879 = ~w22835 & w22878;
assign w22880 = ~w22556 & ~w22608;
assign w22881 = ~w22877 & w47633;
assign w22882 = (w22880 & w22877) | (w22880 & w47634) | (w22877 & w47634);
assign w22883 = ~w22881 & ~w22882;
assign w22884 = ~w22546 & w22594;
assign w22885 = w22585 & ~w22884;
assign w22886 = ~w22207 & w22885;
assign w22887 = ~w22204 & ~w22745;
assign w22888 = w22764 & w22885;
assign w22889 = w22887 & w22888;
assign w22890 = w22599 & ~w22864;
assign w22891 = ~w22886 & ~w22889;
assign w22892 = ~w22890 & ~w22891;
assign w22893 = ~w22206 & w41972;
assign w22894 = ~w22765 & w22893;
assign w22895 = ~w22873 & w41973;
assign w22896 = ~w22894 & ~w22895;
assign w22897 = ~w22877 & w22896;
assign w22898 = ~w22892 & ~w22897;
assign w22899 = w4838 & ~w22880;
assign w22900 = (w22899 & w22877) | (w22899 & w47635) | (w22877 & w47635);
assign w22901 = w4838 & w22880;
assign w22902 = ~w22877 & w47636;
assign w22903 = ~w22900 & ~w22902;
assign w22904 = (w6027 & w22892) | (w6027 & w49013) | (w22892 & w49013);
assign w22905 = w22903 & ~w22904;
assign w22906 = ~w5330 & w22883;
assign w22907 = w22905 & ~w22906;
assign w22908 = ~w22892 & w49014;
assign w22909 = (~w22908 & ~w22905) | (~w22908 & w47637) | (~w22905 & w47637);
assign w22910 = w22871 & ~w22909;
assign w22911 = (w22485 & ~w22416) | (w22485 & w41974) | (~w22416 & w41974);
assign w22912 = w22416 & w22473;
assign w22913 = w22446 & ~w22911;
assign w22914 = w22416 & w41975;
assign w22915 = ~w22304 & w22914;
assign w22916 = ~w22913 & ~w22915;
assign w22917 = ~w22433 & w22451;
assign w22918 = w9195 & w22917;
assign w22919 = w22916 & w22918;
assign w22920 = w9195 & ~w22917;
assign w22921 = ~w22916 & w22920;
assign w22922 = ~w22919 & ~w22921;
assign w22923 = ~w22204 & w22922;
assign w22924 = w9195 & w22432;
assign w22925 = ~w22206 & w49015;
assign w22926 = ~w22835 & w22925;
assign w22927 = ~w22766 & w22923;
assign w22928 = ~w22926 & ~w22927;
assign w22929 = ~w22304 & w22912;
assign w22930 = w22416 & w45258;
assign w22931 = ~w22304 & w22930;
assign w22932 = w10419 & w52252;
assign w22933 = ~w22929 & w22932;
assign w22934 = (w22416 & w49016) | (w22416 & w49017) | (w49016 & w49017);
assign w22935 = ~w22931 & ~w22934;
assign w22936 = ~w22933 & w22935;
assign w22937 = ~w9781 & w22483;
assign w22938 = ~w22204 & w45259;
assign w22939 = ~w9781 & ~w22483;
assign w22940 = ~w21955 & w49018;
assign w22941 = (w22939 & ~w22935) | (w22939 & w41977) | (~w22935 & w41977);
assign w22942 = ~w22203 & w22940;
assign w22943 = ~w22941 & ~w22942;
assign w22944 = ~w22206 & w22940;
assign w22945 = ~w22765 & w22944;
assign w22946 = w22943 & ~w22945;
assign w22947 = ~w22766 & w22938;
assign w22948 = w22946 & ~w22947;
assign w22949 = ~w22928 & w22948;
assign w22950 = w22303 & w22497;
assign w22951 = ~w22273 & w22950;
assign w22952 = ~w22473 & w22497;
assign w22953 = (w22387 & w22473) | (w22387 & w49019) | (w22473 & w49019);
assign w22954 = ~w22366 & ~w22413;
assign w22955 = ~w22413 & w22953;
assign w22956 = (~w22954 & w22951) | (~w22954 & w49020) | (w22951 & w49020);
assign w22957 = ~w22397 & ~w22479;
assign w22958 = w10419 & w22957;
assign w22959 = ~w22956 & w22958;
assign w22960 = w10419 & ~w22957;
assign w22961 = w22956 & w22960;
assign w22962 = ~w22959 & ~w22961;
assign w22963 = ~w22204 & w22962;
assign w22964 = w10419 & w22396;
assign w22965 = ~w22206 & w49021;
assign w22966 = ~w22835 & w22965;
assign w22967 = ~w22766 & w22963;
assign w22968 = ~w22966 & ~w22967;
assign w22969 = w9781 & ~w22483;
assign w22970 = ~w22204 & w45260;
assign w22971 = w9781 & w22483;
assign w22972 = ~w21955 & w49022;
assign w22973 = (w22971 & ~w22935) | (w22971 & w41978) | (~w22935 & w41978);
assign w22974 = ~w22203 & w22972;
assign w22975 = ~w22973 & ~w22974;
assign w22976 = ~w22206 & w22972;
assign w22977 = ~w22765 & w22976;
assign w22978 = w22975 & ~w22977;
assign w22979 = ~w22766 & w22970;
assign w22980 = w22978 & ~w22979;
assign w22981 = ~w22968 & w22980;
assign w22982 = w22949 & ~w22981;
assign w22983 = w22916 & ~w22917;
assign w22984 = ~w22916 & w22917;
assign w22985 = ~w22983 & ~w22984;
assign w22986 = w22432 & ~w22767;
assign w22987 = ~w9195 & ~w22986;
assign w22988 = w22767 & w22985;
assign w22989 = w22987 & ~w22988;
assign w22990 = ~w22982 & ~w22989;
assign w22991 = ~w22507 & ~w22519;
assign w22992 = ~w22501 & w41979;
assign w22993 = ~w22477 & w22992;
assign w22994 = w7924 & ~w22993;
assign w22995 = ~w7924 & w22993;
assign w22996 = ~w22994 & ~w22995;
assign w22997 = ~w22204 & ~w22996;
assign w22998 = ~w7315 & ~w22515;
assign w22999 = (w22998 & w22766) | (w22998 & w41980) | (w22766 & w41980);
assign w23000 = ~w7315 & w22515;
assign w23001 = ~w22766 & w41981;
assign w23002 = ~w22999 & ~w23001;
assign w23003 = w22325 & ~w22519;
assign w23004 = ~w22506 & w23003;
assign w23005 = w22314 & ~w23003;
assign w23006 = ~w23004 & ~w23005;
assign w23007 = w22326 & ~w22519;
assign w23008 = (~w23006 & w22817) | (~w23006 & w49023) | (w22817 & w49023);
assign w23009 = ~w22506 & ~w23003;
assign w23010 = w22817 & w23009;
assign w23011 = w23008 & ~w23010;
assign w23012 = ~w7924 & w22518;
assign w23013 = w23012 & ~w22767;
assign w23014 = ~w7924 & w23011;
assign w23015 = w22767 & w23014;
assign w23016 = ~w23013 & ~w23015;
assign w23017 = w23002 & w23016;
assign w23018 = ~w9195 & w22817;
assign w23019 = w9195 & ~w22817;
assign w23020 = ~w23018 & ~w23019;
assign w23021 = ~w22204 & w23020;
assign w23022 = (w22505 & w22766) | (w22505 & w41982) | (w22766 & w41982);
assign w23023 = ~w22766 & w41983;
assign w23024 = ~w23022 & ~w23023;
assign w23025 = ~w8666 & w23024;
assign w23026 = w23017 & ~w23025;
assign w23027 = ~w22990 & w23026;
assign w23028 = w8666 & w22505;
assign w23029 = (w23028 & w22766) | (w23028 & w41984) | (w22766 & w41984);
assign w23030 = w8666 & ~w22505;
assign w23031 = ~w22766 & w41985;
assign w23032 = ~w23029 & ~w23031;
assign w23033 = w7924 & ~w22518;
assign w23034 = w23033 & ~w22767;
assign w23035 = w7924 & ~w23011;
assign w23036 = w22767 & w23035;
assign w23037 = ~w23034 & ~w23036;
assign w23038 = w23032 & w23037;
assign w23039 = w23017 & ~w23038;
assign w23040 = w22767 & w22852;
assign w23041 = w22848 & ~w23040;
assign w23042 = (~w6769 & ~w22848) | (~w6769 & w41986) | (~w22848 & w41986);
assign w23043 = w7315 & w22515;
assign w23044 = (w23043 & w22766) | (w23043 & w41987) | (w22766 & w41987);
assign w23045 = w7315 & ~w22515;
assign w23046 = ~w22766 & w41988;
assign w23047 = ~w23044 & ~w23046;
assign w23048 = w22834 & w23047;
assign w23049 = ~w23042 & w23048;
assign w23050 = ~w23039 & w23049;
assign w23051 = ~w23027 & w23050;
assign w23052 = ~w23027 & w41989;
assign w23053 = w5330 & w22898;
assign w23054 = (w22892 & w49024) | (w22892 & w49025) | (w49024 & w49025);
assign w23055 = w4430 & w22799;
assign w23056 = ~w22883 & ~w23054;
assign w23057 = ~w23055 & ~w23056;
assign w23058 = ~w22858 & w41990;
assign w23059 = w22907 & w23058;
assign w23060 = (w23057 & ~w23059) | (w23057 & w47638) | (~w23059 & w47638);
assign w23061 = w22910 & ~w23052;
assign w23062 = w23060 & ~w23061;
assign w23063 = ~w22273 & ~w22293;
assign w23064 = ~w16559 & w23063;
assign w23065 = w16559 & ~w23063;
assign w23066 = ~w23064 & ~w23065;
assign w23067 = w22764 & w23066;
assign w23068 = w22887 & w23067;
assign w23069 = ~w22207 & w23066;
assign w23070 = ~w23068 & ~w23069;
assign w23071 = ~w15681 & ~w22282;
assign w23072 = (w23071 & w23068) | (w23071 & w41991) | (w23068 & w41991);
assign w23073 = ~w23068 & w41992;
assign w23074 = ~w23072 & ~w23073;
assign w23075 = w15681 & w22282;
assign w23076 = (w23075 & w23068) | (w23075 & w41993) | (w23068 & w41993);
assign w23077 = w15681 & ~w22282;
assign w23078 = ~w23068 & w41994;
assign w23079 = ~w23076 & ~w23078;
assign w23080 = ~w22261 & ~w22271;
assign w23081 = ~w22270 & ~w22293;
assign w23082 = w23080 & ~w23081;
assign w23083 = ~w23080 & w23081;
assign w23084 = ~w23082 & ~w23083;
assign w23085 = ~w16559 & ~w22269;
assign w23086 = w23085 & ~w22767;
assign w23087 = ~w16559 & w23084;
assign w23088 = w23087 & w22767;
assign w23089 = ~w23086 & ~w23088;
assign w23090 = w23079 & ~w23089;
assign w23091 = ~a[28] & ~a[29];
assign w23092 = ~a[30] & w23091;
assign w23093 = w21801 & ~w23092;
assign w23094 = ~a[31] & ~w23093;
assign w23095 = w20906 & w23094;
assign w23096 = ~w22206 & w49026;
assign w23097 = ~w22835 & w23096;
assign w23098 = (w21952 & ~w21917) | (w21952 & w49027) | (~w21917 & w49027);
assign w23099 = (w21968 & w21921) | (w21968 & w49028) | (w21921 & w49028);
assign w23100 = ~w22205 & w23099;
assign w23101 = ~w21801 & w23091;
assign w23102 = ~a[30] & w23101;
assign w23103 = ~w22205 & w49029;
assign w23104 = ~w22765 & w23103;
assign w23105 = a[31] & w23093;
assign w23106 = ~w22208 & ~w23105;
assign w23107 = w20906 & w23106;
assign w23108 = w20906 & w23102;
assign w23109 = ~w23107 & ~w23108;
assign w23110 = (~w23109 & w22203) | (~w23109 & w49030) | (w22203 & w49030);
assign w23111 = ~w23104 & w23110;
assign w23112 = ~w23097 & ~w23111;
assign w23113 = ~a[32] & ~w21801;
assign w23114 = a[32] & w21801;
assign w23115 = ~w23113 & ~w23114;
assign w23116 = ~w20906 & ~w23102;
assign w23117 = ~w23094 & w23116;
assign w23118 = w23115 & ~w23117;
assign w23119 = a[32] & ~w22208;
assign w23120 = ~w22209 & ~w23119;
assign w23121 = ~w23106 & w23116;
assign w23122 = w23120 & ~w23121;
assign w23123 = (w23122 & w22203) | (w23122 & w49031) | (w22203 & w49031);
assign w23124 = (w23100 & w22745) | (w23100 & w41996) | (w22745 & w41996);
assign w23125 = w23123 & ~w23124;
assign w23126 = ~w22206 & w49032;
assign w23127 = ~w22835 & w23126;
assign w23128 = ~w23125 & ~w23127;
assign w23129 = w23112 & w23128;
assign w23130 = ~w20000 & ~w23129;
assign w23131 = ~w22211 & w22767;
assign w23132 = ~a[33] & w23113;
assign w23133 = a[33] & ~w23113;
assign w23134 = ~w23132 & ~w23133;
assign w23135 = ~w23131 & w23134;
assign w23136 = a[33] & ~w20906;
assign w23137 = ~a[33] & w20906;
assign w23138 = ~w23136 & ~w23137;
assign w23139 = ~w22208 & ~w23136;
assign w23140 = w23113 & ~w23139;
assign w23141 = w21801 & ~w22209;
assign w23142 = ~w23140 & ~w23141;
assign w23143 = w23138 & ~w23142;
assign w23144 = ~w23138 & w23142;
assign w23145 = ~w23143 & ~w23144;
assign w23146 = w22767 & ~w23145;
assign w23147 = ~w23135 & ~w23146;
assign w23148 = ~w23130 & w23147;
assign w23149 = w20000 & w23129;
assign w23150 = w22220 & ~w22233;
assign w23151 = (w22228 & w22766) | (w22228 & w41997) | (w22766 & w41997);
assign w23152 = ~w22766 & w41998;
assign w23153 = ~w23151 & ~w23152;
assign w23154 = w19040 & ~w23153;
assign w23155 = ~w23149 & ~w23154;
assign w23156 = ~w23148 & w23155;
assign w23157 = ~w19040 & w23153;
assign w23158 = ~w19040 & w22235;
assign w23159 = w19040 & ~w22235;
assign w23160 = ~w23158 & ~w23159;
assign w23161 = w22764 & ~w23160;
assign w23162 = w22887 & w23161;
assign w23163 = (~w23160 & w22206) | (~w23160 & w49033) | (w22206 & w49033);
assign w23164 = a[35] & ~w22242;
assign w23165 = ~a[35] & w22242;
assign w23166 = ~w23164 & ~w23165;
assign w23167 = ~w18183 & w23166;
assign w23168 = (w23167 & w23162) | (w23167 & w41999) | (w23162 & w41999);
assign w23169 = ~w18183 & ~w23166;
assign w23170 = ~w23162 & w42000;
assign w23171 = ~w23168 & ~w23170;
assign w23172 = w23074 & w23171;
assign w23173 = ~w23157 & w23172;
assign w23174 = ~w22247 & w22252;
assign w23175 = ~w18183 & w23174;
assign w23176 = w18183 & ~w23174;
assign w23177 = ~w23175 & ~w23176;
assign w23178 = w23177 & w22767;
assign w23179 = w17380 & w22258;
assign w23180 = ~w23178 & w23179;
assign w23181 = w17380 & ~w22258;
assign w23182 = w23178 & w23181;
assign w23183 = ~w23180 & ~w23182;
assign w23184 = ~w23090 & w23183;
assign w23185 = w23173 & w23184;
assign w23186 = ~w23156 & w23185;
assign w23187 = ~w23162 & w42001;
assign w23188 = (w23166 & w23162) | (w23166 & w42002) | (w23162 & w42002);
assign w23189 = ~w23187 & ~w23188;
assign w23190 = w18183 & w23189;
assign w23191 = ~w17380 & ~w22258;
assign w23192 = ~w23178 & w23191;
assign w23193 = ~w17380 & w22258;
assign w23194 = w23178 & w23193;
assign w23195 = ~w23192 & ~w23194;
assign w23196 = w16559 & w22269;
assign w23197 = w23196 & ~w22767;
assign w23198 = w16559 & ~w23084;
assign w23199 = w23198 & w22767;
assign w23200 = ~w23197 & ~w23199;
assign w23201 = w23079 & w23200;
assign w23202 = w23195 & w23201;
assign w23203 = w23183 & w23190;
assign w23204 = w23202 & ~w23203;
assign w23205 = w23074 & ~w23090;
assign w23206 = ~w23204 & w23205;
assign w23207 = ~w23186 & ~w23206;
assign w23208 = ~w22951 & w22953;
assign w23209 = w22365 & w22411;
assign w23210 = (w23209 & w22951) | (w23209 & w45261) | (w22951 & w45261);
assign w23211 = w11870 & ~w22411;
assign w23212 = ~w11870 & w22411;
assign w23213 = ~w23211 & ~w23212;
assign w23214 = w11870 & w23210;
assign w23215 = ~w23210 & ~w23213;
assign w23216 = ~w23214 & ~w23215;
assign w23217 = w20980 & ~w22340;
assign w23218 = ~w20980 & w22340;
assign w23219 = ~w23217 & ~w23218;
assign w23220 = ~w22766 & w42003;
assign w23221 = (w23219 & w22766) | (w23219 & w42004) | (w22766 & w42004);
assign w23222 = ~w23220 & ~w23221;
assign w23223 = w11138 & ~w23222;
assign w23224 = ~w11138 & w23222;
assign w23225 = w21801 & w22329;
assign w23226 = ~w21801 & w22360;
assign w23227 = ~w23225 & ~w23226;
assign w23228 = w21970 & ~w23227;
assign w23229 = ~w22206 & w23228;
assign w23230 = ~w22765 & w23229;
assign w23231 = w22356 & ~w23208;
assign w23232 = w12666 & ~w23231;
assign w23233 = ~w22203 & w23228;
assign w23234 = ~w23227 & ~w23232;
assign w23235 = ~w23233 & ~w23234;
assign w23236 = ~w12666 & w23231;
assign w23237 = ~w22204 & w23236;
assign w23238 = ~w22766 & w23237;
assign w23239 = ~w23230 & w23235;
assign w23240 = ~w23238 & ~w23239;
assign w23241 = ~w23232 & ~w23236;
assign w23242 = w23227 & ~w23241;
assign w23243 = w22767 & w23242;
assign w23244 = ~w23240 & ~w23243;
assign w23245 = (w11870 & w23240) | (w11870 & w42005) | (w23240 & w42005);
assign w23246 = ~w23224 & ~w23245;
assign w23247 = ~w21970 & ~w23208;
assign w23248 = ~w22202 & w49034;
assign w23249 = ~w23247 & ~w23248;
assign w23250 = w20997 & ~w22367;
assign w23251 = ~w20997 & w22367;
assign w23252 = ~w23250 & ~w23251;
assign w23253 = w21970 & w23252;
assign w23254 = ~w22203 & w23253;
assign w23255 = w22356 & ~w23254;
assign w23256 = w22765 & ~w23249;
assign w23257 = w23255 & ~w23256;
assign w23258 = ~w22206 & w23253;
assign w23259 = ~w22765 & w23258;
assign w23260 = ~w22207 & ~w23208;
assign w23261 = ~w23259 & ~w23260;
assign w23262 = w22386 & ~w22952;
assign w23263 = ~w22951 & w23262;
assign w23264 = ~w22356 & ~w23263;
assign w23265 = ~w22372 & ~w23263;
assign w23266 = (~w23265 & w22766) | (~w23265 & w42006) | (w22766 & w42006);
assign w23267 = w23257 & w23261;
assign w23268 = w23266 & ~w23267;
assign w23269 = ~w23267 & w42007;
assign w23270 = ~w23240 & w42008;
assign w23271 = ~w23269 & ~w23270;
assign w23272 = (~w23223 & w23271) | (~w23223 & w47639) | (w23271 & w47639);
assign w23273 = w22386 & w22491;
assign w23274 = w16559 & ~w22282;
assign w23275 = ~w22293 & ~w23274;
assign w23276 = (w23275 & w22261) | (w23275 & w45262) | (w22261 & w45262);
assign w23277 = ~w22454 & w22463;
assign w23278 = ~w23276 & w23277;
assign w23279 = w21125 & ~w22458;
assign w23280 = ~w21125 & w22458;
assign w23281 = ~w23279 & ~w23280;
assign w23282 = w15681 & w23281;
assign w23283 = ~w23278 & ~w23282;
assign w23284 = w22496 & w23283;
assign w23285 = w22470 & ~w23284;
assign w23286 = w23273 & ~w23285;
assign w23287 = ~w23273 & w23285;
assign w23288 = ~w23286 & ~w23287;
assign w23289 = ~w21115 & ~w22381;
assign w23290 = w21115 & w22381;
assign w23291 = ~w23289 & ~w23290;
assign w23292 = w22767 & w23288;
assign w23293 = ~w23291 & ~w22767;
assign w23294 = ~w23292 & ~w23293;
assign w23295 = (~w13384 & w23292) | (~w13384 & w47640) | (w23292 & w47640);
assign w23296 = (w12666 & w23267) | (w12666 & w42009) | (w23267 & w42009);
assign w23297 = ~w23295 & ~w23296;
assign w23298 = w23246 & w23297;
assign w23299 = ~w14766 & w23283;
assign w23300 = w14766 & ~w23283;
assign w23301 = ~w23299 & ~w23300;
assign w23302 = w21101 & ~w22465;
assign w23303 = ~w21101 & w22465;
assign w23304 = ~w23302 & ~w23303;
assign w23305 = ~w22766 & w42010;
assign w23306 = (~w23304 & w22766) | (~w23304 & w42011) | (w22766 & w42011);
assign w23307 = ~w23305 & ~w23306;
assign w23308 = ~w14039 & w23307;
assign w23309 = ~w23292 & w47641;
assign w23310 = ~w23308 & ~w23309;
assign w23311 = ~w22454 & ~w23276;
assign w23312 = ~w15681 & w23311;
assign w23313 = w15681 & ~w23311;
assign w23314 = ~w23312 & ~w23313;
assign w23315 = ~w23314 & w22767;
assign w23316 = w14039 & ~w23304;
assign w23317 = (w23316 & w22766) | (w23316 & w42012) | (w22766 & w42012);
assign w23318 = w14039 & w23304;
assign w23319 = ~w22766 & w42013;
assign w23320 = ~w23317 & ~w23319;
assign w23321 = ~w14766 & ~w23281;
assign w23322 = ~w23315 & w23321;
assign w23323 = w23320 & ~w23322;
assign w23324 = ~w14766 & w23281;
assign w23325 = w23315 & w23324;
assign w23326 = w23323 & ~w23325;
assign w23327 = w23310 & ~w23326;
assign w23328 = w23298 & ~w23327;
assign w23329 = w23272 & ~w23328;
assign w23330 = ~w23207 & ~w23329;
assign w23331 = (~w23281 & ~w22767) | (~w23281 & w45263) | (~w22767 & w45263);
assign w23332 = w22767 & w45264;
assign w23333 = ~w23331 & ~w23332;
assign w23334 = w14766 & w23320;
assign w23335 = w23333 & w23334;
assign w23336 = w23310 & ~w23335;
assign w23337 = w23298 & ~w23336;
assign w23338 = w23272 & ~w23337;
assign w23339 = w22956 & ~w22957;
assign w23340 = ~w22956 & w22957;
assign w23341 = ~w23339 & ~w23340;
assign w23342 = w22767 & ~w23341;
assign w23343 = ~w10419 & ~w23342;
assign w23344 = w22396 & ~w22767;
assign w23345 = w23343 & ~w23344;
assign w23346 = w22949 & ~w23345;
assign w23347 = (w23026 & ~w22990) | (w23026 & w45265) | (~w22990 & w45265);
assign w23348 = w23338 & w23347;
assign w23349 = ~w23330 & w23348;
assign w23350 = w23057 & ~w23059;
assign w23351 = ~w22910 & w23350;
assign w23352 = ~w22815 & ~w23062;
assign w23353 = (~w22815 & ~w23350) | (~w22815 & w47642) | (~w23350 & w47642);
assign w23354 = w23349 & w23353;
assign w23355 = ~w23352 & ~w23354;
assign w23356 = w5392 & ~w23058;
assign w23357 = ~w4056 & ~w22908;
assign w23358 = w22810 & ~w23357;
assign w23359 = ~w23356 & w23358;
assign w23360 = ~w23039 & w23047;
assign w23361 = ~w23027 & w23360;
assign w23362 = ~w5745 & w22829;
assign w23363 = ~w23042 & ~w23362;
assign w23364 = w6264 & ~w23363;
assign w23365 = w23042 & w23362;
assign w23366 = w5392 & ~w23365;
assign w23367 = ~w23364 & w23366;
assign w23368 = w23361 & w23367;
assign w23369 = (w23368 & w23330) | (w23368 & w42014) | (w23330 & w42014);
assign w23370 = w23359 & ~w23369;
assign w23371 = w23355 & ~w23370;
assign w23372 = (w23051 & w23330) | (w23051 & w42015) | (w23330 & w42015);
assign w23373 = w22647 & w22653;
assign w23374 = (~w23373 & w22203) | (~w23373 & w45266) | (w22203 & w45266);
assign w23375 = w22725 & ~w22742;
assign w23376 = w22619 & w42017;
assign w23377 = (w22742 & w22755) | (w22742 & w42018) | (w22755 & w42018);
assign w23378 = w22725 & ~w23377;
assign w23379 = ~w23377 & w45267;
assign w23380 = ~w23376 & w23379;
assign w23381 = (~w22638 & w23376) | (~w22638 & w45268) | (w23376 & w45268);
assign w23382 = w23374 & ~w23381;
assign w23383 = ~w22765 & w42019;
assign w23384 = w23382 & ~w23383;
assign w23385 = w22648 & w22653;
assign w23386 = ~w23380 & w23385;
assign w23387 = w22641 & ~w22642;
assign w23388 = ~w22641 & w22642;
assign w23389 = ~w23387 & ~w23388;
assign w23390 = w22767 & w23386;
assign w23391 = w23389 & ~w22767;
assign w23392 = ~w23390 & ~w23391;
assign w23393 = ~w23384 & w23392;
assign w23394 = (~w2006 & ~w23392) | (~w2006 & w45269) | (~w23392 & w45269);
assign w23395 = (w2006 & w22745) | (w2006 & w45270) | (w22745 & w45270);
assign w23396 = w22767 & ~w23395;
assign w23397 = ~w2006 & w22765;
assign w23398 = w23396 & ~w23397;
assign w23399 = ~w1738 & w22079;
assign w23400 = (w23399 & ~w23396) | (w23399 & w45271) | (~w23396 & w45271);
assign w23401 = ~w1738 & ~w22079;
assign w23402 = w23396 & w45272;
assign w23403 = ~w23400 & ~w23402;
assign w23404 = ~w23394 & w23403;
assign w23405 = w1738 & ~w22079;
assign w23406 = (w23405 & ~w23396) | (w23405 & w45273) | (~w23396 & w45273);
assign w23407 = w1738 & w22079;
assign w23408 = w23396 & w45274;
assign w23409 = ~w23406 & ~w23408;
assign w23410 = w22668 & ~w22688;
assign w23411 = w22723 & ~w22741;
assign w23412 = ~w22705 & ~w23411;
assign w23413 = (w22619 & w49035) | (w22619 & w49036) | (w49035 & w49036);
assign w23414 = (w22620 & w45275) | (w22620 & w45276) | (w45275 & w45276);
assign w23415 = w22685 & ~w23414;
assign w23416 = w2896 & ~w22767;
assign w23417 = w22767 & ~w23415;
assign w23418 = (w23410 & w23417) | (w23410 & w47643) | (w23417 & w47643);
assign w23419 = ~w23417 & w47644;
assign w23420 = ~w23418 & ~w23419;
assign w23421 = ~w22638 & ~w22726;
assign w23422 = ~w23376 & w45277;
assign w23423 = (w23421 & w23376) | (w23421 & w45278) | (w23376 & w45278);
assign w23424 = ~w23422 & ~w23423;
assign w23425 = w22637 & ~w22767;
assign w23426 = w22767 & ~w23424;
assign w23427 = ~w23425 & ~w23426;
assign w23428 = ~w2285 & ~w23427;
assign w23429 = w23420 & w45281;
assign w23430 = ~w23426 & w47645;
assign w23431 = (w2006 & w23383) | (w2006 & w45279) | (w23383 & w45279);
assign w23432 = w23392 & w23431;
assign w23433 = ~w23430 & ~w23432;
assign w23434 = ~w23404 & w23409;
assign w23435 = w23409 & w23433;
assign w23436 = ~w23429 & w23435;
assign w23437 = ~w23434 & ~w23436;
assign w23438 = w23396 & w45280;
assign w23439 = w23396 & ~w23438;
assign w23440 = ~w1738 & ~w22767;
assign w23441 = ~w23439 & ~w23440;
assign w23442 = ~w22135 & ~w22191;
assign w23443 = w1541 & w23442;
assign w23444 = ~w23441 & w23443;
assign w23445 = w1541 & ~w23442;
assign w23446 = w23441 & w23445;
assign w23447 = ~w23444 & ~w23446;
assign w23448 = ~w23437 & w23447;
assign w23449 = w2558 & ~w23420;
assign w23450 = (~w23428 & w23420) | (~w23428 & w45281) | (w23420 & w45281);
assign w23451 = ~w22206 & w49037;
assign w23452 = ~w22835 & w23451;
assign w23453 = ~w22204 & ~w23413;
assign w23454 = ~w22766 & w23453;
assign w23455 = ~w23452 & ~w23454;
assign w23456 = w22685 & w22695;
assign w23457 = ~w2896 & ~w23456;
assign w23458 = ~w23455 & w23457;
assign w23459 = ~w2896 & w23456;
assign w23460 = w23455 & w23459;
assign w23461 = ~w23458 & ~w23460;
assign w23462 = (w22762 & ~w22619) | (w22762 & w42021) | (~w22619 & w42021);
assign w23463 = ~w23462 & w22741;
assign w23464 = w22721 & ~w23463;
assign w23465 = ~w22705 & ~w22722;
assign w23466 = ~w23464 & ~w23465;
assign w23467 = (~w22705 & w22766) | (~w22705 & w42022) | (w22766 & w42022);
assign w23468 = ~w23466 & ~w23467;
assign w23469 = ~w22704 & ~w22767;
assign w23470 = ~w3242 & ~w23469;
assign w23471 = ~w23468 & w23470;
assign w23472 = w23461 & w23471;
assign w23473 = w23455 & ~w23456;
assign w23474 = ~w23455 & w23456;
assign w23475 = ~w23473 & ~w23474;
assign w23476 = w2896 & ~w23475;
assign w23477 = ~w23472 & ~w23476;
assign w23478 = w22721 & ~w22733;
assign w23479 = ~w23462 & w49038;
assign w23480 = (w23478 & w23462) | (w23478 & w49039) | (w23462 & w49039);
assign w23481 = ~w23479 & ~w23480;
assign w23482 = w22732 & ~w22767;
assign w23483 = w22767 & w23481;
assign w23484 = ~w23482 & ~w23483;
assign w23485 = (w3646 & w23483) | (w3646 & w49040) | (w23483 & w49040);
assign w23486 = w23461 & ~w23485;
assign w23487 = (~w23469 & w23467) | (~w23469 & w49041) | (w23467 & w49041);
assign w23488 = w3242 & ~w23487;
assign w23489 = w23486 & ~w23488;
assign w23490 = w23477 & ~w23489;
assign w23491 = ~w23490 & w42023;
assign w23492 = w23448 & ~w23491;
assign w23493 = ~w22814 & w22908;
assign w23494 = ~w5330 & w5745;
assign w23495 = w22860 & ~w23494;
assign w23496 = w23493 & w23495;
assign w23497 = ~w22892 & w49042;
assign w23498 = ~w22814 & w23497;
assign w23499 = ~w3646 & w23484;
assign w23500 = w23477 & w42025;
assign w23501 = w23491 & ~w23500;
assign w23502 = w23448 & ~w23501;
assign w23503 = (w23496 & ~w23448) | (w23496 & w47646) | (~w23448 & w47646);
assign w23504 = (w23502 & w23372) | (w23502 & w47647) | (w23372 & w47647);
assign w23505 = w23371 & w23504;
assign w23506 = w22156 & w22175;
assign w23507 = w22142 & ~w22198;
assign w23508 = w23507 & w50209;
assign w23509 = w1320 & ~w22767;
assign w23510 = w22767 & ~w23508;
assign w23511 = (w23506 & w23510) | (w23506 & w49043) | (w23510 & w49043);
assign w23512 = ~w23510 & w49044;
assign w23513 = ~w23511 & ~w23512;
assign w23514 = w1120 & ~w23513;
assign w23515 = w23441 & ~w23442;
assign w23516 = ~w23441 & w23442;
assign w23517 = ~w23515 & ~w23516;
assign w23518 = ~w1541 & w23517;
assign w23519 = w22133 & w22142;
assign w23520 = w22197 & w52253;
assign w23521 = w1541 & ~w22767;
assign w23522 = w22767 & w49045;
assign w23523 = ~w23521 & ~w23522;
assign w23524 = w23519 & ~w23523;
assign w23525 = ~w23519 & w23523;
assign w23526 = ~w23524 & ~w23525;
assign w23527 = ~w1320 & ~w23526;
assign w23528 = ~w23518 & ~w23527;
assign w23529 = ~w23492 & w23528;
assign w23530 = ~w23492 & w45282;
assign w23531 = w22031 & w22182;
assign w23532 = ~w22137 & w22199;
assign w23533 = ~w22730 & w45283;
assign w23534 = (w42028 & w22745) | (w42028 & w45284) | (w22745 & w45284);
assign w23535 = w23531 & ~w23534;
assign w23536 = w22175 & ~w23531;
assign w23537 = (w42029 & w22745) | (w42029 & w45285) | (w22745 & w45285);
assign w23538 = w1120 & w22182;
assign w23539 = w22031 & ~w23538;
assign w23540 = ~w22767 & w23539;
assign w23541 = w22767 & ~w23537;
assign w23542 = ~w23535 & w23541;
assign w23543 = (w945 & w23542) | (w945 & w45286) | (w23542 & w45286);
assign w23544 = (w42030 & w22745) | (w42030 & w45287) | (w22745 & w45287);
assign w23545 = w22031 & ~w23544;
assign w23546 = w754 & w22186;
assign w23547 = w945 & ~w22204;
assign w23548 = ~w22766 & w23547;
assign w23549 = ~w945 & ~w22204;
assign w23550 = ~w22766 & w23549;
assign w23551 = ~w22766 & w42031;
assign w23552 = ~w23545 & w23551;
assign w23553 = ~w22766 & w42032;
assign w23554 = w23545 & w23553;
assign w23555 = ~w23552 & ~w23554;
assign w23556 = w754 & ~w22186;
assign w23557 = (w23556 & w22766) | (w23556 & w42033) | (w22766 & w42033);
assign w23558 = w23545 & w23557;
assign w23559 = (w23556 & w22766) | (w23556 & w42034) | (w22766 & w42034);
assign w23560 = ~w23545 & w23559;
assign w23561 = ~w23558 & ~w23560;
assign w23562 = w23555 & w23561;
assign w23563 = w23543 & w23562;
assign w23564 = ~w754 & ~w22186;
assign w23565 = ~w22766 & w42035;
assign w23566 = ~w23545 & w23565;
assign w23567 = ~w22766 & w42036;
assign w23568 = w23545 & w23567;
assign w23569 = ~w23566 & ~w23568;
assign w23570 = ~w754 & w22186;
assign w23571 = (w23570 & w22766) | (w23570 & w42037) | (w22766 & w42037);
assign w23572 = w23545 & w23571;
assign w23573 = (w23570 & w22766) | (w23570 & w42038) | (w22766 & w42038);
assign w23574 = ~w23545 & w23573;
assign w23575 = ~w23572 & ~w23574;
assign w23576 = w23569 & w23575;
assign w23577 = w612 & w23576;
assign w23578 = ~w23563 & w23577;
assign w23579 = w945 & ~w23513;
assign w23580 = w23578 & ~w23579;
assign w23581 = ~w23542 & w49046;
assign w23582 = w493 & w23581;
assign w23583 = ~w23545 & w23548;
assign w23584 = w23545 & w23550;
assign w23585 = ~w23583 & ~w23584;
assign w23586 = w22186 & w23585;
assign w23587 = ~w22186 & ~w23585;
assign w23588 = ~w23586 & ~w23587;
assign w23589 = w23578 & w23588;
assign w23590 = ~w23582 & ~w23589;
assign w23591 = ~w1120 & ~w23590;
assign w23592 = ~w23580 & ~w23591;
assign w23593 = w23530 & ~w23592;
assign w23594 = w23359 & ~w23490;
assign w23595 = ~w5330 & ~w23058;
assign w23596 = w23493 & ~w23595;
assign w23597 = ~w23594 & ~w23596;
assign w23598 = w23349 & ~w23597;
assign w23599 = ~w23437 & w23500;
assign w23600 = ~w23051 & w23496;
assign w23601 = w23599 & ~w23600;
assign w23602 = ~w23368 & w23594;
assign w23603 = w23601 & ~w23602;
assign w23604 = ~w23598 & w23603;
assign w23605 = w23355 & w23604;
assign w23606 = w1320 & ~w23519;
assign w23607 = (w23606 & w23522) | (w23606 & w45288) | (w23522 & w45288);
assign w23608 = w1320 & w23519;
assign w23609 = ~w23522 & w45289;
assign w23610 = ~w23607 & ~w23609;
assign w23611 = w945 & w23610;
assign w23612 = w1320 & ~w23611;
assign w23613 = w945 & ~w1541;
assign w23614 = w23526 & ~w23613;
assign w23615 = ~w23518 & w23612;
assign w23616 = ~w23517 & w23614;
assign w23617 = ~w23615 & ~w23616;
assign w23618 = ~w23437 & ~w23491;
assign w23619 = ~w1120 & w23581;
assign w23620 = ~w23618 & w23619;
assign w23621 = ~w23617 & w23620;
assign w23622 = ~w23605 & w23621;
assign w23623 = ~w23527 & ~w23611;
assign w23624 = ~w23447 & w23623;
assign w23625 = w23619 & w23624;
assign w23626 = ~w23542 & w49047;
assign w23627 = w23562 & ~w23626;
assign w23628 = ~w1120 & w23513;
assign w23629 = w23610 & ~w23628;
assign w23630 = ~w23514 & ~w23629;
assign w23631 = ~w945 & w23582;
assign w23632 = (~w23631 & ~w23630) | (~w23631 & w47648) | (~w23630 & w47648);
assign w23633 = w23589 & ~w23627;
assign w23634 = w23632 & ~w23633;
assign w23635 = ~w23625 & w23634;
assign w23636 = w23591 & ~w23610;
assign w23637 = w23635 & ~w23636;
assign w23638 = (w23637 & w23605) | (w23637 & w42039) | (w23605 & w42039);
assign w23639 = (w23593 & ~w23371) | (w23593 & w42040) | (~w23371 & w42040);
assign w23640 = w23638 & ~w23639;
assign w23641 = ~w21818 & w22773;
assign w23642 = ~w22772 & w23641;
assign w23643 = (w21931 & w22772) | (w21931 & w49048) | (w22772 & w49048);
assign w23644 = w21903 & w22767;
assign w23645 = (~w21820 & w22772) | (~w21820 & w47649) | (w22772 & w47649);
assign w23646 = w21903 & w21930;
assign w23647 = w21897 & ~w21898;
assign w23648 = ~w21897 & w21898;
assign w23649 = ~w23647 & ~w23648;
assign w23650 = w23649 & ~w22767;
assign w23651 = (w41967 & w47650) | (w41967 & w47651) | (w47650 & w47651);
assign w23652 = ~w23645 & w23651;
assign w23653 = ~w23650 & ~w23652;
assign w23654 = w23643 & w23644;
assign w23655 = w23653 & ~w23654;
assign w23656 = ~w80 & w23655;
assign w23657 = w57 & w22778;
assign w23658 = ~w23656 & ~w23657;
assign w23659 = ~w23643 & w23644;
assign w23660 = (w21915 & w21916) | (w21915 & ~w22767) | (w21916 & ~w22767);
assign w23661 = w45290 & w22767;
assign w23662 = ~w23660 & ~w23661;
assign w23663 = w23659 & ~w23662;
assign w23664 = ~w23659 & w23662;
assign w23665 = ~w23663 & ~w23664;
assign w23666 = w22778 & w23655;
assign w23667 = (w3 & w23666) | (w3 & w49049) | (w23666 & w49049);
assign w23668 = w23658 & ~w23667;
assign w23669 = (~w22745 & w45291) | (~w22745 & w45292) | (w45291 & w45292);
assign w23670 = ~w22064 & w23669;
assign w23671 = ~w21856 & w22767;
assign w23672 = (w21891 & ~w23669) | (w21891 & w49050) | (~w23669 & w49050);
assign w23673 = w23671 & ~w23672;
assign w23674 = ~w21866 & ~w21918;
assign w23675 = w21865 & ~w22767;
assign w23676 = w23674 & w22767;
assign w23677 = ~w23675 & ~w23676;
assign w23678 = w23673 & w23674;
assign w23679 = ~w23673 & w23677;
assign w23680 = ~w23678 & ~w23679;
assign w23681 = ~w252 & ~w23680;
assign w23682 = ~w57 & ~w22778;
assign w23683 = ~w23681 & ~w23682;
assign w23684 = w23668 & ~w23683;
assign w23685 = w22183 & ~w22187;
assign w23686 = (w42041 & w22745) | (w42041 & w45293) | (w22745 & w45293);
assign w23687 = ~w22040 & ~w22057;
assign w23688 = ~w23686 & w23687;
assign w23689 = ~w21984 & ~w22041;
assign w23690 = ~w21983 & ~w22767;
assign w23691 = (w41967 & w47652) | (w41967 & w47653) | (w47652 & w47653);
assign w23692 = ~w23688 & w23691;
assign w23693 = (w41967 & w47654) | (w41967 & w47655) | (w47654 & w47655);
assign w23694 = w23688 & w23693;
assign w23695 = ~w23692 & ~w23694;
assign w23696 = ~w23690 & w23695;
assign w23697 = w23576 & ~w23696;
assign w23698 = ~w23563 & w23697;
assign w23699 = ~w23578 & ~w23698;
assign w23700 = w21890 & ~w22064;
assign w23701 = (~w41967 & w47656) | (~w41967 & w47657) | (w47656 & w47657);
assign w23702 = w22767 & ~w23669;
assign w23703 = (w23700 & w23702) | (w23700 & w47658) | (w23702 & w47658);
assign w23704 = ~w23702 & w47659;
assign w23705 = ~w23703 & ~w23704;
assign w23706 = w22059 & ~w23686;
assign w23707 = ~w21984 & w22767;
assign w23708 = ~w23706 & w23707;
assign w23709 = w612 & ~w22767;
assign w23710 = ~w23708 & ~w23709;
assign w23711 = ~w22000 & ~w22066;
assign w23712 = ~w19000 & ~w23711;
assign w23713 = ~w23708 & w45294;
assign w23714 = ~w19000 & w23711;
assign w23715 = (w23714 & w23708) | (w23714 & w45295) | (w23708 & w45295);
assign w23716 = ~w23713 & ~w23715;
assign w23717 = w400 & ~w23705;
assign w23718 = w23716 & ~w23717;
assign w23719 = ~w23699 & w23718;
assign w23720 = ~w23627 & w23718;
assign w23721 = ~w23699 & w23720;
assign w23722 = ~w21856 & ~w21868;
assign w23723 = ~w400 & ~w22767;
assign w23724 = w21890 & w22767;
assign w23725 = ~w23670 & w23724;
assign w23726 = ~w23723 & ~w23725;
assign w23727 = w23722 & ~w23726;
assign w23728 = ~w23722 & w23726;
assign w23729 = ~w23727 & ~w23728;
assign w23730 = w351 & w23729;
assign w23731 = (w612 & ~w23695) | (w612 & w45296) | (~w23695 & w45296);
assign w23732 = w493 & ~w23711;
assign w23733 = (w23732 & w23708) | (w23732 & w45297) | (w23708 & w45297);
assign w23734 = w493 & w23711;
assign w23735 = ~w23708 & w45298;
assign w23736 = ~w23733 & ~w23735;
assign w23737 = ~w23731 & w23736;
assign w23738 = w23718 & ~w23737;
assign w23739 = ~w23730 & ~w23738;
assign w23740 = ~w23721 & w23739;
assign w23741 = ~w18997 & w23705;
assign w23742 = w23740 & ~w23741;
assign w23743 = w23630 & w23719;
assign w23744 = w23742 & ~w23743;
assign w23745 = w23742 & w49051;
assign w23746 = w23698 & w23741;
assign w23747 = (w23695 & w32606) | (w23695 & w49052) | (w32606 & w49052);
assign w23748 = w23741 & ~w23747;
assign w23749 = ~w23746 & ~w23748;
assign w23750 = ~w23719 & w23749;
assign w23751 = w23739 & w23750;
assign w23752 = w23530 & ~w23751;
assign w23753 = (w23752 & ~w23371) | (w23752 & w42042) | (~w23371 & w42042);
assign w23754 = w23745 & ~w23753;
assign w23755 = (~w23748 & w23629) | (~w23748 & w47660) | (w23629 & w47660);
assign w23756 = w23698 & w45299;
assign w23757 = w23755 & ~w23756;
assign w23758 = w23683 & w23740;
assign w23759 = w23757 & w23758;
assign w23760 = w23371 & w42043;
assign w23761 = ~w23530 & w23759;
assign w23762 = ~w23684 & w23751;
assign w23763 = ~w23761 & ~w23762;
assign w23764 = ~w23760 & w23763;
assign w23765 = ~w23754 & w23764;
assign w23766 = w23640 & ~w23765;
assign w23767 = w252 & w23680;
assign w23768 = ~w351 & ~w23729;
assign w23769 = ~w23767 & ~w23768;
assign w23770 = w23668 & w23769;
assign w23771 = ~w23684 & ~w23770;
assign w23772 = ~w21946 & ~w21957;
assign w23773 = (w21917 & w23642) | (w21917 & w21932) | (w23642 & w21932);
assign w23774 = w21951 & ~w23773;
assign w23775 = w3 & ~w22767;
assign w23776 = w22767 & w23774;
assign w23777 = ~w23775 & ~w23776;
assign w23778 = w21952 & ~w23773;
assign w23779 = ~w21957 & ~w23778;
assign w23780 = ~w21829 & w21830;
assign w23781 = w21623 & ~w23780;
assign w23782 = w21636 & ~w21829;
assign w23783 = ~w21848 & ~w23782;
assign w23784 = w21848 & ~w21957;
assign w23785 = ~w23778 & w23784;
assign w23786 = ~w42 & ~w23785;
assign w23787 = ~w23781 & w23783;
assign w23788 = ~w23779 & w23787;
assign w23789 = w23786 & ~w23788;
assign w23790 = w42 & w23772;
assign w23791 = ~w23777 & w23790;
assign w23792 = w42 & ~w23772;
assign w23793 = w23777 & w23792;
assign w23794 = ~w23789 & ~w23793;
assign w23795 = ~w23791 & w23794;
assign w23796 = ~w21848 & ~w21946;
assign w23797 = w42 & ~w23796;
assign w23798 = w22767 & w23797;
assign w23799 = ~w23785 & w23798;
assign w23800 = w23774 & ~w23784;
assign w23801 = w23799 & ~w23800;
assign w23802 = ~w23795 & ~w23801;
assign w23803 = ~w23771 & w23802;
assign w23804 = ~w23761 & w45300;
assign w23805 = ~w23760 & w23804;
assign w23806 = ~w23745 & w23803;
assign w23807 = (~w23806 & w23760) | (~w23806 & w45301) | (w23760 & w45301);
assign w23808 = (~w23807 & w23765) | (~w23807 & w45302) | (w23765 & w45302);
assign w23809 = w3 & ~w80;
assign w23810 = ~w23665 & ~w23809;
assign w23811 = w536 & ~w23655;
assign w23812 = ~w23810 & ~w23811;
assign w23813 = w376 & ~w23680;
assign w23814 = w3 & w23655;
assign w23815 = ~w23813 & w23814;
assign w23816 = ~w23812 & ~w23815;
assign w23817 = ~w42 & ~w23772;
assign w23818 = w23777 & w23817;
assign w23819 = ~w42 & w23772;
assign w23820 = ~w23777 & w23819;
assign w23821 = ~w23818 & ~w23820;
assign w23822 = ~w23816 & w23821;
assign w23823 = w22767 & w23643;
assign w23824 = ~w57 & ~w21951;
assign w23825 = ~w23823 & w23824;
assign w23826 = ~w23768 & w47661;
assign w23827 = w23822 & ~w23826;
assign w23828 = w23802 & ~w23827;
assign w23829 = ~w23827 & w47662;
assign w23830 = ~w23750 & ~w23757;
assign w23831 = w23740 & w23822;
assign w23832 = ~w23830 & w23831;
assign w23833 = w23828 & ~w23832;
assign w23834 = ~w23829 & ~w23833;
assign w23835 = w23637 & ~w23833;
assign w23836 = (~w23834 & w23622) | (~w23834 & w42044) | (w23622 & w42044);
assign w23837 = ~w23492 & w49053;
assign w23838 = w23593 & w23829;
assign w23839 = w23828 & w23837;
assign w23840 = ~w23838 & ~w23839;
assign w23841 = ~w23505 & ~w23840;
assign w23842 = ~w23836 & ~w23841;
assign w23843 = ~w23808 & w23842;
assign w23844 = (w23837 & ~w23371) | (w23837 & w42045) | (~w23371 & w42045);
assign w23845 = w23740 & ~w23830;
assign w23846 = ~w23681 & w23845;
assign w23847 = ~w23844 & w23846;
assign w23848 = w23640 & w23847;
assign w23849 = w23530 & w23719;
assign w23850 = ~w23681 & ~w23769;
assign w23851 = w23849 & ~w23850;
assign w23852 = ~w23744 & w23769;
assign w23853 = ~w23681 & ~w23852;
assign w23854 = (w23853 & w23505) | (w23853 & w42046) | (w23505 & w42046);
assign w23855 = ~w23848 & ~w23854;
assign w23856 = ~w23657 & ~w23682;
assign w23857 = ~w23855 & ~w23856;
assign w23858 = w23855 & w23856;
assign w23859 = ~w22778 & ~w23843;
assign w23860 = ~w23857 & ~w23858;
assign w23861 = w23843 & w23860;
assign w23862 = ~w23859 & ~w23861;
assign w23863 = w80 & ~w23862;
assign w23864 = ~w23330 & w23338;
assign w23865 = ~w22968 & ~w23864;
assign w23866 = ~w23345 & ~w23865;
assign w23867 = w22948 & w23866;
assign w23868 = w22980 & ~w23867;
assign w23869 = ~w9195 & ~w23842;
assign w23870 = ~w9195 & ~w23807;
assign w23871 = ~w23766 & w23870;
assign w23872 = ~w23869 & ~w23871;
assign w23873 = w23842 & ~w23868;
assign w23874 = ~w23808 & w23873;
assign w23875 = w23872 & ~w23874;
assign w23876 = ~w22928 & ~w22989;
assign w23877 = ~w8666 & ~w23876;
assign w23878 = w23872 & w45303;
assign w23879 = ~w8666 & w23876;
assign w23880 = (w23879 & ~w23872) | (w23879 & w45304) | (~w23872 & w45304);
assign w23881 = ~w23878 & ~w23880;
assign w23882 = w8666 & ~w23876;
assign w23883 = (w23882 & ~w23872) | (w23882 & w45305) | (~w23872 & w45305);
assign w23884 = w8666 & w23876;
assign w23885 = w23872 & w45306;
assign w23886 = ~w23883 & ~w23885;
assign w23887 = ~w9781 & ~w23842;
assign w23888 = ~w9781 & ~w23807;
assign w23889 = ~w23766 & w23888;
assign w23890 = ~w23887 & ~w23889;
assign w23891 = w23842 & ~w23866;
assign w23892 = ~w23808 & w23891;
assign w23893 = w22948 & w22980;
assign w23894 = ~w9195 & w23893;
assign w23895 = (w23894 & ~w23890) | (w23894 & w45307) | (~w23890 & w45307);
assign w23896 = ~w9195 & ~w23893;
assign w23897 = w23890 & w45308;
assign w23898 = ~w23895 & ~w23897;
assign w23899 = w23886 & w23898;
assign w23900 = w23881 & ~w23899;
assign w23901 = (w14766 & w23186) | (w14766 & w45309) | (w23186 & w45309);
assign w23902 = ~w23186 & w42047;
assign w23903 = (w23333 & w23186) | (w23333 & w45310) | (w23186 & w45310);
assign w23904 = ~w23901 & ~w23903;
assign w23905 = w23320 & ~w23904;
assign w23906 = (w23310 & w23904) | (w23310 & w47663) | (w23904 & w47663);
assign w23907 = w23297 & ~w23906;
assign w23908 = ~w23269 & ~w23907;
assign w23909 = ~w11870 & w23908;
assign w23910 = w23842 & w23909;
assign w23911 = ~w23808 & w23910;
assign w23912 = w23750 & w23758;
assign w23913 = ~w23761 & w47664;
assign w23914 = ~w23760 & w23913;
assign w23915 = w23741 & w23803;
assign w23916 = ~w23640 & w23915;
assign w23917 = ~w23914 & ~w23916;
assign w23918 = w11870 & ~w23908;
assign w23919 = w23842 & w23918;
assign w23920 = w23917 & w23919;
assign w23921 = w11138 & w23244;
assign w23922 = ~w23920 & w23921;
assign w23923 = ~w23911 & w23922;
assign w23924 = ~w23909 & ~w23918;
assign w23925 = w23842 & w45311;
assign w23926 = ~w23808 & w23925;
assign w23927 = w11138 & w23926;
assign w23928 = ~w23923 & ~w23927;
assign w23929 = ~w23223 & ~w23224;
assign w23930 = w23271 & ~w23907;
assign w23931 = ~w23245 & ~w23930;
assign w23932 = w23929 & ~w23931;
assign w23933 = ~w23929 & w23931;
assign w23934 = ~w23932 & ~w23933;
assign w23935 = ~w23222 & ~w23842;
assign w23936 = ~w23222 & ~w23807;
assign w23937 = ~w23766 & w23936;
assign w23938 = ~w23935 & ~w23937;
assign w23939 = w23842 & ~w23934;
assign w23940 = ~w23808 & w23939;
assign w23941 = w23938 & ~w23940;
assign w23942 = (~w10419 & ~w23938) | (~w10419 & w45312) | (~w23938 & w45312);
assign w23943 = w23928 & ~w23942;
assign w23944 = w23244 & ~w23920;
assign w23945 = ~w23911 & w23944;
assign w23946 = ~w11138 & ~w23926;
assign w23947 = ~w23945 & w23946;
assign w23948 = ~w23295 & ~w23906;
assign w23949 = w12666 & ~w23948;
assign w23950 = ~w12666 & w23948;
assign w23951 = ~w23949 & ~w23950;
assign w23952 = w23842 & w23951;
assign w23953 = ~w23808 & w23952;
assign w23954 = w11870 & ~w23268;
assign w23955 = ~w23953 & w23954;
assign w23956 = w11870 & w23268;
assign w23957 = w23953 & w23956;
assign w23958 = ~w23955 & ~w23957;
assign w23959 = ~w23947 & w23958;
assign w23960 = w10419 & w23941;
assign w23961 = w10419 & ~w23842;
assign w23962 = w10419 & ~w23807;
assign w23963 = ~w23766 & w23962;
assign w23964 = ~w23961 & ~w23963;
assign w23965 = w23842 & w23864;
assign w23966 = ~w23808 & w23965;
assign w23967 = w23964 & ~w23966;
assign w23968 = ~w22968 & ~w23345;
assign w23969 = w9781 & ~w23968;
assign w23970 = (w23969 & ~w23964) | (w23969 & w45313) | (~w23964 & w45313);
assign w23971 = w9781 & w23968;
assign w23972 = w23964 & w45314;
assign w23973 = ~w23970 & ~w23972;
assign w23974 = ~w23960 & w23973;
assign w23975 = w23943 & ~w23959;
assign w23976 = w23974 & ~w23975;
assign w23977 = ~w23900 & w23976;
assign w23978 = w14039 & ~w23904;
assign w23979 = ~w14039 & w23904;
assign w23980 = ~w23978 & ~w23979;
assign w23981 = w23842 & ~w23980;
assign w23982 = w23917 & w23981;
assign w23983 = w23307 & ~w23982;
assign w23984 = w23842 & w45315;
assign w23985 = ~w23808 & w23984;
assign w23986 = ~w23983 & ~w23985;
assign w23987 = ~w23983 & w45316;
assign w23988 = (w13384 & w23983) | (w13384 & w45317) | (w23983 & w45317);
assign w23989 = ~w23987 & ~w23988;
assign w23990 = ~w23901 & ~w23902;
assign w23991 = w23917 & w45318;
assign w23992 = ~w23333 & w23990;
assign w23993 = ~w23808 & w47665;
assign w23994 = w23333 & ~w23991;
assign w23995 = ~w23993 & ~w23994;
assign w23996 = (~w14039 & w23994) | (~w14039 & w47666) | (w23994 & w47666);
assign w23997 = w23989 & ~w23996;
assign w23998 = ~w23308 & ~w23905;
assign w23999 = ~w13384 & w23998;
assign w24000 = w13384 & ~w23998;
assign w24001 = ~w23999 & ~w24000;
assign w24002 = w23842 & w24001;
assign w24003 = ~w23640 & w23741;
assign w24004 = (~w23294 & ~w24002) | (~w23294 & w45320) | (~w24002 & w45320);
assign w24005 = ~w23294 & w50210;
assign w24006 = w23808 & w24005;
assign w24007 = ~w24004 & ~w24006;
assign w24008 = w23842 & w47667;
assign w24009 = ~w23808 & w24008;
assign w24010 = w24007 & ~w24009;
assign w24011 = (w12666 & ~w24007) | (w12666 & w47668) | (~w24007 & w47668);
assign w24012 = ~w23987 & ~w24011;
assign w24013 = ~w23997 & w24012;
assign w24014 = w23268 & ~w23953;
assign w24015 = ~w23268 & w23953;
assign w24016 = ~w24014 & ~w24015;
assign w24017 = ~w11870 & ~w24016;
assign w24018 = w24007 & w47669;
assign w24019 = ~w24017 & ~w24018;
assign w24020 = w23943 & w24019;
assign w24021 = ~w24013 & w24020;
assign w24022 = w23977 & ~w24021;
assign w24023 = w23890 & w45321;
assign w24024 = (w23893 & ~w23890) | (w23893 & w45322) | (~w23890 & w45322);
assign w24025 = ~w24023 & ~w24024;
assign w24026 = w9195 & w24025;
assign w24027 = ~w9781 & ~w23968;
assign w24028 = w23964 & w45323;
assign w24029 = ~w9781 & w23968;
assign w24030 = (w24029 & ~w23964) | (w24029 & w45324) | (~w23964 & w45324);
assign w24031 = ~w24028 & ~w24030;
assign w24032 = w23881 & w24031;
assign w24033 = ~w24026 & w24032;
assign w24034 = ~w23900 & ~w24033;
assign w24035 = (~w24034 & ~w23977) | (~w24034 & w45325) | (~w23977 & w45325);
assign w24036 = w14039 & w23995;
assign w24037 = ~w23988 & w24036;
assign w24038 = w24012 & ~w24037;
assign w24039 = w24020 & ~w24038;
assign w24040 = w23977 & ~w24039;
assign w24041 = w21801 & w22767;
assign w24042 = ~w21801 & ~w22767;
assign w24043 = ~w24041 & ~w24042;
assign w24044 = w23842 & ~w24043;
assign w24045 = ~w23808 & w24044;
assign w24046 = a[30] & ~w24045;
assign w24047 = ~w22767 & ~w23842;
assign w24048 = ~w22767 & ~w23807;
assign w24049 = ~w23766 & w24048;
assign w24050 = ~w24047 & ~w24049;
assign w24051 = ~w23092 & ~w24043;
assign w24052 = w23091 & ~w24041;
assign w24053 = ~w24051 & ~w24052;
assign w24054 = w23842 & w24053;
assign w24055 = w23917 & w24054;
assign w24056 = w21801 & ~w23091;
assign w24057 = ~w23102 & ~w24056;
assign w24058 = ~w22767 & ~w24057;
assign w24059 = a[31] & ~w24058;
assign w24060 = ~w24055 & w24059;
assign w24061 = w24050 & w24060;
assign w24062 = ~a[30] & w22767;
assign w24063 = (w24062 & ~w23917) | (w24062 & w45326) | (~w23917 & w45326);
assign w24064 = ~a[31] & ~w24063;
assign w24065 = ~w23753 & w23845;
assign w24066 = w21801 & w23091;
assign w24067 = ~w22767 & w24066;
assign w24068 = ~w23684 & w24067;
assign w24069 = ~w23753 & w45327;
assign w24070 = ~w23101 & ~w24056;
assign w24071 = w22767 & ~w24070;
assign w24072 = ~w23803 & w24067;
assign w24073 = ~w24071 & ~w24072;
assign w24074 = (w24073 & w24003) | (w24073 & w45328) | (w24003 & w45328);
assign w24075 = w24051 & ~w24062;
assign w24076 = w23842 & w24075;
assign w24077 = ~w23808 & w24076;
assign w24078 = ~a[30] & w23842;
assign w24079 = ~w24074 & w24078;
assign w24080 = ~w24077 & ~w24079;
assign w24081 = ~w24046 & w24061;
assign w24082 = w24064 & w24080;
assign w24083 = ~w24081 & ~w24082;
assign w24084 = w23640 & w24065;
assign w24085 = ~w23816 & w24084;
assign w24086 = ~w23684 & w23821;
assign w24087 = w23770 & ~w23845;
assign w24088 = w24086 & ~w24087;
assign w24089 = (w24088 & ~w23753) | (w24088 & w45329) | (~w23753 & w45329);
assign w24090 = (w23849 & ~w23371) | (w23849 & w42048) | (~w23371 & w42048);
assign w24091 = ~w23816 & ~w23826;
assign w24092 = w23744 & ~w23816;
assign w24093 = (~w24091 & w24090) | (~w24091 & w45330) | (w24090 & w45330);
assign w24094 = w24089 & ~w24093;
assign w24095 = w23802 & ~w24094;
assign w24096 = ~w23640 & ~w23754;
assign w24097 = w23803 & w24096;
assign w24098 = ~w24095 & ~w24097;
assign w24099 = w24085 & w24089;
assign w24100 = ~w24098 & ~w24099;
assign w24101 = ~a[26] & ~a[27];
assign w24102 = ~a[28] & w24101;
assign w24103 = w22767 & w24102;
assign w24104 = ~w22767 & ~w24102;
assign w24105 = a[29] & w24104;
assign w24106 = ~w23091 & ~w24105;
assign w24107 = ~w24103 & ~w24106;
assign w24108 = a[30] & ~w23091;
assign w24109 = ~w23092 & ~w24108;
assign w24110 = w21801 & w24107;
assign w24111 = w24109 & ~w24110;
assign w24112 = ~w21801 & ~w24107;
assign w24113 = ~w24111 & ~w24112;
assign w24114 = a[30] & ~w22767;
assign w24115 = ~w24062 & ~w24114;
assign w24116 = ~a[29] & ~w24104;
assign w24117 = ~w24103 & ~w24116;
assign w24118 = ~w21801 & w24115;
assign w24119 = w24117 & ~w24118;
assign w24120 = w21801 & ~w24115;
assign w24121 = ~w24119 & ~w24120;
assign w24122 = w20906 & ~w24113;
assign w24123 = ~w24100 & w24122;
assign w24124 = w20906 & w24121;
assign w24125 = w24100 & w24124;
assign w24126 = ~w24123 & ~w24125;
assign w24127 = w24083 & w24126;
assign w24128 = ~w22204 & w23106;
assign w24129 = ~w23104 & w24128;
assign w24130 = w23116 & ~w24129;
assign w24131 = ~w22767 & w23094;
assign w24132 = w24130 & ~w24131;
assign w24133 = w23112 & ~w24132;
assign w24134 = w23842 & w24133;
assign w24135 = w23917 & w24134;
assign w24136 = ~w22767 & w23115;
assign w24137 = w22767 & w23120;
assign w24138 = ~w24136 & ~w24137;
assign w24139 = ~w24135 & w24138;
assign w24140 = w23842 & w45331;
assign w24141 = ~w23808 & w24140;
assign w24142 = ~w24139 & ~w24141;
assign w24143 = w20000 & ~w24142;
assign w24144 = ~w20906 & ~w24121;
assign w24145 = w24100 & w24144;
assign w24146 = ~w20906 & w24113;
assign w24147 = ~w24100 & w24146;
assign w24148 = ~w24145 & ~w24147;
assign w24149 = ~w24143 & w24148;
assign w24150 = ~w24127 & w24149;
assign w24151 = ~w24139 & w45332;
assign w24152 = ~w23130 & ~w23149;
assign w24153 = w23842 & w24152;
assign w24154 = w23917 & w24153;
assign w24155 = ~w23147 & ~w24154;
assign w24156 = w23842 & w45333;
assign w24157 = ~w23808 & w24156;
assign w24158 = ~w24155 & ~w24157;
assign w24159 = (~w19040 & w24155) | (~w19040 & w45334) | (w24155 & w45334);
assign w24160 = ~w24151 & ~w24159;
assign w24161 = w19040 & w23147;
assign w24162 = ~w23842 & w24161;
assign w24163 = ~w24160 & ~w24162;
assign w24164 = ~w23147 & ~w23149;
assign w24165 = w19040 & ~w23130;
assign w24166 = ~w19040 & ~w23149;
assign w24167 = ~w23148 & w24166;
assign w24168 = ~w24164 & w24165;
assign w24169 = ~w24167 & ~w24168;
assign w24170 = w23842 & w45335;
assign w24171 = ~w23808 & w24170;
assign w24172 = ~w23153 & ~w24171;
assign w24173 = (w23153 & ~w23842) | (w23153 & w45336) | (~w23842 & w45336);
assign w24174 = ~w23808 & ~w24170;
assign w24175 = ~w24173 & w24174;
assign w24176 = ~w24172 & ~w24175;
assign w24177 = ~w18183 & w24176;
assign w24178 = ~w24163 & ~w24177;
assign w24179 = ~w24150 & w24178;
assign w24180 = ~w23156 & ~w23157;
assign w24181 = w23171 & w24180;
assign w24182 = ~w23190 & ~w24181;
assign w24183 = ~w22258 & ~w23178;
assign w24184 = w22258 & w23178;
assign w24185 = ~w24183 & ~w24184;
assign w24186 = ~w23916 & w45337;
assign w24187 = w24185 & ~w24186;
assign w24188 = ~w23808 & ~w24182;
assign w24189 = w24187 & ~w24188;
assign w24190 = ~w17380 & ~w24182;
assign w24191 = w23183 & ~w24182;
assign w24192 = w23195 & ~w24191;
assign w24193 = (w24185 & ~w23842) | (w24185 & w47670) | (~w23842 & w47670);
assign w24194 = w23842 & w45338;
assign w24195 = ~w23808 & w24194;
assign w24196 = ~w24193 & ~w24195;
assign w24197 = ~w24189 & w24196;
assign w24198 = w16559 & w24197;
assign w24199 = w23089 & w23200;
assign w24200 = w24192 & ~w24199;
assign w24201 = ~w24192 & w24199;
assign w24202 = ~w24200 & ~w24201;
assign w24203 = w22269 & ~w22767;
assign w24204 = w22767 & ~w23084;
assign w24205 = ~w24203 & ~w24204;
assign w24206 = ~w23808 & w47671;
assign w24207 = (~w24205 & w23808) | (~w24205 & w47672) | (w23808 & w47672);
assign w24208 = ~w24206 & ~w24207;
assign w24209 = w15681 & ~w24208;
assign w24210 = w22282 & ~w23070;
assign w24211 = ~w22282 & w23070;
assign w24212 = ~w24210 & ~w24211;
assign w24213 = w23074 & w23079;
assign w24214 = w23200 & ~w24201;
assign w24215 = w24213 & ~w24214;
assign w24216 = ~w24213 & w24214;
assign w24217 = ~w24215 & ~w24216;
assign w24218 = ~w23843 & ~w24212;
assign w24219 = w23843 & w24217;
assign w24220 = ~w24218 & ~w24219;
assign w24221 = w14766 & ~w24220;
assign w24222 = ~w24198 & ~w24209;
assign w24223 = ~w24221 & w24222;
assign w24224 = w23171 & ~w23190;
assign w24225 = ~w24180 & w24224;
assign w24226 = (w18183 & ~w23917) | (w18183 & w45339) | (~w23917 & w45339);
assign w24227 = w24225 & ~w24226;
assign w24228 = (w23189 & w23808) | (w23189 & w47673) | (w23808 & w47673);
assign w24229 = ~w24227 & ~w24228;
assign w24230 = w24180 & ~w24224;
assign w24231 = w23843 & w24230;
assign w24232 = w24229 & ~w24231;
assign w24233 = (~w17380 & ~w24229) | (~w17380 & w47674) | (~w24229 & w47674);
assign w24234 = (w23842 & w47675) | (w23842 & w47676) | (w47675 & w47676);
assign w24235 = ~w24171 & w24234;
assign w24236 = ~w24154 & w24161;
assign w24237 = w24164 & w24165;
assign w24238 = w23842 & w24237;
assign w24239 = (~w24238 & w24154) | (~w24238 & w45340) | (w24154 & w45340);
assign w24240 = ~w24235 & w24239;
assign w24241 = (w18183 & ~w23808) | (w18183 & w47675) | (~w23808 & w47675);
assign w24242 = ~w24175 & ~w24241;
assign w24243 = ~w24240 & ~w24242;
assign w24244 = (~w18183 & w24171) | (~w18183 & w47677) | (w24171 & w47677);
assign w24245 = w24236 & ~w24244;
assign w24246 = ~w24243 & ~w24245;
assign w24247 = ~w24233 & w24246;
assign w24248 = w24229 & w47678;
assign w24249 = ~w16559 & ~w24197;
assign w24250 = ~w24248 & ~w24249;
assign w24251 = ~w14766 & w24220;
assign w24252 = ~w15681 & w24208;
assign w24253 = ~w24221 & w24252;
assign w24254 = ~w24251 & ~w24253;
assign w24255 = w24223 & ~w24250;
assign w24256 = w24254 & ~w24255;
assign w24257 = w24223 & w24247;
assign w24258 = ~w24179 & w24257;
assign w24259 = w24256 & ~w24258;
assign w24260 = w24040 & w24259;
assign w24261 = (w24035 & ~w24259) | (w24035 & w45341) | (~w24259 & w45341);
assign w24262 = ~w23428 & ~w23430;
assign w24263 = ~w2558 & w23420;
assign w24264 = ~w23027 & w45342;
assign w24265 = w23596 & w50211;
assign w24266 = w3242 & ~w23499;
assign w24267 = w3242 & w23485;
assign w24268 = (w42049 & w47679) | (w42049 & w47680) | (w47679 & w47680);
assign w24269 = ~w3242 & w23486;
assign w24270 = (w23371 & w45345) | (w23371 & w45346) | (w45345 & w45346);
assign w24271 = w23461 & w23487;
assign w24272 = (~w23371 & w45347) | (~w23371 & w45348) | (w45347 & w45348);
assign w24273 = w24270 & ~w24272;
assign w24274 = (~w24263 & w24273) | (~w24263 & w49054) | (w24273 & w49054);
assign w24275 = ~w24262 & w24274;
assign w24276 = w24262 & ~w24274;
assign w24277 = w23427 & ~w23843;
assign w24278 = w23843 & w49055;
assign w24279 = ~w24277 & ~w24278;
assign w24280 = ~w2006 & w24279;
assign w24281 = w2006 & ~w24279;
assign w24282 = ~w2558 & w24273;
assign w24283 = w2558 & ~w24273;
assign w24284 = ~w24282 & ~w24283;
assign w24285 = (w23420 & ~w23843) | (w23420 & w49056) | (~w23843 & w49056);
assign w24286 = w23843 & w49057;
assign w24287 = ~w24285 & ~w24286;
assign w24288 = w2285 & ~w24287;
assign w24289 = ~w24281 & ~w24288;
assign w24290 = ~w24280 & ~w24289;
assign w24291 = w23447 & ~w23518;
assign w24292 = ~w23605 & ~w23618;
assign w24293 = (w1541 & w23808) | (w1541 & w49058) | (w23808 & w49058);
assign w24294 = ~w23808 & w49059;
assign w24295 = ~w24293 & ~w24294;
assign w24296 = w24291 & w24295;
assign w24297 = ~w24291 & ~w24295;
assign w24298 = ~w24296 & ~w24297;
assign w24299 = w1320 & ~w24298;
assign w24300 = ~w23429 & w23433;
assign w24301 = ~w23394 & w23450;
assign w24302 = ~w23394 & ~w24300;
assign w24303 = (~w24302 & w24273) | (~w24302 & w49060) | (w24273 & w49060);
assign w24304 = w23403 & w23409;
assign w24305 = ~w24303 & ~w24304;
assign w24306 = w23843 & w24305;
assign w24307 = w22079 & ~w23398;
assign w24308 = ~w23438 & ~w24307;
assign w24309 = (w24308 & w23808) | (w24308 & w49061) | (w23808 & w49061);
assign w24310 = w24303 & w24304;
assign w24311 = w23843 & w24310;
assign w24312 = ~w24309 & ~w24311;
assign w24313 = (w1541 & ~w24312) | (w1541 & w49062) | (~w24312 & w49062);
assign w24314 = ~w23430 & ~w23450;
assign w24315 = ~w23394 & ~w23432;
assign w24316 = w24314 & ~w24315;
assign w24317 = ~w24314 & w24315;
assign w24318 = ~w24316 & ~w24317;
assign w24319 = ~w23430 & ~w24263;
assign w24320 = w23450 & w24319;
assign w24321 = (w24318 & ~w24273) | (w24318 & w49063) | (~w24273 & w49063);
assign w24322 = w24273 & w49064;
assign w24323 = ~w24321 & ~w24322;
assign w24324 = (w23393 & w23808) | (w23393 & w49065) | (w23808 & w49065);
assign w24325 = w23843 & ~w24323;
assign w24326 = ~w24324 & ~w24325;
assign w24327 = w1738 & ~w24326;
assign w24328 = ~w24313 & ~w24327;
assign w24329 = ~w24299 & w24328;
assign w24330 = ~w24290 & w24329;
assign w24331 = ~w2285 & w24287;
assign w24332 = w23461 & ~w23476;
assign w24333 = (~w23371 & w49066) | (~w23371 & w49067) | (w49066 & w49067);
assign w24334 = (~w23485 & ~w45344) | (~w23485 & w47681) | (~w45344 & w47681);
assign w24335 = (w47681 & w49068) | (w47681 & w49069) | (w49068 & w49069);
assign w24336 = ~w24333 & ~w24335;
assign w24337 = w24332 & ~w24336;
assign w24338 = ~w24332 & w24336;
assign w24339 = ~w24337 & ~w24338;
assign w24340 = ~w23475 & ~w23843;
assign w24341 = w23843 & w24339;
assign w24342 = ~w24340 & ~w24341;
assign w24343 = w2558 & w24342;
assign w24344 = ~w24280 & ~w24343;
assign w24345 = ~w24281 & w24331;
assign w24346 = w24344 & ~w24345;
assign w24347 = ~w2558 & ~w24342;
assign w24348 = (~w23488 & w23766) | (~w23488 & w45349) | (w23766 & w45349);
assign w24349 = ~w23916 & w49070;
assign w24350 = ~w24348 & ~w24349;
assign w24351 = (~w23487 & ~w23842) | (~w23487 & w49071) | (~w23842 & w49071);
assign w24352 = w23842 & w45350;
assign w24353 = ~w23808 & w24352;
assign w24354 = ~w24351 & ~w24353;
assign w24355 = ~w24350 & w24354;
assign w24356 = w2896 & w24355;
assign w24357 = ~w24347 & ~w24356;
assign w24358 = ~w2896 & ~w24355;
assign w24359 = w23371 & ~w24265;
assign w24360 = w23842 & ~w24359;
assign w24361 = ~w3646 & ~w23842;
assign w24362 = ~w3646 & ~w23807;
assign w24363 = ~w23766 & w24362;
assign w24364 = ~w24361 & ~w24363;
assign w24365 = ~w23808 & w24360;
assign w24366 = ~w23485 & ~w23499;
assign w24367 = w3242 & ~w24366;
assign w24368 = w24364 & w45351;
assign w24369 = w3242 & w24366;
assign w24370 = (w24369 & ~w24364) | (w24369 & w45352) | (~w24364 & w45352);
assign w24371 = ~w24368 & ~w24370;
assign w24372 = ~w24358 & w24371;
assign w24373 = w23349 & ~w23351;
assign w24374 = w23062 & ~w24373;
assign w24375 = ~w23356 & ~w23357;
assign w24376 = ~w23369 & w24375;
assign w24377 = ~w22800 & ~w24265;
assign w24378 = ~w22814 & ~w24374;
assign w24379 = w24377 & ~w24378;
assign w24380 = w24374 & ~w24376;
assign w24381 = w24379 & ~w24380;
assign w24382 = w23842 & w24381;
assign w24383 = ~w23808 & w24382;
assign w24384 = w22809 & ~w24383;
assign w24385 = ~w22809 & w24383;
assign w24386 = ~w24384 & ~w24385;
assign w24387 = ~w3646 & ~w24386;
assign w24388 = ~w3242 & ~w24366;
assign w24389 = (w24388 & ~w24364) | (w24388 & w45353) | (~w24364 & w45353);
assign w24390 = ~w3242 & w24366;
assign w24391 = w24364 & w45354;
assign w24392 = ~w24389 & ~w24391;
assign w24393 = ~w24387 & w24392;
assign w24394 = w24372 & ~w24393;
assign w24395 = w24357 & ~w24394;
assign w24396 = w24346 & ~w24395;
assign w24397 = w24330 & ~w24396;
assign w24398 = w23058 & ~w23372;
assign w24399 = (w23052 & w23330) | (w23052 & w49072) | (w23330 & w49072);
assign w24400 = (w42015 & w47682) | (w42015 & w47683) | (w47682 & w47683);
assign w24401 = ~w24399 & ~w24400;
assign w24402 = ~w5330 & ~w22898;
assign w24403 = ~w24400 & w49073;
assign w24404 = ~w23053 & ~w24403;
assign w24405 = ~w4838 & ~w24404;
assign w24406 = w23054 & ~w24403;
assign w24407 = ~w22883 & ~w24406;
assign w24408 = ~w24405 & ~w24407;
assign w24409 = w4430 & ~w22799;
assign w24410 = ~w4430 & w22799;
assign w24411 = ~w24409 & ~w24410;
assign w24412 = w24408 & w24411;
assign w24413 = ~w24408 & ~w24411;
assign w24414 = ~w24412 & ~w24413;
assign w24415 = (w22799 & w23808) | (w22799 & w49074) | (w23808 & w49074);
assign w24416 = w23843 & w24414;
assign w24417 = ~w24415 & ~w24416;
assign w24418 = ~w24416 & w49075;
assign w24419 = w23842 & w45356;
assign w24420 = ~w23808 & w24419;
assign w24421 = w22883 & ~w24420;
assign w24422 = ~w22883 & w24420;
assign w24423 = ~w24421 & ~w24422;
assign w24424 = ~w4430 & ~w24423;
assign w24425 = ~w24418 & ~w24424;
assign w24426 = ~w22861 & ~w24399;
assign w24427 = ~w24398 & w24426;
assign w24428 = ~w5330 & w22870;
assign w24429 = w23842 & w45357;
assign w24430 = ~w23808 & w24429;
assign w24431 = ~w5330 & ~w22870;
assign w24432 = (w24431 & ~w23842) | (w24431 & w45358) | (~w23842 & w45358);
assign w24433 = ~w23807 & w24431;
assign w24434 = ~w23766 & w24433;
assign w24435 = ~w24432 & ~w24434;
assign w24436 = ~w24430 & w24435;
assign w24437 = w5330 & ~w24401;
assign w24438 = ~w5330 & w24401;
assign w24439 = ~w24437 & ~w24438;
assign w24440 = w23842 & ~w24439;
assign w24441 = w4838 & w22898;
assign w24442 = w23842 & w45359;
assign w24443 = ~w23808 & w24442;
assign w24444 = w4838 & ~w22898;
assign w24445 = (w24444 & ~w23842) | (w24444 & w45360) | (~w23842 & w45360);
assign w24446 = ~w23807 & w24444;
assign w24447 = ~w23766 & w24446;
assign w24448 = ~w24445 & ~w24447;
assign w24449 = ~w24443 & w24448;
assign w24450 = w24436 & w24449;
assign w24451 = w5330 & ~w22870;
assign w24452 = w23842 & w45361;
assign w24453 = ~w23808 & w24452;
assign w24454 = w5330 & w22870;
assign w24455 = (w24454 & ~w23842) | (w24454 & w45362) | (~w23842 & w45362);
assign w24456 = ~w23807 & w24454;
assign w24457 = ~w23766 & w24456;
assign w24458 = ~w24455 & ~w24457;
assign w24459 = ~w24453 & w24458;
assign w24460 = (w23361 & w23330) | (w23361 & w45363) | (w23330 & w45363);
assign w24461 = ~w6769 & ~w24460;
assign w24462 = w6769 & w24460;
assign w24463 = ~w23041 & ~w24462;
assign w24464 = ~w24461 & ~w24463;
assign w24465 = w6264 & ~w24464;
assign w24466 = ~w6264 & w24464;
assign w24467 = ~w24465 & ~w24466;
assign w24468 = w23842 & w24467;
assign w24469 = ~w5745 & ~w22829;
assign w24470 = w23842 & w45364;
assign w24471 = ~w23808 & w24470;
assign w24472 = (w23362 & ~w23842) | (w23362 & w45365) | (~w23842 & w45365);
assign w24473 = w23362 & ~w23807;
assign w24474 = ~w23766 & w24473;
assign w24475 = ~w24472 & ~w24474;
assign w24476 = ~w24471 & w24475;
assign w24477 = w24459 & w24476;
assign w24478 = w24450 & ~w24477;
assign w24479 = ~w23808 & w24440;
assign w24480 = ~w4838 & ~w22898;
assign w24481 = w22908 & ~w24479;
assign w24482 = w24479 & w24480;
assign w24483 = ~w24481 & ~w24482;
assign w24484 = w4430 & ~w22883;
assign w24485 = ~w24420 & w24484;
assign w24486 = w4430 & w22883;
assign w24487 = w24420 & w24486;
assign w24488 = ~w24485 & ~w24487;
assign w24489 = w24483 & w24488;
assign w24490 = ~w24478 & w24489;
assign w24491 = w24425 & ~w24490;
assign w24492 = w4056 & ~w24417;
assign w24493 = ~w24461 & ~w24462;
assign w24494 = w23843 & w24493;
assign w24495 = w23041 & ~w24494;
assign w24496 = ~w23041 & w24494;
assign w24497 = ~w24495 & ~w24496;
assign w24498 = w6264 & w24497;
assign w24499 = ~w24492 & ~w24498;
assign w24500 = ~w24491 & w24499;
assign w24501 = w23346 & w23864;
assign w24502 = w22990 & ~w24501;
assign w24503 = ~w23025 & ~w24502;
assign w24504 = w23032 & ~w24503;
assign w24505 = w23016 & ~w24504;
assign w24506 = w23037 & ~w24505;
assign w24507 = ~w7315 & ~w23842;
assign w24508 = ~w7315 & ~w23807;
assign w24509 = ~w23766 & w24508;
assign w24510 = ~w24507 & ~w24509;
assign w24511 = w23842 & w24506;
assign w24512 = ~w23808 & w24511;
assign w24513 = w23002 & w23047;
assign w24514 = w24510 & w45366;
assign w24515 = (w24513 & ~w24510) | (w24513 & w45367) | (~w24510 & w45367);
assign w24516 = ~w24514 & ~w24515;
assign w24517 = w6769 & w24516;
assign w24518 = ~w6264 & ~w24497;
assign w24519 = ~w24517 & ~w24518;
assign w24520 = w7924 & ~w23842;
assign w24521 = w7924 & ~w23807;
assign w24522 = ~w23766 & w24521;
assign w24523 = ~w24520 & ~w24522;
assign w24524 = w23842 & ~w24504;
assign w24525 = ~w23808 & w24524;
assign w24526 = w24523 & ~w24525;
assign w24527 = w23016 & w23037;
assign w24528 = ~w7315 & ~w24527;
assign w24529 = w24523 & w45368;
assign w24530 = ~w7315 & w24527;
assign w24531 = (w24530 & ~w24523) | (w24530 & w45369) | (~w24523 & w45369);
assign w24532 = ~w24529 & ~w24531;
assign w24533 = ~w23025 & w23032;
assign w24534 = w24502 & ~w24533;
assign w24535 = ~w24502 & w24533;
assign w24536 = ~w24534 & ~w24535;
assign w24537 = ~w23024 & ~w23843;
assign w24538 = w23843 & w24536;
assign w24539 = ~w24537 & ~w24538;
assign w24540 = w7924 & ~w24539;
assign w24541 = w7315 & ~w24527;
assign w24542 = (w24541 & ~w24523) | (w24541 & w45370) | (~w24523 & w45370);
assign w24543 = w7315 & w24527;
assign w24544 = w24523 & w45371;
assign w24545 = ~w24542 & ~w24544;
assign w24546 = ~w6769 & w24513;
assign w24547 = (w24546 & ~w24510) | (w24546 & w45372) | (~w24510 & w45372);
assign w24548 = ~w6769 & ~w24513;
assign w24549 = w24510 & w45373;
assign w24550 = ~w24547 & ~w24549;
assign w24551 = w24545 & w24550;
assign w24552 = w24532 & w24540;
assign w24553 = w24551 & ~w24552;
assign w24554 = w24519 & ~w24553;
assign w24555 = w24500 & ~w24554;
assign w24556 = w24397 & w24555;
assign w24557 = ~w24261 & w24556;
assign w24558 = ~w23808 & w24468;
assign w24559 = ~w22829 & ~w24558;
assign w24560 = w22829 & w24558;
assign w24561 = ~w24559 & ~w24560;
assign w24562 = w5745 & ~w24561;
assign w24563 = w24459 & w24562;
assign w24564 = w24450 & ~w24563;
assign w24565 = (~w24492 & w24490) | (~w24492 & w45374) | (w24490 & w45374);
assign w24566 = w24425 & w24564;
assign w24567 = w24565 & ~w24566;
assign w24568 = ~w7924 & w24539;
assign w24569 = w24532 & ~w24568;
assign w24570 = w24551 & ~w24569;
assign w24571 = w24519 & ~w24570;
assign w24572 = w24500 & ~w24571;
assign w24573 = ~w24567 & ~w24572;
assign w24574 = w24397 & ~w24573;
assign w24575 = w3646 & w24386;
assign w24576 = w24392 & w24575;
assign w24577 = w24372 & ~w24576;
assign w24578 = w24357 & ~w24577;
assign w24579 = w24346 & ~w24578;
assign w24580 = w24330 & ~w24579;
assign w24581 = ~w24325 & w49076;
assign w24582 = (~w1541 & ~w23843) | (~w1541 & w49077) | (~w23843 & w49077);
assign w24583 = w24312 & w24582;
assign w24584 = ~w24581 & ~w24583;
assign w24585 = ~w24313 & ~w24584;
assign w24586 = ~w1320 & w24298;
assign w24587 = ~w23518 & w24292;
assign w24588 = w23447 & ~w24587;
assign w24589 = w1320 & ~w23842;
assign w24590 = w1320 & ~w23807;
assign w24591 = ~w23766 & w24590;
assign w24592 = ~w24589 & ~w24591;
assign w24593 = w23842 & ~w24588;
assign w24594 = ~w23808 & w24593;
assign w24595 = w24592 & ~w24594;
assign w24596 = ~w23527 & w23610;
assign w24597 = (~w24596 & ~w24592) | (~w24596 & w49078) | (~w24592 & w49078);
assign w24598 = w1120 & ~w24597;
assign w24599 = w24595 & w24596;
assign w24600 = w24598 & ~w24599;
assign w24601 = ~w24586 & ~w24600;
assign w24602 = ~w24299 & w24585;
assign w24603 = w24601 & ~w24602;
assign w24604 = w493 & ~w23696;
assign w24605 = (w23530 & ~w23371) | (w23530 & w42051) | (~w23371 & w42051);
assign w24606 = ~w23626 & ~w23630;
assign w24607 = (~w23543 & w24605) | (~w23543 & w42052) | (w24605 & w42052);
assign w24608 = ~w612 & w23562;
assign w24609 = w24606 & w24608;
assign w24610 = ~w24605 & w24609;
assign w24611 = ~w23543 & w23576;
assign w24612 = w24608 & ~w24611;
assign w24613 = w612 & w23588;
assign w24614 = w754 & w24613;
assign w24615 = ~w24612 & ~w24614;
assign w24616 = (w24615 & w24605) | (w24615 & w42053) | (w24605 & w42053);
assign w24617 = w23842 & w24616;
assign w24618 = w23577 & w24607;
assign w24619 = w24617 & ~w24618;
assign w24620 = ~w23808 & w24619;
assign w24621 = w493 & w23696;
assign w24622 = (w24604 & ~w24619) | (w24604 & w45375) | (~w24619 & w45375);
assign w24623 = w24619 & w45376;
assign w24624 = ~w24622 & ~w24623;
assign w24625 = w23562 & w23576;
assign w24626 = w24607 & ~w24625;
assign w24627 = ~w24607 & w24625;
assign w24628 = ~w24626 & ~w24627;
assign w24629 = (w24613 & w23808) | (w24613 & w42054) | (w23808 & w42054);
assign w24630 = w612 & ~w24628;
assign w24631 = w23843 & w24630;
assign w24632 = ~w24629 & ~w24631;
assign w24633 = w24624 & w24632;
assign w24634 = ~w23505 & w23529;
assign w24635 = w23610 & ~w24634;
assign w24636 = w1120 & ~w23842;
assign w24637 = (w1120 & w23805) | (w1120 & w42055) | (w23805 & w42055);
assign w24638 = ~w23766 & w24637;
assign w24639 = ~w24636 & ~w24638;
assign w24640 = w23842 & w24635;
assign w24641 = ~w23808 & w24640;
assign w24642 = w24639 & ~w24641;
assign w24643 = ~w23514 & ~w23628;
assign w24644 = w945 & ~w24643;
assign w24645 = (w24644 & ~w24639) | (w24644 & w45377) | (~w24639 & w45377);
assign w24646 = w945 & w24643;
assign w24647 = w24639 & w45378;
assign w24648 = ~w24645 & ~w24647;
assign w24649 = ~w23630 & ~w24605;
assign w24650 = ~w945 & ~w23842;
assign w24651 = (~w945 & w23805) | (~w945 & w42056) | (w23805 & w42056);
assign w24652 = ~w23766 & w24651;
assign w24653 = ~w24650 & ~w24652;
assign w24654 = w23842 & ~w24649;
assign w24655 = ~w23808 & w24654;
assign w24656 = w24653 & ~w24655;
assign w24657 = ~w23543 & ~w23626;
assign w24658 = w754 & ~w24657;
assign w24659 = (w24658 & ~w24653) | (w24658 & w45379) | (~w24653 & w45379);
assign w24660 = w754 & w24657;
assign w24661 = w24653 & w45380;
assign w24662 = ~w24659 & ~w24661;
assign w24663 = ~w24648 & w24662;
assign w24664 = (w23588 & w23808) | (w23588 & w42057) | (w23808 & w42057);
assign w24665 = ~w23808 & w42058;
assign w24666 = ~w24664 & ~w24665;
assign w24667 = ~w612 & w24666;
assign w24668 = ~w754 & ~w24657;
assign w24669 = w24653 & w45381;
assign w24670 = ~w754 & w24657;
assign w24671 = (w24670 & ~w24653) | (w24670 & w45382) | (~w24653 & w45382);
assign w24672 = ~w24669 & ~w24671;
assign w24673 = ~w24667 & w24672;
assign w24674 = ~w24663 & w24673;
assign w24675 = w24633 & ~w24674;
assign w24676 = w23710 & ~w23711;
assign w24677 = ~w23710 & w23711;
assign w24678 = ~w24676 & ~w24677;
assign w24679 = ~w493 & ~w23731;
assign w24680 = w23576 & ~w23627;
assign w24681 = w23699 & w24679;
assign w24682 = w24679 & ~w24680;
assign w24683 = ~w24605 & w42059;
assign w24684 = ~w24681 & ~w24683;
assign w24685 = w24604 & ~w24612;
assign w24686 = w493 & ~w23640;
assign w24687 = ~w24610 & w24685;
assign w24688 = ~w24686 & ~w24687;
assign w24689 = (~w24678 & ~w23843) | (~w24678 & w42060) | (~w23843 & w42060);
assign w24690 = w23843 & w42061;
assign w24691 = ~w24689 & ~w24690;
assign w24692 = w400 & ~w24691;
assign w24693 = w24619 & w49079;
assign w24694 = ~w493 & ~w24693;
assign w24695 = ~w23696 & ~w24620;
assign w24696 = w24694 & ~w24695;
assign w24697 = ~w24692 & ~w24696;
assign w24698 = (w24697 & w24674) | (w24697 & w42062) | (w24674 & w42062);
assign w24699 = w24603 & w24698;
assign w24700 = ~w24580 & w24699;
assign w24701 = ~w24574 & w24700;
assign w24702 = ~w24557 & w24701;
assign w24703 = ~w24035 & w24555;
assign w24704 = w24040 & w24555;
assign w24705 = w24259 & w24704;
assign w24706 = ~w24703 & ~w24705;
assign w24707 = w24573 & w45383;
assign w24708 = w24706 & w24707;
assign w24709 = (~w23768 & w23753) | (~w23768 & w42063) | (w23753 & w42063);
assign w24710 = w23842 & ~w24709;
assign w24711 = ~w23640 & w42064;
assign w24712 = w24710 & ~w24711;
assign w24713 = w252 & ~w23842;
assign w24714 = (w252 & w23805) | (w252 & w42065) | (w23805 & w42065);
assign w24715 = ~w23766 & w24714;
assign w24716 = ~w24713 & ~w24715;
assign w24717 = ~w23808 & w24712;
assign w24718 = w24716 & ~w24717;
assign w24719 = ~w23681 & ~w23767;
assign w24720 = ~w57 & w24719;
assign w24721 = ~w24718 & w24720;
assign w24722 = ~w57 & ~w24719;
assign w24723 = w24718 & w24722;
assign w24724 = ~w24721 & ~w24723;
assign w24725 = ~w23730 & ~w23768;
assign w24726 = ~w23721 & ~w23738;
assign w24727 = ~w23830 & w24726;
assign w24728 = ~w23844 & w24727;
assign w24729 = (w24725 & w24003) | (w24725 & w42066) | (w24003 & w42066);
assign w24730 = ~w24003 & w42067;
assign w24731 = ~w24729 & ~w24730;
assign w24732 = (w23729 & w23808) | (w23729 & w42068) | (w23808 & w42068);
assign w24733 = w23843 & w24731;
assign w24734 = (~w252 & w24733) | (~w252 & w42069) | (w24733 & w42069);
assign w24735 = w24724 & ~w24734;
assign w24736 = w24678 & w24684;
assign w24737 = w24688 & ~w24736;
assign w24738 = w400 & w23842;
assign w24739 = ~w23808 & w24738;
assign w24740 = ~w24737 & w24739;
assign w24741 = ~w400 & w23842;
assign w24742 = ~w23808 & w24741;
assign w24743 = w24737 & w24742;
assign w24744 = ~w24740 & ~w24743;
assign w24745 = w23705 & w24744;
assign w24746 = ~w23705 & ~w24744;
assign w24747 = ~w24745 & ~w24746;
assign w24748 = w351 & ~w24747;
assign w24749 = ~w945 & w24643;
assign w24750 = (w24749 & ~w24639) | (w24749 & w45384) | (~w24639 & w45384);
assign w24751 = ~w945 & ~w24643;
assign w24752 = w24639 & w45385;
assign w24753 = ~w24750 & ~w24752;
assign w24754 = ~w1120 & ~w24596;
assign w24755 = (w24754 & ~w24592) | (w24754 & w45386) | (~w24592 & w45386);
assign w24756 = ~w1120 & w24596;
assign w24757 = w24592 & w45387;
assign w24758 = ~w24755 & ~w24757;
assign w24759 = w24753 & w24758;
assign w24760 = w24633 & w24662;
assign w24761 = w24759 & w24760;
assign w24762 = w24697 & ~w24761;
assign w24763 = ~w24675 & w24762;
assign w24764 = ~w400 & w24691;
assign w24765 = ~w24763 & ~w24764;
assign w24766 = ~w24763 & w42070;
assign w24767 = w24735 & w24766;
assign w24768 = (w24767 & ~w24706) | (w24767 & w45388) | (~w24706 & w45388);
assign w24769 = ~w24702 & w24768;
assign w24770 = ~w351 & ~w23705;
assign w24771 = w24744 & w24770;
assign w24772 = ~w351 & w23705;
assign w24773 = ~w24744 & w24772;
assign w24774 = ~w24771 & ~w24773;
assign w24775 = w24718 & ~w24719;
assign w24776 = ~w24718 & w24719;
assign w24777 = ~w24775 & ~w24776;
assign w24778 = w57 & w24777;
assign w24779 = ~w24733 & w42071;
assign w24780 = w24724 & w24779;
assign w24781 = ~w24778 & ~w24780;
assign w24782 = w24735 & ~w24774;
assign w24783 = w24781 & ~w24782;
assign w24784 = ~w80 & w23862;
assign w24785 = w24783 & ~w24784;
assign w24786 = (~w23863 & w24769) | (~w23863 & w42072) | (w24769 & w42072);
assign w24787 = ~w23863 & ~w24783;
assign w24788 = w3 & w23842;
assign w24789 = ~w23808 & w24788;
assign w24790 = w80 & ~w23655;
assign w24791 = ~w23658 & ~w24790;
assign w24792 = ~w23854 & ~w24791;
assign w24793 = ~w23656 & w23682;
assign w24794 = ~w24790 & ~w24793;
assign w24795 = ~w23848 & w24792;
assign w24796 = w24794 & ~w24795;
assign w24797 = ~w3 & w23842;
assign w24798 = ~w23808 & w24797;
assign w24799 = w24789 & ~w24796;
assign w24800 = w24796 & w24798;
assign w24801 = ~w24799 & ~w24800;
assign w24802 = (w23745 & w23760) | (w23745 & w42073) | (w23760 & w42073);
assign w24803 = ~w23771 & ~w24802;
assign w24804 = ~w24085 & w24093;
assign w24805 = ~w23766 & w24803;
assign w24806 = ~w24804 & ~w24805;
assign w24807 = ~w23772 & w23777;
assign w24808 = ~w42 & ~w24807;
assign w24809 = w23772 & ~w23777;
assign w24810 = w24808 & ~w24809;
assign w24811 = w23795 & ~w24810;
assign w24812 = w24806 & ~w24811;
assign w24813 = ~w23801 & ~w24810;
assign w24814 = ~w24806 & w24813;
assign w24815 = ~w24812 & ~w24814;
assign w24816 = w42 & w23665;
assign w24817 = w24801 & w24816;
assign w24818 = w42 & ~w23665;
assign w24819 = ~w24801 & w24818;
assign w24820 = ~w24817 & ~w24819;
assign w24821 = ~w24815 & w24820;
assign w24822 = (~w80 & w23808) | (~w80 & w42074) | (w23808 & w42074);
assign w24823 = (~w23682 & ~w23855) | (~w23682 & w42075) | (~w23855 & w42075);
assign w24824 = w23843 & w24823;
assign w24825 = ~w24822 & ~w24824;
assign w24826 = ~w23656 & ~w24790;
assign w24827 = w3 & ~w24826;
assign w24828 = (w24827 & w24824) | (w24827 & w42076) | (w24824 & w42076);
assign w24829 = w3 & w24826;
assign w24830 = ~w24824 & w42077;
assign w24831 = ~w24828 & ~w24830;
assign w24832 = ~w24784 & w24831;
assign w24833 = w24821 & w24832;
assign w24834 = ~w23863 & w24735;
assign w24835 = ~w24748 & w24834;
assign w24836 = w24833 & ~w24835;
assign w24837 = ~w24787 & w24836;
assign w24838 = (~w23821 & ~w24806) | (~w23821 & w42078) | (~w24806 & w42078);
assign w24839 = w24806 & w24810;
assign w24840 = ~w24838 & ~w24839;
assign w24841 = (w23665 & w24795) | (w23665 & w42079) | (w24795 & w42079);
assign w24842 = w24789 & w24841;
assign w24843 = (~w23665 & w24795) | (~w23665 & w42080) | (w24795 & w42080);
assign w24844 = ~w24789 & w24843;
assign w24845 = ~w24842 & ~w24844;
assign w24846 = ~w24795 & w42081;
assign w24847 = ~w24798 & w24846;
assign w24848 = ~w24795 & w42082;
assign w24849 = w24798 & w24848;
assign w24850 = ~w24847 & ~w24849;
assign w24851 = w24845 & w24850;
assign w24852 = ~w24840 & ~w24851;
assign w24853 = ~w3 & w24826;
assign w24854 = (w24853 & w24824) | (w24853 & w42083) | (w24824 & w42083);
assign w24855 = ~w3 & ~w24826;
assign w24856 = ~w24824 & w42084;
assign w24857 = ~w24854 & ~w24856;
assign w24858 = ~w24852 & w24857;
assign w24859 = w24821 & ~w24858;
assign w24860 = ~w24764 & ~w24859;
assign w24861 = ~w24763 & w24860;
assign w24862 = ~w24837 & w24861;
assign w24863 = (w24833 & w24783) | (w24833 & w45389) | (w24783 & w45389);
assign w24864 = (~w24859 & w24787) | (~w24859 & w42085) | (w24787 & w42085);
assign w24865 = ~w24862 & ~w24864;
assign w24866 = ~w24580 & w24603;
assign w24867 = ~w24574 & w24866;
assign w24868 = ~w24837 & ~w24859;
assign w24869 = ~w24698 & ~w24764;
assign w24870 = w24863 & ~w24869;
assign w24871 = w24868 & ~w24870;
assign w24872 = w24867 & ~w24871;
assign w24873 = ~w24557 & w24872;
assign w24874 = (~w24865 & ~w24872) | (~w24865 & w45390) | (~w24872 & w45390);
assign w24875 = w24831 & w24857;
assign w24876 = w24825 & ~w24826;
assign w24877 = ~w24825 & w24826;
assign w24878 = ~w24876 & ~w24877;
assign w24879 = ~w24874 & ~w24878;
assign w24880 = w24874 & w24875;
assign w24881 = w24786 & w24880;
assign w24882 = w24874 & ~w24875;
assign w24883 = ~w24786 & w24882;
assign w24884 = ~w24881 & ~w24883;
assign w24885 = ~w24879 & w24884;
assign w24886 = w23958 & ~w24017;
assign w24887 = ~w24258 & w45391;
assign w24888 = ~w24013 & ~w24018;
assign w24889 = ~w24887 & w24888;
assign w24890 = (w24016 & w24873) | (w24016 & w42086) | (w24873 & w42086);
assign w24891 = w24886 & ~w24889;
assign w24892 = ~w24873 & w42087;
assign w24893 = ~w24890 & ~w24892;
assign w24894 = w24261 & w24867;
assign w24895 = ~w24397 & w24603;
assign w24896 = ~w24567 & w24579;
assign w24897 = ~w24555 & w24603;
assign w24898 = w24896 & w24897;
assign w24899 = ~w24895 & ~w24898;
assign w24900 = w24862 & w24899;
assign w24901 = ~w24894 & w24900;
assign w24902 = (~w24016 & ~w24868) | (~w24016 & w45392) | (~w24868 & w45392);
assign w24903 = ~w24886 & w24889;
assign w24904 = (w24903 & w24901) | (w24903 & w42088) | (w24901 & w42088);
assign w24905 = w11138 & ~w24904;
assign w24906 = w24893 & w24905;
assign w24907 = ~w23926 & ~w23945;
assign w24908 = (~w24907 & w24873) | (~w24907 & w42089) | (w24873 & w42089);
assign w24909 = ~w24013 & w24019;
assign w24910 = (w24258 & w45393) | (w24258 & w45394) | (w45393 & w45394);
assign w24911 = w23928 & ~w23947;
assign w24912 = w24910 & ~w24911;
assign w24913 = ~w23958 & ~w24911;
assign w24914 = (~w24913 & w24862) | (~w24913 & w42091) | (w24862 & w42091);
assign w24915 = ~w24912 & w24914;
assign w24916 = ~w24873 & w24915;
assign w24917 = ~w24908 & ~w24916;
assign w24918 = (~w11138 & ~w24868) | (~w11138 & w45395) | (~w24868 & w45395);
assign w24919 = w23928 & w23959;
assign w24920 = ~w24910 & w24919;
assign w24921 = (w24920 & w24901) | (w24920 & w42092) | (w24901 & w42092);
assign w24922 = ~w10419 & ~w24921;
assign w24923 = ~w24917 & w24922;
assign w24924 = ~w24906 & ~w24923;
assign w24925 = (w24901 & w45396) | (w24901 & w45397) | (w45396 & w45397);
assign w24926 = (w10419 & w24873) | (w10419 & w42093) | (w24873 & w42093);
assign w24927 = ~w24908 & w24926;
assign w24928 = ~w24925 & ~w24927;
assign w24929 = w24893 & ~w24904;
assign w24930 = (~w11138 & ~w24893) | (~w11138 & w45398) | (~w24893 & w45398);
assign w24931 = ~w23996 & ~w24036;
assign w24932 = w24259 & w24931;
assign w24933 = (w24258 & w45399) | (w24258 & w45400) | (w45399 & w45400);
assign w24934 = w12666 & ~w23987;
assign w24935 = ~w12666 & w23987;
assign w24936 = ~w24934 & ~w24935;
assign w24937 = w24933 & ~w24936;
assign w24938 = ~w24933 & w24936;
assign w24939 = ~w24937 & ~w24938;
assign w24940 = (w24010 & w24873) | (w24010 & w45401) | (w24873 & w45401);
assign w24941 = ~w24871 & ~w24901;
assign w24942 = ~w24010 & w24939;
assign w24943 = (w24942 & w24901) | (w24942 & w45402) | (w24901 & w45402);
assign w24944 = (w11870 & w42096) | (w11870 & w24941) | (w42096 & w24941);
assign w24945 = ~w24940 & w24944;
assign w24946 = ~w24924 & w24928;
assign w24947 = w24928 & ~w24945;
assign w24948 = ~w24930 & w24947;
assign w24949 = ~w24946 & ~w24948;
assign w24950 = ~w23989 & w52254;
assign w24951 = ~w24933 & ~w24950;
assign w24952 = w23986 & w24951;
assign w24953 = (w23986 & ~w24868) | (w23986 & w49080) | (~w24868 & w49080);
assign w24954 = (~w24952 & w24901) | (~w24952 & w45405) | (w24901 & w45405);
assign w24955 = ~w24873 & w42098;
assign w24956 = w24954 & ~w24955;
assign w24957 = w12666 & ~w24956;
assign w24958 = ~w24259 & ~w24931;
assign w24959 = ~w24901 & w42099;
assign w24960 = ~w24932 & ~w24958;
assign w24961 = (w24960 & w24901) | (w24960 & w42100) | (w24901 & w42100);
assign w24962 = ~w24959 & ~w24961;
assign w24963 = w13384 & ~w24962;
assign w24964 = w24954 & w42101;
assign w24965 = ~w24963 & ~w24964;
assign w24966 = ~w24957 & ~w24965;
assign w24967 = ~w24940 & ~w24943;
assign w24968 = ~w11870 & ~w24967;
assign w24969 = w24924 & ~w24968;
assign w24970 = ~w24966 & w24969;
assign w24971 = ~w24949 & ~w24970;
assign w24972 = w24526 & ~w24527;
assign w24973 = ~w24526 & w24527;
assign w24974 = ~w24972 & ~w24973;
assign w24975 = (~w24974 & w24873) | (~w24974 & w45406) | (w24873 & w45406);
assign w24976 = (~w24540 & w24022) | (~w24540 & w45407) | (w24022 & w45407);
assign w24977 = w23977 & w47684;
assign w24978 = w24259 & w24977;
assign w24979 = ~w24976 & ~w24978;
assign w24980 = w24545 & ~w24979;
assign w24981 = w24874 & ~w24980;
assign w24982 = ~w24975 & ~w24981;
assign w24983 = ~w24978 & w47685;
assign w24984 = ~w24978 & w45408;
assign w24985 = (~w24901 & w45409) | (~w24901 & w45410) | (w45409 & w45410);
assign w24986 = w6769 & w24985;
assign w24987 = ~w24982 & w24986;
assign w24988 = w7924 & ~w24261;
assign w24989 = ~w7924 & w24261;
assign w24990 = ~w24988 & ~w24989;
assign w24991 = (w24539 & ~w24874) | (w24539 & w42104) | (~w24874 & w42104);
assign w24992 = w24874 & w42105;
assign w24993 = ~w24991 & ~w24992;
assign w24994 = ~w7315 & ~w24993;
assign w24995 = ~w24987 & ~w24994;
assign w24996 = ~w24258 & w45411;
assign w24997 = w23976 & ~w24021;
assign w24998 = w24031 & ~w24997;
assign w24999 = ~w24996 & w47686;
assign w25000 = (w9195 & w24996) | (w9195 & w47687) | (w24996 & w47687);
assign w25001 = ~w24999 & ~w25000;
assign w25002 = (w24025 & ~w24874) | (w24025 & w42107) | (~w24874 & w42107);
assign w25003 = w24874 & w42108;
assign w25004 = ~w25002 & ~w25003;
assign w25005 = ~w8666 & ~w25004;
assign w25006 = w23875 & ~w23876;
assign w25007 = ~w23875 & w23876;
assign w25008 = ~w25006 & ~w25007;
assign w25009 = ~w24556 & w24872;
assign w25010 = w23881 & w23886;
assign w25011 = ~w24026 & w24998;
assign w25012 = ~w24996 & w25011;
assign w25013 = w23898 & ~w25012;
assign w25014 = (w24872 & w47688) | (w24872 & w47689) | (w47688 & w47689);
assign w25015 = ~w25010 & w25013;
assign w25016 = w25010 & ~w25013;
assign w25017 = ~w25015 & ~w25016;
assign w25018 = ~w25014 & w25017;
assign w25019 = ~w24901 & w45412;
assign w25020 = ~w25018 & ~w25019;
assign w25021 = ~w25018 & w45413;
assign w25022 = ~w25005 & ~w25021;
assign w25023 = w24995 & w25022;
assign w25024 = w8666 & w25004;
assign w25025 = w23967 & ~w23968;
assign w25026 = ~w23967 & w23968;
assign w25027 = ~w25025 & ~w25026;
assign w25028 = w23973 & w24031;
assign w25029 = ~w23942 & ~w23960;
assign w25030 = w24919 & w25029;
assign w25031 = ~w24910 & w25030;
assign w25032 = ~w23943 & ~w23960;
assign w25033 = ~w25031 & ~w25032;
assign w25034 = w25028 & ~w25033;
assign w25035 = ~w25028 & w25033;
assign w25036 = ~w24901 & w45414;
assign w25037 = ~w24941 & w42110;
assign w25038 = ~w25036 & ~w25037;
assign w25039 = ~w25037 & w45415;
assign w25040 = ~w25024 & ~w25039;
assign w25041 = ~w24901 & w42111;
assign w25042 = w23959 & ~w24910;
assign w25043 = w23928 & ~w25042;
assign w25044 = (w23941 & w24873) | (w23941 & w42112) | (w24873 & w42112);
assign w25045 = w25029 & ~w25043;
assign w25046 = w24874 & w25045;
assign w25047 = ~w25044 & ~w25046;
assign w25048 = ~w25029 & w25043;
assign w25049 = ~w25041 & w25048;
assign w25050 = w25047 & ~w25049;
assign w25051 = w25047 & w42113;
assign w25052 = (w9195 & w25037) | (w9195 & w45416) | (w25037 & w45416);
assign w25053 = ~w25051 & ~w25052;
assign w25054 = w25040 & ~w25053;
assign w25055 = w25023 & ~w25054;
assign w25056 = ~w24971 & w25055;
assign w25057 = (w9781 & ~w25047) | (w9781 & w42114) | (~w25047 & w42114);
assign w25058 = ~w25052 & w25057;
assign w25059 = w25040 & ~w25058;
assign w25060 = w25023 & ~w25059;
assign w25061 = w7315 & w24993;
assign w25062 = (w7924 & w25018) | (w7924 & w45417) | (w25018 & w45417);
assign w25063 = ~w25061 & ~w25062;
assign w25064 = w24995 & ~w25063;
assign w25065 = w24532 & w24545;
assign w25066 = ~w6769 & w24532;
assign w25067 = w8205 & ~w24974;
assign w25068 = ~w25066 & ~w25067;
assign w25069 = (w42115 & w24978) | (w42115 & w45418) | (w24978 & w45418);
assign w25070 = (w25068 & w42116) | (w25068 & w24979) | (w42116 & w24979);
assign w25071 = ~w25069 & ~w25070;
assign w25072 = (w24516 & ~w24874) | (w24516 & w42117) | (~w24874 & w42117);
assign w25073 = ~w24941 & w42118;
assign w25074 = ~w25073 & w47690;
assign w25075 = ~w24982 & w24985;
assign w25076 = (~w6769 & w24982) | (~w6769 & w47691) | (w24982 & w47691);
assign w25077 = ~w25074 & ~w25076;
assign w25078 = ~w25064 & w25077;
assign w25079 = ~w25060 & w25078;
assign w25080 = ~w25056 & w25079;
assign w25081 = ~w23808 & w24238;
assign w25082 = ~w24236 & ~w25081;
assign w25083 = ~w24150 & ~w24163;
assign w25084 = w25082 & ~w25083;
assign w25085 = ~w18183 & w25084;
assign w25086 = w18183 & ~w25084;
assign w25087 = ~w25085 & ~w25086;
assign w25088 = (~w24176 & ~w24868) | (~w24176 & w47692) | (~w24868 & w47692);
assign w25089 = w24176 & w25087;
assign w25090 = ~w24873 & w42119;
assign w25091 = ~w24176 & ~w25087;
assign w25092 = (~w25091 & w24901) | (~w25091 & w42120) | (w24901 & w42120);
assign w25093 = ~w25090 & w25092;
assign w25094 = ~w17380 & ~w25093;
assign w25095 = ~w24150 & ~w24151;
assign w25096 = w19040 & ~w25095;
assign w25097 = ~w19040 & w25095;
assign w25098 = ~w25096 & ~w25097;
assign w25099 = (w24158 & w24873) | (w24158 & w42121) | (w24873 & w42121);
assign w25100 = ~w24873 & w42122;
assign w25101 = ~w25099 & ~w25100;
assign w25102 = w18183 & ~w25101;
assign w25103 = ~w25094 & ~w25102;
assign w25104 = w19040 & ~w24142;
assign w25105 = ~w24083 & ~w24126;
assign w25106 = ~w21010 & ~w24143;
assign w25107 = ~w25105 & ~w25106;
assign w25108 = ~w24083 & ~w25104;
assign w25109 = w25107 & ~w25108;
assign w25110 = w24126 & w24148;
assign w25111 = ~w24083 & w25110;
assign w25112 = ~w24127 & w24148;
assign w25113 = ~w20000 & w25112;
assign w25114 = ~w24865 & ~w25113;
assign w25115 = ~w24873 & w25114;
assign w25116 = w20000 & ~w25105;
assign w25117 = w19040 & ~w25113;
assign w25118 = ~w25116 & ~w25117;
assign w25119 = w24148 & ~w25104;
assign w25120 = w25109 & ~w25119;
assign w25121 = ~w25095 & ~w25118;
assign w25122 = ~w25120 & ~w25121;
assign w25123 = (~w25122 & w24901) | (~w25122 & w47693) | (w24901 & w47693);
assign w25124 = (w25104 & w24873) | (w25104 & w47694) | (w24873 & w47694);
assign w25125 = ~w25123 & ~w25124;
assign w25126 = w25109 & ~w25111;
assign w25127 = w24941 & w25126;
assign w25128 = w25125 & ~w25127;
assign w25129 = w25103 & w25128;
assign w25130 = w24100 & ~w24117;
assign w25131 = w21801 & ~w25130;
assign w25132 = ~w24100 & ~w24107;
assign w25133 = w25131 & ~w25132;
assign w25134 = ~w24100 & w24113;
assign w25135 = w24100 & ~w24121;
assign w25136 = ~w25134 & ~w25135;
assign w25137 = ~w25133 & ~w25136;
assign w25138 = ~a[28] & w23843;
assign w25139 = ~a[29] & w25138;
assign w25140 = ~w23843 & ~w24116;
assign w25141 = ~w24105 & ~w25140;
assign w25142 = ~w25139 & w25141;
assign w25143 = ~w24103 & ~w25142;
assign w25144 = ~w21801 & ~w25143;
assign w25145 = ~w25133 & ~w25144;
assign w25146 = ~w24100 & w24109;
assign w25147 = w24100 & w24115;
assign w25148 = ~w25146 & ~w25147;
assign w25149 = ~w25145 & ~w25148;
assign w25150 = (~w25148 & ~w24868) | (~w25148 & w47695) | (~w24868 & w47695);
assign w25151 = (~w25149 & w24901) | (~w25149 & w42123) | (w24901 & w42123);
assign w25152 = ~w24941 & w25137;
assign w25153 = w25151 & ~w25152;
assign w25154 = w20906 & ~w25153;
assign w25155 = w22767 & w23843;
assign w25156 = ~w24103 & ~w25155;
assign w25157 = ~w25138 & ~w25156;
assign w25158 = ~w23843 & w24104;
assign w25159 = a[29] & ~w25158;
assign w25160 = ~w25157 & w25159;
assign w25161 = w23843 & ~w24868;
assign w25162 = w24050 & ~w25155;
assign w25163 = ~w24101 & ~w25162;
assign w25164 = ~w25161 & w25163;
assign w25165 = w25160 & ~w25164;
assign w25166 = w22767 & w24863;
assign w25167 = w24868 & ~w25166;
assign w25168 = ~w24869 & w25160;
assign w25169 = ~w25167 & w25168;
assign w25170 = ~w24898 & w45419;
assign w25171 = ~w24894 & w25170;
assign w25172 = w25169 & ~w25171;
assign w25173 = ~w24871 & ~w25138;
assign w25174 = ~w24901 & w25173;
assign w25175 = w24102 & w25162;
assign w25176 = ~w24865 & w25175;
assign w25177 = ~w24873 & w25176;
assign w25178 = ~w25174 & ~w25177;
assign w25179 = ~w25165 & ~w25172;
assign w25180 = w25178 & ~w25179;
assign w25181 = ~w24102 & ~w25138;
assign w25182 = w25162 & w25181;
assign w25183 = ~w24873 & w42124;
assign w25184 = ~a[29] & ~w25183;
assign w25185 = ~w25180 & ~w25184;
assign w25186 = w23091 & w24101;
assign w25187 = ~w25162 & w25186;
assign w25188 = w22767 & w25187;
assign w25189 = ~w24859 & w25187;
assign w25190 = (~w25188 & w24837) | (~w25188 & w42125) | (w24837 & w42125);
assign w25191 = w24765 & ~w25190;
assign w25192 = ~w24708 & w25191;
assign w25193 = ~w22767 & ~w24101;
assign w25194 = w24862 & ~w25193;
assign w25195 = ~w24708 & w25194;
assign w25196 = w24864 & ~w25193;
assign w25197 = w25139 & ~w25196;
assign w25198 = (w25197 & ~w25195) | (w25197 & w45420) | (~w25195 & w45420);
assign w25199 = ~w22767 & ~w24864;
assign w25200 = w25187 & ~w25199;
assign w25201 = (~w25200 & ~w25192) | (~w25200 & w45421) | (~w25192 & w45421);
assign w25202 = ~w25198 & w25201;
assign w25203 = ~w25185 & w25202;
assign w25204 = ~w20906 & ~w25137;
assign w25205 = (~w25204 & w24901) | (~w25204 & w42126) | (w24901 & w42126);
assign w25206 = w25151 & ~w25205;
assign w25207 = ~w21801 & ~w25206;
assign w25208 = ~w25185 & w42127;
assign w25209 = ~w25154 & ~w25208;
assign w25210 = w25202 & ~w25206;
assign w25211 = (~w25207 & w25185) | (~w25207 & w45422) | (w25185 & w45422);
assign w25212 = ~a[24] & ~a[25];
assign w25213 = ~a[26] & w25212;
assign w25214 = w23843 & w25213;
assign w25215 = ~w23843 & ~w25213;
assign w25216 = w24101 & ~w25214;
assign w25217 = a[27] & w25215;
assign w25218 = ~w25216 & ~w25217;
assign w25219 = ~a[27] & ~w25215;
assign w25220 = ~w25214 & ~w25219;
assign w25221 = (w25218 & w24901) | (w25218 & w45423) | (w24901 & w45423);
assign w25222 = ~w24901 & w45424;
assign w25223 = ~w25221 & ~w25222;
assign w25224 = w22767 & ~w25223;
assign w25225 = ~w22767 & w25223;
assign w25226 = a[28] & ~w23843;
assign w25227 = ~w24901 & w49081;
assign w25228 = a[28] & ~w24101;
assign w25229 = ~w24102 & ~w25228;
assign w25230 = (w25229 & w24901) | (w25229 & w49082) | (w24901 & w49082);
assign w25231 = ~w25227 & ~w25230;
assign w25232 = ~w25225 & ~w25231;
assign w25233 = ~w25224 & ~w25232;
assign w25234 = w25129 & ~w25209;
assign w25235 = w25129 & ~w25211;
assign w25236 = ~w25233 & w25235;
assign w25237 = ~w25234 & ~w25236;
assign w25238 = w17380 & w25093;
assign w25239 = (w25110 & w24901) | (w25110 & w42128) | (w24901 & w42128);
assign w25240 = w21009 & ~w24083;
assign w25241 = (~w24901 & w45425) | (~w24901 & w45426) | (w45425 & w45426);
assign w25242 = ~w19040 & w24148;
assign w25243 = w24151 & ~w25242;
assign w25244 = ~w25112 & ~w25243;
assign w25245 = ~w24143 & w25244;
assign w25246 = (w25245 & w24901) | (w25245 & w45427) | (w24901 & w45427);
assign w25247 = w25097 & w25112;
assign w25248 = (w24142 & w24873) | (w24142 & w45428) | (w24873 & w45428);
assign w25249 = w24874 & w25247;
assign w25250 = ~w25248 & ~w25249;
assign w25251 = ~w20000 & ~w24083;
assign w25252 = (~w24901 & w45429) | (~w24901 & w45430) | (w45429 & w45430);
assign w25253 = ~w20000 & w24083;
assign w25254 = (w24901 & w45431) | (w24901 & w45432) | (w45431 & w45432);
assign w25255 = ~w25252 & ~w25254;
assign w25256 = w19040 & w25255;
assign w25257 = ~w25241 & ~w25246;
assign w25258 = w25250 & w25257;
assign w25259 = ~w25256 & ~w25258;
assign w25260 = ~w18183 & w25101;
assign w25261 = ~w25103 & ~w25238;
assign w25262 = ~w25238 & ~w25260;
assign w25263 = ~w25259 & w25262;
assign w25264 = ~w25261 & ~w25263;
assign w25265 = ~w24221 & ~w24251;
assign w25266 = (w24247 & w24150) | (w24247 & w45433) | (w24150 & w45433);
assign w25267 = (~w24198 & w25266) | (~w24198 & w47696) | (w25266 & w47696);
assign w25268 = ~w24252 & ~w25267;
assign w25269 = ~w24209 & ~w25268;
assign w25270 = w25265 & ~w25269;
assign w25271 = ~w25265 & w25269;
assign w25272 = ~w25270 & ~w25271;
assign w25273 = ~w24901 & w45434;
assign w25274 = (w25272 & w24901) | (w25272 & w47697) | (w24901 & w47697);
assign w25275 = ~w25273 & ~w25274;
assign w25276 = ~w14039 & ~w25275;
assign w25277 = ~w15681 & w25267;
assign w25278 = w15681 & ~w25267;
assign w25279 = ~w25277 & ~w25278;
assign w25280 = ~w24208 & w25279;
assign w25281 = w24874 & w25280;
assign w25282 = (~w24901 & w45435) | (~w24901 & w45436) | (w45435 & w45436);
assign w25283 = ~w25281 & ~w25282;
assign w25284 = w14766 & w25283;
assign w25285 = ~w25276 & ~w25284;
assign w25286 = ~w24248 & ~w25266;
assign w25287 = ~w16559 & w25286;
assign w25288 = w16559 & ~w25286;
assign w25289 = ~w25287 & ~w25288;
assign w25290 = (~w24901 & w45437) | (~w24901 & w45438) | (w45437 & w45438);
assign w25291 = (w24901 & w45439) | (w24901 & w45440) | (w45439 & w45440);
assign w25292 = ~w25290 & ~w25291;
assign w25293 = ~w15681 & w25292;
assign w25294 = ~w14766 & ~w25283;
assign w25295 = ~w25293 & ~w25294;
assign w25296 = w15681 & ~w25292;
assign w25297 = ~w24179 & w24246;
assign w25298 = ~w17380 & w25297;
assign w25299 = w24232 & ~w25298;
assign w25300 = (~w25299 & w24901) | (~w25299 & w42130) | (w24901 & w42130);
assign w25301 = w24874 & w25286;
assign w25302 = w25300 & ~w25301;
assign w25303 = w24233 & ~w25297;
assign w25304 = w24248 & ~w25297;
assign w25305 = (~w25303 & w24873) | (~w25303 & w47698) | (w24873 & w47698);
assign w25306 = ~w25302 & w25305;
assign w25307 = ~w25302 & w42132;
assign w25308 = ~w25296 & w25307;
assign w25309 = w25295 & ~w25308;
assign w25310 = w25285 & ~w25309;
assign w25311 = ~w25264 & ~w25310;
assign w25312 = (w16559 & w25302) | (w16559 & w47699) | (w25302 & w47699);
assign w25313 = ~w25296 & ~w25312;
assign w25314 = w25295 & ~w25313;
assign w25315 = w25285 & ~w25314;
assign w25316 = (w25315 & ~w25237) | (w25315 & w42133) | (~w25237 & w42133);
assign w25317 = ~w25274 & w45441;
assign w25318 = ~w13384 & w24962;
assign w25319 = ~w24963 & ~w25318;
assign w25320 = ~w25317 & w25319;
assign w25321 = ~w13384 & w25317;
assign w25322 = ~w24957 & ~w25321;
assign w25323 = w24962 & ~w24964;
assign w25324 = (w25323 & ~w25319) | (w25323 & w47700) | (~w25319 & w47700);
assign w25325 = w25322 & ~w25324;
assign w25326 = ~w24949 & w25325;
assign w25327 = w25079 & w25326;
assign w25328 = ~w25316 & w25327;
assign w25329 = ~w25080 & ~w25328;
assign w25330 = ~w24288 & ~w24331;
assign w25331 = ~w24498 & ~w24571;
assign w25332 = w24035 & ~w25331;
assign w25333 = ~w24260 & w25332;
assign w25334 = (~w24343 & w24577) | (~w24343 & w49083) | (w24577 & w49083);
assign w25335 = (~w24424 & w24478) | (~w24424 & w49084) | (w24478 & w49084);
assign w25336 = w24499 & ~w25335;
assign w25337 = ~w24554 & w25336;
assign w25338 = ~w24395 & w25334;
assign w25339 = w25337 & ~w25338;
assign w25340 = (w25339 & w24260) | (w25339 & w45442) | (w24260 & w45442);
assign w25341 = (w25334 & ~w24567) | (w25334 & w25338) | (~w24567 & w25338);
assign w25342 = (~w25333 & w45443) | (~w25333 & w45444) | (w45443 & w45444);
assign w25343 = (w25333 & w45445) | (w25333 & w45446) | (w45445 & w45446);
assign w25344 = ~w25342 & ~w25343;
assign w25345 = ~w24287 & ~w24874;
assign w25346 = w24874 & ~w25344;
assign w25347 = ~w25345 & ~w25346;
assign w25348 = ~w2006 & w25347;
assign w25349 = ~w24901 & w42135;
assign w25350 = ~w24356 & ~w24394;
assign w25351 = ~w24356 & w52343;
assign w25352 = ~w24343 & ~w24347;
assign w25353 = (~w24342 & w24873) | (~w24342 & w42137) | (w24873 & w42137);
assign w25354 = (w24706 & w49085) | (w24706 & w49086) | (w49085 & w49086);
assign w25355 = w24874 & w25354;
assign w25356 = ~w25353 & ~w25355;
assign w25357 = w25351 & w25352;
assign w25358 = ~w25349 & w25357;
assign w25359 = w25356 & ~w25358;
assign w25360 = (w2285 & ~w25356) | (w2285 & w42138) | (~w25356 & w42138);
assign w25361 = w2006 & ~w25347;
assign w25362 = ~w25360 & ~w25361;
assign w25363 = ~w25348 & ~w25362;
assign w25364 = ~w24280 & ~w24281;
assign w25365 = ~w24279 & ~w24874;
assign w25366 = ~w25364 & w50212;
assign w25367 = (w25340 & w49087) | (w25340 & w49088) | (w49087 & w49088);
assign w25368 = ~w25366 & ~w25367;
assign w25369 = ~w25365 & w25368;
assign w25370 = ~w24901 & w49089;
assign w25371 = ~w25369 & w49090;
assign w25372 = ~w24290 & ~w24396;
assign w25373 = ~w24572 & w24896;
assign w25374 = ~w24705 & w45447;
assign w25375 = (w24706 & w45448) | (w24706 & w45449) | (w45448 & w45449);
assign w25376 = (~w24706 & w45450) | (~w24706 & w45451) | (w45450 & w45451);
assign w25377 = ~w25375 & ~w25376;
assign w25378 = w24874 & w25377;
assign w25379 = (~w24326 & w24901) | (~w24326 & w42140) | (w24901 & w42140);
assign w25380 = (w1541 & ~w25379) | (w1541 & w49091) | (~w25379 & w49091);
assign w25381 = w24326 & ~w25378;
assign w25382 = w25380 & ~w25381;
assign w25383 = ~w25371 & ~w25382;
assign w25384 = ~w25363 & w25383;
assign w25385 = (~w24299 & w24862) | (~w24299 & w49092) | (w24862 & w49092);
assign w25386 = ~w24327 & w25372;
assign w25387 = ~w24585 & ~w24586;
assign w25388 = (w25387 & w25374) | (w25387 & w42141) | (w25374 & w42141);
assign w25389 = ~w24873 & w45452;
assign w25390 = (~w24298 & w24873) | (~w24298 & w42142) | (w24873 & w42142);
assign w25391 = ~w25389 & ~w25390;
assign w25392 = ~w24901 & w42143;
assign w25393 = ~w24299 & ~w24586;
assign w25394 = (~w24585 & w25374) | (~w24585 & w42144) | (w25374 & w42144);
assign w25395 = ~w25393 & ~w25394;
assign w25396 = ~w25392 & w25395;
assign w25397 = ~w25391 & ~w25396;
assign w25398 = (w1120 & w25391) | (w1120 & w42145) | (w25391 & w42145);
assign w25399 = (w24872 & w49093) | (w24872 & w49094) | (w49093 & w49094);
assign w25400 = ~w25389 & ~w25399;
assign w25401 = ~w24600 & w24758;
assign w25402 = w945 & ~w25401;
assign w25403 = (w25402 & w25389) | (w25402 & w42147) | (w25389 & w42147);
assign w25404 = w945 & w25401;
assign w25405 = ~w25389 & w42148;
assign w25406 = ~w25403 & ~w25405;
assign w25407 = ~w25398 & w25406;
assign w25408 = ~w1541 & w24326;
assign w25409 = ~w25378 & w25408;
assign w25410 = w25379 & w45453;
assign w25411 = ~w25409 & ~w25410;
assign w25412 = ~w24896 & w25386;
assign w25413 = ~w24581 & ~w25412;
assign w25414 = w25337 & w25386;
assign w25415 = ~w25333 & w25414;
assign w25416 = w25413 & ~w25415;
assign w25417 = w24874 & w25416;
assign w25418 = ~w24313 & ~w24583;
assign w25419 = ~w1320 & ~w25418;
assign w25420 = ~w25417 & w42150;
assign w25421 = ~w1320 & w25418;
assign w25422 = (w25421 & w25417) | (w25421 & w42151) | (w25417 & w42151);
assign w25423 = ~w25420 & ~w25422;
assign w25424 = w25411 & w25423;
assign w25425 = w25407 & w25424;
assign w25426 = (~w1738 & w25369) | (~w1738 & w49095) | (w25369 & w49095);
assign w25427 = ~w25382 & w25426;
assign w25428 = w25425 & ~w25427;
assign w25429 = ~w25384 & w25428;
assign w25430 = ~w1120 & w25397;
assign w25431 = ~w25417 & w42152;
assign w25432 = (w25418 & w25417) | (w25418 & w42153) | (w25417 & w42153);
assign w25433 = ~w25431 & ~w25432;
assign w25434 = w1320 & w25433;
assign w25435 = ~w25430 & ~w25434;
assign w25436 = w25407 & ~w25435;
assign w25437 = w24648 & w24753;
assign w25438 = ~w24557 & w24867;
assign w25439 = w24758 & ~w24895;
assign w25440 = w25437 & w52255;
assign w25441 = ~w25437 & ~w52255;
assign w25442 = w24642 & ~w24643;
assign w25443 = ~w24642 & w24643;
assign w25444 = ~w25442 & ~w25443;
assign w25445 = ~w24874 & w25444;
assign w25446 = ~w25440 & ~w25441;
assign w25447 = w24874 & w25446;
assign w25448 = ~w25445 & ~w25447;
assign w25449 = w754 & w25448;
assign w25450 = (~w25401 & w25389) | (~w25401 & w49096) | (w25389 & w49096);
assign w25451 = ~w945 & ~w25450;
assign w25452 = w25400 & w25401;
assign w25453 = w25451 & ~w25452;
assign w25454 = ~w25449 & ~w25453;
assign w25455 = ~w25436 & w25454;
assign w25456 = ~w25429 & w25455;
assign w25457 = ~w24498 & ~w24554;
assign w25458 = w24476 & w25457;
assign w25459 = w24436 & w24459;
assign w25460 = w25458 & w25459;
assign w25461 = ~w24562 & ~w25459;
assign w25462 = (w25461 & w25333) | (w25461 & w42155) | (w25333 & w42155);
assign w25463 = w24562 & w25459;
assign w25464 = (~w25463 & w25333) | (~w25463 & w42156) | (w25333 & w42156);
assign w25465 = ~w25462 & w25464;
assign w25466 = w23843 & w24427;
assign w25467 = w22870 & ~w25466;
assign w25468 = ~w22870 & w25466;
assign w25469 = ~w25467 & ~w25468;
assign w25470 = w24874 & w25465;
assign w25471 = (w25469 & w24873) | (w25469 & w42157) | (w24873 & w42157);
assign w25472 = (w4838 & w25470) | (w4838 & w42158) | (w25470 & w42158);
assign w25473 = w24436 & ~w24865;
assign w25474 = ~w24873 & w25473;
assign w25475 = w24459 & w25458;
assign w25476 = (~w24563 & w25333) | (~w24563 & w42159) | (w25333 & w42159);
assign w25477 = ~w24873 & w45454;
assign w25478 = w24449 & w24483;
assign w25479 = ~w4430 & ~w25478;
assign w25480 = w4838 & w25479;
assign w25481 = ~w24865 & w25479;
assign w25482 = (~w25480 & w24873) | (~w25480 & w42160) | (w24873 & w42160);
assign w25483 = ~w4430 & w25478;
assign w25484 = w25476 & w25483;
assign w25485 = w25474 & w25484;
assign w25486 = ~w4838 & w25483;
assign w25487 = (w25486 & w24873) | (w25486 & w42161) | (w24873 & w42161);
assign w25488 = ~w25485 & ~w25487;
assign w25489 = ~w25477 & ~w25482;
assign w25490 = w25488 & ~w25489;
assign w25491 = ~w25472 & w25490;
assign w25492 = ~w25333 & w25457;
assign w25493 = (w24561 & ~w24874) | (w24561 & w42162) | (~w24874 & w42162);
assign w25494 = ~w24562 & ~w25331;
assign w25495 = (~w25494 & w42163) | (~w25494 & w25333) | (w42163 & w25333);
assign w25496 = (w42164 & w24260) | (w42164 & w47701) | (w24260 & w47701);
assign w25497 = ~w25495 & ~w25496;
assign w25498 = w24874 & ~w25497;
assign w25499 = (~w5330 & ~w24874) | (~w5330 & w42165) | (~w24874 & w42165);
assign w25500 = ~w25493 & w25499;
assign w25501 = ~w24517 & ~w24570;
assign w25502 = ~w24553 & w25501;
assign w25503 = (~w25502 & w24260) | (~w25502 & w42167) | (w24260 & w42167);
assign w25504 = ~w6264 & ~w25503;
assign w25505 = (w25504 & w24901) | (w25504 & w42168) | (w24901 & w42168);
assign w25506 = (w6264 & w24862) | (w6264 & w42169) | (w24862 & w42169);
assign w25507 = w25503 & w25506;
assign w25508 = ~w5745 & w24497;
assign w25509 = (w25508 & w24873) | (w25508 & w42170) | (w24873 & w42170);
assign w25510 = ~w25505 & w25509;
assign w25511 = ~w25504 & ~w25507;
assign w25512 = ~w5745 & ~w24497;
assign w25513 = w24874 & w42171;
assign w25514 = ~w25510 & ~w25513;
assign w25515 = ~w25500 & ~w25514;
assign w25516 = w5330 & w24561;
assign w25517 = (w25516 & ~w24874) | (w25516 & w42172) | (~w24874 & w42172);
assign w25518 = w24874 & w47702;
assign w25519 = ~w25517 & ~w25518;
assign w25520 = ~w25470 & w42173;
assign w25521 = w25519 & ~w25520;
assign w25522 = ~w25515 & w25521;
assign w25523 = w25491 & ~w25522;
assign w25524 = ~w24705 & w45455;
assign w25525 = ~w24356 & ~w24358;
assign w25526 = w24371 & ~w24576;
assign w25527 = ~w25525 & w25526;
assign w25528 = w24393 & ~w25524;
assign w25529 = w25527 & ~w25528;
assign w25530 = ~w24901 & w42174;
assign w25531 = w25529 & ~w25530;
assign w25532 = w25525 & ~w25526;
assign w25533 = w24393 & w25525;
assign w25534 = (w25533 & ~w24706) | (w25533 & w42175) | (~w24706 & w42175);
assign w25535 = ~w25532 & ~w25534;
assign w25536 = (w24355 & w24873) | (w24355 & w42176) | (w24873 & w42176);
assign w25537 = w24874 & ~w25535;
assign w25538 = ~w25536 & ~w25537;
assign w25539 = ~w25531 & w25538;
assign w25540 = (~w2558 & ~w25538) | (~w2558 & w42177) | (~w25538 & w42177);
assign w25541 = (w24706 & w45456) | (w24706 & w45457) | (w45456 & w45457);
assign w25542 = w24371 & w24392;
assign w25543 = w2896 & w25542;
assign w25544 = w2896 & ~w25542;
assign w25545 = w25541 & ~w25544;
assign w25546 = w24874 & ~w25545;
assign w25547 = ~w25541 & ~w25543;
assign w25548 = w25546 & ~w25547;
assign w25549 = (w3646 & ~w24706) | (w3646 & w42179) | (~w24706 & w42179);
assign w25550 = ~w3646 & w24573;
assign w25551 = w24706 & w25550;
assign w25552 = ~w25549 & ~w25551;
assign w25553 = ~w3242 & ~w24386;
assign w25554 = (w25553 & ~w24874) | (w25553 & w42180) | (~w24874 & w42180);
assign w25555 = w3242 & w25543;
assign w25556 = ~w3242 & w25544;
assign w25557 = ~w25555 & ~w25556;
assign w25558 = (~w25557 & w24873) | (~w25557 & w42181) | (w24873 & w42181);
assign w25559 = ~w3242 & w24386;
assign w25560 = (w25559 & ~w24706) | (w25559 & w42182) | (~w24706 & w42182);
assign w25561 = ~w25549 & w25560;
assign w25562 = w24874 & w25561;
assign w25563 = ~w25558 & ~w25562;
assign w25564 = ~w25554 & w25563;
assign w25565 = ~w25548 & w25564;
assign w25566 = ~w25540 & w25565;
assign w25567 = (~w4838 & w24873) | (~w4838 & w42183) | (w24873 & w42183);
assign w25568 = ~w25477 & ~w25567;
assign w25569 = w4430 & ~w25478;
assign w25570 = (w25569 & w25477) | (w25569 & w42184) | (w25477 & w42184);
assign w25571 = w4430 & w25478;
assign w25572 = ~w25477 & w42185;
assign w25573 = ~w25570 & ~w25572;
assign w25574 = ~w25331 & ~w25457;
assign w25575 = ~w24424 & w24564;
assign w25576 = w24490 & w25575;
assign w25577 = ~w25574 & w25576;
assign w25578 = ~w24418 & ~w24492;
assign w25579 = ~w25335 & ~w25575;
assign w25580 = w25578 & ~w25579;
assign w25581 = ~w25578 & w25579;
assign w25582 = ~w25580 & ~w25581;
assign w25583 = ~w25333 & w42186;
assign w25584 = (w25582 & w25333) | (w25582 & w42187) | (w25333 & w42187);
assign w25585 = ~w25583 & ~w25584;
assign w25586 = (w24417 & w24873) | (w24417 & w42188) | (w24873 & w42188);
assign w25587 = w24874 & w25585;
assign w25588 = ~w25586 & ~w25587;
assign w25589 = ~w25587 & w42189;
assign w25590 = ~w24478 & w24483;
assign w25591 = ~w24564 & w25590;
assign w25592 = w25457 & w25590;
assign w25593 = (~w25591 & w42190) | (~w25591 & w25333) | (w42190 & w25333);
assign w25594 = ~w24424 & w24488;
assign w25595 = (~w25594 & w24862) | (~w25594 & w47703) | (w24862 & w47703);
assign w25596 = (w25593 & w25009) | (w25593 & w42191) | (w25009 & w42191);
assign w25597 = (w25594 & w24862) | (w25594 & w47704) | (w24862 & w47704);
assign w25598 = ~w25593 & ~w25597;
assign w25599 = (w4056 & ~w24872) | (w4056 & w45458) | (~w24872 & w45458);
assign w25600 = ~w25598 & w25599;
assign w25601 = ~w25596 & w25600;
assign w25602 = (w24423 & w24873) | (w24423 & w42192) | (w24873 & w42192);
assign w25603 = (w24873 & w47705) | (w24873 & w47706) | (w47705 & w47706);
assign w25604 = ~w25601 & ~w25603;
assign w25605 = ~w25589 & w25604;
assign w25606 = w25573 & w25605;
assign w25607 = (w3646 & w25587) | (w3646 & w42193) | (w25587 & w42193);
assign w25608 = ~w24873 & ~w25598;
assign w25609 = ~w25596 & w25608;
assign w25610 = ~w4056 & ~w25602;
assign w25611 = ~w25609 & w25610;
assign w25612 = ~w25607 & ~w25611;
assign w25613 = (~w25589 & w25611) | (~w25589 & w47707) | (w25611 & w47707);
assign w25614 = w25566 & w25606;
assign w25615 = ~w25523 & w25614;
assign w25616 = w25566 & w25613;
assign w25617 = ~w25615 & ~w25616;
assign w25618 = (~w24386 & ~w24874) | (~w24386 & w42194) | (~w24874 & w42194);
assign w25619 = w24874 & w42195;
assign w25620 = ~w25618 & ~w25619;
assign w25621 = w3242 & w25620;
assign w25622 = w24874 & ~w25541;
assign w25623 = ~w2896 & w25542;
assign w25624 = ~w25622 & w42197;
assign w25625 = ~w2896 & ~w25542;
assign w25626 = (w25625 & w25622) | (w25625 & w42198) | (w25622 & w42198);
assign w25627 = ~w25624 & ~w25626;
assign w25628 = ~w25621 & w25627;
assign w25629 = ~w25548 & ~w25558;
assign w25630 = ~w25540 & w25629;
assign w25631 = ~w25628 & w25630;
assign w25632 = w2558 & w25539;
assign w25633 = (~w25632 & w25628) | (~w25632 & w47708) | (w25628 & w47708);
assign w25634 = w25356 & w42199;
assign w25635 = ~w25348 & ~w25634;
assign w25636 = ~w25426 & w25635;
assign w25637 = w25425 & w25636;
assign w25638 = w25633 & w25637;
assign w25639 = w25617 & w25638;
assign w25640 = w25456 & ~w25639;
assign w25641 = ~w24769 & w24783;
assign w25642 = ~w23862 & w52256;
assign w25643 = w24784 & w24874;
assign w25644 = ~w25642 & ~w25643;
assign w25645 = (w23863 & w24901) | (w23863 & w45459) | (w24901 & w45459);
assign w25646 = (w23862 & w24873) | (w23862 & w45460) | (w24873 & w45460);
assign w25647 = ~w25645 & ~w25646;
assign w25648 = (w3 & ~w25647) | (w3 & w49097) | (~w25647 & w49097);
assign w25649 = w25641 & ~w25644;
assign w25650 = w25648 & ~w25649;
assign w25651 = (~w3 & w24769) | (~w3 & w49098) | (w24769 & w49098);
assign w25652 = w25647 & w25651;
assign w25653 = ~w24769 & w49099;
assign w25654 = ~w25644 & w25653;
assign w25655 = ~w25652 & ~w25654;
assign w25656 = (w24766 & w24574) | (w24766 & w45461) | (w24574 & w45461);
assign w25657 = w24556 & w24766;
assign w25658 = ~w24261 & w25657;
assign w25659 = ~w25656 & ~w25658;
assign w25660 = w24774 & ~w24779;
assign w25661 = w24724 & ~w24778;
assign w25662 = ~w24734 & w25661;
assign w25663 = (w25662 & ~w25659) | (w25662 & w42202) | (~w25659 & w42202);
assign w25664 = ~w24901 & w42203;
assign w25665 = w25663 & ~w25664;
assign w25666 = ~w24777 & ~w24874;
assign w25667 = ~w25665 & ~w25666;
assign w25668 = ~w24873 & w42204;
assign w25669 = (~w24734 & ~w25659) | (~w24734 & w42205) | (~w25659 & w42205);
assign w25670 = (w80 & ~w25667) | (w80 & w45462) | (~w25667 & w45462);
assign w25671 = w25655 & ~w25670;
assign w25672 = ~w25650 & ~w25671;
assign w25673 = (w24765 & ~w24706) | (w24765 & w45463) | (~w24706 & w45463);
assign w25674 = ~w24702 & w25673;
assign w25675 = ~w24748 & w24774;
assign w25676 = ~w24865 & ~w25675;
assign w25677 = ~w24873 & w25676;
assign w25678 = ~w25674 & w25677;
assign w25679 = ~w24865 & w25675;
assign w25680 = ~w24873 & w25679;
assign w25681 = w25674 & w25680;
assign w25682 = ~w25678 & ~w25681;
assign w25683 = (~w24747 & w24873) | (~w24747 & w42206) | (w24873 & w42206);
assign w25684 = w252 & ~w25683;
assign w25685 = w25682 & w25684;
assign w25686 = ~w24734 & ~w24779;
assign w25687 = w24774 & w25659;
assign w25688 = w24874 & w25687;
assign w25689 = ~w25688 & w42208;
assign w25690 = (~w25686 & w25688) | (~w25686 & w42209) | (w25688 & w42209);
assign w25691 = ~w25689 & ~w25690;
assign w25692 = (~w57 & ~w25682) | (~w57 & w42210) | (~w25682 & w42210);
assign w25693 = w25691 & ~w25692;
assign w25694 = (~w80 & ~w25668) | (~w80 & w45464) | (~w25668 & w45464);
assign w25695 = w25667 & w25694;
assign w25696 = w25682 & ~w25683;
assign w25697 = w25682 & w42211;
assign w25698 = ~w25695 & ~w25697;
assign w25699 = ~w25693 & w25698;
assign w25700 = ~w25650 & w25699;
assign w25701 = ~w25672 & ~w25700;
assign w25702 = ~w252 & ~w25696;
assign w25703 = ~w25689 & w50347;
assign w25704 = (w57 & w25689) | (w57 & w50348) | (w25689 & w50348);
assign w25705 = ~w25703 & ~w25704;
assign w25706 = ~w25702 & ~w25705;
assign w25707 = ~w25672 & w25706;
assign w25708 = ~w24691 & ~w24874;
assign w25709 = ~w24692 & ~w24764;
assign w25710 = w24691 & ~w24864;
assign w25711 = w24706 & w42212;
assign w25712 = ~w24675 & ~w24696;
assign w25713 = (w25712 & ~w42213) | (w25712 & w45465) | (~w42213 & w45465);
assign w25714 = (w25709 & w24901) | (w25709 & w49100) | (w24901 & w49100);
assign w25715 = w25713 & w25714;
assign w25716 = ~w25709 & ~w25710;
assign w25717 = ~w25713 & w25716;
assign w25718 = ~w25715 & ~w25717;
assign w25719 = ~w25708 & w25718;
assign w25720 = ~w351 & ~w25719;
assign w25721 = (~w24667 & w24901) | (~w24667 & w42214) | (w24901 & w42214);
assign w25722 = w24662 & w24759;
assign w25723 = (w25722 & w24574) | (w25722 & w45466) | (w24574 & w45466);
assign w25724 = w24397 & w42215;
assign w25725 = ~w24261 & w25724;
assign w25726 = ~w25723 & ~w25725;
assign w25727 = ~w24663 & w24672;
assign w25728 = (w25727 & w25726) | (w25727 & w42216) | (w25726 & w42216);
assign w25729 = w24632 & ~w24667;
assign w25730 = ~w24901 & w45467;
assign w25731 = (~w25729 & w24901) | (~w25729 & w42217) | (w24901 & w42217);
assign w25732 = w25728 & w25731;
assign w25733 = ~w25730 & ~w25732;
assign w25734 = w25721 & w47709;
assign w25735 = w25733 & ~w25734;
assign w25736 = w25733 & w47710;
assign w25737 = w493 & ~w24871;
assign w25738 = ~w24901 & w25737;
assign w25739 = ~w25721 & ~w25738;
assign w25740 = (w24632 & w24901) | (w24632 & w42218) | (w24901 & w42218);
assign w25741 = ~w25728 & w25740;
assign w25742 = ~w25739 & ~w25741;
assign w25743 = w24624 & ~w24696;
assign w25744 = w400 & ~w25743;
assign w25745 = ~w25742 & w25744;
assign w25746 = w400 & w25743;
assign w25747 = w25742 & w25746;
assign w25748 = ~w25745 & ~w25747;
assign w25749 = ~w25736 & w25748;
assign w25750 = w24656 & ~w24657;
assign w25751 = ~w24656 & w24657;
assign w25752 = ~w25750 & ~w25751;
assign w25753 = w24662 & w24672;
assign w25754 = w24648 & ~w24759;
assign w25755 = ~w24556 & w24866;
assign w25756 = ~w24261 & ~w25755;
assign w25757 = ~w24867 & w24899;
assign w25758 = w24648 & ~w25757;
assign w25759 = (w25758 & w45468) | (w25758 & w45469) | (w45468 & w45469);
assign w25760 = w25753 & ~w25754;
assign w25761 = (w25760 & ~w25758) | (w25760 & w42220) | (~w25758 & w42220);
assign w25762 = ~w24874 & w25752;
assign w25763 = ~w25761 & ~w25762;
assign w25764 = ~w24901 & w45470;
assign w25765 = (~w25764 & ~w25763) | (~w25764 & w42221) | (~w25763 & w42221);
assign w25766 = w612 & w25765;
assign w25767 = (w493 & ~w25733) | (w493 & w47711) | (~w25733 & w47711);
assign w25768 = ~w25766 & ~w25767;
assign w25769 = w25749 & ~w25768;
assign w25770 = w351 & ~w25708;
assign w25771 = ~w25715 & w45471;
assign w25772 = ~w400 & w25743;
assign w25773 = ~w25742 & w25772;
assign w25774 = ~w400 & ~w25743;
assign w25775 = w25742 & w25774;
assign w25776 = ~w25773 & ~w25775;
assign w25777 = ~w25771 & w25776;
assign w25778 = ~w25769 & w25777;
assign w25779 = (~w25720 & w25769) | (~w25720 & w45472) | (w25769 & w45472);
assign w25780 = w25707 & ~w25779;
assign w25781 = ~w25701 & ~w25780;
assign w25782 = w25640 & ~w25781;
assign w25783 = ~w754 & ~w25448;
assign w25784 = ~w612 & ~w25765;
assign w25785 = ~w25783 & ~w25784;
assign w25786 = w25749 & w25785;
assign w25787 = w25749 & w49101;
assign w25788 = ~w25456 & w25787;
assign w25789 = (~w6264 & w25073) | (~w6264 & w45473) | (w25073 & w45473);
assign w25790 = w24874 & w42222;
assign w25791 = (w24497 & w24873) | (w24497 & w45474) | (w24873 & w45474);
assign w25792 = ~w25505 & w25791;
assign w25793 = ~w25790 & ~w25792;
assign w25794 = ~w25792 & w42223;
assign w25795 = ~w25789 & ~w25794;
assign w25796 = ~w25794 & w45475;
assign w25797 = w25491 & w25612;
assign w25798 = w25796 & w25797;
assign w25799 = (~w25798 & w25615) | (~w25798 & w42224) | (w25615 & w42224);
assign w25800 = w25638 & w25787;
assign w25801 = ~w25799 & w25800;
assign w25802 = ~w25788 & ~w25801;
assign w25803 = (~w25701 & ~w25802) | (~w25701 & w25781) | (~w25802 & w25781);
assign w25804 = ~w25329 & w25782;
assign w25805 = w25803 & ~w25804;
assign w25806 = w24885 & w25805;
assign w25807 = (w24769 & w50007) | (w24769 & w50008) | (w50007 & w50008);
assign w25808 = w24851 & ~w25807;
assign w25809 = ~w24851 & w25807;
assign w25810 = ~w25808 & ~w25809;
assign w25811 = ~w24852 & ~w25810;
assign w25812 = ~w24885 & ~w25805;
assign w25813 = w25811 & w25812;
assign w25814 = ~w25806 & ~w25813;
assign w25815 = ~w42 & w25814;
assign w25816 = (~w42 & ~w24884) | (~w42 & w50009) | (~w24884 & w50009);
assign w25817 = ~w25650 & w25655;
assign w25818 = w25237 & w42225;
assign w25819 = ~w25315 & w25326;
assign w25820 = w25056 & ~w25819;
assign w25821 = ~w25818 & w25820;
assign w25822 = ~w25615 & w42226;
assign w25823 = w25079 & ~w25822;
assign w25824 = w25456 & w25823;
assign w25825 = ~w25821 & w25824;
assign w25826 = ~w3 & w24821;
assign w25827 = (w24769 & w50010) | (w24769 & w50011) | (w50010 & w50011);
assign w25828 = ~w3 & w24851;
assign w25829 = ~w24821 & ~w25828;
assign w25830 = ~w24878 & ~w25829;
assign w25831 = ~w25827 & w25830;
assign w25832 = ~w25809 & ~w25831;
assign w25833 = ~w24885 & ~w25832;
assign w25834 = ~w42 & w25811;
assign w25835 = w42 & ~w25831;
assign w25836 = (w25835 & w24885) | (w25835 & w50012) | (w24885 & w50012);
assign w25837 = ~w25834 & ~w25836;
assign w25838 = w25650 & ~w25816;
assign w25839 = w25699 & ~w25838;
assign w25840 = w25837 & w25839;
assign w25841 = (w25840 & w25801) | (w25840 & w47712) | (w25801 & w47712);
assign w25842 = ~w25825 & w25841;
assign w25843 = ~w25700 & w45476;
assign w25844 = w25837 & ~w25843;
assign w25845 = w25720 & ~w25816;
assign w25846 = w25776 & w50013;
assign w25847 = (~w25845 & w25769) | (~w25845 & w50014) | (w25769 & w50014);
assign w25848 = ~w25701 & ~w25707;
assign w25849 = ~w25847 & ~w25848;
assign w25850 = w25844 & ~w25849;
assign w25851 = ~w25842 & ~w25850;
assign w25852 = w25573 & w25604;
assign w25853 = ~w25522 & w25797;
assign w25854 = w25612 & ~w25852;
assign w25855 = ~w25853 & ~w25854;
assign w25856 = w25823 & w25855;
assign w25857 = ~w25821 & w25856;
assign w25858 = (w25801 & w25821) | (w25801 & w45477) | (w25821 & w45477);
assign w25859 = (~w25779 & w25456) | (~w25779 & w45478) | (w25456 & w45478);
assign w25860 = w25706 & w25859;
assign w25861 = (w25699 & w25858) | (w25699 & w49104) | (w25858 & w49104);
assign w25862 = w3 & ~w25851;
assign w25863 = ~w25842 & w45479;
assign w25864 = ~w25861 & w25863;
assign w25865 = ~w25862 & ~w25864;
assign w25866 = w25817 & ~w25865;
assign w25867 = ~w25817 & w25865;
assign w25868 = ~w25866 & ~w25867;
assign w25869 = (~w25833 & ~w25805) | (~w25833 & w49105) | (~w25805 & w49105);
assign w25870 = w42 & ~w25869;
assign w25871 = ~w25812 & ~w25870;
assign w25872 = ~w25816 & ~w25871;
assign w25873 = ~w25868 & w25872;
assign w25874 = ~w25815 & ~w25873;
assign w25875 = ~w25693 & ~w25697;
assign w25876 = ~w25860 & w25875;
assign w25877 = w25801 & w25875;
assign w25878 = ~w25857 & w25877;
assign w25879 = ~w25876 & ~w25878;
assign w25880 = (w80 & w25842) | (w80 & w45480) | (w25842 & w45480);
assign w25881 = w25851 & ~w25879;
assign w25882 = ~w25670 & ~w25695;
assign w25883 = w3 & ~w25882;
assign w25884 = ~w25881 & w45481;
assign w25885 = w3 & w25882;
assign w25886 = (w25885 & w25881) | (w25885 & w45482) | (w25881 & w45482);
assign w25887 = ~w25884 & ~w25886;
assign w25888 = ~w25685 & ~w25850;
assign w25889 = ~w25842 & w25888;
assign w25890 = ~w25702 & w25859;
assign w25891 = ~w25858 & w25890;
assign w25892 = w25889 & ~w25891;
assign w25893 = (~w57 & w25842) | (~w57 & w45483) | (w25842 & w45483);
assign w25894 = ~w80 & ~w25705;
assign w25895 = (w25894 & w25892) | (w25894 & w45484) | (w25892 & w45484);
assign w25896 = ~w80 & w25705;
assign w25897 = ~w25892 & w45485;
assign w25898 = ~w25895 & ~w25897;
assign w25899 = w25887 & w25898;
assign w25900 = (~w25783 & w25429) | (~w25783 & w45486) | (w25429 & w45486);
assign w25901 = ~w25639 & ~w25900;
assign w25902 = ~w25329 & w25901;
assign w25903 = w25638 & ~w25799;
assign w25904 = (w25786 & w25903) | (w25786 & w45487) | (w25903 & w45487);
assign w25905 = (w25904 & w25329) | (w25904 & w49106) | (w25329 & w49106);
assign w25906 = ~w252 & w25696;
assign w25907 = ~w25720 & w25906;
assign w25908 = w25778 & ~w25905;
assign w25909 = w25907 & ~w25908;
assign w25910 = w25696 & ~w25851;
assign w25911 = ~w25909 & ~w25910;
assign w25912 = w252 & ~w25696;
assign w25913 = ~w25906 & ~w25912;
assign w25914 = w25778 & ~w25913;
assign w25915 = ~w25905 & w25914;
assign w25916 = w25858 & ~w25912;
assign w25917 = w25720 & ~w25913;
assign w25918 = (~w25917 & w25849) | (~w25917 & w45488) | (w25849 & w45488);
assign w25919 = ~w25859 & ~w25912;
assign w25920 = w25918 & ~w25919;
assign w25921 = ~w25842 & w25920;
assign w25922 = ~w25916 & w25921;
assign w25923 = ~w25915 & w25922;
assign w25924 = (~w57 & ~w25922) | (~w57 & w45489) | (~w25922 & w45489);
assign w25925 = w25911 & w25924;
assign w25926 = w80 & w25705;
assign w25927 = (w25926 & w25892) | (w25926 & w45490) | (w25892 & w45490);
assign w25928 = w80 & ~w25705;
assign w25929 = ~w25892 & w45491;
assign w25930 = ~w25927 & ~w25929;
assign w25931 = ~w25925 & w25930;
assign w25932 = ~w3 & ~w25882;
assign w25933 = (w25932 & w25881) | (w25932 & w45492) | (w25881 & w45492);
assign w25934 = ~w3 & w25882;
assign w25935 = ~w25881 & w45493;
assign w25936 = ~w25933 & ~w25935;
assign w25937 = ~w42 & w25817;
assign w25938 = ~w25865 & w25937;
assign w25939 = w25936 & ~w25938;
assign w25940 = ~w42 & ~w25817;
assign w25941 = w25865 & w25940;
assign w25942 = w25939 & ~w25941;
assign w25943 = w25899 & ~w25931;
assign w25944 = w25942 & ~w25943;
assign w25945 = ~w25874 & ~w25944;
assign w25946 = w25911 & ~w25923;
assign w25947 = w57 & ~w25946;
assign w25948 = w25638 & ~w25783;
assign w25949 = ~w25799 & w25948;
assign w25950 = ~w25900 & ~w25949;
assign w25951 = ~w25842 & w45494;
assign w25952 = ~w25902 & ~w25950;
assign w25953 = ~w25851 & w25952;
assign w25954 = ~w25951 & ~w25953;
assign w25955 = ~w25639 & w49108;
assign w25956 = ~w25329 & w25955;
assign w25957 = (~w25765 & w25949) | (~w25765 & w49107) | (w25949 & w49107);
assign w25958 = ~w25902 & w25957;
assign w25959 = ~w25949 & w49108;
assign w25960 = ~w25956 & ~w25959;
assign w25961 = ~w25958 & w25960;
assign w25962 = ~w493 & ~w25961;
assign w25963 = ~w25954 & w25962;
assign w25964 = ~w493 & w25961;
assign w25965 = w25954 & w25964;
assign w25966 = ~w25963 & ~w25965;
assign w25967 = (~w25784 & w25949) | (~w25784 & w45495) | (w25949 & w45495);
assign w25968 = (~w25766 & w25902) | (~w25766 & w49109) | (w25902 & w49109);
assign w25969 = ~w25736 & ~w25767;
assign w25970 = ~w25842 & w45496;
assign w25971 = w25768 & ~w25967;
assign w25972 = w25768 & w25901;
assign w25973 = ~w25329 & w25972;
assign w25974 = ~w25971 & ~w25973;
assign w25975 = ~w25736 & ~w25850;
assign w25976 = ~w25842 & w25975;
assign w25977 = (~w25735 & w25842) | (~w25735 & w45497) | (w25842 & w45497);
assign w25978 = ~w25974 & w25976;
assign w25979 = ~w25977 & ~w25978;
assign w25980 = ~w25968 & w25970;
assign w25981 = w25979 & w45498;
assign w25982 = w25966 & ~w25981;
assign w25983 = w493 & ~w25961;
assign w25984 = w25954 & w25983;
assign w25985 = w493 & w25961;
assign w25986 = ~w25954 & w25985;
assign w25987 = ~w25984 & ~w25986;
assign w25988 = ~w25436 & ~w25453;
assign w25989 = ~w25429 & w25988;
assign w25990 = ~w25903 & w25989;
assign w25991 = ~w25617 & w25989;
assign w25992 = ~w25329 & w25991;
assign w25993 = ~w25990 & ~w25992;
assign w25994 = ~w25449 & ~w25783;
assign w25995 = ~w25850 & ~w25994;
assign w25996 = ~w25842 & w25995;
assign w25997 = (~w25448 & w25842) | (~w25448 & w45499) | (w25842 & w45499);
assign w25998 = ~w25993 & w25996;
assign w25999 = ~w25997 & ~w25998;
assign w26000 = w25851 & w45500;
assign w26001 = w25999 & ~w26000;
assign w26002 = w25999 & w45501;
assign w26003 = w25987 & ~w26002;
assign w26004 = w25742 & ~w25743;
assign w26005 = ~w25742 & w25743;
assign w26006 = ~w26004 & ~w26005;
assign w26007 = (w25776 & w25849) | (w25776 & w49110) | (w25849 & w49110);
assign w26008 = ~w25842 & w26007;
assign w26009 = (~w26006 & w25842) | (~w26006 & w45502) | (w25842 & w45502);
assign w26010 = ~w25842 & w45503;
assign w26011 = ~w26009 & ~w26010;
assign w26012 = w25974 & w25976;
assign w26013 = ~w25769 & ~w25904;
assign w26014 = ~w25769 & w25901;
assign w26015 = ~w25329 & w26014;
assign w26016 = ~w26013 & ~w26015;
assign w26017 = (~w26006 & w25842) | (~w26006 & w45504) | (w25842 & w45504);
assign w26018 = w26016 & ~w26017;
assign w26019 = w26011 & ~w26012;
assign w26020 = ~w26018 & ~w26019;
assign w26021 = w351 & w26020;
assign w26022 = (~w400 & ~w25979) | (~w400 & w45505) | (~w25979 & w45505);
assign w26023 = (~w351 & w25842) | (~w351 & w49111) | (w25842 & w49111);
assign w26024 = w26008 & ~w26016;
assign w26025 = ~w25720 & ~w25771;
assign w26026 = ~w252 & w26025;
assign w26027 = (w26026 & w26024) | (w26026 & w49112) | (w26024 & w49112);
assign w26028 = ~w252 & ~w26025;
assign w26029 = ~w26024 & w49113;
assign w26030 = ~w26027 & ~w26029;
assign w26031 = ~w26022 & w26030;
assign w26032 = ~w26021 & w26031;
assign w26033 = w25982 & ~w26003;
assign w26034 = w26032 & ~w26033;
assign w26035 = ~w351 & w26018;
assign w26036 = (~w351 & ~w25976) | (~w351 & w45506) | (~w25976 & w45506);
assign w26037 = w26011 & w26036;
assign w26038 = ~w26035 & ~w26037;
assign w26039 = w252 & ~w26025;
assign w26040 = (w26039 & w26024) | (w26039 & w49114) | (w26024 & w49114);
assign w26041 = w252 & w26025;
assign w26042 = ~w26024 & w49115;
assign w26043 = ~w26040 & ~w26042;
assign w26044 = w26038 & w26043;
assign w26045 = w26030 & ~w26044;
assign w26046 = (~w25947 & w26044) | (~w25947 & w45507) | (w26044 & w45507);
assign w26047 = ~w26034 & w26046;
assign w26048 = ~w612 & ~w26001;
assign w26049 = w25406 & ~w25453;
assign w26050 = w25411 & ~w25427;
assign w26051 = w25633 & ~w25799;
assign w26052 = w25635 & w26050;
assign w26053 = ~w25384 & w26050;
assign w26054 = w25423 & ~w25434;
assign w26055 = (~w25857 & w50015) | (~w25857 & w50016) | (w50015 & w50016);
assign w26056 = w945 & w25435;
assign w26057 = (~w26056 & w25842) | (~w26056 & w45509) | (w25842 & w45509);
assign w26058 = w945 & ~w25851;
assign w26059 = ~w25842 & w45510;
assign w26060 = ~w26058 & ~w26059;
assign w26061 = ~w26055 & ~w26057;
assign w26062 = (w26049 & ~w26060) | (w26049 & w45511) | (~w26060 & w45511);
assign w26063 = w26060 & w45512;
assign w26064 = ~w26062 & ~w26063;
assign w26065 = ~w754 & w26064;
assign w26066 = ~w26048 & ~w26065;
assign w26067 = w25982 & w26044;
assign w26068 = w25982 & w49666;
assign w26069 = w26066 & w26068;
assign w26070 = ~w26047 & ~w26069;
assign w26071 = ~w25899 & w25936;
assign w26072 = ~w25874 & ~w26071;
assign w26073 = (~w25945 & w26070) | (~w25945 & w45513) | (w26070 & w45513);
assign w26074 = ~w25945 & ~w26047;
assign w26075 = w25815 & ~w25868;
assign w26076 = ~w26072 & ~w26075;
assign w26077 = ~w26074 & ~w26076;
assign w26078 = w26073 & ~w26077;
assign w26079 = (~w24971 & ~w25326) | (~w24971 & w45514) | (~w25326 & w45514);
assign w26080 = ~w25818 & w26079;
assign w26081 = w9781 & ~w26080;
assign w26082 = ~w9781 & w26080;
assign w26083 = ~w26081 & ~w26082;
assign w26084 = (w25050 & ~w25851) | (w25050 & w45515) | (~w25851 & w45515);
assign w26085 = w25851 & w45516;
assign w26086 = ~w26084 & ~w26085;
assign w26087 = w9195 & ~w26086;
assign w26088 = ~w24917 & ~w24921;
assign w26089 = ~w9781 & w26088;
assign w26090 = (~w26089 & w25842) | (~w26089 & w45517) | (w25842 & w45517);
assign w26091 = ~w24945 & w25325;
assign w26092 = ~w24906 & ~w24930;
assign w26093 = ~w24966 & ~w24968;
assign w26094 = ~w24945 & ~w26093;
assign w26095 = w26092 & ~w26094;
assign w26096 = (w26095 & w25316) | (w26095 & w50017) | (w25316 & w50017);
assign w26097 = ~w24923 & w24928;
assign w26098 = w24930 & ~w26097;
assign w26099 = ~w24930 & w26097;
assign w26100 = ~w26098 & ~w26099;
assign w26101 = w26096 & ~w26097;
assign w26102 = ~w26096 & ~w26100;
assign w26103 = ~w26101 & ~w26102;
assign w26104 = w25851 & ~w26103;
assign w26105 = ~w26090 & ~w26104;
assign w26106 = (~w26094 & w25316) | (~w26094 & w50018) | (w25316 & w50018);
assign w26107 = ~w10419 & w26096;
assign w26108 = ~w10419 & ~w26092;
assign w26109 = ~w26106 & w26108;
assign w26110 = ~w26107 & ~w26109;
assign w26111 = ~w10419 & w24929;
assign w26112 = (w26111 & w25842) | (w26111 & w45518) | (w25842 & w45518);
assign w26113 = w25851 & ~w26110;
assign w26114 = ~w26112 & ~w26113;
assign w26115 = ~w26105 & w26114;
assign w26116 = ~w25316 & w25320;
assign w26117 = w12666 & w24963;
assign w26118 = ~w12666 & ~w24963;
assign w26119 = ~w26117 & ~w26118;
assign w26120 = ~w26116 & w26119;
assign w26121 = ~w12666 & w25320;
assign w26122 = ~w25316 & w26121;
assign w26123 = ~w25850 & ~w26122;
assign w26124 = ~w26120 & w26123;
assign w26125 = (w24956 & ~w26124) | (w24956 & w49116) | (~w26124 & w49116);
assign w26126 = w26124 & w49117;
assign w26127 = ~w26125 & ~w26126;
assign w26128 = w11870 & w26127;
assign w26129 = w11870 & w50213;
assign w26130 = (w25316 & w50019) | (w25316 & w50020) | (w50019 & w50020);
assign w26131 = ~w26129 & ~w26130;
assign w26132 = w25851 & ~w26131;
assign w26133 = w11138 & ~w24967;
assign w26134 = (w26133 & ~w25851) | (w26133 & w45519) | (~w25851 & w45519);
assign w26135 = w11138 & w24967;
assign w26136 = w25851 & w45520;
assign w26137 = ~w26134 & ~w26136;
assign w26138 = w26128 & w26137;
assign w26139 = ~w11138 & w24967;
assign w26140 = (w26139 & ~w25851) | (w26139 & w45521) | (~w25851 & w45521);
assign w26141 = ~w11138 & ~w24967;
assign w26142 = w25851 & w45522;
assign w26143 = ~w26140 & ~w26142;
assign w26144 = ~w26092 & ~w26106;
assign w26145 = ~w26096 & ~w26144;
assign w26146 = (w24929 & w25842) | (w24929 & w45523) | (w25842 & w45523);
assign w26147 = w25851 & ~w26145;
assign w26148 = ~w26146 & ~w26147;
assign w26149 = ~w26147 & w45524;
assign w26150 = w26143 & ~w26149;
assign w26151 = ~w26138 & w26150;
assign w26152 = (w26115 & w26138) | (w26115 & w45525) | (w26138 & w45525);
assign w26153 = ~w25851 & ~w26088;
assign w26154 = ~w26104 & ~w26153;
assign w26155 = w9781 & ~w26154;
assign w26156 = ~w9195 & w26086;
assign w26157 = ~w26155 & ~w26156;
assign w26158 = ~w11870 & ~w26127;
assign w26159 = w26137 & ~w26158;
assign w26160 = ~w25316 & ~w25317;
assign w26161 = ~w25850 & ~w26160;
assign w26162 = w25839 & w50021;
assign w26163 = (w26162 & w25801) | (w26162 & w49119) | (w25801 & w49119);
assign w26164 = ~w25825 & w26163;
assign w26165 = ~w25849 & w50022;
assign w26166 = ~w26164 & ~w26165;
assign w26167 = ~w25842 & w26161;
assign w26168 = w26166 & ~w26167;
assign w26169 = ~w12666 & w25319;
assign w26170 = ~w26168 & w26169;
assign w26171 = ~w12666 & ~w25319;
assign w26172 = w26168 & w26171;
assign w26173 = ~w26170 & ~w26172;
assign w26174 = w26115 & w26173;
assign w26175 = w26159 & w26174;
assign w26176 = w26157 & ~w26175;
assign w26177 = (~w26087 & ~w26176) | (~w26087 & w45526) | (~w26176 & w45526);
assign w26178 = ~w25039 & ~w25058;
assign w26179 = ~w25005 & ~w25024;
assign w26180 = w26178 & w26179;
assign w26181 = w25053 & w26180;
assign w26182 = ~w25818 & w45527;
assign w26183 = ~w25005 & ~w25059;
assign w26184 = ~w25021 & ~w25062;
assign w26185 = w26183 & ~w26184;
assign w26186 = ~w26183 & w26184;
assign w26187 = ~w26185 & ~w26186;
assign w26188 = w26182 & w26187;
assign w26189 = ~w26182 & ~w26187;
assign w26190 = ~w26188 & ~w26189;
assign w26191 = (w25020 & w25842) | (w25020 & w45528) | (w25842 & w45528);
assign w26192 = w25851 & w26190;
assign w26193 = ~w26191 & ~w26192;
assign w26194 = w7315 & w26193;
assign w26195 = ~w24994 & ~w25061;
assign w26196 = w25022 & ~w25054;
assign w26197 = (w45529 & w50349) | (w45529 & w50350) | (w50349 & w50350);
assign w26198 = ~w26195 & ~w26197;
assign w26199 = w26195 & w26197;
assign w26200 = w25851 & w50024;
assign w26201 = ~w24993 & ~w25851;
assign w26202 = ~w6769 & ~w26201;
assign w26203 = ~w26200 & w26202;
assign w26204 = ~w26194 & ~w26203;
assign w26205 = ~w25039 & ~w25053;
assign w26206 = w26179 & w26205;
assign w26207 = (~w26206 & w25849) | (~w26206 & w45530) | (w25849 & w45530);
assign w26208 = (w26180 & w25818) | (w26180 & w45531) | (w25818 & w45531);
assign w26209 = w26207 & ~w26208;
assign w26210 = ~w25842 & w26209;
assign w26211 = ~w8666 & w25004;
assign w26212 = w25839 & w50025;
assign w26213 = (w26212 & w25801) | (w26212 & w49120) | (w25801 & w49120);
assign w26214 = ~w25825 & w26213;
assign w26215 = ~w25849 & w50026;
assign w26216 = (w26178 & w25818) | (w26178 & w45532) | (w25818 & w45532);
assign w26217 = ~w26179 & ~w26205;
assign w26218 = (w26217 & w25849) | (w26217 & w45533) | (w25849 & w45533);
assign w26219 = ~w26216 & w26218;
assign w26220 = w25839 & w50027;
assign w26221 = (w26220 & w25801) | (w26220 & w49121) | (w25801 & w49121);
assign w26222 = ~w25825 & w26221;
assign w26223 = ~w25849 & w50028;
assign w26224 = ~w26222 & ~w26223;
assign w26225 = ~w25842 & w26219;
assign w26226 = w26224 & ~w26225;
assign w26227 = ~w26214 & ~w26215;
assign w26228 = ~w26210 & w26227;
assign w26229 = w26226 & ~w26228;
assign w26230 = ~w7924 & w26229;
assign w26231 = (~w7315 & w26192) | (~w7315 & w45534) | (w26192 & w45534);
assign w26232 = (~w26231 & ~w26229) | (~w26231 & w47713) | (~w26229 & w47713);
assign w26233 = w7924 & ~w26229;
assign w26234 = ~w26205 & ~w26216;
assign w26235 = ~w25051 & ~w25057;
assign w26236 = (w26235 & w25818) | (w26235 & w45535) | (w25818 & w45535);
assign w26237 = ~w9195 & w25051;
assign w26238 = w9195 & ~w25051;
assign w26239 = ~w26237 & ~w26238;
assign w26240 = ~w9195 & w26236;
assign w26241 = ~w26236 & ~w26239;
assign w26242 = ~w26240 & ~w26241;
assign w26243 = w25851 & ~w26242;
assign w26244 = ~w8666 & ~w25038;
assign w26245 = (w26244 & ~w25851) | (w26244 & w45536) | (~w25851 & w45536);
assign w26246 = ~w8666 & w26234;
assign w26247 = w25851 & w45537;
assign w26248 = ~w26245 & ~w26247;
assign w26249 = ~w26233 & ~w26248;
assign w26250 = w26232 & ~w26249;
assign w26251 = w26204 & ~w26250;
assign w26252 = ~w26200 & ~w26201;
assign w26253 = w6769 & ~w26252;
assign w26254 = ~w24987 & ~w25076;
assign w26255 = ~w24994 & ~w25063;
assign w26256 = ~w24994 & w26196;
assign w26257 = (w45529 & w50351) | (w45529 & w50352) | (w50351 & w50352);
assign w26258 = ~w26254 & w26257;
assign w26259 = w26254 & ~w26257;
assign w26260 = ~w25075 & ~w25851;
assign w26261 = ~w26258 & ~w26259;
assign w26262 = w25851 & w26261;
assign w26263 = ~w26260 & ~w26262;
assign w26264 = ~w6264 & w26263;
assign w26265 = ~w26253 & ~w26264;
assign w26266 = (w26265 & w26250) | (w26265 & w50030) | (w26250 & w50030);
assign w26267 = (w25319 & ~w26166) | (w25319 & w47714) | (~w26166 & w47714);
assign w26268 = w26166 & w47715;
assign w26269 = ~w26267 & ~w26268;
assign w26270 = w12666 & w26269;
assign w26271 = (w25313 & ~w25237) | (w25313 & w42227) | (~w25237 & w42227);
assign w26272 = w25295 & ~w26271;
assign w26273 = ~w25284 & ~w26272;
assign w26274 = (w14039 & w25842) | (w14039 & w45538) | (w25842 & w45538);
assign w26275 = ~w25842 & w45539;
assign w26276 = ~w26274 & ~w26275;
assign w26277 = ~w25276 & ~w25317;
assign w26278 = ~w13384 & ~w26277;
assign w26279 = ~w26276 & w26278;
assign w26280 = ~w13384 & w26277;
assign w26281 = w26276 & w26280;
assign w26282 = ~w26279 & ~w26281;
assign w26283 = ~w26270 & w26282;
assign w26284 = w26157 & w26283;
assign w26285 = ~w26152 & w26284;
assign w26286 = w26266 & ~w26285;
assign w26287 = w26177 & w26286;
assign w26288 = w8666 & ~w26234;
assign w26289 = w25851 & w45540;
assign w26290 = w8666 & w25038;
assign w26291 = (w26290 & ~w25851) | (w26290 & w45541) | (~w25851 & w45541);
assign w26292 = ~w26289 & ~w26291;
assign w26293 = ~w26233 & w26292;
assign w26294 = w26232 & ~w26293;
assign w26295 = w6264 & ~w26263;
assign w26296 = ~w25074 & ~w25789;
assign w26297 = ~w25064 & ~w25076;
assign w26298 = ~w25060 & w26297;
assign w26299 = ~w25821 & w26298;
assign w26300 = (w6264 & w25842) | (w6264 & w45542) | (w25842 & w45542);
assign w26301 = ~w25842 & w45543;
assign w26302 = ~w26300 & ~w26301;
assign w26303 = ~w26296 & w26302;
assign w26304 = ~w5745 & ~w26303;
assign w26305 = w26296 & ~w26302;
assign w26306 = w26304 & ~w26305;
assign w26307 = w25514 & ~w25794;
assign w26308 = (w26307 & w25328) | (w26307 & w50031) | (w25328 & w50031);
assign w26309 = ~w25328 & w50032;
assign w26310 = ~w26308 & ~w26309;
assign w26311 = (w25793 & w25842) | (w25793 & w50033) | (w25842 & w50033);
assign w26312 = w25851 & w26310;
assign w26313 = ~w26311 & ~w26312;
assign w26314 = ~w26312 & w50034;
assign w26315 = ~w26295 & ~w26306;
assign w26316 = ~w26314 & w26315;
assign w26317 = (w26265 & w26294) | (w26265 & w50030) | (w26294 & w50030);
assign w26318 = w26316 & ~w26317;
assign w26319 = ~w25554 & ~w25562;
assign w26320 = ~w25621 & w26319;
assign w26321 = ~w25853 & w42228;
assign w26322 = (w25798 & w25056) | (w25798 & w45544) | (w25056 & w45544);
assign w26323 = (w26321 & w25328) | (w26321 & w50035) | (w25328 & w50035);
assign w26324 = ~w26320 & ~w26323;
assign w26325 = ~w25853 & w45545;
assign w26326 = ~w26322 & w26325;
assign w26327 = w25327 & w26325;
assign w26328 = ~w25316 & w26327;
assign w26329 = ~w26326 & ~w26328;
assign w26330 = w25620 & ~w25851;
assign w26331 = w25851 & w50036;
assign w26332 = ~w26330 & ~w26331;
assign w26333 = ~w2896 & ~w26332;
assign w26334 = ~w25589 & ~w25607;
assign w26335 = (w25796 & w25056) | (w25796 & w45546) | (w25056 & w45546);
assign w26336 = w25491 & w26335;
assign w26337 = ~w25328 & w26336;
assign w26338 = ~w25523 & w25852;
assign w26339 = (~w25611 & w26337) | (~w25611 & w47717) | (w26337 & w47717);
assign w26340 = ~w26334 & ~w26339;
assign w26341 = w25851 & ~w26340;
assign w26342 = w26334 & w26339;
assign w26343 = w26341 & ~w26342;
assign w26344 = (w25588 & w25842) | (w25588 & w50037) | (w25842 & w50037);
assign w26345 = w3242 & ~w26344;
assign w26346 = ~w26343 & w26345;
assign w26347 = ~w25523 & w25573;
assign w26348 = (w4056 & w26337) | (w4056 & w47718) | (w26337 & w47718);
assign w26349 = ~w26337 & w47719;
assign w26350 = w25851 & w45547;
assign w26351 = ~w25602 & ~w25609;
assign w26352 = w3646 & ~w26351;
assign w26353 = w26350 & w26352;
assign w26354 = w3646 & w26351;
assign w26355 = ~w26350 & w26354;
assign w26356 = ~w26353 & ~w26355;
assign w26357 = ~w26346 & w26356;
assign w26358 = ~w26333 & w26357;
assign w26359 = w25478 & ~w25568;
assign w26360 = ~w25478 & w25568;
assign w26361 = ~w26359 & ~w26360;
assign w26362 = ~w25515 & w25519;
assign w26363 = ~w25472 & ~w25520;
assign w26364 = w26362 & w26363;
assign w26365 = w26335 & w26364;
assign w26366 = ~w25328 & w26365;
assign w26367 = ~w25472 & ~w25522;
assign w26368 = w25490 & w25573;
assign w26369 = w26367 & ~w26368;
assign w26370 = ~w26367 & w26368;
assign w26371 = ~w26369 & ~w26370;
assign w26372 = w26366 & ~w26371;
assign w26373 = ~w26366 & w26371;
assign w26374 = ~w26372 & ~w26373;
assign w26375 = (~w26361 & w25842) | (~w26361 & w45548) | (w25842 & w45548);
assign w26376 = w25851 & ~w26374;
assign w26377 = ~w26375 & ~w26376;
assign w26378 = (~w4056 & w26376) | (~w4056 & w45549) | (w26376 & w45549);
assign w26379 = ~w25328 & w26335;
assign w26380 = (w26362 & w25849) | (w26362 & w45550) | (w25849 & w45550);
assign w26381 = ~w26379 & w26380;
assign w26382 = ~w25842 & w26381;
assign w26383 = w4838 & w25840;
assign w26384 = (w26383 & w25801) | (w26383 & w49122) | (w25801 & w49122);
assign w26385 = ~w25825 & w26384;
assign w26386 = w4838 & w25850;
assign w26387 = ~w26385 & ~w26386;
assign w26388 = ~w26382 & w26387;
assign w26389 = ~w4430 & ~w26363;
assign w26390 = (w26389 & ~w26387) | (w26389 & w47720) | (~w26387 & w47720);
assign w26391 = ~w4430 & w26363;
assign w26392 = w26387 & w47721;
assign w26393 = ~w26390 & ~w26392;
assign w26394 = ~w26378 & w26393;
assign w26395 = (w25795 & w25056) | (w25795 & w45551) | (w25056 & w45551);
assign w26396 = (w25514 & w25328) | (w25514 & w49123) | (w25328 & w49123);
assign w26397 = ~w25493 & ~w25498;
assign w26398 = (w26397 & w25842) | (w26397 & w45552) | (w25842 & w45552);
assign w26399 = ~w25519 & w26396;
assign w26400 = w25851 & w26399;
assign w26401 = ~w26398 & ~w26400;
assign w26402 = ~w5330 & ~w26397;
assign w26403 = ~w26396 & w26402;
assign w26404 = w25851 & w26403;
assign w26405 = w5330 & w26397;
assign w26406 = ~w25514 & ~w26405;
assign w26407 = w26395 & ~w26405;
assign w26408 = ~w25328 & w26407;
assign w26409 = ~w26406 & ~w26408;
assign w26410 = ~w25500 & w25514;
assign w26411 = (w26410 & w25328) | (w26410 & w49124) | (w25328 & w49124);
assign w26412 = w26409 & ~w26411;
assign w26413 = (~w4838 & ~w26409) | (~w4838 & w49125) | (~w26409 & w49125);
assign w26414 = ~w26404 & w26413;
assign w26415 = w26401 & w26414;
assign w26416 = w4430 & w26363;
assign w26417 = (w26416 & ~w26387) | (w26416 & w47722) | (~w26387 & w47722);
assign w26418 = w4430 & ~w26363;
assign w26419 = w26387 & w47723;
assign w26420 = ~w26417 & ~w26419;
assign w26421 = ~w26415 & w26420;
assign w26422 = w26394 & ~w26421;
assign w26423 = ~w26376 & w45553;
assign w26424 = ~w3646 & w26351;
assign w26425 = w26350 & w26424;
assign w26426 = ~w3646 & ~w26351;
assign w26427 = ~w26350 & w26426;
assign w26428 = ~w26423 & ~w26427;
assign w26429 = ~w26425 & w26428;
assign w26430 = ~w26422 & w26429;
assign w26431 = w2896 & w26332;
assign w26432 = ~w26343 & ~w26344;
assign w26433 = ~w3242 & ~w26432;
assign w26434 = ~w26333 & w26433;
assign w26435 = ~w26431 & ~w26434;
assign w26436 = w26358 & ~w26430;
assign w26437 = w26435 & ~w26436;
assign w26438 = w26318 & w26437;
assign w26439 = ~w26287 & w26438;
assign w26440 = ~w25329 & w25640;
assign w26441 = (w25849 & w26440) | (w25849 & w49126) | (w26440 & w49126);
assign w26442 = ~a[26] & w24874;
assign w26443 = w25844 & w26442;
assign w26444 = ~w26441 & w26443;
assign w26445 = w23843 & w24874;
assign w26446 = ~w23843 & ~w24874;
assign w26447 = ~w26445 & ~w26446;
assign w26448 = w25213 & ~w26447;
assign w26449 = ~w25213 & w26447;
assign w26450 = ~w26448 & ~w26449;
assign w26451 = w25851 & ~w26450;
assign w26452 = ~w26444 & ~w26451;
assign w26453 = w25841 & ~w26440;
assign w26454 = (w25212 & w25849) | (w25212 & w49127) | (w25849 & w49127);
assign w26455 = ~a[26] & w26454;
assign w26456 = ~w26453 & w26455;
assign w26457 = (w26442 & w25842) | (w26442 & w45554) | (w25842 & w45554);
assign w26458 = ~w26456 & ~w26457;
assign w26459 = ~w25841 & ~w25850;
assign w26460 = w25640 & ~w25850;
assign w26461 = ~w25329 & w26460;
assign w26462 = ~w26459 & ~w26461;
assign w26463 = (w26461 & w49128) | (w26461 & w49129) | (w49128 & w49129);
assign w26464 = ~w26458 & ~w26463;
assign w26465 = w25851 & w26449;
assign w26466 = ~a[27] & ~w26452;
assign w26467 = a[27] & ~w26465;
assign w26468 = ~w26464 & w26467;
assign w26469 = ~w26466 & ~w26468;
assign w26470 = (w45556 & w25801) | (w45556 & w49130) | (w25801 & w49130);
assign w26471 = ~w26440 & w26470;
assign w26472 = a[26] & ~w26454;
assign w26473 = ~w26471 & ~w26472;
assign w26474 = (w24874 & w25842) | (w24874 & w45557) | (w25842 & w45557);
assign w26475 = ~w26473 & ~w26474;
assign w26476 = w26458 & ~w26475;
assign w26477 = a[24] & ~a[25];
assign w26478 = ~a[22] & ~a[23];
assign w26479 = ~a[24] & w26478;
assign w26480 = ~w24874 & ~w26479;
assign w26481 = w24874 & w26479;
assign w26482 = ~a[25] & ~w26481;
assign w26483 = ~w26480 & ~w26482;
assign w26484 = ~w26480 & ~w26481;
assign w26485 = ~a[25] & w26484;
assign w26486 = ~w26481 & ~w26485;
assign w26487 = ~w26477 & ~w26483;
assign w26488 = (w26487 & w26461) | (w26487 & w47724) | (w26461 & w47724);
assign w26489 = ~w26461 & w47725;
assign w26490 = ~w26488 & ~w26489;
assign w26491 = ~w23843 & ~w26490;
assign w26492 = w26476 & ~w26491;
assign w26493 = w23843 & w26483;
assign w26494 = w23843 & w26477;
assign w26495 = ~w25837 & w26494;
assign w26496 = (~w26495 & w45558) | (~w26495 & w26462) | (w45558 & w26462);
assign w26497 = w23843 & ~w26486;
assign w26498 = ~w26461 & w47726;
assign w26499 = ~w25816 & w26494;
assign w26500 = ~w25805 & w26499;
assign w26501 = ~w26498 & ~w26500;
assign w26502 = w26496 & w26501;
assign w26503 = w26501 & w45559;
assign w26504 = ~w26492 & w26503;
assign w26505 = w26469 & ~w26504;
assign w26506 = ~w25224 & ~w25225;
assign w26507 = ~w25842 & w45560;
assign w26508 = ~w21801 & ~w25231;
assign w26509 = ~w26507 & w26508;
assign w26510 = ~w21801 & w25231;
assign w26511 = w26507 & w26510;
assign w26512 = ~w26509 & ~w26511;
assign w26513 = ~w22767 & w26512;
assign w26514 = w26502 & w26512;
assign w26515 = ~w26492 & w26514;
assign w26516 = ~w26513 & ~w26515;
assign w26517 = ~w26505 & ~w26516;
assign w26518 = w25231 & ~w26507;
assign w26519 = ~w25231 & w26507;
assign w26520 = ~w26518 & ~w26519;
assign w26521 = w21801 & ~w26520;
assign w26522 = ~w21801 & ~w25233;
assign w26523 = w21801 & w25233;
assign w26524 = ~w26522 & ~w26523;
assign w26525 = ~w25850 & w26524;
assign w26526 = ~w25842 & w26525;
assign w26527 = w20906 & w25203;
assign w26528 = (w26527 & w25842) | (w26527 & w45561) | (w25842 & w45561);
assign w26529 = w20906 & ~w25203;
assign w26530 = ~w25842 & w45562;
assign w26531 = ~w26528 & ~w26530;
assign w26532 = ~w25211 & ~w25233;
assign w26533 = w25209 & ~w26532;
assign w26534 = ~w20000 & ~w26533;
assign w26535 = w20000 & w26533;
assign w26536 = ~w26534 & ~w26535;
assign w26537 = ~w25850 & w26536;
assign w26538 = ~w25842 & w26537;
assign w26539 = w24874 & w25111;
assign w26540 = w24083 & ~w25239;
assign w26541 = ~w26539 & ~w26540;
assign w26542 = w19040 & ~w26541;
assign w26543 = (w26542 & w25842) | (w26542 & w45563) | (w25842 & w45563);
assign w26544 = w19040 & w26541;
assign w26545 = ~w25842 & w45564;
assign w26546 = ~w26543 & ~w26545;
assign w26547 = ~w25154 & ~w25206;
assign w26548 = ~w25203 & ~w26522;
assign w26549 = ~w26523 & ~w26548;
assign w26550 = w26547 & ~w26549;
assign w26551 = ~w26547 & w26549;
assign w26552 = ~w26550 & ~w26551;
assign w26553 = w20000 & w25153;
assign w26554 = (w26553 & w25842) | (w26553 & w45565) | (w25842 & w45565);
assign w26555 = w20000 & w26552;
assign w26556 = ~w25842 & w45566;
assign w26557 = ~w26554 & ~w26556;
assign w26558 = w26546 & w26557;
assign w26559 = w25203 & ~w26526;
assign w26560 = ~w25203 & w26526;
assign w26561 = ~w26559 & ~w26560;
assign w26562 = ~w20906 & w26561;
assign w26563 = w26558 & ~w26562;
assign w26564 = w26521 & w26531;
assign w26565 = w26563 & ~w26564;
assign w26566 = ~w26517 & w26565;
assign w26567 = w25237 & w47727;
assign w26568 = (w16559 & ~w25237) | (w16559 & w47728) | (~w25237 & w47728);
assign w26569 = ~w26567 & ~w26568;
assign w26570 = (w25306 & w25842) | (w25306 & w45567) | (w25842 & w45567);
assign w26571 = ~w25842 & w45568;
assign w26572 = ~w26570 & ~w26571;
assign w26573 = ~w15681 & ~w26572;
assign w26574 = ~w25293 & ~w25296;
assign w26575 = (w25237 & w49131) | (w25237 & w49132) | (w49131 & w49132);
assign w26576 = w26574 & w52257;
assign w26577 = ~w26575 & ~w26576;
assign w26578 = (w25292 & w25842) | (w25292 & w45569) | (w25842 & w45569);
assign w26579 = ~w25842 & w45570;
assign w26580 = ~w26578 & ~w26579;
assign w26581 = ~w14766 & ~w26580;
assign w26582 = ~w26573 & ~w26581;
assign w26583 = ~w14766 & ~w25293;
assign w26584 = w14766 & w25293;
assign w26585 = ~w26583 & ~w26584;
assign w26586 = ~w26576 & w26585;
assign w26587 = w26271 & w26583;
assign w26588 = ~w25850 & w49133;
assign w26589 = (w25283 & ~w26588) | (w25283 & w47729) | (~w26588 & w47729);
assign w26590 = w26588 & w47730;
assign w26591 = ~w26589 & ~w26590;
assign w26592 = w14039 & w26591;
assign w26593 = w26582 & ~w26592;
assign w26594 = ~w20000 & ~w25153;
assign w26595 = (w26594 & w25842) | (w26594 & w45571) | (w25842 & w45571);
assign w26596 = ~w20000 & ~w26552;
assign w26597 = ~w25842 & w45572;
assign w26598 = ~w26595 & ~w26597;
assign w26599 = w26531 & w26598;
assign w26600 = w26558 & ~w26599;
assign w26601 = ~w26534 & ~w26541;
assign w26602 = ~w26535 & ~w26601;
assign w26603 = w19040 & ~w26602;
assign w26604 = ~w19040 & ~w26535;
assign w26605 = ~w26601 & w26604;
assign w26606 = ~w25850 & ~w26605;
assign w26607 = ~w26603 & w26606;
assign w26608 = w20000 & ~w25112;
assign w26609 = w25115 & ~w26608;
assign w26610 = w24142 & ~w26609;
assign w26611 = ~w24142 & w26609;
assign w26612 = ~w26610 & ~w26611;
assign w26613 = w26607 & w47731;
assign w26614 = (w26612 & ~w26607) | (w26612 & w47732) | (~w26607 & w47732);
assign w26615 = ~w26613 & ~w26614;
assign w26616 = (~w26541 & w25842) | (~w26541 & w45573) | (w25842 & w45573);
assign w26617 = ~w19040 & ~w26616;
assign w26618 = w26538 & w26541;
assign w26619 = w26617 & ~w26618;
assign w26620 = ~w18183 & w26615;
assign w26621 = ~w26619 & ~w26620;
assign w26622 = ~w26600 & w26621;
assign w26623 = ~w25259 & w26533;
assign w26624 = (w25128 & ~w26533) | (w25128 & w49134) | (~w26533 & w49134);
assign w26625 = w18183 & ~w25259;
assign w26626 = w25101 & ~w25128;
assign w26627 = w26625 & w26626;
assign w26628 = w25102 & w26624;
assign w26629 = (~w26627 & w25850) | (~w26627 & w45574) | (w25850 & w45574);
assign w26630 = w25840 & ~w26627;
assign w26631 = (w26630 & w25801) | (w26630 & w49135) | (w25801 & w49135);
assign w26632 = ~w25825 & w26631;
assign w26633 = w25101 & w25840;
assign w26634 = (w26633 & w25801) | (w26633 & w49136) | (w25801 & w49136);
assign w26635 = ~w25825 & w26634;
assign w26636 = w18183 & w26623;
assign w26637 = ~w18183 & w25128;
assign w26638 = ~w26623 & w26637;
assign w26639 = ~w26636 & ~w26638;
assign w26640 = (w25101 & w25850) | (w25101 & w45575) | (w25850 & w45575);
assign w26641 = ~w26635 & ~w26640;
assign w26642 = ~w26629 & ~w26632;
assign w26643 = w26641 & ~w26642;
assign w26644 = ~w25101 & ~w25128;
assign w26645 = ~w26625 & w26644;
assign w26646 = ~w25842 & w45576;
assign w26647 = ~w25102 & ~w25260;
assign w26648 = w26623 & w26647;
assign w26649 = ~w25850 & w26648;
assign w26650 = ~w26453 & w26649;
assign w26651 = ~w26646 & ~w26650;
assign w26652 = w26643 & w26651;
assign w26653 = (w17380 & ~w26651) | (w17380 & w49137) | (~w26651 & w49137);
assign w26654 = ~w25094 & ~w25238;
assign w26655 = ~w25259 & ~w25260;
assign w26656 = ~w26624 & w26655;
assign w26657 = ~w25102 & ~w26656;
assign w26658 = w26654 & ~w26657;
assign w26659 = ~w26654 & w26657;
assign w26660 = ~w26658 & ~w26659;
assign w26661 = (w25093 & w25842) | (w25093 & w45577) | (w25842 & w45577);
assign w26662 = w25851 & ~w26660;
assign w26663 = ~w26661 & ~w26662;
assign w26664 = (~w16559 & w26662) | (~w16559 & w45578) | (w26662 & w45578);
assign w26665 = (~w26664 & w26652) | (~w26664 & w47733) | (w26652 & w47733);
assign w26666 = w26622 & w26665;
assign w26667 = w26622 & w45579;
assign w26668 = (w26667 & w26517) | (w26667 & w45580) | (w26517 & w45580);
assign w26669 = ~w14766 & w26577;
assign w26670 = w15681 & ~w26669;
assign w26671 = w25851 & ~w26670;
assign w26672 = ~w17230 & ~w25296;
assign w26673 = (w26672 & w25842) | (w26672 & w45581) | (w25842 & w45581);
assign w26674 = ~w26671 & ~w26673;
assign w26675 = w26572 & w26674;
assign w26676 = w14766 & ~w25292;
assign w26677 = (w26676 & w25842) | (w26676 & w45582) | (w25842 & w45582);
assign w26678 = w14766 & ~w26577;
assign w26679 = ~w25842 & w45583;
assign w26680 = ~w26677 & ~w26679;
assign w26681 = ~w14039 & w25283;
assign w26682 = (w26681 & ~w26588) | (w26681 & w47734) | (~w26588 & w47734);
assign w26683 = ~w14039 & ~w25283;
assign w26684 = w26588 & w47735;
assign w26685 = ~w26682 & ~w26684;
assign w26686 = w26680 & w26685;
assign w26687 = ~w26675 & w26686;
assign w26688 = ~w26592 & ~w26687;
assign w26689 = w18183 & ~w26615;
assign w26690 = w16559 & w26663;
assign w26691 = ~w17380 & w26643;
assign w26692 = w26651 & w26691;
assign w26693 = w26691 & w47736;
assign w26694 = ~w26690 & ~w26693;
assign w26695 = ~w26664 & w26689;
assign w26696 = ~w26653 & w26695;
assign w26697 = w26694 & ~w26696;
assign w26698 = w26593 & ~w26697;
assign w26699 = (~w26688 & w26697) | (~w26688 & w50038) | (w26697 & w50038);
assign w26700 = ~w26668 & w26699;
assign w26701 = w26276 & ~w26277;
assign w26702 = ~w26276 & w26277;
assign w26703 = ~w26701 & ~w26702;
assign w26704 = w13384 & ~w26703;
assign w26705 = ~w26251 & w45584;
assign w26706 = w26177 & w26705;
assign w26707 = w26700 & w26706;
assign w26708 = w26439 & ~w26707;
assign w26709 = ~w26404 & ~w26412;
assign w26710 = w26401 & w26709;
assign w26711 = ~w5330 & ~w26313;
assign w26712 = w5745 & w26296;
assign w26713 = ~w26302 & w26712;
assign w26714 = w5745 & ~w26296;
assign w26715 = w26302 & w26714;
assign w26716 = ~w26713 & ~w26715;
assign w26717 = ~w26314 & ~w26716;
assign w26718 = ~w26711 & ~w26717;
assign w26719 = w4838 & ~w26710;
assign w26720 = w26718 & ~w26719;
assign w26721 = w26358 & w26394;
assign w26722 = w26720 & w26721;
assign w26723 = w26437 & ~w26722;
assign w26724 = w25635 & w52258;
assign w26725 = (~w25363 & w25849) | (~w25363 & w50039) | (w25849 & w50039);
assign w26726 = ~w25842 & w26725;
assign w26727 = ~w26724 & w26726;
assign w26728 = (~w1738 & w25842) | (~w1738 & w45586) | (w25842 & w45586);
assign w26729 = ~w25371 & ~w25426;
assign w26730 = ~w26727 & w45587;
assign w26731 = (w26729 & w26727) | (w26729 & w45588) | (w26727 & w45588);
assign w26732 = ~w26730 & ~w26731;
assign w26733 = ~w1541 & w26732;
assign w26734 = ~w25363 & ~w25371;
assign w26735 = ~w26724 & w26734;
assign w26736 = ~w25842 & w45589;
assign w26737 = ~w26735 & w26736;
assign w26738 = (w1541 & w25842) | (w1541 & w50040) | (w25842 & w50040);
assign w26739 = ~w25382 & w25411;
assign w26740 = ~w1320 & ~w26739;
assign w26741 = ~w26737 & w50041;
assign w26742 = ~w1320 & w26739;
assign w26743 = (w26742 & w26737) | (w26742 & w50042) | (w26737 & w50042);
assign w26744 = ~w26741 & ~w26743;
assign w26745 = ~w26733 & w26744;
assign w26746 = (w25857 & w50043) | (w25857 & w50044) | (w50043 & w50044);
assign w26747 = w25433 & ~w25851;
assign w26748 = ~w26055 & ~w26746;
assign w26749 = w25851 & w26748;
assign w26750 = ~w26747 & ~w26749;
assign w26751 = w1120 & w26750;
assign w26752 = (w1120 & w25842) | (w1120 & w50045) | (w25842 & w50045);
assign w26753 = ~w25842 & w45590;
assign w26754 = ~w26055 & w26753;
assign w26755 = ~w25398 & ~w25430;
assign w26756 = w945 & ~w26755;
assign w26757 = (w26756 & w26754) | (w26756 & w50046) | (w26754 & w50046);
assign w26758 = w945 & w26755;
assign w26759 = ~w26754 & w50047;
assign w26760 = ~w26757 & ~w26759;
assign w26761 = ~w26751 & w26760;
assign w26762 = w26745 & w26761;
assign w26763 = ~w25565 & w25627;
assign w26764 = ~w25853 & w45591;
assign w26765 = ~w25628 & ~w26763;
assign w26766 = (~w26763 & ~w25797) | (~w26763 & w45592) | (~w25797 & w45592);
assign w26767 = (~w26765 & ~w26321) | (~w26765 & w45593) | (~w26321 & w45593);
assign w26768 = w25080 & w26764;
assign w26769 = w26767 & ~w26768;
assign w26770 = w25327 & w26764;
assign w26771 = ~w25316 & w26770;
assign w26772 = w2558 & ~w25539;
assign w26773 = (w25540 & ~w26769) | (w25540 & w47737) | (~w26769 & w47737);
assign w26774 = w26769 & w47738;
assign w26775 = ~w26773 & ~w26774;
assign w26776 = w25851 & ~w26775;
assign w26777 = w26769 & w47739;
assign w26778 = (w2558 & ~w26769) | (w2558 & w47740) | (~w26769 & w47740);
assign w26779 = ~w26777 & ~w26778;
assign w26780 = w25851 & w26779;
assign w26781 = w25539 & ~w26780;
assign w26782 = ~w26776 & ~w26781;
assign w26783 = (~w2285 & w26781) | (~w2285 & w45594) | (w26781 & w45594);
assign w26784 = w25627 & w25629;
assign w26785 = (w2896 & w25842) | (w2896 & w45595) | (w25842 & w45595);
assign w26786 = (~w25621 & w25849) | (~w25621 & w45596) | (w25849 & w45596);
assign w26787 = w26329 & w26786;
assign w26788 = ~w25842 & w26787;
assign w26789 = ~w26785 & ~w26788;
assign w26790 = w26784 & ~w26789;
assign w26791 = ~w26784 & w26789;
assign w26792 = ~w26790 & ~w26791;
assign w26793 = w2558 & ~w26792;
assign w26794 = ~w26783 & ~w26793;
assign w26795 = ~w25360 & ~w25634;
assign w26796 = ~w26795 & w52258;
assign w26797 = w26795 & ~w52258;
assign w26798 = ~w26796 & ~w26797;
assign w26799 = w25851 & ~w26798;
assign w26800 = (~w25359 & w25842) | (~w25359 & w50353) | (w25842 & w50353);
assign w26801 = ~w2006 & ~w26800;
assign w26802 = ~w26799 & w26801;
assign w26803 = ~w2006 & ~w25360;
assign w26804 = (w26803 & w25615) | (w26803 & w42230) | (w25615 & w42230);
assign w26805 = w2006 & w25360;
assign w26806 = (~w26805 & ~w25080) | (~w26805 & w49138) | (~w25080 & w49138);
assign w26807 = w25633 & ~w25634;
assign w26808 = (w26803 & w25799) | (w26803 & w42231) | (w25799 & w42231);
assign w26809 = w25327 & w26804;
assign w26810 = ~w25316 & w26809;
assign w26811 = ~w26808 & ~w26810;
assign w26812 = ~w25850 & w26806;
assign w26813 = w26811 & w26812;
assign w26814 = ~w25842 & w26813;
assign w26815 = w2006 & ~w25634;
assign w26816 = ~w25857 & w42232;
assign w26817 = w26814 & ~w26816;
assign w26818 = ~w1738 & w25347;
assign w26819 = (w26818 & ~w26814) | (w26818 & w42233) | (~w26814 & w42233);
assign w26820 = ~w1738 & ~w25347;
assign w26821 = w26814 & w42234;
assign w26822 = ~w26819 & ~w26821;
assign w26823 = ~w26802 & w26822;
assign w26824 = w26794 & w26823;
assign w26825 = w26762 & w26824;
assign w26826 = (w26825 & ~w26437) | (w26825 & w45597) | (~w26437 & w45597);
assign w26827 = (w26826 & w26707) | (w26826 & w42235) | (w26707 & w42235);
assign w26828 = w1738 & ~w25347;
assign w26829 = (w26828 & ~w26814) | (w26828 & w42236) | (~w26814 & w42236);
assign w26830 = w1738 & w25347;
assign w26831 = w26814 & w42237;
assign w26832 = ~w26829 & ~w26831;
assign w26833 = (w26832 & w26802) | (w26832 & w42238) | (w26802 & w42238);
assign w26834 = w1541 & w26729;
assign w26835 = (w26834 & w26727) | (w26834 & w45598) | (w26727 & w45598);
assign w26836 = w1541 & ~w26729;
assign w26837 = ~w26727 & w45599;
assign w26838 = ~w26835 & ~w26837;
assign w26839 = w2285 & ~w26776;
assign w26840 = ~w26781 & w26839;
assign w26841 = ~w2558 & w26784;
assign w26842 = ~w26788 & w26841;
assign w26843 = ~w26785 & w26842;
assign w26844 = ~w2558 & ~w26784;
assign w26845 = w2896 & w26844;
assign w26846 = (w26845 & w25842) | (w26845 & w42239) | (w25842 & w42239);
assign w26847 = w26788 & w26844;
assign w26848 = ~w26846 & ~w26847;
assign w26849 = ~w26843 & w26848;
assign w26850 = ~w26840 & w26849;
assign w26851 = ~w26783 & ~w26850;
assign w26852 = (w25359 & w25842) | (w25359 & w42240) | (w25842 & w42240);
assign w26853 = w2006 & ~w26852;
assign w26854 = w25851 & w26798;
assign w26855 = w26853 & ~w26854;
assign w26856 = w26832 & ~w26855;
assign w26857 = (w49139 & w42238) | (w49139 & w50354) | (w42238 & w50354);
assign w26858 = w26838 & w26856;
assign w26859 = ~w26851 & w26858;
assign w26860 = ~w26857 & ~w26859;
assign w26861 = w26762 & w26860;
assign w26862 = (~w1120 & w26749) | (~w1120 & w42241) | (w26749 & w42241);
assign w26863 = w1320 & ~w26739;
assign w26864 = (w26863 & w26737) | (w26863 & w42242) | (w26737 & w42242);
assign w26865 = w1320 & w26739;
assign w26866 = ~w26737 & w42243;
assign w26867 = ~w26864 & ~w26866;
assign w26868 = ~w26862 & w26867;
assign w26869 = w26761 & ~w26868;
assign w26870 = ~w26754 & w42244;
assign w26871 = (w26755 & w26754) | (w26755 & w42245) | (w26754 & w42245);
assign w26872 = ~w26870 & ~w26871;
assign w26873 = ~w945 & ~w26872;
assign w26874 = w754 & ~w26064;
assign w26875 = ~w26873 & ~w26874;
assign w26876 = ~w26869 & w26875;
assign w26877 = ~w26861 & w26876;
assign w26878 = ~w26077 & w26877;
assign w26879 = (~w42235 & w47741) | (~w42235 & w47742) | (w47741 & w47742);
assign w26880 = (~w26078 & w26827) | (~w26078 & w45600) | (w26827 & w45600);
assign w26881 = (w25987 & w26880) | (w25987 & w50048) | (w26880 & w50048);
assign w26882 = (w26066 & w26861) | (w26066 & w45601) | (w26861 & w45601);
assign w26883 = w26439 & ~w26882;
assign w26884 = (w26066 & w26826) | (w26066 & w26882) | (w26826 & w26882);
assign w26885 = ~w26707 & w26883;
assign w26886 = (w26884 & ~w26883) | (w26884 & w45602) | (~w26883 & w45602);
assign w26887 = ~w26002 & ~w26886;
assign w26888 = ~w26881 & ~w26887;
assign w26889 = ~w26070 & w26826;
assign w26890 = w26826 & w42246;
assign w26891 = ~w26708 & w26890;
assign w26892 = ~w26070 & ~w26877;
assign w26893 = w26074 & ~w26892;
assign w26894 = (~w26076 & w26892) | (~w26076 & w26077) | (w26892 & w26077);
assign w26895 = (~w26894 & w26708) | (~w26894 & w42247) | (w26708 & w42247);
assign w26896 = (w26003 & w26885) | (w26003 & w42248) | (w26885 & w42248);
assign w26897 = ~w26880 & ~w26896;
assign w26898 = ~w25954 & ~w25961;
assign w26899 = w25954 & w25961;
assign w26900 = ~w26898 & ~w26899;
assign w26901 = ~w26897 & w26900;
assign w26902 = w26895 & w26896;
assign w26903 = w493 & w26902;
assign w26904 = ~w26901 & ~w26903;
assign w26905 = ~w26888 & w26904;
assign w26906 = w400 & w26905;
assign w26907 = (~w400 & ~w26904) | (~w400 & w50049) | (~w26904 & w50049);
assign w26908 = (~w45603 & w47743) | (~w45603 & w47744) | (w47743 & w47744);
assign w26909 = ~w26065 & w26877;
assign w26910 = w26909 & ~w26827;
assign w26911 = ~w26065 & ~w26910;
assign w26912 = ~w26908 & ~w26911;
assign w26913 = w26001 & ~w26073;
assign w26914 = ~w26002 & ~w26913;
assign w26915 = w26886 & w26914;
assign w26916 = ~w26078 & ~w26913;
assign w26917 = ~w26879 & w26916;
assign w26918 = ~w26915 & ~w26917;
assign w26919 = ~w26912 & w26918;
assign w26920 = ~w493 & ~w26919;
assign w26921 = ~w26917 & w45604;
assign w26922 = ~w26912 & w26921;
assign w26923 = ~w26065 & ~w26073;
assign w26924 = ~w26910 & ~w26923;
assign w26925 = w26064 & ~w26078;
assign w26926 = ~w26879 & w26925;
assign w26927 = ~w26924 & ~w26926;
assign w26928 = ~w26869 & ~w26873;
assign w26929 = ~w26861 & w26928;
assign w26930 = ~w26826 & w26929;
assign w26931 = w26439 & w26929;
assign w26932 = (~w26930 & ~w26931) | (~w26930 & w45605) | (~w26931 & w45605);
assign w26933 = w26874 & w26932;
assign w26934 = (w42249 & ~w26931) | (w42249 & w47745) | (~w26931 & w47745);
assign w26935 = w26895 & w26934;
assign w26936 = ~w26933 & ~w26935;
assign w26937 = ~w26927 & w26936;
assign w26938 = w612 & ~w26937;
assign w26939 = ~w26922 & ~w26938;
assign w26940 = ~w26920 & ~w26939;
assign w26941 = (~w26907 & w26939) | (~w26907 & w50050) | (w26939 & w50050);
assign w26942 = (w26824 & ~w26437) | (w26824 & w45606) | (~w26437 & w45606);
assign w26943 = (w26942 & w26707) | (w26942 & w42250) | (w26707 & w42250);
assign w26944 = ~w26688 & ~w26704;
assign w26945 = ~w26698 & w26944;
assign w26946 = w26285 & ~w26945;
assign w26947 = w26285 & w26667;
assign w26948 = ~w26566 & w26947;
assign w26949 = ~w26946 & ~w26948;
assign w26950 = w26251 & w26316;
assign w26951 = w26437 & w26950;
assign w26952 = w26437 & w52259;
assign w26953 = (w26949 & w50051) | (w26949 & w50052) | (w50051 & w50052);
assign w26954 = w26745 & w26860;
assign w26955 = w26867 & ~w26954;
assign w26956 = ~w26862 & w26955;
assign w26957 = (w26956 & ~w26943) | (w26956 & w50053) | (~w26943 & w50053);
assign w26958 = w26760 & ~w26873;
assign w26959 = (~w26958 & w26879) | (~w26958 & w45607) | (w26879 & w45607);
assign w26960 = ~w26751 & ~w26957;
assign w26961 = w26959 & ~w26960;
assign w26962 = w26761 & ~w26873;
assign w26963 = ~w26073 & w26889;
assign w26964 = ~w26708 & w26963;
assign w26965 = ~w26073 & ~w26893;
assign w26966 = ~w945 & w26962;
assign w26967 = (w26962 & w26893) | (w26962 & w45608) | (w26893 & w45608);
assign w26968 = ~w26964 & w26967;
assign w26969 = ~w26966 & ~w26968;
assign w26970 = w26872 & w26880;
assign w26971 = ~w26957 & ~w26969;
assign w26972 = ~w26970 & ~w26971;
assign w26973 = ~w26961 & w26972;
assign w26974 = (~w754 & ~w26972) | (~w754 & w42252) | (~w26972 & w42252);
assign w26975 = ~w612 & w26937;
assign w26976 = ~w26920 & ~w26975;
assign w26977 = ~w26974 & w26976;
assign w26978 = (~w26906 & ~w26941) | (~w26906 & w45609) | (~w26941 & w45609);
assign w26979 = (~w26750 & w26957) | (~w26750 & w45610) | (w26957 & w45610);
assign w26980 = ~w26751 & ~w26862;
assign w26981 = ~w26980 & w52260;
assign w26982 = ~w26077 & w50054;
assign w26983 = ~w26827 & w26982;
assign w26984 = ~w26981 & ~w26983;
assign w26985 = (w26955 & ~w26943) | (w26955 & w50055) | (~w26943 & w50055);
assign w26986 = ~w26984 & ~w26985;
assign w26987 = ~w26964 & ~w26965;
assign w26988 = ~w26964 & w42254;
assign w26989 = w26957 & w26988;
assign w26990 = ~w26986 & ~w26989;
assign w26991 = ~w26979 & w26990;
assign w26992 = (~w945 & ~w26990) | (~w945 & w45611) | (~w26990 & w45611);
assign w26993 = w26972 & w42255;
assign w26994 = ~w26992 & ~w26993;
assign w26995 = ~w26940 & w49140;
assign w26996 = (~w26860 & ~w26943) | (~w26860 & w50056) | (~w26943 & w50056);
assign w26997 = w1320 & w26880;
assign w26998 = ~w26880 & ~w26996;
assign w26999 = ~w26733 & w26998;
assign w27000 = ~w26997 & ~w26999;
assign w27001 = w26744 & w26867;
assign w27002 = ~w1120 & ~w27001;
assign w27003 = ~w27000 & w27002;
assign w27004 = ~w1120 & w27001;
assign w27005 = w27000 & w27004;
assign w27006 = ~w27003 & ~w27005;
assign w27007 = ~w26439 & ~w26723;
assign w27008 = w26706 & ~w26723;
assign w27009 = w26700 & w27008;
assign w27010 = ~w27007 & ~w27009;
assign w27011 = ~w26794 & ~w26840;
assign w27012 = ~w26951 & ~w27011;
assign w27013 = w26177 & ~w27011;
assign w27014 = w26949 & w27013;
assign w27015 = ~w27012 & ~w27014;
assign w27016 = ~w27010 & ~w27015;
assign w27017 = ~w26851 & ~w27016;
assign w27018 = ~w2006 & w26880;
assign w27019 = ~w26880 & w27017;
assign w27020 = ~w27018 & ~w27019;
assign w27021 = ~w26802 & ~w26855;
assign w27022 = w1738 & ~w27021;
assign w27023 = ~w27019 & w50057;
assign w27024 = w1738 & w27021;
assign w27025 = (w27024 & w27019) | (w27024 & w50058) | (w27019 & w50058);
assign w27026 = ~w27023 & ~w27025;
assign w27027 = (~w26855 & w26850) | (~w26855 & w50059) | (w26850 & w50059);
assign w27028 = ~w26802 & ~w27027;
assign w27029 = w1738 & w27028;
assign w27030 = w26439 & ~w27029;
assign w27031 = w1738 & ~w26802;
assign w27032 = (w26437 & w49141) | (w26437 & w49142) | (w49141 & w49142);
assign w27033 = w27031 & ~w27032;
assign w27034 = (w27033 & ~w27030) | (w27033 & w47746) | (~w27030 & w47746);
assign w27035 = ~w1738 & ~w27028;
assign w27036 = (w42257 & ~w26437) | (w42257 & w49143) | (~w26437 & w49143);
assign w27037 = w27035 & ~w27036;
assign w27038 = w26439 & w27035;
assign w27039 = (~w27037 & ~w27038) | (~w27037 & w47747) | (~w27038 & w47747);
assign w27040 = ~w27034 & w27039;
assign w27041 = ~w25347 & ~w26817;
assign w27042 = w25347 & w26817;
assign w27043 = ~w27041 & ~w27042;
assign w27044 = w1541 & w27043;
assign w27045 = w27040 & w45612;
assign w27046 = w1541 & ~w27043;
assign w27047 = ~w27040 & w27046;
assign w27048 = ~w26078 & w27046;
assign w27049 = ~w26879 & w27048;
assign w27050 = ~w27047 & ~w27049;
assign w27051 = ~w27045 & w27050;
assign w27052 = ~w26733 & w26838;
assign w27053 = ~w26851 & w26856;
assign w27054 = ~w26833 & ~w27053;
assign w27055 = w27052 & w27054;
assign w27056 = w26439 & ~w27055;
assign w27057 = (~w27054 & w26723) | (~w27054 & w42258) | (w26723 & w42258);
assign w27058 = w27052 & ~w27057;
assign w27059 = ~w26707 & w27056;
assign w27060 = w27058 & ~w27059;
assign w27061 = ~w27052 & ~w27054;
assign w27062 = ~w26942 & w27061;
assign w27063 = w26439 & w27061;
assign w27064 = (~w27062 & ~w27063) | (~w27062 & w45613) | (~w27063 & w45613);
assign w27065 = ~w27060 & w27064;
assign w27066 = w1320 & ~w26732;
assign w27067 = w26880 & w27066;
assign w27068 = ~w27060 & w45614;
assign w27069 = ~w26880 & w27068;
assign w27070 = ~w27067 & ~w27069;
assign w27071 = w27051 & w27070;
assign w27072 = ~w26793 & w26849;
assign w27073 = ~w27007 & w47748;
assign w27074 = w2285 & ~w26793;
assign w27075 = ~w2285 & w26793;
assign w27076 = ~w27074 & ~w27075;
assign w27077 = (w27076 & ~w27010) | (w27076 & w42259) | (~w27010 & w42259);
assign w27078 = w27010 & w42260;
assign w27079 = ~w27077 & ~w27078;
assign w27080 = w2006 & w26782;
assign w27081 = (w27080 & w27079) | (w27080 & w50060) | (w27079 & w50060);
assign w27082 = w2006 & ~w26782;
assign w27083 = ~w27079 & w50061;
assign w27084 = ~w27081 & ~w27083;
assign w27085 = w27071 & w27084;
assign w27086 = w27026 & w27085;
assign w27087 = w27006 & w27086;
assign w27088 = w26393 & ~w26421;
assign w27089 = w26393 & w26720;
assign w27090 = (w27089 & w26707) | (w27089 & w42261) | (w26707 & w42261);
assign w27091 = w4056 & ~w26377;
assign w27092 = ~w27090 & w47749;
assign w27093 = ~w26880 & w27092;
assign w27094 = ~w4056 & w26377;
assign w27095 = (w26423 & w27090) | (w26423 & w47750) | (w27090 & w47750);
assign w27096 = ~w27090 & w47751;
assign w27097 = ~w27095 & ~w27096;
assign w27098 = ~w27093 & w27097;
assign w27099 = (w26378 & w27090) | (w26378 & w47752) | (w27090 & w47752);
assign w27100 = ~w26880 & w27099;
assign w27101 = ~w26078 & w26377;
assign w27102 = ~w26879 & w27101;
assign w27103 = ~w27100 & ~w27102;
assign w27104 = w27098 & w27103;
assign w27105 = ~w3646 & ~w27104;
assign w27106 = (w3646 & w26879) | (w3646 & w45615) | (w26879 & w45615);
assign w27107 = ~w27100 & w27106;
assign w27108 = w27098 & w27107;
assign w27109 = w26393 & w26420;
assign w27110 = (w26720 & w26707) | (w26720 & w42262) | (w26707 & w42262);
assign w27111 = ~w26415 & ~w27110;
assign w27112 = (~w27109 & w27110) | (~w27109 & w47753) | (w27110 & w47753);
assign w27113 = ~w26880 & ~w27112;
assign w27114 = w26363 & ~w26388;
assign w27115 = ~w26363 & w26388;
assign w27116 = ~w27114 & ~w27115;
assign w27117 = ~w26078 & w27116;
assign w27118 = ~w26879 & w27117;
assign w27119 = ~w27113 & ~w27118;
assign w27120 = w27109 & w27111;
assign w27121 = (w4430 & w26964) | (w4430 & w42263) | (w26964 & w42263);
assign w27122 = w27120 & ~w27121;
assign w27123 = (~w4056 & w27121) | (~w4056 & w45616) | (w27121 & w45616);
assign w27124 = ~w27119 & w27123;
assign w27125 = ~w27108 & ~w27124;
assign w27126 = ~w27121 & w45617;
assign w27127 = (w4056 & w26879) | (w4056 & w45618) | (w26879 & w45618);
assign w27128 = ~w27113 & w27127;
assign w27129 = ~w27126 & ~w27128;
assign w27130 = (w26718 & w26707) | (w26718 & w42264) | (w26707 & w42264);
assign w27131 = ~w4838 & w27130;
assign w27132 = w4838 & ~w27130;
assign w27133 = ~w27131 & ~w27132;
assign w27134 = ~w26880 & w27133;
assign w27135 = ~w4430 & ~w26710;
assign w27136 = ~w27134 & w27135;
assign w27137 = ~w4430 & w26710;
assign w27138 = w27134 & w27137;
assign w27139 = ~w27136 & ~w27138;
assign w27140 = w27129 & ~w27139;
assign w27141 = w27125 & ~w27140;
assign w27142 = ~w27105 & ~w27141;
assign w27143 = w26718 & w50062;
assign w27144 = (w27143 & w26287) | (w27143 & w42265) | (w26287 & w42265);
assign w27145 = w26706 & w27143;
assign w27146 = w26700 & w27145;
assign w27147 = ~w27144 & ~w27146;
assign w27148 = ~w27146 & w42266;
assign w27149 = ~w26346 & ~w26433;
assign w27150 = w26430 & w27149;
assign w27151 = w26356 & ~w27149;
assign w27152 = (w27151 & ~w42266) | (w27151 & w45619) | (~w42266 & w45619);
assign w27153 = ~w26356 & w27149;
assign w27154 = (~w27153 & ~w42267) | (~w27153 & w45620) | (~w42267 & w45620);
assign w27155 = ~w27152 & w27154;
assign w27156 = w26432 & w26880;
assign w27157 = ~w26880 & w27155;
assign w27158 = ~w27156 & ~w27157;
assign w27159 = w2896 & w27158;
assign w27160 = ~w26422 & ~w26423;
assign w27161 = (~w3646 & w26422) | (~w3646 & w50063) | (w26422 & w50063);
assign w27162 = ~w27143 & w27160;
assign w27163 = ~w3646 & ~w27162;
assign w27164 = (w27163 & w26707) | (w27163 & w42269) | (w26707 & w42269);
assign w27165 = w26350 & ~w26351;
assign w27166 = ~w26350 & w26351;
assign w27167 = ~w27165 & ~w27166;
assign w27168 = (w27167 & w27148) | (w27167 & w50355) | (w27148 & w50355);
assign w27169 = ~w26078 & w27167;
assign w27170 = ~w26879 & w27169;
assign w27171 = ~w27168 & ~w27170;
assign w27172 = (~w26356 & ~w27147) | (~w26356 & w50064) | (~w27147 & w50064);
assign w27173 = w42266 & w50356;
assign w27174 = w26987 & w27173;
assign w27175 = ~w26880 & w27172;
assign w27176 = ~w27174 & ~w27175;
assign w27177 = w27171 & w27176;
assign w27178 = ~w3242 & ~w27177;
assign w27179 = ~w27159 & ~w27178;
assign w27180 = ~w26333 & ~w26431;
assign w27181 = w26357 & w27143;
assign w27182 = (w26357 & w26422) | (w26357 & w45621) | (w26422 & w45621);
assign w27183 = ~w26433 & ~w27182;
assign w27184 = ~w27181 & w27183;
assign w27185 = (~w42271 & w45622) | (~w42271 & w45623) | (w45622 & w45623);
assign w27186 = (w42271 & w45624) | (w42271 & w45625) | (w45624 & w45625);
assign w27187 = ~w27185 & ~w27186;
assign w27188 = ~w26332 & w26880;
assign w27189 = ~w26880 & w27187;
assign w27190 = ~w27188 & ~w27189;
assign w27191 = ~w2558 & w27190;
assign w27192 = (~w27072 & w27007) | (~w27072 & w47754) | (w27007 & w47754);
assign w27193 = ~w26792 & w26880;
assign w27194 = ~w27073 & ~w27192;
assign w27195 = ~w26880 & w27194;
assign w27196 = ~w27193 & ~w27195;
assign w27197 = w2285 & w27196;
assign w27198 = ~w27191 & ~w27197;
assign w27199 = w27179 & w27198;
assign w27200 = w27142 & w27199;
assign w27201 = ~w27168 & w47755;
assign w27202 = w27176 & w27201;
assign w27203 = w2558 & ~w27190;
assign w27204 = ~w2896 & ~w27158;
assign w27205 = ~w27203 & ~w27204;
assign w27206 = ~w27159 & w27202;
assign w27207 = w27205 & ~w27206;
assign w27208 = w27198 & ~w27207;
assign w27209 = (w26782 & w27079) | (w26782 & w50065) | (w27079 & w50065);
assign w27210 = ~w27079 & w50066;
assign w27211 = ~w27209 & ~w27210;
assign w27212 = ~w2006 & w27211;
assign w27213 = ~w2285 & ~w27196;
assign w27214 = ~w27212 & ~w27213;
assign w27215 = ~w27208 & w27214;
assign w27216 = ~w27200 & w27215;
assign w27217 = (w27021 & w27016) | (w27021 & w42272) | (w27016 & w42272);
assign w27218 = ~w26880 & ~w27217;
assign w27219 = ~w27016 & w50067;
assign w27220 = w27218 & ~w27219;
assign w27221 = ~w26799 & ~w26800;
assign w27222 = w26880 & ~w27221;
assign w27223 = ~w1738 & ~w27222;
assign w27224 = ~w27220 & w27223;
assign w27225 = ~w1541 & ~w27043;
assign w27226 = w27040 & w45626;
assign w27227 = ~w1541 & w27043;
assign w27228 = ~w27040 & w27227;
assign w27229 = ~w26078 & w27227;
assign w27230 = ~w26879 & w27229;
assign w27231 = ~w27228 & ~w27230;
assign w27232 = ~w27226 & w27231;
assign w27233 = (~w1320 & ~w27065) | (~w1320 & w50068) | (~w27065 & w50068);
assign w27234 = ~w26732 & w26880;
assign w27235 = w27233 & ~w27234;
assign w27236 = w27070 & ~w27232;
assign w27237 = ~w27235 & ~w27236;
assign w27238 = w27071 & w27224;
assign w27239 = w27237 & ~w27238;
assign w27240 = w27006 & ~w27239;
assign w27241 = w1120 & ~w27001;
assign w27242 = w27000 & w27241;
assign w27243 = w1120 & w27001;
assign w27244 = ~w27000 & w27243;
assign w27245 = ~w27242 & ~w27244;
assign w27246 = ~w27240 & w27245;
assign w27247 = w27087 & ~w27216;
assign w27248 = w27246 & ~w27247;
assign w27249 = w26990 & w50069;
assign w27250 = w26978 & ~w26995;
assign w27251 = ~w27249 & w26978;
assign w27252 = ~w27247 & w45627;
assign w27253 = ~w27250 & ~w27252;
assign w27254 = ~w26974 & ~w27249;
assign w27255 = w27245 & w27254;
assign w27256 = ~w27240 & w27255;
assign w27257 = w26995 & ~w27256;
assign w27258 = (w26978 & w27256) | (w26978 & w27250) | (w27256 & w27250);
assign w27259 = w26995 & w27087;
assign w27260 = ~w27257 & w42273;
assign w27261 = ~a[24] & w25851;
assign w27262 = a[24] & ~w25851;
assign w27263 = ~w27261 & ~w27262;
assign w27264 = a[24] & ~w26478;
assign w27265 = ~w26479 & ~w27264;
assign w27266 = w26073 & w42274;
assign w27267 = ~w26077 & w42275;
assign w27268 = ~w27266 & w52261;
assign w27269 = (~w27263 & w26964) | (~w27263 & w42276) | (w26964 & w42276);
assign w27270 = w27268 & ~w27269;
assign w27271 = ~a[20] & ~a[21];
assign w27272 = ~a[22] & w27271;
assign w27273 = w25851 & w27272;
assign w27274 = ~w25851 & ~w27272;
assign w27275 = ~a[23] & ~w27274;
assign w27276 = ~w27273 & ~w27275;
assign w27277 = (~w27276 & w26891) | (~w27276 & w42277) | (w26891 & w42277);
assign w27278 = a[23] & w27274;
assign w27279 = ~w26478 & ~w27278;
assign w27280 = w26078 & w27279;
assign w27281 = ~w26077 & w50070;
assign w27282 = (~w27280 & w26827) | (~w27280 & w47758) | (w26827 & w47758);
assign w27283 = ~w27277 & w27282;
assign w27284 = ~w24874 & w27266;
assign w27285 = ~w26077 & w50071;
assign w27286 = ~w26827 & w27285;
assign w27287 = ~w27284 & ~w27286;
assign w27288 = ~w24874 & ~w27263;
assign w27289 = (w27288 & w26964) | (w27288 & w42278) | (w26964 & w42278);
assign w27290 = w27287 & ~w27289;
assign w27291 = w24874 & w27270;
assign w27292 = ~w27283 & w27290;
assign w27293 = ~w27291 & ~w27292;
assign w27294 = a[25] & ~w26484;
assign w27295 = ~w26485 & ~w27294;
assign w27296 = w25851 & ~w27295;
assign w27297 = ~w25851 & w27295;
assign w27298 = ~w27296 & ~w27297;
assign w27299 = a[25] & w27261;
assign w27300 = ~w26072 & w42279;
assign w27301 = w27299 & ~w27300;
assign w27302 = (w27301 & w26892) | (w27301 & w50072) | (w26892 & w50072);
assign w27303 = w26889 & w27301;
assign w27304 = ~w26708 & w27303;
assign w27305 = ~w27302 & ~w27304;
assign w27306 = (~w27298 & w26893) | (~w27298 & w45628) | (w26893 & w45628);
assign w27307 = ~w26964 & w27306;
assign w27308 = w27305 & ~w27307;
assign w27309 = ~a[25] & ~w27261;
assign w27310 = (w27309 & w26964) | (w27309 & w42280) | (w26964 & w42280);
assign w27311 = w27308 & ~w27310;
assign w27312 = ~w22767 & ~w26476;
assign w27313 = w23843 & w26490;
assign w27314 = ~w26491 & ~w27313;
assign w27315 = w27312 & ~w27314;
assign w27316 = ~w26077 & w50073;
assign w27317 = w26073 & w42281;
assign w27318 = w27312 & ~w27317;
assign w27319 = ~w26827 & w27316;
assign w27320 = w27318 & ~w27319;
assign w27321 = w26492 & w26502;
assign w27322 = ~w22767 & w27321;
assign w27323 = w26073 & w42282;
assign w27324 = ~w26077 & w50074;
assign w27325 = ~w26827 & w27324;
assign w27326 = ~w27323 & ~w27325;
assign w27327 = ~w27320 & w27326;
assign w27328 = w27308 & w42283;
assign w27329 = w27327 & ~w27328;
assign w27330 = ~w27293 & w27329;
assign w27331 = ~w26476 & ~w27314;
assign w27332 = w26878 & ~w27331;
assign w27333 = ~w26827 & w27332;
assign w27334 = w26078 & w27321;
assign w27335 = w26878 & w27321;
assign w27336 = (~w27334 & w26827) | (~w27334 & w47759) | (w26827 & w47759);
assign w27337 = ~w26476 & ~w27317;
assign w27338 = ~w27333 & w27337;
assign w27339 = w27336 & ~w27338;
assign w27340 = ~w27338 & w47760;
assign w27341 = w23843 & ~w27323;
assign w27342 = ~w27325 & w27341;
assign w27343 = ~w27320 & w27342;
assign w27344 = ~w27311 & w27343;
assign w27345 = ~w27340 & ~w27344;
assign w27346 = w20906 & w26520;
assign w27347 = ~w26078 & w27346;
assign w27348 = ~w26879 & w27347;
assign w27349 = w26512 & ~w26521;
assign w27350 = ~w26492 & w26502;
assign w27351 = w22767 & ~w27350;
assign w27352 = ~w26505 & ~w27351;
assign w27353 = w27349 & ~w27352;
assign w27354 = ~w27349 & w27352;
assign w27355 = ~w27353 & ~w27354;
assign w27356 = w20906 & w27355;
assign w27357 = w26078 & w27356;
assign w27358 = w26878 & w27356;
assign w27359 = (~w27357 & w26827) | (~w27357 & w47761) | (w26827 & w47761);
assign w27360 = ~w27348 & w27359;
assign w27361 = ~w20000 & ~w26561;
assign w27362 = ~w26078 & w27361;
assign w27363 = ~w26879 & w27362;
assign w27364 = w26531 & ~w26562;
assign w27365 = (~w27364 & w26517) | (~w27364 & w50075) | (w26517 & w50075);
assign w27366 = ~w26517 & w45629;
assign w27367 = ~w27365 & ~w27366;
assign w27368 = ~w20000 & w27367;
assign w27369 = w26078 & w27368;
assign w27370 = w26878 & w27368;
assign w27371 = (~w27369 & w26827) | (~w27369 & w47762) | (w26827 & w47762);
assign w27372 = ~w27363 & w27371;
assign w27373 = w27360 & w27372;
assign w27374 = ~w26504 & ~w27351;
assign w27375 = ~w26077 & w42284;
assign w27376 = (~w42235 & w47763) | (~w42235 & w47764) | (w47763 & w47764);
assign w27377 = w26073 & w42285;
assign w27378 = ~w26469 & w27375;
assign w27379 = ~w26827 & w27378;
assign w27380 = w26469 & ~w27377;
assign w27381 = ~w27376 & w27380;
assign w27382 = ~w26469 & w27377;
assign w27383 = ~w27379 & ~w27382;
assign w27384 = ~w27381 & w27383;
assign w27385 = (~w21801 & ~w27383) | (~w21801 & w47765) | (~w27383 & w47765);
assign w27386 = w27373 & ~w27385;
assign w27387 = w27345 & w27386;
assign w27388 = ~w27330 & w27387;
assign w27389 = ~w26600 & ~w26619;
assign w27390 = (w26517 & w50076) | (w26517 & w50077) | (w50076 & w50077);
assign w27391 = w18183 & w52262;
assign w27392 = ~w27390 & ~w27391;
assign w27393 = ~w26077 & w50078;
assign w27394 = ~w26827 & w27393;
assign w27395 = w26878 & w42288;
assign w27396 = ~w26827 & w27395;
assign w27397 = (~w26615 & ~w42287) | (~w26615 & w50079) | (~w42287 & w50079);
assign w27398 = ~w27394 & w27397;
assign w27399 = w42287 & w50080;
assign w27400 = ~w27396 & ~w27399;
assign w27401 = ~w27398 & w27400;
assign w27402 = ~w17380 & ~w27401;
assign w27403 = w26599 & ~w27366;
assign w27404 = w26557 & ~w27403;
assign w27405 = w26078 & ~w27404;
assign w27406 = w26878 & ~w27404;
assign w27407 = (~w27405 & w26827) | (~w27405 & w47766) | (w26827 & w47766);
assign w27408 = w19040 & ~w26078;
assign w27409 = ~w26879 & w27408;
assign w27410 = w27407 & ~w27409;
assign w27411 = w26546 & ~w26619;
assign w27412 = w18183 & ~w27411;
assign w27413 = ~w27410 & w27412;
assign w27414 = w18183 & w27411;
assign w27415 = w27410 & w27414;
assign w27416 = ~w27413 & ~w27415;
assign w27417 = ~w27402 & w27416;
assign w27418 = w21801 & ~w26469;
assign w27419 = ~w27377 & w27418;
assign w27420 = ~w27376 & w27419;
assign w27421 = w21801 & w26469;
assign w27422 = ~w26077 & w50081;
assign w27423 = ~w26827 & w27422;
assign w27424 = w27377 & w27421;
assign w27425 = ~w27423 & ~w27424;
assign w27426 = ~w27420 & w27425;
assign w27427 = ~w20906 & ~w26520;
assign w27428 = ~w26078 & w27427;
assign w27429 = ~w26879 & w27428;
assign w27430 = ~w20906 & ~w27355;
assign w27431 = w26078 & w27430;
assign w27432 = w26878 & w27430;
assign w27433 = (~w27431 & w26827) | (~w27431 & w47767) | (w26827 & w47767);
assign w27434 = ~w27429 & w27433;
assign w27435 = w27426 & w27434;
assign w27436 = w25153 & ~w25851;
assign w27437 = w25851 & w26552;
assign w27438 = ~w27436 & ~w27437;
assign w27439 = (w26557 & ~w42289) | (w26557 & w45630) | (~w42289 & w45630);
assign w27440 = ~w26077 & w50082;
assign w27441 = (w27439 & w26827) | (w27439 & w47768) | (w26827 & w47768);
assign w27442 = ~w26078 & ~w27438;
assign w27443 = ~w26879 & w27442;
assign w27444 = w27441 & ~w27443;
assign w27445 = w26531 & ~w27366;
assign w27446 = ~w26557 & ~w27445;
assign w27447 = ~w26598 & ~w27445;
assign w27448 = (~w27447 & w26891) | (~w27447 & w42290) | (w26891 & w42290);
assign w27449 = w19040 & w27448;
assign w27450 = ~w27444 & w27449;
assign w27451 = w20000 & w26561;
assign w27452 = w26880 & w27451;
assign w27453 = w20000 & ~w27367;
assign w27454 = ~w26880 & w27453;
assign w27455 = ~w27452 & ~w27454;
assign w27456 = ~w27450 & w27455;
assign w27457 = w27373 & ~w27435;
assign w27458 = w27456 & ~w27457;
assign w27459 = w27417 & w27458;
assign w27460 = ~w27388 & w27459;
assign w27461 = (~w19040 & w27444) | (~w19040 & w45631) | (w27444 & w45631);
assign w27462 = ~w18183 & w27411;
assign w27463 = ~w27410 & w27462;
assign w27464 = ~w18183 & ~w27411;
assign w27465 = w27410 & w27464;
assign w27466 = ~w27463 & ~w27465;
assign w27467 = ~w27461 & w27466;
assign w27468 = w27417 & ~w27467;
assign w27469 = ~w26078 & ~w26652;
assign w27470 = ~w26879 & w27469;
assign w27471 = ~w26653 & ~w26692;
assign w27472 = ~w26689 & w52263;
assign w27473 = w27471 & ~w27472;
assign w27474 = ~w27471 & w27472;
assign w27475 = ~w17380 & w27473;
assign w27476 = (~w27475 & ~w42292) | (~w27475 & w50083) | (~w42292 & w50083);
assign w27477 = ~w26077 & w50179;
assign w27478 = ~w26827 & w27477;
assign w27479 = w27476 & ~w27478;
assign w27480 = w27473 & w26895;
assign w27481 = w27479 & ~w27480;
assign w27482 = ~w27470 & w27481;
assign w27483 = ~w16559 & ~w27482;
assign w27484 = w17380 & w27401;
assign w27485 = ~w27483 & ~w27484;
assign w27486 = ~w27468 & w27485;
assign w27487 = ~w27460 & w27486;
assign w27488 = w26282 & ~w26704;
assign w27489 = ~w26668 & w42293;
assign w27490 = (w27488 & w26668) | (w27488 & w42294) | (w26668 & w42294);
assign w27491 = ~w27489 & ~w27490;
assign w27492 = w26078 & w27491;
assign w27493 = w26878 & w27491;
assign w27494 = (~w27492 & w26827) | (~w27492 & w47769) | (w26827 & w47769);
assign w27495 = ~w26078 & ~w26703;
assign w27496 = ~w26879 & w27495;
assign w27497 = w27494 & ~w27496;
assign w27498 = w12666 & w27497;
assign w27499 = w26173 & ~w26270;
assign w27500 = (w26282 & w26668) | (w26282 & w42295) | (w26668 & w42295);
assign w27501 = ~w27499 & w27500;
assign w27502 = w26078 & ~w27501;
assign w27503 = w26878 & ~w27501;
assign w27504 = (~w27502 & w26827) | (~w27502 & w47770) | (w26827 & w47770);
assign w27505 = ~w26078 & w26269;
assign w27506 = ~w26879 & w27505;
assign w27507 = w27504 & ~w27506;
assign w27508 = w27499 & ~w27500;
assign w27509 = ~w26269 & w27508;
assign w27510 = ~w26894 & w27508;
assign w27511 = (~w27509 & w26891) | (~w27509 & w42296) | (w26891 & w42296);
assign w27512 = (w45632 & w50357) | (w45632 & w42296) | (w50357 & w42296);
assign w27513 = ~w27507 & w27512;
assign w27514 = ~w27498 & ~w27513;
assign w27515 = ~w27507 & w27511;
assign w27516 = (~w11870 & w27507) | (~w11870 & w45633) | (w27507 & w45633);
assign w27517 = w14039 & ~w26580;
assign w27518 = ~w26078 & ~w27517;
assign w27519 = w26565 & w26697;
assign w27520 = ~w26517 & w27519;
assign w27521 = ~w26666 & w26697;
assign w27522 = ~w26573 & ~w27521;
assign w27523 = ~w27520 & w27522;
assign w27524 = w15681 & w26572;
assign w27525 = ~w27523 & ~w27524;
assign w27526 = ~w26581 & w26680;
assign w27527 = w14039 & w27526;
assign w27528 = (w27527 & w27523) | (w27527 & w42297) | (w27523 & w42297);
assign w27529 = w14039 & ~w27526;
assign w27530 = ~w27523 & w42298;
assign w27531 = ~w27528 & ~w27530;
assign w27532 = w26078 & w27531;
assign w27533 = w26878 & w27531;
assign w27534 = ~w26827 & w27533;
assign w27535 = ~w27532 & ~w27534;
assign w27536 = ~w26879 & w27518;
assign w27537 = w27535 & ~w27536;
assign w27538 = ~w13384 & w26591;
assign w27539 = w26582 & ~w27521;
assign w27540 = ~w27520 & w27539;
assign w27541 = ~w26675 & w26680;
assign w27542 = (~w14039 & w27540) | (~w14039 & w42299) | (w27540 & w42299);
assign w27543 = ~w27540 & w42300;
assign w27544 = w26878 & ~w27543;
assign w27545 = w27538 & w27542;
assign w27546 = w27544 & ~w27545;
assign w27547 = ~w27542 & ~w27543;
assign w27548 = (w27538 & ~w26078) | (w27538 & w42301) | (~w26078 & w42301);
assign w27549 = ~w26827 & w27546;
assign w27550 = w27548 & ~w27549;
assign w27551 = ~w13384 & ~w26591;
assign w27552 = w26078 & w42302;
assign w27553 = ~w27542 & w27551;
assign w27554 = w27544 & w27553;
assign w27555 = ~w26827 & w27554;
assign w27556 = ~w27552 & ~w27555;
assign w27557 = ~w27550 & w27556;
assign w27558 = ~w27537 & w27557;
assign w27559 = w13384 & ~w26591;
assign w27560 = w27543 & w27559;
assign w27561 = w26878 & ~w27542;
assign w27562 = ~w27560 & w27561;
assign w27563 = ~w26827 & w27562;
assign w27564 = (w27559 & ~w26078) | (w27559 & w42303) | (~w26078 & w42303);
assign w27565 = ~w27563 & w27564;
assign w27566 = w13384 & w26591;
assign w27567 = w26078 & w42304;
assign w27568 = ~w27542 & w27566;
assign w27569 = w27544 & w27568;
assign w27570 = ~w26827 & w27569;
assign w27571 = ~w27567 & ~w27570;
assign w27572 = ~w27565 & w27571;
assign w27573 = ~w27558 & w27572;
assign w27574 = ~w27520 & w50358;
assign w27575 = (w15681 & w27520) | (w15681 & w50359) | (w27520 & w50359);
assign w27576 = ~w27574 & ~w27575;
assign w27577 = w26078 & ~w27576;
assign w27578 = w26878 & ~w27576;
assign w27579 = ~w26827 & w27578;
assign w27580 = ~w27577 & ~w27579;
assign w27581 = w14766 & ~w26572;
assign w27582 = ~w27580 & w27581;
assign w27583 = w14766 & w26572;
assign w27584 = w27580 & w27583;
assign w27585 = ~w27582 & ~w27584;
assign w27586 = ~w14039 & w26580;
assign w27587 = ~w26078 & ~w27586;
assign w27588 = ~w14039 & ~w27526;
assign w27589 = (w27588 & w27523) | (w27588 & w42305) | (w27523 & w42305);
assign w27590 = ~w14039 & w27526;
assign w27591 = ~w27523 & w42306;
assign w27592 = ~w27589 & ~w27591;
assign w27593 = w26078 & w27592;
assign w27594 = w26878 & w27592;
assign w27595 = ~w26827 & w27594;
assign w27596 = ~w27593 & ~w27595;
assign w27597 = ~w26879 & w27587;
assign w27598 = w27596 & ~w27597;
assign w27599 = w27572 & ~w27598;
assign w27600 = w27585 & w27599;
assign w27601 = ~w27573 & ~w27600;
assign w27602 = ~w12666 & ~w27497;
assign w27603 = ~w27514 & ~w27516;
assign w27604 = ~w27516 & ~w27602;
assign w27605 = (~w27603 & w27601) | (~w27603 & w42307) | (w27601 & w42307);
assign w27606 = ~w26664 & ~w26690;
assign w27607 = ~w26692 & ~w27473;
assign w27608 = w26078 & ~w27607;
assign w27609 = w26878 & ~w27607;
assign w27610 = (~w27608 & w26827) | (~w27608 & w47771) | (w26827 & w47771);
assign w27611 = w16559 & ~w26078;
assign w27612 = ~w26879 & w27611;
assign w27613 = w27610 & ~w27612;
assign w27614 = w27606 & ~w27613;
assign w27615 = ~w27606 & w27613;
assign w27616 = ~w27614 & ~w27615;
assign w27617 = w15681 & w27616;
assign w27618 = w26666 & w27620;
assign w27619 = ~w26566 & w27618;
assign w27620 = w26283 & w26593;
assign w27621 = ~w26697 & w27620;
assign w27622 = w26283 & ~w26944;
assign w27623 = ~w27621 & ~w27622;
assign w27624 = w26173 & w27623;
assign w27625 = ~w27619 & w27624;
assign w27626 = w11870 & ~w27625;
assign w27627 = ~w11870 & w27625;
assign w27628 = ~w27626 & ~w27627;
assign w27629 = w26878 & ~w27628;
assign w27630 = ~w26827 & w27629;
assign w27631 = (w26127 & w27630) | (w26127 & w42308) | (w27630 & w42308);
assign w27632 = ~w27630 & w42309;
assign w27633 = ~w27631 & ~w27632;
assign w27634 = w11138 & ~w27633;
assign w27635 = (w16559 & w26879) | (w16559 & w50084) | (w26879 & w50084);
assign w27636 = w27481 & w27635;
assign w27637 = ~w27634 & ~w27636;
assign w27638 = ~w27617 & w27637;
assign w27639 = ~w27605 & w27638;
assign w27640 = ~w27487 & w27639;
assign w27641 = ~w15681 & ~w27616;
assign w27642 = ~w14766 & w26572;
assign w27643 = (w27642 & w27579) | (w27642 & w50360) | (w27579 & w50360);
assign w27644 = ~w14766 & ~w26572;
assign w27645 = ~w27579 & w50361;
assign w27646 = ~w27643 & ~w27645;
assign w27647 = w27557 & w50362;
assign w27648 = w27514 & w27647;
assign w27649 = ~w27641 & w27648;
assign w27650 = (~w27634 & ~w27648) | (~w27634 & w42310) | (~w27648 & w42310);
assign w27651 = ~w27605 & w27650;
assign w27652 = w26159 & w26173;
assign w27653 = w27623 & w27652;
assign w27654 = ~w27619 & w27653;
assign w27655 = ~w26138 & ~w27654;
assign w27656 = (w26115 & w27654) | (w26115 & w45634) | (w27654 & w45634);
assign w27657 = ~w26155 & ~w27656;
assign w27658 = w9195 & w26086;
assign w27659 = w27657 & w27658;
assign w27660 = ~w26078 & w26086;
assign w27661 = ~w26879 & w27660;
assign w27662 = ~w27659 & ~w27661;
assign w27663 = w9195 & ~w26078;
assign w27664 = ~w26879 & w27663;
assign w27665 = ~w26087 & ~w26156;
assign w27666 = ~w27657 & ~w27665;
assign w27667 = ~w27664 & w27666;
assign w27668 = w26895 & w45635;
assign w27669 = ~w27667 & ~w27668;
assign w27670 = w27662 & w27669;
assign w27671 = (w8666 & ~w27669) | (w8666 & w45636) | (~w27669 & w45636);
assign w27672 = w10419 & ~w26148;
assign w27673 = (~w26148 & ~w42311) | (~w26148 & w45637) | (~w42311 & w45637);
assign w27674 = ~w26077 & w50085;
assign w27675 = ~w26827 & w27674;
assign w27676 = w27673 & ~w27675;
assign w27677 = ~w26138 & w26143;
assign w27678 = ~w27654 & w27677;
assign w27679 = ~w10419 & w26148;
assign w27680 = (~w27679 & w27654) | (~w27679 & w42312) | (w27654 & w42312);
assign w27681 = w26078 & ~w27680;
assign w27682 = w26878 & ~w27680;
assign w27683 = ~w26827 & w27682;
assign w27684 = ~w27681 & ~w27683;
assign w27685 = ~w27654 & w45638;
assign w27686 = w27678 & w27679;
assign w27687 = (~w27686 & ~w42313) | (~w27686 & w45639) | (~w42313 & w45639);
assign w27688 = ~w27676 & w27684;
assign w27689 = (w9781 & w27688) | (w9781 & w45640) | (w27688 & w45640);
assign w27690 = ~w26234 & w26243;
assign w27691 = w25038 & ~w26243;
assign w27692 = ~w27690 & ~w27691;
assign w27693 = w26248 & w26292;
assign w27694 = w26949 & w45641;
assign w27695 = (w27693 & ~w26949) | (w27693 & w45642) | (~w26949 & w45642);
assign w27696 = ~w27694 & ~w27695;
assign w27697 = w7924 & ~w27692;
assign w27698 = w26880 & w27697;
assign w27699 = w7924 & ~w27696;
assign w27700 = ~w26880 & w27699;
assign w27701 = ~w27698 & ~w27700;
assign w27702 = ~w26105 & ~w26155;
assign w27703 = (w27654 & w50086) | (w27654 & w50087) | (w50086 & w50087);
assign w27704 = w27702 & w52264;
assign w27705 = ~w27703 & ~w27704;
assign w27706 = ~w26880 & w27705;
assign w27707 = ~w26078 & w26154;
assign w27708 = ~w26879 & w27707;
assign w27709 = (~w9195 & w26879) | (~w9195 & w45644) | (w26879 & w45644);
assign w27710 = ~w27706 & w27709;
assign w27711 = w27701 & ~w27710;
assign w27712 = ~w27689 & w27711;
assign w27713 = ~w27671 & w27712;
assign w27714 = ~w26078 & ~w26229;
assign w27715 = ~w26879 & w27714;
assign w27716 = ~w26230 & ~w26233;
assign w27717 = (w42314 & ~w26176) | (w42314 & w45645) | (~w26176 & w45645);
assign w27718 = (w26949 & w50088) | (w26949 & w50089) | (w50088 & w50089);
assign w27719 = ~w27716 & w52265;
assign w27720 = ~w27718 & ~w27719;
assign w27721 = ~w26880 & w27720;
assign w27722 = ~w27715 & ~w27721;
assign w27723 = w7315 & ~w27722;
assign w27724 = w24967 & ~w26132;
assign w27725 = ~w24967 & w26132;
assign w27726 = ~w27724 & ~w27725;
assign w27727 = w11138 & ~w27655;
assign w27728 = ~w26964 & w42315;
assign w27729 = ~w26128 & ~w26143;
assign w27730 = (w27729 & ~w27625) | (w27729 & w42316) | (~w27625 & w42316);
assign w27731 = w26878 & w27730;
assign w27732 = ~w26827 & w27731;
assign w27733 = ~w26128 & ~w26137;
assign w27734 = (w27733 & ~w27625) | (w27733 & w42317) | (~w27625 & w42317);
assign w27735 = (w27726 & w27654) | (w27726 & w45647) | (w27654 & w45647);
assign w27736 = ~w27734 & ~w27735;
assign w27737 = w26078 & w27730;
assign w27738 = w27736 & ~w27737;
assign w27739 = ~w27732 & w27738;
assign w27740 = ~w27728 & w27739;
assign w27741 = w27740 & w42318;
assign w27742 = ~w11138 & w27633;
assign w27743 = ~w27741 & ~w27742;
assign w27744 = ~w27723 & w27743;
assign w27745 = w27713 & w27744;
assign w27746 = ~w27651 & w27745;
assign w27747 = ~w27640 & w27746;
assign w27748 = ~w26194 & w26293;
assign w27749 = ~w26194 & ~w26232;
assign w27750 = (w26949 & w50090) | (w26949 & w50091) | (w50090 & w50091);
assign w27751 = w26253 & w27750;
assign w27752 = ~w26880 & w27751;
assign w27753 = w26204 & ~w26232;
assign w27754 = ~w26203 & w27748;
assign w27755 = (w26949 & w50092) | (w26949 & w50093) | (w50092 & w50093);
assign w27756 = w26203 & w27750;
assign w27757 = w26252 & ~w27755;
assign w27758 = ~w27756 & ~w27757;
assign w27759 = ~w6769 & ~w27755;
assign w27760 = w26987 & w27759;
assign w27761 = w27758 & ~w27760;
assign w27762 = w26252 & w26880;
assign w27763 = w27761 & ~w27762;
assign w27764 = ~w26194 & ~w26231;
assign w27765 = w26293 & ~w27764;
assign w27766 = (w27765 & ~w26949) | (w27765 & w42321) | (~w26949 & w42321);
assign w27767 = ~w26230 & w27764;
assign w27768 = w26949 & w42322;
assign w27769 = ~w27766 & ~w27768;
assign w27770 = w26230 & ~w27764;
assign w27771 = ~w26293 & w27764;
assign w27772 = ~w26230 & w27771;
assign w27773 = ~w27770 & ~w27772;
assign w27774 = w27769 & w27773;
assign w27775 = w6769 & ~w26193;
assign w27776 = w26880 & w27775;
assign w27777 = w6769 & ~w27774;
assign w27778 = ~w26880 & w27777;
assign w27779 = ~w27776 & ~w27778;
assign w27780 = w27763 & w42323;
assign w27781 = ~w6264 & ~w27779;
assign w27782 = ~w6264 & ~w27752;
assign w27783 = w27763 & w27782;
assign w27784 = ~w27781 & ~w27783;
assign w27785 = ~w27780 & w27784;
assign w27786 = w26078 & ~w26306;
assign w27787 = ~w26077 & w49144;
assign w27788 = ~w26253 & ~w27753;
assign w27789 = ~w27754 & w27788;
assign w27790 = w27717 & w27788;
assign w27791 = (~w27789 & ~w26949) | (~w27789 & w42324) | (~w26949 & w42324);
assign w27792 = (~w26949 & w49145) | (~w26949 & w49146) | (w49145 & w49146);
assign w27793 = ~w26264 & w26716;
assign w27794 = (w26949 & w50094) | (w26949 & w50095) | (w50094 & w50095);
assign w27795 = (~w47772 & w49147) | (~w47772 & w49148) | (w49147 & w49148);
assign w27796 = ~w5330 & ~w26078;
assign w27797 = ~w26879 & w27796;
assign w27798 = ~w26314 & ~w26711;
assign w27799 = w4838 & w27798;
assign w27800 = (w27799 & w26879) | (w27799 & w49149) | (w26879 & w49149);
assign w27801 = ~w27795 & w27800;
assign w27802 = w4838 & ~w27798;
assign w27803 = ~w26879 & w49150;
assign w27804 = ~w27794 & w27802;
assign w27805 = w27804 & w52266;
assign w27806 = ~w27803 & ~w27805;
assign w27807 = ~w27801 & w27806;
assign w27808 = w26078 & ~w26264;
assign w27809 = ~w26077 & w45648;
assign w27810 = (~w42235 & w47773) | (~w42235 & w47774) | (w47773 & w47774);
assign w27811 = (~w27792 & w27810) | (~w27792 & w45649) | (w27810 & w45649);
assign w27812 = ~w5745 & ~w26078;
assign w27813 = ~w26306 & w26716;
assign w27814 = ~w5330 & ~w27813;
assign w27815 = (w27814 & w26879) | (w27814 & w49151) | (w26879 & w49151);
assign w27816 = ~w27811 & w27815;
assign w27817 = ~w5330 & w27813;
assign w27818 = ~w27792 & w27817;
assign w27819 = (w27818 & w27810) | (w27818 & w49152) | (w27810 & w49152);
assign w27820 = ~w26879 & w49153;
assign w27821 = ~w27819 & ~w27820;
assign w27822 = ~w27816 & w27821;
assign w27823 = w27807 & w27822;
assign w27824 = (w26263 & ~w42325) | (w26263 & w45650) | (~w42325 & w45650);
assign w27825 = ~w27810 & w27824;
assign w27826 = w26295 & ~w27791;
assign w27827 = (w26949 & w45651) | (w26949 & w45652) | (w45651 & w45652);
assign w27828 = (~w27826 & ~w42326) | (~w27826 & w45653) | (~w42326 & w45653);
assign w27829 = w5745 & w27828;
assign w27830 = ~w27811 & ~w27825;
assign w27831 = w27829 & ~w27830;
assign w27832 = w27807 & w49154;
assign w27833 = w27785 & w27832;
assign w27834 = ~w5745 & ~w27828;
assign w27835 = (~w5745 & w27810) | (~w5745 & w45654) | (w27810 & w45654);
assign w27836 = ~w27811 & w27835;
assign w27837 = ~w27834 & ~w27836;
assign w27838 = w5330 & w27813;
assign w27839 = (w27838 & w26879) | (w27838 & w45655) | (w26879 & w45655);
assign w27840 = ~w27811 & w27839;
assign w27841 = w5330 & ~w27813;
assign w27842 = ~w27792 & w27841;
assign w27843 = (w27842 & w27810) | (w27842 & w49155) | (w27810 & w49155);
assign w27844 = ~w26879 & w45656;
assign w27845 = ~w27843 & ~w27844;
assign w27846 = ~w27840 & w27845;
assign w27847 = w27837 & w27846;
assign w27848 = w27823 & ~w27847;
assign w27849 = (~w27848 & ~w27785) | (~w27848 & w42327) | (~w27785 & w42327);
assign w27850 = (~w7315 & w26879) | (~w7315 & w45657) | (w26879 & w45657);
assign w27851 = ~w27721 & w27850;
assign w27852 = ~w7924 & w27692;
assign w27853 = w26880 & w27852;
assign w27854 = ~w7924 & w27696;
assign w27855 = ~w26880 & w27854;
assign w27856 = ~w27853 & ~w27855;
assign w27857 = ~w27851 & w27856;
assign w27858 = ~w27706 & ~w27708;
assign w27859 = w9195 & ~w27858;
assign w27860 = ~w27661 & w45658;
assign w27861 = w27669 & w27860;
assign w27862 = ~w27859 & ~w27861;
assign w27863 = w27669 & w45659;
assign w27864 = ~w8666 & w27701;
assign w27865 = ~w27861 & w45660;
assign w27866 = w27857 & ~w27864;
assign w27867 = ~w27863 & w27866;
assign w27868 = ~w27865 & ~w27867;
assign w27869 = ~w27688 & w45661;
assign w27870 = (~w10419 & ~w27740) | (~w10419 & w42328) | (~w27740 & w42328);
assign w27871 = ~w27869 & ~w27870;
assign w27872 = w27713 & ~w27871;
assign w27873 = ~w27868 & ~w27872;
assign w27874 = ~w27723 & ~w27873;
assign w27875 = ~w27849 & ~w27874;
assign w27876 = ~w27747 & w27875;
assign w27877 = w26193 & w26880;
assign w27878 = ~w26880 & w27774;
assign w27879 = ~w27877 & ~w27878;
assign w27880 = ~w6769 & ~w27879;
assign w27881 = (~w42327 & w49156) | (~w42327 & w49157) | (w49156 & w49157);
assign w27882 = w27761 & w42329;
assign w27883 = w6264 & ~w27882;
assign w27884 = ~w27831 & w27883;
assign w27885 = (w27823 & w27884) | (w27823 & w27848) | (w27884 & w27848);
assign w27886 = w4430 & w26710;
assign w27887 = ~w27134 & w27886;
assign w27888 = w4430 & ~w26710;
assign w27889 = w27134 & w27888;
assign w27890 = ~w27887 & ~w27889;
assign w27891 = w27129 & w27890;
assign w27892 = w27125 & ~w27891;
assign w27893 = ~w27105 & ~w27892;
assign w27894 = (~w27202 & w27892) | (~w27202 & w47775) | (w27892 & w47775);
assign w27895 = ~w27795 & ~w27797;
assign w27896 = ~w4838 & w27798;
assign w27897 = ~w27895 & w27896;
assign w27898 = ~w4838 & ~w27798;
assign w27899 = w27895 & w27898;
assign w27900 = ~w27897 & ~w27899;
assign w27901 = w27198 & w27900;
assign w27902 = w27179 & w27901;
assign w27903 = ~w27894 & w27902;
assign w27904 = ~w27885 & w27903;
assign w27905 = ~w27881 & w27904;
assign w27906 = (w27905 & w27747) | (w27905 & w47776) | (w27747 & w47776);
assign w27907 = ~w27876 & w42330;
assign w27908 = ~w27253 & ~w27907;
assign w27909 = w25931 & ~w26047;
assign w27910 = ~w26892 & w27909;
assign w27911 = (w42331 & w50096) | (w42331 & w50097) | (w50096 & w50097);
assign w27912 = w25868 & ~w27911;
assign w27913 = ~w25814 & ~w25868;
assign w27914 = w27911 & w27913;
assign w27915 = ~w27912 & ~w27914;
assign w27916 = ~w42 & w27915;
assign w27917 = w25887 & w25936;
assign w27918 = ~w3 & w26880;
assign w27919 = (~w42331 & w45664) | (~w42331 & w45665) | (w45664 & w45665);
assign w27920 = ~w26880 & w27919;
assign w27921 = ~w27918 & ~w27920;
assign w27922 = w27917 & ~w27921;
assign w27923 = ~w27917 & w27921;
assign w27924 = ~w27922 & ~w27923;
assign w27925 = ~w25947 & w26078;
assign w27926 = ~w26077 & w45666;
assign w27927 = ~w26827 & w27926;
assign w27928 = ~w27925 & ~w27927;
assign w27929 = ~w26034 & ~w26045;
assign w27930 = ~w25925 & ~w27929;
assign w27931 = (w27930 & w26885) | (w27930 & w45667) | (w26885 & w45667);
assign w27932 = ~w27928 & ~w27931;
assign w27933 = w80 & w26880;
assign w27934 = ~w27932 & ~w27933;
assign w27935 = w25898 & w25930;
assign w27936 = (~w27935 & w27932) | (~w27935 & w50098) | (w27932 & w50098);
assign w27937 = w3 & ~w27936;
assign w27938 = w27934 & w27935;
assign w27939 = w27937 & ~w27938;
assign w27940 = w27916 & w27924;
assign w27941 = w27939 & ~w27940;
assign w27942 = w25871 & ~w27911;
assign w27943 = ~w25868 & ~w27942;
assign w27944 = w42 & ~w27912;
assign w27945 = ~w27943 & w27944;
assign w27946 = w27924 & ~w27945;
assign w27947 = w27924 & w50099;
assign w27948 = ~w27916 & ~w27947;
assign w27949 = ~w27941 & ~w27948;
assign w27950 = ~w25982 & ~w26022;
assign w27951 = w26003 & ~w26022;
assign w27952 = ~w27950 & w52267;
assign w27953 = (~w42334 & w27981) | (~w42334 & w45668) | (w27981 & w45668);
assign w27954 = ~w26077 & w49158;
assign w27955 = (~w27953 & w26827) | (~w27953 & w47777) | (w26827 & w47777);
assign w27956 = ~w26038 & w26078;
assign w27957 = ~w26077 & w45669;
assign w27958 = (~w42235 & w47778) | (~w42235 & w47779) | (w47778 & w47779);
assign w27959 = ~w27956 & ~w27958;
assign w27960 = w252 & ~w26078;
assign w27961 = ~w26879 & w27960;
assign w27962 = w27959 & ~w27961;
assign w27963 = ~w27952 & ~w27955;
assign w27964 = w26030 & w26043;
assign w27965 = w27962 & w50100;
assign w27966 = (w27964 & ~w27962) | (w27964 & w50101) | (~w27962 & w50101);
assign w27967 = ~w27965 & ~w27966;
assign w27968 = ~w57 & ~w27967;
assign w27969 = ~w26021 & w26038;
assign w27970 = w26078 & w27969;
assign w27971 = ~w26077 & w45670;
assign w27972 = (~w42235 & w47780) | (~w42235 & w47781) | (w47780 & w47781);
assign w27973 = ~w27970 & ~w27972;
assign w27974 = w26020 & w26880;
assign w27975 = ~w27952 & ~w27973;
assign w27976 = ~w27974 & ~w27975;
assign w27977 = ~w27958 & w45671;
assign w27978 = w27952 & ~w27977;
assign w27979 = (~w252 & ~w27976) | (~w252 & w45672) | (~w27976 & w45672);
assign w27980 = w252 & ~w27952;
assign w27981 = w252 & ~w26021;
assign w27982 = ~w27958 & w45673;
assign w27983 = ~w27980 & ~w27982;
assign w27984 = w27976 & ~w27983;
assign w27985 = w25966 & ~w26896;
assign w27986 = ~w26880 & w27985;
assign w27987 = ~w400 & ~w26078;
assign w27988 = ~w26879 & w27987;
assign w27989 = ~w25981 & ~w26022;
assign w27990 = w351 & w27989;
assign w27991 = (w27990 & w26879) | (w27990 & w45674) | (w26879 & w45674);
assign w27992 = ~w27986 & w27991;
assign w27993 = w351 & ~w27989;
assign w27994 = w25966 & w27993;
assign w27995 = w27994 & ~w26896;
assign w27996 = ~w26880 & w27995;
assign w27997 = ~w26879 & w45675;
assign w27998 = ~w27996 & ~w27997;
assign w27999 = ~w27992 & w27998;
assign w28000 = ~w27984 & ~w27999;
assign w28001 = ~w27979 & ~w28000;
assign w28002 = ~w27968 & w28001;
assign w28003 = ~w25925 & ~w25947;
assign w28004 = ~w27929 & ~w28003;
assign w28005 = ~w25946 & w26880;
assign w28006 = (w28004 & w26885) | (w28004 & w45677) | (w26885 & w45677);
assign w28007 = ~w26880 & w28006;
assign w28008 = ~w28005 & ~w28007;
assign w28009 = ~w27928 & w45678;
assign w28010 = w28008 & ~w28009;
assign w28011 = ~w80 & ~w28010;
assign w28012 = w57 & ~w27964;
assign w28013 = (w28012 & ~w27962) | (w28012 & w50102) | (~w27962 & w50102);
assign w28014 = w57 & w27964;
assign w28015 = w27962 & w50103;
assign w28016 = ~w28013 & ~w28015;
assign w28017 = ~w28011 & w28016;
assign w28018 = (w28017 & ~w28001) | (w28017 & w50104) | (~w28001 & w50104);
assign w28019 = w80 & w28010;
assign w28020 = ~w3 & ~w27935;
assign w28021 = (w28020 & w27932) | (w28020 & w45679) | (w27932 & w45679);
assign w28022 = ~w3 & w27935;
assign w28023 = ~w27932 & w45680;
assign w28024 = ~w28021 & ~w28023;
assign w28025 = ~w28019 & w28024;
assign w28026 = ~w27940 & w28025;
assign w28027 = ~w27986 & ~w27988;
assign w28028 = ~w351 & w27989;
assign w28029 = ~w28027 & w28028;
assign w28030 = ~w351 & ~w27989;
assign w28031 = w28027 & w28030;
assign w28032 = ~w28029 & ~w28031;
assign w28033 = ~w27984 & w28032;
assign w28034 = w28017 & w28033;
assign w28035 = w28026 & ~w28034;
assign w28036 = ~w28018 & w28035;
assign w28037 = w27949 & ~w28036;
assign w28038 = (w28026 & w28002) | (w28026 & w45681) | (w28002 & w45681);
assign w28039 = w27949 & ~w28038;
assign w28040 = ~w25851 & w26880;
assign w28041 = w25851 & ~w26880;
assign w28042 = ~w28040 & ~w28041;
assign w28043 = w27272 & w28042;
assign w28044 = ~w25851 & w28039;
assign w28045 = w28043 & ~w28044;
assign w28046 = ~w26880 & w28037;
assign w28047 = ~w27907 & w50105;
assign w28048 = w28045 & ~w28047;
assign w28049 = ~w27260 & w28038;
assign w28050 = (w28037 & w27260) | (w28037 & w45682) | (w27260 & w45682);
assign w28051 = (~w27651 & w27487) | (~w27651 & w42335) | (w27487 & w42335);
assign w28052 = (~w42335 & w45683) | (~w42335 & w45684) | (w45683 & w45684);
assign w28053 = ~w27823 & ~w27880;
assign w28054 = w27846 & w45685;
assign w28055 = ~w27884 & w28054;
assign w28056 = ~w28053 & ~w28055;
assign w28057 = ~w27743 & w27871;
assign w28058 = w27713 & ~w28057;
assign w28059 = (~w27723 & w28058) | (~w27723 & w45686) | (w28058 & w45686);
assign w28060 = ~w28056 & w28059;
assign w28061 = ~w27207 & w27901;
assign w28062 = ~w27903 & ~w28061;
assign w28063 = w27216 & w28062;
assign w28064 = w28060 & ~w28063;
assign w28065 = ~w28052 & w28064;
assign w28066 = w27849 & ~w28062;
assign w28067 = w27216 & ~w28066;
assign w28068 = ~w28065 & w28067;
assign w28069 = ~w28050 & ~w28068;
assign w28070 = w27258 & w28037;
assign w28071 = (~w28039 & ~w27258) | (~w28039 & w42336) | (~w27258 & w42336);
assign w28072 = ~a[22] & ~w26880;
assign w28073 = ~w28071 & ~w28072;
assign w28074 = ~w28069 & w28073;
assign w28075 = w27258 & w42337;
assign w28076 = ~w27906 & w28075;
assign w28077 = (~w28050 & ~w28075) | (~w28050 & w49159) | (~w28075 & w49159);
assign w28078 = w25851 & w26895;
assign w28079 = ~w28040 & ~w28078;
assign w28080 = ~w27271 & ~w28079;
assign w28081 = ~w25851 & ~w27271;
assign w28082 = w26880 & w28081;
assign w28083 = ~a[23] & ~w28082;
assign w28084 = a[22] & ~w28079;
assign w28085 = w28083 & ~w28084;
assign w28086 = (w28085 & w28076) | (w28085 & w49160) | (w28076 & w49160);
assign w28087 = ~w28074 & w28086;
assign w28088 = ~w27272 & ~w28072;
assign w28089 = ~w28040 & ~w28081;
assign w28090 = ~w28088 & ~w28089;
assign w28091 = ~w28068 & w50106;
assign w28092 = (~w42336 & w49161) | (~w42336 & w49162) | (w49161 & w49162);
assign w28093 = ~w28065 & w28092;
assign w28094 = (~w28050 & ~w28092) | (~w28050 & w45687) | (~w28092 & w45687);
assign w28095 = w27272 & w28078;
assign w28096 = a[23] & ~w28095;
assign w28097 = w28090 & w28071;
assign w28098 = w28096 & ~w28097;
assign w28099 = w28042 & w28088;
assign w28100 = ~w28076 & w42338;
assign w28101 = w28098 & ~w28100;
assign w28102 = w28072 & ~w28094;
assign w28103 = ~w28048 & w28087;
assign w28104 = w28101 & w49163;
assign w28105 = ~w28103 & ~w28104;
assign w28106 = a[22] & ~w27271;
assign w28107 = ~w27272 & ~w28106;
assign w28108 = ~w28050 & w28107;
assign w28109 = ~w28093 & w28108;
assign w28110 = ~w25851 & ~w28050;
assign w28111 = ~w28068 & w28110;
assign w28112 = a[22] & w26880;
assign w28113 = ~w28072 & ~w28112;
assign w28114 = (~w42336 & w45688) | (~w42336 & w45689) | (w45688 & w45689);
assign w28115 = (~w45689 & w50363) | (~w45689 & w50364) | (w50363 & w50364);
assign w28116 = ~w28093 & w45690;
assign w28117 = (w45689 & w50365) | (w45689 & w50366) | (w50365 & w50366);
assign w28118 = ~w28111 & w28117;
assign w28119 = ~w28116 & ~w28118;
assign w28120 = ~a[18] & ~a[19];
assign w28121 = ~a[20] & w28120;
assign w28122 = ~w26880 & w28121;
assign w28123 = w26880 & ~w28121;
assign w28124 = a[21] & w28123;
assign w28125 = ~w27271 & ~w28124;
assign w28126 = ~a[21] & ~w28123;
assign w28127 = ~w28122 & ~w28126;
assign w28128 = ~w28094 & w28127;
assign w28129 = ~w28122 & ~w28125;
assign w28130 = w28094 & w28129;
assign w28131 = ~w28128 & ~w28130;
assign w28132 = ~w28119 & w28131;
assign w28133 = w25851 & w28107;
assign w28134 = ~w28050 & w28133;
assign w28135 = ~w28093 & w28134;
assign w28136 = (w45689 & w50367) | (w45689 & w50368) | (w50367 & w50368);
assign w28137 = ~w28093 & w45691;
assign w28138 = (w45689 & w50369) | (w45689 & w50370) | (w50369 & w50370);
assign w28139 = ~w28069 & w28138;
assign w28140 = ~w28137 & ~w28139;
assign w28141 = w24874 & ~w27283;
assign w28142 = ~w24874 & w27283;
assign w28143 = ~w28141 & ~w28142;
assign w28144 = w28038 & w28143;
assign w28145 = (w27270 & w28076) | (w27270 & w42339) | (w28076 & w42339);
assign w28146 = ~w27270 & w28143;
assign w28147 = ~w28050 & w28146;
assign w28148 = ~w28093 & w28147;
assign w28149 = ~w28145 & ~w28148;
assign w28150 = (w23843 & w28148) | (w23843 & w45692) | (w28148 & w45692);
assign w28151 = w28140 & ~w28150;
assign w28152 = ~w28132 & w28151;
assign w28153 = ~w28105 & w28152;
assign w28154 = ~w28111 & ~w28115;
assign w28155 = ~w28109 & ~w28154;
assign w28156 = w28131 & ~w28155;
assign w28157 = ~w28069 & w28136;
assign w28158 = (~w24874 & w28093) | (~w24874 & w45693) | (w28093 & w45693);
assign w28159 = ~w28157 & w28158;
assign w28160 = (~w42336 & w49165) | (~w42336 & w49166) | (w49165 & w49166);
assign w28161 = (w28160 & w28068) | (w28160 & w50107) | (w28068 & w50107);
assign w28162 = w27327 & ~w27340;
assign w28163 = (w23843 & w27292) | (w23843 & w50108) | (w27292 & w50108);
assign w28164 = ~w27292 & w50109;
assign w28165 = ~w28163 & ~w28164;
assign w28166 = ~w27311 & w28165;
assign w28167 = ~w28163 & ~w28166;
assign w28168 = w28162 & ~w28167;
assign w28169 = ~w28162 & w28167;
assign w28170 = ~w28168 & ~w28169;
assign w28171 = ~w28036 & w49167;
assign w28172 = (w28170 & w28049) | (w28170 & w45694) | (w28049 & w45694);
assign w28173 = ~w27906 & w42340;
assign w28174 = w28172 & ~w28173;
assign w28175 = (w21801 & w28173) | (w21801 & w45695) | (w28173 & w45695);
assign w28176 = ~w28161 & w28175;
assign w28177 = ~w27384 & ~w28071;
assign w28178 = ~w28069 & w28177;
assign w28179 = ~w27330 & w27345;
assign w28180 = ~w21801 & w28179;
assign w28181 = w21801 & ~w28179;
assign w28182 = ~w28180 & ~w28181;
assign w28183 = w27384 & ~w28182;
assign w28184 = ~w28076 & w42341;
assign w28185 = ~w27384 & w28182;
assign w28186 = ~w20906 & ~w28185;
assign w28187 = (w28186 & w28076) | (w28186 & w49168) | (w28076 & w49168);
assign w28188 = ~w28178 & w28187;
assign w28189 = ~w28176 & ~w28188;
assign w28190 = ~w28148 & w45696;
assign w28191 = w28038 & w28166;
assign w28192 = ~w27260 & w28191;
assign w28193 = w27311 & ~w28165;
assign w28194 = (~w28193 & w28076) | (~w28193 & w42342) | (w28076 & w42342);
assign w28195 = (~w42336 & w49169) | (~w42336 & w49170) | (w49169 & w49170);
assign w28196 = (~w28076 & w49171) | (~w28076 & w49172) | (w49171 & w49172);
assign w28197 = (w49170 & w50371) | (w49170 & w50372) | (w50371 & w50372);
assign w28198 = ~w28069 & w28197;
assign w28199 = ~w28196 & ~w28198;
assign w28200 = ~w28190 & w28199;
assign w28201 = w28189 & w28200;
assign w28202 = ~w28150 & w28159;
assign w28203 = ~w28156 & w28202;
assign w28204 = w28201 & ~w28203;
assign w28205 = ~w28153 & w28204;
assign w28206 = ~w28184 & ~w28185;
assign w28207 = ~w28178 & w28206;
assign w28208 = w20906 & ~w28207;
assign w28209 = (w49166 & w50373) | (w49166 & w50374) | (w50373 & w50374);
assign w28210 = ~w28069 & w28209;
assign w28211 = ~w28173 & w45697;
assign w28212 = ~w28210 & ~w28211;
assign w28213 = (w28195 & w28068) | (w28195 & w50110) | (w28068 & w50110);
assign w28214 = (w28076 & w49173) | (w28076 & w49174) | (w49173 & w49174);
assign w28215 = ~w28213 & w28214;
assign w28216 = w28212 & ~w28215;
assign w28217 = w28189 & ~w28216;
assign w28218 = ~w28208 & ~w28217;
assign w28219 = ~w20906 & ~w28094;
assign w28220 = ~w27330 & w47782;
assign w28221 = w27426 & ~w28220;
assign w28222 = w27360 & w27434;
assign w28223 = w26520 & w26880;
assign w28224 = ~w26880 & w27355;
assign w28225 = ~w28223 & ~w28224;
assign w28226 = ~w28077 & ~w28225;
assign w28227 = ~w28221 & w28222;
assign w28228 = w28077 & w28227;
assign w28229 = ~w28226 & ~w28228;
assign w28230 = w28221 & ~w28222;
assign w28231 = ~w28219 & w28230;
assign w28232 = w28229 & ~w28231;
assign w28233 = ~w20000 & ~w28232;
assign w28234 = w28218 & ~w28233;
assign w28235 = ~w28205 & w28234;
assign w28236 = (~w27461 & w27388) | (~w27461 & w50111) | (w27388 & w50111);
assign w28237 = w27416 & ~w28236;
assign w28238 = ~w28076 & w42343;
assign w28239 = w27410 & ~w27411;
assign w28240 = ~w27410 & w27411;
assign w28241 = ~w28239 & ~w28240;
assign w28242 = ~w28238 & w28241;
assign w28243 = w27416 & w27466;
assign w28244 = w28236 & ~w28243;
assign w28245 = ~w28076 & w42344;
assign w28246 = ~w28236 & w28243;
assign w28247 = ~w28050 & w28246;
assign w28248 = ~w28093 & w28247;
assign w28249 = ~w28245 & ~w28248;
assign w28250 = ~w28242 & w28249;
assign w28251 = w28249 & w50112;
assign w28252 = w27435 & ~w28220;
assign w28253 = w27373 & ~w28252;
assign w28254 = w27455 & ~w28253;
assign w28255 = ~w28037 & ~w28254;
assign w28256 = w28038 & ~w28254;
assign w28257 = ~w27260 & w28256;
assign w28258 = ~w28255 & ~w28257;
assign w28259 = w19040 & w28037;
assign w28260 = ~w27257 & w42345;
assign w28261 = ~w28049 & w28259;
assign w28262 = w28259 & w28260;
assign w28263 = ~w27906 & w28262;
assign w28264 = ~w28261 & ~w28263;
assign w28265 = ~w28076 & ~w28258;
assign w28266 = w28264 & ~w28265;
assign w28267 = ~w27450 & ~w27461;
assign w28268 = w28266 & ~w28267;
assign w28269 = ~w28266 & w28267;
assign w28270 = ~w28268 & ~w28269;
assign w28271 = w18183 & w28270;
assign w28272 = (~w17380 & ~w28249) | (~w17380 & w50113) | (~w28249 & w50113);
assign w28273 = (~w28251 & w28271) | (~w28251 & w42346) | (w28271 & w42346);
assign w28274 = w27372 & w27455;
assign w28275 = w27360 & ~w28252;
assign w28276 = (w20000 & w28076) | (w20000 & w42347) | (w28076 & w42347);
assign w28277 = ~w28076 & w42348;
assign w28278 = ~w28276 & ~w28277;
assign w28279 = w28274 & w28278;
assign w28280 = ~w28274 & ~w28278;
assign w28281 = ~w28279 & ~w28280;
assign w28282 = w19040 & ~w28281;
assign w28283 = w20000 & w28232;
assign w28284 = ~w28282 & ~w28283;
assign w28285 = ~w28273 & w28284;
assign w28286 = ~w28235 & w28285;
assign w28287 = ~w19040 & w28281;
assign w28288 = ~w18183 & ~w28270;
assign w28289 = ~w28287 & ~w28288;
assign w28290 = ~w28251 & w28289;
assign w28291 = ~w28273 & ~w28290;
assign w28292 = ~w28286 & ~w28291;
assign w28293 = ~w27402 & ~w27636;
assign w28294 = w27416 & w28293;
assign w28295 = w27458 & w28294;
assign w28296 = ~w27388 & w28295;
assign w28297 = (~w27636 & w27468) | (~w27636 & w45698) | (w27468 & w45698);
assign w28298 = ~w28296 & ~w28297;
assign w28299 = (w27646 & w27616) | (w27646 & w49175) | (w27616 & w49175);
assign w28300 = w27600 & ~w28299;
assign w28301 = ~w27573 & ~w28300;
assign w28302 = w27600 & ~w27617;
assign w28303 = (w28301 & w28298) | (w28301 & w50114) | (w28298 & w50114);
assign w28304 = ~w27498 & ~w27602;
assign w28305 = w28303 & ~w28304;
assign w28306 = ~w28303 & w28304;
assign w28307 = ~w28305 & ~w28306;
assign w28308 = w27497 & ~w28077;
assign w28309 = (w50115 & w49159) | (w50115 & w50375) | (w49159 & w50375);
assign w28310 = ~w28308 & ~w28309;
assign w28311 = ~w11870 & w28310;
assign w28312 = ~w27513 & ~w27516;
assign w28313 = ~w27602 & ~w28303;
assign w28314 = ~w27498 & ~w28313;
assign w28315 = w28312 & ~w28314;
assign w28316 = (w27515 & w28076) | (w27515 & w42349) | (w28076 & w42349);
assign w28317 = w28077 & ~w28315;
assign w28318 = ~w28316 & ~w28317;
assign w28319 = ~w27498 & ~w28312;
assign w28320 = ~w28313 & w28319;
assign w28321 = w27515 & ~w28071;
assign w28322 = w28320 & ~w28321;
assign w28323 = ~w28050 & w28320;
assign w28324 = ~w28068 & w28323;
assign w28325 = ~w28322 & ~w28324;
assign w28326 = ~w28318 & w28325;
assign w28327 = (w11138 & w28318) | (w11138 & w42350) | (w28318 & w42350);
assign w28328 = ~w28311 & ~w28327;
assign w28329 = w11870 & ~w28310;
assign w28330 = ~w13384 & ~w27537;
assign w28331 = w13384 & w27537;
assign w28332 = ~w28330 & ~w28331;
assign w28333 = (w27585 & ~w27616) | (w27585 & w49176) | (~w27616 & w49176);
assign w28334 = ~w27537 & ~w27598;
assign w28335 = w28332 & ~w28334;
assign w28336 = w28333 & ~w28335;
assign w28337 = (w28336 & w28296) | (w28336 & w47783) | (w28296 & w47783);
assign w28338 = w27585 & ~w28299;
assign w28339 = w28334 & w28338;
assign w28340 = ~w27598 & w28330;
assign w28341 = w28333 & w28340;
assign w28342 = (w28341 & w28296) | (w28341 & w47784) | (w28296 & w47784);
assign w28343 = ~w13384 & w28339;
assign w28344 = ~w28342 & ~w28343;
assign w28345 = w28332 & ~w28339;
assign w28346 = ~w28337 & w28345;
assign w28347 = w28344 & ~w28346;
assign w28348 = ~w26880 & w27547;
assign w28349 = ~w26591 & ~w28348;
assign w28350 = w26591 & w28348;
assign w28351 = ~w28349 & ~w28350;
assign w28352 = (~w28351 & w28076) | (~w28351 & w49177) | (w28076 & w49177);
assign w28353 = w28347 & w28351;
assign w28354 = ~w28050 & w28353;
assign w28355 = ~w28068 & w28354;
assign w28356 = w28071 & w28353;
assign w28357 = ~w28355 & ~w28356;
assign w28358 = (~w12666 & ~w28357) | (~w12666 & w49178) | (~w28357 & w49178);
assign w28359 = ~w28329 & w28358;
assign w28360 = w28328 & ~w28359;
assign w28361 = ~w28318 & w50116;
assign w28362 = ~w27617 & ~w28298;
assign w28363 = w27649 & ~w28362;
assign w28364 = ~w27605 & ~w28363;
assign w28365 = ~w27634 & ~w27742;
assign w28366 = ~w28364 & ~w28365;
assign w28367 = ~w27633 & ~w28077;
assign w28368 = w28077 & w28366;
assign w28369 = ~w28367 & ~w28368;
assign w28370 = ~w27742 & ~w28051;
assign w28371 = (w28370 & w28094) | (w28370 & w50117) | (w28094 & w50117);
assign w28372 = w28369 & ~w28371;
assign w28373 = w28369 & w50118;
assign w28374 = ~w28361 & ~w28373;
assign w28375 = ~w28360 & w28374;
assign w28376 = ~w10419 & ~w28372;
assign w28377 = ~w27741 & ~w27870;
assign w28378 = ~w10419 & ~w28077;
assign w28379 = ~w27651 & w52268;
assign w28380 = w28379 & w28077;
assign w28381 = ~w28378 & ~w28380;
assign w28382 = w28377 & w28381;
assign w28383 = ~w28377 & ~w28381;
assign w28384 = ~w28382 & ~w28383;
assign w28385 = ~w9781 & ~w28384;
assign w28386 = ~w28376 & ~w28385;
assign w28387 = ~w28375 & w28386;
assign w28388 = w28357 & w50119;
assign w28389 = w27525 & ~w27526;
assign w28390 = ~w27525 & w27526;
assign w28391 = ~w28389 & ~w28390;
assign w28392 = ~w26580 & w26880;
assign w28393 = ~w26880 & ~w28391;
assign w28394 = ~w28392 & ~w28393;
assign w28395 = ~w28298 & w28333;
assign w28396 = ~w28338 & ~w28395;
assign w28397 = ~w28334 & w28396;
assign w28398 = w28397 & w50214;
assign w28399 = w28394 & ~w28077;
assign w28400 = ~w28398 & ~w28399;
assign w28401 = w28334 & ~w28396;
assign w28402 = (w28401 & w28094) | (w28401 & w50120) | (w28094 & w50120);
assign w28403 = w28400 & ~w28402;
assign w28404 = w28400 & w50121;
assign w28405 = ~w28388 & ~w28404;
assign w28406 = w28374 & w28405;
assign w28407 = ~w28329 & w28406;
assign w28408 = w14766 & w28038;
assign w28409 = ~w27260 & w28408;
assign w28410 = w26572 & w27580;
assign w28411 = ~w26572 & ~w27580;
assign w28412 = ~w28410 & ~w28411;
assign w28413 = (w28412 & w28076) | (w28412 & w42353) | (w28076 & w42353);
assign w28414 = w28396 & w28077;
assign w28415 = ~w28413 & ~w28414;
assign w28416 = w27585 & w27646;
assign w28417 = ~w27641 & ~w28416;
assign w28418 = ~w28362 & w28417;
assign w28419 = (~w49180 & w50377) | (~w49180 & w50378) | (w50377 & w50378);
assign w28420 = ~w28050 & w28418;
assign w28421 = ~w28068 & w28420;
assign w28422 = ~w28419 & ~w28421;
assign w28423 = ~w28415 & w28422;
assign w28424 = (~w14039 & w28415) | (~w14039 & w42354) | (w28415 & w42354);
assign w28425 = (w13384 & ~w28400) | (w13384 & w50122) | (~w28400 & w50122);
assign w28426 = ~w28424 & ~w28425;
assign w28427 = w15681 & ~w27636;
assign w28428 = (w28427 & w27468) | (w28427 & w50123) | (w27468 & w50123);
assign w28429 = (~w15681 & w27388) | (~w15681 & w42355) | (w27388 & w42355);
assign w28430 = ~w28297 & w28429;
assign w28431 = ~w27388 & w42356;
assign w28432 = ~w28428 & ~w28431;
assign w28433 = ~w28430 & w28432;
assign w28434 = w28038 & ~w28433;
assign w28435 = ~w27260 & w28434;
assign w28436 = (w27616 & w28076) | (w27616 & w42357) | (w28076 & w42357);
assign w28437 = ~w28076 & w42358;
assign w28438 = ~w28436 & ~w28437;
assign w28439 = ~w14766 & w28438;
assign w28440 = ~w28415 & w42359;
assign w28441 = ~w28439 & ~w28440;
assign w28442 = ~w27468 & ~w27484;
assign w28443 = ~w27460 & w28442;
assign w28444 = w16559 & w28443;
assign w28445 = w28038 & ~w28444;
assign w28446 = ~w27260 & w28445;
assign w28447 = (~w27482 & w28076) | (~w27482 & w42360) | (w28076 & w42360);
assign w28448 = ~w16559 & w27487;
assign w28449 = ~w28050 & w28448;
assign w28450 = ~w28093 & w28449;
assign w28451 = ~w28447 & ~w28450;
assign w28452 = w27636 & ~w28443;
assign w28453 = ~w28037 & w28452;
assign w28454 = w28038 & w28452;
assign w28455 = ~w27260 & w28454;
assign w28456 = w27483 & ~w28443;
assign w28457 = (~w28456 & w28076) | (~w28456 & w42361) | (w28076 & w42361);
assign w28458 = w28451 & w28457;
assign w28459 = (~w15681 & ~w28451) | (~w15681 & w45699) | (~w28451 & w45699);
assign w28460 = ~w27402 & ~w27484;
assign w28461 = w27466 & ~w28237;
assign w28462 = w28460 & ~w28461;
assign w28463 = (~w42336 & w49181) | (~w42336 & w49182) | (w49181 & w49182);
assign w28464 = w28462 & ~w28463;
assign w28465 = ~w28050 & w28462;
assign w28466 = ~w28068 & w28465;
assign w28467 = ~w28464 & ~w28466;
assign w28468 = (~w27401 & w28076) | (~w27401 & w42362) | (w28076 & w42362);
assign w28469 = ~w28460 & w28461;
assign w28470 = ~w28076 & w42363;
assign w28471 = ~w28468 & ~w28470;
assign w28472 = w28467 & w28471;
assign w28473 = w16559 & ~w28472;
assign w28474 = ~w28459 & w28473;
assign w28475 = (w42361 & w45700) | (w42361 & w45701) | (w45700 & w45701);
assign w28476 = w28451 & w28475;
assign w28477 = w14766 & ~w28438;
assign w28478 = ~w28476 & ~w28477;
assign w28479 = (~w28424 & w28439) | (~w28424 & w50180) | (w28439 & w50180);
assign w28480 = ~w28424 & w28478;
assign w28481 = ~w28474 & w28480;
assign w28482 = ~w28479 & ~w28481;
assign w28483 = (w28426 & w28481) | (w28426 & w45702) | (w28481 & w45702);
assign w28484 = w28407 & ~w28483;
assign w28485 = w28387 & ~w28484;
assign w28486 = ~w28292 & w28485;
assign w28487 = w9781 & w28384;
assign w28488 = ~w27689 & ~w27869;
assign w28489 = w27743 & w28051;
assign w28490 = ~w27870 & ~w28489;
assign w28491 = (w9781 & w28076) | (w9781 & w42364) | (w28076 & w42364);
assign w28492 = ~w28076 & w42365;
assign w28493 = ~w28491 & ~w28492;
assign w28494 = w28488 & w28493;
assign w28495 = ~w28488 & ~w28493;
assign w28496 = ~w28494 & ~w28495;
assign w28497 = ~w9195 & ~w28496;
assign w28498 = ~w28487 & ~w28497;
assign w28499 = w28387 & ~w28407;
assign w28500 = (w28498 & ~w28387) | (w28498 & w50124) | (~w28387 & w50124);
assign w28501 = w28471 & w49183;
assign w28502 = ~w28459 & ~w28501;
assign w28503 = w28478 & ~w28502;
assign w28504 = w28441 & ~w28503;
assign w28505 = (w28426 & w28503) | (w28426 & w50125) | (w28503 & w50125);
assign w28506 = w28387 & w28505;
assign w28507 = (~w27874 & w27640) | (~w27874 & w42366) | (w27640 & w42366);
assign w28508 = ~w27880 & ~w27883;
assign w28509 = w27785 & ~w27831;
assign w28510 = (~w45704 & w47785) | (~w45704 & w47786) | (w47785 & w47786);
assign w28511 = (w47785 & w49184) | (w47785 & w49185) | (w49184 & w49185);
assign w28512 = w27822 & ~w27847;
assign w28513 = ~w28076 & w42367;
assign w28514 = ~w28076 & w49186;
assign w28515 = w27807 & w27900;
assign w28516 = ~w4430 & w28515;
assign w28517 = (~w28076 & w49187) | (~w28076 & w49188) | (w49187 & w49188);
assign w28518 = ~w28514 & w28517;
assign w28519 = ~w4430 & ~w28515;
assign w28520 = ~w28511 & w28519;
assign w28521 = w28513 & w28520;
assign w28522 = (w28076 & w49189) | (w28076 & w49190) | (w49189 & w49190);
assign w28523 = ~w28521 & ~w28522;
assign w28524 = ~w28518 & w28523;
assign w28525 = w27837 & ~w28510;
assign w28526 = w28077 & w28525;
assign w28527 = w27822 & w27846;
assign w28528 = w4838 & ~w28527;
assign w28529 = (w28528 & w28526) | (w28528 & w42368) | (w28526 & w42368);
assign w28530 = w4838 & w28527;
assign w28531 = ~w28526 & w42369;
assign w28532 = ~w28529 & ~w28531;
assign w28533 = w28524 & w28532;
assign w28534 = w4430 & ~w28515;
assign w28535 = (~w28076 & w49191) | (~w28076 & w49192) | (w49191 & w49192);
assign w28536 = ~w28514 & w28535;
assign w28537 = w4430 & w28515;
assign w28538 = ~w28511 & w28537;
assign w28539 = w28513 & w28538;
assign w28540 = (w28076 & w49193) | (w28076 & w49194) | (w49193 & w49194);
assign w28541 = ~w28539 & ~w28540;
assign w28542 = ~w28536 & w28541;
assign w28543 = ~w28526 & w42370;
assign w28544 = (w28527 & w28526) | (w28527 & w42371) | (w28526 & w42371);
assign w28545 = ~w28543 & ~w28544;
assign w28546 = ~w4838 & ~w28545;
assign w28547 = (~w5745 & w28076) | (~w5745 & w42372) | (w28076 & w42372);
assign w28548 = (~w45704 & w47787) | (~w45704 & w47788) | (w47787 & w47788);
assign w28549 = ~w28076 & w42373;
assign w28550 = ~w28547 & ~w28549;
assign w28551 = ~w27831 & w27837;
assign w28552 = w5330 & ~w28551;
assign w28553 = ~w28550 & w28552;
assign w28554 = w5330 & w28551;
assign w28555 = w28550 & w28554;
assign w28556 = ~w28553 & ~w28555;
assign w28557 = ~w28533 & w28542;
assign w28558 = w28542 & w28556;
assign w28559 = ~w28546 & w28558;
assign w28560 = ~w28557 & ~w28559;
assign w28561 = (~w27260 & w28065) | (~w27260 & w50126) | (w28065 & w50126);
assign w28562 = (w27871 & w27651) | (w27871 & w28057) | (w27651 & w28057);
assign w28563 = w27638 & w27871;
assign w28564 = ~w27605 & w28563;
assign w28565 = ~w27689 & ~w27710;
assign w28566 = (w28565 & w27487) | (w28565 & w42374) | (w27487 & w42374);
assign w28567 = ~w27671 & w27701;
assign w28568 = (w27862 & ~w28566) | (w27862 & w50127) | (~w28566 & w50127);
assign w28569 = w28567 & ~w28568;
assign w28570 = w27851 & ~w28039;
assign w28571 = ~w27723 & ~w28570;
assign w28572 = w27856 & ~w28571;
assign w28573 = ~w28569 & w28572;
assign w28574 = ~w7315 & w28070;
assign w28575 = ~w28561 & w28574;
assign w28576 = w28573 & ~w28575;
assign w28577 = ~w28076 & w42375;
assign w28578 = (w27722 & w28076) | (w27722 & w49195) | (w28076 & w49195);
assign w28579 = ~w28577 & ~w28578;
assign w28580 = (~w6769 & w28579) | (~w6769 & w50128) | (w28579 & w50128);
assign w28581 = ~w6264 & w27882;
assign w28582 = ~w27883 & ~w28581;
assign w28583 = ~w28582 & w50215;
assign w28584 = (w47789 & w49196) | (w47789 & w49197) | (w49196 & w49197);
assign w28585 = ~w27882 & ~w28077;
assign w28586 = w28077 & w42377;
assign w28587 = ~w28585 & ~w28586;
assign w28588 = (~w5745 & w28586) | (~w5745 & w50129) | (w28586 & w50129);
assign w28589 = (~w6769 & w28076) | (~w6769 & w42378) | (w28076 & w42378);
assign w28590 = ~w28577 & ~w28589;
assign w28591 = w27779 & ~w27880;
assign w28592 = w6264 & ~w28591;
assign w28593 = ~w6264 & w28591;
assign w28594 = ~w28592 & ~w28593;
assign w28595 = ~w28577 & w49667;
assign w28596 = (w28594 & w28577) | (w28594 & w49668) | (w28577 & w49668);
assign w28597 = ~w28595 & ~w28596;
assign w28598 = ~w28586 & w50130;
assign w28599 = ~w6264 & ~w28591;
assign w28600 = ~w28577 & w49669;
assign w28601 = (w28593 & w28577) | (w28593 & w49670) | (w28577 & w49670);
assign w28602 = ~w28600 & ~w28601;
assign w28603 = (~w28598 & w28602) | (~w28598 & w49198) | (w28602 & w49198);
assign w28604 = ~w28588 & ~w28597;
assign w28605 = ~w28580 & w28604;
assign w28606 = w28603 & ~w28605;
assign w28607 = ~w28560 & ~w28606;
assign w28608 = w27701 & w27856;
assign w28609 = ~w27671 & ~w27861;
assign w28610 = w28565 & w28609;
assign w28611 = (w28610 & w27487) | (w28610 & w42379) | (w27487 & w42379);
assign w28612 = w27859 & w28609;
assign w28613 = (~w28612 & ~w28611) | (~w28612 & w49199) | (~w28611 & w49199);
assign w28614 = ~w27861 & w28613;
assign w28615 = w28613 & w49671;
assign w28616 = w28608 & ~w28614;
assign w28617 = ~w7924 & w27856;
assign w28618 = w27701 & ~w28617;
assign w28619 = ~w28077 & w28618;
assign w28620 = w28077 & ~w28615;
assign w28621 = ~w28616 & w28620;
assign w28622 = ~w28619 & ~w28621;
assign w28623 = w7315 & w28622;
assign w28624 = ~w27859 & ~w28609;
assign w28625 = (w28624 & ~w28566) | (w28624 & w49672) | (~w28566 & w49672);
assign w28626 = w28613 & ~w28625;
assign w28627 = w27670 & ~w28077;
assign w28628 = w28077 & w28626;
assign w28629 = ~w28627 & ~w28628;
assign w28630 = w7924 & w28629;
assign w28631 = (w27216 & w27876) | (w27216 & w42380) | (w27876 & w42380);
assign w28632 = ~w28050 & ~w28631;
assign w28633 = ~w27858 & ~w28071;
assign w28634 = (~w27689 & w27487) | (~w27689 & w47791) | (w27487 & w47791);
assign w28635 = ~w27710 & ~w27859;
assign w28636 = (~w28635 & ~w28634) | (~w28635 & w49673) | (~w28634 & w49673);
assign w28637 = ~w28632 & w28633;
assign w28638 = ~w28076 & w42381;
assign w28639 = ~w28637 & ~w28638;
assign w28640 = w28566 & w49674;
assign w28641 = ~w28633 & w28640;
assign w28642 = ~w28050 & w28640;
assign w28643 = ~w28068 & w28642;
assign w28644 = ~w28641 & ~w28643;
assign w28645 = ~w28639 & w28644;
assign w28646 = ~w7924 & w27670;
assign w28647 = (w28646 & w28076) | (w28646 & w42382) | (w28076 & w42382);
assign w28648 = ~w7924 & w28626;
assign w28649 = w28077 & w28648;
assign w28650 = ~w28647 & ~w28649;
assign w28651 = ~w28649 & w42383;
assign w28652 = ~w28645 & w28651;
assign w28653 = ~w28630 & ~w28652;
assign w28654 = ~w28623 & w28653;
assign w28655 = (~w7315 & w28621) | (~w7315 & w49675) | (w28621 & w49675);
assign w28656 = ~w28579 & w50131;
assign w28657 = ~w28655 & ~w28656;
assign w28658 = w28603 & w28657;
assign w28659 = ~w28654 & w28658;
assign w28660 = w28607 & ~w28659;
assign w28661 = ~w28506 & w28660;
assign w28662 = w28500 & w28661;
assign w28663 = ~w28486 & w28662;
assign w28664 = w28550 & ~w28551;
assign w28665 = ~w28550 & w28551;
assign w28666 = ~w28664 & ~w28665;
assign w28667 = ~w5330 & ~w28666;
assign w28668 = w28533 & ~w28667;
assign w28669 = ~w28560 & ~w28668;
assign w28670 = ~w28639 & w47792;
assign w28671 = w9195 & ~w28488;
assign w28672 = ~w28492 & w49676;
assign w28673 = w9195 & w28488;
assign w28674 = (w28673 & w28492) | (w28673 & w49677) | (w28492 & w49677);
assign w28675 = ~w28672 & ~w28674;
assign w28676 = ~w28670 & w28675;
assign w28677 = w28650 & w28676;
assign w28678 = w28654 & ~w28677;
assign w28679 = (w28658 & ~w28654) | (w28658 & w50132) | (~w28654 & w50132);
assign w28680 = w28607 & ~w28679;
assign w28681 = (~w28669 & w28679) | (~w28669 & w47793) | (w28679 & w47793);
assign w28682 = ~w28663 & w28681;
assign w28683 = w27216 & w28032;
assign w28684 = w27258 & w49200;
assign w28685 = ~w27259 & w28032;
assign w28686 = w27258 & w28685;
assign w28687 = ~w28684 & ~w28686;
assign w28688 = ~w28686 & w28065;
assign w28689 = ~w28687 & ~w28688;
assign w28690 = (w27999 & w28036) | (w27999 & w49678) | (w28036 & w49678);
assign w28691 = w27999 & w28038;
assign w28692 = (~w28690 & w27260) | (~w28690 & w50379) | (w27260 & w50379);
assign w28693 = ~w28076 & ~w28692;
assign w28694 = ~w28689 & w28693;
assign w28695 = (w252 & w28076) | (w252 & w42384) | (w28076 & w42384);
assign w28696 = ~w27979 & ~w27984;
assign w28697 = w57 & ~w28696;
assign w28698 = (w28697 & w28694) | (w28697 & w49201) | (w28694 & w49201);
assign w28699 = w57 & w28696;
assign w28700 = ~w28694 & w49202;
assign w28701 = ~w28698 & ~w28700;
assign w28702 = w27999 & w28032;
assign w28703 = ~w28037 & ~w28702;
assign w28704 = w28038 & ~w28702;
assign w28705 = ~w27260 & w28704;
assign w28706 = ~w28703 & ~w28705;
assign w28707 = ~w28076 & ~w28706;
assign w28708 = ~w27908 & w28707;
assign w28709 = w27989 & ~w28027;
assign w28710 = ~w27989 & w28027;
assign w28711 = ~w28709 & ~w28710;
assign w28712 = (~w28711 & w28076) | (~w28711 & w42385) | (w28076 & w42385);
assign w28713 = ~w28708 & ~w28712;
assign w28714 = w28077 & w42386;
assign w28715 = (w252 & ~w28713) | (w252 & w42387) | (~w28713 & w42387);
assign w28716 = ~w26906 & ~w26907;
assign w28717 = ~w26974 & ~w26994;
assign w28718 = ~w26940 & ~w26976;
assign w28719 = ~w26940 & ~w28717;
assign w28720 = (~w28718 & w27256) | (~w28718 & w42388) | (w27256 & w42388);
assign w28721 = w27216 & w28720;
assign w28722 = ~w28066 & w28721;
assign w28723 = ~w27086 & w27239;
assign w28724 = w27006 & ~w28723;
assign w28725 = ~w28723 & w42389;
assign w28726 = ~w28723 & w45707;
assign w28727 = w28720 & ~w28726;
assign w28728 = ~w28722 & ~w28727;
assign w28729 = ~w28052 & ~w28727;
assign w28730 = w28064 & w28729;
assign w28731 = ~w28728 & ~w28730;
assign w28732 = ~w28716 & ~w28731;
assign w28733 = w28716 & w28731;
assign w28734 = w28077 & ~w28733;
assign w28735 = ~w26905 & ~w28077;
assign w28736 = ~w351 & ~w28735;
assign w28737 = ~w28732 & w28734;
assign w28738 = w28736 & ~w28737;
assign w28739 = ~w28715 & ~w28738;
assign w28740 = w351 & w28735;
assign w28741 = (w351 & w28731) | (w351 & w45708) | (w28731 & w45708);
assign w28742 = w28734 & w28741;
assign w28743 = ~w28740 & ~w28742;
assign w28744 = ~w26938 & w28725;
assign w28745 = ~w28067 & w28744;
assign w28746 = (~w28745 & ~w28075) | (~w28745 & w49203) | (~w28075 & w49203);
assign w28747 = (~w26975 & w27256) | (~w26975 & w42390) | (w27256 & w42390);
assign w28748 = ~w28037 & w28747;
assign w28749 = w28038 & w28747;
assign w28750 = ~w27260 & w28749;
assign w28751 = ~w28748 & ~w28750;
assign w28752 = ~w28052 & w28744;
assign w28753 = w28064 & w28752;
assign w28754 = ~w28751 & ~w28753;
assign w28755 = (w493 & w28076) | (w493 & w42391) | (w28076 & w42391);
assign w28756 = w28746 & w28754;
assign w28757 = ~w28755 & ~w28756;
assign w28758 = ~w26920 & ~w26922;
assign w28759 = ~w400 & ~w28758;
assign w28760 = (w28759 & w28756) | (w28759 & w42392) | (w28756 & w42392);
assign w28761 = ~w400 & w28758;
assign w28762 = ~w28756 & w42393;
assign w28763 = ~w28760 & ~w28762;
assign w28764 = w28743 & w28763;
assign w28765 = w28739 & ~w28764;
assign w28766 = w28713 & w49204;
assign w28767 = ~w57 & w52269;
assign w28768 = ~w28694 & w49679;
assign w28769 = w28767 & ~w28768;
assign w28770 = (w28701 & w28765) | (w28701 & w45709) | (w28765 & w45709);
assign w28771 = (w26991 & w28076) | (w26991 & w42395) | (w28076 & w42395);
assign w28772 = ~w27881 & w28724;
assign w28773 = w27904 & w28772;
assign w28774 = ~w27876 & w28773;
assign w28775 = (w27248 & w27876) | (w27248 & w42396) | (w27876 & w42396);
assign w28776 = ~w26992 & ~w27249;
assign w28777 = w28775 & ~w28776;
assign w28778 = ~w28775 & w28776;
assign w28779 = w28077 & w42397;
assign w28780 = (~w28771 & ~w42397) | (~w28771 & w49680) | (~w42397 & w49680);
assign w28781 = ~w754 & ~w28780;
assign w28782 = w27006 & w27245;
assign w28783 = w27216 & w27239;
assign w28784 = ~w28723 & w52270;
assign w28785 = ~w28723 & w28782;
assign w28786 = w28785 & w52270;
assign w28787 = w28077 & ~w28786;
assign w28788 = ~w28782 & ~w28784;
assign w28789 = w28787 & ~w28788;
assign w28790 = w27000 & ~w27001;
assign w28791 = ~w27000 & w27001;
assign w28792 = ~w28790 & ~w28791;
assign w28793 = (~w28792 & w28076) | (~w28792 & w42399) | (w28076 & w42399);
assign w28794 = ~w945 & ~w28793;
assign w28795 = ~w28789 & w28794;
assign w28796 = w754 & ~w28771;
assign w28797 = ~w28779 & w28796;
assign w28798 = ~w28795 & ~w28797;
assign w28799 = ~w28781 & ~w28798;
assign w28800 = w27248 & ~w27249;
assign w28801 = (~w26992 & w28774) | (~w26992 & w49681) | (w28774 & w49681);
assign w28802 = ~w26974 & ~w26993;
assign w28803 = w26973 & ~w28071;
assign w28804 = ~w28802 & ~w28803;
assign w28805 = ~w28050 & ~w28802;
assign w28806 = ~w28068 & w28805;
assign w28807 = ~w28804 & ~w28806;
assign w28808 = w28801 & ~w28807;
assign w28809 = w27248 & w27254;
assign w28810 = ~w26974 & w26992;
assign w28811 = (~w28810 & w28774) | (~w28810 & w42400) | (w28774 & w42400);
assign w28812 = w28077 & w28811;
assign w28813 = (~w754 & w28036) | (~w754 & w49682) | (w28036 & w49682);
assign w28814 = ~w754 & w28038;
assign w28815 = ~w27260 & w28814;
assign w28816 = (w26973 & w28076) | (w26973 & w42401) | (w28076 & w42401);
assign w28817 = ~w28812 & ~w28816;
assign w28818 = (w612 & w28812) | (w612 & w42402) | (w28812 & w42402);
assign w28819 = ~w28808 & w28818;
assign w28820 = ~w26938 & ~w26975;
assign w28821 = (~w28717 & w27240) | (~w28717 & w50133) | (w27240 & w50133);
assign w28822 = ~w28725 & ~w28821;
assign w28823 = w27216 & ~w28821;
assign w28824 = ~w28066 & w28823;
assign w28825 = ~w28822 & ~w28824;
assign w28826 = ~w28052 & ~w28822;
assign w28827 = w28064 & w28826;
assign w28828 = ~w28825 & ~w28827;
assign w28829 = ~w28820 & w28828;
assign w28830 = (w28820 & w28827) | (w28820 & w50134) | (w28827 & w50134);
assign w28831 = w28077 & ~w28830;
assign w28832 = w26937 & ~w28077;
assign w28833 = w493 & ~w28832;
assign w28834 = ~w28829 & w28831;
assign w28835 = w28833 & ~w28834;
assign w28836 = ~w28819 & ~w28835;
assign w28837 = ~w28799 & w28836;
assign w28838 = ~w612 & w28801;
assign w28839 = ~w28807 & w28838;
assign w28840 = ~w28812 & w42403;
assign w28841 = ~w28839 & ~w28840;
assign w28842 = ~w493 & w28832;
assign w28843 = (~w493 & ~w28828) | (~w493 & w49683) | (~w28828 & w49683);
assign w28844 = w28831 & w28843;
assign w28845 = ~w28842 & ~w28844;
assign w28846 = w28841 & w28845;
assign w28847 = ~w28835 & ~w28846;
assign w28848 = w400 & ~w28758;
assign w28849 = ~w28756 & w49684;
assign w28850 = w400 & w28758;
assign w28851 = (w28850 & w28756) | (w28850 & w49685) | (w28756 & w49685);
assign w28852 = ~w28849 & ~w28851;
assign w28853 = w28701 & w28852;
assign w28854 = w28739 & w28853;
assign w28855 = ~w28837 & ~w28847;
assign w28856 = w28854 & w28855;
assign w28857 = ~w28770 & ~w28856;
assign w28858 = ~w28002 & w28016;
assign w28859 = ~w27984 & w28016;
assign w28860 = (~w28858 & ~w28689) | (~w28858 & w42404) | (~w28689 & w42404);
assign w28861 = w28010 & ~w28077;
assign w28862 = ~w28011 & ~w28019;
assign w28863 = ~w28076 & w42405;
assign w28864 = ~w28861 & ~w28863;
assign w28865 = w28860 & ~w28864;
assign w28866 = (w28010 & w28076) | (w28010 & w49205) | (w28076 & w49205);
assign w28867 = w28011 & w28094;
assign w28868 = ~w28866 & ~w28867;
assign w28869 = ~w28860 & ~w28868;
assign w28870 = ~w28865 & ~w28869;
assign w28871 = (~w3 & w28869) | (~w3 & w49686) | (w28869 & w49686);
assign w28872 = (w3 & w28864) | (w3 & w42406) | (w28864 & w42406);
assign w28873 = ~w28869 & w28872;
assign w28874 = ~w28076 & w42407;
assign w28875 = ~w27984 & w28689;
assign w28876 = w28874 & ~w28875;
assign w28877 = ~w27968 & w28016;
assign w28878 = w80 & w28877;
assign w28879 = (w28878 & w28876) | (w28878 & w42408) | (w28876 & w42408);
assign w28880 = w80 & ~w28877;
assign w28881 = ~w28876 & w42409;
assign w28882 = ~w28879 & ~w28881;
assign w28883 = ~w28873 & ~w28882;
assign w28884 = ~w28871 & ~w28883;
assign w28885 = ~w28018 & ~w28034;
assign w28886 = (w28002 & w27907) | (w28002 & w45710) | (w27907 & w45710);
assign w28887 = ~w28885 & ~w28886;
assign w28888 = w3 & ~w28077;
assign w28889 = ~w28050 & w50216;
assign w28890 = ~w28887 & w28889;
assign w28891 = ~w28888 & ~w28890;
assign w28892 = ~w27939 & w28024;
assign w28893 = ~w27939 & ~w28025;
assign w28894 = ~w27939 & ~w28885;
assign w28895 = (~w28893 & w28886) | (~w28893 & w49688) | (w28886 & w49688);
assign w28896 = w42 & ~w27924;
assign w28897 = ~w27915 & w27924;
assign w28898 = ~w42 & w28897;
assign w28899 = ~w28896 & ~w28898;
assign w28900 = w28895 & ~w28899;
assign w28901 = ~w27946 & ~w28896;
assign w28902 = ~w28895 & w28901;
assign w28903 = ~w28900 & ~w28902;
assign w28904 = w42 & ~w28892;
assign w28905 = (w28904 & w28890) | (w28904 & w49689) | (w28890 & w49689);
assign w28906 = w28903 & ~w28905;
assign w28907 = w42 & w28892;
assign w28908 = w28891 & w28907;
assign w28909 = w28906 & ~w28908;
assign w28910 = w28891 & ~w28892;
assign w28911 = ~w28891 & w28892;
assign w28912 = ~w28910 & ~w28911;
assign w28913 = w28895 & w28897;
assign w28914 = ~w42 & ~w28913;
assign w28915 = ~w27924 & ~w28895;
assign w28916 = w28914 & ~w28915;
assign w28917 = ~w28884 & w28909;
assign w28918 = ~w28912 & w28916;
assign w28919 = ~w28917 & ~w28918;
assign w28920 = w28857 & w28919;
assign w28921 = ~w27967 & ~w28077;
assign w28922 = ~w80 & ~w28921;
assign w28923 = ~w28875 & w42410;
assign w28924 = w28077 & ~w28877;
assign w28925 = ~w28876 & w28924;
assign w28926 = ~w28925 & w42411;
assign w28927 = ~w28873 & ~w28926;
assign w28928 = ~w28871 & ~w28927;
assign w28929 = w28909 & ~w28928;
assign w28930 = w28919 & ~w28929;
assign w28931 = ~w28920 & ~w28930;
assign w28932 = (~w28793 & ~w28787) | (~w28793 & w49690) | (~w28787 & w49690);
assign w28933 = w945 & ~w28932;
assign w28934 = ~w28781 & ~w28933;
assign w28935 = w28846 & w28934;
assign w28936 = w28854 & w28935;
assign w28937 = ~w28856 & w42412;
assign w28938 = ~w28930 & ~w28937;
assign w28939 = w27084 & ~w28631;
assign w28940 = w27026 & w27051;
assign w28941 = w28939 & w28940;
assign w28942 = w27224 & w28940;
assign w28943 = w27232 & ~w28942;
assign w28944 = ~w28076 & w42413;
assign w28945 = ~w28941 & w28944;
assign w28946 = w1320 & ~w28077;
assign w28947 = w27070 & ~w27235;
assign w28948 = ~w28945 & w49206;
assign w28949 = (w28947 & w28945) | (w28947 & w49207) | (w28945 & w49207);
assign w28950 = ~w28948 & ~w28949;
assign w28951 = w1120 & ~w28950;
assign w28952 = ~w27020 & ~w27021;
assign w28953 = w27020 & w27021;
assign w28954 = ~w28952 & ~w28953;
assign w28955 = w27224 & w28071;
assign w28956 = w27026 & ~w28955;
assign w28957 = ~w28939 & ~w28956;
assign w28958 = ~w1738 & w28954;
assign w28959 = ~w28631 & w45711;
assign w28960 = ~w28957 & ~w28959;
assign w28961 = ~w2341 & ~w27211;
assign w28962 = ~w28954 & ~w28961;
assign w28963 = ~w1738 & w27211;
assign w28964 = w28962 & ~w28963;
assign w28965 = (w28954 & w28076) | (w28954 & w42414) | (w28076 & w42414);
assign w28966 = ~w28631 & w47794;
assign w28967 = ~w28965 & ~w28966;
assign w28968 = (w1541 & ~w28960) | (w1541 & w49691) | (~w28960 & w49691);
assign w28969 = w28960 & w49692;
assign w28970 = w27084 & ~w27212;
assign w28971 = ~w27208 & ~w27213;
assign w28972 = ~w27200 & w28971;
assign w28973 = ~w28066 & w28972;
assign w28974 = w28060 & ~w28062;
assign w28975 = ~w28052 & w28974;
assign w28976 = (w28970 & w28975) | (w28970 & w47795) | (w28975 & w47795);
assign w28977 = ~w28975 & w47796;
assign w28978 = ~w28976 & ~w28977;
assign w28979 = (w27211 & w28076) | (w27211 & w45712) | (w28076 & w45712);
assign w28980 = w28077 & w28978;
assign w28981 = ~w28979 & ~w28980;
assign w28982 = (~w1738 & w28980) | (~w1738 & w45713) | (w28980 & w45713);
assign w28983 = ~w28969 & ~w28982;
assign w28984 = ~w28968 & ~w28983;
assign w28985 = w27051 & w27232;
assign w28986 = ~w27224 & ~w28985;
assign w28987 = w45714 & ~w28631;
assign w28988 = w28986 & ~w28987;
assign w28989 = w27051 & ~w28094;
assign w28990 = w28988 & ~w28989;
assign w28991 = ~w26880 & w27040;
assign w28992 = ~w27043 & ~w28991;
assign w28993 = w27043 & w28991;
assign w28994 = ~w28992 & ~w28993;
assign w28995 = (w28994 & w28076) | (w28994 & w49208) | (w28076 & w49208);
assign w28996 = ~w28945 & ~w28995;
assign w28997 = ~w28990 & ~w28996;
assign w28998 = ~w28996 & w49209;
assign w28999 = ~w28980 & w45715;
assign w29000 = ~w28968 & ~w28999;
assign w29001 = ~w28998 & ~w29000;
assign w29002 = ~w28984 & w29001;
assign w29003 = w1320 & ~w28997;
assign w29004 = ~w1120 & w28950;
assign w29005 = ~w29003 & ~w29004;
assign w29006 = (~w28951 & w29002) | (~w28951 & w49210) | (w29002 & w49210);
assign w29007 = ~w28984 & ~w28998;
assign w29008 = ~w28984 & w49211;
assign w29009 = (w27900 & w28055) | (w27900 & w47797) | (w28055 & w47797);
assign w29010 = w28059 & w29009;
assign w29011 = (w27179 & w27893) | (w27179 & w45716) | (w27893 & w45716);
assign w29012 = w28059 & w47798;
assign w29013 = ~w28052 & w29012;
assign w29014 = (~w27202 & w27141) | (~w27202 & w47775) | (w27141 & w47775);
assign w29015 = w27179 & ~w29014;
assign w29016 = ~w27204 & ~w29015;
assign w29017 = (w27900 & ~w27823) | (w27900 & w49693) | (~w27823 & w49693);
assign w29018 = ~w27833 & w29017;
assign w29019 = ~w27191 & ~w27203;
assign w29020 = (w29019 & ~w29018) | (w29019 & w45717) | (~w29018 & w45717);
assign w29021 = w29016 & w29020;
assign w29022 = (~w27191 & w29013) | (~w27191 & w45718) | (w29013 & w45718);
assign w29023 = ~w27197 & ~w27213;
assign w29024 = (~w29023 & w28036) | (~w29023 & w49694) | (w28036 & w49694);
assign w29025 = w28038 & ~w29023;
assign w29026 = (~w29024 & w27260) | (~w29024 & w50135) | (w27260 & w50135);
assign w29027 = ~w28076 & w49212;
assign w29028 = (w27196 & w28076) | (w27196 & w42416) | (w28076 & w42416);
assign w29029 = ~w29027 & ~w29028;
assign w29030 = w2285 & ~w28094;
assign w29031 = w29022 & w29023;
assign w29032 = (w2006 & w29027) | (w2006 & w42417) | (w29027 & w42417);
assign w29033 = w29022 & w47799;
assign w29034 = ~w29030 & w29033;
assign w29035 = ~w29032 & ~w29034;
assign w29036 = (w29031 & w28094) | (w29031 & w45719) | (w28094 & w45719);
assign w29037 = w29029 & ~w29036;
assign w29038 = w29029 & w45720;
assign w29039 = (~w29018 & w28052) | (~w29018 & w45721) | (w28052 & w45721);
assign w29040 = w29011 & ~w29019;
assign w29041 = ~w29039 & w29040;
assign w29042 = ~w29016 & ~w29019;
assign w29043 = (~w29042 & w29013) | (~w29042 & w45722) | (w29013 & w45722);
assign w29044 = (w27190 & w28076) | (w27190 & w47800) | (w28076 & w47800);
assign w29045 = w28077 & w42418;
assign w29046 = ~w29044 & ~w29045;
assign w29047 = ~w2285 & w29046;
assign w29048 = (w27139 & w27833) | (w27139 & w47801) | (w27833 & w47801);
assign w29049 = w27125 & w29048;
assign w29050 = ~w27178 & w27893;
assign w29051 = ~w29049 & w29050;
assign w29052 = w28059 & w47802;
assign w29053 = ~w28052 & w29052;
assign w29054 = ~w27159 & ~w27204;
assign w29055 = ~w27202 & ~w29054;
assign w29056 = ~w29053 & w47803;
assign w29057 = (w27158 & w28076) | (w27158 & w42419) | (w28076 & w42419);
assign w29058 = w28077 & w29056;
assign w29059 = ~w29057 & ~w29058;
assign w29060 = w28077 & w42420;
assign w29061 = w29059 & ~w29060;
assign w29062 = (~w2558 & ~w29059) | (~w2558 & w42421) | (~w29059 & w42421);
assign w29063 = w29059 & w42422;
assign w29064 = w27893 & ~w29049;
assign w29065 = w28059 & w47804;
assign w29066 = ~w28052 & w29065;
assign w29067 = ~w29064 & ~w29066;
assign w29068 = ~w27178 & ~w27202;
assign w29069 = ~w27142 & ~w27849;
assign w29070 = w27177 & w27900;
assign w29071 = ~w29069 & w29070;
assign w29072 = w29068 & ~w29071;
assign w29073 = ~w28052 & w47805;
assign w29074 = w29072 & ~w29073;
assign w29075 = w29067 & ~w29074;
assign w29076 = (w29068 & w29066) | (w29068 & w47806) | (w29066 & w47806);
assign w29077 = w28077 & ~w29076;
assign w29078 = ~w3242 & ~w27893;
assign w29079 = ~w28076 & w42423;
assign w29080 = ~w29075 & w29077;
assign w29081 = w27177 & ~w29079;
assign w29082 = ~w29080 & ~w29081;
assign w29083 = (~w2896 & w29080) | (~w2896 & w42424) | (w29080 & w42424);
assign w29084 = ~w29063 & ~w29083;
assign w29085 = ~w29062 & ~w29084;
assign w29086 = (w2285 & w29045) | (w2285 & w47807) | (w29045 & w47807);
assign w29087 = (w29035 & w29038) | (w29035 & w47808) | (w29038 & w47808);
assign w29088 = w29035 & ~w29086;
assign w29089 = w29085 & w29088;
assign w29090 = ~w29087 & ~w29089;
assign w29091 = ~w28076 & w42425;
assign w29092 = w27139 & w27890;
assign w29093 = ~w28036 & w45723;
assign w29094 = w28260 & w29093;
assign w29095 = ~w27906 & w29094;
assign w29096 = ~w29039 & w29092;
assign w29097 = ~w28076 & w45724;
assign w29098 = ~w29095 & w42426;
assign w29099 = ~w29091 & w29098;
assign w29100 = (w29092 & w29095) | (w29092 & w42427) | (w29095 & w42427);
assign w29101 = ~w29097 & ~w29100;
assign w29102 = ~w29099 & w29101;
assign w29103 = (w4056 & ~w29101) | (w4056 & w42428) | (~w29101 & w42428);
assign w29104 = ~w27124 & w27129;
assign w29105 = w27890 & ~w29048;
assign w29106 = w27890 & w29010;
assign w29107 = ~w28052 & w29106;
assign w29108 = (w29104 & w29107) | (w29104 & w45725) | (w29107 & w45725);
assign w29109 = ~w29107 & w45726;
assign w29110 = w28077 & w42429;
assign w29111 = ~w27119 & ~w27122;
assign w29112 = (w29111 & w28076) | (w29111 & w45727) | (w28076 & w45727);
assign w29113 = ~w29110 & ~w29112;
assign w29114 = ~w29110 & w45728;
assign w29115 = ~w29103 & ~w29114;
assign w29116 = (w3646 & w29110) | (w3646 & w45729) | (w29110 & w45729);
assign w29117 = ~w27124 & ~w27891;
assign w29118 = ~w27124 & w29048;
assign w29119 = (w29118 & w28052) | (w29118 & w47809) | (w28052 & w47809);
assign w29120 = ~w29117 & ~w29119;
assign w29121 = w28077 & w29120;
assign w29122 = ~w27105 & ~w27108;
assign w29123 = w3242 & ~w29122;
assign w29124 = (w29123 & w29121) | (w29123 & w42430) | (w29121 & w42430);
assign w29125 = w3242 & w29122;
assign w29126 = ~w29121 & w42431;
assign w29127 = ~w29124 & ~w29126;
assign w29128 = ~w29116 & w29127;
assign w29129 = ~w29115 & w29128;
assign w29130 = ~w29121 & w42432;
assign w29131 = (w29122 & w29121) | (w29122 & w42433) | (w29121 & w42433);
assign w29132 = ~w29130 & ~w29131;
assign w29133 = ~w3242 & ~w29132;
assign w29134 = ~w29080 & w42434;
assign w29135 = ~w29062 & ~w29134;
assign w29136 = ~w29133 & w29135;
assign w29137 = ~w29129 & w29136;
assign w29138 = ~w29038 & ~w29088;
assign w29139 = ~w29129 & w49213;
assign w29140 = w29090 & ~w29139;
assign w29141 = w29008 & w29140;
assign w29142 = (~w29006 & ~w29140) | (~w29006 & w49695) | (~w29140 & w49695);
assign w29143 = w28938 & ~w29142;
assign w29144 = ~w28931 & ~w29143;
assign w29145 = ~w28682 & w29144;
assign w29146 = w29008 & w29090;
assign w29147 = w29101 & w47810;
assign w29148 = w29128 & ~w29147;
assign w29149 = ~w29138 & ~w29148;
assign w29150 = w29137 & w29149;
assign w29151 = w28929 & w29006;
assign w29152 = w28929 & ~w29150;
assign w29153 = w29146 & w29152;
assign w29154 = ~w29151 & ~w29153;
assign w29155 = w42412 & w49214;
assign w29156 = ~w29154 & ~w29155;
assign w29157 = ~w28931 & ~w29156;
assign w29158 = ~w29145 & ~w29157;
assign w29159 = ~w28855 & ~w28935;
assign w29160 = (w28852 & w28855) | (w28852 & w45730) | (w28855 & w45730);
assign w29161 = w28763 & ~w29160;
assign w29162 = w29146 & ~w29150;
assign w29163 = w28681 & w29162;
assign w29164 = ~w28855 & ~w29006;
assign w29165 = ~w29141 & w29164;
assign w29166 = (~w29161 & ~w29165) | (~w29161 & w45731) | (~w29165 & w45731);
assign w29167 = ~w29161 & w29163;
assign w29168 = ~w28663 & w29167;
assign w29169 = ~w29166 & ~w29168;
assign w29170 = ~w28738 & w28743;
assign w29171 = ~w351 & ~w28738;
assign w29172 = ~w29145 & w45732;
assign w29173 = ~w29168 & w45733;
assign w29174 = ~w29158 & w29173;
assign w29175 = ~w29172 & ~w29174;
assign w29176 = ~w29145 & w45734;
assign w29177 = (~w29170 & w29168) | (~w29170 & w45735) | (w29168 & w45735);
assign w29178 = ~w29158 & w29177;
assign w29179 = ~w29176 & ~w29178;
assign w29180 = w29175 & w29179;
assign w29181 = ~w28282 & ~w28287;
assign w29182 = ~w28235 & ~w28283;
assign w29183 = w29181 & w29182;
assign w29184 = w28289 & ~w29183;
assign w29185 = ~w28271 & ~w29184;
assign w29186 = w17380 & ~w29185;
assign w29187 = ~w17380 & w29185;
assign w29188 = ~w29186 & ~w29187;
assign w29189 = (w28250 & w29158) | (w28250 & w50380) | (w29158 & w50380);
assign w29190 = ~w29158 & w50381;
assign w29191 = ~w29189 & ~w29190;
assign w29192 = w16559 & w29191;
assign w29193 = ~w28287 & ~w29183;
assign w29194 = ~w18183 & w29193;
assign w29195 = w18183 & ~w29193;
assign w29196 = ~w29194 & ~w29195;
assign w29197 = (~w29196 & w29145) | (~w29196 & w45736) | (w29145 & w45736);
assign w29198 = w28270 & ~w29197;
assign w29199 = ~w28270 & w29197;
assign w29200 = ~w29198 & ~w29199;
assign w29201 = ~w17380 & ~w29200;
assign w29202 = ~w29192 & ~w29201;
assign w29203 = (w28232 & w29156) | (w28232 & w49215) | (w29156 & w49215);
assign w29204 = ~w29145 & w29203;
assign w29205 = ~w28233 & ~w28283;
assign w29206 = ~w28205 & w45737;
assign w29207 = (w29205 & w28205) | (w29205 & w45738) | (w28205 & w45738);
assign w29208 = ~w29206 & ~w29207;
assign w29209 = ~w29143 & w49216;
assign w29210 = ~w28682 & w29209;
assign w29211 = ~w29156 & w49216;
assign w29212 = ~w29210 & ~w29211;
assign w29213 = ~w29204 & w29212;
assign w29214 = w19040 & ~w29213;
assign w29215 = ~w29181 & ~w29182;
assign w29216 = ~w29183 & ~w29215;
assign w29217 = w18183 & ~w28281;
assign w29218 = ~w29145 & w45739;
assign w29219 = w18183 & ~w29216;
assign w29220 = (w29219 & w29145) | (w29219 & w45740) | (w29145 & w45740);
assign w29221 = ~w29218 & ~w29220;
assign w29222 = ~w29214 & w29221;
assign w29223 = ~w19040 & w29213;
assign w29224 = ~w28188 & ~w28208;
assign w29225 = w28194 & ~w28213;
assign w29226 = ~w28156 & w28159;
assign w29227 = ~w28132 & w28140;
assign w29228 = ~w28105 & w29227;
assign w29229 = ~w29226 & ~w29228;
assign w29230 = w22767 & ~w28190;
assign w29231 = (~w28150 & w29228) | (~w28150 & w45741) | (w29228 & w45741);
assign w29232 = w29230 & ~w29231;
assign w29233 = (~w29225 & w29231) | (~w29225 & w49696) | (w29231 & w49696);
assign w29234 = ~w22767 & ~w28150;
assign w29235 = ~w29228 & w45742;
assign w29236 = w29234 & ~w29235;
assign w29237 = (~w28176 & w29235) | (~w28176 & w49697) | (w29235 & w49697);
assign w29238 = ~w29233 & w29237;
assign w29239 = w28212 & ~w29238;
assign w29240 = w29224 & ~w29239;
assign w29241 = ~w29224 & w29239;
assign w29242 = ~w29240 & ~w29241;
assign w29243 = ~w20000 & ~w28207;
assign w29244 = ~w29145 & w45743;
assign w29245 = ~w20000 & w29242;
assign w29246 = (w29245 & w29145) | (w29245 & w49217) | (w29145 & w49217);
assign w29247 = ~w29244 & ~w29246;
assign w29248 = ~w29223 & w29247;
assign w29249 = w29222 & ~w29248;
assign w29250 = w17380 & ~w28270;
assign w29251 = ~w29197 & w29250;
assign w29252 = w17380 & w28270;
assign w29253 = w29197 & w29252;
assign w29254 = ~w29251 & ~w29253;
assign w29255 = ~w29145 & w45744;
assign w29256 = ~w18183 & ~w29255;
assign w29257 = ~w29158 & ~w29216;
assign w29258 = w29256 & ~w29257;
assign w29259 = w29254 & ~w29258;
assign w29260 = ~w29249 & w29259;
assign w29261 = ~w29145 & w50382;
assign w29262 = (w29242 & w29145) | (w29242 & w50383) | (w29145 & w50383);
assign w29263 = ~w29261 & ~w29262;
assign w29264 = w20000 & w29263;
assign w29265 = w29222 & ~w29264;
assign w29266 = (w29202 & ~w29260) | (w29202 & w50384) | (~w29260 & w50384);
assign w29267 = (w28504 & w28290) | (w28504 & w49698) | (w28290 & w49698);
assign w29268 = ~w28286 & w29267;
assign w29269 = ~w28482 & ~w29268;
assign w29270 = ~w13384 & w29269;
assign w29271 = w13384 & ~w29269;
assign w29272 = ~w29270 & ~w29271;
assign w29273 = (w29272 & w29145) | (w29272 & w45745) | (w29145 & w45745);
assign w29274 = w28403 & ~w29273;
assign w29275 = ~w28403 & w29273;
assign w29276 = ~w29274 & ~w29275;
assign w29277 = w12666 & ~w29276;
assign w29278 = ~w28358 & ~w28388;
assign w29279 = ~w28404 & ~w29269;
assign w29280 = ~w28425 & ~w29279;
assign w29281 = ~w29145 & w45746;
assign w29282 = (w29280 & w29145) | (w29280 & w45747) | (w29145 & w45747);
assign w29283 = ~w29281 & ~w29282;
assign w29284 = w29278 & w29283;
assign w29285 = ~w29278 & ~w29283;
assign w29286 = ~w29284 & ~w29285;
assign w29287 = ~w11870 & w29286;
assign w29288 = ~w28424 & ~w28440;
assign w29289 = ~w28439 & ~w28477;
assign w29290 = ~w28476 & w29289;
assign w29291 = w28502 & w50217;
assign w29292 = w29290 & ~w29291;
assign w29293 = w28439 & ~w29288;
assign w29294 = ~w28439 & w29288;
assign w29295 = ~w29293 & ~w29294;
assign w29296 = w29288 & w29292;
assign w29297 = ~w29292 & w29295;
assign w29298 = ~w29296 & ~w29297;
assign w29299 = w28423 & w29158;
assign w29300 = ~w29158 & w29298;
assign w29301 = ~w29299 & ~w29300;
assign w29302 = ~w13384 & ~w29301;
assign w29303 = w13384 & w29295;
assign w29304 = ~w29292 & w29303;
assign w29305 = w13384 & w29288;
assign w29306 = w29292 & w29305;
assign w29307 = ~w29304 & ~w29306;
assign w29308 = ~w29158 & ~w29307;
assign w29309 = w13384 & ~w28423;
assign w29310 = ~w29145 & w45749;
assign w29311 = ~w29308 & ~w29310;
assign w29312 = w28502 & ~w29289;
assign w29313 = w29312 & w50217;
assign w29314 = w28476 & ~w29289;
assign w29315 = ~w29313 & ~w29314;
assign w29316 = ~w29292 & w29315;
assign w29317 = ~w14039 & ~w28438;
assign w29318 = ~w29145 & w45750;
assign w29319 = ~w14039 & ~w29316;
assign w29320 = ~w29158 & w29319;
assign w29321 = ~w29318 & ~w29320;
assign w29322 = w29311 & w29321;
assign w29323 = w14039 & w28438;
assign w29324 = ~w14766 & ~w28458;
assign w29325 = ~w29323 & ~w29324;
assign w29326 = ~w28459 & ~w28476;
assign w29327 = ~w28501 & w50217;
assign w29328 = w29326 & ~w29327;
assign w29329 = ~w29326 & w29327;
assign w29330 = ~w29328 & ~w29329;
assign w29331 = w14039 & w29316;
assign w29332 = ~w14766 & w29330;
assign w29333 = ~w29331 & ~w29332;
assign w29334 = w29158 & w29325;
assign w29335 = ~w29158 & w29333;
assign w29336 = ~w29334 & ~w29335;
assign w29337 = w29322 & w29336;
assign w29338 = ~w29302 & ~w29337;
assign w29339 = ~w16559 & w28250;
assign w29340 = (w29339 & w29158) | (w29339 & w45751) | (w29158 & w45751);
assign w29341 = ~w16559 & ~w28250;
assign w29342 = ~w29158 & w45752;
assign w29343 = ~w29340 & ~w29342;
assign w29344 = ~w28273 & w45753;
assign w29345 = ~w28235 & w29344;
assign w29346 = (~w16559 & w28290) | (~w16559 & w49699) | (w28290 & w49699);
assign w29347 = ~w28286 & w29346;
assign w29348 = ~w28290 & w49700;
assign w29349 = ~w29345 & ~w29348;
assign w29350 = ~w29347 & w29349;
assign w29351 = ~w28931 & ~w29350;
assign w29352 = ~w29143 & w29351;
assign w29353 = ~w28682 & w29352;
assign w29354 = w29157 & ~w29350;
assign w29355 = ~w15681 & w52271;
assign w29356 = ~w29353 & w47811;
assign w29357 = w29355 & ~w29356;
assign w29358 = w29343 & ~w29357;
assign w29359 = w11870 & w29278;
assign w29360 = w29283 & w29359;
assign w29361 = w11870 & ~w29278;
assign w29362 = ~w29283 & w29361;
assign w29363 = ~w29360 & ~w29362;
assign w29364 = w29358 & w29363;
assign w29365 = w29338 & w29364;
assign w29366 = w29277 & ~w29287;
assign w29367 = w29365 & ~w29366;
assign w29368 = ~w29266 & w29367;
assign w29369 = ~w28663 & w29163;
assign w29370 = w28920 & ~w28936;
assign w29371 = w28920 & w29142;
assign w29372 = (~w29370 & w29369) | (~w29370 & w47812) | (w29369 & w47812);
assign w29373 = ~w28122 & ~w28123;
assign w29374 = w28094 & w28120;
assign w29375 = ~a[21] & ~w29374;
assign w29376 = ~w27271 & w28094;
assign w29377 = ~w29375 & ~w29376;
assign w29378 = ~w29373 & ~w29377;
assign w29379 = a[21] & w28077;
assign w29380 = ~a[20] & ~w28930;
assign w29381 = w29379 & ~w29380;
assign w29382 = w29373 & ~w29381;
assign w29383 = ~a[21] & ~w28077;
assign w29384 = ~w29378 & ~w29382;
assign w29385 = ~w29378 & w29383;
assign w29386 = (w29385 & w29145) | (w29385 & w45754) | (w29145 & w45754);
assign w29387 = ~w29384 & ~w29386;
assign w29388 = ~w29378 & w29379;
assign w29389 = ~w29372 & w29388;
assign w29390 = w29387 & ~w29389;
assign w29391 = ~a[20] & w28077;
assign w29392 = a[21] & ~w29391;
assign w29393 = ~a[21] & w29391;
assign w29394 = ~w29392 & ~w29393;
assign w29395 = ~a[21] & w28123;
assign w29396 = w28094 & w29395;
assign w29397 = ~w29145 & w45755;
assign w29398 = (w29396 & w29145) | (w29396 & w45756) | (w29145 & w45756);
assign w29399 = ~w29397 & ~w29398;
assign w29400 = w29390 & w29399;
assign w29401 = ~w25851 & ~w29400;
assign w29402 = (w29142 & w28663) | (w29142 & w45757) | (w28663 & w45757);
assign w29403 = a[18] & ~a[19];
assign w29404 = ~w28931 & w29403;
assign w29405 = ~a[16] & ~a[17];
assign w29406 = ~a[18] & w29405;
assign w29407 = w28077 & w29406;
assign w29408 = ~w29404 & ~w29407;
assign w29409 = w29156 & ~w29407;
assign w29410 = ~w29402 & w29409;
assign w29411 = ~w29408 & ~w29410;
assign w29412 = ~w28077 & ~w29406;
assign w29413 = ~a[19] & ~w29412;
assign w29414 = ~w29157 & w29413;
assign w29415 = ~w29145 & w29414;
assign w29416 = a[19] & ~w29412;
assign w29417 = (w29416 & w28920) | (w29416 & w42437) | (w28920 & w42437);
assign w29418 = ~w29143 & w29417;
assign w29419 = ~w28682 & w29418;
assign w29420 = w29157 & w29416;
assign w29421 = ~w29419 & ~w29420;
assign w29422 = ~w29415 & w29421;
assign w29423 = ~w29411 & w29422;
assign w29424 = ~w26880 & ~w29423;
assign w29425 = w29422 & w45758;
assign w29426 = ~w28663 & w45759;
assign w29427 = w28937 & ~w29426;
assign w29428 = a[20] & ~w28120;
assign w29429 = ~w28121 & ~w29428;
assign w29430 = ~w28931 & w29429;
assign w29431 = w29156 & ~w29402;
assign w29432 = ~w29427 & w29431;
assign w29433 = w29430 & ~w29432;
assign w29434 = a[20] & ~w28077;
assign w29435 = ~w29391 & ~w29434;
assign w29436 = w29158 & w29435;
assign w29437 = ~w29433 & ~w29436;
assign w29438 = ~w29425 & ~w29437;
assign w29439 = ~w29424 & ~w29438;
assign w29440 = ~w29401 & ~w29439;
assign w29441 = ~w29232 & ~w29236;
assign w29442 = (w29441 & w29145) | (w29441 & w45760) | (w29145 & w45760);
assign w29443 = ~w21801 & w29225;
assign w29444 = ~w29442 & w29443;
assign w29445 = ~w21801 & ~w29225;
assign w29446 = w29442 & w29445;
assign w29447 = w28149 & ~w29143;
assign w29448 = w23843 & ~w29229;
assign w29449 = ~w23843 & w29229;
assign w29450 = ~w29448 & ~w29449;
assign w29451 = (~w29450 & w29145) | (~w29450 & w45761) | (w29145 & w45761);
assign w29452 = w22767 & ~w28149;
assign w29453 = ~w29451 & w29452;
assign w29454 = w22767 & w29447;
assign w29455 = w29451 & w29454;
assign w29456 = ~w29453 & ~w29455;
assign w29457 = ~w29444 & ~w29446;
assign w29458 = w29456 & w29457;
assign w29459 = ~w29226 & w29227;
assign w29460 = (w29459 & w29145) | (w29459 & w45762) | (w29145 & w45762);
assign w29461 = w23843 & w28105;
assign w29462 = ~w29460 & w29461;
assign w29463 = w23843 & ~w28105;
assign w29464 = w29460 & w29463;
assign w29465 = ~w29462 & ~w29464;
assign w29466 = ~w22767 & ~w29447;
assign w29467 = w29451 & w29466;
assign w29468 = ~w22767 & w28149;
assign w29469 = ~w29451 & w29468;
assign w29470 = ~w29467 & ~w29469;
assign w29471 = ~w29465 & w29470;
assign w29472 = w29458 & ~w29471;
assign w29473 = w25851 & w29399;
assign w29474 = w29390 & w29473;
assign w29475 = ~w28069 & w28114;
assign w29476 = ~w28109 & ~w29475;
assign w29477 = ~w28135 & ~w28157;
assign w29478 = ~w28155 & w29477;
assign w29479 = ~w28131 & ~w29478;
assign w29480 = w28156 & w29477;
assign w29481 = ~w29479 & ~w29480;
assign w29482 = w29158 & ~w29476;
assign w29483 = ~w29158 & w29481;
assign w29484 = ~w29482 & ~w29483;
assign w29485 = w24874 & ~w29484;
assign w29486 = ~w29474 & ~w29485;
assign w29487 = w29472 & w29486;
assign w29488 = ~w29440 & w29487;
assign w29489 = ~w24874 & w29484;
assign w29490 = ~w23843 & ~w28105;
assign w29491 = ~w29460 & w29490;
assign w29492 = ~w23843 & w28105;
assign w29493 = w29460 & w29492;
assign w29494 = ~w29491 & ~w29493;
assign w29495 = w29470 & w29494;
assign w29496 = w29458 & ~w29495;
assign w29497 = w29225 & ~w29442;
assign w29498 = ~w29225 & w29442;
assign w29499 = ~w29497 & ~w29498;
assign w29500 = w21801 & w29499;
assign w29501 = ~w28161 & ~w28174;
assign w29502 = ~w29233 & ~w29236;
assign w29503 = ~w21801 & w29502;
assign w29504 = w21801 & ~w29502;
assign w29505 = ~w29503 & ~w29504;
assign w29506 = (w29505 & w29145) | (w29505 & w45763) | (w29145 & w45763);
assign w29507 = w29501 & ~w29506;
assign w29508 = ~w29501 & w29506;
assign w29509 = ~w29507 & ~w29508;
assign w29510 = ~w20906 & ~w29509;
assign w29511 = ~w29500 & ~w29510;
assign w29512 = ~w29496 & w29511;
assign w29513 = w29472 & w29489;
assign w29514 = w29512 & ~w29513;
assign w29515 = ~w29488 & w29514;
assign w29516 = w20906 & w29509;
assign w29517 = w29260 & ~w29516;
assign w29518 = w29367 & w29517;
assign w29519 = ~w29515 & w29518;
assign w29520 = ~w29368 & ~w29519;
assign w29521 = ~w28630 & w28650;
assign w29522 = w8666 & ~w28645;
assign w29523 = ~w28375 & ~w28376;
assign w29524 = w28385 & ~w28497;
assign w29525 = w28483 & ~w29524;
assign w29526 = w29523 & w29525;
assign w29527 = ~w29268 & w29526;
assign w29528 = ~w28676 & ~w29522;
assign w29529 = ~w28499 & w45764;
assign w29530 = (~w29528 & w29527) | (~w29528 & w45765) | (w29527 & w45765);
assign w29531 = w29521 & ~w29530;
assign w29532 = ~w29521 & w29530;
assign w29533 = ~w29531 & ~w29532;
assign w29534 = ~w29145 & w45766;
assign w29535 = ~w29158 & w29533;
assign w29536 = ~w29534 & ~w29535;
assign w29537 = w7315 & w29536;
assign w29538 = w28653 & w50218;
assign w29539 = ~w28623 & ~w28655;
assign w29540 = ~w29538 & w29539;
assign w29541 = w29538 & ~w29539;
assign w29542 = w28622 & w29158;
assign w29543 = ~w29158 & w45768;
assign w29544 = ~w29542 & ~w29543;
assign w29545 = ~w6769 & ~w29544;
assign w29546 = ~w29537 & ~w29545;
assign w29547 = ~w28670 & ~w29522;
assign w29548 = (w28675 & w29527) | (w28675 & w45769) | (w29527 & w45769);
assign w29549 = w29547 & ~w29548;
assign w29550 = ~w29547 & w29548;
assign w29551 = ~w29549 & ~w29550;
assign w29552 = ~w29145 & w45770;
assign w29553 = ~w29158 & ~w29551;
assign w29554 = (w7924 & w29553) | (w7924 & w45771) | (w29553 & w45771);
assign w29555 = w28407 & w29268;
assign w29556 = w28485 & ~w29555;
assign w29557 = ~w28487 & ~w29556;
assign w29558 = (~w29557 & w29145) | (~w29557 & w45772) | (w29145 & w45772);
assign w29559 = (~w9195 & w29156) | (~w9195 & w49218) | (w29156 & w49218);
assign w29560 = ~w28497 & w28675;
assign w29561 = w8666 & w29560;
assign w29562 = (w29561 & w29145) | (w29561 & w49219) | (w29145 & w49219);
assign w29563 = ~w29558 & w29562;
assign w29564 = w8666 & ~w29560;
assign w29565 = ~w29145 & w49220;
assign w29566 = ~w29557 & w29564;
assign w29567 = ~w29158 & w29566;
assign w29568 = ~w29565 & ~w29567;
assign w29569 = ~w29563 & w29568;
assign w29570 = ~w29554 & w29569;
assign w29571 = ~w8666 & ~w29560;
assign w29572 = (w29571 & w29145) | (w29571 & w49221) | (w29145 & w49221);
assign w29573 = ~w29558 & w29572;
assign w29574 = ~w8666 & w29560;
assign w29575 = ~w29145 & w49222;
assign w29576 = ~w29557 & w29574;
assign w29577 = ~w29158 & w29576;
assign w29578 = ~w29575 & ~w29577;
assign w29579 = ~w29573 & w29578;
assign w29580 = ~w28385 & ~w28487;
assign w29581 = ~w28484 & w29523;
assign w29582 = ~w29555 & w29581;
assign w29583 = w29580 & ~w29582;
assign w29584 = ~w29580 & w29582;
assign w29585 = ~w29583 & ~w29584;
assign w29586 = ~w29145 & w45773;
assign w29587 = ~w29158 & ~w29585;
assign w29588 = ~w29587 & w45774;
assign w29589 = w29579 & ~w29588;
assign w29590 = w29570 & ~w29589;
assign w29591 = (~w7315 & w29535) | (~w7315 & w45775) | (w29535 & w45775);
assign w29592 = ~w29553 & w45776;
assign w29593 = ~w29591 & ~w29592;
assign w29594 = ~w29590 & w29593;
assign w29595 = ~w28358 & w28483;
assign w29596 = ~w29268 & w29595;
assign w29597 = ~w28358 & ~w28405;
assign w29598 = ~w28329 & ~w29597;
assign w29599 = (w29598 & w29268) | (w29598 & w45777) | (w29268 & w45777);
assign w29600 = ~w29599 & w47813;
assign w29601 = (w11138 & w29599) | (w11138 & w47814) | (w29599 & w47814);
assign w29602 = ~w29600 & ~w29601;
assign w29603 = (w28326 & w29158) | (w28326 & w45778) | (w29158 & w45778);
assign w29604 = ~w29158 & w45779;
assign w29605 = ~w29603 & ~w29604;
assign w29606 = w10419 & ~w29605;
assign w29607 = ~w29145 & w45780;
assign w29608 = ~w29596 & ~w29597;
assign w29609 = (w29608 & w29145) | (w29608 & w45781) | (w29145 & w45781);
assign w29610 = ~w29607 & ~w29609;
assign w29611 = ~w28311 & ~w28329;
assign w29612 = ~w11138 & w29611;
assign w29613 = ~w29610 & w29612;
assign w29614 = ~w11138 & ~w29611;
assign w29615 = w29610 & w29614;
assign w29616 = ~w29613 & ~w29615;
assign w29617 = ~w29606 & w29616;
assign w29618 = ~w10419 & w29605;
assign w29619 = ~w28373 & ~w28376;
assign w29620 = (~w28361 & w29599) | (~w28361 & w47815) | (w29599 & w47815);
assign w29621 = w29619 & ~w29620;
assign w29622 = ~w29619 & w29620;
assign w29623 = ~w29621 & ~w29622;
assign w29624 = ~w29145 & w47816;
assign w29625 = ~w29158 & ~w29623;
assign w29626 = ~w29624 & ~w29625;
assign w29627 = (~w9781 & w29625) | (~w9781 & w47817) | (w29625 & w47817);
assign w29628 = ~w29618 & ~w29627;
assign w29629 = ~w29617 & w29628;
assign w29630 = ~w29625 & w47818;
assign w29631 = (~w9195 & w29587) | (~w9195 & w47819) | (w29587 & w47819);
assign w29632 = w29570 & w45782;
assign w29633 = ~w29629 & w29632;
assign w29634 = w29594 & ~w29633;
assign w29635 = w29546 & ~w29634;
assign w29636 = (w29635 & w29519) | (w29635 & w45783) | (w29519 & w45783);
assign w29637 = w29546 & w29633;
assign w29638 = w6769 & w29544;
assign w29639 = ~w29546 & ~w29638;
assign w29640 = w29593 & ~w29638;
assign w29641 = ~w29590 & w29640;
assign w29642 = ~w29639 & ~w29641;
assign w29643 = w15681 & w28472;
assign w29644 = (w29643 & w29353) | (w29643 & w42438) | (w29353 & w42438);
assign w29645 = w15681 & ~w28472;
assign w29646 = ~w29353 & w42439;
assign w29647 = ~w29644 & ~w29646;
assign w29648 = w14766 & w28458;
assign w29649 = ~w29145 & w45784;
assign w29650 = w14766 & ~w29330;
assign w29651 = ~w29158 & w29650;
assign w29652 = ~w29649 & ~w29651;
assign w29653 = w29647 & w29652;
assign w29654 = w29322 & w29653;
assign w29655 = ~w29277 & ~w29654;
assign w29656 = w29338 & w29655;
assign w29657 = ~w12666 & w29276;
assign w29658 = (w29363 & w29656) | (w29363 & w45785) | (w29656 & w45785);
assign w29659 = w29610 & ~w29611;
assign w29660 = ~w29610 & w29611;
assign w29661 = ~w29659 & ~w29660;
assign w29662 = w11138 & w29661;
assign w29663 = ~w29606 & w29662;
assign w29664 = w29628 & ~w29663;
assign w29665 = ~w29637 & ~w29642;
assign w29666 = ~w29642 & w29664;
assign w29667 = ~w29658 & w29666;
assign w29668 = ~w29665 & ~w29667;
assign w29669 = ~w29145 & w47820;
assign w29670 = ~w29158 & w45786;
assign w29671 = ~w28580 & ~w28656;
assign w29672 = ~w29670 & w47821;
assign w29673 = (w29671 & w29670) | (w29671 & w47822) | (w29670 & w47822);
assign w29674 = ~w29672 & ~w29673;
assign w29675 = ~w6264 & w29674;
assign w29676 = (~w29675 & w29667) | (~w29675 & w45787) | (w29667 & w45787);
assign w29677 = ~w29636 & w29676;
assign w29678 = (w4430 & w29156) | (w4430 & w49223) | (w29156 & w49223);
assign w29679 = ~w29145 & w29678;
assign w29680 = (w28556 & ~w28606) | (w28556 & w45788) | (~w28606 & w45788);
assign w29681 = ~w28667 & w28679;
assign w29682 = w29680 & ~w29681;
assign w29683 = ~w28654 & w28657;
assign w29684 = w29680 & ~w29683;
assign w29685 = w28500 & w29684;
assign w29686 = ~w29527 & w29685;
assign w29687 = ~w29682 & ~w29686;
assign w29688 = (~w28546 & w29686) | (~w28546 & w45789) | (w29686 & w45789);
assign w29689 = w28532 & ~w29688;
assign w29690 = ~w29158 & w29689;
assign w29691 = ~w29679 & ~w29690;
assign w29692 = w28524 & w28542;
assign w29693 = w4056 & ~w29692;
assign w29694 = (w29693 & w29690) | (w29693 & w45790) | (w29690 & w45790);
assign w29695 = w4056 & w29692;
assign w29696 = ~w29690 & w45791;
assign w29697 = ~w29694 & ~w29696;
assign w29698 = w4056 & w29145;
assign w29699 = w28682 & w29157;
assign w29700 = ~w4056 & w29699;
assign w29701 = ~w29698 & ~w29700;
assign w29702 = ~w3646 & w29102;
assign w29703 = ~w29701 & w29702;
assign w29704 = ~w3646 & ~w29102;
assign w29705 = w29701 & w29704;
assign w29706 = ~w29703 & ~w29705;
assign w29707 = w28532 & ~w28546;
assign w29708 = ~w29686 & w45792;
assign w29709 = w4430 & ~w29708;
assign w29710 = ~w29687 & ~w29707;
assign w29711 = w29709 & ~w29710;
assign w29712 = ~w28545 & w29679;
assign w29713 = ~w29158 & w29711;
assign w29714 = ~w29712 & ~w29713;
assign w29715 = w29706 & w29714;
assign w29716 = w29697 & w29715;
assign w29717 = w6264 & ~w29674;
assign w29718 = ~w28506 & w28654;
assign w29719 = w28500 & w29718;
assign w29720 = ~w28486 & w29719;
assign w29721 = w28657 & ~w28678;
assign w29722 = ~w28580 & w29721;
assign w29723 = ~w29720 & w29722;
assign w29724 = ~w28580 & ~w28597;
assign w29725 = w28580 & w28597;
assign w29726 = ~w29724 & ~w29725;
assign w29727 = w29721 & w29724;
assign w29728 = ~w29720 & w29727;
assign w29729 = ~w29723 & w29726;
assign w29730 = ~w29728 & ~w29729;
assign w29731 = w28590 & ~w28591;
assign w29732 = ~w28590 & w28591;
assign w29733 = ~w29731 & ~w29732;
assign w29734 = ~w29158 & w29730;
assign w29735 = w29158 & w29733;
assign w29736 = ~w29734 & ~w29735;
assign w29737 = ~w5745 & ~w29736;
assign w29738 = w28602 & ~w29724;
assign w29739 = ~w28588 & ~w28598;
assign w29740 = w29738 & ~w29739;
assign w29741 = ~w29738 & w29739;
assign w29742 = ~w29740 & ~w29741;
assign w29743 = ~w29720 & w45793;
assign w29744 = (w29742 & w29720) | (w29742 & w45794) | (w29720 & w45794);
assign w29745 = ~w29743 & ~w29744;
assign w29746 = ~w29145 & w45795;
assign w29747 = ~w29158 & ~w29745;
assign w29748 = ~w29746 & ~w29747;
assign w29749 = w5330 & w29748;
assign w29750 = ~w29737 & ~w29749;
assign w29751 = w28556 & ~w28667;
assign w29752 = ~w29527 & w45796;
assign w29753 = w28679 & ~w29752;
assign w29754 = ~w28606 & ~w29753;
assign w29755 = w29751 & ~w29754;
assign w29756 = ~w29751 & w29754;
assign w29757 = ~w29755 & ~w29756;
assign w29758 = ~w28666 & w29158;
assign w29759 = ~w29158 & ~w29757;
assign w29760 = ~w29758 & ~w29759;
assign w29761 = ~w4838 & w29760;
assign w29762 = w29750 & ~w29761;
assign w29763 = ~w29717 & w29762;
assign w29764 = w29716 & w29763;
assign w29765 = ~w29083 & ~w29134;
assign w29766 = ~w29129 & ~w29133;
assign w29767 = w29765 & w29766;
assign w29768 = ~w29083 & ~w29767;
assign w29769 = ~w29062 & ~w29063;
assign w29770 = w29768 & ~w29769;
assign w29771 = ~w29768 & w29769;
assign w29772 = ~w29770 & ~w29771;
assign w29773 = (w29148 & w28560) | (w29148 & w45797) | (w28560 & w45797);
assign w29774 = ~w28680 & w45798;
assign w29775 = ~w28680 & w47823;
assign w29776 = ~w28663 & w29775;
assign w29777 = (w29772 & w28663) | (w29772 & w45799) | (w28663 & w45799);
assign w29778 = ~w28663 & w45800;
assign w29779 = ~w29777 & ~w29778;
assign w29780 = ~w29158 & ~w29779;
assign w29781 = (w29061 & w29156) | (w29061 & w49224) | (w29156 & w49224);
assign w29782 = ~w29145 & w29781;
assign w29783 = (w2285 & w29145) | (w2285 & w49225) | (w29145 & w49225);
assign w29784 = ~w29780 & w29783;
assign w29785 = ~w29765 & ~w29766;
assign w29786 = ~w29767 & ~w29785;
assign w29787 = (w29786 & w28663) | (w29786 & w45801) | (w28663 & w45801);
assign w29788 = (~w2558 & w28663) | (~w2558 & w47824) | (w28663 & w47824);
assign w29789 = ~w29787 & w29788;
assign w29790 = ~w2558 & w29082;
assign w29791 = ~w29145 & w45802;
assign w29792 = ~w29158 & w29789;
assign w29793 = ~w29791 & ~w29792;
assign w29794 = ~w29784 & w29793;
assign w29795 = ~w29780 & ~w29782;
assign w29796 = ~w2285 & ~w29795;
assign w29797 = ~w29794 & ~w29796;
assign w29798 = ~w29114 & ~w29116;
assign w29799 = (~w29103 & w28663) | (~w29103 & w45803) | (w28663 & w45803);
assign w29800 = ~w29147 & ~w29799;
assign w29801 = ~w29798 & ~w29800;
assign w29802 = ~w29147 & w29798;
assign w29803 = ~w29799 & w29802;
assign w29804 = ~w29158 & ~w29803;
assign w29805 = ~w29801 & w29804;
assign w29806 = w29113 & w29158;
assign w29807 = ~w29805 & ~w29806;
assign w29808 = (~w3242 & w29805) | (~w3242 & w45804) | (w29805 & w45804);
assign w29809 = ~w29116 & ~w29147;
assign w29810 = w28681 & w29809;
assign w29811 = ~w29115 & ~w29116;
assign w29812 = (~w29811 & w28663) | (~w29811 & w45805) | (w28663 & w45805);
assign w29813 = w29127 & ~w29133;
assign w29814 = w29812 & ~w29813;
assign w29815 = ~w29812 & w29813;
assign w29816 = ~w29814 & ~w29815;
assign w29817 = ~w29145 & w45806;
assign w29818 = w2896 & ~w29817;
assign w29819 = ~w29158 & ~w29816;
assign w29820 = w29818 & ~w29819;
assign w29821 = ~w29808 & ~w29820;
assign w29822 = ~w29797 & w29821;
assign w29823 = w29764 & w29822;
assign w29824 = ~w28968 & ~w28969;
assign w29825 = ~w28680 & w45807;
assign w29826 = ~w28982 & ~w28999;
assign w29827 = ~w29140 & w29826;
assign w29828 = (w29827 & w28663) | (w29827 & w45808) | (w28663 & w45808);
assign w29829 = ~w29145 & w45809;
assign w29830 = ~w28982 & ~w29828;
assign w29831 = ~w29158 & w29830;
assign w29832 = (w29824 & w29831) | (w29824 & w45810) | (w29831 & w45810);
assign w29833 = ~w29831 & w45811;
assign w29834 = ~w29832 & ~w29833;
assign w29835 = w1320 & w29834;
assign w29836 = ~w28998 & ~w29003;
assign w29837 = w29000 & ~w29140;
assign w29838 = (w29837 & w28663) | (w29837 & w45812) | (w28663 & w45812);
assign w29839 = ~w28984 & ~w29838;
assign w29840 = ~w29145 & w45813;
assign w29841 = ~w29158 & w29839;
assign w29842 = ~w29840 & ~w29841;
assign w29843 = (w29836 & w29841) | (w29836 & w45814) | (w29841 & w45814);
assign w29844 = ~w1120 & ~w29843;
assign w29845 = ~w29836 & w29842;
assign w29846 = w29844 & ~w29845;
assign w29847 = ~w29835 & ~w29846;
assign w29848 = ~w28680 & w47825;
assign w29849 = w29140 & ~w29826;
assign w29850 = ~w29827 & ~w29849;
assign w29851 = ~w28663 & w45815;
assign w29852 = (w29850 & w28663) | (w29850 & w45816) | (w28663 & w45816);
assign w29853 = ~w29851 & ~w29852;
assign w29854 = ~w29145 & w45817;
assign w29855 = ~w29158 & ~w29853;
assign w29856 = ~w29854 & ~w29855;
assign w29857 = ~w1541 & ~w29856;
assign w29858 = ~w1320 & w29824;
assign w29859 = (w29858 & w29831) | (w29858 & w45818) | (w29831 & w45818);
assign w29860 = ~w1320 & ~w29824;
assign w29861 = ~w29831 & w45819;
assign w29862 = ~w29859 & ~w29861;
assign w29863 = ~w29857 & w29862;
assign w29864 = (~w29037 & w29156) | (~w29037 & w49226) | (w29156 & w49226);
assign w29865 = ~w29145 & w29864;
assign w29866 = ~w28680 & w45820;
assign w29867 = ~w29085 & ~w29137;
assign w29868 = ~w29086 & ~w29867;
assign w29869 = ~w29047 & w29868;
assign w29870 = w29866 & w29869;
assign w29871 = ~w28663 & w29870;
assign w29872 = w29035 & ~w29038;
assign w29873 = ~w29047 & ~w29868;
assign w29874 = w29872 & ~w29873;
assign w29875 = ~w29872 & w29873;
assign w29876 = ~w29874 & ~w29875;
assign w29877 = w29871 & ~w29876;
assign w29878 = ~w29871 & w29876;
assign w29879 = ~w29877 & ~w29878;
assign w29880 = ~w29158 & w29879;
assign w29881 = (w1738 & w29880) | (w1738 & w45821) | (w29880 & w45821);
assign w29882 = ~w29855 & w47826;
assign w29883 = ~w29881 & ~w29882;
assign w29884 = ~w28680 & w47827;
assign w29885 = w2285 & ~w29867;
assign w29886 = ~w2285 & w29867;
assign w29887 = ~w29885 & ~w29886;
assign w29888 = ~w28663 & w45822;
assign w29889 = (w29887 & w28663) | (w29887 & w45823) | (w28663 & w45823);
assign w29890 = ~w29888 & ~w29889;
assign w29891 = ~w29158 & w29890;
assign w29892 = (w29046 & w29158) | (w29046 & w45824) | (w29158 & w45824);
assign w29893 = ~w29158 & w45825;
assign w29894 = ~w29892 & ~w29893;
assign w29895 = (~w1738 & w29145) | (~w1738 & w49227) | (w29145 & w49227);
assign w29896 = ~w29880 & w29895;
assign w29897 = (w2006 & w29880) | (w2006 & w49228) | (w29880 & w49228);
assign w29898 = w29894 & w29897;
assign w29899 = w29883 & ~w29898;
assign w29900 = w29863 & ~w29899;
assign w29901 = w29847 & ~w29900;
assign w29902 = ~w29145 & w45826;
assign w29903 = ~w29141 & w45827;
assign w29904 = ~w28933 & ~w29903;
assign w29905 = ~w28933 & w29163;
assign w29906 = ~w28663 & w29905;
assign w29907 = ~w29904 & ~w29906;
assign w29908 = ~w28781 & ~w28797;
assign w29909 = ~w29906 & w45828;
assign w29910 = ~w29158 & ~w29909;
assign w29911 = ~w29907 & w29908;
assign w29912 = w29910 & ~w29911;
assign w29913 = (~w29902 & ~w29910) | (~w29902 & w45829) | (~w29910 & w45829);
assign w29914 = w612 & ~w29913;
assign w29915 = (~w945 & w28920) | (~w945 & w45830) | (w28920 & w45830);
assign w29916 = w28932 & ~w29915;
assign w29917 = ~w28932 & w29915;
assign w29918 = ~w29916 & ~w29917;
assign w29919 = ~w28931 & w42440;
assign w29920 = w28932 & w29919;
assign w29921 = ~w28932 & ~w29919;
assign w29922 = w29402 & ~w29918;
assign w29923 = ~w29402 & ~w29920;
assign w29924 = ~w29921 & w29923;
assign w29925 = ~w29922 & ~w29924;
assign w29926 = ~w29924 & w45831;
assign w29927 = ~w612 & ~w29902;
assign w29928 = ~w29912 & w29927;
assign w29929 = ~w29926 & ~w29928;
assign w29930 = ~w29914 & ~w29929;
assign w29931 = ~w29002 & ~w29003;
assign w29932 = ~w29140 & w29931;
assign w29933 = (w29932 & w28663) | (w29932 & w45832) | (w28663 & w45832);
assign w29934 = ~w29003 & ~w29007;
assign w29935 = ~w29933 & ~w29934;
assign w29936 = ~w29145 & w45833;
assign w29937 = ~w29158 & w29935;
assign w29938 = ~w28951 & ~w29004;
assign w29939 = w945 & ~w29938;
assign w29940 = ~w29937 & w45834;
assign w29941 = w945 & w29938;
assign w29942 = (w29941 & w29937) | (w29941 & w45835) | (w29937 & w45835);
assign w29943 = ~w29940 & ~w29942;
assign w29944 = w29836 & w29839;
assign w29945 = ~w29158 & ~w29944;
assign w29946 = ~w29836 & ~w29839;
assign w29947 = w29945 & ~w29946;
assign w29948 = ~w28997 & w29158;
assign w29949 = w1120 & ~w29948;
assign w29950 = ~w29947 & w29949;
assign w29951 = w29943 & ~w29950;
assign w29952 = ~w29930 & w29951;
assign w29953 = ~w29937 & w45836;
assign w29954 = (w29938 & w29937) | (w29938 & w45837) | (w29937 & w45837);
assign w29955 = ~w29953 & ~w29954;
assign w29956 = ~w945 & w29955;
assign w29957 = w754 & ~w29925;
assign w29958 = ~w29956 & ~w29957;
assign w29959 = ~w29914 & w29958;
assign w29960 = ~w29930 & ~w29959;
assign w29961 = ~w29901 & w29952;
assign w29962 = ~w29960 & ~w29961;
assign w29963 = w29823 & w29962;
assign w29964 = ~w28819 & w28841;
assign w29965 = w28934 & w29964;
assign w29966 = ~w28799 & ~w29964;
assign w29967 = w29142 & w29966;
assign w29968 = w28799 & w29964;
assign w29969 = ~w28934 & w29966;
assign w29970 = ~w29968 & ~w29969;
assign w29971 = (w29970 & w29369) | (w29970 & w45838) | (w29369 & w45838);
assign w29972 = ~w29402 & w29965;
assign w29973 = ~w29158 & w45839;
assign w29974 = ~w28808 & ~w28817;
assign w29975 = ~w29145 & w45840;
assign w29976 = ~w493 & ~w29975;
assign w29977 = ~w29973 & w29976;
assign w29978 = ~w28819 & ~w29968;
assign w29979 = ~w29965 & w29978;
assign w29980 = w29163 & ~w29979;
assign w29981 = (w29965 & w29141) | (w29965 & w45841) | (w29141 & w45841);
assign w29982 = w29978 & ~w29981;
assign w29983 = ~w28663 & w29980;
assign w29984 = w29982 & ~w29983;
assign w29985 = ~w29158 & w29984;
assign w29986 = (~w493 & w29156) | (~w493 & w49229) | (w29156 & w49229);
assign w29987 = ~w28835 & w28845;
assign w29988 = w400 & w29987;
assign w29989 = (w29988 & w29145) | (w29988 & w49230) | (w29145 & w49230);
assign w29990 = ~w29985 & w29989;
assign w29991 = w400 & ~w29987;
assign w29992 = ~w29983 & w45842;
assign w29993 = ~w29158 & w29992;
assign w29994 = ~w29145 & w49231;
assign w29995 = ~w29993 & ~w29994;
assign w29996 = ~w29990 & w29995;
assign w29997 = ~w29977 & w29996;
assign w29998 = ~w29159 & ~w29165;
assign w29999 = ~w29150 & ~w29159;
assign w30000 = w29146 & w29999;
assign w30001 = w28681 & w30000;
assign w30002 = ~w28663 & w30001;
assign w30003 = ~w29998 & ~w30002;
assign w30004 = w28763 & w28852;
assign w30005 = ~w30002 & w45843;
assign w30006 = ~w29158 & ~w30005;
assign w30007 = ~w30003 & ~w30004;
assign w30008 = w30006 & ~w30007;
assign w30009 = w28757 & ~w28758;
assign w30010 = ~w28757 & w28758;
assign w30011 = ~w30009 & ~w30010;
assign w30012 = ~w29145 & w45844;
assign w30013 = w351 & ~w30012;
assign w30014 = ~w30008 & w30013;
assign w30015 = ~w400 & ~w29987;
assign w30016 = (w30015 & w29145) | (w30015 & w49232) | (w29145 & w49232);
assign w30017 = ~w29985 & w30016;
assign w30018 = ~w400 & w29987;
assign w30019 = ~w29983 & w45845;
assign w30020 = ~w29158 & w30019;
assign w30021 = ~w29145 & w49233;
assign w30022 = ~w30020 & ~w30021;
assign w30023 = ~w30017 & w30022;
assign w30024 = ~w30014 & w30023;
assign w30025 = (~w30012 & ~w30006) | (~w30012 & w45846) | (~w30006 & w45846);
assign w30026 = ~w351 & ~w30025;
assign w30027 = w252 & w29180;
assign w30028 = ~w30026 & ~w30027;
assign w30029 = ~w29997 & w30024;
assign w30030 = w30028 & ~w30029;
assign w30031 = ~w29973 & ~w29975;
assign w30032 = w493 & ~w30031;
assign w30033 = w29996 & w30032;
assign w30034 = w30024 & ~w30033;
assign w30035 = w30030 & ~w30034;
assign w30036 = w28857 & w28884;
assign w30037 = w29142 & w30036;
assign w30038 = ~w28928 & ~w29155;
assign w30039 = (w30038 & w29369) | (w30038 & w47828) | (w29369 & w47828);
assign w30040 = w28912 & w30039;
assign w30041 = ~w28912 & ~w28916;
assign w30042 = ~w30039 & w30041;
assign w30043 = ~w30040 & ~w30042;
assign w30044 = w3 & w28926;
assign w30045 = (~w30044 & w28920) | (~w30044 & w42441) | (w28920 & w42441);
assign w30046 = ~w29143 & w30045;
assign w30047 = ~w28682 & w30046;
assign w30048 = ~w29156 & w49234;
assign w30049 = ~w30047 & ~w30048;
assign w30050 = ~w28856 & w42442;
assign w30051 = w42442 & w49235;
assign w30052 = w29142 & w30051;
assign w30053 = w28857 & w42443;
assign w30054 = ~w30052 & ~w30053;
assign w30055 = w29163 & ~w30053;
assign w30056 = ~w28663 & w30055;
assign w30057 = ~w30054 & ~w30056;
assign w30058 = ~w3 & ~w28926;
assign w30059 = (w30058 & ~w28857) | (w30058 & w42444) | (~w28857 & w42444);
assign w30060 = w29142 & w30050;
assign w30061 = w29163 & w30059;
assign w30062 = ~w28663 & w30061;
assign w30063 = w30059 & ~w30060;
assign w30064 = ~w30062 & ~w30063;
assign w30065 = ~w30057 & w30064;
assign w30066 = ~w30049 & w30065;
assign w30067 = w28870 & ~w30066;
assign w30068 = ~w28870 & w30066;
assign w30069 = ~w30067 & ~w30068;
assign w30070 = ~w42 & w30043;
assign w30071 = w30069 & w30070;
assign w30072 = ~w28765 & ~w28766;
assign w30073 = w28739 & w28852;
assign w30074 = ~w29165 & w47829;
assign w30075 = w30000 & w42445;
assign w30076 = ~w28663 & w30075;
assign w30077 = ~w30076 & w47830;
assign w30078 = ~w29158 & w30077;
assign w30079 = (w57 & w29156) | (w57 & w49236) | (w29156 & w49236);
assign w30080 = ~w29145 & w30079;
assign w30081 = w28701 & ~w28769;
assign w30082 = w80 & ~w30081;
assign w30083 = (w30082 & w29145) | (w30082 & w49237) | (w29145 & w49237);
assign w30084 = ~w30078 & w30083;
assign w30085 = w80 & w30081;
assign w30086 = ~w29145 & w49238;
assign w30087 = w30072 & w30085;
assign w30088 = ~w30076 & w47831;
assign w30089 = ~w29158 & w30088;
assign w30090 = ~w30086 & ~w30089;
assign w30091 = ~w30084 & w30090;
assign w30092 = ~w80 & ~w29157;
assign w30093 = ~w29145 & w30092;
assign w30094 = w28882 & ~w28926;
assign w30095 = ~w3 & w30094;
assign w30096 = (w30095 & w30093) | (w30095 & w47832) | (w30093 & w47832);
assign w30097 = ~w3 & ~w30094;
assign w30098 = ~w30093 & w47833;
assign w30099 = ~w30096 & ~w30098;
assign w30100 = w30091 & w30099;
assign w30101 = ~w30071 & w30100;
assign w30102 = ~w252 & ~w29180;
assign w30103 = ~w29145 & w42446;
assign w30104 = (~w28738 & w29168) | (~w28738 & w47834) | (w29168 & w47834);
assign w30105 = (w28743 & w29145) | (w28743 & w42447) | (w29145 & w42447);
assign w30106 = ~w28715 & ~w28766;
assign w30107 = ~w57 & w30106;
assign w30108 = w30103 & w30107;
assign w30109 = (w30107 & w29169) | (w30107 & w42448) | (w29169 & w42448);
assign w30110 = w30105 & w30109;
assign w30111 = ~w30108 & ~w30110;
assign w30112 = ~w30104 & w30105;
assign w30113 = ~w57 & ~w30106;
assign w30114 = ~w30103 & w30113;
assign w30115 = ~w30112 & w30114;
assign w30116 = w30111 & ~w30115;
assign w30117 = ~w30102 & w30116;
assign w30118 = (~w30043 & ~w30069) | (~w30043 & w42449) | (~w30069 & w42449);
assign w30119 = ~w28912 & ~w30039;
assign w30120 = ~w30040 & ~w30119;
assign w30121 = ~w29145 & w47835;
assign w30122 = w42 & ~w30121;
assign w30123 = (w30122 & ~w30069) | (w30122 & w42450) | (~w30069 & w42450);
assign w30124 = ~w30118 & ~w30123;
assign w30125 = ~w30093 & w47836;
assign w30126 = (w30094 & w30093) | (w30094 & w47837) | (w30093 & w47837);
assign w30127 = ~w30125 & ~w30126;
assign w30128 = w3 & w30127;
assign w30129 = ~w30071 & w30128;
assign w30130 = w30124 & ~w30129;
assign w30131 = ~w30078 & ~w30080;
assign w30132 = ~w80 & ~w30081;
assign w30133 = (w30132 & w30078) | (w30132 & w47838) | (w30078 & w47838);
assign w30134 = ~w80 & w30081;
assign w30135 = ~w30078 & w47839;
assign w30136 = ~w30133 & ~w30135;
assign w30137 = ~w30103 & ~w30112;
assign w30138 = w57 & ~w30106;
assign w30139 = (w30138 & w30112) | (w30138 & w47840) | (w30112 & w47840);
assign w30140 = w57 & w30106;
assign w30141 = ~w30112 & w47841;
assign w30142 = ~w30139 & ~w30141;
assign w30143 = w30136 & w30142;
assign w30144 = w30101 & ~w30143;
assign w30145 = w30130 & ~w30144;
assign w30146 = w30101 & w30117;
assign w30147 = ~w30035 & w30146;
assign w30148 = w30145 & ~w30147;
assign w30149 = w29963 & ~w30148;
assign w30150 = ~w29677 & w30149;
assign w30151 = w5745 & w29726;
assign w30152 = (w30151 & w29720) | (w30151 & w42451) | (w29720 & w42451);
assign w30153 = w5745 & ~w28597;
assign w30154 = ~w29720 & w42452;
assign w30155 = ~w30152 & ~w30154;
assign w30156 = ~w29158 & ~w30155;
assign w30157 = w5745 & ~w29733;
assign w30158 = (w30157 & w29156) | (w30157 & w49239) | (w29156 & w49239);
assign w30159 = ~w29145 & w30158;
assign w30160 = (w5330 & w29145) | (w5330 & w49240) | (w29145 & w49240);
assign w30161 = ~w30156 & w30160;
assign w30162 = w23494 & w29726;
assign w30163 = (w30162 & w29720) | (w30162 & w42453) | (w29720 & w42453);
assign w30164 = w23494 & ~w28597;
assign w30165 = ~w29720 & w42454;
assign w30166 = ~w30163 & ~w30165;
assign w30167 = ~w29145 & w49241;
assign w30168 = ~w29158 & ~w30166;
assign w30169 = ~w30167 & ~w30168;
assign w30170 = w29748 & w30169;
assign w30171 = ~w30161 & ~w30170;
assign w30172 = (~w4838 & w30170) | (~w4838 & w42455) | (w30170 & w42455);
assign w30173 = (w4838 & w30156) | (w4838 & w49242) | (w30156 & w49242);
assign w30174 = ~w30170 & w30173;
assign w30175 = w29760 & ~w30174;
assign w30176 = ~w30172 & ~w30175;
assign w30177 = ~w29145 & w42456;
assign w30178 = (w29687 & w29145) | (w29687 & w42457) | (w29145 & w42457);
assign w30179 = ~w30177 & ~w30178;
assign w30180 = w29707 & ~w30179;
assign w30181 = ~w29707 & w30179;
assign w30182 = ~w30180 & ~w30181;
assign w30183 = ~w4430 & ~w30182;
assign w30184 = ~w4056 & ~w29692;
assign w30185 = (w30184 & w29145) | (w30184 & w49243) | (w29145 & w49243);
assign w30186 = ~w29690 & w30185;
assign w30187 = ~w4056 & w29692;
assign w30188 = ~w29145 & w49244;
assign w30189 = w28532 & w30187;
assign w30190 = (w30189 & w29687) | (w30189 & w42458) | (w29687 & w42458);
assign w30191 = ~w29158 & w30190;
assign w30192 = ~w30188 & ~w30191;
assign w30193 = ~w30186 & w30192;
assign w30194 = w3646 & ~w29102;
assign w30195 = ~w29702 & ~w30194;
assign w30196 = w29701 & ~w30195;
assign w30197 = ~w29701 & w30195;
assign w30198 = ~w30196 & ~w30197;
assign w30199 = w30193 & ~w30198;
assign w30200 = w29706 & ~w30199;
assign w30201 = ~w30183 & ~w30200;
assign w30202 = ~w30176 & w30201;
assign w30203 = ~w29716 & ~w30200;
assign w30204 = w29822 & ~w30203;
assign w30205 = ~w30202 & w30204;
assign w30206 = ~w2006 & ~w29046;
assign w30207 = w29891 & w30206;
assign w30208 = ~w2006 & w29046;
assign w30209 = (w30208 & w29158) | (w30208 & w45847) | (w29158 & w45847);
assign w30210 = ~w29896 & ~w30209;
assign w30211 = ~w30207 & w30210;
assign w30212 = w29883 & ~w30211;
assign w30213 = w29863 & ~w30212;
assign w30214 = w29847 & ~w30213;
assign w30215 = (w3242 & ~w29158) | (w3242 & w42459) | (~w29158 & w42459);
assign w30216 = ~w29805 & w30215;
assign w30217 = ~w29145 & w42460;
assign w30218 = ~w2896 & ~w30217;
assign w30219 = ~w29158 & w29816;
assign w30220 = w30218 & ~w30219;
assign w30221 = ~w30216 & ~w30220;
assign w30222 = ~w29776 & ~w29787;
assign w30223 = (w2558 & w29158) | (w2558 & w45848) | (w29158 & w45848);
assign w30224 = w29082 & w29158;
assign w30225 = w30223 & ~w30224;
assign w30226 = ~w29784 & w30225;
assign w30227 = ~w29796 & ~w30226;
assign w30228 = w29794 & ~w29820;
assign w30229 = ~w30221 & w30228;
assign w30230 = w30227 & ~w30229;
assign w30231 = w29952 & w30230;
assign w30232 = ~w30214 & w30231;
assign w30233 = ~w30205 & w30232;
assign w30234 = w29962 & ~w30233;
assign w30235 = ~w30030 & w30146;
assign w30236 = ~w30235 & w30145;
assign w30237 = (w30236 & w30233) | (w30236 & w49245) | (w30233 & w49245);
assign w30238 = (~w30148 & w30234) | (~w30148 & w42461) | (w30234 & w42461);
assign w30239 = (~w30238 & w29677) | (~w30238 & w42462) | (w29677 & w42462);
assign w30240 = w29180 & w30239;
assign w30241 = ~w30027 & ~w30102;
assign w30242 = ~w29963 & ~w30234;
assign w30243 = (w30034 & w30234) | (w30034 & w49246) | (w30234 & w49246);
assign w30244 = w29677 & w29997;
assign w30245 = w30243 & ~w30244;
assign w30246 = ~w30205 & w30230;
assign w30247 = w29952 & ~w30214;
assign w30248 = (w30247 & w45849) | (w30247 & w45850) | (w45849 & w45850);
assign w30249 = w29962 & ~w30246;
assign w30250 = w30248 & ~w30249;
assign w30251 = (w30241 & w30245) | (w30241 & w42464) | (w30245 & w42464);
assign w30252 = ~w30239 & ~w30251;
assign w30253 = ~w30245 & w42465;
assign w30254 = w57 & w30240;
assign w30255 = (w57 & w30245) | (w57 & w47842) | (w30245 & w47842);
assign w30256 = w30252 & w30255;
assign w30257 = ~w30254 & ~w30256;
assign w30258 = ~w29677 & w29963;
assign w30259 = (w30250 & w29677) | (w30250 & w42466) | (w29677 & w42466);
assign w30260 = w30023 & ~w30033;
assign w30261 = ~w30239 & w50136;
assign w30262 = ~w30014 & ~w30026;
assign w30263 = w252 & ~w30262;
assign w30264 = (w30263 & w30261) | (w30263 & w45851) | (w30261 & w45851);
assign w30265 = w252 & w30262;
assign w30266 = ~w30261 & w45852;
assign w30267 = ~w30264 & ~w30266;
assign w30268 = w30257 & w30267;
assign w30269 = ~w57 & ~w30240;
assign w30270 = w30252 & ~w30253;
assign w30271 = w30269 & ~w30270;
assign w30272 = ~w400 & ~w30238;
assign w30273 = ~w30150 & w30272;
assign w30274 = ~w29977 & w30238;
assign w30275 = w29963 & w42467;
assign w30276 = ~w29677 & w30275;
assign w30277 = ~w30274 & ~w30276;
assign w30278 = w29677 & ~w30234;
assign w30279 = (~w30032 & w30234) | (~w30032 & w49247) | (w30234 & w49247);
assign w30280 = ~w30278 & w30279;
assign w30281 = ~w30277 & ~w30280;
assign w30282 = ~w30273 & ~w30281;
assign w30283 = w29996 & w30023;
assign w30284 = ~w351 & w30283;
assign w30285 = (w30284 & w30281) | (w30284 & w42468) | (w30281 & w42468);
assign w30286 = ~w30148 & w30234;
assign w30287 = ~w493 & w30236;
assign w30288 = ~w29977 & ~w30032;
assign w30289 = w400 & ~w30288;
assign w30290 = (w30289 & w30150) | (w30289 & w42469) | (w30150 & w42469);
assign w30291 = w400 & w30288;
assign w30292 = ~w30150 & w42470;
assign w30293 = ~w30290 & ~w30292;
assign w30294 = ~w351 & ~w30283;
assign w30295 = (w30294 & w30150) | (w30294 & w42471) | (w30150 & w42471);
assign w30296 = ~w30281 & w30295;
assign w30297 = w30293 & ~w30296;
assign w30298 = ~w30285 & w30297;
assign w30299 = ~w29926 & w30238;
assign w30300 = w29963 & w42472;
assign w30301 = ~w29677 & w30300;
assign w30302 = ~w30299 & ~w30301;
assign w30303 = w29951 & ~w30214;
assign w30304 = w29958 & ~w30303;
assign w30305 = w30246 & ~w30304;
assign w30306 = w29677 & w30305;
assign w30307 = w29847 & w29899;
assign w30308 = ~w29823 & w30246;
assign w30309 = w29958 & w50219;
assign w30310 = ~w30306 & w30309;
assign w30311 = ~w30302 & ~w30310;
assign w30312 = w612 & ~w30238;
assign w30313 = ~w30150 & w30312;
assign w30314 = ~w29914 & ~w29928;
assign w30315 = w493 & ~w30314;
assign w30316 = (w30315 & w30311) | (w30315 & w42474) | (w30311 & w42474);
assign w30317 = ~w400 & w30288;
assign w30318 = (w30317 & w30150) | (w30317 & w42475) | (w30150 & w42475);
assign w30319 = ~w400 & ~w30288;
assign w30320 = ~w30150 & w42476;
assign w30321 = ~w30318 & ~w30320;
assign w30322 = w493 & w30314;
assign w30323 = (w30322 & w30150) | (w30322 & w42477) | (w30150 & w42477);
assign w30324 = ~w30311 & w30323;
assign w30325 = w30321 & ~w30324;
assign w30326 = ~w30316 & w30325;
assign w30327 = ~w30281 & w42478;
assign w30328 = w351 & ~w30327;
assign w30329 = ~w30282 & w30283;
assign w30330 = w30328 & ~w30329;
assign w30331 = w30298 & ~w30326;
assign w30332 = ~w30330 & ~w30331;
assign w30333 = ~w493 & ~w30314;
assign w30334 = ~w30311 & w42479;
assign w30335 = ~w493 & w30314;
assign w30336 = (w30335 & w30311) | (w30335 & w42480) | (w30311 & w42480);
assign w30337 = ~w30334 & ~w30336;
assign w30338 = w30298 & w30337;
assign w30339 = ~w29797 & w29901;
assign w30340 = (w30339 & ~w30246) | (w30339 & w47843) | (~w30246 & w47843);
assign w30341 = (w30340 & ~w29677) | (w30340 & w42481) | (~w29677 & w42481);
assign w30342 = (~w29956 & w30341) | (~w29956 & w47844) | (w30341 & w47844);
assign w30343 = ~w754 & ~w30239;
assign w30344 = ~w30239 & w30342;
assign w30345 = ~w29925 & ~w30343;
assign w30346 = w29925 & w30343;
assign w30347 = ~w30345 & ~w30346;
assign w30348 = ~w30344 & w30347;
assign w30349 = ~w29958 & ~w30239;
assign w30350 = ~w29926 & ~w30349;
assign w30351 = w30342 & ~w30350;
assign w30352 = w612 & ~w30351;
assign w30353 = ~w30348 & w30352;
assign w30354 = w30338 & w30353;
assign w30355 = w30332 & ~w30354;
assign w30356 = ~w30261 & w45853;
assign w30357 = (w30262 & w30261) | (w30262 & w45854) | (w30261 & w45854);
assign w30358 = ~w30356 & ~w30357;
assign w30359 = ~w252 & ~w30358;
assign w30360 = ~w30268 & ~w30271;
assign w30361 = ~w30271 & ~w30359;
assign w30362 = (~w30360 & ~w30355) | (~w30360 & w42482) | (~w30355 & w42482);
assign w30363 = (w30030 & w30278) | (w30030 & w42483) | (w30278 & w42483);
assign w30364 = w30117 & ~w30363;
assign w30365 = ~w42 & ~w30069;
assign w30366 = w30128 & w30365;
assign w30367 = w30143 & ~w30366;
assign w30368 = ~w30100 & ~w30128;
assign w30369 = w30365 & ~w30368;
assign w30370 = ~w30364 & w30367;
assign w30371 = w30369 & ~w30370;
assign w30372 = w30100 & ~w30143;
assign w30373 = w30100 & w30117;
assign w30374 = ~w30043 & w30372;
assign w30375 = ~w30043 & w30373;
assign w30376 = ~w30363 & w30375;
assign w30377 = ~w30374 & ~w30376;
assign w30378 = ~w30043 & w30128;
assign w30379 = w30069 & ~w30378;
assign w30380 = ~w42 & w30379;
assign w30381 = w30377 & w30380;
assign w30382 = ~w30371 & ~w30381;
assign w30383 = w30091 & ~w30239;
assign w30384 = w3 & w30239;
assign w30385 = ~w30383 & ~w30384;
assign w30386 = w30143 & ~w30384;
assign w30387 = ~w30364 & w30386;
assign w30388 = ~w30385 & ~w30387;
assign w30389 = w30099 & ~w30128;
assign w30390 = w30388 & ~w30389;
assign w30391 = ~w30388 & w30389;
assign w30392 = ~w30390 & ~w30391;
assign w30393 = ~w30382 & w30392;
assign w30394 = w42 & ~w30389;
assign w30395 = w30388 & w30394;
assign w30396 = w42 & w30389;
assign w30397 = ~w30388 & w30396;
assign w30398 = ~w30395 & ~w30397;
assign w30399 = ~w30363 & w30373;
assign w30400 = ~w30372 & ~w30399;
assign w30401 = ~w30128 & w30400;
assign w30402 = w42 & ~w30069;
assign w30403 = w30143 & ~w30364;
assign w30404 = w30128 & w30402;
assign w30405 = w30100 & w30402;
assign w30406 = ~w30403 & w30405;
assign w30407 = ~w30404 & ~w30406;
assign w30408 = w30365 & w30401;
assign w30409 = w30407 & ~w30408;
assign w30410 = w30398 & w30409;
assign w30411 = ~w42 & w30100;
assign w30412 = w126 & w30127;
assign w30413 = ~w30411 & ~w30412;
assign w30414 = w30143 & ~w30412;
assign w30415 = ~w30364 & w30414;
assign w30416 = ~w30413 & ~w30415;
assign w30417 = w30069 & ~w30128;
assign w30418 = ~w30124 & w30417;
assign w30419 = w30400 & w30418;
assign w30420 = ~w30416 & ~w30419;
assign w30421 = w30382 & ~w30420;
assign w30422 = w30091 & w30136;
assign w30423 = ~w30239 & ~w30422;
assign w30424 = w30142 & ~w30364;
assign w30425 = w30423 & ~w30424;
assign w30426 = w30143 & w30383;
assign w30427 = ~w30364 & w30426;
assign w30428 = w30081 & ~w30131;
assign w30429 = ~w30081 & w30131;
assign w30430 = ~w30428 & ~w30429;
assign w30431 = w30239 & w30430;
assign w30432 = ~w30427 & ~w30431;
assign w30433 = ~w30425 & w30432;
assign w30434 = ~w3 & w30433;
assign w30435 = ~w30421 & w30434;
assign w30436 = w30410 & w30435;
assign w30437 = ~w30106 & w30137;
assign w30438 = w30106 & ~w30137;
assign w30439 = ~w30437 & ~w30438;
assign w30440 = ~w30439 & ~w30239;
assign w30441 = w57 & ~w30440;
assign w30442 = ~w30102 & ~w30363;
assign w30443 = ~w30116 & ~w30239;
assign w30444 = w30142 & ~w30443;
assign w30445 = w57 & w30035;
assign w30446 = ~w30234 & w30445;
assign w30447 = (w30446 & w29677) | (w30446 & w42484) | (w29677 & w42484);
assign w30448 = w30239 & w30439;
assign w30449 = ~w30239 & w30447;
assign w30450 = ~w30439 & w30449;
assign w30451 = ~w30448 & ~w30450;
assign w30452 = w30442 & ~w30444;
assign w30453 = w30451 & ~w30452;
assign w30454 = ~w30441 & ~w30442;
assign w30455 = w30116 & w30454;
assign w30456 = w30453 & ~w30455;
assign w30457 = w80 & w30456;
assign w30458 = ~w30393 & ~w30457;
assign w30459 = ~w30436 & w30458;
assign w30460 = ~w30362 & w30459;
assign w30461 = w30410 & ~w30421;
assign w30462 = w3 & ~w30433;
assign w30463 = (~w80 & ~w30453) | (~w80 & w47845) | (~w30453 & w47845);
assign w30464 = ~w30462 & ~w30463;
assign w30465 = ~w30434 & ~w30464;
assign w30466 = w30461 & ~w30465;
assign w30467 = ~w30393 & ~w30466;
assign w30468 = ~w30460 & ~w30467;
assign w30469 = ~w29950 & ~w30214;
assign w30470 = w30307 & w50220;
assign w30471 = w30469 & ~w30470;
assign w30472 = w29943 & ~w29956;
assign w30473 = w29955 & w30239;
assign w30474 = ~w30472 & ~w30239;
assign w30475 = w30471 & w30474;
assign w30476 = w30472 & ~w30239;
assign w30477 = ~w30471 & w30476;
assign w30478 = ~w30475 & ~w30477;
assign w30479 = ~w30473 & w30478;
assign w30480 = w754 & ~w30479;
assign w30481 = w29899 & w50220;
assign w30482 = ~w29835 & ~w30239;
assign w30483 = w30213 & ~w30481;
assign w30484 = w30482 & ~w30483;
assign w30485 = w1120 & w30239;
assign w30486 = ~w29846 & ~w29950;
assign w30487 = ~w945 & w30486;
assign w30488 = (w30487 & w30484) | (w30487 & w47846) | (w30484 & w47846);
assign w30489 = ~w945 & ~w30486;
assign w30490 = ~w30484 & w47847;
assign w30491 = ~w30488 & ~w30490;
assign w30492 = ~w30480 & w30491;
assign w30493 = w945 & ~w30486;
assign w30494 = (w30493 & w30484) | (w30493 & w47848) | (w30484 & w47848);
assign w30495 = w945 & w30486;
assign w30496 = ~w30484 & w47849;
assign w30497 = ~w30494 & ~w30496;
assign w30498 = w29834 & w30239;
assign w30499 = ~w29835 & w29862;
assign w30500 = ~w30498 & ~w30499;
assign w30501 = ~w29857 & ~w30212;
assign w30502 = ~w30481 & w30501;
assign w30503 = w30500 & ~w30502;
assign w30504 = ~w29835 & ~w30498;
assign w30505 = ~w30484 & w30504;
assign w30506 = ~w30503 & ~w30505;
assign w30507 = (w1120 & w30505) | (w1120 & w47850) | (w30505 & w47850);
assign w30508 = w30497 & ~w30507;
assign w30509 = w30492 & ~w30508;
assign w30510 = w30268 & w30338;
assign w30511 = ~w754 & w30479;
assign w30512 = (~w612 & w30348) | (~w612 & w47851) | (w30348 & w47851);
assign w30513 = ~w30511 & ~w30512;
assign w30514 = w30510 & w30513;
assign w30515 = w30464 & w30514;
assign w30516 = w30461 & w30515;
assign w30517 = ~w30509 & w30516;
assign w30518 = ~w30468 & ~w30517;
assign w30519 = ~a[14] & ~a[15];
assign w30520 = ~a[16] & w30519;
assign w30521 = ~w29158 & w30520;
assign w30522 = w29158 & ~w30520;
assign w30523 = w29405 & ~w30521;
assign w30524 = a[17] & w30522;
assign w30525 = ~w30523 & ~w30524;
assign w30526 = w30238 & ~w30525;
assign w30527 = w29963 & w42485;
assign w30528 = ~w29677 & w30527;
assign w30529 = ~w30526 & ~w30528;
assign w30530 = a[17] & ~w30521;
assign w30531 = ~w30522 & ~w30530;
assign w30532 = w30236 & ~w30531;
assign w30533 = ~w30234 & w30532;
assign w30534 = ~w30533 & w42486;
assign w30535 = w29963 & w45855;
assign w30536 = ~w29677 & w30535;
assign w30537 = ~w30534 & ~w30536;
assign w30538 = a[19] & ~w29158;
assign w30539 = ~a[19] & w29158;
assign w30540 = ~w30538 & ~w30539;
assign w30541 = w28077 & w30540;
assign w30542 = ~w28077 & ~w30540;
assign w30543 = ~w30541 & ~w30542;
assign w30544 = w29406 & ~w30543;
assign w30545 = ~w29406 & w30543;
assign w30546 = ~w30544 & ~w30545;
assign w30547 = w26880 & ~w30546;
assign w30548 = w29963 & w42487;
assign w30549 = ~w29677 & w30548;
assign w30550 = w30238 & w30547;
assign w30551 = ~w30549 & ~w30550;
assign w30552 = ~a[18] & ~w30540;
assign w30553 = ~w29403 & ~w30552;
assign w30554 = w26880 & w30553;
assign w30555 = ~w30238 & w30554;
assign w30556 = ~w30150 & w30555;
assign w30557 = w30551 & ~w30556;
assign w30558 = a[18] & ~w29405;
assign w30559 = ~w29406 & ~w30558;
assign w30560 = (w30559 & w30147) | (w30559 & w47852) | (w30147 & w47852);
assign w30561 = ~w30030 & w30117;
assign w30562 = w30143 & ~w30561;
assign w30563 = w30130 & w30562;
assign w30564 = ~w30234 & w30563;
assign w30565 = w29963 & w30560;
assign w30566 = ~w29677 & w30565;
assign w30567 = (w30560 & w30234) | (w30560 & w47853) | (w30234 & w47853);
assign w30568 = ~w30566 & ~w30567;
assign w30569 = ~w28077 & ~w30525;
assign w30570 = a[18] & ~w29158;
assign w30571 = ~a[18] & w29158;
assign w30572 = ~w30570 & ~w30571;
assign w30573 = ~w30238 & ~w30572;
assign w30574 = ~w30150 & w30573;
assign w30575 = ~w28077 & ~w30531;
assign w30576 = ~a[19] & ~w30575;
assign w30577 = ~w30150 & w42488;
assign w30578 = ~w30543 & ~w30569;
assign w30579 = (w30578 & w30566) | (w30578 & w42489) | (w30566 & w42489);
assign w30580 = ~w30577 & ~w30579;
assign w30581 = w30529 & ~w30537;
assign w30582 = w30557 & w30581;
assign w30583 = w30580 & ~w30582;
assign w30584 = w30568 & ~w30574;
assign w30585 = w30569 & ~w30239;
assign w30586 = w30575 & w30239;
assign w30587 = ~w30585 & ~w30586;
assign w30588 = ~w26880 & ~w30584;
assign w30589 = w30587 & w30588;
assign w30590 = w24874 & w29400;
assign w30591 = ~w30238 & ~w30590;
assign w30592 = ~w29401 & ~w29474;
assign w30593 = w29439 & ~w30592;
assign w30594 = ~w29439 & w30592;
assign w30595 = ~w30593 & ~w30594;
assign w30596 = w24874 & w30595;
assign w30597 = w30238 & ~w30596;
assign w30598 = w29963 & w42490;
assign w30599 = ~w29677 & w30598;
assign w30600 = ~w30597 & ~w30599;
assign w30601 = ~w30150 & w30591;
assign w30602 = w30600 & ~w30601;
assign w30603 = (w24874 & w29440) | (w24874 & w42491) | (w29440 & w42491);
assign w30604 = ~w29440 & w42492;
assign w30605 = ~w30603 & ~w30604;
assign w30606 = (w30605 & w30147) | (w30605 & w47854) | (w30147 & w47854);
assign w30607 = w29963 & w30606;
assign w30608 = ~w29677 & w30607;
assign w30609 = w23843 & ~w29484;
assign w30610 = (w30609 & w30237) | (w30609 & w42493) | (w30237 & w42493);
assign w30611 = ~w30608 & w30610;
assign w30612 = w23843 & w29484;
assign w30613 = w29963 & w42494;
assign w30614 = ~w29677 & w30613;
assign w30615 = ~w30237 & w42494;
assign w30616 = ~w30614 & ~w30615;
assign w30617 = ~w30611 & w30616;
assign w30618 = ~w30602 & w30617;
assign w30619 = ~w26880 & ~w30553;
assign w30620 = ~w30238 & ~w30619;
assign w30621 = ~w26880 & w30546;
assign w30622 = w30238 & ~w30621;
assign w30623 = w29963 & w47855;
assign w30624 = ~w29677 & w30623;
assign w30625 = ~w30622 & ~w30624;
assign w30626 = ~w30150 & w30620;
assign w30627 = w30625 & ~w30626;
assign w30628 = ~w29424 & ~w29425;
assign w30629 = (w30628 & w30147) | (w30628 & w42495) | (w30147 & w42495);
assign w30630 = w29963 & w30629;
assign w30631 = ~w29677 & w30630;
assign w30632 = (w30629 & w30234) | (w30629 & w42496) | (w30234 & w42496);
assign w30633 = w25851 & ~w29437;
assign w30634 = ~w30632 & w30633;
assign w30635 = ~w30631 & w30634;
assign w30636 = w25851 & w29437;
assign w30637 = w29963 & w47856;
assign w30638 = ~w29677 & w30637;
assign w30639 = w30632 & w30636;
assign w30640 = ~w30638 & ~w30639;
assign w30641 = ~w30635 & w30640;
assign w30642 = ~w30627 & w30641;
assign w30643 = w30618 & w30642;
assign w30644 = w30583 & ~w30589;
assign w30645 = w30643 & w30644;
assign w30646 = ~w24874 & ~w29400;
assign w30647 = ~w30238 & ~w30646;
assign w30648 = ~w24874 & ~w30595;
assign w30649 = w30238 & ~w30648;
assign w30650 = w29963 & w42497;
assign w30651 = ~w29677 & w30650;
assign w30652 = ~w30649 & ~w30651;
assign w30653 = ~w30150 & w30647;
assign w30654 = w30652 & ~w30653;
assign w30655 = ~w25851 & w29437;
assign w30656 = ~w30632 & w30655;
assign w30657 = ~w30631 & w30656;
assign w30658 = ~w25851 & ~w29437;
assign w30659 = w29963 & w42498;
assign w30660 = ~w29677 & w30659;
assign w30661 = w30632 & w30658;
assign w30662 = ~w30660 & ~w30661;
assign w30663 = ~w30657 & w30662;
assign w30664 = ~w30654 & w30663;
assign w30665 = w30618 & ~w30664;
assign w30666 = (w29484 & w30608) | (w29484 & w42499) | (w30608 & w42499);
assign w30667 = ~w30608 & w42500;
assign w30668 = ~w30666 & ~w30667;
assign w30669 = ~w23843 & w30668;
assign w30670 = ~w30665 & ~w30669;
assign w30671 = w28105 & ~w29460;
assign w30672 = ~w28105 & w29460;
assign w30673 = ~w30671 & ~w30672;
assign w30674 = w29465 & w29494;
assign w30675 = (~w29489 & w29440) | (~w29489 & w42501) | (w29440 & w42501);
assign w30676 = w30674 & ~w30675;
assign w30677 = ~w30674 & w30675;
assign w30678 = w30673 & w30239;
assign w30679 = ~w30676 & ~w30677;
assign w30680 = w30679 & ~w30239;
assign w30681 = ~w30678 & ~w30680;
assign w30682 = ~w22767 & ~w30681;
assign w30683 = ~w30665 & w42502;
assign w30684 = ~w30645 & w30683;
assign w30685 = ~w29447 & w29451;
assign w30686 = w28149 & ~w29451;
assign w30687 = ~w30685 & ~w30686;
assign w30688 = w29494 & ~w30676;
assign w30689 = w22767 & ~w30688;
assign w30690 = ~w22767 & w30688;
assign w30691 = ~w30689 & ~w30690;
assign w30692 = ~w30691 & ~w30239;
assign w30693 = w30687 & ~w30692;
assign w30694 = ~w30687 & w30692;
assign w30695 = ~w30693 & ~w30694;
assign w30696 = ~w21801 & ~w30695;
assign w30697 = w29457 & ~w29500;
assign w30698 = w29470 & w30688;
assign w30699 = w29456 & ~w30698;
assign w30700 = w30697 & ~w30699;
assign w30701 = ~w30697 & w30699;
assign w30702 = ~w30700 & ~w30701;
assign w30703 = ~w29499 & w30239;
assign w30704 = ~w30239 & w30702;
assign w30705 = ~w30703 & ~w30704;
assign w30706 = (w20906 & w30704) | (w20906 & w45856) | (w30704 & w45856);
assign w30707 = ~w29496 & ~w29500;
assign w30708 = w29472 & ~w30675;
assign w30709 = w30707 & ~w30708;
assign w30710 = w20906 & ~w30709;
assign w30711 = ~w20906 & w30709;
assign w30712 = ~w30710 & ~w30711;
assign w30713 = ~w30712 & ~w30239;
assign w30714 = ~w20000 & ~w29509;
assign w30715 = w30713 & w30714;
assign w30716 = ~w20000 & w29509;
assign w30717 = ~w30713 & w30716;
assign w30718 = ~w30715 & ~w30717;
assign w30719 = ~w30706 & w30718;
assign w30720 = ~w30696 & w30719;
assign w30721 = w29247 & ~w29264;
assign w30722 = ~w29515 & ~w29516;
assign w30723 = w30721 & ~w30722;
assign w30724 = ~w30721 & w30722;
assign w30725 = ~w30723 & ~w30724;
assign w30726 = w29263 & w30239;
assign w30727 = ~w30725 & ~w30239;
assign w30728 = ~w30726 & ~w30727;
assign w30729 = ~w19040 & w30728;
assign w30730 = w22767 & w30681;
assign w30731 = ~w30729 & ~w30730;
assign w30732 = w30720 & w30731;
assign w30733 = ~w30684 & w30732;
assign w30734 = w21801 & ~w30687;
assign w30735 = ~w30692 & w30734;
assign w30736 = w21801 & w30687;
assign w30737 = w30692 & w30736;
assign w30738 = ~w30735 & ~w30737;
assign w30739 = ~w30704 & w45857;
assign w30740 = w30738 & ~w30739;
assign w30741 = w30719 & ~w30740;
assign w30742 = ~w29214 & ~w29223;
assign w30743 = (~w29264 & w29515) | (~w29264 & w42503) | (w29515 & w42503);
assign w30744 = w29247 & ~w30743;
assign w30745 = w30742 & ~w30744;
assign w30746 = ~w30742 & w30744;
assign w30747 = ~w30745 & ~w30746;
assign w30748 = ~w29213 & w30239;
assign w30749 = ~w30747 & ~w30239;
assign w30750 = ~w30748 & ~w30749;
assign w30751 = w18183 & ~w30750;
assign w30752 = ~w19040 & w29158;
assign w30753 = ~w29158 & w29182;
assign w30754 = ~w30752 & ~w30753;
assign w30755 = w29181 & ~w30754;
assign w30756 = ~w29181 & w30754;
assign w30757 = ~w30755 & ~w30756;
assign w30758 = w29221 & ~w29258;
assign w30759 = w29248 & ~w30743;
assign w30760 = ~w29214 & ~w30759;
assign w30761 = w30758 & ~w30760;
assign w30762 = ~w30758 & w30760;
assign w30763 = ~w30761 & ~w30762;
assign w30764 = w30757 & w30239;
assign w30765 = ~w30239 & ~w30763;
assign w30766 = ~w30764 & ~w30765;
assign w30767 = ~w30765 & w45858;
assign w30768 = ~w30751 & ~w30767;
assign w30769 = w19040 & ~w30728;
assign w30770 = w20000 & ~w29509;
assign w30771 = ~w30713 & w30770;
assign w30772 = w20000 & w29509;
assign w30773 = w30713 & w30772;
assign w30774 = ~w30771 & ~w30773;
assign w30775 = ~w30769 & w30774;
assign w30776 = w30729 & w30768;
assign w30777 = w30768 & w30775;
assign w30778 = ~w30741 & w30777;
assign w30779 = ~w30776 & ~w30778;
assign w30780 = ~w30733 & ~w30779;
assign w30781 = ~w29287 & w29363;
assign w30782 = ~w29202 & w29358;
assign w30783 = ~w29265 & w29358;
assign w30784 = w29260 & w30783;
assign w30785 = ~w30782 & ~w30784;
assign w30786 = w29260 & w42504;
assign w30787 = (w29338 & ~w30785) | (w29338 & w42505) | (~w30785 & w42505);
assign w30788 = w29338 & w30786;
assign w30789 = ~w29515 & w30788;
assign w30790 = ~w30787 & ~w30789;
assign w30791 = (~w29277 & w30789) | (~w29277 & w42506) | (w30789 & w42506);
assign w30792 = ~w29657 & ~w30791;
assign w30793 = w30781 & ~w30792;
assign w30794 = ~w30781 & w30792;
assign w30795 = ~w30793 & ~w30794;
assign w30796 = w29286 & w30239;
assign w30797 = ~w30239 & w30795;
assign w30798 = ~w30796 & ~w30797;
assign w30799 = (w11138 & w30797) | (w11138 & w45859) | (w30797 & w45859);
assign w30800 = (w30237 & w29677) | (w30237 & w42507) | (w29677 & w42507);
assign w30801 = (~w12666 & w30789) | (~w12666 & w42508) | (w30789 & w42508);
assign w30802 = ~w30148 & ~w30801;
assign w30803 = w12666 & w30790;
assign w30804 = w30802 & ~w30803;
assign w30805 = w29276 & w30237;
assign w30806 = ~w30258 & w30805;
assign w30807 = w30802 & w50385;
assign w30808 = ~w30800 & w30807;
assign w30809 = w29276 & ~w30804;
assign w30810 = ~w30806 & ~w30809;
assign w30811 = ~w30808 & w30810;
assign w30812 = (~w11870 & ~w30810) | (~w11870 & w42509) | (~w30810 & w42509);
assign w30813 = ~w30799 & ~w30812;
assign w30814 = ~w29302 & w29311;
assign w30815 = ~w29515 & w30786;
assign w30816 = (~w29336 & w30815) | (~w29336 & w42510) | (w30815 & w42510);
assign w30817 = w29321 & ~w30816;
assign w30818 = w30814 & ~w30817;
assign w30819 = ~w30814 & w30817;
assign w30820 = ~w30818 & ~w30819;
assign w30821 = w29301 & w30239;
assign w30822 = ~w30239 & w30820;
assign w30823 = ~w30821 & ~w30822;
assign w30824 = (~w12666 & w30822) | (~w12666 & w45860) | (w30822 & w45860);
assign w30825 = w30810 & w42511;
assign w30826 = w30824 & ~w30825;
assign w30827 = w30813 & ~w30826;
assign w30828 = w30785 & w42512;
assign w30829 = ~w30815 & w30828;
assign w30830 = (w14766 & ~w30785) | (w14766 & w42513) | (~w30785 & w42513);
assign w30831 = w14766 & w30786;
assign w30832 = ~w29515 & w30831;
assign w30833 = ~w30830 & ~w30832;
assign w30834 = ~w28458 & w29158;
assign w30835 = ~w29158 & w29330;
assign w30836 = ~w30834 & ~w30835;
assign w30837 = ~w30832 & w42514;
assign w30838 = ~w30829 & ~w30837;
assign w30839 = w14039 & ~w30838;
assign w30840 = ~w14039 & w30838;
assign w30841 = ~w30839 & ~w30840;
assign w30842 = ~w30239 & w30841;
assign w30843 = w28438 & w29158;
assign w30844 = ~w29158 & w29316;
assign w30845 = ~w30843 & ~w30844;
assign w30846 = w30842 & w30845;
assign w30847 = ~w30842 & ~w30845;
assign w30848 = ~w30846 & ~w30847;
assign w30849 = ~w13384 & ~w30848;
assign w30850 = ~w11138 & w30798;
assign w30851 = ~w30822 & w47857;
assign w30852 = ~w30825 & ~w30851;
assign w30853 = w30813 & ~w30852;
assign w30854 = ~w30850 & ~w30853;
assign w30855 = w30827 & w30849;
assign w30856 = w30854 & ~w30855;
assign w30857 = ~w18183 & w30750;
assign w30858 = ~w30767 & w30857;
assign w30859 = w17380 & ~w30766;
assign w30860 = ~w30858 & ~w30859;
assign w30861 = ~w29222 & ~w29258;
assign w30862 = ~w29264 & ~w30861;
assign w30863 = ~w29249 & ~w29258;
assign w30864 = w29265 & w29516;
assign w30865 = w30863 & ~w30864;
assign w30866 = (w30865 & ~w29515) | (w30865 & w42515) | (~w29515 & w42515);
assign w30867 = w17380 & ~w30866;
assign w30868 = ~w17380 & w30866;
assign w30869 = ~w30867 & ~w30868;
assign w30870 = ~w30148 & w30869;
assign w30871 = ~w29200 & w30237;
assign w30872 = ~w30258 & w30871;
assign w30873 = w29200 & w30870;
assign w30874 = ~w30800 & w30873;
assign w30875 = ~w29200 & ~w30870;
assign w30876 = ~w30872 & ~w30875;
assign w30877 = ~w30874 & w30876;
assign w30878 = (w29343 & w30147) | (w29343 & w42516) | (w30147 & w42516);
assign w30879 = (w29266 & w29515) | (w29266 & w42517) | (w29515 & w42517);
assign w30880 = w30878 & ~w30879;
assign w30881 = w29254 & w30866;
assign w30882 = ~w29201 & ~w30881;
assign w30883 = w29192 & ~w30882;
assign w30884 = w30880 & ~w30883;
assign w30885 = ~w30148 & ~w30882;
assign w30886 = ~w29191 & w30237;
assign w30887 = ~w30258 & w30886;
assign w30888 = ~w29191 & ~w30878;
assign w30889 = ~w30885 & w30888;
assign w30890 = ~w30887 & ~w30889;
assign w30891 = ~w30800 & w30884;
assign w30892 = w30890 & ~w30891;
assign w30893 = ~w16559 & w30877;
assign w30894 = ~w15681 & ~w30892;
assign w30895 = ~w30893 & ~w30894;
assign w30896 = w30860 & w30895;
assign w30897 = ~w30829 & w30833;
assign w30898 = w30149 & w30897;
assign w30899 = ~w29677 & w30898;
assign w30900 = (~w30836 & w30899) | (~w30836 & w42518) | (w30899 & w42518);
assign w30901 = ~w30899 & w42519;
assign w30902 = ~w30900 & ~w30901;
assign w30903 = w14039 & w30902;
assign w30904 = ~w30237 & w30880;
assign w30905 = w29963 & w30880;
assign w30906 = ~w29677 & w30905;
assign w30907 = ~w30904 & ~w30906;
assign w30908 = w15681 & ~w30238;
assign w30909 = ~w30150 & w30908;
assign w30910 = w30907 & ~w30909;
assign w30911 = ~w29357 & w29647;
assign w30912 = ~w14766 & w30911;
assign w30913 = ~w30910 & w30912;
assign w30914 = ~w14766 & ~w30911;
assign w30915 = w30910 & w30914;
assign w30916 = ~w30913 & ~w30915;
assign w30917 = ~w30903 & w30916;
assign w30918 = ~w14039 & ~w30902;
assign w30919 = w13384 & w30845;
assign w30920 = (w30919 & w30239) | (w30919 & w47858) | (w30239 & w47858);
assign w30921 = w13384 & ~w30845;
assign w30922 = ~w30239 & w47859;
assign w30923 = ~w30920 & ~w30922;
assign w30924 = ~w30918 & w30923;
assign w30925 = ~w30917 & w30924;
assign w30926 = w30827 & w30925;
assign w30927 = w30896 & ~w30926;
assign w30928 = w30856 & w30927;
assign w30929 = ~w30780 & w30928;
assign w30930 = w30910 & ~w30911;
assign w30931 = ~w30910 & w30911;
assign w30932 = ~w30930 & ~w30931;
assign w30933 = w14766 & w30932;
assign w30934 = (w16559 & ~w30876) | (w16559 & w42520) | (~w30876 & w42520);
assign w30935 = w30890 & w42521;
assign w30936 = ~w30934 & ~w30935;
assign w30937 = ~w30894 & ~w30936;
assign w30938 = ~w30933 & ~w30937;
assign w30939 = (w30917 & w30937) | (w30917 & w45861) | (w30937 & w45861);
assign w30940 = w30827 & w30924;
assign w30941 = ~w30939 & w30940;
assign w30942 = w30856 & ~w30941;
assign w30943 = ~w30929 & ~w30942;
assign w30944 = ~w29537 & ~w29591;
assign w30945 = ~w29368 & ~w29658;
assign w30946 = ~w29519 & w30945;
assign w30947 = ~w29590 & ~w29592;
assign w30948 = (w30946 & w47860) | (w30946 & w47861) | (w47860 & w47861);
assign w30949 = w30944 & ~w30948;
assign w30950 = ~w30944 & w30948;
assign w30951 = ~w30949 & ~w30950;
assign w30952 = w29536 & w30239;
assign w30953 = ~w30239 & ~w30951;
assign w30954 = ~w30952 & ~w30953;
assign w30955 = ~w6769 & ~w30954;
assign w30956 = ~w29629 & ~w29630;
assign w30957 = ~w29631 & w30956;
assign w30958 = w29569 & w29579;
assign w30959 = (w30946 & w47862) | (w30946 & w47863) | (w47862 & w47863);
assign w30960 = ~w7924 & w30239;
assign w30961 = ~w30239 & w45864;
assign w30962 = ~w30960 & ~w30961;
assign w30963 = ~w29554 & ~w29592;
assign w30964 = w30962 & ~w30963;
assign w30965 = ~w30962 & w30963;
assign w30966 = ~w30964 & ~w30965;
assign w30967 = w7315 & ~w30966;
assign w30968 = ~w30955 & ~w30967;
assign w30969 = ~w8666 & w29579;
assign w30970 = w29569 & ~w30969;
assign w30971 = ~w30958 & w50221;
assign w30972 = ~w30970 & w30239;
assign w30973 = ~w30239 & w45865;
assign w30974 = ~w30972 & ~w30973;
assign w30975 = (w7924 & w30973) | (w7924 & w49248) | (w30973 & w49248);
assign w30976 = (w30956 & ~w30946) | (w30956 & w47864) | (~w30946 & w47864);
assign w30977 = w30976 & ~w30239;
assign w30978 = (w42462 & w45866) | (w42462 & w45867) | (w45866 & w45867);
assign w30979 = ~w30977 & ~w30978;
assign w30980 = ~w29588 & ~w29631;
assign w30981 = w8666 & w30980;
assign w30982 = (w30981 & w30977) | (w30981 & w45868) | (w30977 & w45868);
assign w30983 = w8666 & ~w30980;
assign w30984 = ~w30977 & w45869;
assign w30985 = ~w30982 & ~w30984;
assign w30986 = ~w30975 & w30985;
assign w30987 = ~w9781 & w29617;
assign w30988 = w11648 & w29605;
assign w30989 = (w30946 & w45870) | (w30946 & w45871) | (w45870 & w45871);
assign w30990 = w9781 & ~w29618;
assign w30991 = (w30946 & w45872) | (w30946 & w45873) | (w45872 & w45873);
assign w30992 = w30989 & ~w30991;
assign w30993 = (w29626 & w30239) | (w29626 & w45874) | (w30239 & w45874);
assign w30994 = (w30946 & w47865) | (w30946 & w47866) | (w47865 & w47866);
assign w30995 = ~w30239 & w45875;
assign w30996 = ~w30993 & ~w30995;
assign w30997 = ~w9195 & ~w30996;
assign w30998 = ~w11138 & w30946;
assign w30999 = w11138 & ~w30946;
assign w31000 = ~w30998 & ~w30999;
assign w31001 = ~w30148 & w31000;
assign w31002 = ~w10419 & ~w29661;
assign w31003 = w31000 & w42526;
assign w31004 = ~w30800 & w31003;
assign w31005 = ~w10419 & w29661;
assign w31006 = (w31005 & ~w31000) | (w31005 & w42527) | (~w31000 & w42527);
assign w31007 = w30237 & w31005;
assign w31008 = ~w30258 & w31007;
assign w31009 = ~w31006 & ~w31008;
assign w31010 = ~w31004 & w31009;
assign w31011 = w29616 & ~w29662;
assign w31012 = ~w29606 & ~w29618;
assign w31013 = w29616 & ~w31012;
assign w31014 = ~w29616 & w31012;
assign w31015 = ~w31013 & ~w31014;
assign w31016 = w30946 & w42528;
assign w31017 = (w31015 & ~w30946) | (w31015 & w42529) | (~w30946 & w42529);
assign w31018 = ~w31016 & ~w31017;
assign w31019 = ~w9781 & w29605;
assign w31020 = w31019 & w30239;
assign w31021 = ~w9781 & w31018;
assign w31022 = ~w30239 & w31021;
assign w31023 = ~w31020 & ~w31022;
assign w31024 = w31010 & w31023;
assign w31025 = w9781 & ~w29605;
assign w31026 = w31025 & w30239;
assign w31027 = w9781 & ~w31018;
assign w31028 = ~w30239 & w31027;
assign w31029 = ~w31026 & ~w31028;
assign w31030 = (w31029 & ~w31010) | (w31029 & w42530) | (~w31010 & w42530);
assign w31031 = ~w30997 & w31030;
assign w31032 = w9195 & w30996;
assign w31033 = ~w8666 & ~w30980;
assign w31034 = (w31033 & w30977) | (w31033 & w45876) | (w30977 & w45876);
assign w31035 = ~w8666 & w30980;
assign w31036 = ~w30977 & w45877;
assign w31037 = ~w31034 & ~w31036;
assign w31038 = ~w31032 & w31037;
assign w31039 = (w30986 & w31031) | (w30986 & w45878) | (w31031 & w45878);
assign w31040 = ~w7924 & w30974;
assign w31041 = ~w7315 & ~w30963;
assign w31042 = ~w30962 & w31041;
assign w31043 = ~w7315 & w30963;
assign w31044 = w30962 & w31043;
assign w31045 = ~w31042 & ~w31044;
assign w31046 = ~w31040 & w31045;
assign w31047 = ~w31039 & w31046;
assign w31048 = w30968 & ~w31047;
assign w31049 = ~w30929 & w42531;
assign w31050 = w10419 & w29661;
assign w31051 = w31000 & w42532;
assign w31052 = ~w30800 & w31051;
assign w31053 = w10419 & ~w29661;
assign w31054 = (w31053 & ~w31000) | (w31053 & w42533) | (~w31000 & w42533);
assign w31055 = w30237 & w31053;
assign w31056 = ~w30258 & w31055;
assign w31057 = ~w31054 & ~w31056;
assign w31058 = ~w31052 & w31057;
assign w31059 = (w31023 & ~w31058) | (w31023 & w42534) | (~w31058 & w42534);
assign w31060 = ~w30997 & ~w31059;
assign w31061 = w30986 & w31060;
assign w31062 = w31046 & ~w31061;
assign w31063 = ~w31039 & w31062;
assign w31064 = w29691 & ~w29692;
assign w31065 = ~w29691 & w29692;
assign w31066 = ~w31064 & ~w31065;
assign w31067 = ~w31066 & w30239;
assign w31068 = w29714 & ~w30183;
assign w31069 = w30176 & w31068;
assign w31070 = (~w31069 & w29634) | (~w31069 & w42535) | (w29634 & w42535);
assign w31071 = ~w29368 & ~w31069;
assign w31072 = ~w29519 & w31071;
assign w31073 = ~w31070 & ~w31072;
assign w31074 = w29676 & ~w31073;
assign w31075 = ~w29763 & ~w30176;
assign w31076 = w31068 & ~w31075;
assign w31077 = (w31076 & w31073) | (w31076 & w47867) | (w31073 & w47867);
assign w31078 = w29697 & w30193;
assign w31079 = ~w30183 & ~w31078;
assign w31080 = (w31079 & w42536) | (w31079 & w31074) | (w42536 & w31074);
assign w31081 = ~w30239 & ~w31080;
assign w31082 = w30183 & w31078;
assign w31083 = w31076 & w31078;
assign w31084 = (~w31082 & w42537) | (~w31082 & w31074) | (w42537 & w31074);
assign w31085 = w3646 & w31067;
assign w31086 = w3646 & w31084;
assign w31087 = w31081 & w31086;
assign w31088 = ~w31085 & ~w31087;
assign w31089 = ~w30176 & ~w31068;
assign w31090 = (w31089 & w29634) | (w31089 & w42538) | (w29634 & w42538);
assign w31091 = ~w29368 & w31089;
assign w31092 = ~w29519 & w31091;
assign w31093 = ~w31090 & ~w31092;
assign w31094 = ~w29763 & w31089;
assign w31095 = (~w31094 & w31093) | (~w31094 & w47868) | (w31093 & w47868);
assign w31096 = ~w30182 & w30239;
assign w31097 = ~w31077 & w31095;
assign w31098 = ~w30239 & w31097;
assign w31099 = ~w31096 & ~w31098;
assign w31100 = (~w4056 & w31098) | (~w4056 & w42539) | (w31098 & w42539);
assign w31101 = w31088 & ~w31100;
assign w31102 = ~w30156 & ~w30159;
assign w31103 = ~w29737 & w31102;
assign w31104 = ~w29717 & w31103;
assign w31105 = ~w5330 & w31104;
assign w31106 = ~w29677 & w31105;
assign w31107 = ~w30161 & w30169;
assign w31108 = (~w31107 & w29634) | (~w31107 & w42540) | (w29634 & w42540);
assign w31109 = ~w29368 & ~w31107;
assign w31110 = ~w29519 & w31109;
assign w31111 = ~w31108 & ~w31110;
assign w31112 = ~w31104 & ~w31107;
assign w31113 = (~w31112 & w31111) | (~w31112 & w47869) | (w31111 & w47869);
assign w31114 = ~w31106 & w31113;
assign w31115 = ~w30239 & w31114;
assign w31116 = w4838 & ~w29748;
assign w31117 = (w31116 & ~w31114) | (w31116 & w42541) | (~w31114 & w42541);
assign w31118 = w4838 & w29748;
assign w31119 = w31114 & w42542;
assign w31120 = ~w31117 & ~w31119;
assign w31121 = (~w30174 & w29634) | (~w30174 & w42543) | (w29634 & w42543);
assign w31122 = ~w29368 & ~w30174;
assign w31123 = ~w29519 & w31122;
assign w31124 = ~w31121 & ~w31123;
assign w31125 = ~w29717 & w29750;
assign w31126 = ~w30171 & ~w31125;
assign w31127 = ~w29637 & w30172;
assign w31128 = ~w29368 & w30172;
assign w31129 = ~w29519 & w31128;
assign w31130 = ~w31127 & ~w31129;
assign w31131 = w4838 & ~w31126;
assign w31132 = (w31131 & w31124) | (w31131 & w47870) | (w31124 & w47870);
assign w31133 = ~w4838 & w31126;
assign w31134 = (~w31133 & w31130) | (~w31133 & w47871) | (w31130 & w47871);
assign w31135 = ~w31132 & w31134;
assign w31136 = ~w30239 & w31135;
assign w31137 = ~w4430 & ~w29760;
assign w31138 = (w31137 & ~w31135) | (w31137 & w42544) | (~w31135 & w42544);
assign w31139 = ~w4430 & w29760;
assign w31140 = w31135 & w42545;
assign w31141 = ~w31138 & ~w31140;
assign w31142 = w31120 & w31141;
assign w31143 = w31101 & w31142;
assign w31144 = w29674 & ~w30238;
assign w31145 = ~w30150 & w31144;
assign w31146 = ~w29675 & ~w29717;
assign w31147 = ~w29634 & w42546;
assign w31148 = (w31147 & w29519) | (w31147 & w45879) | (w29519 & w45879);
assign w31149 = (w31146 & w29667) | (w31146 & w45880) | (w29667 & w45880);
assign w31150 = ~w29636 & w31149;
assign w31151 = ~w29667 & w45881;
assign w31152 = ~w31148 & ~w31151;
assign w31153 = ~w31150 & w31152;
assign w31154 = ~w30150 & w42547;
assign w31155 = w5745 & ~w31153;
assign w31156 = ~w30239 & w31155;
assign w31157 = ~w31154 & ~w31156;
assign w31158 = ~w29675 & ~w31103;
assign w31159 = (w31158 & w29667) | (w31158 & w45882) | (w29667 & w45882);
assign w31160 = ~w29636 & w31159;
assign w31161 = w29717 & ~w31103;
assign w31162 = ~w31160 & ~w31161;
assign w31163 = ~w29677 & w31104;
assign w31164 = w31162 & ~w31163;
assign w31165 = ~w30239 & ~w31164;
assign w31166 = ~w29736 & ~w30238;
assign w31167 = ~w30150 & w31166;
assign w31168 = (~w5330 & w30150) | (~w5330 & w42548) | (w30150 & w42548);
assign w31169 = ~w31165 & w31168;
assign w31170 = w31157 & ~w31169;
assign w31171 = ~w30239 & ~w31153;
assign w31172 = (~w5745 & w30150) | (~w5745 & w42549) | (w30150 & w42549);
assign w31173 = ~w31171 & w31172;
assign w31174 = (~w29537 & w29633) | (~w29537 & w31175) | (w29633 & w31175);
assign w31175 = (~w29537 & w29590) | (~w29537 & w42550) | (w29590 & w42550);
assign w31176 = w29664 & ~w31175;
assign w31177 = ~w29658 & w31176;
assign w31178 = w31174 & w31177;
assign w31179 = ~w29545 & ~w29638;
assign w31180 = w31174 & ~w31179;
assign w31181 = ~w31174 & w31179;
assign w31182 = ~w31180 & ~w31181;
assign w31183 = w29520 & w45883;
assign w31184 = (~w31182 & ~w29520) | (~w31182 & w45884) | (~w29520 & w45884);
assign w31185 = ~w31183 & ~w31184;
assign w31186 = w6264 & ~w29544;
assign w31187 = w31186 & w30239;
assign w31188 = w6264 & w31185;
assign w31189 = ~w30239 & w31188;
assign w31190 = ~w31187 & ~w31189;
assign w31191 = ~w31173 & w31190;
assign w31192 = w31170 & ~w31191;
assign w31193 = ~w31165 & ~w31167;
assign w31194 = (w5330 & w31165) | (w5330 & w42551) | (w31165 & w42551);
assign w31195 = ~w4838 & w29748;
assign w31196 = (w31195 & ~w31114) | (w31195 & w42552) | (~w31114 & w42552);
assign w31197 = ~w4838 & ~w29748;
assign w31198 = w31114 & w42553;
assign w31199 = ~w31196 & ~w31198;
assign w31200 = ~w31194 & w31199;
assign w31201 = ~w31192 & w31200;
assign w31202 = w31081 & w31084;
assign w31203 = ~w31067 & ~w31202;
assign w31204 = ~w3646 & w31203;
assign w31205 = ~w31098 & w42554;
assign w31206 = w4430 & w29760;
assign w31207 = (w31206 & ~w31135) | (w31206 & w42555) | (~w31135 & w42555);
assign w31208 = w4430 & ~w29760;
assign w31209 = w31135 & w42556;
assign w31210 = ~w31207 & ~w31209;
assign w31211 = ~w31205 & w31210;
assign w31212 = w31101 & ~w31211;
assign w31213 = ~w31204 & ~w31212;
assign w31214 = w31143 & ~w31201;
assign w31215 = w31213 & ~w31214;
assign w31216 = w30968 & w31215;
assign w31217 = ~w31063 & w31216;
assign w31218 = ~w1120 & w30506;
assign w31219 = w30497 & w31218;
assign w31220 = w30492 & ~w31219;
assign w31221 = w2006 & w30246;
assign w31222 = (w31221 & w29677) | (w31221 & w42557) | (w29677 & w42557);
assign w31223 = ~w30239 & ~w31222;
assign w31224 = (~w2006 & ~w30246) | (~w2006 & w47872) | (~w30246 & w47872);
assign w31225 = (w31224 & ~w29677) | (w31224 & w42558) | (~w29677 & w42558);
assign w31226 = ~w30239 & w45885;
assign w31227 = w29894 & ~w31226;
assign w31228 = ~w29894 & w31226;
assign w31229 = ~w31227 & ~w31228;
assign w31230 = w1738 & ~w31229;
assign w31231 = w29894 & ~w31225;
assign w31232 = w31223 & ~w31231;
assign w31233 = ~w29881 & ~w29896;
assign w31234 = w1541 & w31233;
assign w31235 = (w31234 & w31232) | (w31234 & w45886) | (w31232 & w45886);
assign w31236 = w1541 & ~w31233;
assign w31237 = ~w31232 & w45887;
assign w31238 = ~w31235 & ~w31237;
assign w31239 = ~w31230 & w31238;
assign w31240 = ~w1738 & w31229;
assign w31241 = ~w29808 & ~w30203;
assign w31242 = ~w30202 & w31241;
assign w31243 = ~w29675 & ~w31242;
assign w31244 = ~w29668 & w31243;
assign w31245 = ~w29636 & w31244;
assign w31246 = ~w30202 & ~w30203;
assign w31247 = ~w29764 & ~w31246;
assign w31248 = w29821 & ~w31247;
assign w31249 = (w31248 & ~w31244) | (w31248 & w47873) | (~w31244 & w47873);
assign w31250 = ~w29820 & ~w30221;
assign w31251 = ~w30225 & ~w31250;
assign w31252 = (w31251 & w31245) | (w31251 & w42559) | (w31245 & w42559);
assign w31253 = ~w2285 & w30239;
assign w31254 = ~w30239 & ~w31252;
assign w31255 = w29793 & w31254;
assign w31256 = (~w31253 & ~w31254) | (~w31253 & w47874) | (~w31254 & w47874);
assign w31257 = ~w29784 & ~w29796;
assign w31258 = w2006 & w31257;
assign w31259 = ~w31256 & w31258;
assign w31260 = w2006 & ~w31257;
assign w31261 = w31256 & w31260;
assign w31262 = ~w31259 & ~w31261;
assign w31263 = ~w31240 & ~w31262;
assign w31264 = w31239 & ~w31263;
assign w31265 = w30238 & ~w31250;
assign w31266 = w29963 & w42560;
assign w31267 = ~w29677 & w31266;
assign w31268 = ~w31265 & ~w31267;
assign w31269 = ~w31249 & ~w31268;
assign w31270 = w29793 & ~w30225;
assign w31271 = ~w2285 & ~w31270;
assign w31272 = (w31271 & w30150) | (w31271 & w42561) | (w30150 & w42561);
assign w31273 = ~w31269 & w31272;
assign w31274 = ~w2285 & w31270;
assign w31275 = (w31274 & w31245) | (w31274 & w42562) | (w31245 & w42562);
assign w31276 = ~w31268 & w31275;
assign w31277 = ~w30150 & w42563;
assign w31278 = ~w31276 & ~w31277;
assign w31279 = ~w31273 & w31278;
assign w31280 = w2285 & ~w31270;
assign w31281 = (w31280 & w31245) | (w31280 & w42564) | (w31245 & w42564);
assign w31282 = ~w31268 & w31281;
assign w31283 = ~w30150 & w42565;
assign w31284 = ~w31282 & ~w31283;
assign w31285 = w2285 & w31270;
assign w31286 = (w31285 & w30150) | (w31285 & w42566) | (w30150 & w42566);
assign w31287 = ~w31269 & w31286;
assign w31288 = w31284 & ~w31287;
assign w31289 = (~w29808 & w31246) | (~w29808 & w47875) | (w31246 & w47875);
assign w31290 = ~w30216 & ~w31289;
assign w31291 = ~w31242 & w42567;
assign w31292 = ~w29668 & w31291;
assign w31293 = ~w29636 & w31292;
assign w31294 = (~w31290 & ~w31292) | (~w31290 & w47876) | (~w31292 & w47876);
assign w31295 = ~w2896 & ~w30238;
assign w31296 = ~w30150 & w31295;
assign w31297 = ~w29820 & ~w30220;
assign w31298 = ~w2558 & w31297;
assign w31299 = (w42568 & ~w31292) | (w42568 & w47877) | (~w31292 & w47877);
assign w31300 = ~w30239 & w31299;
assign w31301 = ~w30150 & w42569;
assign w31302 = ~w31300 & ~w31301;
assign w31303 = ~w30239 & w31294;
assign w31304 = ~w2558 & ~w31297;
assign w31305 = (w31304 & w30150) | (w31304 & w42570) | (w30150 & w42570);
assign w31306 = ~w31303 & w31305;
assign w31307 = w31302 & ~w31306;
assign w31308 = w31288 & w31307;
assign w31309 = w31279 & ~w31308;
assign w31310 = w2558 & w31297;
assign w31311 = (w31310 & w30150) | (w31310 & w42571) | (w30150 & w42571);
assign w31312 = ~w31303 & w31311;
assign w31313 = w2558 & ~w31297;
assign w31314 = ~w31290 & w31313;
assign w31315 = ~w31293 & w31314;
assign w31316 = ~w30239 & w31315;
assign w31317 = ~w30150 & w42572;
assign w31318 = ~w31316 & ~w31317;
assign w31319 = ~w31312 & w31318;
assign w31320 = w31279 & w31319;
assign w31321 = w31288 & ~w31320;
assign w31322 = w29764 & w30202;
assign w31323 = ~w3242 & w31246;
assign w31324 = w3242 & ~w31246;
assign w31325 = ~w31323 & ~w31324;
assign w31326 = ~w29677 & w42573;
assign w31327 = (~w31325 & w29677) | (~w31325 & w42574) | (w29677 & w42574);
assign w31328 = ~w31326 & ~w31327;
assign w31329 = ~w30239 & ~w31328;
assign w31330 = w2896 & ~w29807;
assign w31331 = ~w31329 & w31330;
assign w31332 = w2896 & w29807;
assign w31333 = w31329 & w31332;
assign w31334 = ~w31331 & ~w31333;
assign w31335 = ~w30193 & w30198;
assign w31336 = ~w30199 & ~w31335;
assign w31337 = ~w31078 & ~w31336;
assign w31338 = w30238 & ~w31337;
assign w31339 = w29963 & w42575;
assign w31340 = ~w29677 & w31339;
assign w31341 = ~w31338 & ~w31340;
assign w31342 = ~w30183 & w30199;
assign w31343 = (w31342 & w31074) | (w31342 & w42576) | (w31074 & w42576);
assign w31344 = ~w31341 & ~w31343;
assign w31345 = w30198 & ~w31084;
assign w31346 = w29102 & ~w29701;
assign w31347 = ~w29102 & w29701;
assign w31348 = ~w31346 & ~w31347;
assign w31349 = ~w31348 & w30239;
assign w31350 = (~w31349 & ~w31344) | (~w31349 & w42577) | (~w31344 & w42577);
assign w31351 = ~w2896 & ~w29807;
assign w31352 = ~w3242 & ~w31351;
assign w31353 = w31352 & ~w30239;
assign w31354 = ~w31328 & w31353;
assign w31355 = (~w31246 & w29677) | (~w31246 & w42578) | (w29677 & w42578);
assign w31356 = ~w2896 & w29807;
assign w31357 = ~w3242 & ~w31356;
assign w31358 = (w31357 & w30239) | (w31357 & w47878) | (w30239 & w47878);
assign w31359 = ~w31354 & ~w31358;
assign w31360 = ~w31350 & ~w31359;
assign w31361 = w31334 & ~w31360;
assign w31362 = ~w31321 & ~w31361;
assign w31363 = ~w31309 & ~w31362;
assign w31364 = w31264 & w31363;
assign w31365 = w31220 & w31364;
assign w31366 = w31217 & w31365;
assign w31367 = ~w31049 & w31366;
assign w31368 = ~w1541 & ~w31233;
assign w31369 = (w31368 & w31232) | (w31368 & w45888) | (w31232 & w45888);
assign w31370 = ~w1541 & w31233;
assign w31371 = ~w31232 & w45889;
assign w31372 = ~w31369 & ~w31371;
assign w31373 = w1320 & w31372;
assign w31374 = ~w29881 & ~w29898;
assign w31375 = w31374 & ~w30239;
assign w31376 = w30211 & w30230;
assign w31377 = (w31376 & w31245) | (w31376 & w45890) | (w31245 & w45890);
assign w31378 = w31375 & ~w31377;
assign w31379 = ~w1541 & w30239;
assign w31380 = ~w29857 & ~w29882;
assign w31381 = ~w31378 & w47879;
assign w31382 = (w31380 & w31378) | (w31380 & w47880) | (w31378 & w47880);
assign w31383 = ~w31381 & ~w31382;
assign w31384 = ~w31232 & w45891;
assign w31385 = (w31233 & w31232) | (w31233 & w45892) | (w31232 & w45892);
assign w31386 = ~w31384 & ~w31385;
assign w31387 = ~w31383 & ~w31386;
assign w31388 = ~w31373 & ~w31387;
assign w31389 = ~w2006 & ~w31257;
assign w31390 = (w31389 & w31255) | (w31389 & w45893) | (w31255 & w45893);
assign w31391 = ~w2006 & w31257;
assign w31392 = ~w31255 & w45894;
assign w31393 = ~w31390 & ~w31392;
assign w31394 = ~w31240 & w31393;
assign w31395 = w31239 & ~w31394;
assign w31396 = ~w31388 & ~w31395;
assign w31397 = ~w30509 & w31396;
assign w31398 = w6769 & w30954;
assign w31399 = ~w29544 & w30239;
assign w31400 = ~w6264 & ~w31399;
assign w31401 = ~w30239 & w31185;
assign w31402 = w31400 & ~w31401;
assign w31403 = ~w31398 & ~w31402;
assign w31404 = w31170 & w31403;
assign w31405 = w31143 & w31404;
assign w31406 = w31215 & ~w31405;
assign w31407 = w3242 & w31350;
assign w31408 = ~w31329 & w31356;
assign w31409 = w31329 & w31351;
assign w31410 = ~w31408 & ~w31409;
assign w31411 = w31308 & w31334;
assign w31412 = ~w31407 & w31410;
assign w31413 = w31411 & ~w31412;
assign w31414 = ~w31321 & ~w31413;
assign w31415 = ~w31406 & w31414;
assign w31416 = w31220 & ~w31397;
assign w31417 = w31365 & ~w31415;
assign w31418 = ~w31416 & ~w31417;
assign w31419 = ~w31417 & w42580;
assign w31420 = ~w31367 & w31419;
assign w31421 = w30518 & ~w31420;
assign w31422 = ~w29856 & ~w31378;
assign w31423 = w1541 & ~w31422;
assign w31424 = w29856 & w31378;
assign w31425 = w31423 & ~w31424;
assign w31426 = w1320 & ~w31383;
assign w31427 = ~w31229 & w31425;
assign w31428 = ~w1738 & w31262;
assign w31429 = w31427 & ~w31428;
assign w31430 = w31363 & ~w31429;
assign w31431 = w31256 & ~w31257;
assign w31432 = ~w31256 & w31257;
assign w31433 = ~w31431 & ~w31432;
assign w31434 = w2339 & w31433;
assign w31435 = w31427 & ~w31434;
assign w31436 = (w31435 & w31415) | (w31435 & w42581) | (w31415 & w42581);
assign w31437 = ~w31321 & w31393;
assign w31438 = ~w31413 & w31427;
assign w31439 = (~w31429 & ~w31438) | (~w31429 & w42582) | (~w31438 & w42582);
assign w31440 = (w31393 & w31362) | (w31393 & w31461) | (w31362 & w31461);
assign w31441 = ~w31214 & w42583;
assign w31442 = ~w31440 & w31441;
assign w31443 = ~w31439 & ~w31442;
assign w31444 = (w30968 & ~w31062) | (w30968 & w45895) | (~w31062 & w45895);
assign w31445 = ~w30856 & w31047;
assign w31446 = w31444 & ~w31445;
assign w31447 = ~w31443 & w31446;
assign w31448 = w30896 & w30917;
assign w31449 = (w31448 & w30733) | (w31448 & w42584) | (w30733 & w42584);
assign w31450 = w30924 & ~w30939;
assign w31451 = ~w30827 & ~w30850;
assign w31452 = w31046 & ~w31451;
assign w31453 = ~w31039 & w31452;
assign w31454 = w31450 & w31453;
assign w31455 = ~w31449 & w31454;
assign w31456 = ~w31426 & ~w31436;
assign w31457 = ~w31426 & ~w31455;
assign w31458 = w31447 & w31457;
assign w31459 = ~w31456 & ~w31458;
assign w31460 = w31262 & w31361;
assign w31461 = w31309 & w31393;
assign w31462 = w31460 & ~w31461;
assign w31463 = w31217 & w31462;
assign w31464 = ~w31049 & w31463;
assign w31465 = w31262 & ~w31414;
assign w31466 = w31406 & w31462;
assign w31467 = ~w31465 & ~w31466;
assign w31468 = w1738 & w31393;
assign w31469 = ~w31466 & w42585;
assign w31470 = w31425 & w31469;
assign w31471 = ~w31464 & w31470;
assign w31472 = ~w31459 & ~w31471;
assign w31473 = w30517 & w31418;
assign w31474 = ~w31367 & w31473;
assign w31475 = (~w30468 & ~w31473) | (~w30468 & w42586) | (~w31473 & w42586);
assign w31476 = w31472 & w31475;
assign w31477 = (~w31421 & ~w31472) | (~w31421 & w42587) | (~w31472 & w42587);
assign w31478 = ~w31049 & w31217;
assign w31479 = ~w31425 & ~w31426;
assign w31480 = w30508 & ~w31479;
assign w31481 = w31220 & ~w31480;
assign w31482 = w31264 & ~w31414;
assign w31483 = w31397 & ~w31482;
assign w31484 = (~w31406 & w31483) | (~w31406 & w47881) | (w31483 & w47881);
assign w31485 = ~w31478 & w31484;
assign w31486 = (w31481 & ~w31483) | (w31481 & w47882) | (~w31483 & w47882);
assign w31487 = (w31486 & w31478) | (w31486 & w49249) | (w31478 & w49249);
assign w31488 = ~w30856 & w31453;
assign w31489 = w31444 & ~w31488;
assign w31490 = ~w31455 & w31489;
assign w31491 = (w31436 & ~w31490) | (w31436 & w45896) | (~w31490 & w45896);
assign w31492 = ~w30353 & ~w30513;
assign w31493 = w30510 & ~w31492;
assign w31494 = ~w31464 & w31469;
assign w31495 = (~w1320 & w31417) | (~w1320 & w42588) | (w31417 & w42588);
assign w31496 = ~w1320 & w31366;
assign w31497 = ~w31049 & w31496;
assign w31498 = ~w31495 & ~w31497;
assign w31499 = w31487 & ~w31491;
assign w31500 = ~w30509 & w31493;
assign w31501 = (w31500 & w31498) | (w31500 & w42589) | (w31498 & w42589);
assign w31502 = ~w31499 & w31501;
assign w31503 = ~w31487 & w47883;
assign w31504 = ~w31502 & ~w31503;
assign w31505 = ~w30362 & ~w31477;
assign w31506 = w31504 & w31505;
assign w31507 = ~w30456 & w31477;
assign w31508 = ~w30457 & ~w30463;
assign w31509 = ~w31477 & w31508;
assign w31510 = ~w31507 & ~w31509;
assign w31511 = w31506 & ~w31510;
assign w31512 = ~w31506 & w31510;
assign w31513 = ~w31511 & ~w31512;
assign w31514 = w3 & w31513;
assign w31515 = (~w30509 & w31498) | (~w30509 & w42590) | (w31498 & w42590);
assign w31516 = ~w31499 & w31515;
assign w31517 = (w30355 & w31487) | (w30355 & w47884) | (w31487 & w47884);
assign w31518 = w30337 & ~w31492;
assign w31519 = w30298 & w31518;
assign w31520 = w30332 & ~w31519;
assign w31521 = (~w31520 & w31516) | (~w31520 & w47885) | (w31516 & w47885);
assign w31522 = w30267 & ~w31477;
assign w31523 = w30267 & ~w30359;
assign w31524 = ~w31477 & ~w31523;
assign w31525 = w30358 & w31477;
assign w31526 = ~w31521 & w31524;
assign w31527 = ~w31525 & ~w31526;
assign w31528 = ~w30359 & w31522;
assign w31529 = w31521 & w31528;
assign w31530 = w31527 & ~w31529;
assign w31531 = w57 & ~w31530;
assign w31532 = ~w57 & ~w31421;
assign w31533 = ~w31476 & w31532;
assign w31534 = w30355 & ~w30359;
assign w31535 = (w31436 & ~w42591) | (w31436 & w45896) | (~w42591 & w45896);
assign w31536 = (~w45896 & w47886) | (~w45896 & w47887) | (w47886 & w47887);
assign w31537 = ~w30353 & w31486;
assign w31538 = ~w31485 & w31537;
assign w31539 = ~w31536 & ~w31538;
assign w31540 = w31487 & ~w31535;
assign w31541 = ~w30509 & w31519;
assign w31542 = (w31541 & w31498) | (w31541 & w42592) | (w31498 & w42592);
assign w31543 = ~w31540 & w31542;
assign w31544 = ~w31538 & w47888;
assign w31545 = ~w31543 & ~w31544;
assign w31546 = ~w31522 & ~w31533;
assign w31547 = (w31534 & w31476) | (w31534 & w42593) | (w31476 & w42593);
assign w31548 = w31545 & w31547;
assign w31549 = ~w31546 & ~w31548;
assign w31550 = w30257 & ~w30271;
assign w31551 = w31549 & ~w31550;
assign w31552 = ~w31549 & w31550;
assign w31553 = ~w31551 & ~w31552;
assign w31554 = ~w80 & w31553;
assign w31555 = ~w31531 & ~w31554;
assign w31556 = ~w3 & ~w31513;
assign w31557 = w80 & w31550;
assign w31558 = ~w31549 & w31557;
assign w31559 = w80 & ~w31550;
assign w31560 = w31549 & w31559;
assign w31561 = ~w31558 & ~w31560;
assign w31562 = ~w31556 & w31561;
assign w31563 = ~w30799 & ~w30850;
assign w31564 = ~w31449 & w31450;
assign w31565 = ~w30849 & ~w31564;
assign w31566 = ~w30824 & ~w31565;
assign w31567 = ~w30851 & ~w31566;
assign w31568 = ~w30825 & w31567;
assign w31569 = ~w30812 & ~w31568;
assign w31570 = ~w11138 & w31477;
assign w31571 = ~w31477 & w31569;
assign w31572 = ~w31570 & ~w31571;
assign w31573 = w31563 & ~w31572;
assign w31574 = ~w31563 & w31572;
assign w31575 = ~w31573 & ~w31574;
assign w31576 = w10419 & w31575;
assign w31577 = ~w30780 & w30896;
assign w31578 = ~w30937 & ~w31577;
assign w31579 = w30916 & ~w30933;
assign w31580 = w14039 & ~w31579;
assign w31581 = (w31580 & w31476) | (w31580 & w42594) | (w31476 & w42594);
assign w31582 = ~w31477 & ~w31578;
assign w31583 = w31581 & ~w31582;
assign w31584 = w14039 & w31579;
assign w31585 = ~w31476 & w42595;
assign w31586 = ~w31578 & w31584;
assign w31587 = ~w31477 & w31586;
assign w31588 = ~w31585 & ~w31587;
assign w31589 = ~w31583 & w31588;
assign w31590 = ~w30903 & ~w30918;
assign w31591 = w30938 & ~w31577;
assign w31592 = w30916 & ~w31591;
assign w31593 = w31590 & ~w31592;
assign w31594 = ~w31590 & w31592;
assign w31595 = ~w31593 & ~w31594;
assign w31596 = ~w13384 & w30902;
assign w31597 = w31477 & w31596;
assign w31598 = ~w13384 & w31595;
assign w31599 = ~w31477 & w31598;
assign w31600 = ~w31597 & ~w31599;
assign w31601 = w31589 & w31600;
assign w31602 = w30902 & w31477;
assign w31603 = ~w31477 & w31595;
assign w31604 = ~w31602 & ~w31603;
assign w31605 = w13384 & w31604;
assign w31606 = ~w30849 & w30923;
assign w31607 = ~w30918 & ~w30939;
assign w31608 = ~w31449 & w31607;
assign w31609 = w31606 & ~w31608;
assign w31610 = ~w31606 & w31608;
assign w31611 = ~w31609 & ~w31610;
assign w31612 = w30848 & w31477;
assign w31613 = ~w31477 & w31611;
assign w31614 = ~w31612 & ~w31613;
assign w31615 = ~w12666 & ~w31614;
assign w31616 = ~w31605 & ~w31615;
assign w31617 = w12666 & w31614;
assign w31618 = w12666 & ~w31565;
assign w31619 = ~w12666 & w31565;
assign w31620 = ~w31618 & ~w31619;
assign w31621 = ~w31477 & w31620;
assign w31622 = w11870 & w30823;
assign w31623 = (w31622 & w31477) | (w31622 & w47889) | (w31477 & w47889);
assign w31624 = w11870 & ~w30823;
assign w31625 = ~w31477 & w47890;
assign w31626 = ~w31623 & ~w31625;
assign w31627 = ~w31617 & w31626;
assign w31628 = w11870 & ~w31567;
assign w31629 = ~w11870 & w31567;
assign w31630 = ~w31628 & ~w31629;
assign w31631 = (w30811 & w31477) | (w30811 & w47891) | (w31477 & w47891);
assign w31632 = ~w31477 & w47892;
assign w31633 = ~w31631 & ~w31632;
assign w31634 = ~w11138 & ~w31633;
assign w31635 = w31627 & ~w31634;
assign w31636 = ~w31601 & w31616;
assign w31637 = w31635 & ~w31636;
assign w31638 = w10419 & w31477;
assign w31639 = w30943 & ~w31477;
assign w31640 = ~w31638 & ~w31639;
assign w31641 = w31010 & w31058;
assign w31642 = ~w9781 & ~w31641;
assign w31643 = w31640 & w31642;
assign w31644 = ~w9781 & w31641;
assign w31645 = ~w31640 & w31644;
assign w31646 = ~w31643 & ~w31645;
assign w31647 = ~w11870 & ~w30823;
assign w31648 = (w31647 & w31477) | (w31647 & w47893) | (w31477 & w47893);
assign w31649 = ~w11870 & w30823;
assign w31650 = ~w31477 & w47894;
assign w31651 = ~w31648 & ~w31650;
assign w31652 = w11138 & ~w30811;
assign w31653 = (w31652 & w31477) | (w31652 & w47895) | (w31477 & w47895);
assign w31654 = w11138 & w30811;
assign w31655 = ~w31477 & w47896;
assign w31656 = ~w31653 & ~w31655;
assign w31657 = w31651 & w31656;
assign w31658 = ~w31634 & ~w31657;
assign w31659 = ~w30780 & w30860;
assign w31660 = ~w16559 & w31659;
assign w31661 = w16559 & ~w31659;
assign w31662 = ~w31660 & ~w31661;
assign w31663 = ~w30468 & ~w31662;
assign w31664 = ~w31474 & w31663;
assign w31665 = w31472 & w31664;
assign w31666 = (w30877 & w31665) | (w30877 & w42596) | (w31665 & w42596);
assign w31667 = ~w31665 & w42597;
assign w31668 = ~w31666 & ~w31667;
assign w31669 = w15681 & w30877;
assign w31670 = (w31669 & w31665) | (w31669 & w42598) | (w31665 & w42598);
assign w31671 = w15681 & ~w30877;
assign w31672 = ~w31665 & w42599;
assign w31673 = ~w31670 & ~w31672;
assign w31674 = (~w30730 & w30645) | (~w30730 & w42600) | (w30645 & w42600);
assign w31675 = w30720 & w31674;
assign w31676 = ~w30751 & w30775;
assign w31677 = ~w30741 & w31676;
assign w31678 = ~w31675 & w31677;
assign w31679 = w30729 & ~w30751;
assign w31680 = ~w30857 & ~w31679;
assign w31681 = ~w31678 & w31680;
assign w31682 = w17380 & ~w31681;
assign w31683 = ~w17380 & w31681;
assign w31684 = ~w31682 & ~w31683;
assign w31685 = ~w30468 & w31684;
assign w31686 = ~w31474 & w31685;
assign w31687 = w31472 & w31686;
assign w31688 = w31421 & w31684;
assign w31689 = ~w31687 & ~w31688;
assign w31690 = ~w16559 & w30766;
assign w31691 = (w31690 & w31687) | (w31690 & w42601) | (w31687 & w42601);
assign w31692 = ~w16559 & ~w30766;
assign w31693 = ~w31687 & w42602;
assign w31694 = ~w31691 & ~w31693;
assign w31695 = ~w15681 & w31668;
assign w31696 = w31673 & ~w31694;
assign w31697 = ~w31695 & ~w31696;
assign w31698 = w16559 & ~w30766;
assign w31699 = (w31698 & w31687) | (w31698 & w42603) | (w31687 & w42603);
assign w31700 = w16559 & w30766;
assign w31701 = ~w31687 & w42604;
assign w31702 = ~w31699 & ~w31701;
assign w31703 = w31673 & w31702;
assign w31704 = ~w30893 & w31659;
assign w31705 = ~w30934 & ~w31704;
assign w31706 = ~w15681 & w31705;
assign w31707 = w15681 & ~w31705;
assign w31708 = ~w31706 & ~w31707;
assign w31709 = ~w14766 & ~w30892;
assign w31710 = (w31709 & w31477) | (w31709 & w47897) | (w31477 & w47897);
assign w31711 = ~w14766 & w30892;
assign w31712 = ~w31477 & w47898;
assign w31713 = ~w31710 & ~w31712;
assign w31714 = ~w31703 & w31713;
assign w31715 = w31697 & w31714;
assign w31716 = (w30892 & w31477) | (w30892 & w47899) | (w31477 & w47899);
assign w31717 = ~w31477 & w47900;
assign w31718 = ~w31716 & ~w31717;
assign w31719 = w14766 & ~w31718;
assign w31720 = w31576 & w31646;
assign w31721 = w31646 & ~w31719;
assign w31722 = ~w31715 & w31721;
assign w31723 = ~w31720 & ~w31722;
assign w31724 = w31646 & ~w31658;
assign w31725 = ~w31637 & w31724;
assign w31726 = w31723 & ~w31725;
assign w31727 = w11977 & ~w30798;
assign w31728 = ~w11977 & w30798;
assign w31729 = ~w31727 & ~w31728;
assign w31730 = w31572 & w31729;
assign w31731 = ~w31572 & ~w31729;
assign w31732 = ~w31730 & ~w31731;
assign w31733 = ~w31658 & w31732;
assign w31734 = ~w31637 & w31733;
assign w31735 = w31616 & w31657;
assign w31736 = ~w14766 & w31578;
assign w31737 = w14766 & ~w31578;
assign w31738 = ~w31736 & ~w31737;
assign w31739 = (w30932 & w31477) | (w30932 & w47901) | (w31477 & w47901);
assign w31740 = ~w31477 & w47902;
assign w31741 = ~w31739 & ~w31740;
assign w31742 = ~w14039 & w31600;
assign w31743 = ~w31741 & w31742;
assign w31744 = w31732 & ~w31743;
assign w31745 = w31735 & w31744;
assign w31746 = ~w31576 & ~w31745;
assign w31747 = ~w31734 & w31746;
assign w31748 = ~w31726 & ~w31747;
assign w31749 = ~w30696 & w31674;
assign w31750 = w30740 & ~w31749;
assign w31751 = ~w30706 & ~w31750;
assign w31752 = ~w20000 & w31751;
assign w31753 = w20000 & ~w31751;
assign w31754 = ~w31752 & ~w31753;
assign w31755 = w29509 & ~w30713;
assign w31756 = ~w29509 & w30713;
assign w31757 = ~w31755 & ~w31756;
assign w31758 = ~w19040 & w31757;
assign w31759 = ~w31754 & w31758;
assign w31760 = ~w31477 & w31759;
assign w31761 = ~w19040 & ~w31757;
assign w31762 = w31754 & w31761;
assign w31763 = (~w31762 & w31476) | (~w31762 & w42605) | (w31476 & w42605);
assign w31764 = ~w31760 & w31763;
assign w31765 = w30738 & ~w31749;
assign w31766 = w20906 & ~w31765;
assign w31767 = ~w20906 & w31765;
assign w31768 = ~w31766 & ~w31767;
assign w31769 = ~w20000 & w30705;
assign w31770 = ~w31768 & w31769;
assign w31771 = ~w31477 & w31770;
assign w31772 = ~w20000 & ~w30705;
assign w31773 = w31768 & w31772;
assign w31774 = (~w31773 & w31476) | (~w31773 & w42606) | (w31476 & w42606);
assign w31775 = ~w31771 & w31774;
assign w31776 = w31764 & w31775;
assign w31777 = ~w30645 & w30670;
assign w31778 = w22767 & ~w31777;
assign w31779 = ~w22767 & w31777;
assign w31780 = ~w31778 & ~w31779;
assign w31781 = ~w21801 & w31674;
assign w31782 = ~w31780 & w31781;
assign w31783 = ~w31477 & w31782;
assign w31784 = ~w21801 & w30681;
assign w31785 = w31780 & w31784;
assign w31786 = (~w31785 & w31476) | (~w31785 & w42607) | (w31476 & w42607);
assign w31787 = ~w31783 & w31786;
assign w31788 = w21801 & ~w31674;
assign w31789 = ~w31781 & ~w31788;
assign w31790 = w20906 & w30695;
assign w31791 = ~w31789 & w31790;
assign w31792 = ~w31477 & w31791;
assign w31793 = w20906 & ~w30695;
assign w31794 = w31789 & w31793;
assign w31795 = (~w31794 & w31476) | (~w31794 & w42608) | (w31476 & w42608);
assign w31796 = ~w31792 & w31795;
assign w31797 = w31787 & w31796;
assign w31798 = w31776 & w31797;
assign w31799 = (w30517 & w31498) | (w30517 & w42609) | (w31498 & w42609);
assign w31800 = ~w31499 & w31799;
assign w31801 = (w45896 & w47903) | (w45896 & w47904) | (w47903 & w47904);
assign w31802 = ~w30627 & w30644;
assign w31803 = w25851 & ~w31802;
assign w31804 = ~w25851 & w31802;
assign w31805 = ~w31803 & ~w31804;
assign w31806 = w30629 & ~w30800;
assign w31807 = w29437 & ~w31806;
assign w31808 = ~w29437 & w31806;
assign w31809 = ~w31807 & ~w31808;
assign w31810 = w31805 & ~w31809;
assign w31811 = ~w31804 & ~w31810;
assign w31812 = ~w30654 & w31811;
assign w31813 = ~w24874 & w31812;
assign w31814 = ~w30468 & w31813;
assign w31815 = (w31814 & w31487) | (w31814 & w47905) | (w31487 & w47905);
assign w31816 = w29400 & w30239;
assign w31817 = ~w30239 & w30595;
assign w31818 = ~w31816 & ~w31817;
assign w31819 = w31812 & w31818;
assign w31820 = (~w31819 & w31476) | (~w31819 & w42610) | (w31476 & w42610);
assign w31821 = ~w31800 & w31815;
assign w31822 = w31820 & ~w31821;
assign w31823 = ~w30602 & ~w30654;
assign w31824 = ~w31811 & ~w31823;
assign w31825 = (w31824 & w31476) | (w31824 & w42611) | (w31476 & w42611);
assign w31826 = w23843 & ~w31825;
assign w31827 = w31822 & w31826;
assign w31828 = w30617 & ~w30669;
assign w31829 = ~w30602 & ~w31812;
assign w31830 = w31828 & ~w31829;
assign w31831 = ~w31828 & w31829;
assign w31832 = ~w31830 & ~w31831;
assign w31833 = ~w30668 & w31477;
assign w31834 = ~w31477 & w31832;
assign w31835 = ~w31833 & ~w31834;
assign w31836 = w22767 & ~w31835;
assign w31837 = ~w31827 & ~w31836;
assign w31838 = w31798 & w31837;
assign w31839 = ~w30468 & w31810;
assign w31840 = (w31839 & ~w31473) | (w31839 & w42612) | (~w31473 & w42612);
assign w31841 = w31472 & w31840;
assign w31842 = w31421 & w31810;
assign w31843 = ~w30362 & ~w30457;
assign w31844 = ~w30362 & w47906;
assign w31845 = w30466 & ~w31844;
assign w31846 = ~w30509 & w31845;
assign w31847 = (w31846 & w31498) | (w31846 & w42613) | (w31498 & w42613);
assign w31848 = ~w31540 & w31847;
assign w31849 = ~w31487 & w31535;
assign w31850 = ~w31487 & w47907;
assign w31851 = ~w31848 & ~w31850;
assign w31852 = ~w30468 & w31805;
assign w31853 = ~w31841 & w47908;
assign w31854 = ~w31841 & w42614;
assign w31855 = w31851 & w31854;
assign w31856 = ~w31853 & ~w31855;
assign w31857 = (~w24874 & w31855) | (~w24874 & w47909) | (w31855 & w47909);
assign w31858 = w31822 & ~w31825;
assign w31859 = (~w23843 & ~w31822) | (~w23843 & w47910) | (~w31822 & w47910);
assign w31860 = ~w31857 & ~w31859;
assign w31861 = ~w22767 & w31835;
assign w31862 = ~w31477 & ~w31780;
assign w31863 = w21801 & ~w30681;
assign w31864 = (w31863 & w31477) | (w31863 & w47911) | (w31477 & w47911);
assign w31865 = w21801 & w30681;
assign w31866 = ~w31477 & w47912;
assign w31867 = ~w31864 & ~w31866;
assign w31868 = ~w31861 & w31867;
assign w31869 = ~w20906 & ~w30695;
assign w31870 = ~w31789 & w31869;
assign w31871 = ~w31477 & w31870;
assign w31872 = ~w20906 & w30695;
assign w31873 = w31789 & w31872;
assign w31874 = (~w31873 & w31476) | (~w31873 & w42615) | (w31476 & w42615);
assign w31875 = ~w31871 & w31874;
assign w31876 = w20000 & w30705;
assign w31877 = w31768 & w31876;
assign w31878 = (~w31877 & w31476) | (~w31877 & w42616) | (w31476 & w42616);
assign w31879 = w31753 & ~w31768;
assign w31880 = ~w31477 & w31879;
assign w31881 = w31878 & ~w31880;
assign w31882 = w31875 & w31881;
assign w31883 = w31776 & ~w31882;
assign w31884 = w19040 & w31757;
assign w31885 = (w31884 & w31477) | (w31884 & w47913) | (w31477 & w47913);
assign w31886 = w19040 & ~w31757;
assign w31887 = ~w31477 & w47914;
assign w31888 = ~w31885 & ~w31887;
assign w31889 = ~w30729 & ~w30769;
assign w31890 = ~w30741 & w30774;
assign w31891 = ~w31675 & w31890;
assign w31892 = w31889 & w31891;
assign w31893 = ~w30729 & ~w31892;
assign w31894 = ~w18183 & w31893;
assign w31895 = w18183 & ~w31893;
assign w31896 = ~w31894 & ~w31895;
assign w31897 = ~w17380 & w30750;
assign w31898 = ~w31896 & w31897;
assign w31899 = ~w31477 & w31898;
assign w31900 = ~w17380 & ~w30750;
assign w31901 = (w31900 & w31420) | (w31900 & w47915) | (w31420 & w47915);
assign w31902 = w31896 & w31900;
assign w31903 = (~w31902 & w31476) | (~w31902 & w42617) | (w31476 & w42617);
assign w31904 = ~w31899 & w31903;
assign w31905 = w31889 & ~w31891;
assign w31906 = ~w31889 & w31891;
assign w31907 = ~w31905 & ~w31906;
assign w31908 = w18183 & ~w30728;
assign w31909 = w31477 & w31908;
assign w31910 = w18183 & w31907;
assign w31911 = ~w31477 & w31910;
assign w31912 = ~w31909 & ~w31911;
assign w31913 = w31904 & w31912;
assign w31914 = w31888 & w31913;
assign w31915 = ~w31883 & w31914;
assign w31916 = w31798 & ~w31868;
assign w31917 = w31915 & ~w31916;
assign w31918 = w31838 & ~w31860;
assign w31919 = w31917 & ~w31918;
assign w31920 = ~a[16] & ~w30239;
assign w31921 = ~w29158 & w30239;
assign w31922 = w29158 & ~w30239;
assign w31923 = ~w31921 & ~w31922;
assign w31924 = w30520 & w31923;
assign w31925 = ~w30520 & ~w31920;
assign w31926 = ~w31923 & w31925;
assign w31927 = ~w31924 & ~w31926;
assign w31928 = w30239 & ~w30518;
assign w31929 = w31924 & ~w31928;
assign w31930 = w29158 & ~w30519;
assign w31931 = ~w30468 & ~w31930;
assign w31932 = w31920 & ~w31931;
assign w31933 = a[17] & ~w31932;
assign w31934 = ~w31929 & w31933;
assign w31935 = w31421 & w31926;
assign w31936 = w31934 & ~w31935;
assign w31937 = w31472 & w47916;
assign w31938 = w31936 & ~w31937;
assign w31939 = (w31920 & w31848) | (w31920 & w47917) | (w31848 & w47917);
assign w31940 = w31938 & ~w31939;
assign w31941 = w31515 & ~w31540;
assign w31942 = (~w31849 & ~w31515) | (~w31849 & w49250) | (~w31515 & w49250);
assign w31943 = w30520 & ~w31923;
assign w31944 = ~w30468 & w31943;
assign w31945 = ~w31941 & w47918;
assign w31946 = ~a[16] & ~w29158;
assign w31947 = w30468 & w31946;
assign w31948 = ~w30520 & w31923;
assign w31949 = ~w31947 & w31948;
assign w31950 = (w31949 & w31487) | (w31949 & w47919) | (w31487 & w47919);
assign w31951 = ~w31920 & w31927;
assign w31952 = ~a[17] & ~w31951;
assign w31953 = ~w31845 & w31944;
assign w31954 = w31952 & ~w31953;
assign w31955 = (~w31920 & w31420) | (~w31920 & w47920) | (w31420 & w47920);
assign w31956 = (w31954 & w31476) | (w31954 & w42618) | (w31476 & w42618);
assign w31957 = ~w31800 & w31950;
assign w31958 = w31956 & ~w31957;
assign w31959 = ~w31945 & w31958;
assign w31960 = ~w31940 & ~w31959;
assign w31961 = ~w31959 & w47921;
assign w31962 = a[16] & ~w30519;
assign w31963 = ~w30520 & ~w31962;
assign w31964 = ~w30468 & w31963;
assign w31965 = a[16] & w30239;
assign w31966 = ~w31920 & ~w31965;
assign w31967 = ~w30516 & w31964;
assign w31968 = (~w31967 & w31476) | (~w31967 & w42619) | (w31476 & w42619);
assign w31969 = (w31964 & w31487) | (w31964 & w47922) | (w31487 & w47922);
assign w31970 = ~w31516 & w31969;
assign w31971 = w31968 & ~w31970;
assign w31972 = ~a[15] & ~w30468;
assign w31973 = ~a[12] & ~a[13];
assign w31974 = ~a[14] & w31973;
assign w31975 = w30239 & ~w31974;
assign w31976 = ~w31845 & w31972;
assign w31977 = ~w31975 & ~w31976;
assign w31978 = (a[15] & w31420) | (a[15] & w47923) | (w31420 & w47923);
assign w31979 = (w31977 & w31476) | (w31977 & w42620) | (w31476 & w42620);
assign w31980 = (w31972 & w31487) | (w31972 & w47924) | (w31487 & w47924);
assign w31981 = ~w31516 & w31980;
assign w31982 = w31979 & ~w31981;
assign w31983 = ~w30239 & w31974;
assign w31984 = a[14] & w31972;
assign w31985 = ~w31983 & ~w31984;
assign w31986 = ~w31849 & ~w31985;
assign w31987 = ~w31845 & w31984;
assign w31988 = ~w31983 & ~w31987;
assign w31989 = (w31988 & w31941) | (w31988 & w49251) | (w31941 & w49251);
assign w31990 = ~w31982 & w31989;
assign w31991 = w29158 & w31971;
assign w31992 = ~w31990 & ~w31991;
assign w31993 = ~w29158 & ~w31971;
assign w31994 = ~w31992 & ~w31993;
assign w31995 = ~w31961 & w31994;
assign w31996 = ~w30581 & w30587;
assign w31997 = ~w30468 & w31996;
assign w31998 = (w31997 & ~w31473) | (w31997 & w42621) | (~w31473 & w42621);
assign w31999 = w31472 & w31998;
assign w32000 = w31421 & w31996;
assign w32001 = ~w31999 & ~w32000;
assign w32002 = w26880 & ~w30584;
assign w32003 = (w32002 & w31999) | (w32002 & w42622) | (w31999 & w42622);
assign w32004 = w26880 & w30584;
assign w32005 = ~w31999 & w42623;
assign w32006 = ~w32003 & ~w32005;
assign w32007 = ~w30239 & ~w30546;
assign w32008 = w30239 & w30553;
assign w32009 = ~w32007 & ~w32008;
assign w32010 = w30557 & ~w30627;
assign w32011 = ~w30584 & w30587;
assign w32012 = ~w30581 & ~w32011;
assign w32013 = w32010 & ~w32012;
assign w32014 = ~w32010 & w32012;
assign w32015 = ~w32013 & ~w32014;
assign w32016 = ~w25851 & ~w32015;
assign w32017 = ~w31477 & w32016;
assign w32018 = ~w25851 & ~w32009;
assign w32019 = w31477 & w32018;
assign w32020 = ~w32017 & ~w32019;
assign w32021 = w32006 & w32020;
assign w32022 = w24874 & w32006;
assign w32023 = w31856 & w32022;
assign w32024 = ~w32021 & ~w32023;
assign w32025 = (~w28077 & w31959) | (~w28077 & w47925) | (w31959 & w47925);
assign w32026 = ~w32024 & ~w32025;
assign w32027 = ~w31995 & w32026;
assign w32028 = ~w31855 & w47926;
assign w32029 = w31477 & w32009;
assign w32030 = ~w31477 & w32015;
assign w32031 = ~w32029 & ~w32030;
assign w32032 = w25851 & ~w32031;
assign w32033 = ~w26880 & w30584;
assign w32034 = (w32033 & w31999) | (w32033 & w42624) | (w31999 & w42624);
assign w32035 = ~w31999 & w42625;
assign w32036 = ~w32034 & ~w32035;
assign w32037 = w32020 & ~w32036;
assign w32038 = ~w32032 & ~w32037;
assign w32039 = ~w32028 & w32038;
assign w32040 = w31838 & w32039;
assign w32041 = ~w32027 & w32040;
assign w32042 = w31919 & ~w32041;
assign w32043 = ~w31637 & ~w31658;
assign w32044 = (~w30750 & w31477) | (~w30750 & w47927) | (w31477 & w47927);
assign w32045 = ~w31477 & w47928;
assign w32046 = ~w32044 & ~w32045;
assign w32047 = w17380 & w32046;
assign w32048 = w30728 & w31477;
assign w32049 = ~w31477 & ~w31907;
assign w32050 = ~w32048 & ~w32049;
assign w32051 = ~w18183 & ~w32050;
assign w32052 = w31904 & w32051;
assign w32053 = ~w32047 & ~w32052;
assign w32054 = w31697 & w31713;
assign w32055 = w32053 & w32054;
assign w32056 = ~w31576 & w32055;
assign w32057 = ~w32043 & w32056;
assign w32058 = ~w32042 & w32057;
assign w32059 = w31748 & ~w32058;
assign w32060 = w31141 & w31210;
assign w32061 = w31404 & ~w31490;
assign w32062 = w31201 & ~w32061;
assign w32063 = w31120 & ~w32062;
assign w32064 = w32060 & ~w32063;
assign w32065 = ~w32060 & w32063;
assign w32066 = ~w32064 & ~w32065;
assign w32067 = ~w29760 & ~w31136;
assign w32068 = w29760 & w31136;
assign w32069 = ~w32067 & ~w32068;
assign w32070 = ~w31477 & ~w32066;
assign w32071 = w31477 & w32069;
assign w32072 = ~w32070 & ~w32071;
assign w32073 = ~w4056 & w32072;
assign w32074 = (w31404 & w31049) | (w31404 & w47929) | (w31049 & w47929);
assign w32075 = w29748 & ~w31115;
assign w32076 = ~w29748 & w31115;
assign w32077 = ~w32075 & ~w32076;
assign w32078 = ~w32074 & ~w32077;
assign w32079 = ~w30517 & ~w32074;
assign w32080 = ~w31420 & ~w32061;
assign w32081 = (~w32080 & ~w31472) | (~w32080 & w42626) | (~w31472 & w42626);
assign w32082 = ~w4838 & ~w30468;
assign w32083 = (w32082 & w31472) | (w32082 & w42627) | (w31472 & w42627);
assign w32084 = ~w32081 & w32083;
assign w32085 = ~w31192 & ~w31194;
assign w32086 = ~w4838 & w32078;
assign w32087 = w32085 & ~w32086;
assign w32088 = (w32087 & w32084) | (w32087 & w47930) | (w32084 & w47930);
assign w32089 = w31120 & w31199;
assign w32090 = ~w32074 & w32085;
assign w32091 = ~w32089 & ~w32090;
assign w32092 = w31477 & ~w32077;
assign w32093 = ~w31477 & w32091;
assign w32094 = ~w32092 & ~w32093;
assign w32095 = ~w4430 & w32094;
assign w32096 = ~w32088 & w32095;
assign w32097 = ~w32073 & ~w32096;
assign w32098 = w4430 & w32087;
assign w32099 = (w32098 & w32084) | (w32098 & w47931) | (w32084 & w47931);
assign w32100 = ~w31169 & ~w31194;
assign w32101 = w31403 & ~w31490;
assign w32102 = (w31191 & w31490) | (w31191 & w45897) | (w31490 & w45897);
assign w32103 = w31157 & ~w32102;
assign w32104 = w32100 & ~w32103;
assign w32105 = ~w32100 & w32103;
assign w32106 = ~w32104 & ~w32105;
assign w32107 = ~w31477 & w32106;
assign w32108 = w31193 & ~w31421;
assign w32109 = ~w31476 & w32108;
assign w32110 = (~w4838 & w31476) | (~w4838 & w42628) | (w31476 & w42628);
assign w32111 = ~w32107 & w32110;
assign w32112 = w4430 & ~w32077;
assign w32113 = w31477 & w32112;
assign w32114 = w4430 & w32091;
assign w32115 = ~w31477 & w32114;
assign w32116 = ~w32113 & ~w32115;
assign w32117 = ~w32111 & w32116;
assign w32118 = ~w32099 & w32117;
assign w32119 = w31157 & ~w31173;
assign w32120 = w31190 & ~w32101;
assign w32121 = w32119 & ~w32120;
assign w32122 = ~w32119 & w32120;
assign w32123 = ~w32121 & ~w32122;
assign w32124 = ~w31145 & ~w31171;
assign w32125 = w31477 & w32124;
assign w32126 = ~w31477 & w32123;
assign w32127 = ~w32125 & ~w32126;
assign w32128 = ~w5330 & w32127;
assign w32129 = ~w32107 & ~w32109;
assign w32130 = w4838 & ~w32129;
assign w32131 = ~w32128 & ~w32130;
assign w32132 = w32118 & ~w32131;
assign w32133 = w32097 & ~w32132;
assign w32134 = w31088 & ~w31204;
assign w32135 = w31142 & w31404;
assign w32136 = w31142 & ~w31201;
assign w32137 = w31210 & ~w32136;
assign w32138 = ~w31205 & w32137;
assign w32139 = (w32138 & w31490) | (w32138 & w45898) | (w31490 & w45898);
assign w32140 = ~w31100 & ~w32139;
assign w32141 = w32134 & ~w32140;
assign w32142 = ~w32134 & w32140;
assign w32143 = ~w32141 & ~w32142;
assign w32144 = ~w31203 & w31477;
assign w32145 = ~w31477 & w32143;
assign w32146 = ~w32144 & ~w32145;
assign w32147 = ~w3242 & w32146;
assign w32148 = ~w31406 & ~w31478;
assign w32149 = ~w3242 & w32148;
assign w32150 = w3242 & ~w32148;
assign w32151 = ~w32149 & ~w32150;
assign w32152 = ~w2896 & w31350;
assign w32153 = (w32152 & w31477) | (w32152 & w47932) | (w31477 & w47932);
assign w32154 = ~w2896 & ~w31350;
assign w32155 = ~w31477 & w47933;
assign w32156 = ~w32153 & ~w32155;
assign w32157 = w32147 & w32156;
assign w32158 = w29807 & ~w31329;
assign w32159 = ~w29807 & w31329;
assign w32160 = ~w32158 & ~w32159;
assign w32161 = w31334 & w31410;
assign w32162 = ~w3242 & ~w31350;
assign w32163 = w31406 & ~w32162;
assign w32164 = ~w31407 & ~w32163;
assign w32165 = w31217 & ~w32162;
assign w32166 = ~w31049 & w32165;
assign w32167 = w32164 & ~w32166;
assign w32168 = w32161 & ~w32167;
assign w32169 = ~w32161 & w32167;
assign w32170 = ~w32168 & ~w32169;
assign w32171 = w31477 & ~w32160;
assign w32172 = ~w31477 & w32170;
assign w32173 = ~w32171 & ~w32172;
assign w32174 = ~w2558 & w32173;
assign w32175 = w2896 & ~w31350;
assign w32176 = (w32175 & w31477) | (w32175 & w47934) | (w31477 & w47934);
assign w32177 = w2896 & w31350;
assign w32178 = ~w31477 & w47935;
assign w32179 = ~w32176 & ~w32178;
assign w32180 = ~w32174 & w32179;
assign w32181 = ~w32157 & w32180;
assign w32182 = w4056 & ~w32072;
assign w32183 = ~w31100 & ~w31205;
assign w32184 = (w32137 & w31490) | (w32137 & w45899) | (w31490 & w45899);
assign w32185 = w32183 & ~w32184;
assign w32186 = (w31490 & w45900) | (w31490 & w45901) | (w45900 & w45901);
assign w32187 = ~w32185 & ~w32186;
assign w32188 = ~w31477 & ~w32187;
assign w32189 = ~w3646 & ~w32188;
assign w32190 = ~w31099 & w31477;
assign w32191 = w32189 & ~w32190;
assign w32192 = ~w32182 & ~w32191;
assign w32193 = w3646 & ~w31099;
assign w32194 = w31477 & w32193;
assign w32195 = (w3646 & w32185) | (w3646 & w45902) | (w32185 & w45902);
assign w32196 = ~w31477 & w32195;
assign w32197 = ~w32194 & ~w32196;
assign w32198 = ~w3242 & w32197;
assign w32199 = ~w32146 & ~w32198;
assign w32200 = w3242 & ~w32197;
assign w32201 = w32156 & ~w32200;
assign w32202 = ~w32199 & w32201;
assign w32203 = w31307 & w31319;
assign w32204 = (w31334 & w32166) | (w31334 & w45903) | (w32166 & w45903);
assign w32205 = w31410 & ~w32204;
assign w32206 = w32203 & w32205;
assign w32207 = ~w32203 & ~w32205;
assign w32208 = ~w31477 & w45904;
assign w32209 = ~w31296 & ~w31303;
assign w32210 = ~w31297 & w32209;
assign w32211 = w31297 & ~w32209;
assign w32212 = ~w32210 & ~w32211;
assign w32213 = w31477 & ~w32212;
assign w32214 = ~w32208 & ~w32213;
assign w32215 = w2285 & ~w32214;
assign w32216 = w2558 & ~w32173;
assign w32217 = (~w2285 & ~w31477) | (~w2285 & w45905) | (~w31477 & w45905);
assign w32218 = ~w32208 & w32217;
assign w32219 = ~w32216 & ~w32218;
assign w32220 = ~w31477 & w45906;
assign w32221 = ~w2285 & w31477;
assign w32222 = ~w32220 & ~w32221;
assign w32223 = w31279 & w31288;
assign w32224 = ~w2006 & ~w32223;
assign w32225 = ~w32222 & w32224;
assign w32226 = ~w2006 & w32223;
assign w32227 = w32222 & w32226;
assign w32228 = ~w32225 & ~w32227;
assign w32229 = ~w32215 & ~w32219;
assign w32230 = w32228 & ~w32229;
assign w32231 = w32181 & ~w32202;
assign w32232 = w32230 & ~w32231;
assign w32233 = w32181 & w32192;
assign w32234 = ~w32133 & w32233;
assign w32235 = w32232 & ~w32234;
assign w32236 = w5330 & ~w32127;
assign w32237 = w32118 & w32192;
assign w32238 = w32181 & w32237;
assign w32239 = w32237 & w45907;
assign w32240 = ~w30800 & w31001;
assign w32241 = w29661 & ~w32240;
assign w32242 = ~w29661 & w32240;
assign w32243 = ~w32241 & ~w32242;
assign w32244 = ~w30943 & w31641;
assign w32245 = w30943 & ~w31641;
assign w32246 = w31477 & ~w32243;
assign w32247 = ~w32244 & ~w32245;
assign w32248 = ~w31477 & w32247;
assign w32249 = ~w32246 & ~w32248;
assign w32250 = w9781 & w32249;
assign w32251 = w31023 & w31029;
assign w32252 = w9781 & w31477;
assign w32253 = w31010 & ~w32244;
assign w32254 = ~w31477 & w32253;
assign w32255 = ~w32252 & ~w32254;
assign w32256 = w32251 & ~w32255;
assign w32257 = ~w32251 & w32255;
assign w32258 = ~w32256 & ~w32257;
assign w32259 = ~w9195 & w32258;
assign w32260 = ~w32250 & ~w32259;
assign w32261 = w30943 & ~w31030;
assign w32262 = ~w31059 & ~w32261;
assign w32263 = ~w9195 & ~w31024;
assign w32264 = w32262 & ~w32263;
assign w32265 = ~w9195 & ~w31030;
assign w32266 = w30996 & ~w32265;
assign w32267 = ~w32264 & ~w32266;
assign w32268 = ~w30996 & w32265;
assign w32269 = ~w30996 & ~w31421;
assign w32270 = (~w32268 & w31476) | (~w32268 & w42629) | (w31476 & w42629);
assign w32271 = ~w31477 & ~w32267;
assign w32272 = w32270 & ~w32271;
assign w32273 = w30997 & ~w31059;
assign w32274 = ~w30943 & w32273;
assign w32275 = ~w31477 & w32274;
assign w32276 = w31032 & w32262;
assign w32277 = w8666 & ~w32276;
assign w32278 = ~w32275 & w32277;
assign w32279 = ~w32272 & w32278;
assign w32280 = (~w31032 & ~w31030) | (~w31032 & w45908) | (~w31030 & w45908);
assign w32281 = ~w30856 & w32280;
assign w32282 = w30940 & w32280;
assign w32283 = ~w30939 & w32282;
assign w32284 = ~w32281 & ~w32283;
assign w32285 = ~w31060 & w32280;
assign w32286 = (~w32285 & w30929) | (~w32285 & w42630) | (w30929 & w42630);
assign w32287 = w30985 & w31037;
assign w32288 = w32286 & ~w32287;
assign w32289 = ~w32286 & w32287;
assign w32290 = ~w32288 & ~w32289;
assign w32291 = w30979 & ~w30980;
assign w32292 = ~w30979 & w30980;
assign w32293 = ~w32291 & ~w32292;
assign w32294 = ~w31477 & ~w32290;
assign w32295 = w31477 & w32293;
assign w32296 = ~w32294 & ~w32295;
assign w32297 = w7924 & w32296;
assign w32298 = ~w32279 & ~w32297;
assign w32299 = ~w6264 & ~w31421;
assign w32300 = ~w31476 & w32299;
assign w32301 = ~w31398 & ~w31490;
assign w32302 = w31421 & ~w32301;
assign w32303 = ~w30468 & ~w32301;
assign w32304 = ~w31474 & w32303;
assign w32305 = w31472 & w32304;
assign w32306 = ~w32302 & ~w32305;
assign w32307 = ~w32300 & w32306;
assign w32308 = w31190 & ~w31402;
assign w32309 = ~w5745 & w32308;
assign w32310 = ~w32307 & w32309;
assign w32311 = ~w5745 & ~w32308;
assign w32312 = w32307 & w32311;
assign w32313 = ~w32310 & ~w32312;
assign w32314 = ~w30943 & w31061;
assign w32315 = w31047 & ~w32314;
assign w32316 = ~w30967 & ~w32315;
assign w32317 = ~w30955 & ~w31398;
assign w32318 = w32316 & ~w32317;
assign w32319 = ~w32316 & w32317;
assign w32320 = ~w32318 & ~w32319;
assign w32321 = ~w30954 & w31477;
assign w32322 = ~w31477 & w32320;
assign w32323 = ~w32321 & ~w32322;
assign w32324 = w6264 & ~w32323;
assign w32325 = w32313 & ~w32324;
assign w32326 = ~w30967 & w31045;
assign w32327 = ~w31039 & ~w32326;
assign w32328 = ~w31040 & w32327;
assign w32329 = ~w32314 & w32328;
assign w32330 = w31045 & ~w31421;
assign w32331 = ~w32315 & w32326;
assign w32332 = (~w32331 & w31476) | (~w32331 & w42631) | (w31476 & w42631);
assign w32333 = ~w32329 & w32332;
assign w32334 = w30966 & w31477;
assign w32335 = ~w6769 & ~w32334;
assign w32336 = ~w32333 & w32335;
assign w32337 = ~w30468 & w30985;
assign w32338 = w31037 & ~w32286;
assign w32339 = w32337 & ~w32338;
assign w32340 = ~w31474 & w32339;
assign w32341 = w31472 & w32340;
assign w32342 = w31421 & w32339;
assign w32343 = ~w32341 & ~w32342;
assign w32344 = ~w7924 & ~w31421;
assign w32345 = ~w31476 & w32344;
assign w32346 = w32343 & ~w32345;
assign w32347 = ~w30975 & ~w31040;
assign w32348 = w7315 & w32347;
assign w32349 = ~w32346 & w32348;
assign w32350 = w7315 & ~w32347;
assign w32351 = w32346 & w32350;
assign w32352 = ~w32349 & ~w32351;
assign w32353 = ~w32336 & w32352;
assign w32354 = w32325 & w32353;
assign w32355 = w32298 & w32354;
assign w32356 = w32260 & w32355;
assign w32357 = w32222 & ~w32223;
assign w32358 = ~w32222 & w32223;
assign w32359 = ~w32357 & ~w32358;
assign w32360 = ~w2006 & ~w32215;
assign w32361 = ~w32359 & ~w32360;
assign w32362 = (w31415 & w31049) | (w31415 & w45909) | (w31049 & w45909);
assign w32363 = w31363 & ~w32362;
assign w32364 = w31262 & w31393;
assign w32365 = w32363 & ~w32364;
assign w32366 = ~w32363 & w32364;
assign w32367 = ~w32365 & ~w32366;
assign w32368 = ~w31433 & w31477;
assign w32369 = ~w31477 & w32367;
assign w32370 = ~w32368 & ~w32369;
assign w32371 = w1738 & ~w32370;
assign w32372 = w2006 & ~w32214;
assign w32373 = w2285 & w32372;
assign w32374 = ~w32371 & ~w32373;
assign w32375 = ~w32361 & w32374;
assign w32376 = w32355 & w45910;
assign w32377 = w32235 & ~w32239;
assign w32378 = w32376 & ~w32377;
assign w32379 = ~w32059 & w32378;
assign w32380 = ~w31539 & ~w31941;
assign w32381 = (w31518 & w31941) | (w31518 & w45911) | (w31941 & w45911);
assign w32382 = w30326 & ~w32381;
assign w32383 = w351 & w31477;
assign w32384 = w30293 & ~w31477;
assign w32385 = ~w32382 & w32384;
assign w32386 = ~w32383 & ~w32385;
assign w32387 = ~w30285 & ~w30296;
assign w32388 = ~w30330 & w32387;
assign w32389 = w32386 & ~w32388;
assign w32390 = ~w32386 & w32388;
assign w32391 = ~w32389 & ~w32390;
assign w32392 = ~w252 & w32391;
assign w32393 = ~w7924 & ~w32296;
assign w32394 = ~w7315 & ~w32347;
assign w32395 = ~w32346 & w32394;
assign w32396 = ~w7315 & w32347;
assign w32397 = w32346 & w32396;
assign w32398 = ~w32395 & ~w32397;
assign w32399 = ~w32393 & w32398;
assign w32400 = w9195 & w32251;
assign w32401 = ~w32255 & w32400;
assign w32402 = w9195 & ~w32251;
assign w32403 = w32255 & w32402;
assign w32404 = ~w32401 & ~w32403;
assign w32405 = ~w32275 & ~w32276;
assign w32406 = ~w32272 & w32405;
assign w32407 = ~w8666 & ~w32406;
assign w32408 = w32404 & ~w32407;
assign w32409 = w32399 & w32408;
assign w32410 = ~w32298 & w32399;
assign w32411 = w6769 & w32334;
assign w32412 = w6769 & ~w32329;
assign w32413 = w32332 & w32412;
assign w32414 = ~w32411 & ~w32413;
assign w32415 = ~w6264 & ~w32414;
assign w32416 = ~w32323 & ~w32415;
assign w32417 = w6264 & w32414;
assign w32418 = w32313 & ~w32417;
assign w32419 = ~w32416 & w32418;
assign w32420 = w32307 & ~w32308;
assign w32421 = ~w32307 & w32308;
assign w32422 = ~w32420 & ~w32421;
assign w32423 = w5745 & w32422;
assign w32424 = ~w32419 & ~w32423;
assign w32425 = w32354 & ~w32410;
assign w32426 = ~w32409 & w32425;
assign w32427 = w32424 & ~w32426;
assign w32428 = ~w32235 & w32375;
assign w32429 = w32239 & w32375;
assign w32430 = ~w32427 & w32429;
assign w32431 = ~w32428 & ~w32430;
assign w32432 = ~w30316 & ~w30324;
assign w32433 = w30337 & w32432;
assign w32434 = ~w30468 & ~w31492;
assign w32435 = (w32434 & ~w31473) | (w32434 & w42632) | (~w31473 & w42632);
assign w32436 = w31472 & w32435;
assign w32437 = w31421 & ~w31492;
assign w32438 = ~w32436 & ~w32437;
assign w32439 = ~w32380 & ~w32438;
assign w32440 = w493 & w31477;
assign w32441 = ~w32439 & ~w32440;
assign w32442 = w32433 & ~w32441;
assign w32443 = ~w32433 & w32441;
assign w32444 = ~w32442 & ~w32443;
assign w32445 = ~w30480 & ~w30511;
assign w32446 = ~w30468 & w30491;
assign w32447 = (w32446 & ~w31473) | (w32446 & w42633) | (~w31473 & w42633);
assign w32448 = w31472 & w32447;
assign w32449 = w30491 & w31421;
assign w32450 = ~w32448 & ~w32449;
assign w32451 = ~w31218 & ~w31396;
assign w32452 = w31415 & ~w32451;
assign w32453 = ~w31364 & w31396;
assign w32454 = ~w31218 & ~w32453;
assign w32455 = ~w31478 & w32452;
assign w32456 = w32454 & ~w32455;
assign w32457 = (w30508 & ~w31472) | (w30508 & w42634) | (~w31472 & w42634);
assign w32458 = ~w32450 & ~w32457;
assign w32459 = (w32445 & w32458) | (w32445 & w42635) | (w32458 & w42635);
assign w32460 = ~w32458 & w42636;
assign w32461 = ~w32459 & ~w32460;
assign w32462 = w493 & ~w32461;
assign w32463 = (w400 & w32461) | (w400 & w18997) | (w32461 & w18997);
assign w32464 = w32444 & ~w32463;
assign w32465 = w612 & w31477;
assign w32466 = ~w30468 & ~w30511;
assign w32467 = (w32466 & ~w31473) | (w32466 & w42637) | (~w31473 & w42637);
assign w32468 = w31472 & w32467;
assign w32469 = ~w30511 & w31421;
assign w32470 = ~w32468 & ~w32469;
assign w32471 = ~w31942 & ~w32470;
assign w32472 = ~w30353 & ~w30512;
assign w32473 = w400 & ~w32472;
assign w32474 = ~w32471 & w45912;
assign w32475 = w400 & w32472;
assign w32476 = (w32475 & w32471) | (w32475 & w45913) | (w32471 & w45913);
assign w32477 = ~w32474 & ~w32476;
assign w32478 = ~w612 & ~w32477;
assign w32479 = ~w612 & w32461;
assign w32480 = ~w493 & ~w32472;
assign w32481 = (w32480 & ~w31477) | (w32480 & w45914) | (~w31477 & w45914);
assign w32482 = ~w32471 & w32481;
assign w32483 = ~w493 & w32472;
assign w32484 = w31477 & w45915;
assign w32485 = (w32483 & w32468) | (w32483 & w42638) | (w32468 & w42638);
assign w32486 = ~w31942 & w32485;
assign w32487 = ~w32484 & ~w32486;
assign w32488 = ~w32482 & w32487;
assign w32489 = w400 & ~w32433;
assign w32490 = (w32489 & ~w31477) | (w32489 & w45916) | (~w31477 & w45916);
assign w32491 = ~w32439 & w32490;
assign w32492 = w400 & w32433;
assign w32493 = (w32492 & w32436) | (w32492 & w42639) | (w32436 & w42639);
assign w32494 = ~w32380 & w32493;
assign w32495 = w31477 & w45917;
assign w32496 = ~w32494 & ~w32495;
assign w32497 = ~w32491 & w32496;
assign w32498 = w32488 & w32497;
assign w32499 = ~w32479 & w32498;
assign w32500 = ~w32478 & w32499;
assign w32501 = ~w32464 & ~w32500;
assign w32502 = w30293 & w30321;
assign w32503 = w400 & w31477;
assign w32504 = ~w31477 & w32432;
assign w32505 = ~w32381 & w32504;
assign w32506 = ~w32503 & ~w32505;
assign w32507 = w32502 & ~w32506;
assign w32508 = ~w32502 & w32506;
assign w32509 = ~w32507 & ~w32508;
assign w32510 = w351 & ~w32509;
assign w32511 = w493 & ~w32472;
assign w32512 = (w32511 & w32471) | (w32511 & w45918) | (w32471 & w45918);
assign w32513 = w493 & w32472;
assign w32514 = ~w32471 & w45919;
assign w32515 = ~w32512 & ~w32514;
assign w32516 = w612 & ~w32461;
assign w32517 = w32515 & ~w32516;
assign w32518 = w32477 & w32498;
assign w32519 = ~w32517 & w32518;
assign w32520 = ~w32510 & ~w32519;
assign w32521 = w30491 & w30497;
assign w32522 = ~w945 & w31477;
assign w32523 = (~w30507 & ~w31472) | (~w30507 & w42640) | (~w31472 & w42640);
assign w32524 = ~w31477 & w32523;
assign w32525 = ~w32522 & ~w32524;
assign w32526 = w32521 & ~w32525;
assign w32527 = ~w32521 & w32525;
assign w32528 = ~w32526 & ~w32527;
assign w32529 = w754 & w32528;
assign w32530 = ~w754 & ~w32528;
assign w32531 = w31394 & w31467;
assign w32532 = ~w31464 & w32531;
assign w32533 = w31239 & ~w32532;
assign w32534 = ~w31388 & ~w32533;
assign w32535 = w31476 & ~w32534;
assign w32536 = w1120 & w31477;
assign w32537 = ~w32535 & ~w32536;
assign w32538 = ~w30507 & ~w31218;
assign w32539 = (w945 & ~w32537) | (w945 & w45920) | (~w32537 & w45920);
assign w32540 = ~w32537 & w32538;
assign w32541 = w32539 & ~w32540;
assign w32542 = ~w32530 & ~w32541;
assign w32543 = ~w32529 & ~w32542;
assign w32544 = ~w1738 & w32370;
assign w32545 = ~w31230 & ~w32532;
assign w32546 = ~w31477 & ~w32545;
assign w32547 = w31428 & w32363;
assign w32548 = ~w31434 & ~w31494;
assign w32549 = ~w32547 & w32548;
assign w32550 = ~w31477 & w45921;
assign w32551 = (w31229 & w31477) | (w31229 & w45922) | (w31477 & w45922);
assign w32552 = ~w32550 & ~w32551;
assign w32553 = ~w1541 & ~w32552;
assign w32554 = ~w32544 & ~w32553;
assign w32555 = w31372 & ~w32533;
assign w32556 = ~w1320 & ~w32555;
assign w32557 = w31373 & ~w32533;
assign w32558 = ~w31477 & ~w32557;
assign w32559 = w1120 & w31383;
assign w32560 = (w32559 & ~w32558) | (w32559 & w45923) | (~w32558 & w45923);
assign w32561 = w1120 & ~w31383;
assign w32562 = w32558 & w45924;
assign w32563 = ~w32560 & ~w32562;
assign w32564 = w1541 & w31477;
assign w32565 = ~w32546 & ~w32564;
assign w32566 = w31238 & w31372;
assign w32567 = ~w1320 & ~w32566;
assign w32568 = w32565 & w32567;
assign w32569 = ~w1320 & w32566;
assign w32570 = ~w32565 & w32569;
assign w32571 = ~w32568 & ~w32570;
assign w32572 = w32563 & w32571;
assign w32573 = w32554 & w32572;
assign w32574 = ~w32543 & w32573;
assign w32575 = w32501 & w32520;
assign w32576 = w32574 & ~w32575;
assign w32577 = w32431 & w32576;
assign w32578 = w252 & ~w32391;
assign w32579 = ~w351 & w32509;
assign w32580 = ~w32578 & ~w32579;
assign w32581 = ~w32392 & ~w32580;
assign w32582 = w32431 & w42641;
assign w32583 = w1541 & w32552;
assign w32584 = w1320 & ~w32566;
assign w32585 = ~w32565 & w32584;
assign w32586 = w1320 & w32566;
assign w32587 = w32565 & w32586;
assign w32588 = ~w32585 & ~w32587;
assign w32589 = ~w32583 & w32588;
assign w32590 = w32572 & ~w32589;
assign w32591 = ~w1120 & ~w31383;
assign w32592 = (w32591 & ~w32558) | (w32591 & w45925) | (~w32558 & w45925);
assign w32593 = ~w1120 & w31383;
assign w32594 = w32558 & w45926;
assign w32595 = ~w32592 & ~w32594;
assign w32596 = ~w945 & w32538;
assign w32597 = ~w32537 & w32596;
assign w32598 = ~w945 & ~w32538;
assign w32599 = w32537 & w32598;
assign w32600 = ~w32597 & ~w32599;
assign w32601 = w32595 & w32600;
assign w32602 = ~w32529 & w32601;
assign w32603 = ~w32590 & w32602;
assign w32604 = ~w32543 & ~w32603;
assign w32605 = ~w32501 & w32604;
assign w32606 = w400 & ~w612;
assign w32607 = w32464 & ~w32606;
assign w32608 = w32520 & ~w32607;
assign w32609 = ~w32605 & w32608;
assign w32610 = w32580 & ~w32609;
assign w32611 = ~w32392 & ~w32610;
assign w32612 = ~w32379 & w32582;
assign w32613 = w32611 & ~w32612;
assign w32614 = ~w57 & w31530;
assign w32615 = ~w32612 & w45927;
assign w32616 = ~w31514 & ~w31562;
assign w32617 = ~w31514 & w31555;
assign w32618 = (w32617 & w32612) | (w32617 & w47936) | (w32612 & w47936);
assign w32619 = ~w32616 & ~w32618;
assign w32620 = ~w31531 & ~w32614;
assign w32621 = ~w31554 & w31561;
assign w32622 = w32620 & w32621;
assign w32623 = ~w31555 & w31561;
assign w32624 = ~w31514 & ~w31556;
assign w32625 = w32623 & ~w32624;
assign w32626 = ~w32623 & w32624;
assign w32627 = ~w32625 & ~w32626;
assign w32628 = ~w32612 & w47937;
assign w32629 = (w32627 & w32612) | (w32627 & w47938) | (w32612 & w47938);
assign w32630 = ~w32628 & ~w32629;
assign w32631 = w32619 & ~w32630;
assign w32632 = w42 & ~w32631;
assign w32633 = ~w30434 & ~w30462;
assign w32634 = w3 & w31477;
assign w32635 = w30463 & ~w31477;
assign w32636 = ~w32634 & ~w32635;
assign w32637 = ~w31477 & w31843;
assign w32638 = w31504 & w32637;
assign w32639 = w32636 & ~w32638;
assign w32640 = w32633 & ~w32639;
assign w32641 = ~w32633 & w32639;
assign w32642 = ~w32640 & ~w32641;
assign w32643 = ~w30434 & w31843;
assign w32644 = ~w30465 & ~w32643;
assign w32645 = (~w32644 & w31487) | (~w32644 & w45929) | (w31487 & w45929);
assign w32646 = ~w30515 & ~w32644;
assign w32647 = (~w32646 & w31516) | (~w32646 & w45930) | (w31516 & w45930);
assign w32648 = ~w30069 & ~w30401;
assign w32649 = w30392 & ~w32648;
assign w32650 = w30377 & w30379;
assign w32651 = w32649 & ~w32650;
assign w32652 = ~w30392 & w32647;
assign w32653 = ~w32647 & w32651;
assign w32654 = ~w32652 & ~w32653;
assign w32655 = ~w42 & ~w32654;
assign w32656 = w32619 & w32655;
assign w32657 = ~w32642 & ~w32656;
assign w32658 = w32619 & w32642;
assign w32659 = w42 & w32642;
assign w32660 = ~w30419 & w32649;
assign w32661 = ~w42 & w30392;
assign w32662 = w30398 & ~w32661;
assign w32663 = ~w32660 & w32662;
assign w32664 = w32647 & w32663;
assign w32665 = w30382 & ~w32662;
assign w32666 = ~w32647 & w32665;
assign w32667 = ~w32664 & ~w32666;
assign w32668 = (w32667 & ~w31513) | (w32667 & w45931) | (~w31513 & w45931);
assign w32669 = ~w32659 & w32668;
assign w32670 = w42 & ~w31513;
assign w32671 = w32669 & w32670;
assign w32672 = ~w32619 & w32671;
assign w32673 = ~w1 & ~w31513;
assign w32674 = w32659 & w32673;
assign w32675 = ~w32623 & w32674;
assign w32676 = w31561 & w32615;
assign w32677 = w32675 & ~w32676;
assign w32678 = ~w32672 & ~w32677;
assign w32679 = ~w42 & w32658;
assign w32680 = w32678 & ~w32679;
assign w32681 = ~w32632 & w32657;
assign w32682 = w32680 & ~w32681;
assign w32683 = ~w42 & w32654;
assign w32684 = ~w32642 & w32683;
assign w32685 = w31562 & ~w32684;
assign w32686 = ~w32669 & ~w32684;
assign w32687 = ~w31555 & w32685;
assign w32688 = ~w32686 & ~w32687;
assign w32689 = ~w32614 & w32685;
assign w32690 = ~w32392 & w32689;
assign w32691 = ~w32580 & w32690;
assign w32692 = w32688 & ~w32691;
assign w32693 = w32577 & w32692;
assign w32694 = ~w32379 & w32693;
assign w32695 = w32688 & ~w32690;
assign w32696 = w32609 & ~w32695;
assign w32697 = w32692 & ~w32696;
assign w32698 = (~w32697 & ~w32693) | (~w32697 & w42642) | (~w32693 & w42642);
assign w32699 = ~w31531 & w32698;
assign w32700 = ~w32615 & w32699;
assign w32701 = (w32621 & w32700) | (w32621 & w45932) | (w32700 & w45932);
assign w32702 = ~w32700 & w45933;
assign w32703 = ~w32701 & ~w32702;
assign w32704 = ~w3 & w32703;
assign w32705 = w31513 & ~w32698;
assign w32706 = w32630 & w32698;
assign w32707 = ~w32705 & ~w32706;
assign w32708 = ~w42 & w32707;
assign w32709 = ~w32704 & ~w32708;
assign w32710 = ~w32682 & ~w32709;
assign w32711 = ~w32613 & w32698;
assign w32712 = ~w57 & ~w32698;
assign w32713 = ~w32711 & ~w32712;
assign w32714 = w32620 & ~w32713;
assign w32715 = ~w32620 & w32713;
assign w32716 = ~w32714 & ~w32715;
assign w32717 = ~w80 & ~w32716;
assign w32718 = w3 & ~w32703;
assign w32719 = ~w32717 & ~w32718;
assign w32720 = ~w32682 & w32719;
assign w32721 = w351 & w32509;
assign w32722 = ~w351 & ~w32509;
assign w32723 = (~w32721 & w32694) | (~w32721 & w42643) | (w32694 & w42643);
assign w32724 = ~w32501 & w32574;
assign w32725 = ~w32430 & w42644;
assign w32726 = ~w32605 & ~w32607;
assign w32727 = ~w32725 & w32726;
assign w32728 = w32378 & w32726;
assign w32729 = ~w32059 & w32728;
assign w32730 = ~w32727 & ~w32729;
assign w32731 = ~w32519 & ~w32730;
assign w32732 = w32698 & w32731;
assign w32733 = ~w32723 & ~w32732;
assign w32734 = (~w32579 & w32694) | (~w32579 & w42645) | (w32694 & w42645);
assign w32735 = w32698 & ~w32731;
assign w32736 = ~w32734 & ~w32735;
assign w32737 = ~w32733 & ~w32736;
assign w32738 = w252 & ~w32737;
assign w32739 = ~w32379 & w32577;
assign w32740 = ~w32392 & ~w32578;
assign w32741 = ~w32579 & ~w32609;
assign w32742 = ~w32740 & ~w32741;
assign w32743 = ~w32697 & w32742;
assign w32744 = ~w32694 & w32743;
assign w32745 = ~w32579 & w32739;
assign w32746 = w32744 & ~w32745;
assign w32747 = ~w32391 & ~w32698;
assign w32748 = ~w32746 & ~w32747;
assign w32749 = ~w32392 & w32711;
assign w32750 = w32748 & ~w32749;
assign w32751 = (w57 & ~w32748) | (w57 & w42646) | (~w32748 & w42646);
assign w32752 = ~w32738 & ~w32751;
assign w32753 = ~w252 & w32737;
assign w32754 = ~w32430 & w42647;
assign w32755 = ~w612 & ~w32604;
assign w32756 = ~w32754 & w32755;
assign w32757 = w32378 & w32755;
assign w32758 = ~w32059 & w32757;
assign w32759 = ~w32756 & ~w32758;
assign w32760 = ~w32543 & w45934;
assign w32761 = ~w32430 & w42648;
assign w32762 = w612 & w32604;
assign w32763 = (w32461 & ~w32604) | (w32461 & w32479) | (~w32604 & w32479);
assign w32764 = ~w32761 & w32763;
assign w32765 = w32378 & w32763;
assign w32766 = ~w32059 & w32765;
assign w32767 = ~w32764 & ~w32766;
assign w32768 = w32759 & w32767;
assign w32769 = (w32515 & ~w32768) | (w32515 & w45935) | (~w32768 & w45935);
assign w32770 = (w32444 & w32694) | (w32444 & w42649) | (w32694 & w42649);
assign w32771 = ~w32694 & w42650;
assign w32772 = ~w32770 & ~w32771;
assign w32773 = (w32444 & w32694) | (w32444 & w42651) | (w32694 & w42651);
assign w32774 = ~w32694 & w42652;
assign w32775 = ~w32773 & ~w32774;
assign w32776 = ~w32769 & w32772;
assign w32777 = w32769 & w32775;
assign w32778 = ~w32776 & ~w32777;
assign w32779 = w351 & w32778;
assign w32780 = ~w32753 & ~w32779;
assign w32781 = w32752 & ~w32780;
assign w32782 = w80 & w32716;
assign w32783 = w32748 & w45936;
assign w32784 = ~w32782 & ~w32783;
assign w32785 = ~w351 & ~w32778;
assign w32786 = w32752 & ~w32785;
assign w32787 = w32784 & ~w32786;
assign w32788 = ~w32781 & w32787;
assign w32789 = w32720 & ~w32788;
assign w32790 = (~w32710 & w32788) | (~w32710 & w45962) | (w32788 & w45962);
assign w32791 = w493 & ~w32698;
assign w32792 = w32698 & w32768;
assign w32793 = ~w32791 & ~w32792;
assign w32794 = w32488 & w32515;
assign w32795 = ~w400 & ~w32794;
assign w32796 = ~w32793 & w32795;
assign w32797 = ~w400 & w32794;
assign w32798 = w32793 & w32797;
assign w32799 = ~w32796 & ~w32798;
assign w32800 = w612 & w32754;
assign w32801 = ~w32379 & w32800;
assign w32802 = w32759 & ~w32801;
assign w32803 = w32698 & w32802;
assign w32804 = w493 & w32461;
assign w32805 = (w32462 & ~w32803) | (w32462 & w45937) | (~w32803 & w45937);
assign w32806 = w32803 & w45938;
assign w32807 = ~w32805 & ~w32806;
assign w32808 = w32799 & w32807;
assign w32809 = ~w493 & w32461;
assign w32810 = (w32809 & ~w32803) | (w32809 & w45939) | (~w32803 & w45939);
assign w32811 = ~w493 & ~w32461;
assign w32812 = w32803 & w45940;
assign w32813 = ~w32810 & ~w32812;
assign w32814 = ~w32430 & w42653;
assign w32815 = ~w32377 & w45941;
assign w32816 = ~w32059 & w32815;
assign w32817 = (w32589 & w32430) | (w32589 & w45942) | (w32430 & w45942);
assign w32818 = ~w32816 & ~w32817;
assign w32819 = ~w32572 & w32601;
assign w32820 = ~w32541 & ~w32819;
assign w32821 = ~w32697 & w32820;
assign w32822 = ~w32694 & w32821;
assign w32823 = w32601 & ~w32818;
assign w32824 = w32822 & ~w32823;
assign w32825 = ~w32529 & ~w32530;
assign w32826 = w612 & ~w32825;
assign w32827 = (w32826 & w32824) | (w32826 & w42654) | (w32824 & w42654);
assign w32828 = w612 & w32825;
assign w32829 = ~w32824 & w42655;
assign w32830 = ~w32827 & ~w32829;
assign w32831 = w32813 & ~w32830;
assign w32832 = w32808 & ~w32831;
assign w32833 = ~w1120 & ~w32698;
assign w32834 = ~w32816 & w45943;
assign w32835 = w32698 & w32834;
assign w32836 = ~w32833 & ~w32835;
assign w32837 = w32563 & w32595;
assign w32838 = ~w945 & w32837;
assign w32839 = w32836 & w32838;
assign w32840 = ~w945 & ~w32837;
assign w32841 = ~w32836 & w32840;
assign w32842 = ~w32839 & ~w32841;
assign w32843 = w32595 & ~w32697;
assign w32844 = ~w32694 & w32843;
assign w32845 = w32572 & w32818;
assign w32846 = w32844 & ~w32845;
assign w32847 = w945 & ~w32698;
assign w32848 = ~w32846 & ~w32847;
assign w32849 = ~w32541 & w32600;
assign w32850 = w754 & w32849;
assign w32851 = (w32850 & w32846) | (w32850 & w42656) | (w32846 & w42656);
assign w32852 = w754 & ~w32849;
assign w32853 = ~w32846 & w42657;
assign w32854 = ~w32851 & ~w32853;
assign w32855 = w32842 & w32854;
assign w32856 = w945 & ~w32837;
assign w32857 = w32836 & w32856;
assign w32858 = w945 & w32837;
assign w32859 = ~w32836 & w32858;
assign w32860 = ~w32857 & ~w32859;
assign w32861 = (~w32583 & w32379) | (~w32583 & w45944) | (w32379 & w45944);
assign w32862 = w1320 & ~w32698;
assign w32863 = w32698 & ~w32861;
assign w32864 = ~w32862 & ~w32863;
assign w32865 = w32571 & w32588;
assign w32866 = ~w1120 & ~w32865;
assign w32867 = ~w32864 & w32866;
assign w32868 = ~w1120 & w32865;
assign w32869 = w32864 & w32868;
assign w32870 = ~w32867 & ~w32869;
assign w32871 = w32860 & ~w32870;
assign w32872 = w32855 & ~w32871;
assign w32873 = w32832 & w32872;
assign w32874 = w32355 & w42658;
assign w32875 = ~w31748 & w32874;
assign w32876 = w32057 & w32874;
assign w32877 = ~w32042 & w32876;
assign w32878 = ~w32875 & ~w32877;
assign w32879 = ~w32133 & w32192;
assign w32880 = (w32202 & w32133) | (w32202 & w45945) | (w32133 & w45945);
assign w32881 = w32181 & ~w32880;
assign w32882 = w32219 & ~w32881;
assign w32883 = (w32239 & w32426) | (w32239 & w45946) | (w32426 & w45946);
assign w32884 = w32882 & ~w32883;
assign w32885 = ~w32215 & w32238;
assign w32886 = ~w32878 & w32885;
assign w32887 = ~w32215 & ~w32884;
assign w32888 = (~w2006 & w32886) | (~w2006 & w45947) | (w32886 & w45947);
assign w32889 = w32698 & ~w32888;
assign w32890 = ~w32886 & w45948;
assign w32891 = w32359 & ~w32890;
assign w32892 = w32889 & ~w32891;
assign w32893 = ~w32370 & ~w32698;
assign w32894 = ~w32371 & ~w32544;
assign w32895 = w32698 & w32894;
assign w32896 = ~w32893 & ~w32895;
assign w32897 = w32892 & w32896;
assign w32898 = ~w32892 & ~w32896;
assign w32899 = ~w32897 & ~w32898;
assign w32900 = w1541 & ~w32899;
assign w32901 = ~w32430 & w45949;
assign w32902 = ~w32379 & w32901;
assign w32903 = (~w1541 & w32379) | (~w1541 & w45950) | (w32379 & w45950);
assign w32904 = w32698 & ~w32903;
assign w32905 = w1541 & w32902;
assign w32906 = w32904 & ~w32905;
assign w32907 = w1320 & w32552;
assign w32908 = (w32907 & ~w32904) | (w32907 & w45951) | (~w32904 & w45951);
assign w32909 = w1320 & ~w32552;
assign w32910 = w32904 & w45952;
assign w32911 = ~w32908 & ~w32910;
assign w32912 = w32889 & w32891;
assign w32913 = w32698 & w45953;
assign w32914 = w32889 & w45954;
assign w32915 = w1738 & ~w32359;
assign w32916 = ~w32913 & w32915;
assign w32917 = ~w32914 & ~w32916;
assign w32918 = w32911 & w32917;
assign w32919 = ~w32900 & w32918;
assign w32920 = ~w32216 & ~w32881;
assign w32921 = (~w32236 & w32426) | (~w32236 & w42659) | (w32426 & w42659);
assign w32922 = ~w32238 & w32920;
assign w32923 = w32920 & ~w32921;
assign w32924 = (~w32922 & ~w32878) | (~w32922 & w45955) | (~w32878 & w45955);
assign w32925 = ~w32215 & ~w32218;
assign w32926 = w32924 & ~w32925;
assign w32927 = ~w32924 & w32925;
assign w32928 = ~w32926 & ~w32927;
assign w32929 = w32214 & ~w32698;
assign w32930 = w32698 & ~w32928;
assign w32931 = ~w32929 & ~w32930;
assign w32932 = ~w2006 & ~w32931;
assign w32933 = (~w2285 & w32698) | (~w2285 & w45956) | (w32698 & w45956);
assign w32934 = w2006 & w32698;
assign w32935 = w32928 & w32934;
assign w32936 = w32933 & ~w32935;
assign w32937 = (w32237 & ~w32878) | (w32237 & w45957) | (~w32878 & w45957);
assign w32938 = w32880 & ~w32937;
assign w32939 = ~w32157 & ~w32938;
assign w32940 = ~w32174 & ~w32216;
assign w32941 = (w32940 & w32698) | (w32940 & w45958) | (w32698 & w45958);
assign w32942 = w32179 & w32698;
assign w32943 = w32939 & w32942;
assign w32944 = w32941 & ~w32943;
assign w32945 = w32936 & w32944;
assign w32946 = ~w32932 & ~w32945;
assign w32947 = w32179 & ~w32940;
assign w32948 = w32216 & ~w32698;
assign w32949 = w32698 & w32947;
assign w32950 = w32939 & w32949;
assign w32951 = ~w32948 & ~w32950;
assign w32952 = w32936 & ~w32951;
assign w32953 = ~w1738 & w32359;
assign w32954 = ~w32913 & w32953;
assign w32955 = ~w1738 & ~w32359;
assign w32956 = w32913 & w32955;
assign w32957 = ~w32954 & ~w32956;
assign w32958 = ~w32952 & w32957;
assign w32959 = w32946 & w32958;
assign w32960 = w32552 & ~w32906;
assign w32961 = ~w32552 & w32906;
assign w32962 = ~w32960 & ~w32961;
assign w32963 = ~w1320 & w32962;
assign w32964 = ~w1541 & w32899;
assign w32965 = w32899 & w45959;
assign w32966 = ~w32963 & ~w32965;
assign w32967 = w32919 & ~w32959;
assign w32968 = w32966 & ~w32967;
assign w32969 = w1120 & ~w32865;
assign w32970 = w32864 & w32969;
assign w32971 = w1120 & w32865;
assign w32972 = ~w32864 & w32971;
assign w32973 = ~w32970 & ~w32972;
assign w32974 = w32860 & w32973;
assign w32975 = ~w754 & w50222;
assign w32976 = w32848 & ~w32849;
assign w32977 = w32975 & ~w32976;
assign w32978 = w32855 & ~w32974;
assign w32979 = ~w32977 & ~w32978;
assign w32980 = ~w32793 & ~w32794;
assign w32981 = w400 & ~w32980;
assign w32982 = w32793 & w32794;
assign w32983 = w32981 & ~w32982;
assign w32984 = ~w32824 & w42660;
assign w32985 = (w32825 & w32824) | (w32825 & w42661) | (w32824 & w42661);
assign w32986 = ~w32984 & ~w32985;
assign w32987 = ~w612 & ~w32986;
assign w32988 = (w32813 & w32986) | (w32813 & w45961) | (w32986 & w45961);
assign w32989 = w32808 & ~w32988;
assign w32990 = ~w32983 & ~w32989;
assign w32991 = w32832 & ~w32979;
assign w32992 = w32990 & ~w32991;
assign w32993 = w32873 & ~w32968;
assign w32994 = w32992 & ~w32993;
assign w32995 = ~w32781 & w32784;
assign w32996 = (~w32710 & w32995) | (~w32710 & w45962) | (w32995 & w45962);
assign w32997 = ~w32994 & w32996;
assign w32998 = (~w32790 & w32994) | (~w32790 & w47939) | (w32994 & w47939);
assign w32999 = ~w29158 & w31990;
assign w33000 = w29158 & ~w31990;
assign w33001 = ~w32999 & ~w33000;
assign w33002 = (w31971 & w32694) | (w31971 & w42662) | (w32694 & w42662);
assign w33003 = ~w32694 & w42663;
assign w33004 = ~w33002 & ~w33003;
assign w33005 = w28077 & w33004;
assign w33006 = ~w30239 & ~w31477;
assign w33007 = w30239 & ~w31973;
assign w33008 = w31974 & w33006;
assign w33009 = ~w33007 & ~w33008;
assign w33010 = w32696 & w33009;
assign w33011 = ~w32739 & w33010;
assign w33012 = ~a[14] & ~w31477;
assign w33013 = (w33009 & w32691) | (w33009 & w45963) | (w32691 & w45963);
assign w33014 = w33012 & ~w33013;
assign w33015 = (w33014 & w32739) | (w33014 & w45964) | (w32739 & w45964);
assign w33016 = ~w31975 & ~w31983;
assign w33017 = w31477 & ~w33016;
assign w33018 = ~w33006 & ~w33012;
assign w33019 = ~w33017 & w33018;
assign w33020 = ~a[15] & ~w29158;
assign w33021 = (w33020 & w32694) | (w33020 & w42664) | (w32694 & w42664);
assign w33022 = ~w33015 & w33021;
assign w33023 = a[15] & ~w29158;
assign w33024 = w33014 & w33023;
assign w33025 = ~w33011 & w33024;
assign w33026 = ~w32694 & w42665;
assign w33027 = ~w33025 & ~w33026;
assign w33028 = ~w33022 & w33027;
assign w33029 = ~w33005 & w33028;
assign w33030 = ~w28077 & w31971;
assign w33031 = (w33030 & w32694) | (w33030 & w42666) | (w32694 & w42666);
assign w33032 = ~w28077 & ~w31971;
assign w33033 = ~w32694 & w42667;
assign w33034 = ~w33031 & ~w33033;
assign w33035 = ~w31961 & ~w32025;
assign w33036 = w31994 & ~w33035;
assign w33037 = ~w31994 & w33035;
assign w33038 = ~w33036 & ~w33037;
assign w33039 = w26880 & ~w31960;
assign w33040 = ~w32698 & w33039;
assign w33041 = w26880 & ~w33038;
assign w33042 = w32698 & w33041;
assign w33043 = ~w33040 & ~w33042;
assign w33044 = w33034 & w33043;
assign w33045 = ~a[10] & ~a[11];
assign w33046 = ~a[12] & w33045;
assign w33047 = w31477 & ~w33046;
assign w33048 = ~a[13] & ~w33047;
assign w33049 = ~w31477 & w33046;
assign w33050 = ~w33048 & ~w33049;
assign w33051 = ~w31477 & w33045;
assign w33052 = a[13] & w33047;
assign w33053 = ~w31973 & ~w33052;
assign w33054 = ~w33051 & ~w33053;
assign w33055 = w30239 & w33050;
assign w33056 = ~w32698 & w33055;
assign w33057 = w30239 & w33054;
assign w33058 = w32698 & w33057;
assign w33059 = ~w33056 & ~w33058;
assign w33060 = a[14] & w31477;
assign w33061 = a[14] & ~w31973;
assign w33062 = ~w31974 & ~w33061;
assign w33063 = ~w33012 & ~w33060;
assign w33064 = ~w32698 & w33063;
assign w33065 = w32698 & w33062;
assign w33066 = ~w33064 & ~w33065;
assign w33067 = (~w30239 & w32698) | (~w30239 & w45965) | (w32698 & w45965);
assign w33068 = w32698 & w33054;
assign w33069 = w33067 & ~w33068;
assign w33070 = w33059 & ~w33066;
assign w33071 = ~w33069 & ~w33070;
assign w33072 = a[15] & w29158;
assign w33073 = (w33072 & w32694) | (w33072 & w42668) | (w32694 & w42668);
assign w33074 = ~w33015 & w33073;
assign w33075 = ~a[15] & w29158;
assign w33076 = w33014 & w33075;
assign w33077 = ~w33011 & w33076;
assign w33078 = ~w32694 & w42669;
assign w33079 = ~w33077 & ~w33078;
assign w33080 = ~w33074 & w33079;
assign w33081 = ~w33029 & w33044;
assign w33082 = w33044 & w33080;
assign w33083 = ~w33071 & w33082;
assign w33084 = ~w33081 & ~w33083;
assign w33085 = ~w31995 & ~w32025;
assign w33086 = w26880 & ~w33085;
assign w33087 = ~w31995 & w45966;
assign w33088 = ~w33086 & ~w33087;
assign w33089 = w30584 & ~w32001;
assign w33090 = ~w30584 & w32001;
assign w33091 = ~w33089 & ~w33090;
assign w33092 = w32698 & w47940;
assign w33093 = (w33091 & ~w32698) | (w33091 & w47941) | (~w32698 & w47941);
assign w33094 = ~w33092 & ~w33093;
assign w33095 = w25851 & w33094;
assign w33096 = w31960 & ~w32698;
assign w33097 = w32698 & w33038;
assign w33098 = ~w33096 & ~w33097;
assign w33099 = ~w26880 & ~w33098;
assign w33100 = ~w33095 & ~w33099;
assign w33101 = w33084 & w33100;
assign w33102 = ~w33087 & w33091;
assign w33103 = ~w33086 & ~w33102;
assign w33104 = w25851 & ~w33103;
assign w33105 = ~w25851 & w33103;
assign w33106 = ~w33104 & ~w33105;
assign w33107 = (w32031 & ~w32698) | (w32031 & w45967) | (~w32698 & w45967);
assign w33108 = w32698 & w45968;
assign w33109 = ~w33107 & ~w33108;
assign w33110 = ~w24874 & ~w33109;
assign w33111 = ~w31857 & ~w32028;
assign w33112 = ~w32020 & ~w33111;
assign w33113 = w32032 & w33111;
assign w33114 = ~w33112 & ~w33113;
assign w33115 = w32020 & w33111;
assign w33116 = w33103 & w33115;
assign w33117 = ~w32032 & ~w33111;
assign w33118 = ~w33103 & w33117;
assign w33119 = ~w33116 & ~w33118;
assign w33120 = w33114 & w33119;
assign w33121 = ~w23843 & ~w31856;
assign w33122 = ~w32698 & w33121;
assign w33123 = ~w23843 & ~w33120;
assign w33124 = w32698 & w33123;
assign w33125 = ~w33122 & ~w33124;
assign w33126 = ~w33110 & w33125;
assign w33127 = w31856 & ~w32698;
assign w33128 = w32698 & w33120;
assign w33129 = ~w33127 & ~w33128;
assign w33130 = w23843 & ~w33129;
assign w33131 = ~w32027 & w32039;
assign w33132 = ~w31857 & ~w33131;
assign w33133 = w23843 & ~w33132;
assign w33134 = ~w23843 & w33132;
assign w33135 = ~w33133 & ~w33134;
assign w33136 = w32698 & ~w33135;
assign w33137 = w22767 & ~w31858;
assign w33138 = w32698 & w45969;
assign w33139 = w22767 & w31858;
assign w33140 = (w33139 & ~w32698) | (w33139 & w45970) | (~w32698 & w45970);
assign w33141 = ~w33138 & ~w33140;
assign w33142 = ~w33130 & w33141;
assign w33143 = ~w33126 & w33142;
assign w33144 = ~w25851 & ~w33094;
assign w33145 = w30681 & ~w31862;
assign w33146 = ~w30681 & w31862;
assign w33147 = ~w33145 & ~w33146;
assign w33148 = w31787 & w31867;
assign w33149 = ~w31827 & w32039;
assign w33150 = ~w32027 & w33149;
assign w33151 = ~w31827 & ~w31860;
assign w33152 = ~w33150 & ~w33151;
assign w33153 = ~w31861 & w33152;
assign w33154 = ~w31836 & ~w33153;
assign w33155 = w33148 & ~w33154;
assign w33156 = ~w33148 & w33154;
assign w33157 = ~w33155 & ~w33156;
assign w33158 = ~w32698 & w33147;
assign w33159 = w32698 & ~w33157;
assign w33160 = ~w33158 & ~w33159;
assign w33161 = ~w20906 & ~w33160;
assign w33162 = ~w31477 & ~w31789;
assign w33163 = w30695 & ~w33162;
assign w33164 = ~w30695 & w33162;
assign w33165 = ~w33163 & ~w33164;
assign w33166 = w31796 & w31875;
assign w33167 = w31836 & w31867;
assign w33168 = w31868 & ~w33151;
assign w33169 = (w33168 & w32027) | (w33168 & w47942) | (w32027 & w47942);
assign w33170 = ~w33167 & ~w33169;
assign w33171 = w31787 & w33170;
assign w33172 = w33166 & ~w33171;
assign w33173 = ~w33166 & w33171;
assign w33174 = ~w33172 & ~w33173;
assign w33175 = ~w32698 & ~w33165;
assign w33176 = w32698 & ~w33174;
assign w33177 = ~w33175 & ~w33176;
assign w33178 = w20000 & ~w33177;
assign w33179 = ~w33161 & ~w33178;
assign w33180 = ~w23843 & w31477;
assign w33181 = ~w31477 & w31829;
assign w33182 = ~w33180 & ~w33181;
assign w33183 = w31828 & ~w33182;
assign w33184 = ~w31828 & w33182;
assign w33185 = ~w33183 & ~w33184;
assign w33186 = ~w31836 & ~w31861;
assign w33187 = w33152 & ~w33186;
assign w33188 = ~w33152 & w33186;
assign w33189 = ~w33187 & ~w33188;
assign w33190 = ~w32698 & ~w33185;
assign w33191 = w32698 & ~w33189;
assign w33192 = ~w33190 & ~w33191;
assign w33193 = w21801 & w33192;
assign w33194 = ~w22767 & ~w31858;
assign w33195 = (w33194 & ~w32698) | (w33194 & w45971) | (~w32698 & w45971);
assign w33196 = ~w22767 & w31858;
assign w33197 = w32698 & w45972;
assign w33198 = ~w33195 & ~w33197;
assign w33199 = ~w33193 & w33198;
assign w33200 = w33179 & w33199;
assign w33201 = ~w33144 & w33200;
assign w33202 = ~w33143 & w33201;
assign w33203 = ~w33101 & w33202;
assign w33204 = w24874 & w33125;
assign w33205 = w33109 & w33204;
assign w33206 = w33142 & ~w33205;
assign w33207 = ~w20000 & w33177;
assign w33208 = ~w21801 & ~w33192;
assign w33209 = w20906 & w33160;
assign w33210 = ~w33208 & ~w33209;
assign w33211 = w33179 & ~w33210;
assign w33212 = ~w33207 & ~w33211;
assign w33213 = w33200 & ~w33206;
assign w33214 = w33212 & ~w33213;
assign w33215 = w31764 & w31888;
assign w33216 = w31775 & w31881;
assign w33217 = ~w31875 & w33216;
assign w33218 = w31797 & w33216;
assign w33219 = w33170 & w33218;
assign w33220 = ~w33217 & ~w33219;
assign w33221 = w31881 & w33220;
assign w33222 = w33215 & ~w33221;
assign w33223 = ~w33215 & w33221;
assign w33224 = ~w33222 & ~w33223;
assign w33225 = ~w19040 & w31764;
assign w33226 = w31888 & ~w33225;
assign w33227 = (~w18183 & w32698) | (~w18183 & w47943) | (w32698 & w47943);
assign w33228 = w32698 & w33224;
assign w33229 = w33227 & ~w33228;
assign w33230 = w31912 & ~w32051;
assign w33231 = ~w31883 & w31888;
assign w33232 = w31798 & ~w33167;
assign w33233 = (w33232 & w33150) | (w33232 & w45973) | (w33150 & w45973);
assign w33234 = w33231 & ~w33233;
assign w33235 = ~w33230 & ~w33234;
assign w33236 = w33230 & w33231;
assign w33237 = ~w33233 & w33236;
assign w33238 = ~w33235 & ~w33237;
assign w33239 = w17380 & w33238;
assign w33240 = ~w17380 & ~w33238;
assign w33241 = w17380 & ~w32050;
assign w33242 = ~w17380 & w32050;
assign w33243 = ~w33241 & ~w33242;
assign w33244 = ~w32698 & w33243;
assign w33245 = w32698 & w47944;
assign w33246 = ~w33244 & ~w33245;
assign w33247 = ~w33229 & ~w33246;
assign w33248 = w32050 & ~w32698;
assign w33249 = w32698 & ~w33238;
assign w33250 = ~w33248 & ~w33249;
assign w33251 = ~w17380 & ~w33250;
assign w33252 = w31904 & ~w32047;
assign w33253 = ~w32051 & ~w33237;
assign w33254 = w33252 & ~w33253;
assign w33255 = ~w33252 & w33253;
assign w33256 = ~w33254 & ~w33255;
assign w33257 = w32046 & ~w32698;
assign w33258 = w32698 & w33256;
assign w33259 = ~w33257 & ~w33258;
assign w33260 = w16559 & w33259;
assign w33261 = w30766 & ~w31689;
assign w33262 = ~w30766 & w31689;
assign w33263 = ~w33261 & ~w33262;
assign w33264 = ~w31919 & w32053;
assign w33265 = w32040 & w32053;
assign w33266 = ~w32027 & w33265;
assign w33267 = ~w33264 & ~w33266;
assign w33268 = w31694 & w31702;
assign w33269 = w33267 & w33268;
assign w33270 = ~w33267 & ~w33268;
assign w33271 = ~w32698 & ~w33263;
assign w33272 = ~w33269 & ~w33270;
assign w33273 = w32698 & w33272;
assign w33274 = ~w33271 & ~w33273;
assign w33275 = w15681 & w33274;
assign w33276 = ~w33251 & ~w33260;
assign w33277 = ~w33275 & w33276;
assign w33278 = w33276 & w47945;
assign w33279 = w31797 & w33170;
assign w33280 = w31875 & ~w33216;
assign w33281 = ~w33279 & w33280;
assign w33282 = w33220 & ~w33281;
assign w33283 = ~w31477 & ~w31768;
assign w33284 = w30705 & ~w33283;
assign w33285 = ~w30705 & w33283;
assign w33286 = ~w33284 & ~w33285;
assign w33287 = w32698 & ~w33282;
assign w33288 = ~w32698 & w33286;
assign w33289 = ~w33287 & ~w33288;
assign w33290 = ~w19040 & ~w33289;
assign w33291 = ~w15681 & ~w33274;
assign w33292 = ~w16559 & ~w33259;
assign w33293 = ~w33291 & ~w33292;
assign w33294 = ~w33275 & ~w33293;
assign w33295 = (~w33290 & w33293) | (~w33290 & w45974) | (w33293 & w45974);
assign w33296 = ~w33278 & w33295;
assign w33297 = w33214 & w33296;
assign w33298 = ~w33203 & w33297;
assign w33299 = w19040 & w33289;
assign w33300 = (w18183 & w32698) | (w18183 & w47946) | (w32698 & w47946);
assign w33301 = w32698 & ~w33224;
assign w33302 = w33300 & ~w33301;
assign w33303 = ~w33299 & ~w33302;
assign w33304 = w33247 & ~w33303;
assign w33305 = w33277 & ~w33304;
assign w33306 = ~w33294 & ~w33305;
assign w33307 = ~w31919 & w32055;
assign w33308 = w32040 & w32055;
assign w33309 = ~w32027 & w33308;
assign w33310 = ~w33307 & ~w33309;
assign w33311 = ~w31715 & ~w31719;
assign w33312 = ~w14039 & ~w31741;
assign w33313 = w33311 & ~w33312;
assign w33314 = w33310 & w33313;
assign w33315 = w31589 & ~w33314;
assign w33316 = w31600 & ~w31605;
assign w33317 = w33315 & ~w33316;
assign w33318 = ~w33315 & w33316;
assign w33319 = ~w33317 & ~w33318;
assign w33320 = w31604 & ~w32698;
assign w33321 = w32698 & ~w33319;
assign w33322 = ~w33320 & ~w33321;
assign w33323 = ~w12666 & ~w33322;
assign w33324 = w12666 & w33322;
assign w33325 = w33310 & w33311;
assign w33326 = w31589 & ~w33312;
assign w33327 = w33325 & ~w33326;
assign w33328 = ~w33325 & w33326;
assign w33329 = ~w33327 & ~w33328;
assign w33330 = ~w14039 & w31741;
assign w33331 = w31589 & ~w33330;
assign w33332 = w32698 & w33329;
assign w33333 = ~w32698 & w33331;
assign w33334 = ~w33332 & ~w33333;
assign w33335 = ~w13384 & w33334;
assign w33336 = ~w33324 & ~w33335;
assign w33337 = ~w15681 & w31694;
assign w33338 = w15681 & ~w31694;
assign w33339 = ~w33337 & ~w33338;
assign w33340 = w33267 & w45975;
assign w33341 = (~w33339 & ~w33267) | (~w33339 & w45976) | (~w33267 & w45976);
assign w33342 = ~w33340 & ~w33341;
assign w33343 = (~w31668 & w32694) | (~w31668 & w42670) | (w32694 & w42670);
assign w33344 = w31668 & w32520;
assign w33345 = ~w32695 & w33344;
assign w33346 = ~w33342 & w33345;
assign w33347 = ~w32730 & w33346;
assign w33348 = (w31668 & w32691) | (w31668 & w45977) | (w32691 & w45977);
assign w33349 = ~w33342 & w33348;
assign w33350 = (~w33349 & w32730) | (~w33349 & w45978) | (w32730 & w45978);
assign w33351 = ~w33343 & w33350;
assign w33352 = (w31697 & ~w33267) | (w31697 & w45979) | (~w33267 & w45979);
assign w33353 = w31713 & ~w31719;
assign w33354 = ~w33352 & ~w33353;
assign w33355 = ~w31719 & ~w33325;
assign w33356 = ~w33354 & ~w33355;
assign w33357 = w14039 & w31718;
assign w33358 = ~w32698 & w33357;
assign w33359 = w14039 & ~w33356;
assign w33360 = w32698 & w33359;
assign w33361 = ~w33358 & ~w33360;
assign w33362 = ~w33351 & w33361;
assign w33363 = w14766 & w33362;
assign w33364 = w13384 & w33329;
assign w33365 = w32698 & w33364;
assign w33366 = w13384 & w33331;
assign w33367 = ~w32698 & w33366;
assign w33368 = ~w33365 & ~w33367;
assign w33369 = ~w14039 & ~w31718;
assign w33370 = ~w32698 & w33369;
assign w33371 = ~w14039 & w33356;
assign w33372 = w32698 & w33371;
assign w33373 = ~w33370 & ~w33372;
assign w33374 = w33368 & w33373;
assign w33375 = ~w33323 & ~w33336;
assign w33376 = ~w33323 & w33374;
assign w33377 = ~w33363 & w33376;
assign w33378 = ~w33375 & ~w33377;
assign w33379 = ~w31616 & ~w31617;
assign w33380 = w31601 & ~w31617;
assign w33381 = (w33380 & ~w33310) | (w33380 & w45980) | (~w33310 & w45980);
assign w33382 = ~w33379 & ~w33381;
assign w33383 = w11870 & ~w33382;
assign w33384 = ~w11870 & w33382;
assign w33385 = ~w33383 & ~w33384;
assign w33386 = w30823 & ~w31621;
assign w33387 = ~w30823 & w31621;
assign w33388 = ~w33386 & ~w33387;
assign w33389 = w32698 & w45981;
assign w33390 = (w33388 & ~w32698) | (w33388 & w45982) | (~w32698 & w45982);
assign w33391 = ~w33389 & ~w33390;
assign w33392 = w11138 & ~w33391;
assign w33393 = ~w31615 & ~w31617;
assign w33394 = (w31601 & ~w33310) | (w31601 & w45983) | (~w33310 & w45983);
assign w33395 = ~w31605 & ~w33394;
assign w33396 = w33393 & ~w33395;
assign w33397 = ~w33393 & w33395;
assign w33398 = ~w33396 & ~w33397;
assign w33399 = w31614 & ~w32698;
assign w33400 = w32698 & ~w33398;
assign w33401 = ~w33399 & ~w33400;
assign w33402 = ~w11870 & w33401;
assign w33403 = ~w33392 & ~w33402;
assign w33404 = ~w33378 & w33403;
assign w33405 = ~w33306 & w33404;
assign w33406 = ~w33298 & w33405;
assign w33407 = ~w31748 & w32260;
assign w33408 = w32057 & w32260;
assign w33409 = ~w32042 & w33408;
assign w33410 = ~w33407 & ~w33409;
assign w33411 = w32352 & ~w32410;
assign w33412 = ~w32336 & w33411;
assign w33413 = (w33412 & ~w33410) | (w33412 & w45984) | (~w33410 & w45984);
assign w33414 = ~w6264 & w33413;
assign w33415 = w32416 & ~w33414;
assign w33416 = w32417 & ~w33413;
assign w33417 = w32698 & ~w33416;
assign w33418 = ~w33415 & w33417;
assign w33419 = (w32422 & ~w32698) | (w32422 & w45985) | (~w32698 & w45985);
assign w33420 = w32698 & w45986;
assign w33421 = ~w33419 & ~w33420;
assign w33422 = w33418 & ~w33421;
assign w33423 = ~w33418 & w33421;
assign w33424 = ~w33422 & ~w33423;
assign w33425 = w5330 & ~w33424;
assign w33426 = w33415 & w33417;
assign w33427 = (w32323 & ~w33417) | (w32323 & w45987) | (~w33417 & w45987);
assign w33428 = ~w33426 & ~w33427;
assign w33429 = ~w5745 & w33428;
assign w33430 = (w33411 & ~w33410) | (w33411 & w45988) | (~w33410 & w45988);
assign w33431 = ~w32336 & w32414;
assign w33432 = ~w33430 & w33431;
assign w33433 = w33430 & ~w33431;
assign w33434 = w32698 & w45989;
assign w33435 = ~w32333 & ~w32334;
assign w33436 = ~w32698 & w33435;
assign w33437 = ~w33434 & ~w33436;
assign w33438 = w6264 & ~w33437;
assign w33439 = w32352 & w32398;
assign w33440 = ~w32298 & ~w32393;
assign w33441 = ~w32393 & w32408;
assign w33442 = (~w33440 & ~w33410) | (~w33440 & w45990) | (~w33410 & w45990);
assign w33443 = w33439 & w33442;
assign w33444 = ~w33439 & ~w33442;
assign w33445 = ~w7315 & w32398;
assign w33446 = w32352 & ~w33445;
assign w33447 = ~w32698 & w33446;
assign w33448 = w32698 & w45991;
assign w33449 = ~w33447 & ~w33448;
assign w33450 = ~w6769 & w33449;
assign w33451 = ~w33438 & ~w33450;
assign w33452 = ~w33429 & w33451;
assign w33453 = ~w33425 & w33452;
assign w33454 = ~w14766 & ~w33349;
assign w33455 = ~w33347 & w33454;
assign w33456 = ~w33343 & w33455;
assign w33457 = w33361 & ~w33456;
assign w33458 = w33374 & ~w33457;
assign w33459 = w33336 & ~w33458;
assign w33460 = w33403 & ~w33459;
assign w33461 = ~w33378 & w33460;
assign w33462 = ~w32059 & ~w32250;
assign w33463 = w9195 & ~w32698;
assign w33464 = w32698 & w33462;
assign w33465 = ~w33463 & ~w33464;
assign w33466 = ~w32259 & w32404;
assign w33467 = w8666 & ~w33466;
assign w33468 = w33465 & w33467;
assign w33469 = w8666 & w33466;
assign w33470 = ~w33465 & w33469;
assign w33471 = ~w33468 & ~w33470;
assign w33472 = w8666 & ~w32406;
assign w33473 = (~w33472 & ~w33410) | (~w33472 & w45992) | (~w33410 & w45992);
assign w33474 = w32408 & w33410;
assign w33475 = ~w33473 & ~w33474;
assign w33476 = w32698 & w33475;
assign w33477 = w33410 & w45993;
assign w33478 = (~w8666 & ~w33410) | (~w8666 & w45994) | (~w33410 & w45994);
assign w33479 = ~w33477 & ~w33478;
assign w33480 = w32698 & w33479;
assign w33481 = ~w32406 & ~w33477;
assign w33482 = w32698 & w45995;
assign w33483 = w7924 & ~w33481;
assign w33484 = ~w33480 & w33483;
assign w33485 = ~w33482 & ~w33484;
assign w33486 = ~w32279 & w32408;
assign w33487 = w7924 & ~w32279;
assign w33488 = ~w7924 & w32279;
assign w33489 = ~w33487 & ~w33488;
assign w33490 = w33410 & w45996;
assign w33491 = (w33489 & ~w33410) | (w33489 & w45997) | (~w33410 & w45997);
assign w33492 = ~w33490 & ~w33491;
assign w33493 = w7315 & w32296;
assign w33494 = (w33493 & ~w32698) | (w33493 & w45998) | (~w32698 & w45998);
assign w33495 = w7315 & ~w32296;
assign w33496 = w32698 & w45999;
assign w33497 = ~w33494 & ~w33496;
assign w33498 = w33485 & w33497;
assign w33499 = w33471 & w33498;
assign w33500 = w11870 & ~w33401;
assign w33501 = ~w11138 & ~w33388;
assign w33502 = (w33501 & ~w32698) | (w33501 & w46000) | (~w32698 & w46000);
assign w33503 = ~w11138 & w33388;
assign w33504 = w32698 & w46001;
assign w33505 = ~w33502 & ~w33504;
assign w33506 = ~w33500 & w33505;
assign w33507 = ~w33392 & ~w33506;
assign w33508 = (~w31576 & w31637) | (~w31576 & w47947) | (w31637 & w47947);
assign w33509 = w31745 & w33311;
assign w33510 = w33508 & w33509;
assign w33511 = w33310 & w33510;
assign w33512 = w31646 & ~w32250;
assign w33513 = ~w31734 & w46002;
assign w33514 = (w33512 & w31734) | (w33512 & w46003) | (w31734 & w46003);
assign w33515 = ~w33513 & ~w33514;
assign w33516 = w33310 & w47948;
assign w33517 = ~w33511 & ~w33515;
assign w33518 = ~w33516 & ~w33517;
assign w33519 = ~w32697 & w33518;
assign w33520 = ~w32694 & w33519;
assign w33521 = ~w9195 & w32249;
assign w33522 = ~w32698 & w33521;
assign w33523 = ~w32694 & w42671;
assign w33524 = ~w33522 & ~w33523;
assign w33525 = w31735 & ~w31743;
assign w33526 = w33310 & w46004;
assign w33527 = w33310 & w33509;
assign w33528 = ~w31734 & ~w33527;
assign w33529 = ~w31732 & ~w32043;
assign w33530 = ~w33526 & w33529;
assign w33531 = w33528 & ~w33530;
assign w33532 = w9781 & w31575;
assign w33533 = ~w32698 & w33532;
assign w33534 = w9781 & w33531;
assign w33535 = w32698 & w33534;
assign w33536 = ~w33533 & ~w33535;
assign w33537 = w33524 & w33536;
assign w33538 = ~w31634 & w31656;
assign w33539 = ~w31627 & w31651;
assign w33540 = w31601 & ~w33539;
assign w33541 = w31626 & w33379;
assign w33542 = w31651 & ~w33541;
assign w33543 = (w33540 & ~w33310) | (w33540 & w46005) | (~w33310 & w46005);
assign w33544 = w33542 & ~w33543;
assign w33545 = w33538 & ~w33544;
assign w33546 = ~w33538 & w33544;
assign w33547 = ~w33545 & ~w33546;
assign w33548 = w32698 & ~w33547;
assign w33549 = ~w31633 & ~w32698;
assign w33550 = ~w33548 & ~w33549;
assign w33551 = w10419 & ~w33550;
assign w33552 = w33537 & ~w33551;
assign w33553 = ~w33507 & w33552;
assign w33554 = w33499 & w33553;
assign w33555 = ~w33461 & w33554;
assign w33556 = w33453 & w33555;
assign w33557 = ~w33406 & w33556;
assign w33558 = ~w32200 & w32698;
assign w33559 = ~w32199 & ~w32879;
assign w33560 = ~w32937 & w33559;
assign w33561 = ~w32147 & ~w33560;
assign w33562 = w33558 & ~w33561;
assign w33563 = w32156 & w32179;
assign w33564 = ~w33562 & w46006;
assign w33565 = (w33563 & w33562) | (w33563 & w46007) | (w33562 & w46007);
assign w33566 = ~w33564 & ~w33565;
assign w33567 = w2558 & ~w33566;
assign w33568 = w32131 & ~w32921;
assign w33569 = w32097 & ~w32118;
assign w33570 = (~w33569 & ~w32878) | (~w33569 & w46008) | (~w32878 & w46008);
assign w33571 = (~w32878 & w50386) | (~w32878 & w50387) | (w50386 & w50387);
assign w33572 = ~w32198 & ~w33571;
assign w33573 = w32698 & w47949;
assign w33574 = w32698 & w46009;
assign w33575 = ~w33573 & ~w33574;
assign w33576 = (~w46010 & w47950) | (~w46010 & w47951) | (w47950 & w47951);
assign w33577 = w32146 & w33575;
assign w33578 = w33576 & ~w33577;
assign w33579 = ~w33567 & ~w33578;
assign w33580 = w32072 & ~w32698;
assign w33581 = w32698 & w46011;
assign w33582 = ~w33580 & ~w33581;
assign w33583 = w32878 & w33568;
assign w33584 = w32118 & ~w33583;
assign w33585 = ~w32073 & ~w32182;
assign w33586 = w32698 & ~w33585;
assign w33587 = ~w32096 & ~w33584;
assign w33588 = w33586 & ~w33587;
assign w33589 = w33582 & ~w33588;
assign w33590 = w3646 & ~w33589;
assign w33591 = w3646 & ~w32698;
assign w33592 = w32698 & w46012;
assign w33593 = ~w33591 & ~w33592;
assign w33594 = ~w32191 & w32197;
assign w33595 = w3242 & ~w33594;
assign w33596 = ~w33593 & w33595;
assign w33597 = w3242 & w33594;
assign w33598 = w33593 & w33597;
assign w33599 = ~w33596 & ~w33598;
assign w33600 = ~w33590 & w33599;
assign w33601 = ~w4430 & ~w32111;
assign w33602 = (w33601 & ~w32878) | (w33601 & w46013) | (~w32878 & w46013);
assign w33603 = w4430 & w32111;
assign w33604 = (~w33603 & ~w32878) | (~w33603 & w46014) | (~w32878 & w46014);
assign w33605 = ~w33602 & w33604;
assign w33606 = ~w32088 & w32094;
assign w33607 = w32698 & w46015;
assign w33608 = (w33606 & ~w32698) | (w33606 & w46016) | (~w32698 & w46016);
assign w33609 = ~w33607 & ~w33608;
assign w33610 = w4056 & w33609;
assign w33611 = (~w3646 & ~w33586) | (~w3646 & w46017) | (~w33586 & w46017);
assign w33612 = w33582 & w33611;
assign w33613 = ~w33610 & ~w33612;
assign w33614 = w32878 & w46018;
assign w33615 = ~w32111 & ~w32130;
assign w33616 = ~w33614 & w33615;
assign w33617 = w32698 & ~w33616;
assign w33618 = w33614 & ~w33615;
assign w33619 = ~w32698 & w46019;
assign w33620 = ~w4430 & ~w33618;
assign w33621 = w33617 & w33620;
assign w33622 = ~w33619 & ~w33621;
assign w33623 = ~w4056 & ~w33606;
assign w33624 = w32698 & w46020;
assign w33625 = ~w4056 & w33606;
assign w33626 = (w33625 & ~w32698) | (w33625 & w46021) | (~w32698 & w46021);
assign w33627 = ~w33624 & ~w33626;
assign w33628 = w33622 & w33627;
assign w33629 = w33613 & ~w33628;
assign w33630 = w33600 & ~w33629;
assign w33631 = w33579 & w33630;
assign w33632 = ~w10419 & w31633;
assign w33633 = (~w33632 & w32694) | (~w33632 & w42672) | (w32694 & w42672);
assign w33634 = ~w33548 & ~w33633;
assign w33635 = ~w9781 & ~w31575;
assign w33636 = ~w32698 & w33635;
assign w33637 = ~w9781 & ~w33531;
assign w33638 = w32698 & w33637;
assign w33639 = ~w33636 & ~w33638;
assign w33640 = ~w33634 & w33639;
assign w33641 = w33537 & ~w33640;
assign w33642 = ~w8666 & ~w33466;
assign w33643 = ~w33465 & w33642;
assign w33644 = (w9195 & w32694) | (w9195 & w42673) | (w32694 & w42673);
assign w33645 = w32249 & ~w32698;
assign w33646 = w33644 & ~w33645;
assign w33647 = ~w8666 & w33466;
assign w33648 = ~w33462 & w33647;
assign w33649 = w32698 & w33648;
assign w33650 = ~w9195 & w33647;
assign w33651 = ~w32698 & w33650;
assign w33652 = ~w33649 & ~w33651;
assign w33653 = ~w33646 & w33652;
assign w33654 = ~w33643 & w33653;
assign w33655 = ~w33641 & w33654;
assign w33656 = w33499 & ~w33655;
assign w33657 = (~w33481 & ~w32698) | (~w33481 & w46022) | (~w32698 & w46022);
assign w33658 = (~w7924 & ~w32698) | (~w7924 & w46023) | (~w32698 & w46023);
assign w33659 = ~w33657 & w33658;
assign w33660 = ~w7315 & w32296;
assign w33661 = ~w33495 & ~w33660;
assign w33662 = w32698 & w46024;
assign w33663 = (w33661 & ~w32698) | (w33661 & w46025) | (~w32698 & w46025);
assign w33664 = ~w33662 & ~w33663;
assign w33665 = ~w33659 & w33664;
assign w33666 = w33497 & ~w33665;
assign w33667 = w6769 & ~w33449;
assign w33668 = ~w33666 & ~w33667;
assign w33669 = ~w33656 & w33668;
assign w33670 = ~w33434 & w42674;
assign w33671 = w33417 & w46026;
assign w33672 = w5745 & w32323;
assign w33673 = (w33672 & ~w33417) | (w33672 & w46027) | (~w33417 & w46027);
assign w33674 = ~w33671 & ~w33673;
assign w33675 = ~w33670 & w33674;
assign w33676 = ~w33429 & ~w33675;
assign w33677 = w32356 & w32427;
assign w33678 = ~w32059 & w33677;
assign w33679 = ~w32128 & ~w32236;
assign w33680 = w32427 & ~w33679;
assign w33681 = ~w32427 & w33679;
assign w33682 = ~w33680 & ~w33681;
assign w33683 = ~w32059 & w42675;
assign w33684 = ~w33678 & ~w33682;
assign w33685 = ~w33683 & ~w33684;
assign w33686 = w32127 & ~w32698;
assign w33687 = w32698 & w33685;
assign w33688 = ~w33686 & ~w33687;
assign w33689 = w4838 & ~w33688;
assign w33690 = ~w5330 & w33424;
assign w33691 = (~w33689 & ~w33424) | (~w33689 & w42676) | (~w33424 & w42676);
assign w33692 = ~w33425 & w33676;
assign w33693 = w33691 & ~w33692;
assign w33694 = w33453 & ~w33669;
assign w33695 = w33693 & ~w33694;
assign w33696 = ~w33694 & w46028;
assign w33697 = (w33696 & w33406) | (w33696 & w46029) | (w33406 & w46029);
assign w33698 = ~w2558 & w33566;
assign w33699 = ~w4838 & w33688;
assign w33700 = w32698 & w46030;
assign w33701 = (w4430 & w32698) | (w4430 & w42677) | (w32698 & w42677);
assign w33702 = ~w33700 & w33701;
assign w33703 = ~w33699 & ~w33702;
assign w33704 = w33628 & ~w33703;
assign w33705 = w33613 & ~w33704;
assign w33706 = w33600 & ~w33705;
assign w33707 = ~w3242 & w33594;
assign w33708 = (w33707 & w33592) | (w33707 & w42678) | (w33592 & w42678);
assign w33709 = ~w3242 & ~w33594;
assign w33710 = ~w33592 & w42679;
assign w33711 = ~w33708 & ~w33710;
assign w33712 = w2896 & ~w32146;
assign w33713 = (w33712 & w33573) | (w33712 & w46031) | (w33573 & w46031);
assign w33714 = w2896 & w32146;
assign w33715 = ~w33573 & w46032;
assign w33716 = ~w33713 & ~w33715;
assign w33717 = w33711 & w33716;
assign w33718 = ~w33579 & ~w33698;
assign w33719 = ~w33698 & w33717;
assign w33720 = ~w33706 & w33719;
assign w33721 = ~w33718 & ~w33720;
assign w33722 = ~w32944 & w32951;
assign w33723 = w2285 & w33722;
assign w33724 = w2006 & w32931;
assign w33725 = (~w33724 & ~w33722) | (~w33724 & w46033) | (~w33722 & w46033);
assign w33726 = w32919 & w33725;
assign w33727 = w32873 & w33726;
assign w33728 = ~w33721 & w33727;
assign w33729 = w32996 & w33728;
assign w33730 = ~w33697 & w33729;
assign w33731 = w32998 & ~w33730;
assign w33732 = w32864 & ~w32865;
assign w33733 = ~w32864 & w32865;
assign w33734 = ~w33732 & ~w33733;
assign w33735 = ~w33730 & w42680;
assign w33736 = (w33726 & w33720) | (w33726 & w47952) | (w33720 & w47952);
assign w33737 = w32968 & ~w33736;
assign w33738 = w33695 & w42681;
assign w33739 = ~w33557 & w33738;
assign w33740 = (~w33737 & w33557) | (~w33737 & w47953) | (w33557 & w47953);
assign w33741 = w32870 & w32973;
assign w33742 = (~w33741 & w33739) | (~w33741 & w42682) | (w33739 & w42682);
assign w33743 = ~w33731 & ~w33742;
assign w33744 = w33740 & w33741;
assign w33745 = w33743 & ~w33744;
assign w33746 = (~w33735 & ~w33743) | (~w33735 & w42683) | (~w33743 & w42683);
assign w33747 = ~w32682 & w32707;
assign w33748 = w32786 & w32994;
assign w33749 = (w33728 & w33557) | (w33728 & w42684) | (w33557 & w42684);
assign w33750 = w33748 & ~w33749;
assign w33751 = (w32995 & w33749) | (w32995 & w46034) | (w33749 & w46034);
assign w33752 = (~w32717 & w33730) | (~w32717 & w42685) | (w33730 & w42685);
assign w33753 = ~w33751 & w33752;
assign w33754 = ~w33730 & w47954;
assign w33755 = ~w32704 & ~w32718;
assign w33756 = ~w33753 & w47955;
assign w33757 = (w33755 & w33753) | (w33755 & w47956) | (w33753 & w47956);
assign w33758 = ~w33756 & ~w33757;
assign w33759 = ~w42 & w33758;
assign w33760 = (w33749 & w49701) | (w33749 & w49702) | (w49701 & w49702);
assign w33761 = w32707 & ~w33760;
assign w33762 = ~w32707 & w33760;
assign w33763 = ~w33761 & ~w33762;
assign w33764 = ~w33747 & w33763;
assign w33765 = w33759 & ~w33764;
assign w33766 = ~w32717 & ~w32782;
assign w33767 = ~w32781 & ~w32783;
assign w33768 = ~w33731 & ~w33750;
assign w33769 = w33767 & w33768;
assign w33770 = (w33766 & w33769) | (w33766 & w47959) | (w33769 & w47959);
assign w33771 = ~w33769 & w47960;
assign w33772 = ~w33770 & ~w33771;
assign w33773 = ~w3 & ~w33772;
assign w33774 = w42 & ~w33758;
assign w33775 = w42 & ~w32707;
assign w33776 = ~w32657 & w32707;
assign w33777 = ~w42 & ~w32658;
assign w33778 = w33776 & w33777;
assign w33779 = ~w33775 & ~w33778;
assign w33780 = w33760 & ~w33779;
assign w33781 = ~w33747 & w33779;
assign w33782 = ~w33760 & w33781;
assign w33783 = ~w33780 & ~w33782;
assign w33784 = (w33783 & w33758) | (w33783 & w49703) | (w33758 & w49703);
assign w33785 = w3 & w33772;
assign w33786 = w33784 & ~w33785;
assign w33787 = w32750 & w33731;
assign w33788 = w32830 & w32872;
assign w33789 = (w42686 & w33557) | (w42686 & w47961) | (w33557 & w47961);
assign w33790 = ~w32738 & ~w32785;
assign w33791 = (w32830 & w32978) | (w32830 & w46035) | (w32978 & w46035);
assign w33792 = w32988 & ~w33791;
assign w33793 = ~w33791 & w49704;
assign w33794 = ~w32808 & ~w32983;
assign w33795 = ~w32779 & ~w33794;
assign w33796 = w33790 & ~w33795;
assign w33797 = ~w32753 & ~w33796;
assign w33798 = w33790 & w33793;
assign w33799 = w33797 & w52272;
assign w33800 = ~w32751 & ~w32783;
assign w33801 = ~w33799 & w33800;
assign w33802 = ~w33731 & ~w33801;
assign w33803 = w33799 & ~w33800;
assign w33804 = (~w33787 & ~w33802) | (~w33787 & w49705) | (~w33802 & w49705);
assign w33805 = ~w57 & ~w33731;
assign w33806 = w80 & ~w33805;
assign w33807 = ~w32832 & ~w32983;
assign w33808 = ~w32779 & ~w33807;
assign w33809 = (w42687 & w33557) | (w42687 & w47962) | (w33557 & w47962);
assign w33810 = ~w33739 & w46037;
assign w33811 = ~w33793 & w33808;
assign w33812 = ~w32785 & ~w33811;
assign w33813 = (w33812 & w33730) | (w33812 & w42688) | (w33730 & w42688);
assign w33814 = ~w33810 & w33813;
assign w33815 = ~w32738 & ~w32753;
assign w33816 = ~w57 & ~w33815;
assign w33817 = (w33816 & w33814) | (w33816 & w46038) | (w33814 & w46038);
assign w33818 = ~w57 & w33815;
assign w33819 = ~w33814 & w46039;
assign w33820 = ~w33817 & ~w33819;
assign w33821 = w32750 & ~w33799;
assign w33822 = (~w32750 & w33730) | (~w32750 & w47963) | (w33730 & w47963);
assign w33823 = w33799 & w33822;
assign w33824 = ~w33821 & ~w33823;
assign w33825 = ~w80 & w33824;
assign w33826 = ~w33820 & ~w33825;
assign w33827 = ~w57 & w32737;
assign w33828 = w33787 & w33827;
assign w33829 = ~w57 & w80;
assign w33830 = ~w33824 & w33829;
assign w33831 = ~w33828 & ~w33830;
assign w33832 = ~w33826 & w33831;
assign w33833 = ~w33804 & w33806;
assign w33834 = w33832 & ~w33833;
assign w33835 = ~w33789 & w33792;
assign w33836 = ~w32779 & ~w32785;
assign w33837 = ~w32983 & ~w33836;
assign w33838 = (w33837 & w33730) | (w33837 & w49706) | (w33730 & w49706);
assign w33839 = (w32808 & w33789) | (w32808 & w49707) | (w33789 & w49707);
assign w33840 = w33838 & ~w33839;
assign w33841 = (w351 & w33730) | (w351 & w47964) | (w33730 & w47964);
assign w33842 = ~w32778 & ~w33841;
assign w33843 = ~w33814 & ~w33842;
assign w33844 = ~w33840 & ~w33843;
assign w33845 = ~w33843 & w49708;
assign w33846 = ~w33814 & w46040;
assign w33847 = (w33815 & w33814) | (w33815 & w46041) | (w33814 & w46041);
assign w33848 = ~w33846 & ~w33847;
assign w33849 = w57 & ~w33848;
assign w33850 = ~w33845 & ~w33849;
assign w33851 = ~w80 & w33804;
assign w33852 = w33850 & ~w33851;
assign w33853 = w33834 & ~w33852;
assign w33854 = (w33786 & ~w33853) | (w33786 & w49709) | (~w33853 & w49709);
assign w33855 = ~w33765 & ~w33854;
assign w33856 = a[12] & ~w33045;
assign w33857 = ~w33046 & ~w33856;
assign w33858 = ~a[12] & w32698;
assign w33859 = a[12] & ~w32698;
assign w33860 = ~w33858 & ~w33859;
assign w33861 = ~w31477 & w33857;
assign w33862 = (w33861 & w33730) | (w33861 & w42689) | (w33730 & w42689);
assign w33863 = ~w31477 & w33860;
assign w33864 = ~w33730 & w42690;
assign w33865 = ~w33862 & ~w33864;
assign w33866 = ~a[8] & ~a[9];
assign w33867 = ~a[10] & w33866;
assign w33868 = ~w32698 & ~w33867;
assign w33869 = w32698 & w33867;
assign w33870 = a[11] & w33868;
assign w33871 = ~w33045 & ~w33870;
assign w33872 = ~w33869 & ~w33871;
assign w33873 = (~w33872 & w33730) | (~w33872 & w42691) | (w33730 & w42691);
assign w33874 = ~a[11] & ~w33868;
assign w33875 = ~w33730 & w42692;
assign w33876 = ~w33873 & ~w33875;
assign w33877 = w31477 & ~w33860;
assign w33878 = w31477 & ~w33857;
assign w33879 = ~w30239 & ~w33878;
assign w33880 = (w33879 & w33730) | (w33879 & w42693) | (w33730 & w42693);
assign w33881 = ~w30239 & ~w33877;
assign w33882 = ~w33730 & w42694;
assign w33883 = ~w33880 & ~w33882;
assign w33884 = ~w30239 & ~w33865;
assign w33885 = ~w33876 & ~w33883;
assign w33886 = ~w33884 & ~w33885;
assign w33887 = ~w31477 & w32698;
assign w33888 = w31477 & ~w32698;
assign w33889 = ~w33887 & ~w33888;
assign w33890 = w33046 & ~w33889;
assign w33891 = a[13] & ~w33890;
assign w33892 = a[13] & ~w32698;
assign w33893 = ~w33730 & w42695;
assign w33894 = ~w33891 & ~w33893;
assign w33895 = ~w33730 & w42696;
assign w33896 = ~w33046 & w33889;
assign w33897 = (~w33896 & w33730) | (~w33896 & w42697) | (w33730 & w42697);
assign w33898 = ~w33895 & ~w33897;
assign w33899 = ~w33047 & ~w33051;
assign w33900 = w32698 & w33899;
assign w33901 = (~w42698 & w46042) | (~w42698 & w46043) | (w46042 & w46043);
assign w33902 = ~w32790 & w33858;
assign w33903 = ~w33890 & ~w33896;
assign w33904 = ~w33902 & w33903;
assign w33905 = ~a[13] & ~w33904;
assign w33906 = ~w33895 & ~w33901;
assign w33907 = w33905 & w33906;
assign w33908 = ~w33894 & ~w33898;
assign w33909 = ~w33907 & ~w33908;
assign w33910 = w33886 & ~w33909;
assign w33911 = w33059 & ~w33069;
assign w33912 = (w33911 & w33730) | (w33911 & w42699) | (w33730 & w42699);
assign w33913 = w33066 & ~w33912;
assign w33914 = ~w33066 & w33912;
assign w33915 = ~w33913 & ~w33914;
assign w33916 = w29158 & ~w33915;
assign w33917 = ~w33730 & w42700;
assign w33918 = (w33878 & w33730) | (w33878 & w42701) | (w33730 & w42701);
assign w33919 = ~w33917 & ~w33918;
assign w33920 = w30239 & w33865;
assign w33921 = ~w33876 & w33919;
assign w33922 = w33920 & ~w33921;
assign w33923 = ~w33916 & ~w33922;
assign w33924 = ~w33910 & w33923;
assign w33925 = ~w33005 & w33034;
assign w33926 = w33028 & w33080;
assign w33927 = ~w33071 & w33926;
assign w33928 = w33028 & ~w33927;
assign w33929 = w33925 & ~w33928;
assign w33930 = ~w33925 & w33928;
assign w33931 = ~w33929 & ~w33930;
assign w33932 = ~w33730 & w42702;
assign w33933 = (~w33931 & w33730) | (~w33931 & w42703) | (w33730 & w42703);
assign w33934 = ~w33932 & ~w33933;
assign w33935 = ~w26880 & w33934;
assign w33936 = w26880 & ~w33934;
assign w33937 = ~w29158 & w33926;
assign w33938 = ~w32997 & w42704;
assign w33939 = (~w33927 & w32997) | (~w33927 & w42705) | (w32997 & w42705);
assign w33940 = w33728 & w46044;
assign w33941 = ~w33697 & w33940;
assign w33942 = ~w33939 & ~w33941;
assign w33943 = ~w33730 & w33938;
assign w33944 = w33942 & ~w33943;
assign w33945 = w33071 & ~w33926;
assign w33946 = (w33945 & w32997) | (w33945 & w42706) | (w32997 & w42706);
assign w33947 = w33728 & w46045;
assign w33948 = ~w33697 & w33947;
assign w33949 = ~w33946 & ~w33948;
assign w33950 = ~w32997 & w42707;
assign w33951 = ~w33730 & w33950;
assign w33952 = w33949 & ~w33951;
assign w33953 = ~w33944 & w33952;
assign w33954 = ~w28077 & ~w33953;
assign w33955 = ~w33936 & ~w33954;
assign w33956 = w28077 & w33953;
assign w33957 = ~w29158 & ~w33066;
assign w33958 = ~w33912 & w33957;
assign w33959 = ~w29158 & w33066;
assign w33960 = w33912 & w33959;
assign w33961 = ~w33958 & ~w33960;
assign w33962 = ~w33956 & w33961;
assign w33963 = w33955 & ~w33962;
assign w33964 = ~w33935 & ~w33963;
assign w33965 = ~w33924 & w33964;
assign w33966 = (~w33935 & w33954) | (~w33935 & w42708) | (w33954 & w42708);
assign w33967 = w33043 & ~w33099;
assign w33968 = ~w33005 & w33928;
assign w33969 = w33034 & ~w33968;
assign w33970 = w33967 & ~w33969;
assign w33971 = ~w33967 & w33969;
assign w33972 = ~w33970 & ~w33971;
assign w33973 = (w33972 & w32997) | (w33972 & w42709) | (w32997 & w42709);
assign w33974 = w33729 & w33972;
assign w33975 = ~w33697 & w33974;
assign w33976 = ~w33973 & ~w33975;
assign w33977 = ~w32997 & w42710;
assign w33978 = ~w33730 & w33977;
assign w33979 = w33976 & ~w33978;
assign w33980 = ~w33095 & ~w33144;
assign w33981 = w33084 & ~w33099;
assign w33982 = w33980 & ~w33981;
assign w33983 = ~w33980 & w33981;
assign w33984 = ~w33982 & ~w33983;
assign w33985 = ~w24874 & ~w33094;
assign w33986 = ~w33730 & w42711;
assign w33987 = ~w24874 & ~w33984;
assign w33988 = (w33987 & w33730) | (w33987 & w42712) | (w33730 & w42712);
assign w33989 = ~w33986 & ~w33988;
assign w33990 = (~w25851 & ~w33976) | (~w25851 & w49710) | (~w33976 & w49710);
assign w33991 = w33989 & ~w33990;
assign w33992 = ~w33966 & w33991;
assign w33993 = w24874 & w33109;
assign w33994 = (w33084 & w47965) | (w33084 & w47966) | (w47965 & w47966);
assign w33995 = w33126 & ~w33994;
assign w33996 = ~w33130 & ~w33995;
assign w33997 = ~w22767 & ~w33996;
assign w33998 = w31858 & ~w33136;
assign w33999 = ~w31858 & w33136;
assign w34000 = ~w33998 & ~w33999;
assign w34001 = w22767 & w33996;
assign w34002 = w33997 & ~w34000;
assign w34003 = ~w34001 & ~w34002;
assign w34004 = ~w33997 & w34000;
assign w34005 = ~w32997 & w42714;
assign w34006 = (~w34004 & w33730) | (~w34004 & w42715) | (w33730 & w42715);
assign w34007 = ~w33731 & ~w34003;
assign w34008 = w34006 & ~w34007;
assign w34009 = w33142 & ~w33995;
assign w34010 = w33198 & w34009;
assign w34011 = (w34010 & w33730) | (w34010 & w42716) | (w33730 & w42716);
assign w34012 = w21801 & ~w34011;
assign w34013 = ~w34008 & w34012;
assign w34014 = (w33084 & w47967) | (w33084 & w47968) | (w47967 & w47968);
assign w34015 = ~w24874 & w52273;
assign w34016 = ~w34014 & ~w34015;
assign w34017 = w33728 & w47969;
assign w34018 = ~w33697 & w34017;
assign w34019 = ~w33109 & ~w34016;
assign w34020 = w33728 & w47970;
assign w34021 = ~w33697 & w34020;
assign w34022 = ~w34021 & w42719;
assign w34023 = ~w34018 & w42720;
assign w34024 = w34022 & ~w34023;
assign w34025 = ~w33110 & ~w33993;
assign w34026 = ~w26447 & ~w34025;
assign w34027 = w23843 & ~w33110;
assign w34028 = w34027 & w52273;
assign w34029 = ~w34026 & ~w34028;
assign w34030 = ~w23843 & w33994;
assign w34031 = w34029 & ~w34030;
assign w34032 = w33728 & w47971;
assign w34033 = ~w33697 & w34032;
assign w34034 = ~w22767 & ~w33129;
assign w34035 = (w34034 & w34033) | (w34034 & w42722) | (w34033 & w42722);
assign w34036 = ~w22767 & w33129;
assign w34037 = ~w34033 & w42723;
assign w34038 = ~w34035 & ~w34037;
assign w34039 = ~w34024 & w34038;
assign w34040 = ~w34013 & w34039;
assign w34041 = w33198 & ~w34009;
assign w34042 = ~w33193 & ~w33208;
assign w34043 = w34041 & ~w34042;
assign w34044 = ~w34041 & w34042;
assign w34045 = ~w34043 & ~w34044;
assign w34046 = w33192 & w33731;
assign w34047 = ~w33731 & w34045;
assign w34048 = ~w34046 & ~w34047;
assign w34049 = ~w20906 & ~w34048;
assign w34050 = ~w33161 & ~w33210;
assign w34051 = ~w33161 & w33199;
assign w34052 = ~w34009 & w34051;
assign w34053 = ~w34050 & ~w34052;
assign w34054 = ~w33178 & ~w33207;
assign w34055 = ~w34053 & w34054;
assign w34056 = w34053 & ~w34054;
assign w34057 = ~w33731 & w42724;
assign w34058 = w33177 & w33731;
assign w34059 = (w19040 & ~w33731) | (w19040 & w42725) | (~w33731 & w42725);
assign w34060 = ~w34057 & w34059;
assign w34061 = (w20906 & w32997) | (w20906 & w42726) | (w32997 & w42726);
assign w34062 = w33728 & w46046;
assign w34063 = ~w33697 & w34062;
assign w34064 = ~w34061 & ~w34063;
assign w34065 = w33199 & ~w34009;
assign w34066 = ~w33208 & ~w34065;
assign w34067 = w21801 & ~w32698;
assign w34068 = w32698 & w33154;
assign w34069 = ~w34067 & ~w34068;
assign w34070 = w33148 & w34069;
assign w34071 = ~w33148 & ~w34069;
assign w34072 = ~w34070 & ~w34071;
assign w34073 = w20000 & w34072;
assign w34074 = w20000 & ~w34072;
assign w34075 = w34066 & w34073;
assign w34076 = ~w34064 & w34075;
assign w34077 = w34066 & w34074;
assign w34078 = w34064 & w34077;
assign w34079 = ~w34076 & ~w34078;
assign w34080 = (~w20906 & w32997) | (~w20906 & w42727) | (w32997 & w42727);
assign w34081 = w33728 & w46047;
assign w34082 = ~w33697 & w34081;
assign w34083 = ~w34080 & ~w34082;
assign w34084 = ~w34066 & w34073;
assign w34085 = ~w34083 & w34084;
assign w34086 = ~w34066 & w34074;
assign w34087 = w34083 & w34086;
assign w34088 = ~w34085 & ~w34087;
assign w34089 = w34079 & w34088;
assign w34090 = ~w34060 & w34089;
assign w34091 = ~w34049 & w34090;
assign w34092 = w34040 & w34091;
assign w34093 = w33992 & w34092;
assign w34094 = ~w33965 & w34093;
assign w34095 = (w33129 & w34033) | (w33129 & w42728) | (w34033 & w42728);
assign w34096 = ~w34033 & w42729;
assign w34097 = ~w34095 & ~w34096;
assign w34098 = w22767 & ~w34097;
assign w34099 = (~w34011 & w34007) | (~w34011 & w42730) | (w34007 & w42730);
assign w34100 = ~w34013 & w34098;
assign w34101 = ~w21801 & ~w34099;
assign w34102 = ~w34100 & ~w34101;
assign w34103 = w20906 & w34048;
assign w34104 = ~w34066 & w34072;
assign w34105 = ~w34083 & w34104;
assign w34106 = ~w34066 & ~w34072;
assign w34107 = w34083 & w34106;
assign w34108 = ~w34105 & ~w34107;
assign w34109 = w34066 & w34072;
assign w34110 = ~w34064 & w34109;
assign w34111 = w34066 & ~w34072;
assign w34112 = w34064 & w34111;
assign w34113 = ~w34110 & ~w34112;
assign w34114 = w34108 & w34113;
assign w34115 = ~w20000 & w34114;
assign w34116 = ~w34103 & ~w34115;
assign w34117 = w34091 & ~w34102;
assign w34118 = w34090 & ~w34116;
assign w34119 = ~w34117 & ~w34118;
assign w34120 = w33976 & w46048;
assign w34121 = w33989 & w34120;
assign w34122 = (w23843 & w34021) | (w23843 & w42731) | (w34021 & w42731);
assign w34123 = w23843 & w33109;
assign w34124 = ~w34018 & w42732;
assign w34125 = ~w34122 & ~w34124;
assign w34126 = w24874 & w33094;
assign w34127 = ~w33730 & w42733;
assign w34128 = w24874 & w33984;
assign w34129 = (w34128 & w33730) | (w34128 & w42734) | (w33730 & w42734);
assign w34130 = ~w34127 & ~w34129;
assign w34131 = w34125 & w34130;
assign w34132 = ~w34121 & w34131;
assign w34133 = w34040 & ~w34132;
assign w34134 = w34091 & w34133;
assign w34135 = w19040 & ~w32698;
assign w34136 = w32698 & ~w33221;
assign w34137 = ~w34135 & ~w34136;
assign w34138 = w33215 & ~w34137;
assign w34139 = ~w33215 & w34137;
assign w34140 = ~w34138 & ~w34139;
assign w34141 = ~w33229 & ~w33302;
assign w34142 = w33214 & ~w33290;
assign w34143 = ~w33203 & w34142;
assign w34144 = (w34141 & w34143) | (w34141 & w47972) | (w34143 & w47972);
assign w34145 = ~w34143 & w47973;
assign w34146 = ~w34144 & ~w34145;
assign w34147 = ~w33730 & w42735;
assign w34148 = (w34146 & w33730) | (w34146 & w42736) | (w33730 & w42736);
assign w34149 = ~w34147 & ~w34148;
assign w34150 = ~w17380 & ~w34149;
assign w34151 = ~w33203 & w33214;
assign w34152 = ~w33290 & ~w33299;
assign w34153 = w34151 & ~w34152;
assign w34154 = ~w34151 & w34152;
assign w34155 = ~w34153 & ~w34154;
assign w34156 = ~w33730 & w42737;
assign w34157 = (w34155 & w33730) | (w34155 & w42738) | (w33730 & w42738);
assign w34158 = ~w34156 & ~w34157;
assign w34159 = ~w18183 & ~w34158;
assign w34160 = ~w34150 & w34159;
assign w34161 = w17380 & w34149;
assign w34162 = ~w34057 & ~w34058;
assign w34163 = ~w19040 & ~w34162;
assign w34164 = ~w34160 & ~w34163;
assign w34165 = ~w34161 & w34164;
assign w34166 = ~w34134 & w34165;
assign w34167 = w34119 & w34166;
assign w34168 = ~w34094 & w34167;
assign w34169 = w33247 & w34143;
assign w34170 = ~w33251 & ~w33304;
assign w34171 = (w34170 & ~w34143) | (w34170 & w42739) | (~w34143 & w42739);
assign w34172 = ~w33260 & ~w33292;
assign w34173 = w34171 & ~w34172;
assign w34174 = ~w34171 & w34172;
assign w34175 = ~w34173 & ~w34174;
assign w34176 = w15681 & w33259;
assign w34177 = ~w33730 & w42740;
assign w34178 = w15681 & w34175;
assign w34179 = ~w33731 & w34178;
assign w34180 = ~w34177 & ~w34179;
assign w34181 = ~w15681 & ~w33259;
assign w34182 = w16559 & ~w33250;
assign w34183 = ~w34181 & w34182;
assign w34184 = ~w15681 & w33259;
assign w34185 = w34171 & w34184;
assign w34186 = w16559 & ~w34185;
assign w34187 = w33246 & w33303;
assign w34188 = ~w34143 & w34187;
assign w34189 = w33229 & w33246;
assign w34190 = ~w33304 & ~w34189;
assign w34191 = ~w34169 & ~w34188;
assign w34192 = w34190 & w34191;
assign w34193 = ~w34171 & w34181;
assign w34194 = w34192 & ~w34193;
assign w34195 = ~w33730 & w42741;
assign w34196 = w34186 & w34194;
assign w34197 = (~w34195 & ~w34196) | (~w34195 & w47974) | (~w34196 & w47974);
assign w34198 = w34180 & w34197;
assign w34199 = w14039 & w14302;
assign w34200 = ~w14766 & w34199;
assign w34201 = (~w11870 & ~w34198) | (~w11870 & w42742) | (~w34198 & w42742);
assign w34202 = ~w33323 & ~w33324;
assign w34203 = w33361 & w33373;
assign w34204 = (w14766 & w33298) | (w14766 & w42743) | (w33298 & w42743);
assign w34205 = ~w33298 & w42744;
assign w34206 = (~w33351 & w33298) | (~w33351 & w47975) | (w33298 & w47975);
assign w34207 = w34203 & ~w34204;
assign w34208 = ~w34206 & w34207;
assign w34209 = ~w33335 & w33368;
assign w34210 = ~w33731 & w42745;
assign w34211 = w12666 & w33731;
assign w34212 = (w33335 & w33730) | (w33335 & w42746) | (w33730 & w42746);
assign w34213 = ~w34211 & ~w34212;
assign w34214 = (w34202 & ~w34213) | (w34202 & w42747) | (~w34213 & w42747);
assign w34215 = w34213 & w42748;
assign w34216 = ~w34214 & ~w34215;
assign w34217 = ~w34201 & w34216;
assign w34218 = w18183 & w34158;
assign w34219 = ~w34161 & w34218;
assign w34220 = ~w34150 & ~w34219;
assign w34221 = ~w33334 & w33731;
assign w34222 = ~w34210 & ~w34221;
assign w34223 = ~w33731 & w42749;
assign w34224 = w34222 & ~w34223;
assign w34225 = ~w12666 & ~w34224;
assign w34226 = w12666 & ~w34223;
assign w34227 = w34222 & w34226;
assign w34228 = ~w34204 & ~w34206;
assign w34229 = w34203 & w34228;
assign w34230 = ~w31718 & ~w32698;
assign w34231 = w32698 & w33356;
assign w34232 = ~w34230 & ~w34231;
assign w34233 = ~w34203 & ~w34228;
assign w34234 = w33731 & w34232;
assign w34235 = ~w33731 & w42750;
assign w34236 = ~w34234 & ~w34235;
assign w34237 = w13384 & w34236;
assign w34238 = ~w34227 & w34237;
assign w34239 = ~w34225 & ~w34238;
assign w34240 = ~w33402 & ~w33500;
assign w34241 = (w33459 & w33298) | (w33459 & w42751) | (w33298 & w42751);
assign w34242 = ~w33378 & ~w34241;
assign w34243 = w34240 & ~w34242;
assign w34244 = ~w34240 & w34242;
assign w34245 = ~w34243 & ~w34244;
assign w34246 = w33401 & w33731;
assign w34247 = ~w33731 & w34245;
assign w34248 = ~w34246 & ~w34247;
assign w34249 = w11138 & ~w34248;
assign w34250 = ~w11870 & w34202;
assign w34251 = (w34250 & ~w34213) | (w34250 & w42752) | (~w34213 & w42752);
assign w34252 = ~w11870 & ~w34202;
assign w34253 = w34213 & w42753;
assign w34254 = ~w34251 & ~w34253;
assign w34255 = ~w34249 & w34254;
assign w34256 = w34239 & w34255;
assign w34257 = ~w33275 & ~w33291;
assign w34258 = ~w33292 & w34257;
assign w34259 = ~w33260 & w34171;
assign w34260 = w34258 & ~w34259;
assign w34261 = ~w33260 & ~w34257;
assign w34262 = ~w34174 & w34261;
assign w34263 = ~w34260 & ~w34262;
assign w34264 = ~w33730 & w42754;
assign w34265 = ~w33731 & w34263;
assign w34266 = ~w34264 & ~w34265;
assign w34267 = ~w34265 & w42755;
assign w34268 = ~w34198 & ~w34267;
assign w34269 = ~w34204 & ~w34205;
assign w34270 = (w34269 & w33730) | (w34269 & w42756) | (w33730 & w42756);
assign w34271 = w33351 & ~w34270;
assign w34272 = ~w33351 & w34269;
assign w34273 = (w34272 & w33730) | (w34272 & w42757) | (w33730 & w42757);
assign w34274 = ~w14039 & ~w34273;
assign w34275 = ~w34271 & w34274;
assign w34276 = (w14766 & w34265) | (w14766 & w42758) | (w34265 & w42758);
assign w34277 = ~w34275 & ~w34276;
assign w34278 = ~w34268 & w34277;
assign w34279 = w34220 & w34278;
assign w34280 = w34217 & w34220;
assign w34281 = w34256 & w34279;
assign w34282 = ~w34280 & ~w34281;
assign w34283 = ~w34168 & ~w34282;
assign w34284 = ~w33392 & w33505;
assign w34285 = ~w33378 & ~w33402;
assign w34286 = w34285 & ~w34241;
assign w34287 = ~w33500 & ~w34286;
assign w34288 = w34284 & ~w34287;
assign w34289 = ~w34284 & w34287;
assign w34290 = w33391 & w33731;
assign w34291 = ~w33731 & w42759;
assign w34292 = ~w34290 & ~w34291;
assign w34293 = w10419 & ~w34292;
assign w34294 = ~w16559 & w33250;
assign w34295 = ~w33730 & w42760;
assign w34296 = ~w16559 & ~w34192;
assign w34297 = ~w33731 & w34296;
assign w34298 = ~w34295 & ~w34297;
assign w34299 = ~w33730 & w42761;
assign w34300 = ~w15681 & ~w34175;
assign w34301 = ~w33731 & w34300;
assign w34302 = ~w34299 & ~w34301;
assign w34303 = w34298 & w34302;
assign w34304 = (~w34267 & w34303) | (~w34267 & w42762) | (w34303 & w42762);
assign w34305 = w34278 & ~w34304;
assign w34306 = ~w13384 & ~w34236;
assign w34307 = ~w34271 & ~w34273;
assign w34308 = w14039 & ~w34307;
assign w34309 = ~w34227 & ~w34306;
assign w34310 = ~w34308 & w34309;
assign w34311 = ~w34305 & w34310;
assign w34312 = ~w11138 & w34248;
assign w34313 = ~w11870 & w34303;
assign w34314 = w34217 & ~w34313;
assign w34315 = ~w34312 & ~w34314;
assign w34316 = w34256 & ~w34311;
assign w34317 = w34315 & ~w34316;
assign w34318 = ~w34316 & w42763;
assign w34319 = ~w34283 & w34318;
assign w34320 = ~w33438 & ~w33670;
assign w34321 = w33405 & w33669;
assign w34322 = ~w33298 & w34321;
assign w34323 = (w34320 & w34322) | (w34320 & w42765) | (w34322 & w42765);
assign w34324 = ~w34322 & w42766;
assign w34325 = ~w34323 & ~w34324;
assign w34326 = ~w5745 & ~w33437;
assign w34327 = ~w33730 & w42767;
assign w34328 = ~w5745 & w34325;
assign w34329 = ~w33731 & w34328;
assign w34330 = ~w34327 & ~w34329;
assign w34331 = ~w33450 & ~w33667;
assign w34332 = ~w33656 & ~w33666;
assign w34333 = w33405 & w34332;
assign w34334 = ~w33298 & w34333;
assign w34335 = (w34331 & w34334) | (w34331 & w42768) | (w34334 & w42768);
assign w34336 = ~w34334 & w42769;
assign w34337 = ~w34335 & ~w34336;
assign w34338 = w6264 & w33449;
assign w34339 = ~w33730 & w42770;
assign w34340 = w6264 & w34337;
assign w34341 = ~w33731 & w34340;
assign w34342 = ~w34339 & ~w34341;
assign w34343 = w34330 & w34342;
assign w34344 = w6769 & w33664;
assign w34345 = w6769 & ~w33664;
assign w34346 = w7315 & w34344;
assign w34347 = ~w7315 & w34345;
assign w34348 = ~w34346 & ~w34347;
assign w34349 = w33471 & ~w33655;
assign w34350 = w33405 & ~w34349;
assign w34351 = ~w33298 & w34350;
assign w34352 = ~w33507 & w42771;
assign w34353 = (~w34349 & w33461) | (~w34349 & w42772) | (w33461 & w42772);
assign w34354 = (~w33659 & w34351) | (~w33659 & w42773) | (w34351 & w42773);
assign w34355 = (w34351 & w47976) | (w34351 & w47977) | (w47976 & w47977);
assign w34356 = w34345 & ~w34354;
assign w34357 = ~w34355 & ~w34356;
assign w34358 = ~w33730 & w42774;
assign w34359 = ~w33731 & ~w34357;
assign w34360 = ~w34358 & ~w34359;
assign w34361 = ~w6264 & ~w33449;
assign w34362 = ~w33730 & w42775;
assign w34363 = ~w6264 & ~w34337;
assign w34364 = ~w33731 & w34363;
assign w34365 = ~w34362 & ~w34364;
assign w34366 = w34360 & w34365;
assign w34367 = w34343 & ~w34366;
assign w34368 = ~w33429 & w33674;
assign w34369 = (~w33670 & w34322) | (~w33670 & w47978) | (w34322 & w47978);
assign w34370 = ~w34368 & ~w34369;
assign w34371 = w34368 & w34369;
assign w34372 = ~w33731 & w42777;
assign w34373 = (~w5330 & ~w33731) | (~w5330 & w42778) | (~w33731 & w42778);
assign w34374 = ~w34372 & w34373;
assign w34375 = ~w33730 & w42779;
assign w34376 = w5745 & ~w34375;
assign w34377 = ~w33731 & w34325;
assign w34378 = w34376 & ~w34377;
assign w34379 = ~w34374 & ~w34378;
assign w34380 = ~w34367 & w34379;
assign w34381 = ~w33730 & w42780;
assign w34382 = (w34354 & w33730) | (w34354 & w42781) | (w33730 & w42781);
assign w34383 = ~w34381 & ~w34382;
assign w34384 = ~w6769 & w33664;
assign w34385 = w34383 & w34384;
assign w34386 = ~w6769 & ~w33664;
assign w34387 = ~w34383 & w34386;
assign w34388 = ~w34385 & ~w34387;
assign w34389 = w34343 & w34388;
assign w34390 = w34380 & ~w34389;
assign w34391 = (w33452 & w33555) | (w33452 & w42782) | (w33555 & w42782);
assign w34392 = (~w33676 & w34322) | (~w33676 & w42783) | (w34322 & w42783);
assign w34393 = ~w33690 & w34392;
assign w34394 = ~w33425 & ~w34393;
assign w34395 = ~w33730 & w42784;
assign w34396 = ~w33731 & w34394;
assign w34397 = ~w33689 & ~w33699;
assign w34398 = w4430 & ~w34397;
assign w34399 = ~w34396 & w42785;
assign w34400 = w4430 & w34397;
assign w34401 = (w34400 & w34396) | (w34400 & w42786) | (w34396 & w42786);
assign w34402 = ~w34399 & ~w34401;
assign w34403 = ~w5745 & w33731;
assign w34404 = ~w33731 & w34369;
assign w34405 = ~w34403 & ~w34404;
assign w34406 = w34368 & ~w34405;
assign w34407 = ~w34368 & w34405;
assign w34408 = ~w34406 & ~w34407;
assign w34409 = w5330 & w34408;
assign w34410 = ~w4430 & ~w34397;
assign w34411 = (w34410 & w34396) | (w34410 & w42787) | (w34396 & w42787);
assign w34412 = ~w4430 & w34397;
assign w34413 = ~w34396 & w42788;
assign w34414 = ~w34411 & ~w34413;
assign w34415 = ~w33425 & ~w33690;
assign w34416 = w34392 & ~w34415;
assign w34417 = ~w34392 & w34415;
assign w34418 = ~w34416 & ~w34417;
assign w34419 = w33424 & w33731;
assign w34420 = ~w33731 & w34418;
assign w34421 = ~w34419 & ~w34420;
assign w34422 = ~w4838 & w34421;
assign w34423 = w33622 & ~w33703;
assign w34424 = (~w34423 & w33557) | (~w34423 & w42789) | (w33557 & w42789);
assign w34425 = ~w33610 & w33627;
assign w34426 = ~w33702 & w34425;
assign w34427 = (w33557 & w47979) | (w33557 & w47980) | (w47979 & w47980);
assign w34428 = w34425 & ~w34424;
assign w34429 = ~w33731 & ~w34428;
assign w34430 = ~w33731 & w42790;
assign w34431 = ~w33730 & w42791;
assign w34432 = w3646 & ~w34431;
assign w34433 = ~w34430 & w34432;
assign w34434 = ~w33695 & ~w33699;
assign w34435 = w33555 & w42792;
assign w34436 = ~w33406 & w34435;
assign w34437 = ~w34436 & w42793;
assign w34438 = ~w34424 & ~w34437;
assign w34439 = w4838 & ~w32698;
assign w34440 = w32698 & ~w33614;
assign w34441 = ~w34439 & ~w34440;
assign w34442 = w33615 & ~w34441;
assign w34443 = ~w33615 & w34441;
assign w34444 = ~w34442 & ~w34443;
assign w34445 = ~w32997 & w42794;
assign w34446 = ~w33730 & w34445;
assign w34447 = (~w33622 & w34436) | (~w33622 & w47981) | (w34436 & w47981);
assign w34448 = ~w34446 & ~w34447;
assign w34449 = ~w33731 & w34438;
assign w34450 = w34448 & ~w34449;
assign w34451 = w4056 & w34450;
assign w34452 = ~w3646 & w34431;
assign w34453 = ~w3646 & ~w34427;
assign w34454 = w34429 & w34453;
assign w34455 = ~w34452 & ~w34454;
assign w34456 = ~w34451 & w34455;
assign w34457 = ~w34433 & ~w34456;
assign w34458 = w34414 & w34422;
assign w34459 = ~w34457 & ~w34458;
assign w34460 = w34402 & ~w34409;
assign w34461 = ~w34390 & w34459;
assign w34462 = w34460 & w34461;
assign w34463 = ~w33461 & ~w33507;
assign w34464 = ~w33641 & ~w33646;
assign w34465 = ~w33643 & w33652;
assign w34466 = w33471 & w34465;
assign w34467 = w34464 & ~w34466;
assign w34468 = ~w34464 & w34466;
assign w34469 = ~w34467 & ~w34468;
assign w34470 = (~w34469 & w33406) | (~w34469 & w42795) | (w33406 & w42795);
assign w34471 = ~w33406 & w42796;
assign w34472 = ~w33465 & ~w33466;
assign w34473 = w33465 & w33466;
assign w34474 = ~w34472 & ~w34473;
assign w34475 = ~w33730 & w42797;
assign w34476 = w7924 & ~w34475;
assign w34477 = ~w34470 & ~w34471;
assign w34478 = ~w33731 & w34477;
assign w34479 = w34476 & ~w34478;
assign w34480 = ~w33461 & w42798;
assign w34481 = w33536 & w33640;
assign w34482 = ~w34480 & w34481;
assign w34483 = w33405 & w34481;
assign w34484 = ~w33298 & w34483;
assign w34485 = w33524 & ~w33646;
assign w34486 = ~w33536 & ~w34485;
assign w34487 = w33536 & w34485;
assign w34488 = ~w34486 & ~w34487;
assign w34489 = ~w8666 & w34485;
assign w34490 = (w34489 & w34484) | (w34489 & w42799) | (w34484 & w42799);
assign w34491 = ~w8666 & w34488;
assign w34492 = ~w34484 & w42800;
assign w34493 = ~w34490 & ~w34492;
assign w34494 = ~w33634 & ~w34480;
assign w34495 = w33405 & ~w33634;
assign w34496 = ~w33298 & w34495;
assign w34497 = ~w34494 & ~w34496;
assign w34498 = ~w31575 & ~w32698;
assign w34499 = w32698 & ~w33531;
assign w34500 = ~w34498 & ~w34499;
assign w34501 = ~w34496 & w42801;
assign w34502 = ~w9781 & w34500;
assign w34503 = (w34502 & w34496) | (w34502 & w42802) | (w34496 & w42802);
assign w34504 = ~w34501 & ~w34503;
assign w34505 = w34493 & w34504;
assign w34506 = ~w33731 & ~w34505;
assign w34507 = w9781 & ~w32249;
assign w34508 = w31646 & ~w34507;
assign w34509 = ~w32698 & w34508;
assign w34510 = ~w33520 & ~w34509;
assign w34511 = ~w8666 & w34510;
assign w34512 = w34500 & ~w34511;
assign w34513 = ~w32997 & w42803;
assign w34514 = ~w34496 & w42804;
assign w34515 = ~w9195 & ~w34514;
assign w34516 = w9781 & ~w34500;
assign w34517 = ~w34497 & w34516;
assign w34518 = w34515 & ~w34517;
assign w34519 = ~w33730 & w34513;
assign w34520 = w34518 & ~w34519;
assign w34521 = (w34485 & w34484) | (w34485 & w42805) | (w34484 & w42805);
assign w34522 = ~w34484 & w42806;
assign w34523 = ~w34521 & ~w34522;
assign w34524 = w8666 & ~w34510;
assign w34525 = ~w33730 & w42807;
assign w34526 = w8666 & w34523;
assign w34527 = ~w33731 & w34526;
assign w34528 = ~w34525 & ~w34527;
assign w34529 = ~w34506 & w34520;
assign w34530 = w34528 & ~w34529;
assign w34531 = ~w7924 & w34477;
assign w34532 = ~w33731 & w34531;
assign w34533 = ~w7924 & ~w34474;
assign w34534 = ~w33730 & w42808;
assign w34535 = ~w34532 & ~w34534;
assign w34536 = (w34535 & ~w34530) | (w34535 & w42809) | (~w34530 & w42809);
assign w34537 = ~w33476 & ~w33657;
assign w34538 = (w7924 & w34351) | (w7924 & w47982) | (w34351 & w47982);
assign w34539 = ~w34351 & w47983;
assign w34540 = ~w34538 & ~w34539;
assign w34541 = (w34537 & w33731) | (w34537 & w42810) | (w33731 & w42810);
assign w34542 = ~w33731 & w42811;
assign w34543 = ~w34541 & ~w34542;
assign w34544 = w7315 & w34543;
assign w34545 = (w9781 & w34496) | (w9781 & w42812) | (w34496 & w42812);
assign w34546 = ~w34496 & w42813;
assign w34547 = ~w34545 & ~w34546;
assign w34548 = w9195 & ~w34500;
assign w34549 = ~w34547 & w34548;
assign w34550 = ~w34511 & ~w34548;
assign w34551 = ~w33730 & w42814;
assign w34552 = w9195 & w34500;
assign w34553 = w34547 & w34552;
assign w34554 = w34493 & ~w34553;
assign w34555 = (w34463 & w33298) | (w34463 & w42815) | (w33298 & w42815);
assign w34556 = ~w33551 & ~w33634;
assign w34557 = w34555 & ~w34556;
assign w34558 = ~w34555 & w34556;
assign w34559 = ~w34557 & ~w34558;
assign w34560 = ~w9781 & w33550;
assign w34561 = ~w33730 & w42816;
assign w34562 = ~w9781 & ~w34559;
assign w34563 = ~w33731 & w34562;
assign w34564 = ~w34561 & ~w34563;
assign w34565 = ~w33731 & ~w34554;
assign w34566 = w34564 & ~w34565;
assign w34567 = ~w34549 & ~w34551;
assign w34568 = w34535 & w34567;
assign w34569 = w34566 & w34568;
assign w34570 = ~w34544 & ~w34569;
assign w34571 = ~w34536 & w34570;
assign w34572 = ~w7315 & ~w34543;
assign w34573 = ~w34367 & w42817;
assign w34574 = ~w34571 & w34573;
assign w34575 = w34462 & ~w34574;
assign w34576 = w4838 & ~w34421;
assign w34577 = ~w4056 & ~w34450;
assign w34578 = ~w34433 & ~w34577;
assign w34579 = w34414 & w34578;
assign w34580 = w34402 & w34576;
assign w34581 = w34579 & ~w34580;
assign w34582 = ~w34457 & ~w34581;
assign w34583 = ~w10419 & w34292;
assign w34584 = ~w34293 & ~w34312;
assign w34585 = ~w34583 & ~w34584;
assign w34586 = ~w34249 & ~w34583;
assign w34587 = w34254 & w34586;
assign w34588 = ~w34585 & ~w34587;
assign w34589 = ~w34582 & ~w34588;
assign w34590 = ~w34575 & w34589;
assign w34591 = ~w34319 & w34590;
assign w34592 = w32807 & w32813;
assign w34593 = ~w32987 & ~w33791;
assign w34594 = ~w33730 & w49711;
assign w34595 = ~w33731 & w42818;
assign w34596 = (w34592 & w34595) | (w34592 & w49712) | (w34595 & w49712);
assign w34597 = ~w34595 & w49713;
assign w34598 = ~w34596 & ~w34597;
assign w34599 = w400 & ~w34598;
assign w34600 = ~w33730 & w49714;
assign w34601 = (w32807 & w33730) | (w32807 & w42819) | (w33730 & w42819);
assign w34602 = ~w33835 & w34601;
assign w34603 = w32799 & ~w32983;
assign w34604 = ~w34602 & w49715;
assign w34605 = (w34603 & w34602) | (w34603 & w49716) | (w34602 & w49716);
assign w34606 = ~w34604 & ~w34605;
assign w34607 = ~w351 & w34606;
assign w34608 = ~w34599 & ~w34607;
assign w34609 = w32979 & ~w33809;
assign w34610 = w32830 & ~w32987;
assign w34611 = w32986 & w33731;
assign w34612 = (~w34610 & w33730) | (~w34610 & w42820) | (w33730 & w42820);
assign w34613 = w34609 & w34612;
assign w34614 = (w34610 & w33730) | (w34610 & w42821) | (w33730 & w42821);
assign w34615 = ~w34609 & w34614;
assign w34616 = ~w34613 & ~w34615;
assign w34617 = ~w34611 & w34616;
assign w34618 = w34616 & w49717;
assign w34619 = (w32842 & w33730) | (w32842 & w42822) | (w33730 & w42822);
assign w34620 = (w32974 & w33739) | (w32974 & w46049) | (w33739 & w46049);
assign w34621 = w34619 & ~w34620;
assign w34622 = ~w33730 & w47984;
assign w34623 = w32854 & ~w32977;
assign w34624 = w612 & w34623;
assign w34625 = (w34624 & w34621) | (w34624 & w49718) | (w34621 & w49718);
assign w34626 = w612 & ~w34623;
assign w34627 = ~w34621 & w49719;
assign w34628 = ~w34625 & ~w34627;
assign w34629 = (w493 & ~w34616) | (w493 & w49720) | (~w34616 & w49720);
assign w34630 = ~w400 & ~w34592;
assign w34631 = (w34630 & w34595) | (w34630 & w49721) | (w34595 & w49721);
assign w34632 = ~w400 & w34592;
assign w34633 = ~w34595 & w49722;
assign w34634 = ~w34631 & ~w34633;
assign w34635 = ~w34629 & w34634;
assign w34636 = ~w34618 & ~w34628;
assign w34637 = w34635 & ~w34636;
assign w34638 = ~w945 & w33746;
assign w34639 = w945 & w32860;
assign w34640 = w32842 & ~w34639;
assign w34641 = w32842 & w32860;
assign w34642 = w32973 & ~w34641;
assign w34643 = ~w33730 & w47985;
assign w34644 = ~w33731 & w42823;
assign w34645 = ~w34643 & ~w34644;
assign w34646 = w32860 & w34621;
assign w34647 = w34645 & ~w34646;
assign w34648 = w754 & ~w34647;
assign w34649 = ~w34638 & ~w34648;
assign w34650 = ~w754 & w34647;
assign w34651 = ~w612 & ~w34623;
assign w34652 = (w34651 & w34621) | (w34651 & w47986) | (w34621 & w47986);
assign w34653 = ~w612 & w34623;
assign w34654 = ~w34621 & w47987;
assign w34655 = ~w34652 & ~w34654;
assign w34656 = ~w34650 & w34655;
assign w34657 = ~w34650 & w49723;
assign w34658 = ~w34649 & w34657;
assign w34659 = w34637 & ~w34658;
assign w34660 = (w34608 & w34658) | (w34608 & w47988) | (w34658 & w47988);
assign w34661 = ~w252 & ~w33844;
assign w34662 = w351 & ~w34606;
assign w34663 = ~w34661 & ~w34662;
assign w34664 = ~w34660 & w34663;
assign w34665 = w34637 & ~w34657;
assign w34666 = ~w32997 & w42824;
assign w34667 = ~w33730 & w34666;
assign w34668 = ~w33610 & ~w33628;
assign w34669 = w33590 & w33711;
assign w34670 = ~w33590 & ~w33705;
assign w34671 = w33711 & ~w34670;
assign w34672 = w33599 & w52274;
assign w34673 = ~w33731 & w34672;
assign w34674 = ~w34667 & ~w34673;
assign w34675 = ~w33578 & w33716;
assign w34676 = ~w2558 & ~w34675;
assign w34677 = (w34676 & w34673) | (w34676 & w42827) | (w34673 & w42827);
assign w34678 = ~w2558 & w34675;
assign w34679 = ~w34673 & w42828;
assign w34680 = ~w34677 & ~w34679;
assign w34681 = w33555 & w42829;
assign w34682 = ~w33406 & w34681;
assign w34683 = (w33705 & ~w33695) | (w33705 & w42830) | (~w33695 & w42830);
assign w34684 = ~w34682 & w42831;
assign w34685 = w33717 & ~w34684;
assign w34686 = ~w33599 & w33716;
assign w34687 = ~w33578 & ~w34686;
assign w34688 = (w34687 & w32997) | (w34687 & w42832) | (w32997 & w42832);
assign w34689 = w33728 & w47989;
assign w34690 = ~w33697 & w34689;
assign w34691 = ~w34688 & ~w34690;
assign w34692 = ~w33730 & w42833;
assign w34693 = ~w34685 & ~w34691;
assign w34694 = ~w34692 & ~w34693;
assign w34695 = ~w33567 & ~w33698;
assign w34696 = w2285 & ~w34695;
assign w34697 = (w34696 & w34693) | (w34696 & w42834) | (w34693 & w42834);
assign w34698 = w2285 & w34695;
assign w34699 = ~w34693 & w42835;
assign w34700 = ~w34697 & ~w34699;
assign w34701 = w34680 & w34700;
assign w34702 = w33599 & w33711;
assign w34703 = ~w33590 & ~w34702;
assign w34704 = ~w34682 & w42836;
assign w34705 = w33590 & w34702;
assign w34706 = w33695 & w42837;
assign w34707 = ~w34670 & w34702;
assign w34708 = (w34707 & w33557) | (w34707 & w42838) | (w33557 & w42838);
assign w34709 = w33593 & ~w33594;
assign w34710 = ~w33593 & w33594;
assign w34711 = ~w34709 & ~w34710;
assign w34712 = ~w33730 & w42839;
assign w34713 = ~w34704 & ~w34708;
assign w34714 = ~w33731 & w34713;
assign w34715 = ~w34712 & ~w34714;
assign w34716 = (~w2896 & w34714) | (~w2896 & w42840) | (w34714 & w42840);
assign w34717 = w2558 & ~w34675;
assign w34718 = (w34717 & w33730) | (w34717 & w42841) | (w33730 & w42841);
assign w34719 = ~w34673 & w34718;
assign w34720 = w2558 & w34675;
assign w34721 = ~w33730 & w42842;
assign w34722 = w33599 & w34720;
assign w34723 = w34722 & w52274;
assign w34724 = ~w33731 & w34723;
assign w34725 = ~w34721 & ~w34724;
assign w34726 = ~w34719 & w34725;
assign w34727 = ~w34716 & w34726;
assign w34728 = ~w34714 & w42843;
assign w34729 = ~w33610 & ~w33704;
assign w34730 = w33555 & w47990;
assign w34731 = ~w33406 & w34730;
assign w34732 = ~w34731 & w42845;
assign w34733 = (w3646 & w34731) | (w3646 & w42846) | (w34731 & w42846);
assign w34734 = ~w34732 & ~w34733;
assign w34735 = ~w33731 & w34734;
assign w34736 = w3242 & ~w33589;
assign w34737 = (w34736 & w33731) | (w34736 & w42847) | (w33731 & w42847);
assign w34738 = w3242 & w33589;
assign w34739 = ~w33731 & w42848;
assign w34740 = ~w34737 & ~w34739;
assign w34741 = ~w34728 & ~w34740;
assign w34742 = w34727 & ~w34741;
assign w34743 = w34701 & ~w34742;
assign w34744 = ~w32359 & ~w32913;
assign w34745 = ~w32912 & ~w34744;
assign w34746 = ~w33730 & w42849;
assign w34747 = ~w32932 & ~w33725;
assign w34748 = w33556 & ~w33721;
assign w34749 = ~w33406 & w34748;
assign w34750 = ~w33696 & ~w33721;
assign w34751 = w32917 & w32957;
assign w34752 = w32946 & ~w32952;
assign w34753 = ~w34751 & w34752;
assign w34754 = (w34753 & w42850) | (w34753 & w52275) | (w42850 & w52275);
assign w34755 = ~w34747 & w34751;
assign w34756 = ~w34749 & w46050;
assign w34757 = w34755 & ~w34756;
assign w34758 = ~w33731 & ~w34754;
assign w34759 = ~w34757 & w34758;
assign w34760 = (~w34746 & ~w34758) | (~w34746 & w42851) | (~w34758 & w42851);
assign w34761 = ~w1541 & ~w34760;
assign w34762 = ~w2285 & ~w33722;
assign w34763 = ~w33720 & w46051;
assign w34764 = w33631 & ~w34762;
assign w34765 = w33695 & w34764;
assign w34766 = ~w34763 & ~w34765;
assign w34767 = ~w34749 & ~w34766;
assign w34768 = ~w33723 & ~w34767;
assign w34769 = ~w32932 & ~w33724;
assign w34770 = ~w34767 & w42852;
assign w34771 = (w34769 & w34767) | (w34769 & w47991) | (w34767 & w47991);
assign w34772 = ~w33731 & ~w34770;
assign w34773 = ~w34771 & w34772;
assign w34774 = ~w34773 & w42853;
assign w34775 = ~w34761 & ~w34774;
assign w34776 = ~w2285 & ~w34695;
assign w34777 = ~w34693 & w42854;
assign w34778 = ~w2285 & w34695;
assign w34779 = (w34778 & w34693) | (w34778 & w42855) | (w34693 & w42855);
assign w34780 = ~w34777 & ~w34779;
assign w34781 = w32917 & ~w32959;
assign w34782 = ~w33720 & w47992;
assign w34783 = w33631 & ~w34781;
assign w34784 = w33695 & w34783;
assign w34785 = ~w34782 & ~w34784;
assign w34786 = ~w34755 & ~w34781;
assign w34787 = ~w34749 & ~w34785;
assign w34788 = ~w34786 & ~w34787;
assign w34789 = ~w33730 & w42856;
assign w34790 = ~w33731 & w34788;
assign w34791 = ~w34789 & ~w34790;
assign w34792 = ~w32900 & ~w32964;
assign w34793 = ~w1320 & ~w34792;
assign w34794 = (w34793 & w34790) | (w34793 & w42857) | (w34790 & w42857);
assign w34795 = ~w1320 & w34792;
assign w34796 = (w34795 & w34787) | (w34795 & w42858) | (w34787 & w42858);
assign w34797 = ~w33731 & w34796;
assign w34798 = w1541 & w34795;
assign w34799 = ~w33730 & w42859;
assign w34800 = ~w34797 & ~w34799;
assign w34801 = w2285 & w33727;
assign w34802 = w32789 & ~w34801;
assign w34803 = w32994 & w34802;
assign w34804 = w32996 & ~w34803;
assign w34805 = ~w34749 & w46052;
assign w34806 = (w33722 & w34803) | (w33722 & w42860) | (w34803 & w42860);
assign w34807 = ~w34805 & ~w34806;
assign w34808 = ~w2285 & w33722;
assign w34809 = (w34808 & w34749) | (w34808 & w47993) | (w34749 & w47993);
assign w34810 = w34807 & ~w34809;
assign w34811 = w2285 & ~w33722;
assign w34812 = (~w34811 & w34749) | (~w34811 & w46053) | (w34749 & w46053);
assign w34813 = ~w34767 & w34804;
assign w34814 = ~w34812 & w34813;
assign w34815 = (~w2006 & ~w34813) | (~w2006 & w46054) | (~w34813 & w46054);
assign w34816 = w34810 & w34815;
assign w34817 = w34800 & ~w34816;
assign w34818 = ~w34794 & w34817;
assign w34819 = w34780 & w34818;
assign w34820 = w34775 & w34819;
assign w34821 = ~w34743 & w34820;
assign w34822 = ~w33730 & w42861;
assign w34823 = w32911 & ~w32963;
assign w34824 = ~w32900 & w52276;
assign w34825 = ~w34823 & ~w34824;
assign w34826 = ~w33731 & ~w34825;
assign w34827 = w34823 & w34824;
assign w34828 = w34826 & ~w34827;
assign w34829 = ~w34822 & ~w34828;
assign w34830 = ~w1120 & w34829;
assign w34831 = w1541 & ~w34746;
assign w34832 = ~w34759 & w34831;
assign w34833 = ~w34775 & ~w34832;
assign w34834 = (w1738 & w34773) | (w1738 & w42863) | (w34773 & w42863);
assign w34835 = w34810 & ~w34814;
assign w34836 = (w2006 & ~w34810) | (w2006 & w42864) | (~w34810 & w42864);
assign w34837 = ~w34832 & ~w34836;
assign w34838 = ~w34834 & w34837;
assign w34839 = ~w34794 & w34800;
assign w34840 = (w34839 & ~w34837) | (w34839 & w42865) | (~w34837 & w42865);
assign w34841 = ~w34833 & w34840;
assign w34842 = ~w34791 & ~w34792;
assign w34843 = w34791 & w34792;
assign w34844 = ~w34842 & ~w34843;
assign w34845 = w1320 & w34844;
assign w34846 = ~w3242 & w33589;
assign w34847 = (w34846 & w33731) | (w34846 & w42866) | (w33731 & w42866);
assign w34848 = ~w3242 & ~w33589;
assign w34849 = ~w33731 & w42867;
assign w34850 = ~w34847 & ~w34849;
assign w34851 = ~w34728 & w34850;
assign w34852 = w34727 & ~w34851;
assign w34853 = w34701 & ~w34852;
assign w34854 = ~w34853 & w42868;
assign w34855 = ~w34841 & ~w34845;
assign w34856 = ~w34854 & w34855;
assign w34857 = w34628 & ~w34830;
assign w34858 = ~w34821 & w34857;
assign w34859 = w34856 & w34858;
assign w34860 = ~w945 & ~w34822;
assign w34861 = ~w33735 & ~w34822;
assign w34862 = (~w34860 & w33745) | (~w34860 & w42869) | (w33745 & w42869);
assign w34863 = w945 & ~w33746;
assign w34864 = ~w34828 & ~w34862;
assign w34865 = ~w1120 & ~w34863;
assign w34866 = ~w34864 & ~w34865;
assign w34867 = w34628 & w34866;
assign w34868 = w34608 & ~w34867;
assign w34869 = ~w34665 & w34868;
assign w34870 = ~w34859 & w34869;
assign w34871 = (w34664 & w34859) | (w34664 & w49724) | (w34859 & w49724);
assign w34872 = ~w33550 & w33731;
assign w34873 = ~w33731 & w34559;
assign w34874 = ~w34872 & ~w34873;
assign w34875 = w9781 & ~w34874;
assign w34876 = w34569 & w34875;
assign w34877 = ~w34536 & ~w34876;
assign w34878 = ~w34876 & w42870;
assign w34879 = w34574 & ~w34878;
assign w34880 = w34462 & ~w34879;
assign w34881 = ~w34582 & ~w34880;
assign w34882 = ~w34852 & w42871;
assign w34883 = w34821 & ~w34882;
assign w34884 = ~w34830 & ~w34845;
assign w34885 = ~w34841 & w34884;
assign w34886 = w34608 & ~w34866;
assign w34887 = ~w34665 & w34886;
assign w34888 = (w34887 & w34883) | (w34887 & w49725) | (w34883 & w49725);
assign w34889 = ~w34881 & ~w34888;
assign w34890 = ~w33765 & ~w33773;
assign w34891 = w33784 & ~w34890;
assign w34892 = w33834 & ~w34891;
assign w34893 = ~w33765 & ~w33786;
assign w34894 = (w33784 & w33786) | (w33784 & w49726) | (w33786 & w49726);
assign w34895 = ~w34892 & w34894;
assign w34896 = w34664 & ~w34895;
assign w34897 = (w34896 & w34889) | (w34896 & w47994) | (w34889 & w47994);
assign w34898 = ~w34319 & w49727;
assign w34899 = w34897 & ~w34898;
assign w34900 = (~w33855 & w34898) | (~w33855 & w47995) | (w34898 & w47995);
assign w34901 = w1120 & ~w34829;
assign w34902 = ~w34575 & w42872;
assign w34903 = ~w34319 & w34902;
assign w34904 = w34821 & w34881;
assign w34905 = ~w34903 & ~w34904;
assign w34906 = ~w34830 & w34856;
assign w34907 = ~w34903 & w42873;
assign w34908 = ~w34901 & ~w34907;
assign w34909 = ~w34638 & ~w34863;
assign w34910 = w34908 & ~w34909;
assign w34911 = ~w34908 & w34909;
assign w34912 = ~w33746 & w34900;
assign w34913 = ~w34910 & ~w34911;
assign w34914 = ~w34900 & w34913;
assign w34915 = ~w34912 & ~w34914;
assign w34916 = ~w34881 & w34995;
assign w34917 = ~w34591 & w34916;
assign w34918 = ~w33855 & ~w34871;
assign w34919 = (w34918 & w34591) | (w34918 & w49728) | (w34591 & w49728);
assign w34920 = (~w34591 & w49729) | (~w34591 & w49730) | (w49729 & w49730);
assign w34921 = (~w33954 & w33924) | (~w33954 & w49731) | (w33924 & w49731);
assign w34922 = ~w33956 & w34921;
assign w34923 = w34920 & w34922;
assign w34924 = ~w33924 & w33961;
assign w34925 = w33956 & w34924;
assign w34926 = (w34925 & w42875) | (w34925 & w34899) | (w42875 & w34899);
assign w34927 = w28077 & w34922;
assign w34928 = w33954 & w34924;
assign w34929 = ~w34927 & ~w34928;
assign w34930 = ~w33855 & ~w33953;
assign w34931 = (w34930 & w34898) | (w34930 & w47996) | (w34898 & w47996);
assign w34932 = w34929 & ~w34931;
assign w34933 = ~w34923 & ~w34926;
assign w34934 = w34932 & w34933;
assign w34935 = ~w33935 & ~w33936;
assign w34936 = w34921 & ~w34935;
assign w34937 = ~w34921 & w34935;
assign w34938 = ~w34936 & ~w34937;
assign w34939 = w25851 & w33934;
assign w34940 = (w42876 & w34898) | (w42876 & w47997) | (w34898 & w47997);
assign w34941 = w25851 & ~w34938;
assign w34942 = (w34941 & w42877) | (w34941 & w34899) | (w42877 & w34899);
assign w34943 = ~w34940 & ~w34942;
assign w34944 = w34933 & w47998;
assign w34945 = w34943 & ~w34944;
assign w34946 = ~w33966 & ~w34937;
assign w34947 = w25851 & w34946;
assign w34948 = ~w25851 & ~w34946;
assign w34949 = ~w34947 & ~w34948;
assign w34950 = (~w48000 & w49732) | (~w48000 & w49733) | (w49732 & w49733);
assign w34951 = (w48000 & w49734) | (w48000 & w49735) | (w49734 & w49735);
assign w34952 = ~w34950 & ~w34951;
assign w34953 = w24874 & w34952;
assign w34954 = ~w23843 & ~w34953;
assign w34955 = w34945 & w34954;
assign w34956 = (w42879 & w34898) | (w42879 & w48001) | (w34898 & w48001);
assign w34957 = (w34938 & w42880) | (w34938 & w34899) | (w42880 & w34899);
assign w34958 = ~w34956 & ~w34957;
assign w34959 = ~w25851 & ~w34958;
assign w34960 = ~w33094 & w33731;
assign w34961 = ~w33731 & ~w33984;
assign w34962 = ~w34960 & ~w34961;
assign w34963 = w33979 & ~w34948;
assign w34964 = ~w34947 & ~w34963;
assign w34965 = w24874 & ~w34964;
assign w34966 = (~w34965 & w34899) | (~w34965 & w42881) | (w34899 & w42881);
assign w34967 = ~w25851 & w34938;
assign w34968 = w24874 & ~w34967;
assign w34969 = w33979 & w34947;
assign w34970 = ~w34968 & ~w34969;
assign w34971 = ~w34959 & w34962;
assign w34972 = w34966 & ~w34970;
assign w34973 = ~w34971 & ~w34972;
assign w34974 = w26880 & w34943;
assign w34975 = ~w34934 & w34974;
assign w34976 = ~w24874 & ~w34963;
assign w34977 = w34962 & ~w34976;
assign w34978 = w34966 & w34977;
assign w34979 = ~w24874 & w34950;
assign w34980 = ~w34978 & ~w34979;
assign w34981 = ~w34975 & w34980;
assign w34982 = ~w34973 & w34981;
assign w34983 = ~w34947 & w34976;
assign w34984 = (w34899 & w48002) | (w34899 & w48003) | (w48002 & w48003);
assign w34985 = w34962 & ~w34984;
assign w34986 = ~w34962 & w34984;
assign w34987 = ~w34985 & ~w34986;
assign w34988 = ~w34954 & ~w34987;
assign w34989 = ~w34982 & ~w34988;
assign w34990 = ~w32698 & w33731;
assign w34991 = w32698 & ~w33731;
assign w34992 = ~w34990 & ~w34991;
assign w34993 = w33867 & ~w34992;
assign w34994 = (~w34871 & w34591) | (~w34871 & w49736) | (w34591 & w49736);
assign w34995 = w34664 & ~w34888;
assign w34996 = ~w34575 & ~w34582;
assign w34997 = ~a[11] & w33731;
assign w34998 = ~w34893 & w34997;
assign w34999 = (w34994 & w48004) | (w34994 & w48005) | (w48004 & w48005);
assign w35000 = ~a[11] & ~w34993;
assign w35001 = ~w34999 & ~w35000;
assign w35002 = ~w34892 & ~w34893;
assign w35003 = ~a[10] & ~w33731;
assign w35004 = (~w34591 & w49737) | (~w34591 & w49738) | (w49737 & w49738);
assign w35005 = ~w33867 & w34992;
assign w35006 = (~w35003 & ~w35004) | (~w35003 & w48006) | (~w35004 & w48006);
assign w35007 = w33852 & ~w34893;
assign w35008 = (w48007 & w34591) | (w48007 & w49739) | (w34591 & w49739);
assign w35009 = ~w32698 & ~w33866;
assign w35010 = w35003 & ~w35009;
assign w35011 = ~w35002 & w35010;
assign w35012 = ~w35008 & w35011;
assign w35013 = ~w35006 & ~w35012;
assign w35014 = ~w34993 & ~w35005;
assign w35015 = (~w35014 & w34920) | (~w35014 & w48008) | (w34920 & w48008);
assign w35016 = ~w33855 & w35003;
assign w35017 = ~w35004 & w35016;
assign w35018 = ~w35015 & ~w35017;
assign w35019 = ~w35001 & ~w35013;
assign w35020 = a[11] & ~w35018;
assign w35021 = ~w35019 & ~w35020;
assign w35022 = (w34917 & w49252) | (w34917 & w49253) | (w49252 & w49253);
assign w35023 = ~a[6] & ~a[7];
assign w35024 = ~a[8] & w35023;
assign w35025 = w33731 & ~w35024;
assign w35026 = (~w34898 & w48009) | (~w34898 & w48010) | (w48009 & w48010);
assign w35027 = ~w33731 & w35024;
assign w35028 = a[9] & ~w35025;
assign w35029 = ~w34895 & w35028;
assign w35030 = ~w35027 & w52277;
assign w35031 = ~w35022 & w35026;
assign w35032 = w35030 & ~w35031;
assign w35033 = a[10] & ~w33866;
assign w35034 = ~w33867 & ~w35033;
assign w35035 = ~w34895 & w35034;
assign w35036 = w34995 & w35035;
assign w35037 = (w35036 & w34917) | (w35036 & w42885) | (w34917 & w42885);
assign w35038 = a[10] & w33731;
assign w35039 = ~w35003 & ~w35038;
assign w35040 = (w42886 & w34591) | (w42886 & w49740) | (w34591 & w49740);
assign w35041 = w34895 & w35039;
assign w35042 = ~w33854 & ~w34895;
assign w35043 = w35034 & w35042;
assign w35044 = ~w35041 & ~w35043;
assign w35045 = ~w35037 & ~w35040;
assign w35046 = w35044 & w35045;
assign w35047 = (w35037 & w49741) | (w35037 & w49742) | (w49741 & w49742);
assign w35048 = ~w35037 & w49743;
assign w35049 = ~w31477 & ~w35048;
assign w35050 = w35032 & ~w35047;
assign w35051 = w35049 & ~w35050;
assign w35052 = w35021 & ~w35051;
assign w35053 = w31477 & ~w35047;
assign w35054 = ~w35032 & ~w35048;
assign w35055 = w35053 & ~w35054;
assign w35056 = ~w33855 & ~w34995;
assign w35057 = ~w34895 & ~w35056;
assign w35058 = ~w33731 & w33857;
assign w35059 = w33731 & w33860;
assign w35060 = ~w35058 & ~w35059;
assign w35061 = (w35060 & w34919) | (w35060 & w48014) | (w34919 & w48014);
assign w35062 = ~w31477 & w33876;
assign w35063 = w31477 & ~w33876;
assign w35064 = ~w35062 & ~w35063;
assign w35065 = w35004 & ~w35056;
assign w35066 = w35060 & w35064;
assign w35067 = ~w35060 & ~w35064;
assign w35068 = w35004 & w48015;
assign w35069 = ~w35066 & ~w35068;
assign w35070 = ~w35061 & w35069;
assign w35071 = w30239 & ~w35070;
assign w35072 = ~w35055 & ~w35071;
assign w35073 = ~w35052 & w35072;
assign w35074 = (w42887 & w34898) | (w42887 & w48016) | (w34898 & w48016);
assign w35075 = ~w33916 & w33961;
assign w35076 = ~w33910 & ~w33922;
assign w35077 = ~w35075 & ~w35076;
assign w35078 = w35075 & w35076;
assign w35079 = ~w35077 & ~w35078;
assign w35080 = (w35079 & w35004) | (w35079 & w48017) | (w35004 & w48017);
assign w35081 = ~w35074 & ~w35080;
assign w35082 = w28077 & ~w35081;
assign w35083 = ~w30239 & ~w35061;
assign w35084 = w35069 & w35083;
assign w35085 = w33886 & ~w33922;
assign w35086 = (~w33909 & w34919) | (~w33909 & w48018) | (w34919 & w48018);
assign w35087 = ~w29158 & ~w35086;
assign w35088 = w33909 & w35085;
assign w35089 = w35065 & w35088;
assign w35090 = w35087 & ~w35089;
assign w35091 = ~w35084 & ~w35090;
assign w35092 = ~w35082 & w35091;
assign w35093 = ~w35073 & w35092;
assign w35094 = (w33909 & w34919) | (w33909 & w48019) | (w34919 & w48019);
assign w35095 = w33910 & ~w33922;
assign w35096 = ~w35056 & w35095;
assign w35097 = w35004 & w35096;
assign w35098 = (w29158 & ~w35004) | (w29158 & w48020) | (~w35004 & w48020);
assign w35099 = ~w35094 & w35098;
assign w35100 = (~w48016 & w49744) | (~w48016 & w49745) | (w49744 & w49745);
assign w35101 = ~w35080 & w35100;
assign w35102 = ~w35099 & ~w35101;
assign w35103 = ~w35082 & ~w35102;
assign w35104 = ~w34955 & ~w34989;
assign w35105 = (~w35103 & w34982) | (~w35103 & w48021) | (w34982 & w48021);
assign w35106 = ~w35093 & w35105;
assign w35107 = ~w35104 & ~w35106;
assign w35108 = (~w34959 & w34934) | (~w34959 & w48022) | (w34934 & w48022);
assign w35109 = ~w35103 & w35108;
assign w35110 = w23843 & w34952;
assign w35111 = w35108 & w49746;
assign w35112 = (w35111 & w35073) | (w35111 & w48023) | (w35073 & w48023);
assign w35113 = ~w34024 & w34125;
assign w35114 = (w47995 & w49747) | (w47995 & w49748) | (w49747 & w49748);
assign w35115 = ~w34966 & ~w35114;
assign w35116 = w34962 & w34984;
assign w35117 = ~w35115 & ~w35116;
assign w35118 = w35113 & ~w35117;
assign w35119 = ~w35113 & w35117;
assign w35120 = ~w35118 & ~w35119;
assign w35121 = w22767 & w35120;
assign w35122 = ~w34945 & ~w34959;
assign w35123 = ~w24874 & ~w35122;
assign w35124 = w35110 & ~w35123;
assign w35125 = ~w35121 & ~w35124;
assign w35126 = ~w35112 & w35125;
assign w35127 = w35107 & w35126;
assign w35128 = w35092 & ~w35122;
assign w35129 = ~w35073 & w35128;
assign w35130 = ~w35109 & ~w35122;
assign w35131 = ~w35073 & w35091;
assign w35132 = w26445 & ~w26880;
assign w35133 = w28077 & w35132;
assign w35134 = w34958 & w35133;
assign w35135 = ~w35099 & w35134;
assign w35136 = (w35135 & w35073) | (w35135 & w48024) | (w35073 & w48024);
assign w35137 = (w26445 & w35109) | (w26445 & w49749) | (w35109 & w49749);
assign w35138 = ~w35129 & w35137;
assign w35139 = ~w35136 & ~w35138;
assign w35140 = w34180 & w34302;
assign w35141 = ~w34168 & w34220;
assign w35142 = ~w33250 & w33731;
assign w35143 = ~w33731 & w34192;
assign w35144 = ~w35142 & ~w35143;
assign w35145 = w16559 & ~w35144;
assign w35146 = ~w34168 & w49750;
assign w35147 = w34298 & ~w35146;
assign w35148 = w35140 & ~w35147;
assign w35149 = ~w35140 & w35147;
assign w35150 = ~w35148 & ~w35149;
assign w35151 = w33259 & w33731;
assign w35152 = ~w33731 & w34175;
assign w35153 = ~w35151 & ~w35152;
assign w35154 = ~w34900 & ~w35150;
assign w35155 = (w47995 & w49751) | (w47995 & w49752) | (w49751 & w49752);
assign w35156 = ~w35154 & ~w35155;
assign w35157 = w14766 & ~w35156;
assign w35158 = w14039 & ~w35157;
assign w35159 = (~w42889 & w46055) | (~w42889 & w46056) | (w46055 & w46056);
assign w35160 = (w34102 & w35159) | (w34102 & w49753) | (w35159 & w49753);
assign w35161 = w20906 & ~w35160;
assign w35162 = ~w20906 & w35160;
assign w35163 = ~w35161 & ~w35162;
assign w35164 = ~w33853 & w34891;
assign w35165 = w20906 & w35164;
assign w35166 = w34048 & ~w35165;
assign w35167 = ~w34048 & ~w35163;
assign w35168 = ~w33855 & ~w34048;
assign w35169 = (~w35167 & w34899) | (~w35167 & w42890) | (w34899 & w42890);
assign w35170 = w35163 & w35166;
assign w35171 = w35004 & w35170;
assign w35172 = w35169 & ~w35171;
assign w35173 = ~w20000 & w35172;
assign w35174 = ~w34103 & w35160;
assign w35175 = ~w34049 & ~w35160;
assign w35176 = ~w20000 & ~w34103;
assign w35177 = ~w35175 & w35176;
assign w35178 = w20000 & ~w34049;
assign w35179 = ~w35174 & w35178;
assign w35180 = ~w35177 & ~w35179;
assign w35181 = ~w34114 & w50223;
assign w35182 = w34114 & ~w35180;
assign w35183 = ~w34919 & w48025;
assign w35184 = (w34919 & w48026) | (w34919 & w48027) | (w48026 & w48027);
assign w35185 = ~w35181 & w35184;
assign w35186 = ~w35173 & ~w35185;
assign w35187 = ~w34895 & w35160;
assign w35188 = ~w34024 & ~w35159;
assign w35189 = ~w34098 & ~w35188;
assign w35190 = w34038 & ~w35189;
assign w35191 = ~w34013 & w35187;
assign w35192 = w35187 & w35190;
assign w35193 = (~w35191 & w35056) | (~w35191 & w48028) | (w35056 & w48028);
assign w35194 = ~w21801 & ~w35190;
assign w35195 = ~w34099 & ~w35194;
assign w35196 = w21801 & w35190;
assign w35197 = w35195 & ~w35196;
assign w35198 = ~w33855 & ~w34099;
assign w35199 = (w35198 & w34898) | (w35198 & w48029) | (w34898 & w48029);
assign w35200 = ~w35197 & ~w35199;
assign w35201 = w35200 & w42893;
assign w35202 = w20000 & ~w35172;
assign w35203 = ~w35201 & ~w35202;
assign w35204 = w35186 & ~w35203;
assign w35205 = ~w34060 & ~w34163;
assign w35206 = w34116 & ~w35175;
assign w35207 = w34089 & ~w35206;
assign w35208 = w35205 & ~w35207;
assign w35209 = ~w35205 & w35207;
assign w35210 = ~w35208 & ~w35209;
assign w35211 = ~w33855 & w50224;
assign w35212 = ~w34900 & ~w35210;
assign w35213 = ~w35211 & ~w35212;
assign w35214 = w18183 & w35213;
assign w35215 = ~w35181 & ~w35183;
assign w35216 = w19040 & ~w35215;
assign w35217 = ~w35214 & ~w35216;
assign w35218 = ~w35204 & w35217;
assign w35219 = ~w34134 & ~w34163;
assign w35220 = w34119 & w35219;
assign w35221 = ~w34094 & w35220;
assign w35222 = ~w18183 & ~w35221;
assign w35223 = w18183 & w35221;
assign w35224 = ~w35222 & ~w35223;
assign w35225 = (w35224 & w42894) | (w35224 & w34899) | (w42894 & w34899);
assign w35226 = w34158 & ~w35225;
assign w35227 = ~w34158 & w35225;
assign w35228 = ~w35226 & ~w35227;
assign w35229 = ~w17380 & ~w35228;
assign w35230 = w34298 & ~w35145;
assign w35231 = w35141 & ~w35230;
assign w35232 = ~w35141 & w35230;
assign w35233 = ~w35231 & ~w35232;
assign w35234 = (w42895 & w34898) | (w42895 & w48030) | (w34898 & w48030);
assign w35235 = (w35233 & w34899) | (w35233 & w42896) | (w34899 & w42896);
assign w35236 = ~w35234 & ~w35235;
assign w35237 = (w15681 & w35235) | (w15681 & w48031) | (w35235 & w48031);
assign w35238 = ~w34150 & ~w34161;
assign w35239 = (~w34158 & ~w35221) | (~w34158 & w34159) | (~w35221 & w34159);
assign w35240 = ~w35222 & ~w35239;
assign w35241 = w35238 & ~w35240;
assign w35242 = ~w35238 & w35240;
assign w35243 = ~w35241 & ~w35242;
assign w35244 = ~w34899 & w42897;
assign w35245 = ~w34900 & w35243;
assign w35246 = ~w35244 & ~w35245;
assign w35247 = ~w35245 & w42898;
assign w35248 = ~w35237 & ~w35247;
assign w35249 = ~w35229 & w35248;
assign w35250 = (w20906 & ~w35200) | (w20906 & w42899) | (~w35200 & w42899);
assign w35251 = w34038 & ~w34098;
assign w35252 = w35188 & ~w35251;
assign w35253 = ~w35188 & w35251;
assign w35254 = ~w35252 & ~w35253;
assign w35255 = (w42900 & w34898) | (w42900 & w48032) | (w34898 & w48032);
assign w35256 = (w35254 & w42901) | (w35254 & w34899) | (w42901 & w34899);
assign w35257 = ~w35255 & ~w35256;
assign w35258 = ~w21801 & w35257;
assign w35259 = ~w35250 & ~w35258;
assign w35260 = w35186 & w35259;
assign w35261 = w35249 & ~w35260;
assign w35262 = w35218 & w35261;
assign w35263 = (~w18183 & w35212) | (~w18183 & w49755) | (w35212 & w49755);
assign w35264 = w17380 & w35228;
assign w35265 = ~w35263 & ~w35264;
assign w35266 = w35249 & ~w35265;
assign w35267 = ~w35262 & ~w35266;
assign w35268 = ~w35154 & w49756;
assign w35269 = ~w35235 & w48033;
assign w35270 = (~w16559 & w35245) | (~w16559 & w42902) | (w35245 & w42902);
assign w35271 = (~w35237 & w35270) | (~w35237 & w50137) | (w35270 & w50137);
assign w35272 = ~w35268 & ~w35271;
assign w35273 = ~w35262 & w48034;
assign w35274 = w35158 & ~w35273;
assign w35275 = w35139 & ~w35274;
assign w35276 = ~w22767 & ~w35120;
assign w35277 = w21801 & ~w35257;
assign w35278 = ~w35276 & ~w35277;
assign w35279 = w35218 & w35278;
assign w35280 = ~w35249 & ~w35271;
assign w35281 = w35279 & ~w35280;
assign w35282 = w35273 & ~w35281;
assign w35283 = w35158 & ~w35282;
assign w35284 = w35127 & w35275;
assign w35285 = w35283 & ~w35284;
assign w35286 = ~w34275 & ~w34308;
assign w35287 = ~w34268 & ~w34276;
assign w35288 = w34304 & ~w35141;
assign w35289 = w35287 & ~w35288;
assign w35290 = w14039 & w34900;
assign w35291 = ~w34900 & w35289;
assign w35292 = ~w35290 & ~w35291;
assign w35293 = w35286 & w35292;
assign w35294 = ~w35286 & ~w35292;
assign w35295 = ~w35293 & ~w35294;
assign w35296 = ~w13384 & ~w35295;
assign w35297 = (~w35296 & w35284) | (~w35296 & w48035) | (w35284 & w48035);
assign w35298 = ~w14039 & ~w35268;
assign w35299 = ~w35271 & w35298;
assign w35300 = ~w34267 & ~w34276;
assign w35301 = w34180 & ~w35147;
assign w35302 = w34302 & ~w35301;
assign w35303 = w35300 & ~w35302;
assign w35304 = ~w35300 & w35302;
assign w35305 = w34266 & w34900;
assign w35306 = ~w34900 & ~w35303;
assign w35307 = ~w35304 & w35306;
assign w35308 = ~w35305 & ~w35307;
assign w35309 = ~w14039 & w14766;
assign w35310 = ~w35156 & w35309;
assign w35311 = ~w35308 & ~w35310;
assign w35312 = (w35311 & w35262) | (w35311 & w48036) | (w35262 & w48036);
assign w35313 = ~w34237 & ~w34306;
assign w35314 = ~w34305 & ~w34308;
assign w35315 = (w35314 & w34168) | (w35314 & w48037) | (w34168 & w48037);
assign w35316 = w35313 & ~w35315;
assign w35317 = ~w35313 & w35315;
assign w35318 = ~w35316 & ~w35317;
assign w35319 = ~w34236 & w34900;
assign w35320 = ~w34900 & w35318;
assign w35321 = ~w35319 & ~w35320;
assign w35322 = w12666 & ~w35321;
assign w35323 = ~w35312 & ~w35322;
assign w35324 = w35281 & w35311;
assign w35325 = w35323 & ~w35324;
assign w35326 = w35139 & w35323;
assign w35327 = w35127 & w35326;
assign w35328 = ~w35325 & ~w35327;
assign w35329 = ~w34430 & ~w34431;
assign w35330 = (~w34588 & w34283) | (~w34588 & w42903) | (w34283 & w42903);
assign w35331 = (~w34283 & w48038) | (~w34283 & w48039) | (w48038 & w48039);
assign w35332 = ~w34390 & ~w34409;
assign w35333 = (w34283 & w49757) | (w34283 & w49758) | (w49757 & w49758);
assign w35334 = w35332 & ~w35333;
assign w35335 = ~w34422 & w35334;
assign w35336 = w34414 & ~w34576;
assign w35337 = ~w35335 & w35336;
assign w35338 = w34402 & ~w34450;
assign w35339 = ~w35337 & w35338;
assign w35340 = ~w34577 & ~w35339;
assign w35341 = ~w4056 & w34402;
assign w35342 = ~w35337 & w35341;
assign w35343 = w35340 & ~w35342;
assign w35344 = w35329 & ~w35343;
assign w35345 = w34402 & ~w35337;
assign w35346 = ~w3242 & ~w35329;
assign w35347 = w34450 & w34900;
assign w35348 = ~w35346 & ~w35347;
assign w35349 = w34451 & ~w35345;
assign w35350 = w35348 & ~w35349;
assign w35351 = w3242 & w35329;
assign w35352 = w35340 & ~w35351;
assign w35353 = w34900 & ~w35352;
assign w35354 = ~w3242 & w35329;
assign w35355 = w34451 & w35351;
assign w35356 = ~w3646 & ~w35355;
assign w35357 = ~w34450 & ~w35354;
assign w35358 = w35342 & w35357;
assign w35359 = w35356 & ~w35358;
assign w35360 = ~w35353 & w35359;
assign w35361 = ~w35344 & w35350;
assign w35362 = w35360 & ~w35361;
assign w35363 = ~w34900 & ~w35342;
assign w35364 = w35340 & w35363;
assign w35365 = (~w47995 & w49759) | (~w47995 & w49760) | (w49759 & w49760);
assign w35366 = w35329 & ~w35365;
assign w35367 = ~w35329 & w35365;
assign w35368 = ~w35366 & ~w35367;
assign w35369 = w35346 & w35368;
assign w35370 = ~w35364 & w35369;
assign w35371 = (~w34881 & w34319) | (~w34881 & w42904) | (w34319 & w42904);
assign w35372 = w34740 & w34850;
assign w35373 = w35371 & ~w35372;
assign w35374 = ~w35371 & w35372;
assign w35375 = ~w35373 & ~w35374;
assign w35376 = w33589 & ~w34735;
assign w35377 = ~w33589 & w34735;
assign w35378 = ~w35376 & ~w35377;
assign w35379 = ~w34900 & ~w35375;
assign w35380 = w34900 & w35378;
assign w35381 = ~w35379 & ~w35380;
assign w35382 = w2896 & w35381;
assign w35383 = w35354 & ~w35365;
assign w35384 = w35364 & w35383;
assign w35385 = ~w35382 & ~w35384;
assign w35386 = ~w35370 & w35385;
assign w35387 = ~w35362 & w35386;
assign w35388 = w4056 & ~w35345;
assign w35389 = w35363 & ~w35388;
assign w35390 = w34450 & ~w35389;
assign w35391 = ~w34450 & w35389;
assign w35392 = ~w35390 & ~w35391;
assign w35393 = ~w34900 & ~w35339;
assign w35394 = ~w34450 & ~w35393;
assign w35395 = w35354 & ~w35394;
assign w35396 = w35346 & ~w35393;
assign w35397 = w3646 & ~w35396;
assign w35398 = ~w35395 & w35397;
assign w35399 = w35392 & w35398;
assign w35400 = ~w2896 & ~w35381;
assign w35401 = w3242 & ~w35368;
assign w35402 = ~w35364 & w35401;
assign w35403 = w3242 & w35368;
assign w35404 = w35364 & w35403;
assign w35405 = ~w35402 & ~w35404;
assign w35406 = ~w35400 & w35405;
assign w35407 = ~w35399 & w35406;
assign w35408 = ~w35382 & ~w35407;
assign w35409 = ~w35387 & ~w35408;
assign w35410 = ~w34544 & ~w34572;
assign w35411 = w34569 & w35330;
assign w35412 = w34877 & ~w35411;
assign w35413 = (w35412 & w34899) | (w35412 & w42906) | (w34899 & w42906);
assign w35414 = (w35410 & w35413) | (w35410 & w48041) | (w35413 & w48041);
assign w35415 = ~w35413 & w48042;
assign w35416 = ~w35414 & ~w35415;
assign w35417 = ~w6769 & ~w35416;
assign w35418 = w9916 & ~w34874;
assign w35419 = ~w34293 & ~w35418;
assign w35420 = ~w34316 & w42907;
assign w35421 = w34564 & ~w34588;
assign w35422 = ~w34875 & ~w35421;
assign w35423 = ~w9195 & ~w35422;
assign w35424 = (w35423 & w34283) | (w35423 & w42908) | (w34283 & w42908);
assign w35425 = w9195 & ~w34875;
assign w35426 = ~w34293 & w35425;
assign w35427 = ~w34316 & w42909;
assign w35428 = ~w34283 & w35427;
assign w35429 = ~w33731 & w34547;
assign w35430 = ~w34500 & ~w35429;
assign w35431 = w34500 & w35429;
assign w35432 = ~w35430 & ~w35431;
assign w35433 = w9195 & w35422;
assign w35434 = w35432 & ~w35433;
assign w35435 = ~w35428 & w35434;
assign w35436 = (w8666 & w35435) | (w8666 & w42910) | (w35435 & w42910);
assign w35437 = (~w35436 & w34899) | (~w35436 & w42911) | (w34899 & w42911);
assign w35438 = ~w35435 & w42912;
assign w35439 = w33731 & ~w34510;
assign w35440 = ~w33731 & w34523;
assign w35441 = ~w35439 & ~w35440;
assign w35442 = (~w35441 & ~w42912) | (~w35441 & w46057) | (~w42912 & w46057);
assign w35443 = ~w7924 & w34900;
assign w35444 = (w42911 & w46058) | (w42911 & w46059) | (w46058 & w46059);
assign w35445 = ~w35443 & ~w35444;
assign w35446 = ~w34479 & w34535;
assign w35447 = w7315 & w35446;
assign w35448 = (w35447 & w35444) | (w35447 & w48043) | (w35444 & w48043);
assign w35449 = w7315 & ~w35446;
assign w35450 = ~w35444 & w48044;
assign w35451 = ~w35448 & ~w35450;
assign w35452 = ~w35417 & w35451;
assign w35453 = (~w35433 & w34283) | (~w35433 & w42913) | (w34283 & w42913);
assign w35454 = ~w35424 & w35453;
assign w35455 = ~w33855 & w35454;
assign w35456 = ~w34899 & w35455;
assign w35457 = w35432 & ~w35454;
assign w35458 = ~w35432 & w35454;
assign w35459 = ~w35457 & ~w35458;
assign w35460 = ~w34899 & w42914;
assign w35461 = ~w35456 & w35459;
assign w35462 = ~w35460 & ~w35461;
assign w35463 = (~w8666 & w35461) | (~w8666 & w42915) | (w35461 & w42915);
assign w35464 = ~w35436 & ~w35438;
assign w35465 = ~w34900 & w35464;
assign w35466 = ~w7924 & w35442;
assign w35467 = w35437 & w35466;
assign w35468 = ~w7924 & w35441;
assign w35469 = (w35468 & w34900) | (w35468 & w42916) | (w34900 & w42916);
assign w35470 = ~w35467 & ~w35469;
assign w35471 = ~w35463 & w35470;
assign w35472 = (~w42917 & w46060) | (~w42917 & w46061) | (w46060 & w46061);
assign w35473 = ~w35441 & w35465;
assign w35474 = w35472 & ~w35473;
assign w35475 = ~w35471 & ~w35474;
assign w35476 = ~w7315 & ~w35446;
assign w35477 = ~w35445 & w35476;
assign w35478 = ~w7315 & w35446;
assign w35479 = w35445 & w35478;
assign w35480 = ~w35477 & ~w35479;
assign w35481 = ~w35475 & w35480;
assign w35482 = ~w34293 & ~w34583;
assign w35483 = ~w34283 & w34317;
assign w35484 = ~w34249 & ~w35483;
assign w35485 = w35482 & ~w35484;
assign w35486 = ~w35482 & w35484;
assign w35487 = ~w35485 & ~w35486;
assign w35488 = ~w34899 & w42918;
assign w35489 = ~w34900 & ~w35487;
assign w35490 = ~w35488 & ~w35489;
assign w35491 = ~w35489 & w42919;
assign w35492 = w9781 & ~w35330;
assign w35493 = (w34283 & w48045) | (w34283 & w48046) | (w48045 & w48046);
assign w35494 = ~w35492 & ~w35493;
assign w35495 = (~w35494 & w34899) | (~w35494 & w42920) | (w34899 & w42920);
assign w35496 = w9195 & w34874;
assign w35497 = (~w34899 & w48047) | (~w34899 & w48048) | (w48047 & w48048);
assign w35498 = w9195 & ~w34874;
assign w35499 = (w34899 & w48049) | (w34899 & w48050) | (w48049 & w48050);
assign w35500 = ~w35497 & ~w35499;
assign w35501 = ~w35491 & w35500;
assign w35502 = (w9781 & w35489) | (w9781 & w42921) | (w35489 & w42921);
assign w35503 = ~w34249 & ~w34312;
assign w35504 = (w34311 & w34168) | (w34311 & w42922) | (w34168 & w42922);
assign w35505 = w34239 & w34254;
assign w35506 = ~w35504 & w35505;
assign w35507 = (w34313 & w34168) | (w34313 & w42923) | (w34168 & w42923);
assign w35508 = w34217 & ~w35507;
assign w35509 = ~w35506 & ~w35508;
assign w35510 = w35503 & ~w35509;
assign w35511 = ~w35503 & w35509;
assign w35512 = ~w35510 & ~w35511;
assign w35513 = ~w34899 & w42924;
assign w35514 = ~w34900 & ~w35512;
assign w35515 = ~w35513 & ~w35514;
assign w35516 = (~w10419 & w35514) | (~w10419 & w42925) | (w35514 & w42925);
assign w35517 = ~w35502 & w35516;
assign w35518 = w35501 & ~w35517;
assign w35519 = ~w35461 & w42926;
assign w35520 = ~w9195 & ~w34874;
assign w35521 = (~w34899 & w48051) | (~w34899 & w48052) | (w48051 & w48052);
assign w35522 = ~w9195 & w34874;
assign w35523 = (w34899 & w48053) | (w34899 & w48054) | (w48053 & w48054);
assign w35524 = ~w35521 & ~w35523;
assign w35525 = ~w35519 & w35524;
assign w35526 = ~w35474 & w35525;
assign w35527 = ~w35518 & w35526;
assign w35528 = (w35452 & ~w35481) | (w35452 & w46062) | (~w35481 & w46062);
assign w35529 = w34360 & w34388;
assign w35530 = ~w34571 & ~w34572;
assign w35531 = ~w34899 & w42927;
assign w35532 = ~w35331 & w35530;
assign w35533 = (w35532 & w34899) | (w35532 & w42928) | (w34899 & w42928);
assign w35534 = ~w35531 & ~w35533;
assign w35535 = w35529 & ~w35534;
assign w35536 = ~w35529 & w35534;
assign w35537 = ~w35535 & ~w35536;
assign w35538 = ~w6264 & ~w35537;
assign w35539 = w6769 & w35416;
assign w35540 = ~w35538 & ~w35539;
assign w35541 = (~w46062 & w48055) | (~w46062 & w48056) | (w48055 & w48056);
assign w35542 = ~w35514 & w42929;
assign w35543 = ~w35502 & ~w35542;
assign w35544 = w35501 & ~w35543;
assign w35545 = w35526 & ~w35544;
assign w35546 = (w34239 & ~w34311) | (w34239 & w52278) | (~w34311 & w52278);
assign w35547 = ~w11870 & w35546;
assign w35548 = ~w34201 & ~w35507;
assign w35549 = ~w35546 & w35548;
assign w35550 = ~w35547 & ~w35549;
assign w35551 = (~w34899 & w48057) | (~w34899 & w48058) | (w48057 & w48058);
assign w35552 = (w34899 & w48059) | (w34899 & w48060) | (w48059 & w48060);
assign w35553 = ~w35551 & ~w35552;
assign w35554 = ~w11138 & w35553;
assign w35555 = w11138 & ~w35553;
assign w35556 = ~w34225 & ~w34227;
assign w35557 = ~w34237 & ~w35315;
assign w35558 = ~w34306 & ~w35557;
assign w35559 = w35556 & ~w35558;
assign w35560 = ~w35556 & w35558;
assign w35561 = ~w35559 & ~w35560;
assign w35562 = (w47995 & w49761) | (w47995 & w49762) | (w49761 & w49762);
assign w35563 = ~w34900 & w35561;
assign w35564 = ~w35562 & ~w35563;
assign w35565 = (w11870 & w35563) | (w11870 & w49763) | (w35563 & w49763);
assign w35566 = ~w35555 & w35565;
assign w35567 = ~w35554 & ~w35566;
assign w35568 = w35452 & w35567;
assign w35569 = w35481 & ~w35545;
assign w35570 = (w35568 & ~w35481) | (w35568 & w50138) | (~w35481 & w50138);
assign w35571 = w35541 & ~w35570;
assign w35572 = w34402 & w34414;
assign w35573 = ~w34576 & ~w34900;
assign w35574 = ~w35335 & w35573;
assign w35575 = w4430 & w34900;
assign w35576 = ~w35574 & ~w35575;
assign w35577 = w35572 & ~w35576;
assign w35578 = ~w35572 & w35576;
assign w35579 = ~w35577 & ~w35578;
assign w35580 = w34330 & ~w34378;
assign w35581 = w34388 & w34878;
assign w35582 = w35581 & ~w35330;
assign w35583 = w34388 & ~w35530;
assign w35584 = w34360 & ~w35583;
assign w35585 = w34365 & w35584;
assign w35586 = ~w35582 & w35585;
assign w35587 = w34342 & ~w35586;
assign w35588 = ~w34900 & w35587;
assign w35589 = ~w35588 & w42931;
assign w35590 = (~w35580 & w35588) | (~w35580 & w42932) | (w35588 & w42932);
assign w35591 = ~w35589 & ~w35590;
assign w35592 = ~w5330 & ~w35591;
assign w35593 = w33449 & w33731;
assign w35594 = ~w33731 & w34337;
assign w35595 = ~w35593 & ~w35594;
assign w35596 = w34342 & w35586;
assign w35597 = w34342 & w34365;
assign w35598 = ~w35582 & w35584;
assign w35599 = ~w35597 & ~w35598;
assign w35600 = w34900 & ~w35595;
assign w35601 = ~w34900 & w49764;
assign w35602 = ~w35600 & ~w35601;
assign w35603 = ~w5745 & ~w35602;
assign w35604 = w5330 & w35591;
assign w35605 = w6264 & w35537;
assign w35606 = ~w35604 & ~w35605;
assign w35607 = ~w35592 & w35603;
assign w35608 = w35606 & ~w35607;
assign w35609 = ~w35579 & w35608;
assign w35610 = (w35609 & ~w35541) | (w35609 & w50139) | (~w35541 & w50139);
assign w35611 = ~w35409 & w35610;
assign w35612 = (w35611 & w35327) | (w35611 & w48061) | (w35327 & w48061);
assign w35613 = w35297 & w35612;
assign w35614 = w13384 & w35295;
assign w35615 = ~w12666 & w35321;
assign w35616 = ~w35322 & ~w35615;
assign w35617 = ~w35614 & w35616;
assign w35618 = ~w35322 & ~w35617;
assign w35619 = w35609 & w35618;
assign w35620 = ~w35571 & w35619;
assign w35621 = w5745 & w35602;
assign w35622 = ~w35604 & w35621;
assign w35623 = ~w35592 & ~w35622;
assign w35624 = w5372 & w35623;
assign w35625 = ~w35579 & ~w35624;
assign w35626 = w4056 & ~w35625;
assign w35627 = ~w35620 & w35626;
assign w35628 = ~w11870 & w35564;
assign w35629 = ~w35555 & ~w35628;
assign w35630 = ~w35569 & w46063;
assign w35631 = w35541 & ~w35630;
assign w35632 = w35609 & ~w35631;
assign w35633 = (~w35408 & w35631) | (~w35408 & w49765) | (w35631 & w49765);
assign w35634 = (~w35409 & ~w35627) | (~w35409 & w49766) | (~w35627 & w49766);
assign w35635 = ~w4056 & ~w35579;
assign w35636 = ~w35387 & ~w35400;
assign w35637 = w35407 & ~w35635;
assign w35638 = ~w35636 & ~w35637;
assign w35639 = ~w34343 & ~w34378;
assign w35640 = ~w34378 & w35585;
assign w35641 = ~w34374 & ~w34409;
assign w35642 = w34408 & w34900;
assign w35643 = ~w34900 & w42933;
assign w35644 = ~w34900 & w42934;
assign w35645 = ~w35643 & ~w35644;
assign w35646 = ~w35642 & w35645;
assign w35647 = w35645 & w49767;
assign w35648 = ~w35592 & ~w35647;
assign w35649 = ~w35622 & w35648;
assign w35650 = (w35649 & w35569) | (w35649 & w46064) | (w35569 & w46064);
assign w35651 = w35541 & w35650;
assign w35652 = ~w4838 & ~w35646;
assign w35653 = ~w35608 & w35649;
assign w35654 = ~w34422 & ~w34576;
assign w35655 = w4838 & w34900;
assign w35656 = ~w34900 & w35334;
assign w35657 = ~w35655 & ~w35656;
assign w35658 = w35654 & w35657;
assign w35659 = ~w35654 & ~w35657;
assign w35660 = ~w35658 & ~w35659;
assign w35661 = w4430 & w35660;
assign w35662 = ~w35653 & w46065;
assign w35663 = ~w35651 & w35662;
assign w35664 = ~w4430 & ~w35660;
assign w35665 = (~w35664 & w35651) | (~w35664 & w46066) | (w35651 & w46066);
assign w35666 = ~w35653 & w52279;
assign w35667 = ~w35618 & ~w35664;
assign w35668 = ~w35666 & w35667;
assign w35669 = ~w35665 & ~w35668;
assign w35670 = ~w35638 & ~w35669;
assign w35671 = (~w35670 & w35613) | (~w35670 & w46067) | (w35613 & w46067);
assign w35672 = ~w2006 & w33731;
assign w35673 = ~w33731 & w34768;
assign w35674 = ~w35672 & ~w35673;
assign w35675 = w34769 & ~w35674;
assign w35676 = ~w34769 & w35674;
assign w35677 = ~w35675 & ~w35676;
assign w35678 = ~w34774 & ~w34834;
assign w35679 = ~w34716 & ~w34851;
assign w35680 = w34701 & ~w35679;
assign w35681 = w35371 & w35680;
assign w35682 = ~w34743 & w34780;
assign w35683 = ~w34816 & w35682;
assign w35684 = (w35371 & w49768) | (w35371 & w49769) | (w49768 & w49769);
assign w35685 = w35678 & ~w35684;
assign w35686 = ~w35678 & w35684;
assign w35687 = w34900 & ~w35677;
assign w35688 = ~w35685 & ~w35686;
assign w35689 = ~w34900 & w35688;
assign w35690 = ~w35687 & ~w35689;
assign w35691 = ~w1541 & w35690;
assign w35692 = w34680 & ~w34852;
assign w35693 = ~w34742 & w35692;
assign w35694 = (w34591 & w46069) | (w34591 & w46070) | (w46069 & w46070);
assign w35695 = w2006 & w35682;
assign w35696 = ~w35681 & w35695;
assign w35697 = ~w34900 & ~w35696;
assign w35698 = ~w2006 & w34700;
assign w35699 = ~w35694 & w35698;
assign w35700 = (w34835 & ~w35697) | (w34835 & w42936) | (~w35697 & w42936);
assign w35701 = ~w34900 & w46071;
assign w35702 = ~w35700 & ~w35701;
assign w35703 = ~w1738 & ~w35702;
assign w35704 = ~w35691 & ~w35703;
assign w35705 = w34700 & w34780;
assign w35706 = w35705 & w50225;
assign w35707 = (w34591 & w46072) | (w34591 & w46073) | (w46072 & w46073);
assign w35708 = w34694 & ~w34695;
assign w35709 = ~w34694 & w34695;
assign w35710 = ~w35708 & ~w35709;
assign w35711 = ~w34899 & w46074;
assign w35712 = ~w34900 & w42938;
assign w35713 = ~w35711 & ~w35712;
assign w35714 = (~w2006 & w35712) | (~w2006 & w46075) | (w35712 & w46075);
assign w35715 = ~w34716 & w34740;
assign w35716 = ~w35371 & w35715;
assign w35717 = w34680 & w34726;
assign w35718 = ~w35679 & w35717;
assign w35719 = ~w35716 & w35718;
assign w35720 = w34674 & ~w34675;
assign w35721 = ~w34674 & w34675;
assign w35722 = ~w35720 & ~w35721;
assign w35723 = ~w34900 & w35719;
assign w35724 = ~w34899 & w42939;
assign w35725 = ~w35723 & ~w35724;
assign w35726 = ~w34900 & w42940;
assign w35727 = w35725 & ~w35726;
assign w35728 = w35725 & w42941;
assign w35729 = ~w35714 & ~w35728;
assign w35730 = ~w34716 & ~w34728;
assign w35731 = (w35371 & w49770) | (w35371 & w49771) | (w49770 & w49771);
assign w35732 = ~w35730 & w52280;
assign w35733 = ~w34900 & w46077;
assign w35734 = ~w34715 & w34900;
assign w35735 = (~w2558 & ~w34900) | (~w2558 & w46078) | (~w34900 & w46078);
assign w35736 = ~w35733 & w35735;
assign w35737 = (w2285 & ~w35725) | (w2285 & w42942) | (~w35725 & w42942);
assign w35738 = ~w35736 & ~w35737;
assign w35739 = w35729 & ~w35738;
assign w35740 = w2006 & w35713;
assign w35741 = ~w35700 & w46079;
assign w35742 = ~w35740 & ~w35741;
assign w35743 = ~w35739 & w35742;
assign w35744 = ~w35733 & ~w35734;
assign w35745 = w2558 & ~w35744;
assign w35746 = ~w35737 & w35745;
assign w35747 = w35729 & ~w35746;
assign w35748 = w35743 & ~w35747;
assign w35749 = (w35704 & ~w35743) | (w35704 & w46080) | (~w35743 & w46080);
assign w35750 = (~w35312 & ~w35281) | (~w35312 & w46081) | (~w35281 & w46081);
assign w35751 = ~w35138 & w48062;
assign w35752 = (~w35750 & ~w35127) | (~w35750 & w48063) | (~w35127 & w48063);
assign w35753 = ~w35285 & ~w35752;
assign w35754 = w35322 & w35649;
assign w35755 = ~w35296 & w52281;
assign w35756 = ~w35638 & w35665;
assign w35757 = w35755 & ~w35756;
assign w35758 = w35753 & w35757;
assign w35759 = ~w35612 & ~w35634;
assign w35760 = w35758 & ~w35759;
assign w35761 = w35749 & ~w35760;
assign w35762 = ~w35671 & w35761;
assign w35763 = w35704 & ~w35743;
assign w35764 = w1541 & ~w35690;
assign w35765 = ~w34761 & ~w34832;
assign w35766 = ~w1541 & w34900;
assign w35767 = (~w34834 & w34899) | (~w34834 & w46083) | (w34899 & w46083);
assign w35768 = ~w35685 & w35767;
assign w35769 = ~w35766 & ~w35768;
assign w35770 = w35765 & ~w35769;
assign w35771 = ~w35765 & w35769;
assign w35772 = ~w35770 & ~w35771;
assign w35773 = w1320 & ~w35772;
assign w35774 = ~w35764 & ~w35773;
assign w35775 = ~w35763 & w35774;
assign w35776 = ~w34830 & ~w34901;
assign w35777 = w34856 & w34905;
assign w35778 = ~w34900 & w35777;
assign w35779 = (w35776 & w35778) | (w35776 & w46085) | (w35778 & w46085);
assign w35780 = ~w35778 & w46086;
assign w35781 = ~w35779 & ~w35780;
assign w35782 = ~w945 & ~w35781;
assign w35783 = (~w34833 & w34899) | (~w34833 & w42943) | (w34899 & w42943);
assign w35784 = (w35371 & w49772) | (w35371 & w49773) | (w49772 & w49773);
assign w35785 = w35783 & ~w35784;
assign w35786 = w34839 & ~w34845;
assign w35787 = w34845 & w34900;
assign w35788 = w35783 & w46087;
assign w35789 = (w35786 & w34899) | (w35786 & w46088) | (w34899 & w46088);
assign w35790 = ~w35785 & w35789;
assign w35791 = ~w35790 & w46089;
assign w35792 = ~w1120 & ~w35791;
assign w35793 = ~w35782 & ~w35792;
assign w35794 = w945 & w35781;
assign w35795 = w754 & ~w35794;
assign w35796 = ~w35793 & w35795;
assign w35797 = w35775 & ~w35796;
assign w35798 = w35638 & w35775;
assign w35799 = ~w1320 & w35772;
assign w35800 = w1120 & w35791;
assign w35801 = ~w35799 & ~w35800;
assign w35802 = ~w35665 & w35755;
assign w35803 = w35753 & w35802;
assign w35804 = ~w35798 & w35801;
assign w35805 = ~w35669 & w35801;
assign w35806 = ~w35803 & w35805;
assign w35807 = (~w35804 & w35803) | (~w35804 & w46090) | (w35803 & w46090);
assign w35808 = w35793 & w35807;
assign w35809 = w35795 & ~w35808;
assign w35810 = (w35797 & ~w35761) | (w35797 & w46091) | (~w35761 & w46091);
assign w35811 = w35809 & ~w35810;
assign w35812 = (w35775 & ~w35761) | (w35775 & w46092) | (~w35761 & w46092);
assign w35813 = w3 & w34900;
assign w35814 = (w34917 & w49774) | (w34917 & w49775) | (w49774 & w49775);
assign w35815 = ~w33804 & ~w35814;
assign w35816 = w80 & w52282;
assign w35817 = ~w34900 & ~w35816;
assign w35818 = ~w35815 & w35817;
assign w35819 = ~w35813 & ~w35818;
assign w35820 = ~w33773 & ~w33785;
assign w35821 = w35819 & ~w35820;
assign w35822 = ~w35819 & w35820;
assign w35823 = ~w35821 & ~w35822;
assign w35824 = w42 & w35823;
assign w35825 = ~w33759 & ~w33774;
assign w35826 = ~w33773 & ~w35816;
assign w35827 = ~w35815 & w35826;
assign w35828 = ~w33785 & ~w35827;
assign w35829 = ~w33747 & ~w33763;
assign w35830 = w42 & ~w35829;
assign w35831 = ~w35825 & ~w35828;
assign w35832 = w35825 & ~w35830;
assign w35833 = w35828 & w35832;
assign w35834 = ~w35831 & ~w35833;
assign w35835 = ~w35824 & w35834;
assign w35836 = ~w33765 & ~w35835;
assign w35837 = ~w35814 & w35817;
assign w35838 = w33804 & ~w35837;
assign w35839 = ~w33804 & w35837;
assign w35840 = ~w35838 & ~w35839;
assign w35841 = w3 & ~w35840;
assign w35842 = w33820 & ~w33849;
assign w35843 = (w35842 & w34917) | (w35842 & w46094) | (w34917 & w46094);
assign w35844 = ~w34917 & w46095;
assign w35845 = ~w33848 & w34900;
assign w35846 = ~w35843 & ~w35844;
assign w35847 = ~w34900 & w35846;
assign w35848 = ~w35847 & w49776;
assign w35849 = (~w80 & w35847) | (~w80 & w49777) | (w35847 & w49777);
assign w35850 = ~w33845 & ~w34661;
assign w35851 = ~w34660 & ~w34870;
assign w35852 = ~w34660 & ~w34888;
assign w35853 = ~w34662 & w35852;
assign w35854 = (w35853 & w35371) | (w35853 & w49778) | (w35371 & w49778);
assign w35855 = ~w34900 & w35854;
assign w35856 = ~w35855 & w42948;
assign w35857 = (~w35850 & w35855) | (~w35850 & w42949) | (w35855 & w42949);
assign w35858 = ~w35856 & ~w35857;
assign w35859 = w57 & ~w35858;
assign w35860 = (~w35848 & w35859) | (~w35848 & w46096) | (w35859 & w46096);
assign w35861 = ~w35841 & ~w35860;
assign w35862 = ~w34599 & w34634;
assign w35863 = w34657 & ~w34867;
assign w35864 = w34589 & w35863;
assign w35865 = ~w34575 & w35864;
assign w35866 = ~w34859 & w35865;
assign w35867 = w34881 & w42950;
assign w35868 = ~w34319 & w35866;
assign w35869 = w34657 & ~w34866;
assign w35870 = (w35869 & w34883) | (w35869 & w49779) | (w34883 & w49779);
assign w35871 = ~w34649 & w34656;
assign w35872 = w34628 & ~w35871;
assign w35873 = ~w34618 & ~w35872;
assign w35874 = ~w34629 & ~w35873;
assign w35875 = ~w35870 & w35874;
assign w35876 = ~w35868 & w42951;
assign w35877 = ~w35862 & ~w35876;
assign w35878 = ~w34599 & w34659;
assign w35879 = ~w35870 & w35878;
assign w35880 = ~w35868 & w42952;
assign w35881 = (w46098 & ~w42953) | (w46098 & w49780) | (~w42953 & w49780);
assign w35882 = ~w34618 & ~w34629;
assign w35883 = (~w34898 & w48064) | (~w34898 & w48065) | (w48064 & w48065);
assign w35884 = (~w34917 & w49254) | (~w34917 & w49255) | (w49254 & w49255);
assign w35885 = ~w35883 & ~w35884;
assign w35886 = w34628 & ~w34656;
assign w35887 = ~w34866 & ~w35886;
assign w35888 = (w35887 & w34903) | (w35887 & w46099) | (w34903 & w46099);
assign w35889 = w35872 & ~w35888;
assign w35890 = (w42955 & w34898) | (w42955 & w48066) | (w34898 & w48066);
assign w35891 = ~w35883 & ~w35890;
assign w35892 = (w400 & w35888) | (w400 & w49256) | (w35888 & w49256);
assign w35893 = ~w35885 & w35892;
assign w35894 = ~w35888 & w49257;
assign w35895 = w35891 & w35894;
assign w35896 = ~w35893 & ~w35895;
assign w35897 = (w42953 & w49781) | (w42953 & w49782) | (w49781 & w49782);
assign w35898 = (w42956 & w34898) | (w42956 & w49258) | (w34898 & w49258);
assign w35899 = ~w34599 & ~w35880;
assign w35900 = ~w34900 & w35899;
assign w35901 = ~w35898 & ~w35900;
assign w35902 = ~w34607 & ~w34662;
assign w35903 = w252 & ~w35902;
assign w35904 = ~w35900 & w42957;
assign w35905 = w252 & w35902;
assign w35906 = (w35905 & w35900) | (w35905 & w42958) | (w35900 & w42958);
assign w35907 = ~w35904 & ~w35906;
assign w35908 = ~w35897 & w35907;
assign w35909 = ~w35881 & ~w35896;
assign w35910 = w35908 & ~w35909;
assign w35911 = ~w34648 & ~w34650;
assign w35912 = (~w34866 & w34903) | (~w34866 & w46101) | (w34903 & w46101);
assign w35913 = ~w34638 & ~w35912;
assign w35914 = ~w35911 & w35913;
assign w35915 = w35911 & ~w35913;
assign w35916 = ~w34647 & w34900;
assign w35917 = ~w35914 & ~w35915;
assign w35918 = ~w34900 & w35917;
assign w35919 = ~w35916 & ~w35918;
assign w35920 = ~w612 & w35919;
assign w35921 = (~w34898 & w48067) | (~w34898 & w48068) | (w48067 & w48068);
assign w35922 = w34649 & ~w35912;
assign w35923 = w35921 & ~w35922;
assign w35924 = (w612 & w33854) | (w612 & w49259) | (w33854 & w49259);
assign w35925 = w34628 & w34655;
assign w35926 = (w42960 & w34898) | (w42960 & w48069) | (w34898 & w48069);
assign w35927 = (~w34898 & w48070) | (~w34898 & w48071) | (w48070 & w48071);
assign w35928 = ~w35926 & ~w35927;
assign w35929 = w35923 & ~w35928;
assign w35930 = ~w35923 & w35928;
assign w35931 = ~w35929 & ~w35930;
assign w35932 = ~w493 & ~w35931;
assign w35933 = w35910 & ~w35920;
assign w35934 = ~w35932 & w35933;
assign w35935 = w35861 & w35934;
assign w35936 = ~w35836 & w35935;
assign w35937 = w493 & w35931;
assign w35938 = (w34903 & w49783) | (w34903 & w49784) | (w49783 & w49784);
assign w35939 = ~w35884 & w48072;
assign w35940 = ~w35888 & w42963;
assign w35941 = ~w35891 & w35940;
assign w35942 = ~w35939 & ~w35941;
assign w35943 = ~w35881 & w35942;
assign w35944 = ~w35937 & w35943;
assign w35945 = w35910 & ~w35944;
assign w35946 = ~w57 & w35858;
assign w35947 = ~w35848 & ~w35946;
assign w35948 = ~w35900 & w42964;
assign w35949 = ~w252 & ~w35948;
assign w35950 = ~w35901 & w35902;
assign w35951 = w35949 & ~w35950;
assign w35952 = w35947 & ~w35951;
assign w35953 = ~w35945 & w35952;
assign w35954 = w35861 & ~w35953;
assign w35955 = ~w3 & w35840;
assign w35956 = ~w42 & ~w35823;
assign w35957 = ~w35955 & ~w35956;
assign w35958 = ~w35954 & w35957;
assign w35959 = ~w35836 & ~w35958;
assign w35960 = (w612 & w35918) | (w612 & w42965) | (w35918 & w42965);
assign w35961 = (~w754 & w34914) | (~w754 & w49260) | (w34914 & w49260);
assign w35962 = ~w35794 & ~w35800;
assign w35963 = ~w35960 & w35961;
assign w35964 = w35962 & ~w35963;
assign w35965 = w35793 & w35799;
assign w35966 = w35964 & ~w35965;
assign w35967 = ~w35793 & ~w35794;
assign w35968 = w754 & w34915;
assign w35969 = ~w35960 & ~w35968;
assign w35970 = ~w35793 & w42966;
assign w35971 = w35969 & ~w35970;
assign w35972 = (w35971 & w35775) | (w35971 & w46102) | (w35775 & w46102);
assign w35973 = ~w35959 & w35972;
assign w35974 = w35749 & w35966;
assign w35975 = ~w35638 & w35974;
assign w35976 = ~w35936 & ~w35959;
assign w35977 = w35973 & ~w35975;
assign w35978 = ~w35976 & ~w35977;
assign w35979 = (w35627 & w49785) | (w35627 & w49786) | (w49785 & w49786);
assign w35980 = (~w35978 & w35613) | (~w35978 & w42968) | (w35613 & w42968);
assign w35981 = ~w35664 & w35974;
assign w35982 = ~w35663 & w35981;
assign w35983 = w35973 & ~w35982;
assign w35984 = ~w35618 & w35649;
assign w35985 = (w35984 & w35631) | (w35984 & w46103) | (w35631 & w46103);
assign w35986 = w35981 & w35985;
assign w35987 = w35983 & ~w35986;
assign w35988 = w35973 & w48073;
assign w35989 = w35753 & w35988;
assign w35990 = ~w35987 & ~w35989;
assign w35991 = ~w35634 & w35978;
assign w35992 = ~w35613 & w35991;
assign w35993 = ~w35990 & ~w35992;
assign w35994 = ~w35980 & ~w35993;
assign w35995 = (~w35794 & w35806) | (~w35794 & w42969) | (w35806 & w42969);
assign w35996 = ~w35994 & w35995;
assign w35997 = ~w35812 & w35996;
assign w35998 = ~w754 & ~w35967;
assign w35999 = (~w35998 & w35993) | (~w35998 & w42970) | (w35993 & w42970);
assign w36000 = ~w35997 & ~w35999;
assign w36001 = ~w612 & ~w34915;
assign w36002 = (w36001 & w36000) | (w36001 & w42971) | (w36000 & w42971);
assign w36003 = ~w612 & w34915;
assign w36004 = ~w36000 & w42972;
assign w36005 = ~w36002 & ~w36004;
assign w36006 = w612 & w34915;
assign w36007 = (w36006 & w36000) | (w36006 & w42973) | (w36000 & w42973);
assign w36008 = w612 & ~w34915;
assign w36009 = ~w36000 & w42974;
assign w36010 = ~w36007 & ~w36009;
assign w36011 = w36005 & w36010;
assign w36012 = ~w35993 & w42975;
assign w36013 = ~w35025 & ~w35027;
assign w36014 = ~w34900 & ~w36013;
assign w36015 = w34900 & w36013;
assign w36016 = ~w36014 & ~w36015;
assign w36017 = (~w36016 & w35993) | (~w36016 & w42976) | (w35993 & w42976);
assign w36018 = ~w36012 & ~w36017;
assign w36019 = a[9] & ~w36018;
assign w36020 = w35661 & w35974;
assign w36021 = (~w36020 & w35989) | (~w36020 & w42977) | (w35989 & w42977);
assign w36022 = ~w35980 & ~w36021;
assign w36023 = (w36014 & ~w35991) | (w36014 & w48074) | (~w35991 & w48074);
assign w36024 = ~w36022 & w36023;
assign w36025 = ~w35665 & w35973;
assign w36026 = (w36025 & w35613) | (w36025 & w42978) | (w35613 & w42978);
assign w36027 = (w35668 & ~w35297) | (w35668 & w42979) | (~w35297 & w42979);
assign w36028 = ~w35978 & w36015;
assign w36029 = ~a[9] & ~w36028;
assign w36030 = w36015 & ~w36027;
assign w36031 = w36026 & w36030;
assign w36032 = w36029 & ~w36031;
assign w36033 = ~w36012 & ~w36024;
assign w36034 = w36032 & w36033;
assign w36035 = ~w36019 & ~w36034;
assign w36036 = w32698 & ~w35032;
assign w36037 = ~w32698 & w35032;
assign w36038 = ~w36036 & ~w36037;
assign w36039 = w31477 & w35046;
assign w36040 = w36039 & w52283;
assign w36041 = w31477 & ~w35046;
assign w36042 = (w35993 & w49787) | (w35993 & w49788) | (w49787 & w49788);
assign w36043 = ~w36040 & ~w36042;
assign w36044 = ~a[4] & ~a[5];
assign w36045 = ~a[6] & w36044;
assign w36046 = ~a[7] & w36045;
assign w36047 = ~a[8] & w33731;
assign w36048 = ~a[8] & ~w33731;
assign w36049 = w34900 & ~w36048;
assign w36050 = a[7] & ~w36045;
assign w36051 = a[8] & w33731;
assign w36052 = ~w35024 & ~w36051;
assign w36053 = w36049 & w36050;
assign w36054 = w36052 & ~w36053;
assign w36055 = w36046 & ~w36047;
assign w36056 = ~w34900 & w36055;
assign w36057 = ~w36054 & ~w36056;
assign w36058 = w36046 & ~w36051;
assign w36059 = w36049 & ~w36058;
assign w36060 = ~w34900 & w36047;
assign w36061 = ~w36050 & ~w36060;
assign w36062 = ~w33731 & ~w35022;
assign w36063 = ~w36061 & ~w36062;
assign w36064 = (~w36057 & w35993) | (~w36057 & w42981) | (w35993 & w42981);
assign w36065 = ~w36059 & ~w36063;
assign w36066 = ~w35993 & w42982;
assign w36067 = ~w36064 & ~w36066;
assign w36068 = ~w32698 & w36067;
assign w36069 = w32698 & ~w36067;
assign w36070 = ~w31477 & ~w35046;
assign w36071 = w36070 & w52283;
assign w36072 = ~w31477 & w35046;
assign w36073 = (w35993 & w49789) | (w35993 & w49790) | (w49789 & w49790);
assign w36074 = ~w36071 & ~w36073;
assign w36075 = ~w35051 & ~w35055;
assign w36076 = ~w30239 & ~w35021;
assign w36077 = w36076 & w52284;
assign w36078 = ~w30239 & w35021;
assign w36079 = (w35993 & w49791) | (w35993 & w49792) | (w49791 & w49792);
assign w36080 = ~w36077 & ~w36079;
assign w36081 = w36074 & w36080;
assign w36082 = w36043 & w36069;
assign w36083 = w36081 & ~w36082;
assign w36084 = w36043 & ~w36068;
assign w36085 = ~w36035 & w36084;
assign w36086 = w36083 & ~w36085;
assign w36087 = ~w35073 & ~w35084;
assign w36088 = ~w35094 & ~w35097;
assign w36089 = ~w29158 & ~w36088;
assign w36090 = ~w35992 & w36089;
assign w36091 = ~w36022 & w36090;
assign w36092 = (w36087 & w36091) | (w36087 & w46104) | (w36091 & w46104);
assign w36093 = ~w35099 & ~w36087;
assign w36094 = (w29158 & w35993) | (w29158 & w42984) | (w35993 & w42984);
assign w36095 = ~w36088 & ~w36094;
assign w36096 = (~w36093 & w35993) | (~w36093 & w46105) | (w35993 & w46105);
assign w36097 = ~w36095 & ~w36096;
assign w36098 = ~w36092 & ~w36097;
assign w36099 = (~w28077 & w36097) | (~w28077 & w46106) | (w36097 & w46106);
assign w36100 = ~w35052 & ~w35055;
assign w36101 = ~w30239 & w36100;
assign w36102 = w30239 & ~w36100;
assign w36103 = ~w36101 & ~w36102;
assign w36104 = w35070 & w52285;
assign w36105 = (w35993 & w49793) | (w35993 & w49794) | (w49793 & w49794);
assign w36106 = ~w36104 & ~w36105;
assign w36107 = w29158 & w36106;
assign w36108 = w35021 & w52284;
assign w36109 = (w35993 & w49795) | (w35993 & w49796) | (w49795 & w49796);
assign w36110 = ~w36108 & ~w36109;
assign w36111 = w30239 & ~w36110;
assign w36112 = ~w36107 & ~w36111;
assign w36113 = ~w36099 & w36112;
assign w36114 = ~w36086 & w36113;
assign w36115 = w28077 & w36098;
assign w36116 = ~w29158 & ~w36106;
assign w36117 = ~w36099 & w36116;
assign w36118 = ~w36115 & ~w36117;
assign w36119 = ~w36114 & w36118;
assign w36120 = ~w35093 & ~w35103;
assign w36121 = w26880 & ~w36120;
assign w36122 = ~w26880 & w36120;
assign w36123 = ~w36121 & ~w36122;
assign w36124 = w34934 & w52286;
assign w36125 = (w35993 & w49797) | (w35993 & w49798) | (w49797 & w49798);
assign w36126 = ~w36124 & ~w36125;
assign w36127 = ~w25851 & w36126;
assign w36128 = ~w35082 & ~w35101;
assign w36129 = ~w35993 & w42987;
assign w36130 = ~w35099 & ~w35131;
assign w36131 = (w36130 & w35993) | (w36130 & w42988) | (w35993 & w42988);
assign w36132 = ~w36129 & ~w36131;
assign w36133 = w36128 & w36132;
assign w36134 = ~w36128 & ~w36132;
assign w36135 = ~w36133 & ~w36134;
assign w36136 = w25851 & w34934;
assign w36137 = w36136 & w52286;
assign w36138 = w25851 & ~w34934;
assign w36139 = (w35993 & w49799) | (w35993 & w49800) | (w49799 & w49800);
assign w36140 = ~w36137 & ~w36139;
assign w36141 = w26880 & w36140;
assign w36142 = (~w36127 & ~w36135) | (~w36127 & w49801) | (~w36135 & w49801);
assign w36143 = ~w35129 & w50388;
assign w36144 = (~w24874 & w35129) | (~w24874 & w50389) | (w35129 & w50389);
assign w36145 = ~w36143 & ~w36144;
assign w36146 = w34952 & w52287;
assign w36147 = (w35993 & w49802) | (w35993 & w49803) | (w49802 & w49803);
assign w36148 = ~w36146 & ~w36147;
assign w36149 = w23843 & ~w36148;
assign w36150 = ~w23843 & w36148;
assign w36151 = ~w34934 & ~w36122;
assign w36152 = ~w36121 & ~w36151;
assign w36153 = ~w35993 & w42990;
assign w36154 = (w36152 & w35993) | (w36152 & w42991) | (w35993 & w42991);
assign w36155 = ~w36153 & ~w36154;
assign w36156 = w34943 & ~w34959;
assign w36157 = ~w24874 & ~w36156;
assign w36158 = w36155 & w36157;
assign w36159 = ~w24874 & w36156;
assign w36160 = ~w36155 & w36159;
assign w36161 = ~w36158 & ~w36160;
assign w36162 = (~w36149 & ~w36161) | (~w36149 & w49804) | (~w36161 & w49804);
assign w36163 = w36142 & ~w36162;
assign w36164 = w35127 & w35139;
assign w36165 = ~w35276 & ~w36164;
assign w36166 = ~w35258 & ~w35277;
assign w36167 = w36165 & ~w36166;
assign w36168 = ~w36165 & w36166;
assign w36169 = ~w36167 & ~w36168;
assign w36170 = ~w35993 & w42992;
assign w36171 = (~w36169 & w35993) | (~w36169 & w42993) | (w35993 & w42993);
assign w36172 = ~w36170 & ~w36171;
assign w36173 = ~w20906 & w36172;
assign w36174 = ~w35112 & ~w35124;
assign w36175 = w35139 & w36174;
assign w36176 = w35107 & w36175;
assign w36177 = ~w35121 & ~w35276;
assign w36178 = w36176 & ~w36177;
assign w36179 = ~w36176 & w36177;
assign w36180 = ~w36178 & ~w36179;
assign w36181 = ~w35993 & w42994;
assign w36182 = (~w36180 & w35993) | (~w36180 & w42995) | (w35993 & w42995);
assign w36183 = ~w36181 & ~w36182;
assign w36184 = ~w21801 & w36183;
assign w36185 = w21801 & ~w36183;
assign w36186 = ~w36184 & ~w36185;
assign w36187 = w34952 & ~w36144;
assign w36188 = ~w23843 & ~w36143;
assign w36189 = ~w36187 & w36188;
assign w36190 = w36175 & ~w36189;
assign w36191 = (w36190 & w35993) | (w36190 & w42996) | (w35993 & w42996);
assign w36192 = w22767 & ~w34987;
assign w36193 = w36192 & ~w36191;
assign w36194 = w22767 & w34987;
assign w36195 = (w35993 & w49805) | (w35993 & w49806) | (w49805 & w49806);
assign w36196 = ~w36193 & ~w36195;
assign w36197 = ~w22767 & w34987;
assign w36198 = w36197 & ~w36191;
assign w36199 = ~w22767 & ~w34987;
assign w36200 = (w35993 & w49807) | (w35993 & w49808) | (w49807 & w49808);
assign w36201 = ~w36198 & ~w36200;
assign w36202 = w36196 & w36201;
assign w36203 = w36186 & w36202;
assign w36204 = w36186 & w49809;
assign w36205 = w20906 & ~w36172;
assign w36206 = ~w36184 & w36196;
assign w36207 = ~w36173 & ~w36185;
assign w36208 = ~w36206 & w36207;
assign w36209 = ~w36205 & ~w36208;
assign w36210 = ~w36204 & w36209;
assign w36211 = w36163 & ~w36210;
assign w36212 = (w24874 & ~w36155) | (w24874 & w46107) | (~w36155 & w46107);
assign w36213 = ~w36155 & w36156;
assign w36214 = w36212 & ~w36213;
assign w36215 = ~w36149 & ~w36214;
assign w36216 = ~w26880 & w36128;
assign w36217 = w36132 & w36216;
assign w36218 = w36140 & ~w36217;
assign w36219 = ~w26880 & ~w36128;
assign w36220 = ~w36132 & w36219;
assign w36221 = w36218 & ~w36220;
assign w36222 = ~w36127 & w36161;
assign w36223 = ~w36221 & w36222;
assign w36224 = w36215 & ~w36223;
assign w36225 = w36203 & w46108;
assign w36226 = ~w36224 & w36225;
assign w36227 = ~w35201 & ~w35250;
assign w36228 = ~w35258 & ~w35278;
assign w36229 = w35139 & ~w35258;
assign w36230 = w35127 & w36229;
assign w36231 = ~w36228 & ~w36230;
assign w36232 = w20906 & w35994;
assign w36233 = ~w35994 & w36231;
assign w36234 = ~w36232 & ~w36233;
assign w36235 = w36227 & w36234;
assign w36236 = ~w36227 & ~w36234;
assign w36237 = ~w36235 & ~w36236;
assign w36238 = ~w20000 & ~w36237;
assign w36239 = w36209 & ~w36238;
assign w36240 = ~w36226 & w36239;
assign w36241 = ~w36119 & w36211;
assign w36242 = w36240 & ~w36241;
assign w36243 = w35186 & ~w35250;
assign w36244 = (w36243 & w36230) | (w36243 & w42997) | (w36230 & w42997);
assign w36245 = ~w35214 & ~w35263;
assign w36246 = ~w35204 & ~w35216;
assign w36247 = w36245 & w36246;
assign w36248 = ~w36244 & w36247;
assign w36249 = ~w35229 & ~w35264;
assign w36250 = w35263 & ~w36249;
assign w36251 = ~w35263 & w36249;
assign w36252 = ~w36250 & ~w36251;
assign w36253 = w36248 & w36249;
assign w36254 = ~w36248 & w36252;
assign w36255 = ~w36253 & ~w36254;
assign w36256 = ~w35993 & w42998;
assign w36257 = (w36255 & w35993) | (w36255 & w42999) | (w35993 & w42999);
assign w36258 = ~w36256 & ~w36257;
assign w36259 = ~w16559 & ~w36258;
assign w36260 = ~w35237 & ~w35269;
assign w36261 = ~w35229 & ~w35247;
assign w36262 = ~w35270 & ~w36261;
assign w36263 = (w35279 & ~w35127) | (w35279 & w43000) | (~w35127 & w43000);
assign w36264 = ~w35247 & ~w35270;
assign w36265 = w35218 & ~w35260;
assign w36266 = w35265 & ~w36265;
assign w36267 = w36264 & w36266;
assign w36268 = ~w36263 & w36267;
assign w36269 = ~w36262 & ~w36268;
assign w36270 = w36260 & ~w36269;
assign w36271 = ~w36260 & w36269;
assign w36272 = ~w36270 & ~w36271;
assign w36273 = ~w14766 & w35236;
assign w36274 = ~w35993 & w43001;
assign w36275 = ~w14766 & ~w36272;
assign w36276 = ~w35994 & w36275;
assign w36277 = ~w36274 & ~w36276;
assign w36278 = ~w36263 & w36266;
assign w36279 = ~w35229 & ~w36278;
assign w36280 = w36264 & ~w36279;
assign w36281 = ~w36264 & w36279;
assign w36282 = ~w36280 & ~w36281;
assign w36283 = ~w15681 & ~w35246;
assign w36284 = ~w35993 & w43002;
assign w36285 = ~w15681 & ~w36282;
assign w36286 = ~w35994 & w36285;
assign w36287 = ~w36284 & ~w36286;
assign w36288 = w36277 & w36287;
assign w36289 = ~w36259 & w36288;
assign w36290 = ~w36244 & w36246;
assign w36291 = ~w36245 & ~w36290;
assign w36292 = ~w36248 & ~w36291;
assign w36293 = ~w35993 & w43003;
assign w36294 = (w36292 & w35993) | (w36292 & w43004) | (w35993 & w43004);
assign w36295 = ~w36293 & ~w36294;
assign w36296 = ~w17380 & w36295;
assign w36297 = w17380 & ~w35213;
assign w36298 = ~w35993 & w43005;
assign w36299 = w17380 & w36292;
assign w36300 = ~w35994 & w36299;
assign w36301 = ~w36298 & ~w36300;
assign w36302 = ~w35185 & ~w35216;
assign w36303 = ~w35173 & ~w35203;
assign w36304 = ~w35173 & ~w35250;
assign w36305 = (w36304 & w36230) | (w36304 & w43006) | (w36230 & w43006);
assign w36306 = ~w36303 & ~w36305;
assign w36307 = w36302 & ~w36306;
assign w36308 = ~w36302 & w36306;
assign w36309 = ~w36307 & ~w36308;
assign w36310 = ~w18183 & w35215;
assign w36311 = ~w35993 & w43007;
assign w36312 = ~w18183 & ~w36309;
assign w36313 = ~w35994 & w36312;
assign w36314 = ~w36311 & ~w36313;
assign w36315 = w36301 & w36314;
assign w36316 = ~w36296 & ~w36315;
assign w36317 = w18183 & ~w35215;
assign w36318 = ~w35993 & w43008;
assign w36319 = w18183 & w36309;
assign w36320 = ~w35994 & w36319;
assign w36321 = ~w36318 & ~w36320;
assign w36322 = ~w35173 & ~w35202;
assign w36323 = (~w35250 & w36230) | (~w35250 & w43009) | (w36230 & w43009);
assign w36324 = ~w35201 & ~w36323;
assign w36325 = w36322 & ~w36324;
assign w36326 = ~w36322 & w36324;
assign w36327 = ~w36325 & ~w36326;
assign w36328 = w19040 & ~w35172;
assign w36329 = ~w35993 & w43010;
assign w36330 = w19040 & w36327;
assign w36331 = ~w35994 & w36330;
assign w36332 = ~w36329 & ~w36331;
assign w36333 = w36321 & w36332;
assign w36334 = ~w36296 & w36333;
assign w36335 = ~w36316 & ~w36334;
assign w36336 = w36289 & w36335;
assign w36337 = w36289 & w36315;
assign w36338 = w15681 & w35246;
assign w36339 = ~w35993 & w43011;
assign w36340 = w15681 & w36282;
assign w36341 = ~w35994 & w36340;
assign w36342 = ~w36339 & ~w36341;
assign w36343 = w16559 & ~w35228;
assign w36344 = ~w35993 & w43012;
assign w36345 = w16559 & ~w36255;
assign w36346 = ~w35994 & w36345;
assign w36347 = ~w36344 & ~w36346;
assign w36348 = w36342 & w36347;
assign w36349 = w36288 & ~w36348;
assign w36350 = ~w35993 & w43013;
assign w36351 = (w36272 & w35993) | (w36272 & w43014) | (w35993 & w43014);
assign w36352 = ~w36350 & ~w36351;
assign w36353 = w14766 & ~w36352;
assign w36354 = w35267 & ~w35271;
assign w36355 = w35249 & w36263;
assign w36356 = w36354 & ~w36355;
assign w36357 = ~w14766 & w36356;
assign w36358 = w14766 & ~w36356;
assign w36359 = ~w36357 & ~w36358;
assign w36360 = (~w36359 & w35993) | (~w36359 & w43015) | (w35993 & w43015);
assign w36361 = ~w14039 & ~w35156;
assign w36362 = ~w36360 & w36361;
assign w36363 = ~w14039 & w35156;
assign w36364 = w36360 & w36363;
assign w36365 = ~w36362 & ~w36364;
assign w36366 = ~w36353 & w36365;
assign w36367 = ~w36349 & w36366;
assign w36368 = ~w36337 & w36367;
assign w36369 = ~w36336 & w36368;
assign w36370 = ~w35157 & ~w36356;
assign w36371 = w35298 & ~w36370;
assign w36372 = ~w35285 & ~w36371;
assign w36373 = (w35308 & w35994) | (w35308 & w43016) | (w35994 & w43016);
assign w36374 = ~w35994 & w43017;
assign w36375 = ~w36373 & ~w36374;
assign w36376 = ~w13384 & w36375;
assign w36377 = w35156 & ~w36360;
assign w36378 = ~w35156 & w36360;
assign w36379 = ~w36377 & ~w36378;
assign w36380 = w14039 & ~w36379;
assign w36381 = ~w36376 & ~w36380;
assign w36382 = ~w35172 & w35994;
assign w36383 = ~w35994 & w36327;
assign w36384 = ~w36382 & ~w36383;
assign w36385 = ~w19040 & w36384;
assign w36386 = w36381 & ~w36385;
assign w36387 = ~w36369 & w36386;
assign w36388 = ~w35618 & w35629;
assign w36389 = w35567 & ~w36388;
assign w36390 = (w35567 & w35327) | (w35567 & w50390) | (w35327 & w50390);
assign w36391 = w35297 & w36390;
assign w36392 = w35471 & w35518;
assign w36393 = (w35543 & w36391) | (w35543 & w43018) | (w36391 & w43018);
assign w36394 = w36392 & ~w36393;
assign w36395 = ~w35475 & ~w35526;
assign w36396 = w35451 & ~w36395;
assign w36397 = ~w36394 & w36396;
assign w36398 = (w35480 & w35993) | (w35480 & w43019) | (w35993 & w43019);
assign w36399 = ~w36397 & w36398;
assign w36400 = w35451 & w35480;
assign w36401 = ~w36395 & ~w36400;
assign w36402 = w35445 & ~w35446;
assign w36403 = ~w35445 & w35446;
assign w36404 = ~w36402 & ~w36403;
assign w36405 = ~w35993 & w46109;
assign w36406 = ~w35994 & w43020;
assign w36407 = ~w36405 & ~w36406;
assign w36408 = w36398 & w46110;
assign w36409 = w36407 & ~w36408;
assign w36410 = (w6769 & ~w36407) | (w6769 & w46111) | (~w36407 & w46111);
assign w36411 = w35470 & ~w35474;
assign w36412 = ~w35518 & w35525;
assign w36413 = w35525 & w35543;
assign w36414 = (w36413 & w36391) | (w36413 & w43021) | (w36391 & w43021);
assign w36415 = ~w36412 & ~w36414;
assign w36416 = (w43022 & w35993) | (w43022 & w50391) | (w35993 & w50391);
assign w36417 = ~w35993 & w46112;
assign w36418 = (~w36411 & w36416) | (~w36411 & w46113) | (w36416 & w46113);
assign w36419 = (w35993 & w48075) | (w35993 & w48076) | (w48075 & w48076);
assign w36420 = ~w36416 & w36419;
assign w36421 = (~w7315 & w36416) | (~w7315 & w48077) | (w36416 & w48077);
assign w36422 = ~w36418 & w36421;
assign w36423 = ~w36410 & ~w36422;
assign w36424 = ~w36411 & w36415;
assign w36425 = ~w35993 & w46114;
assign w36426 = (~w35463 & w35993) | (~w35463 & w43024) | (w35993 & w43024);
assign w36427 = w36424 & w36426;
assign w36428 = ~w36425 & ~w36427;
assign w36429 = (w7315 & ~w36428) | (w7315 & w50392) | (~w36428 & w50392);
assign w36430 = ~w35463 & ~w35519;
assign w36431 = w35524 & ~w36430;
assign w36432 = ~w35993 & w46115;
assign w36433 = ~w35994 & w43025;
assign w36434 = ~w36432 & ~w36433;
assign w36435 = ~w35994 & w46116;
assign w36436 = w36434 & ~w36435;
assign w36437 = w36434 & w46117;
assign w36438 = ~w36429 & ~w36437;
assign w36439 = w36423 & ~w36438;
assign w36440 = w36407 & w46118;
assign w36441 = ~w35993 & w46119;
assign w36442 = ~w36399 & ~w36441;
assign w36443 = ~w35417 & ~w35539;
assign w36444 = w6264 & ~w36443;
assign w36445 = (w36444 & w36399) | (w36444 & w46120) | (w36399 & w46120);
assign w36446 = w6264 & w36443;
assign w36447 = ~w36399 & w46121;
assign w36448 = ~w36445 & ~w36447;
assign w36449 = ~w36440 & w36448;
assign w36450 = w34874 & ~w35495;
assign w36451 = ~w34874 & w35495;
assign w36452 = ~w36450 & ~w36451;
assign w36453 = w35994 & w36452;
assign w36454 = w35500 & w35524;
assign w36455 = ~w35516 & ~w36389;
assign w36456 = ~w35491 & ~w35502;
assign w36457 = ~w35542 & w36456;
assign w36458 = (w36457 & w36391) | (w36457 & w43026) | (w36391 & w43026);
assign w36459 = ~w35491 & ~w36458;
assign w36460 = w36454 & w36459;
assign w36461 = ~w36454 & ~w36459;
assign w36462 = ~w35994 & w46122;
assign w36463 = ~w36453 & ~w36462;
assign w36464 = w8666 & ~w36463;
assign w36465 = ~w36437 & ~w36464;
assign w36466 = w36449 & w36465;
assign w36467 = ~w36439 & w36466;
assign w36468 = (~w35542 & w36391) | (~w35542 & w43027) | (w36391 & w43027);
assign w36469 = ~w36456 & ~w36468;
assign w36470 = w35490 & w35994;
assign w36471 = ~w35994 & w43028;
assign w36472 = ~w36470 & ~w36471;
assign w36473 = w9195 & ~w36472;
assign w36474 = ~w8666 & w36463;
assign w36475 = ~w36473 & ~w36474;
assign w36476 = ~w35554 & ~w35555;
assign w36477 = ~w35618 & ~w35628;
assign w36478 = ~w35565 & ~w36477;
assign w36479 = ~w35328 & ~w35565;
assign w36480 = w35297 & w36479;
assign w36481 = (w36476 & w36480) | (w36476 & w43029) | (w36480 & w43029);
assign w36482 = ~w36480 & w43030;
assign w36483 = ~w36481 & ~w36482;
assign w36484 = ~w35993 & w43031;
assign w36485 = ~w35994 & w36483;
assign w36486 = ~w36484 & ~w36485;
assign w36487 = (~w10419 & w36485) | (~w10419 & w43032) | (w36485 & w43032);
assign w36488 = ~w35516 & ~w35542;
assign w36489 = ~w36391 & w43033;
assign w36490 = (w36488 & w36391) | (w36488 & w43034) | (w36391 & w43034);
assign w36491 = ~w35993 & w46123;
assign w36492 = ~w36489 & ~w36490;
assign w36493 = ~w35994 & w36492;
assign w36494 = ~w36491 & ~w36493;
assign w36495 = (~w9781 & w36493) | (~w9781 & w46124) | (w36493 & w46124);
assign w36496 = ~w36487 & ~w36495;
assign w36497 = (~w35618 & ~w35297) | (~w35618 & w43035) | (~w35297 & w43035);
assign w36498 = w35322 & w35614;
assign w36499 = w11870 & w36497;
assign w36500 = ~w11870 & ~w36498;
assign w36501 = ~w36497 & w36500;
assign w36502 = ~w36499 & ~w36501;
assign w36503 = ~w35994 & w36502;
assign w36504 = ~w35296 & ~w35614;
assign w36505 = w35614 & ~w35616;
assign w36506 = ~w35617 & ~w36505;
assign w36507 = w35753 & w43036;
assign w36508 = (w36506 & ~w35753) | (w36506 & w43037) | (~w35753 & w43037);
assign w36509 = ~w36507 & ~w36508;
assign w36510 = ~w11870 & w35321;
assign w36511 = ~w35993 & w43038;
assign w36512 = ~w11870 & w36509;
assign w36513 = ~w35994 & w36512;
assign w36514 = ~w36511 & ~w36513;
assign w36515 = w11138 & ~w35564;
assign w36516 = w36503 & w36515;
assign w36517 = w11138 & w35564;
assign w36518 = (w36517 & w35994) | (w36517 & w43039) | (w35994 & w43039);
assign w36519 = w36514 & ~w36518;
assign w36520 = ~w36516 & w36519;
assign w36521 = w36496 & w36520;
assign w36522 = w35321 & w35994;
assign w36523 = ~w35994 & w36509;
assign w36524 = ~w36522 & ~w36523;
assign w36525 = w11870 & w36524;
assign w36526 = ~w13384 & w35753;
assign w36527 = w13384 & ~w35753;
assign w36528 = ~w36526 & ~w36527;
assign w36529 = (~w36528 & w35993) | (~w36528 & w43040) | (w35993 & w43040);
assign w36530 = w35295 & ~w36529;
assign w36531 = ~w35295 & w36529;
assign w36532 = ~w36530 & ~w36531;
assign w36533 = w12666 & w36532;
assign w36534 = ~w36525 & ~w36533;
assign w36535 = w36521 & ~w36534;
assign w36536 = ~w9195 & w36472;
assign w36537 = w9781 & w36494;
assign w36538 = ~w36536 & ~w36537;
assign w36539 = ~w36485 & w43041;
assign w36540 = ~w11138 & ~w35564;
assign w36541 = (w36540 & w35994) | (w36540 & w43042) | (w35994 & w43042);
assign w36542 = ~w11138 & w35564;
assign w36543 = ~w35994 & w43043;
assign w36544 = ~w36541 & ~w36543;
assign w36545 = ~w36539 & w36544;
assign w36546 = w36496 & ~w36545;
assign w36547 = w36538 & ~w36546;
assign w36548 = ~w36535 & w36547;
assign w36549 = ~w12666 & ~w36532;
assign w36550 = w36520 & w46125;
assign w36551 = w36548 & ~w36550;
assign w36552 = (w36475 & ~w36548) | (w36475 & w43044) | (~w36548 & w43044);
assign w36553 = ~w7924 & ~w36436;
assign w36554 = ~w36429 & w36553;
assign w36555 = w36423 & ~w36554;
assign w36556 = w36449 & ~w36555;
assign w36557 = w13384 & ~w36375;
assign w36558 = ~w36381 & ~w36557;
assign w36559 = ~w36349 & ~w36353;
assign w36560 = w36365 & ~w36557;
assign w36561 = w36559 & w36560;
assign w36562 = ~w36336 & w36561;
assign w36563 = ~w36558 & ~w36562;
assign w36564 = w20000 & w36237;
assign w36565 = w36386 & w36564;
assign w36566 = ~w36369 & w36565;
assign w36567 = ~w36563 & ~w36566;
assign w36568 = ~w36556 & w36567;
assign w36569 = w36467 & ~w36552;
assign w36570 = w36568 & ~w36569;
assign w36571 = w36242 & w36387;
assign w36572 = w36570 & ~w36571;
assign w36573 = (~w36535 & w46126) | (~w36535 & w46127) | (w46126 & w46127);
assign w36574 = w36467 & w36573;
assign w36575 = ~w36556 & ~w36574;
assign w36576 = (~w36575 & ~w36570) | (~w36575 & w43046) | (~w36570 & w43046);
assign w36577 = (~w35799 & w35762) | (~w35799 & w43047) | (w35762 & w43047);
assign w36578 = ~w35792 & ~w35800;
assign w36579 = (~w36578 & w35993) | (~w36578 & w43048) | (w35993 & w43048);
assign w36580 = ~w35993 & w43049;
assign w36581 = ~w36579 & ~w36580;
assign w36582 = ~w35993 & w43050;
assign w36583 = ~w36577 & ~w36581;
assign w36584 = ~w36579 & ~w36582;
assign w36585 = w36577 & w36584;
assign w36586 = ~w36583 & ~w36585;
assign w36587 = ~w945 & w36586;
assign w36588 = (~w35807 & w35762) | (~w35807 & w43051) | (w35762 & w43051);
assign w36589 = ~w35792 & ~w35994;
assign w36590 = ~w36588 & w36589;
assign w36591 = w945 & w35994;
assign w36592 = ~w35782 & ~w35794;
assign w36593 = w754 & ~w36592;
assign w36594 = ~w36591 & w36593;
assign w36595 = ~w36590 & w36594;
assign w36596 = w35793 & w35795;
assign w36597 = ~w35994 & w36596;
assign w36598 = ~w36588 & w36597;
assign w36599 = w754 & ~w35781;
assign w36600 = w36591 & w36599;
assign w36601 = ~w36598 & ~w36600;
assign w36602 = ~w36595 & w36601;
assign w36603 = ~w36587 & w36602;
assign w36604 = ~w35671 & ~w35760;
assign w36605 = ~w35671 & w43052;
assign w36606 = ~w35739 & ~w35740;
assign w36607 = ~w1738 & w35994;
assign w36608 = (w36606 & w35993) | (w36606 & w43053) | (w35993 & w43053);
assign w36609 = ~w36605 & w36608;
assign w36610 = ~w36607 & ~w36609;
assign w36611 = ~w35703 & ~w35741;
assign w36612 = w1541 & w36611;
assign w36613 = ~w36610 & w36612;
assign w36614 = w1541 & ~w36611;
assign w36615 = w36610 & w36614;
assign w36616 = ~w36613 & ~w36615;
assign w36617 = ~w35763 & ~w35764;
assign w36618 = (w36617 & ~w35761) | (w36617 & w46128) | (~w35761 & w46128);
assign w36619 = ~w35994 & w36618;
assign w36620 = ~w35993 & w43054;
assign w36621 = ~w35773 & ~w35799;
assign w36622 = ~w1120 & ~w36621;
assign w36623 = ~w36620 & w36622;
assign w36624 = ~w36619 & w36623;
assign w36625 = ~w35994 & ~w36618;
assign w36626 = ~w35993 & w43055;
assign w36627 = ~w1120 & w36621;
assign w36628 = ~w36626 & w36627;
assign w36629 = ~w36625 & w36628;
assign w36630 = ~w36624 & ~w36629;
assign w36631 = ~w35703 & ~w35748;
assign w36632 = (w36631 & w35993) | (w36631 & w43056) | (w35993 & w43056);
assign w36633 = ~w35669 & ~w35803;
assign w36634 = ~w35653 & ~w35747;
assign w36635 = ~w35651 & w36634;
assign w36636 = ~w35638 & ~w36635;
assign w36637 = w35755 & ~w36636;
assign w36638 = ~w35985 & w36635;
assign w36639 = ~w35638 & ~w36638;
assign w36640 = w35753 & w36637;
assign w36641 = w36639 & ~w36640;
assign w36642 = (w35743 & w35613) | (w35743 & w43057) | (w35613 & w43057);
assign w36643 = w36633 & w36641;
assign w36644 = w36642 & ~w36643;
assign w36645 = w36632 & ~w36644;
assign w36646 = ~w35993 & w43058;
assign w36647 = ~w35691 & ~w35764;
assign w36648 = w1320 & w36647;
assign w36649 = ~w36646 & w36648;
assign w36650 = ~w36645 & w36649;
assign w36651 = w1320 & ~w36647;
assign w36652 = (w36651 & w36643) | (w36651 & w43059) | (w36643 & w43059);
assign w36653 = w36632 & w36652;
assign w36654 = w35764 & w36626;
assign w36655 = ~w36653 & ~w36654;
assign w36656 = ~w36650 & w36655;
assign w36657 = w36630 & w36656;
assign w36658 = w36616 & w36657;
assign w36659 = w36603 & w36658;
assign w36660 = ~w36590 & ~w36591;
assign w36661 = ~w754 & ~w36592;
assign w36662 = ~w36660 & w36661;
assign w36663 = ~w754 & w36592;
assign w36664 = w36660 & w36663;
assign w36665 = ~w36662 & ~w36664;
assign w36666 = ~w35728 & ~w35737;
assign w36667 = ~w35736 & ~w36666;
assign w36668 = ~w35728 & w35978;
assign w36669 = (w36668 & ~w36026) | (w36668 & w46129) | (~w36026 & w46129);
assign w36670 = w36667 & ~w36669;
assign w36671 = ~w35671 & w49261;
assign w36672 = w36670 & ~w36671;
assign w36673 = ~w35728 & ~w35738;
assign w36674 = (~w36673 & w35993) | (~w36673 & w43060) | (w35993 & w43060);
assign w36675 = ~w35728 & ~w35745;
assign w36676 = ~w35671 & w43061;
assign w36677 = w36674 & ~w36676;
assign w36678 = (~w2285 & w35993) | (~w2285 & w43062) | (w35993 & w43062);
assign w36679 = ~w35727 & ~w36678;
assign w36680 = ~w36677 & ~w36679;
assign w36681 = ~w36672 & ~w36680;
assign w36682 = ~w36680 & w46130;
assign w36683 = ~w35993 & w46131;
assign w36684 = ~w36677 & ~w36683;
assign w36685 = ~w35714 & ~w35740;
assign w36686 = w1738 & w36685;
assign w36687 = (w36686 & w36677) | (w36686 & w46132) | (w36677 & w46132);
assign w36688 = w1738 & ~w36685;
assign w36689 = ~w36677 & w46133;
assign w36690 = ~w36687 & ~w36689;
assign w36691 = ~w36682 & w36690;
assign w36692 = ~w35736 & ~w35745;
assign w36693 = ~w35994 & w36604;
assign w36694 = (w36692 & w36693) | (w36692 & w43064) | (w36693 & w43064);
assign w36695 = ~w36693 & w43065;
assign w36696 = ~w36694 & ~w36695;
assign w36697 = ~w2285 & ~w36696;
assign w36698 = (~w2006 & w36680) | (~w2006 & w46134) | (w36680 & w46134);
assign w36699 = ~w36697 & ~w36698;
assign w36700 = w36691 & ~w36699;
assign w36701 = ~w1738 & ~w36685;
assign w36702 = ~w36684 & w36701;
assign w36703 = ~w1738 & w36685;
assign w36704 = w36684 & w36703;
assign w36705 = ~w36702 & ~w36704;
assign w36706 = ~w1541 & ~w36611;
assign w36707 = ~w36610 & w36706;
assign w36708 = ~w1541 & w36611;
assign w36709 = w36610 & w36708;
assign w36710 = ~w36707 & ~w36709;
assign w36711 = w36705 & w36710;
assign w36712 = (w36665 & ~w36658) | (w36665 & w43066) | (~w36658 & w43066);
assign w36713 = w36665 & w36711;
assign w36714 = ~w36700 & w36713;
assign w36715 = ~w36712 & ~w36714;
assign w36716 = w945 & ~w36586;
assign w36717 = ~w1320 & ~w36647;
assign w36718 = ~w36646 & w36717;
assign w36719 = ~w36645 & w36718;
assign w36720 = ~w1320 & w36647;
assign w36721 = w36646 & w36720;
assign w36722 = (w36720 & w36643) | (w36720 & w43067) | (w36643 & w43067);
assign w36723 = w36632 & w36722;
assign w36724 = ~w36721 & ~w36723;
assign w36725 = ~w36719 & w36724;
assign w36726 = w1120 & w36621;
assign w36727 = ~w36620 & w36726;
assign w36728 = ~w36619 & w36727;
assign w36729 = w1120 & ~w36621;
assign w36730 = ~w36626 & w36729;
assign w36731 = ~w36625 & w36730;
assign w36732 = ~w36728 & ~w36731;
assign w36733 = w36725 & w36732;
assign w36734 = w36630 & ~w36733;
assign w36735 = (~w36716 & w36733) | (~w36716 & w43068) | (w36733 & w43068);
assign w36736 = w36603 & ~w36735;
assign w36737 = ~w35931 & w35994;
assign w36738 = ~w35920 & w35974;
assign w36739 = ~w35760 & w36738;
assign w36740 = ~w35920 & ~w35972;
assign w36741 = ~w35932 & ~w35937;
assign w36742 = (w43069 & ~w36739) | (w43069 & w46135) | (~w36739 & w46135);
assign w36743 = (w36739 & w46136) | (w36739 & w46137) | (w46136 & w46137);
assign w36744 = ~w36742 & ~w36743;
assign w36745 = ~w35994 & ~w36744;
assign w36746 = (~w36737 & w36744) | (~w36737 & w49262) | (w36744 & w49262);
assign w36747 = w400 & ~w36746;
assign w36748 = ~w35937 & ~w36740;
assign w36749 = (w36739 & w46138) | (w36739 & w46139) | (w46138 & w46139);
assign w36750 = w35896 & w35942;
assign w36751 = (w36750 & w35993) | (w36750 & w43072) | (w35993 & w43072);
assign w36752 = w35885 & ~w35889;
assign w36753 = w35889 & ~w35891;
assign w36754 = ~w36752 & ~w36753;
assign w36755 = ~w35993 & w43073;
assign w36756 = ~w36751 & ~w36755;
assign w36757 = ~w35993 & w43074;
assign w36758 = ~w36751 & ~w36757;
assign w36759 = ~w36749 & w36756;
assign w36760 = w36749 & ~w36758;
assign w36761 = ~w36759 & ~w36760;
assign w36762 = ~w351 & ~w36761;
assign w36763 = w35896 & ~w35932;
assign w36764 = w35942 & ~w36763;
assign w36765 = w35942 & w36748;
assign w36766 = (w36739 & w46140) | (w36739 & w46141) | (w46140 & w46141);
assign w36767 = ~w35881 & ~w35897;
assign w36768 = w400 & w34900;
assign w36769 = ~w34900 & w35876;
assign w36770 = ~w36768 & ~w36769;
assign w36771 = w35862 & w36770;
assign w36772 = ~w35862 & ~w36770;
assign w36773 = ~w36771 & ~w36772;
assign w36774 = w35994 & w36773;
assign w36775 = (~w36767 & w35993) | (~w36767 & w46142) | (w35993 & w46142);
assign w36776 = w36766 & w36775;
assign w36777 = ~w36774 & ~w36776;
assign w36778 = (w36767 & w35993) | (w36767 & w46143) | (w35993 & w46143);
assign w36779 = ~w36766 & w36778;
assign w36780 = (w252 & w36766) | (w252 & w49263) | (w36766 & w49263);
assign w36781 = w36777 & w36780;
assign w36782 = ~w36762 & ~w36781;
assign w36783 = ~w36747 & w36782;
assign w36784 = ~w35993 & w43076;
assign w36785 = ~w34915 & ~w36784;
assign w36786 = ~w35811 & w36785;
assign w36787 = ~w35999 & ~w36784;
assign w36788 = ~w35997 & w36787;
assign w36789 = ~w36786 & ~w36788;
assign w36790 = ~w35920 & ~w35960;
assign w36791 = ~w493 & ~w36790;
assign w36792 = (w36791 & w36788) | (w36791 & w46144) | (w36788 & w46144);
assign w36793 = ~w493 & w36790;
assign w36794 = ~w36788 & w46145;
assign w36795 = ~w36792 & ~w36794;
assign w36796 = w36005 & w36795;
assign w36797 = w36783 & w36796;
assign w36798 = ~w36736 & w36797;
assign w36799 = ~w36715 & w36798;
assign w36800 = w36777 & ~w36779;
assign w36801 = ~w252 & ~w36800;
assign w36802 = w351 & w36761;
assign w36803 = ~w400 & ~w36737;
assign w36804 = ~w36745 & w36803;
assign w36805 = ~w36802 & ~w36804;
assign w36806 = w36782 & ~w36805;
assign w36807 = ~w36801 & ~w36806;
assign w36808 = w493 & w36790;
assign w36809 = (w36808 & w36788) | (w36808 & w46146) | (w36788 & w46146);
assign w36810 = w493 & ~w36790;
assign w36811 = ~w36788 & w46147;
assign w36812 = ~w36809 & ~w36811;
assign w36813 = w36010 & w36812;
assign w36814 = w36795 & ~w36813;
assign w36815 = ~w36813 & w43077;
assign w36816 = w36807 & ~w36815;
assign w36817 = ~w36799 & w36816;
assign w36818 = ~w35328 & w35610;
assign w36819 = w35297 & w36818;
assign w36820 = w35627 & ~w35632;
assign w36821 = ~w36819 & w36820;
assign w36822 = (~w35635 & w35668) | (~w35635 & w43078) | (w35668 & w43078);
assign w36823 = (w36822 & ~w35753) | (w36822 & w46148) | (~w35753 & w46148);
assign w36824 = ~w36821 & ~w36823;
assign w36825 = ~w36821 & w46149;
assign w36826 = ~w35994 & ~w36825;
assign w36827 = ~w3646 & ~w36824;
assign w36828 = (~w36821 & w46150) | (~w36821 & w46151) | (w46150 & w46151);
assign w36829 = ~w35994 & w46152;
assign w36830 = w35364 & ~w35368;
assign w36831 = ~w35364 & w35368;
assign w36832 = ~w36830 & ~w36831;
assign w36833 = ~w3242 & ~w36832;
assign w36834 = w35405 & ~w36833;
assign w36835 = ~w36829 & w43080;
assign w36836 = (w36834 & w36829) | (w36834 & w43081) | (w36829 & w43081);
assign w36837 = ~w36835 & ~w36836;
assign w36838 = w2896 & w36837;
assign w36839 = w36826 & w43082;
assign w36840 = w2896 & ~w36833;
assign w36841 = ~w2896 & w36833;
assign w36842 = ~w36840 & ~w36841;
assign w36843 = (~w36842 & w35993) | (~w36842 & w43083) | (w35993 & w43083);
assign w36844 = w35381 & ~w36843;
assign w36845 = ~w35381 & w36843;
assign w36846 = ~w36844 & ~w36845;
assign w36847 = w36839 & ~w36846;
assign w36848 = ~w36839 & w36846;
assign w36849 = ~w36847 & ~w36848;
assign w36850 = ~w2558 & w36849;
assign w36851 = ~w36838 & ~w36850;
assign w36852 = ~w2896 & ~w36837;
assign w36853 = (w35392 & ~w36826) | (w35392 & w46153) | (~w36826 & w46153);
assign w36854 = w36826 & w46154;
assign w36855 = ~w36853 & ~w36854;
assign w36856 = w3242 & ~w36855;
assign w36857 = ~w36852 & ~w36856;
assign w36858 = w2558 & ~w36849;
assign w36859 = (~w36858 & ~w36851) | (~w36858 & w46155) | (~w36851 & w46155);
assign w36860 = w36442 & ~w36443;
assign w36861 = (w36443 & w36399) | (w36443 & w46156) | (w36399 & w46156);
assign w36862 = ~w36860 & ~w36861;
assign w36863 = (~w6264 & w36860) | (~w6264 & w46157) | (w36860 & w46157);
assign w36864 = ~w35538 & ~w35605;
assign w36865 = ~w35528 & ~w35539;
assign w36866 = w35570 & ~w36388;
assign w36867 = w36865 & ~w36866;
assign w36868 = ~w35328 & w35570;
assign w36869 = w35297 & w36868;
assign w36870 = ~w36869 & w43084;
assign w36871 = (w36864 & w36869) | (w36864 & w43085) | (w36869 & w43085);
assign w36872 = ~w35993 & w46158;
assign w36873 = ~w36870 & ~w36871;
assign w36874 = ~w35994 & w36873;
assign w36875 = ~w36872 & ~w36874;
assign w36876 = w5745 & ~w36875;
assign w36877 = ~w36863 & ~w36876;
assign w36878 = ~w35592 & ~w35604;
assign w36879 = ~w35571 & ~w35605;
assign w36880 = ~w35603 & w36879;
assign w36881 = ~w35618 & w35631;
assign w36882 = w36880 & ~w36881;
assign w36883 = ~w35621 & ~w36882;
assign w36884 = ~w35328 & w36880;
assign w36885 = w35297 & w36884;
assign w36886 = ~w36885 & w43086;
assign w36887 = (w36878 & w36885) | (w36878 & w43087) | (w36885 & w43087);
assign w36888 = ~w35993 & w46159;
assign w36889 = ~w36886 & ~w36887;
assign w36890 = ~w35994 & w36889;
assign w36891 = ~w36888 & ~w36890;
assign w36892 = (w4838 & w36890) | (w4838 & w46160) | (w36890 & w46160);
assign w36893 = (w36881 & ~w35297) | (w36881 & w43088) | (~w35297 & w43088);
assign w36894 = w36879 & ~w36893;
assign w36895 = ~w35603 & ~w35621;
assign w36896 = ~w5330 & w36895;
assign w36897 = ~w36894 & w36896;
assign w36898 = ~w35994 & w36897;
assign w36899 = ~w5745 & w36896;
assign w36900 = ~w35993 & w43089;
assign w36901 = ~w36898 & ~w36900;
assign w36902 = ~w5330 & ~w36895;
assign w36903 = w5745 & w36902;
assign w36904 = ~w35993 & w43090;
assign w36905 = w36894 & w36902;
assign w36906 = ~w35994 & w36905;
assign w36907 = ~w36904 & ~w36906;
assign w36908 = w36901 & w36907;
assign w36909 = ~w36892 & w36908;
assign w36910 = ~w35647 & ~w35652;
assign w36911 = w35623 & ~w36910;
assign w36912 = ~w35623 & w36910;
assign w36913 = ~w36911 & ~w36912;
assign w36914 = w36878 & w36895;
assign w36915 = w36894 & w36914;
assign w36916 = ~w36913 & ~w36915;
assign w36917 = w36913 & w36914;
assign w36918 = w36894 & w36917;
assign w36919 = ~w35994 & ~w36918;
assign w36920 = ~w36916 & w36919;
assign w36921 = ~w35993 & w43091;
assign w36922 = (~w36921 & ~w36919) | (~w36921 & w43092) | (~w36919 & w43092);
assign w36923 = ~w4430 & ~w36922;
assign w36924 = w36909 & ~w36923;
assign w36925 = w36877 & w36924;
assign w36926 = ~w4056 & ~w35665;
assign w36927 = ~w36027 & w36926;
assign w36928 = ~w35803 & w43093;
assign w36929 = ~w36927 & ~w36928;
assign w36930 = ~w4056 & ~w35661;
assign w36931 = w35666 & w36930;
assign w36932 = w35579 & ~w36931;
assign w36933 = (w35579 & w35994) | (w35579 & w43094) | (w35994 & w43094);
assign w36934 = ~w35994 & w43095;
assign w36935 = ~w36933 & ~w36934;
assign w36936 = w3646 & w36935;
assign w36937 = ~w35661 & ~w35664;
assign w36938 = w35649 & w36937;
assign w36939 = ~w36880 & w36938;
assign w36940 = w36881 & w36938;
assign w36941 = (w36940 & ~w35297) | (w36940 & w43096) | (~w35297 & w43096);
assign w36942 = ~w36939 & ~w36941;
assign w36943 = ~w35604 & ~w35652;
assign w36944 = ~w36937 & w36943;
assign w36945 = w36880 & w36944;
assign w36946 = ~w35647 & ~w36943;
assign w36947 = ~w35652 & ~w36937;
assign w36948 = ~w35649 & w36947;
assign w36949 = w36937 & w36946;
assign w36950 = ~w36948 & ~w36949;
assign w36951 = ~w36945 & w36950;
assign w36952 = w36881 & w36950;
assign w36953 = (w36952 & ~w35297) | (w36952 & w43097) | (~w35297 & w43097);
assign w36954 = ~w36951 & ~w36953;
assign w36955 = ~w35993 & w43098;
assign w36956 = w36942 & ~w36954;
assign w36957 = ~w35994 & w36956;
assign w36958 = ~w36955 & ~w36957;
assign w36959 = ~w36957 & w43099;
assign w36960 = ~w3646 & w35579;
assign w36961 = (w36960 & w35994) | (w36960 & w43100) | (w35994 & w43100);
assign w36962 = ~w3646 & ~w36932;
assign w36963 = ~w35994 & w43101;
assign w36964 = ~w36961 & ~w36963;
assign w36965 = w36959 & w36964;
assign w36966 = ~w36936 & ~w36965;
assign w36967 = w36925 & w36966;
assign w36968 = w36859 & w36967;
assign w36969 = (w35946 & w35993) | (w35946 & w43102) | (w35993 & w43102);
assign w36970 = ~w35859 & ~w36969;
assign w36971 = w35934 & w35974;
assign w36972 = ~w35760 & w36971;
assign w36973 = w35934 & ~w35972;
assign w36974 = ~w35945 & ~w35951;
assign w36975 = ~w36973 & w36974;
assign w36976 = (w36975 & ~w36972) | (w36975 & w46161) | (~w36972 & w46161);
assign w36977 = (w36972 & w46162) | (w36972 & w46163) | (w46162 & w46163);
assign w36978 = (~w35946 & w35993) | (~w35946 & w43104) | (w35993 & w43104);
assign w36979 = ~w36977 & w36978;
assign w36980 = w35858 & ~w36978;
assign w36981 = ~w36970 & w46164;
assign w36982 = (~w80 & w36978) | (~w80 & w46165) | (w36978 & w46165);
assign w36983 = ~w36979 & w36982;
assign w36984 = ~w36981 & ~w36983;
assign w36985 = ~w35993 & w46166;
assign w36986 = ~w35848 & ~w35849;
assign w36987 = w3 & w36986;
assign w36988 = ~w36985 & w36987;
assign w36989 = ~w36979 & w36988;
assign w36990 = w3 & ~w36986;
assign w36991 = (w35993 & w49810) | (w35993 & w49811) | (w49810 & w49811);
assign w36992 = ~w36977 & w36991;
assign w36993 = w36985 & w36990;
assign w36994 = ~w36992 & ~w36993;
assign w36995 = ~w36989 & w36994;
assign w36996 = w36984 & w36995;
assign w36997 = (w80 & w36970) | (w80 & w46167) | (w36970 & w46167);
assign w36998 = ~w36979 & ~w36980;
assign w36999 = w36997 & ~w36998;
assign w37000 = w35943 & w36748;
assign w37001 = (w37000 & ~w36739) | (w37000 & w46168) | (~w36739 & w46168);
assign w37002 = w35943 & ~w36763;
assign w37003 = ~w35897 & ~w37002;
assign w37004 = ~w252 & w35994;
assign w37005 = (w37003 & w35993) | (w37003 & w43105) | (w35993 & w43105);
assign w37006 = ~w37001 & w37005;
assign w37007 = ~w37004 & ~w37006;
assign w37008 = w35907 & ~w35951;
assign w37009 = ~w57 & ~w37008;
assign w37010 = (w37009 & w37006) | (w37009 & w43106) | (w37006 & w43106);
assign w37011 = ~w57 & w37008;
assign w37012 = ~w37006 & w43107;
assign w37013 = ~w37010 & ~w37012;
assign w37014 = ~w36999 & w37013;
assign w37015 = (~w36985 & w36977) | (~w36985 & w49264) | (w36977 & w49264);
assign w37016 = ~w3 & w36986;
assign w37017 = ~w37015 & w37016;
assign w37018 = ~w3 & ~w36986;
assign w37019 = w37015 & w37018;
assign w37020 = ~w37017 & ~w37019;
assign w37021 = ~w35860 & w50226;
assign w37022 = ~w35993 & w46170;
assign w37023 = ~w35841 & ~w35955;
assign w37024 = (w37023 & w35993) | (w37023 & w46171) | (w35993 & w46171);
assign w37025 = ~w37022 & ~w37024;
assign w37026 = ~w35993 & w46172;
assign w37027 = ~w37024 & ~w37026;
assign w37028 = w37021 & ~w37025;
assign w37029 = ~w37021 & w37027;
assign w37030 = ~w37028 & ~w37029;
assign w37031 = ~w42 & w37030;
assign w37032 = w37020 & ~w37031;
assign w37033 = w36996 & ~w37014;
assign w37034 = w37032 & ~w37033;
assign w37035 = (~w37008 & w37006) | (~w37008 & w49265) | (w37006 & w49265);
assign w37036 = w57 & ~w37035;
assign w37037 = w37007 & w37008;
assign w37038 = w37036 & ~w37037;
assign w37039 = w36996 & ~w37038;
assign w37040 = w37034 & ~w37039;
assign w37041 = w35861 & w50226;
assign w37042 = ~w35955 & ~w37041;
assign w37043 = w35834 & w35840;
assign w37044 = w42 & ~w37043;
assign w37045 = ~w35823 & ~w37044;
assign w37046 = ~w37042 & ~w37045;
assign w37047 = ~w35824 & ~w37046;
assign w37048 = w35836 & w35956;
assign w37049 = w37042 & w37048;
assign w37050 = w37047 & ~w37049;
assign w37051 = w42 & w35841;
assign w37052 = ~w37021 & w37051;
assign w37053 = w37050 & ~w37052;
assign w37054 = w35824 & w35955;
assign w37055 = w37021 & w37054;
assign w37056 = ~w37053 & ~w37055;
assign w37057 = ~w37040 & ~w37056;
assign w37058 = w36968 & w37057;
assign w37059 = ~w36817 & w37058;
assign w37060 = ~w36576 & w37059;
assign w37061 = ~w36700 & w36711;
assign w37062 = w2285 & w36696;
assign w37063 = ~w36682 & ~w36698;
assign w37064 = w37062 & w37063;
assign w37065 = w36691 & ~w37064;
assign w37066 = w37061 & ~w37065;
assign w37067 = w36736 & w36813;
assign w37068 = w36659 & w36813;
assign w37069 = ~w37066 & w37068;
assign w37070 = ~w37067 & ~w37069;
assign w37071 = w36807 & w37034;
assign w37072 = ~w36874 & w46173;
assign w37073 = w5330 & w36895;
assign w37074 = w5745 & w37073;
assign w37075 = ~w35993 & w43109;
assign w37076 = w36894 & w37073;
assign w37077 = ~w35994 & w37076;
assign w37078 = ~w37075 & ~w37077;
assign w37079 = w5330 & ~w36895;
assign w37080 = ~w36894 & w37079;
assign w37081 = ~w35994 & w37080;
assign w37082 = ~w5745 & w37079;
assign w37083 = ~w35993 & w43110;
assign w37084 = ~w37081 & ~w37083;
assign w37085 = w37078 & w37084;
assign w37086 = ~w37072 & w37085;
assign w37087 = w36909 & ~w37086;
assign w37088 = (w4056 & w36957) | (w4056 & w43111) | (w36957 & w43111);
assign w37089 = w36964 & ~w37088;
assign w37090 = ~w36890 & w46174;
assign w37091 = w4430 & ~w36921;
assign w37092 = ~w36920 & w37091;
assign w37093 = ~w37090 & ~w37092;
assign w37094 = w36923 & w37089;
assign w37095 = w36966 & ~w37094;
assign w37096 = w37089 & w37093;
assign w37097 = ~w37087 & w37096;
assign w37098 = w37095 & ~w37097;
assign w37099 = ~w3242 & w36855;
assign w37100 = ~w37098 & w43112;
assign w37101 = w36859 & ~w37100;
assign w37102 = ~w36815 & w37071;
assign w37103 = (w37057 & w36799) | (w37057 & w43113) | (w36799 & w43113);
assign w37104 = w37071 & ~w37101;
assign w37105 = ~w37070 & w37104;
assign w37106 = w37103 & ~w37105;
assign w37107 = ~w37060 & ~w37106;
assign w37108 = w612 & ~w37107;
assign w37109 = ~w36968 & ~w37101;
assign w37110 = ~w36575 & ~w37101;
assign w37111 = (w37110 & ~w36570) | (w37110 & w46175) | (~w36570 & w46175);
assign w37112 = (~w37109 & w36572) | (~w37109 & w43114) | (w36572 & w43114);
assign w37113 = w36658 & ~w37066;
assign w37114 = w36603 & w37113;
assign w37115 = (~w36572 & w46176) | (~w36572 & w46177) | (w46176 & w46177);
assign w37116 = ~w36715 & ~w36736;
assign w37117 = ~w37060 & w46178;
assign w37118 = ~w37115 & w37117;
assign w37119 = ~w37108 & ~w37118;
assign w37120 = w36011 & ~w37119;
assign w37121 = ~w36011 & w37119;
assign w37122 = ~w37120 & ~w37121;
assign w37123 = w493 & w37122;
assign w37124 = w36005 & w37116;
assign w37125 = ~w37115 & w37124;
assign w37126 = w36010 & ~w37125;
assign w37127 = w36795 & w36812;
assign w37128 = w36789 & ~w36790;
assign w37129 = ~w36789 & w36790;
assign w37130 = ~w37128 & ~w37129;
assign w37131 = ~w37107 & w37130;
assign w37132 = w37107 & w37127;
assign w37133 = ~w37126 & w37132;
assign w37134 = w37107 & ~w37127;
assign w37135 = w37126 & w37134;
assign w37136 = ~w37133 & ~w37135;
assign w37137 = ~w37131 & w37136;
assign w37138 = ~w400 & w37137;
assign w37139 = ~w37123 & ~w37138;
assign w37140 = ~w36734 & w37061;
assign w37141 = (w37140 & w37101) | (w37140 & w46179) | (w37101 & w46179);
assign w37142 = ~w36734 & ~w37113;
assign w37143 = ~w36587 & ~w36716;
assign w37144 = (w46181 & w49266) | (w46181 & w49267) | (w49266 & w49267);
assign w37145 = w37143 & w52288;
assign w37146 = ~w37144 & ~w37145;
assign w37147 = ~w36586 & ~w37107;
assign w37148 = w37107 & ~w37146;
assign w37149 = ~w37147 & ~w37148;
assign w37150 = w754 & w37149;
assign w37151 = ~w754 & ~w37107;
assign w37152 = ~w36716 & w37141;
assign w37153 = ~w37111 & w37152;
assign w37154 = w36735 & ~w37113;
assign w37155 = ~w36587 & ~w37154;
assign w37156 = ~w37060 & w46182;
assign w37157 = ~w37153 & w37156;
assign w37158 = ~w37151 & ~w37157;
assign w37159 = w36602 & w36665;
assign w37160 = w612 & w37159;
assign w37161 = ~w37158 & w37160;
assign w37162 = w612 & ~w37159;
assign w37163 = w37158 & w37162;
assign w37164 = ~w37161 & ~w37163;
assign w37165 = ~w37150 & w37164;
assign w37166 = w36616 & w36710;
assign w37167 = ~w36700 & w36705;
assign w37168 = (w37167 & w37101) | (w37167 & w46183) | (w37101 & w46183);
assign w37169 = w37166 & w37168;
assign w37170 = w36705 & ~w37065;
assign w37171 = w37166 & w37170;
assign w37172 = w36616 & ~w37171;
assign w37173 = (w37172 & w37111) | (w37172 & w43116) | (w37111 & w43116);
assign w37174 = w36656 & w37173;
assign w37175 = w36725 & ~w37174;
assign w37176 = (w46181 & w49268) | (w46181 & w49269) | (w49268 & w49269);
assign w37177 = ~w36619 & ~w36620;
assign w37178 = w36621 & ~w37177;
assign w37179 = ~w36621 & w37177;
assign w37180 = ~w37178 & ~w37179;
assign w37181 = (~w37180 & w37060) | (~w37180 & w46184) | (w37060 & w46184);
assign w37182 = w36630 & w36733;
assign w37183 = ~w37113 & w37182;
assign w37184 = ~w37060 & w46185;
assign w37185 = w37061 & w37182;
assign w37186 = w37112 & w37185;
assign w37187 = w37184 & ~w37186;
assign w37188 = ~w37181 & ~w37187;
assign w37189 = ~w37176 & ~w37181;
assign w37190 = ~w37175 & w37189;
assign w37191 = ~w37188 & ~w37190;
assign w37192 = ~w945 & w37191;
assign w37193 = w37165 & ~w37192;
assign w37194 = w37139 & w37193;
assign w37195 = ~w37170 & w50227;
assign w37196 = (~w37171 & w37111) | (~w37171 & w43118) | (w37111 & w43118);
assign w37197 = w37107 & w37196;
assign w37198 = (w46187 & w49270) | (w46187 & w49271) | (w49270 & w49271);
assign w37199 = w37197 & ~w37198;
assign w37200 = w36610 & ~w36611;
assign w37201 = ~w36610 & w36611;
assign w37202 = ~w37200 & ~w37201;
assign w37203 = (~w37202 & w37060) | (~w37202 & w46188) | (w37060 & w46188);
assign w37204 = ~w1320 & ~w37203;
assign w37205 = ~w37199 & w37204;
assign w37206 = w36656 & w36725;
assign w37207 = w37172 & w37206;
assign w37208 = (w37207 & w37111) | (w37207 & w43119) | (w37111 & w43119);
assign w37209 = ~w36645 & ~w36646;
assign w37210 = w36647 & ~w37209;
assign w37211 = ~w36647 & w37209;
assign w37212 = ~w37210 & ~w37211;
assign w37213 = w37107 & ~w37208;
assign w37214 = (~w37212 & w37060) | (~w37212 & w46189) | (w37060 & w46189);
assign w37215 = ~w37213 & ~w37214;
assign w37216 = ~w37106 & ~w37206;
assign w37217 = ~w37060 & w37216;
assign w37218 = ~w37173 & w37217;
assign w37219 = (w1120 & ~w37217) | (w1120 & w46190) | (~w37217 & w46190);
assign w37220 = ~w37215 & w37219;
assign w37221 = ~w37205 & ~w37220;
assign w37222 = ~w37215 & ~w37218;
assign w37223 = (~w1120 & w37215) | (~w1120 & w46191) | (w37215 & w46191);
assign w37224 = ~w37221 & ~w37223;
assign w37225 = (~w36697 & w37101) | (~w36697 & w46192) | (w37101 & w46192);
assign w37226 = (~w37064 & w37111) | (~w37064 & w43120) | (w37111 & w43120);
assign w37227 = w37107 & w37226;
assign w37228 = w37107 & w46193;
assign w37229 = (~w1738 & w37060) | (~w1738 & w46194) | (w37060 & w46194);
assign w37230 = w36690 & w36705;
assign w37231 = w1541 & ~w37230;
assign w37232 = ~w37229 & w37231;
assign w37233 = ~w37228 & w37232;
assign w37234 = w1541 & w37230;
assign w37235 = ~w36682 & w37234;
assign w37236 = w37107 & w46195;
assign w37237 = w37229 & w37234;
assign w37238 = ~w37236 & ~w37237;
assign w37239 = ~w37233 & w37238;
assign w37240 = (w1541 & w37060) | (w1541 & w46196) | (w37060 & w46196);
assign w37241 = w37107 & ~w37195;
assign w37242 = w1320 & ~w37166;
assign w37243 = (w37242 & w37241) | (w37242 & w46197) | (w37241 & w46197);
assign w37244 = w1320 & w37166;
assign w37245 = ~w37241 & w46198;
assign w37246 = ~w37243 & ~w37245;
assign w37247 = w37239 & w37246;
assign w37248 = ~w37223 & w37247;
assign w37249 = (w36681 & w37060) | (w36681 & w46199) | (w37060 & w46199);
assign w37250 = ~w37062 & ~w37063;
assign w37251 = w1738 & w37249;
assign w37252 = w1738 & w52289;
assign w37253 = w37227 & w37252;
assign w37254 = ~w37251 & ~w37253;
assign w37255 = ~w36697 & ~w37062;
assign w37256 = (w37255 & w37101) | (w37255 & w46202) | (w37101 & w46202);
assign w37257 = (w37256 & w36572) | (w37256 & w43122) | (w36572 & w43122);
assign w37258 = w37106 & w37255;
assign w37259 = ~w37257 & ~w37258;
assign w37260 = ~w2285 & w37106;
assign w37261 = ~w36817 & w43123;
assign w37262 = ~w36576 & w37261;
assign w37263 = ~w37260 & ~w37262;
assign w37264 = ~w36817 & w43124;
assign w37265 = ~w36576 & w37264;
assign w37266 = w36697 & w37106;
assign w37267 = ~w37265 & ~w37266;
assign w37268 = ~w37106 & ~w37255;
assign w37269 = ~w37112 & w37268;
assign w37270 = w37267 & ~w37269;
assign w37271 = ~w37259 & w37263;
assign w37272 = w37270 & ~w37271;
assign w37273 = w37250 & w37259;
assign w37274 = w37227 & ~w37273;
assign w37275 = ~w1738 & ~w37249;
assign w37276 = ~w37274 & w37275;
assign w37277 = ~w2006 & ~w37272;
assign w37278 = w37254 & w37277;
assign w37279 = ~w37276 & ~w37278;
assign w37280 = ~w37228 & ~w37229;
assign w37281 = ~w1541 & ~w37230;
assign w37282 = ~w37280 & w37281;
assign w37283 = ~w1541 & w37230;
assign w37284 = w37280 & w37283;
assign w37285 = ~w37282 & ~w37284;
assign w37286 = w37279 & w37285;
assign w37287 = (~w37224 & w37286) | (~w37224 & w38190) | (w37286 & w38190);
assign w37288 = w945 & ~w37191;
assign w37289 = ~w754 & ~w37149;
assign w37290 = ~w37288 & ~w37289;
assign w37291 = w37165 & ~w37290;
assign w37292 = w37158 & ~w37159;
assign w37293 = ~w37158 & w37159;
assign w37294 = ~w37292 & ~w37293;
assign w37295 = ~w493 & ~w37122;
assign w37296 = ~w612 & w37294;
assign w37297 = ~w37295 & ~w37296;
assign w37298 = ~w37291 & w37297;
assign w37299 = w37139 & ~w37298;
assign w37300 = w400 & ~w37137;
assign w37301 = w36795 & w37124;
assign w37302 = ~w37115 & w37301;
assign w37303 = ~w36814 & ~w37302;
assign w37304 = ~w36747 & ~w36804;
assign w37305 = ~w36746 & ~w37107;
assign w37306 = w37107 & ~w37304;
assign w37307 = w37303 & w37306;
assign w37308 = ~w37305 & ~w37307;
assign w37309 = w37107 & w37304;
assign w37310 = ~w37303 & w37309;
assign w37311 = w37308 & ~w37310;
assign w37312 = ~w351 & ~w37311;
assign w37313 = ~w37300 & ~w37312;
assign w37314 = ~w37299 & w37313;
assign w37315 = w37194 & ~w37287;
assign w37316 = w37314 & ~w37315;
assign w37317 = ~w36099 & ~w36115;
assign w37318 = ~w36086 & ~w36111;
assign w37319 = ~w36107 & ~w36116;
assign w37320 = w37318 & w37319;
assign w37321 = ~w36116 & ~w37320;
assign w37322 = w37317 & ~w37321;
assign w37323 = ~w37317 & w37321;
assign w37324 = ~w37322 & ~w37323;
assign w37325 = ~w26880 & w37324;
assign w37326 = ~w37106 & ~w37325;
assign w37327 = ~w26880 & w36098;
assign w37328 = w37106 & ~w37327;
assign w37329 = ~w36817 & w43125;
assign w37330 = ~w36576 & w37329;
assign w37331 = ~w37328 & ~w37330;
assign w37332 = ~w37060 & w37326;
assign w37333 = w37331 & ~w37332;
assign w37334 = ~w26880 & ~w36119;
assign w37335 = w26880 & w36119;
assign w37336 = ~w37334 & ~w37335;
assign w37337 = ~w37106 & w37336;
assign w37338 = ~w37060 & w37337;
assign w37339 = w36135 & ~w37338;
assign w37340 = ~w36135 & w37338;
assign w37341 = ~w37339 & ~w37340;
assign w37342 = ~w25851 & ~w37333;
assign w37343 = w37341 & ~w37342;
assign w37344 = w25851 & w37333;
assign w37345 = ~w37343 & ~w37344;
assign w37346 = ~w36127 & w36140;
assign w37347 = ~w36135 & ~w37335;
assign w37348 = ~w37334 & ~w37347;
assign w37349 = w37346 & ~w37348;
assign w37350 = ~w37346 & w37348;
assign w37351 = ~w37349 & ~w37350;
assign w37352 = (~w36126 & w37060) | (~w36126 & w46203) | (w37060 & w46203);
assign w37353 = ~w37060 & w46204;
assign w37354 = ~w37352 & ~w37353;
assign w37355 = w24874 & ~w37354;
assign w37356 = ~w36035 & ~w36068;
assign w37357 = ~w36069 & ~w37356;
assign w37358 = w36043 & ~w37357;
assign w37359 = w36074 & ~w37358;
assign w37360 = ~w30239 & w37359;
assign w37361 = w30239 & ~w37359;
assign w37362 = ~w37360 & ~w37361;
assign w37363 = ~w37106 & ~w37362;
assign w37364 = ~w37060 & w37363;
assign w37365 = ~w29158 & w36110;
assign w37366 = ~w37364 & w37365;
assign w37367 = ~w29158 & ~w36110;
assign w37368 = w37364 & w37367;
assign w37369 = ~w37366 & ~w37368;
assign w37370 = w37318 & ~w37319;
assign w37371 = ~w37318 & w37319;
assign w37372 = ~w37370 & ~w37371;
assign w37373 = w28077 & ~w36106;
assign w37374 = (w37373 & w37060) | (w37373 & w46205) | (w37060 & w46205);
assign w37375 = w28077 & ~w37372;
assign w37376 = ~w37060 & w46206;
assign w37377 = ~w37374 & ~w37376;
assign w37378 = w37369 & w37377;
assign w37379 = ~w37355 & w37378;
assign w37380 = w37345 & w37379;
assign w37381 = ~a[2] & ~a[3];
assign w37382 = ~a[4] & w37381;
assign w37383 = w35994 & ~w37382;
assign w37384 = ~w35994 & w37382;
assign w37385 = a[5] & ~w37384;
assign w37386 = ~w37383 & ~w37385;
assign w37387 = a[5] & w37383;
assign w37388 = ~w36044 & ~w37387;
assign w37389 = w34900 & ~w37384;
assign w37390 = ~w37388 & w37389;
assign w37391 = w34900 & ~w37386;
assign w37392 = (w37391 & w37060) | (w37391 & w46207) | (w37060 & w46207);
assign w37393 = ~w37060 & w46208;
assign w37394 = ~w37392 & ~w37393;
assign w37395 = ~a[6] & ~w35994;
assign w37396 = a[6] & w35994;
assign w37397 = ~w37395 & ~w37396;
assign w37398 = a[6] & ~w36044;
assign w37399 = (w37397 & w37060) | (w37397 & w46209) | (w37060 & w46209);
assign w37400 = ~w36045 & ~w37398;
assign w37401 = ~w37060 & w46210;
assign w37402 = ~w37399 & ~w37401;
assign w37403 = w37394 & ~w37402;
assign w37404 = ~w34900 & w37384;
assign w37405 = ~w37106 & ~w37404;
assign w37406 = ~w34900 & w37386;
assign w37407 = ~w37060 & w37405;
assign w37408 = w37406 & ~w37407;
assign w37409 = ~w34900 & w37388;
assign w37410 = ~w37060 & w46211;
assign w37411 = ~w37408 & ~w37410;
assign w37412 = w35023 & ~w35994;
assign w37413 = a[7] & ~w37395;
assign w37414 = ~w37412 & ~w37413;
assign w37415 = ~a[7] & ~w35994;
assign w37416 = a[7] & w35994;
assign w37417 = ~w37415 & ~w37416;
assign w37418 = w34900 & ~w37417;
assign w37419 = ~w34900 & w37417;
assign w37420 = ~w37418 & ~w37419;
assign w37421 = ~w36045 & w37420;
assign w37422 = w36045 & ~w37420;
assign w37423 = ~w37421 & ~w37422;
assign w37424 = ~w33731 & w37414;
assign w37425 = (w37424 & w37060) | (w37424 & w46212) | (w37060 & w46212);
assign w37426 = ~w33731 & ~w37423;
assign w37427 = ~w37060 & w46213;
assign w37428 = ~w37425 & ~w37427;
assign w37429 = w37411 & w37428;
assign w37430 = ~w37403 & w37429;
assign w37431 = ~w34900 & w35994;
assign w37432 = ~w37412 & ~w37431;
assign w37433 = a[8] & ~w37432;
assign w37434 = ~a[8] & w37432;
assign w37435 = ~w37433 & ~w37434;
assign w37436 = a[6] & w37415;
assign w37437 = ~w37418 & ~w37421;
assign w37438 = ~w37436 & ~w37437;
assign w37439 = ~w33731 & w37438;
assign w37440 = w33731 & ~w37438;
assign w37441 = ~w37439 & ~w37440;
assign w37442 = ~w37106 & ~w37441;
assign w37443 = ~w37060 & w37442;
assign w37444 = w37435 & ~w37443;
assign w37445 = ~w37435 & w37443;
assign w37446 = ~w37444 & ~w37445;
assign w37447 = ~w32698 & ~w37446;
assign w37448 = ~w36068 & ~w36069;
assign w37449 = ~w37106 & w37448;
assign w37450 = ~w37060 & w37449;
assign w37451 = w31477 & w36035;
assign w37452 = ~w37450 & w37451;
assign w37453 = w31477 & ~w36035;
assign w37454 = w37450 & w37453;
assign w37455 = ~w37452 & ~w37454;
assign w37456 = w33731 & ~w37414;
assign w37457 = (w37456 & w37060) | (w37456 & w46214) | (w37060 & w46214);
assign w37458 = w33731 & w37423;
assign w37459 = ~w37060 & w46215;
assign w37460 = ~w37457 & ~w37459;
assign w37461 = w37455 & w37460;
assign w37462 = ~w37447 & w37461;
assign w37463 = ~w37430 & w37462;
assign w37464 = ~w31477 & w36074;
assign w37465 = w36043 & ~w37464;
assign w37466 = w36043 & w36074;
assign w37467 = w37357 & ~w37466;
assign w37468 = ~w37357 & w37466;
assign w37469 = ~w37467 & ~w37468;
assign w37470 = ~w37107 & w37465;
assign w37471 = w37107 & w37469;
assign w37472 = ~w37470 & ~w37471;
assign w37473 = ~w30239 & ~w37472;
assign w37474 = w32698 & ~w37435;
assign w37475 = ~w37443 & w37474;
assign w37476 = w32698 & w37435;
assign w37477 = w37443 & w37476;
assign w37478 = ~w37475 & ~w37477;
assign w37479 = ~w31477 & ~w36035;
assign w37480 = ~w37450 & w37479;
assign w37481 = ~w31477 & w36035;
assign w37482 = w37450 & w37481;
assign w37483 = ~w37480 & ~w37482;
assign w37484 = w37478 & w37483;
assign w37485 = w37455 & ~w37484;
assign w37486 = ~w37473 & ~w37485;
assign w37487 = ~w37463 & w37486;
assign w37488 = w37380 & w37487;
assign w37489 = w30239 & w37472;
assign w37490 = ~w36110 & ~w37364;
assign w37491 = w36110 & w37364;
assign w37492 = ~w37490 & ~w37491;
assign w37493 = w29158 & ~w37492;
assign w37494 = ~w37489 & ~w37493;
assign w37495 = w37380 & ~w37494;
assign w37496 = w26880 & ~w37324;
assign w37497 = ~w37106 & ~w37496;
assign w37498 = w26880 & ~w36098;
assign w37499 = w37106 & ~w37498;
assign w37500 = ~w36817 & w43126;
assign w37501 = ~w36576 & w37500;
assign w37502 = ~w37499 & ~w37501;
assign w37503 = ~w37060 & w37497;
assign w37504 = w37502 & ~w37503;
assign w37505 = ~w28077 & w37372;
assign w37506 = ~w37106 & ~w37505;
assign w37507 = ~w28077 & w36106;
assign w37508 = w37106 & ~w37507;
assign w37509 = ~w36817 & w43127;
assign w37510 = ~w36576 & w37509;
assign w37511 = ~w37508 & ~w37510;
assign w37512 = ~w37060 & w37506;
assign w37513 = w37511 & ~w37512;
assign w37514 = ~w37504 & ~w37513;
assign w37515 = ~w25851 & w36135;
assign w37516 = ~w37338 & w37515;
assign w37517 = ~w25851 & ~w36135;
assign w37518 = w37338 & w37517;
assign w37519 = ~w37516 & ~w37518;
assign w37520 = w37514 & w37519;
assign w37521 = ~w37355 & ~w37520;
assign w37522 = w37345 & w37521;
assign w37523 = ~w24874 & w37354;
assign w37524 = ~w36114 & w46216;
assign w37525 = (w24874 & w37060) | (w24874 & w46217) | (w37060 & w46217);
assign w37526 = w36142 & ~w37524;
assign w37527 = ~w37060 & w46218;
assign w37528 = ~w37525 & ~w37527;
assign w37529 = w36161 & ~w36214;
assign w37530 = ~w23843 & ~w37529;
assign w37531 = w37528 & w37530;
assign w37532 = ~w23843 & w37529;
assign w37533 = ~w37528 & w37532;
assign w37534 = ~w37531 & ~w37533;
assign w37535 = ~w37523 & w37534;
assign w37536 = ~w37522 & w37535;
assign w37537 = ~w37495 & w37536;
assign w37538 = ~w37488 & w37537;
assign w37539 = ~w36119 & w36163;
assign w37540 = ~w36150 & ~w36224;
assign w37541 = (w36203 & w37539) | (w36203 & w46219) | (w37539 & w46219);
assign w37542 = ~w36173 & ~w36205;
assign w37543 = ~w36185 & ~w36206;
assign w37544 = w37542 & ~w37543;
assign w37545 = ~w37542 & w37543;
assign w37546 = ~w37544 & ~w37545;
assign w37547 = w37541 & ~w37546;
assign w37548 = ~w37541 & w37546;
assign w37549 = ~w37547 & ~w37548;
assign w37550 = ~w20000 & ~w36172;
assign w37551 = (w37550 & w37060) | (w37550 & w46220) | (w37060 & w46220);
assign w37552 = ~w20000 & w37549;
assign w37553 = ~w37060 & w46221;
assign w37554 = ~w37551 & ~w37553;
assign w37555 = w36196 & ~w37540;
assign w37556 = ~w37539 & w37555;
assign w37557 = w36201 & ~w37556;
assign w37558 = w36186 & ~w37557;
assign w37559 = ~w36186 & w37557;
assign w37560 = ~w37558 & ~w37559;
assign w37561 = w20906 & w36183;
assign w37562 = (w37561 & w37060) | (w37561 & w46222) | (w37060 & w46222);
assign w37563 = w20906 & ~w37560;
assign w37564 = w37107 & w37563;
assign w37565 = ~w37562 & ~w37564;
assign w37566 = w37554 & w37565;
assign w37567 = w20000 & w36172;
assign w37568 = (w37567 & w37060) | (w37567 & w46223) | (w37060 & w46223);
assign w37569 = w20000 & ~w37549;
assign w37570 = ~w37060 & w46224;
assign w37571 = ~w37568 & ~w37570;
assign w37572 = ~w37539 & w46225;
assign w37573 = w36142 & w36161;
assign w37574 = ~w36150 & w36202;
assign w37575 = ~w36215 & w37574;
assign w37576 = w37573 & w37574;
assign w37577 = ~w37524 & w37576;
assign w37578 = ~w37575 & ~w37577;
assign w37579 = ~w37572 & w37578;
assign w37580 = ~w21801 & w37579;
assign w37581 = ~w34987 & ~w36191;
assign w37582 = w34987 & w36191;
assign w37583 = ~w37581 & ~w37582;
assign w37584 = ~w21801 & ~w37583;
assign w37585 = w37106 & ~w37584;
assign w37586 = ~w36817 & w43128;
assign w37587 = ~w36576 & w37586;
assign w37588 = ~w37585 & ~w37587;
assign w37589 = ~w37106 & ~w37580;
assign w37590 = ~w37060 & w37589;
assign w37591 = w37588 & ~w37590;
assign w37592 = ~w37524 & w37573;
assign w37593 = ~w36214 & ~w37592;
assign w37594 = ~w36149 & ~w36150;
assign w37595 = ~w22767 & ~w37594;
assign w37596 = w37593 & w37595;
assign w37597 = ~w22767 & w37594;
assign w37598 = ~w37593 & w37597;
assign w37599 = ~w37596 & ~w37598;
assign w37600 = ~w22767 & w36148;
assign w37601 = ~w36817 & w43129;
assign w37602 = ~w36576 & w37601;
assign w37603 = w37106 & w37600;
assign w37604 = ~w37602 & ~w37603;
assign w37605 = ~w37106 & ~w37599;
assign w37606 = ~w37060 & w37605;
assign w37607 = w37604 & ~w37606;
assign w37608 = ~w37591 & ~w37607;
assign w37609 = w36215 & ~w37592;
assign w37610 = w21801 & w37572;
assign w37611 = w21801 & w37574;
assign w37612 = ~w37609 & w37611;
assign w37613 = ~w37610 & ~w37612;
assign w37614 = w21801 & w37583;
assign w37615 = w37106 & ~w37614;
assign w37616 = ~w36817 & w49272;
assign w37617 = ~w36576 & w37616;
assign w37618 = ~w37615 & ~w37617;
assign w37619 = ~w37106 & w37613;
assign w37620 = ~w37060 & w37619;
assign w37621 = w37618 & ~w37620;
assign w37622 = ~w20906 & ~w36186;
assign w37623 = ~w37557 & w37622;
assign w37624 = ~w20906 & w36186;
assign w37625 = w37557 & w37624;
assign w37626 = ~w37623 & ~w37625;
assign w37627 = ~w37106 & w37626;
assign w37628 = ~w20906 & ~w36183;
assign w37629 = w37106 & ~w37628;
assign w37630 = ~w36817 & w49273;
assign w37631 = ~w36576 & w37630;
assign w37632 = ~w37629 & ~w37631;
assign w37633 = ~w37060 & w37627;
assign w37634 = w37632 & ~w37633;
assign w37635 = ~w37621 & ~w37634;
assign w37636 = (w37571 & ~w37565) | (w37571 & w46226) | (~w37565 & w46226);
assign w37637 = w37571 & ~w37608;
assign w37638 = w37635 & w37637;
assign w37639 = ~w37636 & ~w37638;
assign w37640 = ~w36242 & ~w36564;
assign w37641 = w36332 & ~w36385;
assign w37642 = w37640 & ~w37641;
assign w37643 = ~w37640 & w37641;
assign w37644 = ~w37642 & ~w37643;
assign w37645 = (w36384 & w37060) | (w36384 & w46227) | (w37060 & w46227);
assign w37646 = ~w37060 & w46228;
assign w37647 = ~w37645 & ~w37646;
assign w37648 = w18183 & w37647;
assign w37649 = ~w18183 & ~w37647;
assign w37650 = ~w36238 & ~w36564;
assign w37651 = ~w36173 & w37541;
assign w37652 = w36209 & ~w37651;
assign w37653 = w37650 & ~w37652;
assign w37654 = ~w37650 & w37652;
assign w37655 = ~w37653 & ~w37654;
assign w37656 = (w36237 & w37060) | (w36237 & w46229) | (w37060 & w46229);
assign w37657 = w37107 & ~w37655;
assign w37658 = ~w37656 & ~w37657;
assign w37659 = (w19040 & w37657) | (w19040 & w46230) | (w37657 & w46230);
assign w37660 = ~w37649 & w37659;
assign w37661 = ~w37648 & ~w37660;
assign w37662 = ~w37639 & w37661;
assign w37663 = w37538 & w37662;
assign w37664 = w37528 & ~w37529;
assign w37665 = ~w37528 & w37529;
assign w37666 = ~w37664 & ~w37665;
assign w37667 = w23843 & w37666;
assign w37668 = w37593 & ~w37594;
assign w37669 = ~w37593 & w37594;
assign w37670 = ~w37668 & ~w37669;
assign w37671 = (w36148 & w37060) | (w36148 & w46231) | (w37060 & w46231);
assign w37672 = ~w37060 & w46232;
assign w37673 = ~w37671 & ~w37672;
assign w37674 = w22767 & w37673;
assign w37675 = w37591 & ~w37634;
assign w37676 = w37566 & w46233;
assign w37677 = ~w37667 & w37676;
assign w37678 = w37662 & ~w37677;
assign w37679 = ~w35215 & w35994;
assign w37680 = ~w35994 & w36309;
assign w37681 = ~w37679 & ~w37680;
assign w37682 = w36314 & w36321;
assign w37683 = (~w36385 & w36242) | (~w36385 & w46234) | (w36242 & w46234);
assign w37684 = w36332 & ~w37683;
assign w37685 = w37682 & ~w37684;
assign w37686 = ~w37682 & w37684;
assign w37687 = ~w37685 & ~w37686;
assign w37688 = ~w37107 & ~w37681;
assign w37689 = w37107 & w37687;
assign w37690 = ~w37688 & ~w37689;
assign w37691 = w17380 & w37690;
assign w37692 = ~w19040 & w37658;
assign w37693 = ~w37648 & w37692;
assign w37694 = ~w37649 & ~w37693;
assign w37695 = ~w37691 & w37694;
assign w37696 = ~w37678 & w37695;
assign w37697 = w36514 & ~w36525;
assign w37698 = ~w36533 & ~w36549;
assign w37699 = ~w36369 & w46235;
assign w37700 = w36242 & w37699;
assign w37701 = ~w36567 & w37698;
assign w37702 = (~w36549 & w36567) | (~w36549 & w43130) | (w36567 & w43130);
assign w37703 = ~w37700 & w37702;
assign w37704 = w37697 & ~w37703;
assign w37705 = ~w37697 & w37703;
assign w37706 = (~w36524 & w37060) | (~w36524 & w46236) | (w37060 & w46236);
assign w37707 = ~w37704 & ~w37705;
assign w37708 = w37107 & w37707;
assign w37709 = (w11138 & w37708) | (w11138 & w46237) | (w37708 & w46237);
assign w37710 = w36289 & w36296;
assign w37711 = w36559 & ~w37710;
assign w37712 = ~w36337 & w37711;
assign w37713 = w36333 & w37711;
assign w37714 = w36385 & w37713;
assign w37715 = ~w36564 & w37713;
assign w37716 = (~w37714 & w36242) | (~w37714 & w46238) | (w36242 & w46238);
assign w37717 = ~w37712 & w37716;
assign w37718 = w36560 & ~w37698;
assign w37719 = ~w37717 & w37718;
assign w37720 = w36558 & ~w37698;
assign w37721 = ~w37701 & ~w37720;
assign w37722 = ~w37700 & w37721;
assign w37723 = ~w37719 & w37722;
assign w37724 = (~w36532 & w37060) | (~w36532 & w46239) | (w37060 & w46239);
assign w37725 = w37107 & w37723;
assign w37726 = ~w37724 & ~w37725;
assign w37727 = ~w11138 & w36514;
assign w37728 = (~w11870 & w37703) | (~w11870 & w37731) | (w37703 & w37731);
assign w37729 = ~w11138 & w37705;
assign w37730 = w37728 & ~w37729;
assign w37731 = ~w11870 & ~w37727;
assign w37732 = (w37731 & w37060) | (w37731 & w46240) | (w37060 & w46240);
assign w37733 = w37107 & w37730;
assign w37734 = ~w37732 & ~w37733;
assign w37735 = ~w37726 & ~w37734;
assign w37736 = ~w37709 & ~w37735;
assign w37737 = ~w36380 & ~w37712;
assign w37738 = w37716 & w37737;
assign w37739 = w36365 & ~w37738;
assign w37740 = ~w36376 & ~w36557;
assign w37741 = w37739 & w37740;
assign w37742 = ~w37739 & ~w37740;
assign w37743 = w37107 & w46241;
assign w37744 = w36375 & ~w37107;
assign w37745 = (~w12666 & w37107) | (~w12666 & w46242) | (w37107 & w46242);
assign w37746 = ~w37743 & w37745;
assign w37747 = w36365 & ~w36380;
assign w37748 = w37717 & ~w37747;
assign w37749 = ~w37717 & w37747;
assign w37750 = ~w37748 & ~w37749;
assign w37751 = (~w36379 & w37060) | (~w36379 & w46243) | (w37060 & w46243);
assign w37752 = w37107 & w37750;
assign w37753 = ~w37751 & ~w37752;
assign w37754 = ~w37752 & w46244;
assign w37755 = ~w37746 & ~w37754;
assign w37756 = w37736 & w37755;
assign w37757 = ~w36316 & ~w36385;
assign w37758 = (w37757 & w36242) | (w37757 & w46245) | (w36242 & w46245);
assign w37759 = ~w36335 & ~w37758;
assign w37760 = ~w36259 & ~w37759;
assign w37761 = w36348 & ~w37760;
assign w37762 = w36287 & ~w37761;
assign w37763 = w36277 & ~w36353;
assign w37764 = ~w37060 & w46246;
assign w37765 = (w36352 & w37060) | (w36352 & w46247) | (w37060 & w46247);
assign w37766 = ~w37764 & ~w37765;
assign w37767 = w37107 & ~w37762;
assign w37768 = w37766 & ~w37767;
assign w37769 = ~w37762 & w37764;
assign w37770 = w14039 & ~w37769;
assign w37771 = ~w37768 & w37770;
assign w37772 = ~w13384 & ~w37753;
assign w37773 = ~w37771 & ~w37772;
assign w37774 = ~w37743 & ~w37744;
assign w37775 = w12666 & ~w37774;
assign w37776 = ~w37725 & w46248;
assign w37777 = ~w37708 & w46249;
assign w37778 = ~w37776 & ~w37777;
assign w37779 = ~w37775 & w37778;
assign w37780 = w37756 & ~w37773;
assign w37781 = w37736 & ~w37779;
assign w37782 = ~w37780 & ~w37781;
assign w37783 = ~w36259 & w36347;
assign w37784 = w37759 & w37783;
assign w37785 = ~w37759 & ~w37783;
assign w37786 = ~w36258 & ~w37107;
assign w37787 = ~w37784 & ~w37785;
assign w37788 = w37107 & w37787;
assign w37789 = ~w37786 & ~w37788;
assign w37790 = ~w15681 & ~w37789;
assign w37791 = (w15681 & w37060) | (w15681 & w46250) | (w37060 & w46250);
assign w37792 = ~w36259 & ~w37784;
assign w37793 = w37107 & w37792;
assign w37794 = ~w37791 & ~w37793;
assign w37795 = w36287 & w36342;
assign w37796 = w14766 & ~w37795;
assign w37797 = (w37796 & w37793) | (w37796 & w46251) | (w37793 & w46251);
assign w37798 = w14766 & w37795;
assign w37799 = ~w37793 & w46252;
assign w37800 = ~w37797 & ~w37799;
assign w37801 = ~w36296 & w36301;
assign w37802 = w36333 & ~w37683;
assign w37803 = w36314 & ~w37802;
assign w37804 = w37801 & ~w37803;
assign w37805 = ~w37801 & w37803;
assign w37806 = ~w37804 & ~w37805;
assign w37807 = ~w36295 & ~w37107;
assign w37808 = w37107 & w37806;
assign w37809 = ~w37807 & ~w37808;
assign w37810 = ~w16559 & ~w37809;
assign w37811 = ~w14766 & w37795;
assign w37812 = (w37811 & w37793) | (w37811 & w46253) | (w37793 & w46253);
assign w37813 = ~w14766 & ~w37795;
assign w37814 = ~w37793 & w46254;
assign w37815 = ~w37812 & ~w37814;
assign w37816 = ~w37810 & w37815;
assign w37817 = w37790 & w37800;
assign w37818 = w37816 & ~w37817;
assign w37819 = ~w37780 & w46255;
assign w37820 = w37696 & w37819;
assign w37821 = ~w37663 & w37820;
assign w37822 = ~w37768 & ~w37769;
assign w37823 = ~w14039 & ~w37822;
assign w37824 = w15681 & w37789;
assign w37825 = w37815 & w37824;
assign w37826 = w37800 & ~w37825;
assign w37827 = ~w37823 & w37826;
assign w37828 = w37773 & ~w37827;
assign w37829 = ~w17380 & ~w37690;
assign w37830 = w16559 & w37809;
assign w37831 = ~w37829 & ~w37830;
assign w37832 = w37818 & ~w37831;
assign w37833 = w37756 & ~w37832;
assign w37834 = ~w37828 & w37833;
assign w37835 = w37782 & ~w37834;
assign w37836 = ~w37821 & ~w37835;
assign w37837 = ~w36422 & ~w36429;
assign w37838 = (w36573 & ~w36567) | (w36573 & w43131) | (~w36567 & w43131);
assign w37839 = w36387 & w36573;
assign w37840 = w36242 & w37839;
assign w37841 = ~w37838 & ~w37840;
assign w37842 = ~w36437 & ~w36553;
assign w37843 = w36465 & w36551;
assign w37844 = ~w36553 & ~w37843;
assign w37845 = ~w37841 & w37842;
assign w37846 = (w37844 & w37841) | (w37844 & w46256) | (w37841 & w46256);
assign w37847 = w37837 & w37846;
assign w37848 = ~w36410 & ~w36440;
assign w37849 = ~w36429 & w37848;
assign w37850 = ~w37847 & w37849;
assign w37851 = ~w36410 & ~w37850;
assign w37852 = w36448 & ~w36863;
assign w37853 = w37107 & ~w37852;
assign w37854 = ~w37851 & w37853;
assign w37855 = w37107 & w37852;
assign w37856 = w37851 & w37855;
assign w37857 = ~w37854 & ~w37856;
assign w37858 = ~w36862 & ~w37107;
assign w37859 = ~w5745 & ~w37858;
assign w37860 = w37857 & w37859;
assign w37861 = ~w36429 & ~w37847;
assign w37862 = ~w37848 & ~w37861;
assign w37863 = w37107 & ~w37850;
assign w37864 = ~w37862 & w37863;
assign w37865 = ~w36409 & ~w37107;
assign w37866 = w6264 & ~w37865;
assign w37867 = ~w37864 & w37866;
assign w37868 = ~w37860 & ~w37867;
assign w37869 = ~w37864 & ~w37865;
assign w37870 = ~w6264 & ~w37869;
assign w37871 = ~w37837 & ~w37846;
assign w37872 = ~w37847 & ~w37871;
assign w37873 = w37107 & ~w37872;
assign w37874 = ~w7315 & ~w36422;
assign w37875 = ~w36429 & ~w37874;
assign w37876 = (w37875 & w37060) | (w37875 & w46257) | (w37060 & w46257);
assign w37877 = ~w37873 & ~w37876;
assign w37878 = w6769 & ~w37877;
assign w37879 = ~w37870 & ~w37878;
assign w37880 = w37868 & ~w37879;
assign w37881 = ~w36576 & ~w36863;
assign w37882 = ~w36876 & ~w37072;
assign w37883 = (w37882 & w36576) | (w37882 & w46258) | (w36576 & w46258);
assign w37884 = w37107 & ~w37883;
assign w37885 = w37881 & ~w37882;
assign w37886 = w37884 & ~w37885;
assign w37887 = ~w36875 & ~w37107;
assign w37888 = ~w37886 & ~w37887;
assign w37889 = ~w5330 & ~w37888;
assign w37890 = w37857 & ~w37858;
assign w37891 = w5745 & ~w37890;
assign w37892 = ~w37889 & ~w37891;
assign w37893 = ~w37880 & w37892;
assign w37894 = w37841 & ~w37842;
assign w37895 = ~w37845 & ~w37894;
assign w37896 = (w36436 & w37060) | (w36436 & w46259) | (w37060 & w46259);
assign w37897 = w37107 & ~w37895;
assign w37898 = ~w37896 & ~w37897;
assign w37899 = (w7315 & w37897) | (w7315 & w46260) | (w37897 & w46260);
assign w37900 = ~w6769 & ~w37876;
assign w37901 = ~w37873 & w37900;
assign w37902 = ~w37899 & ~w37901;
assign w37903 = ~w37867 & w37902;
assign w37904 = ~w37860 & w37903;
assign w37905 = ~w7315 & w37898;
assign w37906 = ~w36464 & ~w36474;
assign w37907 = w36520 & ~w36549;
assign w37908 = (w37907 & w36567) | (w37907 & w43132) | (w36567 & w43132);
assign w37909 = ~w37700 & w37908;
assign w37910 = w35564 & ~w36503;
assign w37911 = ~w35564 & w36503;
assign w37912 = ~w37910 & ~w37911;
assign w37913 = w11138 & ~w37912;
assign w37914 = w36525 & ~w37913;
assign w37915 = w36545 & ~w37914;
assign w37916 = ~w36473 & ~w36538;
assign w37917 = w37915 & ~w37916;
assign w37918 = ~w36496 & w36538;
assign w37919 = ~w36473 & ~w37918;
assign w37920 = (w37919 & w37909) | (w37919 & w46261) | (w37909 & w46261);
assign w37921 = ~w37906 & w37920;
assign w37922 = w37906 & ~w37920;
assign w37923 = w36463 & ~w37107;
assign w37924 = w37107 & w46262;
assign w37925 = ~w37923 & ~w37924;
assign w37926 = ~w7924 & ~w37925;
assign w37927 = ~w37905 & ~w37926;
assign w37928 = w7924 & w37925;
assign w37929 = ~w36473 & ~w36536;
assign w37930 = (w36496 & w37909) | (w36496 & w46263) | (w37909 & w46263);
assign w37931 = ~w36537 & ~w37930;
assign w37932 = w37929 & ~w37931;
assign w37933 = ~w36537 & ~w37929;
assign w37934 = ~w37930 & w37933;
assign w37935 = w36472 & ~w37107;
assign w37936 = w37107 & ~w37934;
assign w37937 = ~w37932 & w37936;
assign w37938 = ~w37935 & ~w37937;
assign w37939 = ~w8666 & w37938;
assign w37940 = ~w37928 & w37939;
assign w37941 = w37927 & ~w37940;
assign w37942 = ~w36817 & w43133;
assign w37943 = ~w36576 & w37942;
assign w37944 = w37106 & w37912;
assign w37945 = ~w37943 & ~w37944;
assign w37946 = w36544 & ~w37913;
assign w37947 = ~w36514 & ~w37946;
assign w37948 = w36514 & w37946;
assign w37949 = ~w37947 & ~w37948;
assign w37950 = ~w37703 & w46264;
assign w37951 = (~w37949 & w37703) | (~w37949 & w46265) | (w37703 & w46265);
assign w37952 = ~w37950 & ~w37951;
assign w37953 = w37107 & w37952;
assign w37954 = w37945 & ~w37953;
assign w37955 = (w9781 & w37953) | (w9781 & w46266) | (w37953 & w46266);
assign w37956 = ~w9781 & w37945;
assign w37957 = ~w37953 & w37956;
assign w37958 = w36544 & ~w37914;
assign w37959 = ~w37909 & w37958;
assign w37960 = ~w37106 & ~w37959;
assign w37961 = ~w37060 & w37960;
assign w37962 = w36486 & ~w37961;
assign w37963 = ~w36486 & w37961;
assign w37964 = ~w37962 & ~w37963;
assign w37965 = ~w37957 & ~w37964;
assign w37966 = ~w36495 & ~w36537;
assign w37967 = w37915 & ~w37966;
assign w37968 = ~w36487 & w37966;
assign w37969 = (w37968 & w37909) | (w37968 & w46267) | (w37909 & w46267);
assign w37970 = w36487 & ~w37966;
assign w37971 = (~w37970 & w37909) | (~w37970 & w46268) | (w37909 & w46268);
assign w37972 = ~w37969 & w37971;
assign w37973 = (~w36494 & w37060) | (~w36494 & w46269) | (w37060 & w46269);
assign w37974 = w37107 & ~w37972;
assign w37975 = ~w37973 & ~w37974;
assign w37976 = (w9195 & w37974) | (w9195 & w46270) | (w37974 & w46270);
assign w37977 = ~w37060 & w46271;
assign w37978 = w36486 & ~w37977;
assign w37979 = ~w36486 & w37977;
assign w37980 = ~w37978 & ~w37979;
assign w37981 = ~w9781 & w10419;
assign w37982 = w37980 & w37981;
assign w37983 = ~w37976 & ~w37982;
assign w37984 = ~w37965 & w46272;
assign w37985 = w37983 & ~w37984;
assign w37986 = ~w9195 & w37975;
assign w37987 = (w8666 & w37937) | (w8666 & w46273) | (w37937 & w46273);
assign w37988 = ~w37928 & ~w37987;
assign w37989 = ~w37986 & w37988;
assign w37990 = ~w37985 & w37989;
assign w37991 = w37941 & ~w37990;
assign w37992 = w37904 & ~w37991;
assign w37993 = w37893 & ~w37992;
assign w37994 = w36556 & ~w37098;
assign w37995 = w36467 & ~w37098;
assign w37996 = w36573 & w37995;
assign w37997 = ~w37994 & ~w37996;
assign w37998 = (~w37997 & ~w36570) | (~w37997 & w43134) | (~w36570 & w43134);
assign w37999 = ~w36967 & ~w37098;
assign w38000 = ~w36856 & ~w37099;
assign w38001 = ~w37999 & w38000;
assign w38002 = ~w37998 & w38001;
assign w38003 = (~w37099 & w37998) | (~w37099 & w46274) | (w37998 & w46274);
assign w38004 = ~w36838 & ~w36852;
assign w38005 = w38003 & ~w38004;
assign w38006 = ~w38003 & w38004;
assign w38007 = w36837 & ~w37107;
assign w38008 = ~w38005 & ~w38006;
assign w38009 = w37107 & w38008;
assign w38010 = ~w38007 & ~w38009;
assign w38011 = ~w2558 & ~w38010;
assign w38012 = w36555 & w36925;
assign w38013 = ~w36936 & w36965;
assign w38014 = w38012 & ~w38013;
assign w38015 = w37841 & w38014;
assign w38016 = ~w36936 & w36964;
assign w38017 = ~w36439 & w36449;
assign w38018 = w36925 & ~w38017;
assign w38019 = ~w37087 & w37093;
assign w38020 = ~w36923 & ~w38019;
assign w38021 = ~w38018 & ~w38020;
assign w38022 = ~w36959 & ~w37088;
assign w38023 = ~w38018 & w46275;
assign w38024 = ~w36959 & ~w38023;
assign w38025 = ~w36959 & ~w38016;
assign w38026 = w38012 & w38025;
assign w38027 = w37841 & w38026;
assign w38028 = w38016 & ~w38024;
assign w38029 = ~w38015 & w38028;
assign w38030 = ~w38016 & w38024;
assign w38031 = ~w38027 & ~w38030;
assign w38032 = ~w38029 & w38031;
assign w38033 = w37107 & w38032;
assign w38034 = ~w36817 & w43135;
assign w38035 = ~w36576 & w38034;
assign w38036 = w36935 & w37106;
assign w38037 = ~w38035 & ~w38036;
assign w38038 = ~w3242 & w38037;
assign w38039 = ~w38033 & w38038;
assign w38040 = (~w38000 & w37996) | (~w38000 & w46276) | (w37996 & w46276);
assign w38041 = w37999 & ~w38000;
assign w38042 = (~w38041 & w36572) | (~w38041 & w43136) | (w36572 & w43136);
assign w38043 = ~w38002 & w38042;
assign w38044 = w37107 & ~w38043;
assign w38045 = ~w36855 & w37106;
assign w38046 = ~w36817 & w43137;
assign w38047 = ~w36576 & w38046;
assign w38048 = ~w38045 & ~w38047;
assign w38049 = w2896 & w38048;
assign w38050 = ~w38044 & w38049;
assign w38051 = ~w38039 & ~w38050;
assign w38052 = ~w2896 & ~w36855;
assign w38053 = ~w2896 & ~w37106;
assign w38054 = ~w37060 & w38053;
assign w38055 = ~w38052 & ~w38054;
assign w38056 = w37107 & w38043;
assign w38057 = ~w38055 & ~w38056;
assign w38058 = ~w38033 & w38037;
assign w38059 = (w3242 & w38033) | (w3242 & w46277) | (w38033 & w46277);
assign w38060 = w38012 & w38021;
assign w38061 = w38021 & ~w38022;
assign w38062 = ~w38021 & w38022;
assign w38063 = ~w38061 & ~w38062;
assign w38064 = w37841 & w46278;
assign w38065 = (~w38063 & ~w37841) | (~w38063 & w50393) | (~w37841 & w50393);
assign w38066 = ~w38064 & ~w38065;
assign w38067 = w37107 & w38066;
assign w38068 = ~w36958 & w37106;
assign w38069 = ~w36817 & w43138;
assign w38070 = ~w36576 & w38069;
assign w38071 = ~w38068 & ~w38070;
assign w38072 = w3646 & w38071;
assign w38073 = ~w38067 & w38072;
assign w38074 = ~w38051 & ~w38057;
assign w38075 = ~w38057 & ~w38073;
assign w38076 = ~w38059 & w38075;
assign w38077 = ~w38074 & ~w38076;
assign w38078 = w2558 & w38010;
assign w38079 = w2558 & ~w37107;
assign w38080 = ~w36838 & ~w37106;
assign w38081 = ~w37060 & w38080;
assign w38082 = ~w38006 & w38081;
assign w38083 = ~w38079 & ~w38082;
assign w38084 = ~w36850 & ~w36858;
assign w38085 = ~w2285 & w38084;
assign w38086 = w38083 & w38085;
assign w38087 = ~w2285 & ~w38084;
assign w38088 = ~w38083 & w38087;
assign w38089 = ~w38086 & ~w38088;
assign w38090 = ~w38078 & w38089;
assign w38091 = ~w38011 & w38077;
assign w38092 = w38090 & ~w38091;
assign w38093 = ~w36877 & w37086;
assign w38094 = w36909 & ~w38093;
assign w38095 = (w36570 & w46279) | (w36570 & w46280) | (w46279 & w46280);
assign w38096 = (~w36891 & w37060) | (~w36891 & w46281) | (w37060 & w46281);
assign w38097 = ~w37090 & w38095;
assign w38098 = w37107 & w38097;
assign w38099 = ~w38096 & ~w38098;
assign w38100 = w36908 & ~w38093;
assign w38101 = (w36570 & w46282) | (w36570 & w46283) | (w46282 & w46283);
assign w38102 = ~w36892 & ~w37090;
assign w38103 = ~w38101 & ~w38102;
assign w38104 = w37107 & w38103;
assign w38105 = (w4430 & ~w37107) | (w4430 & w46284) | (~w37107 & w46284);
assign w38106 = (~w4056 & ~w38099) | (~w4056 & w46285) | (~w38099 & w46285);
assign w38107 = w4430 & w36922;
assign w38108 = ~w36923 & ~w38107;
assign w38109 = (~w4430 & w37060) | (~w4430 & w43141) | (w37060 & w43141);
assign w38110 = ~w37090 & ~w38095;
assign w38111 = w37107 & w38110;
assign w38112 = ~w38111 & w43142;
assign w38113 = (~w38108 & w38111) | (~w38108 & w43143) | (w38111 & w43143);
assign w38114 = ~w38112 & ~w38113;
assign w38115 = ~w38106 & w38114;
assign w38116 = ~w38067 & w38071;
assign w38117 = ~w3646 & ~w38116;
assign w38118 = w38051 & ~w38117;
assign w38119 = ~w38115 & w38118;
assign w38120 = w38099 & ~w38104;
assign w38121 = w38099 & w43144;
assign w38122 = w4430 & w38121;
assign w38123 = ~w38011 & ~w38122;
assign w38124 = w38119 & w38123;
assign w38125 = w38092 & ~w38124;
assign w38126 = w37107 & w46286;
assign w38127 = w5330 & ~w37107;
assign w38128 = ~w38126 & ~w38127;
assign w38129 = w36908 & w37085;
assign w38130 = w4838 & ~w38129;
assign w38131 = ~w38126 & w43145;
assign w38132 = w4838 & w38129;
assign w38133 = (w38132 & w38126) | (w38132 & w43146) | (w38126 & w43146);
assign w38134 = ~w38131 & ~w38133;
assign w38135 = w4430 & w38134;
assign w38136 = ~w38120 & ~w38135;
assign w38137 = ~w4056 & ~w38114;
assign w38138 = w38134 & ~w38137;
assign w38139 = w38092 & w43147;
assign w38140 = ~w38125 & ~w38139;
assign w38141 = w37993 & ~w38140;
assign w38142 = w37836 & w38141;
assign w38143 = w10419 & ~w37957;
assign w38144 = ~w37976 & w38143;
assign w38145 = ~w37955 & w37980;
assign w38146 = w38144 & ~w38145;
assign w38147 = w36539 & w37958;
assign w38148 = ~w37909 & w38147;
assign w38149 = ~w37106 & w38148;
assign w38150 = ~w37060 & w38149;
assign w38151 = w9781 & ~w38150;
assign w38152 = w10419 & ~w36486;
assign w38153 = (w38152 & w37060) | (w38152 & w43148) | (w37060 & w43148);
assign w38154 = w38151 & ~w38153;
assign w38155 = w36487 & ~w37961;
assign w38156 = ~w36487 & ~w36539;
assign w38157 = w37961 & w38156;
assign w38158 = ~w38155 & ~w38157;
assign w38159 = w38154 & w38158;
assign w38160 = ~w37976 & w38159;
assign w38161 = ~w37986 & ~w38160;
assign w38162 = ~w38146 & w38161;
assign w38163 = w37927 & ~w37939;
assign w38164 = ~w38162 & w38163;
assign w38165 = w37927 & ~w37988;
assign w38166 = w37904 & ~w38165;
assign w38167 = ~w38164 & w38166;
assign w38168 = w37893 & ~w38167;
assign w38169 = w5330 & w37888;
assign w38170 = w38128 & ~w38129;
assign w38171 = ~w38128 & w38129;
assign w38172 = ~w38170 & ~w38171;
assign w38173 = ~w4838 & w38172;
assign w38174 = ~w38169 & ~w38173;
assign w38175 = (w38174 & ~w38092) | (w38174 & w46287) | (~w38092 & w46287);
assign w38176 = ~w38168 & w38175;
assign w38177 = ~w38140 & ~w38176;
assign w38178 = w2285 & w38084;
assign w38179 = ~w37107 & w43149;
assign w38180 = w38081 & w38178;
assign w38181 = ~w38006 & w38180;
assign w38182 = ~w38179 & ~w38181;
assign w38183 = w2285 & ~w38084;
assign w38184 = (w38183 & w37107) | (w38183 & w43150) | (w37107 & w43150);
assign w38185 = ~w38082 & w38184;
assign w38186 = w2006 & w37272;
assign w38187 = ~w38185 & ~w38186;
assign w38188 = w37254 & w38182;
assign w38189 = w38187 & w38188;
assign w38190 = ~w37224 & ~w37248;
assign w38191 = ~w37224 & ~w38189;
assign w38192 = w37286 & w38191;
assign w38193 = ~w38190 & ~w38192;
assign w38194 = w37194 & w38193;
assign w38195 = ~w37299 & ~w38194;
assign w38196 = ~w38177 & ~w38195;
assign w38197 = ~w38142 & w38196;
assign w38198 = w36807 & ~w37070;
assign w38199 = ~w36817 & ~w37057;
assign w38200 = (w38199 & w37112) | (w38199 & w43151) | (w37112 & w43151);
assign w38201 = (~w57 & w37060) | (~w57 & w43152) | (w37060 & w43152);
assign w38202 = ~w38200 & ~w38201;
assign w38203 = w37013 & ~w37038;
assign w38204 = w80 & ~w38203;
assign w38205 = ~w80 & w38203;
assign w38206 = ~w38204 & ~w38205;
assign w38207 = w38202 & ~w38206;
assign w38208 = ~w38202 & w38206;
assign w38209 = ~w38207 & ~w38208;
assign w38210 = w80 & w38209;
assign w38211 = ~w36817 & ~w37038;
assign w38212 = (w38211 & w37112) | (w38211 & w43153) | (w37112 & w43153);
assign w38213 = ~w80 & ~w37107;
assign w38214 = ~w37060 & w43154;
assign w38215 = ~w38212 & w38214;
assign w38216 = ~w38213 & ~w38215;
assign w38217 = w36984 & ~w36999;
assign w38218 = w38216 & ~w38217;
assign w38219 = ~w38216 & w38217;
assign w38220 = ~w38218 & ~w38219;
assign w38221 = w3 & w38220;
assign w38222 = ~w3 & ~w38220;
assign w38223 = ~w37020 & w37030;
assign w38224 = w37014 & ~w38223;
assign w38225 = ~w38212 & w38224;
assign w38226 = ~w36996 & w37020;
assign w38227 = ~w42 & w37050;
assign w38228 = w37030 & ~w38227;
assign w38229 = w37014 & w37020;
assign w38230 = w38226 & ~w38228;
assign w38231 = ~w38228 & w38229;
assign w38232 = ~w38212 & w38231;
assign w38233 = ~w38230 & ~w38232;
assign w38234 = w37030 & ~w38226;
assign w38235 = ~w38225 & w38234;
assign w38236 = w38233 & ~w38235;
assign w38237 = ~w42 & ~w38236;
assign w38238 = w36984 & w37107;
assign w38239 = w37014 & ~w38212;
assign w38240 = w38238 & ~w38239;
assign w38241 = (~w3 & w37060) | (~w3 & w43155) | (w37060 & w43155);
assign w38242 = w36995 & w37020;
assign w38243 = w38241 & ~w38242;
assign w38244 = ~w38241 & w38242;
assign w38245 = ~w38243 & ~w38244;
assign w38246 = w38240 & ~w38245;
assign w38247 = ~w38240 & w38245;
assign w38248 = ~w38246 & ~w38247;
assign w38249 = w38237 & w38248;
assign w38250 = ~w38222 & ~w38249;
assign w38251 = w38210 & ~w38221;
assign w38252 = w38250 & ~w38251;
assign w38253 = (w351 & w37303) | (w351 & w43156) | (w37303 & w43156);
assign w38254 = w37308 & w38253;
assign w38255 = ~w36762 & ~w36802;
assign w38256 = w36804 & ~w38255;
assign w38257 = ~w36814 & ~w38256;
assign w38258 = ~w36747 & ~w38255;
assign w38259 = (w38257 & w37115) | (w38257 & w43157) | (w37115 & w43157);
assign w38260 = w38258 & ~w38259;
assign w38261 = (~w36761 & w37060) | (~w36761 & w43158) | (w37060 & w43158);
assign w38262 = ~w252 & ~w38261;
assign w38263 = ~w36747 & w37107;
assign w38264 = ~w37303 & w38263;
assign w38265 = ~w36762 & w36805;
assign w38266 = w37107 & ~w38265;
assign w38267 = w38260 & w38262;
assign w38268 = w38262 & ~w38266;
assign w38269 = ~w38264 & w38268;
assign w38270 = ~w38267 & ~w38269;
assign w38271 = ~w38254 & w38270;
assign w38272 = w36747 & ~w36802;
assign w38273 = ~w36762 & ~w38272;
assign w38274 = w36805 & ~w36814;
assign w38275 = w37301 & w38273;
assign w38276 = (w38275 & w37112) | (w38275 & w43159) | (w37112 & w43159);
assign w38277 = w38273 & ~w38274;
assign w38278 = ~w38276 & ~w38277;
assign w38279 = ~w37060 & w43160;
assign w38280 = w36800 & ~w38279;
assign w38281 = w36801 & w37107;
assign w38282 = ~w38280 & ~w38281;
assign w38283 = ~w37060 & w43161;
assign w38284 = w36800 & ~w38283;
assign w38285 = ~w36800 & w38283;
assign w38286 = w38278 & w38282;
assign w38287 = ~w38278 & ~w38284;
assign w38288 = ~w38285 & w38287;
assign w38289 = ~w38286 & ~w38288;
assign w38290 = ~w57 & ~w38289;
assign w38291 = w38271 & ~w38290;
assign w38292 = w38252 & w38291;
assign w38293 = ~w35994 & w37107;
assign w38294 = w35994 & ~w37107;
assign w38295 = ~w38293 & ~w38294;
assign w38296 = ~w37382 & w38295;
assign w38297 = w37381 & ~w38295;
assign w38298 = ~w38296 & ~w38297;
assign w38299 = w42 & ~w38248;
assign w38300 = ~w42 & w38236;
assign w38301 = w42 & w37107;
assign w38302 = ~w38236 & w38301;
assign w38303 = ~w38300 & ~w38302;
assign w38304 = ~w38299 & w38303;
assign w38305 = w57 & w38289;
assign w38306 = w38260 & ~w38261;
assign w38307 = ~w38261 & ~w38266;
assign w38308 = ~w38264 & w38307;
assign w38309 = ~w38306 & ~w38308;
assign w38310 = w57 & w36801;
assign w38311 = w37107 & w38310;
assign w38312 = ~w36781 & ~w38311;
assign w38313 = ~w38278 & w38285;
assign w38314 = ~w377 & ~w38313;
assign w38315 = w38278 & ~w38312;
assign w38316 = w38314 & ~w38315;
assign w38317 = w38309 & ~w38316;
assign w38318 = ~w38305 & ~w38317;
assign w38319 = ~w80 & w38209;
assign w38320 = w36781 & w38261;
assign w38321 = ~w38319 & ~w38320;
assign w38322 = ~w38221 & w38321;
assign w38323 = w38318 & w38322;
assign w38324 = w38252 & ~w38323;
assign w38325 = w38304 & ~w38324;
assign w38326 = w36044 & w37107;
assign w38327 = w38325 & w38326;
assign w38328 = w38292 & w38298;
assign w38329 = w38327 & w52290;
assign w38330 = ~w38252 & w38304;
assign w38331 = ~w38291 & w38304;
assign w38332 = w38323 & w38331;
assign w38333 = ~w38330 & ~w38332;
assign w38334 = ~w38195 & w38333;
assign w38335 = ~w38177 & w38334;
assign w38336 = ~w38142 & w38335;
assign w38337 = (w38292 & ~w37314) | (w38292 & w43163) | (~w37314 & w43163);
assign w38338 = w38325 & ~w38337;
assign w38339 = ~w38336 & w38338;
assign w38340 = ~a[4] & w37107;
assign w38341 = ~a[3] & a[4];
assign w38342 = ~w38293 & ~w38341;
assign w38343 = ~a[0] & ~a[1];
assign w38344 = ~a[2] & w38343;
assign w38345 = ~w38294 & w38344;
assign w38346 = ~w38342 & w38345;
assign w38347 = a[4] & w38293;
assign w38348 = ~w38346 & ~w38347;
assign w38349 = a[3] & ~w38344;
assign w38350 = ~a[3] & w38344;
assign w38351 = w35994 & ~w38350;
assign w38352 = ~a[4] & ~w38351;
assign w38353 = w37107 & ~w38349;
assign w38354 = ~w38352 & ~w38353;
assign w38355 = ~a[3] & w38293;
assign w38356 = ~w38340 & ~w38354;
assign w38357 = ~w38355 & ~w38356;
assign w38358 = w38348 & w38357;
assign w38359 = w34900 & w38358;
assign w38360 = a[5] & ~w38340;
assign w38361 = ~w38359 & ~w38360;
assign w38362 = ~a[4] & ~w38294;
assign w38363 = w38349 & ~w38362;
assign w38364 = a[4] & w35994;
assign w38365 = ~w37382 & ~w38364;
assign w38366 = ~w38363 & w38365;
assign w38367 = w38348 & ~w38366;
assign w38368 = w37382 & ~w38295;
assign w38369 = ~w38296 & ~w38368;
assign w38370 = w35994 & ~w37381;
assign w38371 = a[5] & ~w38370;
assign w38372 = ~w35994 & w37381;
assign w38373 = w38371 & ~w38372;
assign w38374 = w38340 & w38373;
assign w38375 = ~a[5] & ~w38369;
assign w38376 = w38360 & w38369;
assign w38377 = ~w38375 & ~w38376;
assign w38378 = ~w38374 & w38377;
assign w38379 = w34900 & w38367;
assign w38380 = w38378 & ~w38379;
assign w38381 = ~w38336 & w43164;
assign w38382 = (w38380 & w38336) | (w38380 & w43165) | (w38336 & w43165);
assign w38383 = ~w38381 & ~w38382;
assign w38384 = ~w37107 & w37414;
assign w38385 = w37107 & ~w37423;
assign w38386 = ~w38384 & ~w38385;
assign w38387 = w32698 & ~w38386;
assign w38388 = ~w33731 & ~w37402;
assign w38389 = ~w38387 & ~w38388;
assign w38390 = ~w34900 & ~w38358;
assign w38391 = w38389 & ~w38390;
assign w38392 = ~w37394 & w37402;
assign w38393 = w37429 & w38387;
assign w38394 = ~w33731 & ~w38392;
assign w38395 = ~w38393 & ~w38394;
assign w38396 = w37411 & ~w38387;
assign w38397 = ~w33731 & ~w38396;
assign w38398 = w37403 & ~w38397;
assign w38399 = ~w38395 & ~w38398;
assign w38400 = w37402 & ~w38387;
assign w38401 = ~w34900 & ~w38367;
assign w38402 = w37411 & w38399;
assign w38403 = ~w38401 & ~w38402;
assign w38404 = w38399 & ~w38400;
assign w38405 = ~w38404 & w52291;
assign w38406 = ~w38336 & w48078;
assign w38407 = w38405 & ~w38406;
assign w38408 = ~w38329 & ~w38383;
assign w38409 = w38407 & ~w38408;
assign w38410 = ~w37402 & ~w37411;
assign w38411 = ~w38386 & ~w38392;
assign w38412 = w34990 & ~w38411;
assign w38413 = ~w37403 & w37411;
assign w38414 = ~w37428 & ~w38413;
assign w38415 = w33731 & ~w38410;
assign w38416 = w32698 & ~w38415;
assign w38417 = ~w38414 & ~w38416;
assign w38418 = ~w37430 & w38417;
assign w38419 = ~w38412 & ~w38418;
assign w38420 = ~w37460 & w38410;
assign w38421 = ~w38419 & ~w38420;
assign w38422 = ~w32698 & w38386;
assign w38423 = w33731 & w38400;
assign w38424 = ~w38422 & ~w38423;
assign w38425 = ~w37460 & w38392;
assign w38426 = ~w38336 & w46288;
assign w38427 = ~w38425 & ~w38426;
assign w38428 = ~w38339 & w38421;
assign w38429 = w38427 & ~w38428;
assign w38430 = ~w37430 & w37460;
assign w38431 = w32698 & ~w38430;
assign w38432 = ~w32698 & w38430;
assign w38433 = ~w38431 & ~w38432;
assign w38434 = ~w37446 & w52292;
assign w38435 = (w38336 & w46289) | (w38336 & w46290) | (w46289 & w46290);
assign w38436 = ~w38434 & ~w38435;
assign w38437 = w33731 & w38413;
assign w38438 = w38431 & ~w38437;
assign w38439 = ~w38339 & w38438;
assign w38440 = ~w31477 & w38436;
assign w38441 = ~w38439 & ~w38440;
assign w38442 = ~w38409 & w38429;
assign w38443 = w38441 & ~w38442;
assign w38444 = ~w37473 & ~w37489;
assign w38445 = ~w37463 & ~w37485;
assign w38446 = w38444 & ~w38445;
assign w38447 = ~w38444 & w38445;
assign w38448 = ~w38446 & ~w38447;
assign w38449 = ~w37487 & ~w37489;
assign w38450 = ~w29158 & w38449;
assign w38451 = w29158 & ~w38449;
assign w38452 = ~w38450 & ~w38451;
assign w38453 = (w38452 & w38336) | (w38452 & w43168) | (w38336 & w43168);
assign w38454 = ~w30239 & ~w38448;
assign w38455 = (w38336 & w46291) | (w38336 & w46292) | (w46291 & w46292);
assign w38456 = ~w38336 & w43169;
assign w38457 = (w38448 & w38336) | (w38448 & w43170) | (w38336 & w43170);
assign w38458 = ~w38456 & ~w38457;
assign w38459 = w29158 & w38458;
assign w38460 = ~w28077 & w37492;
assign w38461 = w38455 & w38460;
assign w38462 = ~w28077 & ~w37492;
assign w38463 = ~w38455 & w38462;
assign w38464 = ~w38459 & w46293;
assign w38465 = w37478 & ~w38430;
assign w38466 = ~w37447 & ~w38465;
assign w38467 = ~w31477 & w38466;
assign w38468 = w31477 & ~w38466;
assign w38469 = ~w38467 & ~w38468;
assign w38470 = w36035 & ~w37450;
assign w38471 = ~w36035 & w37450;
assign w38472 = ~w38470 & ~w38471;
assign w38473 = (w38336 & w46294) | (w38336 & w46295) | (w46294 & w46295);
assign w38474 = w38472 & w52293;
assign w38475 = ~w38473 & ~w38474;
assign w38476 = w31477 & ~w38436;
assign w38477 = w30239 & w38475;
assign w38478 = ~w38476 & ~w38477;
assign w38479 = w38464 & w38478;
assign w38480 = ~w38443 & w38479;
assign w38481 = ~w29158 & ~w38458;
assign w38482 = ~w30239 & ~w38475;
assign w38483 = ~w38481 & ~w38482;
assign w38484 = w37377 & ~w37513;
assign w38485 = (w37369 & w37487) | (w37369 & w43172) | (w37487 & w43172);
assign w38486 = ~w38336 & w46296;
assign w38487 = (w38485 & w38336) | (w38485 & w43173) | (w38336 & w43173);
assign w38488 = ~w38486 & ~w38487;
assign w38489 = (~w38484 & w38486) | (~w38484 & w43174) | (w38486 & w43174);
assign w38490 = ~w26880 & ~w38489;
assign w38491 = w38484 & w38488;
assign w38492 = w38490 & ~w38491;
assign w38493 = w36098 & ~w37107;
assign w38494 = w37107 & w37324;
assign w38495 = ~w38493 & ~w38494;
assign w38496 = ~w37333 & ~w37504;
assign w38497 = (w37487 & w37378) | (w37487 & w46297) | (w37378 & w46297);
assign w38498 = ~w37513 & ~w38497;
assign w38499 = w38496 & ~w38498;
assign w38500 = ~w38496 & w38498;
assign w38501 = ~w38499 & ~w38500;
assign w38502 = (~w38336 & w46298) | (~w38336 & w46299) | (w46298 & w46299);
assign w38503 = ~w38336 & w48079;
assign w38504 = w38502 & ~w38503;
assign w38505 = w37514 & ~w38497;
assign w38506 = ~w37333 & ~w38505;
assign w38507 = w25851 & ~w38506;
assign w38508 = ~w25851 & w38506;
assign w38509 = ~w38507 & ~w38508;
assign w38510 = (w38509 & w38336) | (w38509 & w43176) | (w38336 & w43176);
assign w38511 = w24874 & w37341;
assign w38512 = (~w38336 & w46300) | (~w38336 & w46301) | (w46300 & w46301);
assign w38513 = w24874 & ~w37341;
assign w38514 = (w38336 & w46302) | (w38336 & w46303) | (w46302 & w46303);
assign w38515 = ~w38512 & ~w38514;
assign w38516 = ~w38504 & w38515;
assign w38517 = (w38336 & w46304) | (w38336 & w46305) | (w46304 & w46305);
assign w38518 = w28077 & ~w38517;
assign w38519 = ~w37492 & ~w38453;
assign w38520 = w38518 & ~w38519;
assign w38521 = w38516 & ~w38520;
assign w38522 = ~w38492 & w38521;
assign w38523 = w38464 & ~w38483;
assign w38524 = w38522 & ~w38523;
assign w38525 = ~w37810 & ~w37831;
assign w38526 = (~w38525 & w37663) | (~w38525 & w43178) | (w37663 & w43178);
assign w38527 = (w37663 & w46306) | (w37663 & w46307) | (w46306 & w46307);
assign w38528 = ~w14766 & ~w37824;
assign w38529 = ~w37790 & ~w38526;
assign w38530 = w38528 & ~w38529;
assign w38531 = w14766 & ~w37790;
assign w38532 = ~w38527 & w38531;
assign w38533 = ~w38530 & ~w38532;
assign w38534 = w37794 & ~w37795;
assign w38535 = ~w37794 & w37795;
assign w38536 = ~w38534 & ~w38535;
assign w38537 = ~w38339 & w43179;
assign w38538 = (w38536 & w38339) | (w38536 & w43180) | (w38339 & w43180);
assign w38539 = ~w38537 & ~w38538;
assign w38540 = w14039 & w38539;
assign w38541 = ~w37810 & ~w37830;
assign w38542 = (w37663 & w46308) | (w37663 & w46309) | (w46308 & w46309);
assign w38543 = w38541 & w52294;
assign w38544 = ~w38542 & ~w38543;
assign w38545 = ~w38336 & w43183;
assign w38546 = (w38544 & w38336) | (w38544 & w43184) | (w38336 & w43184);
assign w38547 = ~w38545 & ~w38546;
assign w38548 = w14766 & ~w37789;
assign w38549 = (w38336 & w46310) | (w38336 & w46311) | (w46310 & w46311);
assign w38550 = w38547 & ~w38549;
assign w38551 = w15681 & ~w37789;
assign w38552 = (w38336 & w46312) | (w38336 & w46313) | (w46312 & w46313);
assign w38553 = ~w17230 & ~w38552;
assign w38554 = ~w38550 & ~w38553;
assign w38555 = ~w15681 & w38526;
assign w38556 = (~w38555 & w38336) | (~w38555 & w43185) | (w38336 & w43185);
assign w38557 = w14766 & w37789;
assign w38558 = ~w38556 & w38557;
assign w38559 = w14766 & w37790;
assign w38560 = w38556 & w38559;
assign w38561 = ~w38558 & ~w38560;
assign w38562 = w37824 & w52295;
assign w38563 = w14766 & ~w38526;
assign w38564 = ~w37809 & ~w38563;
assign w38565 = ~w38336 & w43186;
assign w38566 = ~w38544 & ~w38563;
assign w38567 = (w38566 & w38336) | (w38566 & w46314) | (w38336 & w46314);
assign w38568 = ~w38565 & ~w38567;
assign w38569 = w38562 & w38568;
assign w38570 = w38561 & ~w38569;
assign w38571 = (~w38540 & ~w38570) | (~w38540 & w43187) | (~w38570 & w43187);
assign w38572 = w37826 & w37831;
assign w38573 = (w38572 & w37678) | (w38572 & w46315) | (w37678 & w46315);
assign w38574 = w37662 & w38572;
assign w38575 = w37538 & w38574;
assign w38576 = ~w38573 & ~w38575;
assign w38577 = ~w37818 & w37826;
assign w38578 = ~w37771 & ~w38577;
assign w38579 = (w38575 & w46316) | (w38575 & w46317) | (w46316 & w46317);
assign w38580 = ~w13384 & w38579;
assign w38581 = w13384 & ~w37771;
assign w38582 = ~w38579 & w38581;
assign w38583 = ~w38580 & ~w38582;
assign w38584 = (w37753 & w38339) | (w37753 & w43189) | (w38339 & w43189);
assign w38585 = ~w37753 & ~w37823;
assign w38586 = (w38575 & w46318) | (w38575 & w46319) | (w46318 & w46319);
assign w38587 = ~w37772 & ~w38586;
assign w38588 = ~w38580 & ~w38587;
assign w38589 = (w38588 & w38336) | (w38588 & w46320) | (w38336 & w46320);
assign w38590 = ~w37746 & ~w37775;
assign w38591 = ~w38580 & w38587;
assign w38592 = ~w38336 & w43191;
assign w38593 = (w38591 & w38336) | (w38591 & w46321) | (w38336 & w46321);
assign w38594 = ~w38592 & ~w38593;
assign w38595 = ~w11870 & ~w37775;
assign w38596 = w37746 & ~w38587;
assign w38597 = w38595 & ~w38596;
assign w38598 = ~w38593 & w43192;
assign w38599 = ~w11870 & ~w38590;
assign w38600 = (w38599 & w38593) | (w38599 & w43193) | (w38593 & w43193);
assign w38601 = ~w38598 & ~w38600;
assign w38602 = (~w12666 & w38584) | (~w12666 & w46322) | (w38584 & w46322);
assign w38603 = w38601 & ~w38602;
assign w38604 = w38576 & ~w38577;
assign w38605 = ~w37771 & ~w37823;
assign w38606 = w38604 & ~w38605;
assign w38607 = ~w38604 & w38605;
assign w38608 = ~w38606 & ~w38607;
assign w38609 = ~w38336 & w46323;
assign w38610 = ~w38339 & w38608;
assign w38611 = ~w14039 & ~w38539;
assign w38612 = ~w38610 & w46324;
assign w38613 = ~w38611 & ~w38612;
assign w38614 = w38603 & w38613;
assign w38615 = ~w38571 & w38614;
assign w38616 = (w22767 & w37538) | (w22767 & w43194) | (w37538 & w43194);
assign w38617 = ~w37673 & ~w38616;
assign w38618 = ~w37538 & w43195;
assign w38619 = (~w37621 & w37538) | (~w37621 & w46325) | (w37538 & w46325);
assign w38620 = ~w38617 & w38619;
assign w38621 = w20906 & ~w37591;
assign w38622 = ~w38620 & w38621;
assign w38623 = ~w20906 & w38620;
assign w38624 = w37107 & ~w37579;
assign w38625 = ~w37107 & w37583;
assign w38626 = ~w38624 & ~w38625;
assign w38627 = w38623 & w38626;
assign w38628 = ~w38622 & ~w38627;
assign w38629 = ~w36183 & ~w37107;
assign w38630 = w37107 & w37560;
assign w38631 = ~w38629 & ~w38630;
assign w38632 = w20000 & w38631;
assign w38633 = ~w38628 & w38632;
assign w38634 = w20000 & ~w38631;
assign w38635 = ~w20906 & w37591;
assign w38636 = ~w38622 & ~w38635;
assign w38637 = ~w38623 & ~w38634;
assign w38638 = w38636 & ~w38637;
assign w38639 = ~w37621 & ~w38635;
assign w38640 = ~w38634 & w38639;
assign w38641 = ~w38621 & ~w38640;
assign w38642 = ~w38617 & ~w38618;
assign w38643 = w38641 & ~w38642;
assign w38644 = ~w37591 & ~w38620;
assign w38645 = w37565 & ~w37634;
assign w38646 = w20000 & ~w38645;
assign w38647 = ~w38644 & ~w38646;
assign w38648 = ~w20000 & ~w37634;
assign w38649 = ~w36172 & ~w37107;
assign w38650 = w37107 & w37549;
assign w38651 = ~w38649 & ~w38650;
assign w38652 = ~w38648 & w38651;
assign w38653 = ~w19040 & w38652;
assign w38654 = ~w38645 & ~w38653;
assign w38655 = ~w20000 & ~w38654;
assign w38656 = ~w37566 & ~w38648;
assign w38657 = ~w38651 & ~w38656;
assign w38658 = ~w37565 & ~w37571;
assign w38659 = ~w38657 & ~w38658;
assign w38660 = ~w19040 & ~w38659;
assign w38661 = ~w38655 & ~w38660;
assign w38662 = w21009 & ~w38651;
assign w38663 = w38645 & ~w38662;
assign w38664 = ~w38653 & w38663;
assign w38665 = ~w38644 & w38664;
assign w38666 = ~w38647 & w38661;
assign w38667 = ~w38665 & ~w38666;
assign w38668 = ~w38638 & ~w38643;
assign w38669 = ~w38633 & w38668;
assign w38670 = ~w38667 & ~w38669;
assign w38671 = w37565 & ~w37591;
assign w38672 = ~w38620 & w38671;
assign w38673 = ~w37634 & ~w38672;
assign w38674 = w19040 & w38651;
assign w38675 = w18183 & ~w37658;
assign w38676 = ~w38674 & ~w38675;
assign w38677 = ~w20421 & ~w37554;
assign w38678 = ~w37692 & w38677;
assign w38679 = w21010 & ~w38676;
assign w38680 = ~w38678 & ~w38679;
assign w38681 = ~w37691 & ~w37829;
assign w38682 = (w38681 & w37663) | (w38681 & w43196) | (w37663 & w43196);
assign w38683 = ~w37663 & w43197;
assign w38684 = ~w38682 & ~w38683;
assign w38685 = w16559 & ~w38684;
assign w38686 = (~w38685 & w38336) | (~w38685 & w43198) | (w38336 & w43198);
assign w38687 = (~w37639 & w37538) | (~w37639 & w43199) | (w37538 & w43199);
assign w38688 = (w37538 & w46326) | (w37538 & w46327) | (w46326 & w46327);
assign w38689 = ~w37692 & ~w38688;
assign w38690 = ~w37648 & ~w37649;
assign w38691 = ~w37658 & w38674;
assign w38692 = w37692 & ~w38687;
assign w38693 = ~w38691 & ~w38692;
assign w38694 = w18183 & ~w38693;
assign w38695 = ~w17380 & w38690;
assign w38696 = ~w38689 & w38695;
assign w38697 = ~w17380 & ~w38690;
assign w38698 = w38689 & w38697;
assign w38699 = ~w38694 & ~w38698;
assign w38700 = ~w38696 & w38699;
assign w38701 = ~w38673 & ~w38680;
assign w38702 = w38686 & w46328;
assign w38703 = ~w37659 & ~w37692;
assign w38704 = w19040 & w37554;
assign w38705 = w18183 & w38703;
assign w38706 = ~w38704 & ~w38705;
assign w38707 = w37571 & ~w38706;
assign w38708 = w38673 & w38707;
assign w38709 = w37520 & ~w38497;
assign w38710 = w37345 & ~w38709;
assign w38711 = w37355 & ~w38710;
assign w38712 = ~w23843 & ~w38711;
assign w38713 = w37523 & w38507;
assign w38714 = ~w37355 & ~w37523;
assign w38715 = ~w38507 & w38714;
assign w38716 = w38712 & ~w38715;
assign w38717 = ~w38713 & w38716;
assign w38718 = w21801 & ~w37673;
assign w38719 = ~w22767 & ~w37666;
assign w38720 = ~w38616 & ~w38618;
assign w38721 = ~w38719 & w38720;
assign w38722 = w38718 & ~w38721;
assign w38723 = w21801 & w37673;
assign w38724 = (w38723 & w37538) | (w38723 & w46329) | (w37538 & w46329);
assign w38725 = w37534 & ~w37667;
assign w38726 = ~w37522 & ~w37523;
assign w38727 = ~w37495 & w38726;
assign w38728 = ~w37488 & w38727;
assign w38729 = w38725 & w38728;
assign w38730 = ~w38724 & ~w38729;
assign w38731 = ~w22767 & ~w38725;
assign w38732 = ~w38728 & w38731;
assign w38733 = ~w38616 & ~w38730;
assign w38734 = ~w38732 & ~w38733;
assign w38735 = ~w38722 & w38734;
assign w38736 = ~w26445 & w37341;
assign w38737 = ~w37355 & w38736;
assign w38738 = w38509 & w38737;
assign w38739 = ~w38708 & ~w38717;
assign w38740 = w38735 & ~w38738;
assign w38741 = w38739 & w38740;
assign w38742 = w38702 & w38741;
assign w38743 = ~w38670 & w38742;
assign w38744 = ~w38718 & ~w38719;
assign w38745 = ~w20000 & w38631;
assign w38746 = ~w19040 & ~w38651;
assign w38747 = ~w38745 & ~w38746;
assign w38748 = ~w20906 & ~w38626;
assign w38749 = ~w38634 & ~w38748;
assign w38750 = w38747 & ~w38749;
assign w38751 = w38676 & ~w38750;
assign w38752 = ~w23843 & w37354;
assign w38753 = ~w17380 & w37647;
assign w38754 = w16559 & ~w37690;
assign w38755 = ~w38753 & ~w38754;
assign w38756 = w38744 & w38751;
assign w38757 = ~w38752 & w38755;
assign w38758 = w38756 & w38757;
assign w38759 = w38339 & w38758;
assign w38760 = ~w38743 & ~w38759;
assign w38761 = w26880 & w38484;
assign w38762 = ~w38485 & w38761;
assign w38763 = ~w25851 & w38501;
assign w38764 = ~w38762 & ~w38763;
assign w38765 = ~w25851 & w38495;
assign w38766 = w28077 & w38761;
assign w38767 = ~w38765 & ~w38766;
assign w38768 = (w38764 & w38336) | (w38764 & w46330) | (w38336 & w46330);
assign w38769 = ~w38336 & w46331;
assign w38770 = ~w38768 & ~w38769;
assign w38771 = w26880 & ~w38484;
assign w38772 = (w38771 & w38486) | (w38771 & w43200) | (w38486 & w43200);
assign w38773 = ~w38770 & ~w38772;
assign w38774 = ~w24874 & ~w37341;
assign w38775 = ~w38510 & w38774;
assign w38776 = (~w38775 & ~w38516) | (~w38775 & w46332) | (~w38516 & w46332);
assign w38777 = ~w38760 & w38776;
assign w38778 = w38615 & w38777;
assign w38779 = ~w38480 & w38524;
assign w38780 = w38778 & ~w38779;
assign w38781 = ~w38711 & w38728;
assign w38782 = w23843 & ~w38781;
assign w38783 = ~w23843 & w38728;
assign w38784 = w23843 & w37354;
assign w38785 = w38710 & w38784;
assign w38786 = ~w38783 & ~w38785;
assign w38787 = ~w37666 & w38786;
assign w38788 = w22767 & ~w38787;
assign w38789 = w22767 & ~w37666;
assign w38790 = ~w26445 & ~w38789;
assign w38791 = ~w38786 & w38790;
assign w38792 = w38735 & ~w38791;
assign w38793 = ~w38782 & ~w38788;
assign w38794 = w38792 & ~w38793;
assign w38795 = ~w21801 & w38617;
assign w38796 = w21801 & ~w38618;
assign w38797 = ~w38617 & w38796;
assign w38798 = ~w38795 & ~w38797;
assign w38799 = ~w21801 & ~w38618;
assign w38800 = w20906 & ~w38626;
assign w38801 = ~w38799 & ~w38800;
assign w38802 = ~w21801 & w37673;
assign w38803 = w20906 & w38626;
assign w38804 = w38798 & w38803;
assign w38805 = ~w38720 & w38802;
assign w38806 = ~w38804 & ~w38805;
assign w38807 = ~w38798 & ~w38801;
assign w38808 = w38806 & ~w38807;
assign w38809 = w38702 & ~w38708;
assign w38810 = ~w38670 & w38809;
assign w38811 = ~w38667 & w38808;
assign w38812 = ~w38794 & w38811;
assign w38813 = w38810 & ~w38812;
assign w38814 = (~w38336 & w46333) | (~w38336 & w46334) | (w46333 & w46334);
assign w38815 = ~w38562 & ~w38814;
assign w38816 = w37790 & w38556;
assign w38817 = w38815 & ~w38816;
assign w38818 = ~w14766 & ~w38552;
assign w38819 = w38817 & w38818;
assign w38820 = ~w17380 & ~w37647;
assign w38821 = ~w37648 & ~w38820;
assign w38822 = ~w38688 & w38821;
assign w38823 = ~w38687 & ~w38703;
assign w38824 = w38822 & ~w38823;
assign w38825 = w17380 & ~w37658;
assign w38826 = w38690 & w38825;
assign w38827 = w37658 & ~w38753;
assign w38828 = ~w20421 & ~w37648;
assign w38829 = w38827 & ~w38828;
assign w38830 = w38826 & ~w38687;
assign w38831 = (w37538 & w46335) | (w37538 & w46336) | (w46335 & w46336);
assign w38832 = ~w38830 & ~w38831;
assign w38833 = ~w37658 & ~w38687;
assign w38834 = w19040 & w37647;
assign w38835 = w17380 & ~w38834;
assign w38836 = ~w38690 & w38835;
assign w38837 = ~w38833 & w38836;
assign w38838 = w38832 & ~w38837;
assign w38839 = ~w16559 & w38684;
assign w38840 = ~w38839 & w46337;
assign w38841 = w38686 & ~w38840;
assign w38842 = w23843 & ~w37354;
assign w38843 = w22767 & w37666;
assign w38844 = ~w38842 & ~w38843;
assign w38845 = ~w38802 & ~w38803;
assign w38846 = w38747 & w38845;
assign w38847 = w38744 & ~w38844;
assign w38848 = w38846 & ~w38847;
assign w38849 = w17380 & ~w37647;
assign w38850 = ~w18183 & w37658;
assign w38851 = ~w38849 & ~w38850;
assign w38852 = w38751 & ~w38848;
assign w38853 = w38851 & ~w38852;
assign w38854 = ~w16559 & w37690;
assign w38855 = w38755 & ~w38853;
assign w38856 = ~w38854 & ~w38855;
assign w38857 = ~w38336 & w46338;
assign w38858 = ~w38841 & ~w38857;
assign w38859 = ~w15681 & w38547;
assign w38860 = w38858 & ~w38859;
assign w38861 = ~w38540 & w38860;
assign w38862 = ~w38819 & w38861;
assign w38863 = ~w38813 & w38862;
assign w38864 = w38615 & ~w38863;
assign w38865 = ~w37746 & ~w38591;
assign w38866 = ~w37775 & ~w37776;
assign w38867 = ~w38865 & w38866;
assign w38868 = ~w11870 & ~w37726;
assign w38869 = ~w11138 & w38339;
assign w38870 = (~w38868 & w38336) | (~w38868 & w46339) | (w38336 & w46339);
assign w38871 = ~w38867 & w38870;
assign w38872 = ~w38869 & ~w38871;
assign w38873 = ~w37709 & ~w37777;
assign w38874 = ~w10419 & ~w37836;
assign w38875 = ~w37821 & w46340;
assign w38876 = (~w38875 & w38336) | (~w38875 & w43201) | (w38336 & w43201);
assign w38877 = (w38336 & w46341) | (w38336 & w46342) | (w46341 & w46342);
assign w38878 = w37954 & ~w38877;
assign w38879 = ~w37954 & w38877;
assign w38880 = ~w38878 & ~w38879;
assign w38881 = w9781 & w38880;
assign w38882 = w10419 & w38873;
assign w38883 = w38872 & w38882;
assign w38884 = w10419 & ~w38873;
assign w38885 = ~w38872 & w38884;
assign w38886 = ~w38881 & ~w38885;
assign w38887 = ~w38883 & w38886;
assign w38888 = ~w38584 & w46343;
assign w38889 = (~w13384 & w38610) | (~w13384 & w48080) | (w38610 & w48080);
assign w38890 = ~w38888 & ~w38889;
assign w38891 = ~w38593 & w43202;
assign w38892 = w11870 & ~w38891;
assign w38893 = ~w38590 & ~w38594;
assign w38894 = w38892 & ~w38893;
assign w38895 = ~w38336 & w46344;
assign w38896 = (~w37775 & w38336) | (~w37775 & w43203) | (w38336 & w43203);
assign w38897 = ~w38865 & w38896;
assign w38898 = ~w38895 & ~w38897;
assign w38899 = ~w37776 & ~w38868;
assign w38900 = ~w11138 & w38899;
assign w38901 = (w38900 & w38897) | (w38900 & w46345) | (w38897 & w46345);
assign w38902 = ~w11138 & ~w38899;
assign w38903 = ~w38897 & w46346;
assign w38904 = ~w38901 & ~w38903;
assign w38905 = ~w38894 & w38904;
assign w38906 = w38603 & ~w38890;
assign w38907 = w38905 & ~w38906;
assign w38908 = w38887 & w38907;
assign w38909 = ~w38864 & w38908;
assign w38910 = ~w38780 & w38909;
assign w38911 = ~w38897 & w46347;
assign w38912 = w11138 & ~w38911;
assign w38913 = ~w38898 & w38899;
assign w38914 = w38912 & ~w38913;
assign w38915 = ~w10419 & ~w38873;
assign w38916 = w38872 & w38915;
assign w38917 = ~w10419 & w38873;
assign w38918 = ~w38872 & w38917;
assign w38919 = ~w38916 & ~w38918;
assign w38920 = ~w38914 & w38919;
assign w38921 = w38887 & ~w38920;
assign w38922 = ~w7924 & w37938;
assign w38923 = (w37821 & w46348) | (w37821 & w46349) | (w46348 & w46349);
assign w38924 = w8666 & ~w38923;
assign w38925 = ~w8666 & ~w37975;
assign w38926 = ~w38924 & ~w38925;
assign w38927 = w38922 & ~w38926;
assign w38928 = w4838 & ~w37888;
assign w38929 = ~w5330 & ~w37890;
assign w38930 = ~w38928 & ~w38929;
assign w38931 = ~w7315 & ~w37925;
assign w38932 = w6769 & w37898;
assign w38933 = ~w38931 & ~w38932;
assign w38934 = w6264 & w37877;
assign w38935 = ~w6769 & ~w37898;
assign w38936 = ~w38934 & ~w38935;
assign w38937 = ~w38933 & w38936;
assign w38938 = ~w6264 & ~w37877;
assign w38939 = w5745 & ~w37869;
assign w38940 = ~w38938 & ~w38939;
assign w38941 = ~w38937 & w38940;
assign w38942 = ~w38922 & ~w38925;
assign w38943 = w38930 & w38941;
assign w38944 = w38942 & w38943;
assign w38945 = ~w38336 & w46350;
assign w38946 = ~w38927 & ~w38945;
assign w38947 = ~w8666 & ~w38942;
assign w38948 = w11648 & w37964;
assign w38949 = ~w37982 & ~w38948;
assign w38950 = (~w37954 & w43205) | (~w37954 & w37836) | (w43205 & w37836);
assign w38951 = (w37821 & w46351) | (w37821 & w46352) | (w46351 & w46352);
assign w38952 = ~w38950 & w38951;
assign w38953 = w38949 & ~w38952;
assign w38954 = w9195 & ~w38953;
assign w38955 = ~w9195 & w38949;
assign w38956 = ~w38952 & w38955;
assign w38957 = ~w37939 & ~w38162;
assign w38958 = (~w37987 & w38162) | (~w37987 & w43207) | (w38162 & w43207);
assign w38959 = (w38162 & w37988) | (w38162 & w46353) | (w37988 & w46353);
assign w38960 = (w38959 & w37821) | (w38959 & w46354) | (w37821 & w46354);
assign w38961 = w37990 & ~w38957;
assign w38962 = w37941 & ~w38961;
assign w38963 = ~w37899 & w52296;
assign w38964 = w6769 & w38938;
assign w38965 = w38963 & w38964;
assign w38966 = ~w6769 & w38938;
assign w38967 = ~w38963 & w38966;
assign w38968 = ~w38965 & ~w38967;
assign w38969 = ~w37986 & w38947;
assign w38970 = w38956 & w38969;
assign w38971 = w38968 & ~w38970;
assign w38972 = w38947 & w38954;
assign w38973 = w38971 & ~w38972;
assign w38974 = w37736 & ~w37939;
assign w38975 = ~w37985 & ~w37986;
assign w38976 = w38974 & ~w38975;
assign w38977 = w38958 & ~w38976;
assign w38978 = w37779 & w38958;
assign w38979 = ~w38865 & w38978;
assign w38980 = ~w38977 & ~w38979;
assign w38981 = ~w37899 & ~w37905;
assign w38982 = ~w37926 & ~w38931;
assign w38983 = w38981 & ~w38982;
assign w38984 = w6769 & ~w38983;
assign w38985 = ~w38981 & w38982;
assign w38986 = w38984 & ~w38985;
assign w38987 = ~w37926 & ~w37928;
assign w38988 = ~w7315 & w38987;
assign w38989 = ~w38986 & ~w38988;
assign w38990 = w6769 & ~w38963;
assign w38991 = w38934 & ~w38990;
assign w38992 = (w37836 & w46355) | (w37836 & w46356) | (w46355 & w46356);
assign w38993 = ~w6769 & ~w38992;
assign w38994 = w6841 & ~w37877;
assign w38995 = ~w38963 & w38994;
assign w38996 = ~w38993 & ~w38995;
assign w38997 = ~w7545 & ~w37926;
assign w38998 = ~w37940 & w38997;
assign w38999 = ~w38961 & w38998;
assign w39000 = w7315 & w37877;
assign w39001 = ~w8258 & ~w37901;
assign w39002 = ~w39000 & ~w39001;
assign w39003 = ~w6769 & w38981;
assign w39004 = w6264 & ~w39002;
assign w39005 = ~w39003 & ~w39004;
assign w39006 = ~w38960 & w38999;
assign w39007 = w39005 & ~w39006;
assign w39008 = ~w38991 & w38996;
assign w39009 = ~w39007 & ~w39008;
assign w39010 = ~w37898 & w37928;
assign w39011 = w6769 & ~w39010;
assign w39012 = ~w37928 & w38981;
assign w39013 = w39011 & ~w39012;
assign w39014 = ~w7315 & ~w38987;
assign w39015 = ~w39013 & ~w39014;
assign w39016 = ~w38980 & w39015;
assign w39017 = ~w39009 & ~w39016;
assign w39018 = w38980 & w38989;
assign w39019 = w39017 & ~w39018;
assign w39020 = ~w8666 & w37975;
assign w39021 = w9195 & w39020;
assign w39022 = w38953 & w39021;
assign w39023 = ~w9195 & w39020;
assign w39024 = ~w38953 & w39023;
assign w39025 = ~w39022 & ~w39024;
assign w39026 = ~w37867 & ~w37870;
assign w39027 = w37927 & ~w38959;
assign w39028 = w37902 & ~w39027;
assign w39029 = (w39028 & w37821) | (w39028 & w46357) | (w37821 & w46357);
assign w39030 = w37902 & ~w37991;
assign w39031 = ~w39027 & w39030;
assign w39032 = ~w37878 & ~w39031;
assign w39033 = ~w39029 & w39032;
assign w39034 = (w39026 & w39029) | (w39026 & w43209) | (w39029 & w43209);
assign w39035 = ~w39029 & w43210;
assign w39036 = ~w39034 & ~w39035;
assign w39037 = w7545 & w37877;
assign w39038 = ~w38963 & w39037;
assign w39039 = ~w6264 & w37901;
assign w39040 = w38963 & w39039;
assign w39041 = ~w39038 & ~w39040;
assign w39042 = w5745 & w39036;
assign w39043 = w39041 & ~w39042;
assign w39044 = ~w7924 & ~w37938;
assign w39045 = ~w38924 & w39044;
assign w39046 = ~w8666 & ~w38956;
assign w39047 = w39045 & ~w39046;
assign w39048 = w38946 & w39025;
assign w39049 = w39043 & ~w39047;
assign w39050 = w39048 & w39049;
assign w39051 = w37879 & ~w39030;
assign w39052 = (w39051 & w37836) | (w39051 & w43211) | (w37836 & w43211);
assign w39053 = w37868 & ~w39052;
assign w39054 = ~w37891 & ~w39053;
assign w39055 = w4838 & w37888;
assign w39056 = w37860 & ~w39055;
assign w39057 = ~w37860 & ~w37891;
assign w39058 = ~w37860 & w38928;
assign w39059 = ~w5330 & ~w39058;
assign w39060 = ~w37867 & ~w39057;
assign w39061 = ~w39052 & w39060;
assign w39062 = w39059 & ~w39061;
assign w39063 = w39054 & ~w39056;
assign w39064 = w39062 & ~w39063;
assign w39065 = w5330 & ~w39055;
assign w39066 = ~w39054 & w39065;
assign w39067 = w5330 & ~w38928;
assign w39068 = w39054 & w39067;
assign w39069 = ~w39066 & ~w39068;
assign w39070 = ~w39064 & w39069;
assign w39071 = w38973 & ~w39070;
assign w39072 = w39050 & w39071;
assign w39073 = ~w39019 & w39072;
assign w39074 = w38339 & w38946;
assign w39075 = w38973 & w39074;
assign w39076 = ~w39073 & ~w39075;
assign w39077 = ~w38159 & w38949;
assign w39078 = ~w9781 & w38339;
assign w39079 = w38876 & ~w38950;
assign w39080 = ~w39078 & ~w39079;
assign w39081 = w39077 & ~w39080;
assign w39082 = ~w39077 & w39080;
assign w39083 = ~w39081 & ~w39082;
assign w39084 = ~w9781 & ~w38880;
assign w39085 = w9195 & w39083;
assign w39086 = ~w39084 & ~w39085;
assign w39087 = ~w38921 & ~w39076;
assign w39088 = w39086 & w39087;
assign w39089 = ~w38910 & w39088;
assign w39090 = ~w38115 & ~w38117;
assign w39091 = ~w38073 & ~w39090;
assign w39092 = ~w37821 & w46358;
assign w39093 = ~w38168 & w38174;
assign w39094 = (~w38136 & w39092) | (~w38136 & w43212) | (w39092 & w43212);
assign w39095 = ~w4430 & ~w38134;
assign w39096 = (~w39095 & w39092) | (~w39095 & w43213) | (w39092 & w43213);
assign w39097 = w39094 & w39096;
assign w39098 = ~w38073 & ~w38137;
assign w39099 = w39097 & w39098;
assign w39100 = ~w39091 & ~w39099;
assign w39101 = w3242 & ~w38339;
assign w39102 = (~w3242 & w38336) | (~w3242 & w46359) | (w38336 & w46359);
assign w39103 = ~w39100 & w39101;
assign w39104 = w39100 & w39102;
assign w39105 = ~w39103 & ~w39104;
assign w39106 = (~w38115 & w38336) | (~w38115 & w46360) | (w38336 & w46360);
assign w39107 = ~w38137 & w39097;
assign w39108 = w39106 & ~w39107;
assign w39109 = ~w38073 & ~w38117;
assign w39110 = ~w38336 & w46361;
assign w39111 = (w39109 & w38336) | (w39109 & w46362) | (w38336 & w46362);
assign w39112 = ~w39110 & ~w39111;
assign w39113 = w39108 & w39109;
assign w39114 = ~w39108 & w39112;
assign w39115 = ~w39113 & ~w39114;
assign w39116 = ~w3242 & ~w39115;
assign w39117 = w2896 & w38058;
assign w39118 = w39105 & w39117;
assign w39119 = w2896 & ~w38058;
assign w39120 = ~w39105 & w39119;
assign w39121 = ~w39116 & ~w39120;
assign w39122 = ~w39118 & w39121;
assign w39123 = ~w2896 & ~w38058;
assign w39124 = ~w38059 & w39091;
assign w39125 = ~w38039 & ~w39124;
assign w39126 = ~w38059 & w39098;
assign w39127 = w39097 & w39126;
assign w39128 = w39125 & ~w39127;
assign w39129 = ~w38044 & w38048;
assign w39130 = w2558 & ~w39129;
assign w39131 = w38339 & w39130;
assign w39132 = w2896 & w39130;
assign w39133 = ~w39128 & w39132;
assign w39134 = ~w39131 & ~w39133;
assign w39135 = ~w38050 & ~w38057;
assign w39136 = w2558 & ~w39135;
assign w39137 = ~w38339 & w39136;
assign w39138 = w3278 & w39129;
assign w39139 = w39102 & w39138;
assign w39140 = ~w39100 & w39139;
assign w39141 = w39128 & w39137;
assign w39142 = ~w39140 & ~w39141;
assign w39143 = w39134 & w39142;
assign w39144 = w39105 & w39123;
assign w39145 = w39143 & ~w39144;
assign w39146 = ~w2896 & w38058;
assign w39147 = ~w39105 & w39146;
assign w39148 = w39145 & ~w39147;
assign w39149 = (~w2285 & w38336) | (~w2285 & w43214) | (w38336 & w43214);
assign w39150 = ~w38077 & ~w38137;
assign w39151 = ~w38136 & w39150;
assign w39152 = ~w38078 & w39151;
assign w39153 = (w39152 & w39092) | (w39152 & w43215) | (w39092 & w43215);
assign w39154 = w39096 & w39153;
assign w39155 = ~w38077 & ~w38119;
assign w39156 = ~w38078 & w39155;
assign w39157 = ~w38011 & ~w39156;
assign w39158 = ~w39154 & w39157;
assign w39159 = (w2285 & w38336) | (w2285 & w43216) | (w38336 & w43216);
assign w39160 = w39149 & ~w39158;
assign w39161 = w39158 & w39159;
assign w39162 = ~w39160 & ~w39161;
assign w39163 = w1738 & w37272;
assign w39164 = ~w39162 & ~w39163;
assign w39165 = w38083 & ~w38084;
assign w39166 = ~w38083 & w38084;
assign w39167 = ~w39165 & ~w39166;
assign w39168 = w2285 & ~w39167;
assign w39169 = ~w2006 & ~w39168;
assign w39170 = ~w38142 & w43217;
assign w39171 = ~w38339 & ~w39170;
assign w39172 = ~w38339 & w43218;
assign w39173 = w2798 & ~w39158;
assign w39174 = w39172 & ~w39173;
assign w39175 = ~w38142 & w43219;
assign w39176 = (w2006 & w38142) | (w2006 & w46363) | (w38142 & w46363);
assign w39177 = ~w38339 & w46364;
assign w39178 = (~w37272 & ~w39171) | (~w37272 & w43220) | (~w39171 & w43220);
assign w39179 = w39167 & w39177;
assign w39180 = ~w39162 & w39179;
assign w39181 = (w39171 & w39163) | (w39171 & w46365) | (w39163 & w46365);
assign w39182 = ~w39174 & w39181;
assign w39183 = ~w39180 & ~w39182;
assign w39184 = w2006 & ~w39167;
assign w39185 = ~w39164 & w39184;
assign w39186 = w39183 & ~w39185;
assign w39187 = (w39151 & w39092) | (w39151 & w43221) | (w39092 & w43221);
assign w39188 = w39096 & w39187;
assign w39189 = ~w39155 & ~w39188;
assign w39190 = (~w2558 & w38336) | (~w2558 & w46366) | (w38336 & w46366);
assign w39191 = w39189 & w39190;
assign w39192 = (w2558 & w38336) | (w2558 & w46367) | (w38336 & w46367);
assign w39193 = ~w39189 & w39192;
assign w39194 = ~w39191 & ~w39193;
assign w39195 = ~w2558 & w39129;
assign w39196 = ~w38010 & ~w39195;
assign w39197 = w2285 & ~w39196;
assign w39198 = w38010 & w39194;
assign w39199 = w39197 & ~w39198;
assign w39200 = ~w3277 & ~w38057;
assign w39201 = ~w39128 & ~w39200;
assign w39202 = ~w2558 & w38057;
assign w39203 = w39189 & ~w39202;
assign w39204 = ~w38339 & ~w39203;
assign w39205 = ~w39201 & w39204;
assign w39206 = w2285 & ~w38010;
assign w39207 = ~w39195 & ~w39206;
assign w39208 = ~w39191 & w39207;
assign w39209 = ~w39205 & ~w39208;
assign w39210 = ~w39199 & ~w39209;
assign w39211 = w39186 & w39210;
assign w39212 = ~w39122 & w39148;
assign w39213 = w39211 & ~w39212;
assign w39214 = ~w38339 & ~w38956;
assign w39215 = ~w38954 & w39214;
assign w39216 = w37975 & w39215;
assign w39217 = w8666 & ~w39216;
assign w39218 = ~w37975 & ~w39215;
assign w39219 = w39217 & ~w39218;
assign w39220 = ~w9195 & ~w39083;
assign w39221 = ~w39219 & ~w39220;
assign w39222 = ~w37939 & ~w37987;
assign w39223 = w37925 & ~w37987;
assign w39224 = ~w37925 & w37987;
assign w39225 = ~w39223 & ~w39224;
assign w39226 = w7924 & ~w39225;
assign w39227 = w7315 & ~w39226;
assign w39228 = w7315 & ~w39225;
assign w39229 = ~w7924 & ~w39228;
assign w39230 = ~w38923 & w39222;
assign w39231 = ~w39222 & ~w39227;
assign w39232 = w38923 & w39231;
assign w39233 = ~w39230 & ~w39232;
assign w39234 = ~w39229 & w39233;
assign w39235 = w7315 & ~w37939;
assign w39236 = ~w38987 & w39235;
assign w39237 = ~w38923 & w39236;
assign w39238 = ~w3646 & w38114;
assign w39239 = ~w38121 & ~w39238;
assign w39240 = w38339 & w39239;
assign w39241 = w7315 & w37925;
assign w39242 = w7924 & ~w37938;
assign w39243 = ~w39241 & ~w39242;
assign w39244 = w38936 & w39243;
assign w39245 = w38941 & ~w39244;
assign w39246 = ~w5745 & w37869;
assign w39247 = w5330 & w37890;
assign w39248 = ~w39246 & ~w39247;
assign w39249 = ~w39245 & w39248;
assign w39250 = w38930 & ~w39249;
assign w39251 = ~w4838 & w37888;
assign w39252 = ~w39250 & ~w39251;
assign w39253 = w39240 & w39252;
assign w39254 = ~w39070 & ~w39253;
assign w39255 = w38968 & w39043;
assign w39256 = w39254 & w39255;
assign w39257 = ~w39234 & ~w39237;
assign w39258 = ~w39009 & w39257;
assign w39259 = w39256 & ~w39258;
assign w39260 = w4056 & ~w39097;
assign w39261 = ~w4056 & w39097;
assign w39262 = ~w39260 & ~w39261;
assign w39263 = w4056 & ~w39094;
assign w39264 = w39096 & w39263;
assign w39265 = ~w38339 & ~w39264;
assign w39266 = ~w3646 & ~w38114;
assign w39267 = ~w39262 & w39266;
assign w39268 = w39265 & ~w39267;
assign w39269 = ~w37889 & ~w38169;
assign w39270 = w37975 & w38164;
assign w39271 = ~w37991 & ~w39270;
assign w39272 = ~w38960 & ~w39271;
assign w39273 = w37904 & ~w39272;
assign w39274 = ~w37880 & ~w37891;
assign w39275 = ~w39273 & w39274;
assign w39276 = ~w39269 & ~w39275;
assign w39277 = ~w4838 & ~w39276;
assign w39278 = w39269 & w39275;
assign w39279 = w39277 & ~w39278;
assign w39280 = w39268 & ~w39279;
assign w39281 = ~w6264 & w38939;
assign w39282 = (~w37867 & w39029) | (~w37867 & w43222) | (w39029 & w43222);
assign w39283 = ~w39281 & ~w39282;
assign w39284 = w39057 & w39283;
assign w39285 = w5330 & ~w39284;
assign w39286 = ~w39057 & ~w39283;
assign w39287 = w39285 & ~w39286;
assign w39288 = ~w39026 & ~w39033;
assign w39289 = ~w5745 & ~w39288;
assign w39290 = ~w37867 & w39052;
assign w39291 = w39289 & ~w39290;
assign w39292 = ~w39287 & ~w39291;
assign w39293 = ~w39092 & w39093;
assign w39294 = w38135 & ~w39293;
assign w39295 = w39096 & ~w39294;
assign w39296 = w39238 & ~w39263;
assign w39297 = w38121 & ~w39295;
assign w39298 = ~w39296 & ~w39297;
assign w39299 = ~w39261 & ~w39298;
assign w39300 = w38134 & ~w38173;
assign w39301 = ~w38168 & ~w38169;
assign w39302 = ~w39092 & w39301;
assign w39303 = (w39302 & w38336) | (w39302 & w46368) | (w38336 & w46368);
assign w39304 = ~w39303 & w43224;
assign w39305 = (~w39300 & w39303) | (~w39300 & w43225) | (w39303 & w43225);
assign w39306 = ~w39304 & ~w39305;
assign w39307 = w4430 & w39306;
assign w39308 = ~w39299 & ~w39307;
assign w39309 = w39254 & ~w39292;
assign w39310 = w39308 & ~w39309;
assign w39311 = ~w39253 & ~w39280;
assign w39312 = w39310 & ~w39311;
assign w39313 = ~w39019 & w39259;
assign w39314 = w39312 & ~w39313;
assign w39315 = ~w39076 & ~w39221;
assign w39316 = w39314 & ~w39315;
assign w39317 = w39213 & w39316;
assign w39318 = ~w39089 & w39317;
assign w39319 = ~w38339 & w39295;
assign w39320 = w38120 & ~w39319;
assign w39321 = ~w4056 & ~w39320;
assign w39322 = ~w38120 & w39319;
assign w39323 = w39321 & ~w39322;
assign w39324 = ~w4430 & ~w39306;
assign w39325 = ~w39323 & ~w39324;
assign w39326 = w39268 & ~w39299;
assign w39327 = ~w39240 & ~w39326;
assign w39328 = ~w39325 & ~w39327;
assign w39329 = ~w39123 & ~w39130;
assign w39330 = w38339 & w39329;
assign w39331 = ~w39262 & ~w39330;
assign w39332 = ~w38114 & ~w38339;
assign w39333 = ~w39262 & w39332;
assign w39334 = w3646 & ~w39333;
assign w39335 = w38114 & ~w39331;
assign w39336 = w39334 & ~w39335;
assign w39337 = w3242 & w39115;
assign w39338 = ~w39336 & ~w39337;
assign w39339 = w39148 & ~w39328;
assign w39340 = w39338 & w39339;
assign w39341 = w39213 & ~w39340;
assign w39342 = w252 & w38309;
assign w39343 = w38270 & ~w39342;
assign w39344 = (~w38254 & w38197) | (~w38254 & w46369) | (w38197 & w46369);
assign w39345 = ~w39343 & w39344;
assign w39346 = w39343 & ~w39344;
assign w39347 = ~w38309 & w38339;
assign w39348 = ~w39345 & ~w39346;
assign w39349 = ~w38339 & w39348;
assign w39350 = ~w39347 & ~w39349;
assign w39351 = ~w39342 & w52297;
assign w39352 = ~w38290 & ~w38305;
assign w39353 = ~w39351 & w39352;
assign w39354 = w39351 & ~w39352;
assign w39355 = w38289 & w38339;
assign w39356 = ~w39353 & ~w39354;
assign w39357 = ~w38339 & w39356;
assign w39358 = ~w39355 & ~w39357;
assign w39359 = ~w57 & ~w39350;
assign w39360 = w80 & w39358;
assign w39361 = ~w39359 & ~w39360;
assign w39362 = w37193 & ~w37287;
assign w39363 = w37298 & ~w39362;
assign w39364 = (w39363 & w38142) | (w39363 & w43227) | (w38142 & w43227);
assign w39365 = (~w37300 & w39364) | (~w37300 & w46370) | (w39364 & w46370);
assign w39366 = ~w37312 & ~w38254;
assign w39367 = ~w39365 & w39366;
assign w39368 = w39365 & ~w39366;
assign w39369 = ~w37311 & w38339;
assign w39370 = ~w39367 & ~w39368;
assign w39371 = ~w38339 & w39370;
assign w39372 = ~w39369 & ~w39371;
assign w39373 = w57 & w39350;
assign w39374 = w252 & ~w39372;
assign w39375 = ~w39373 & ~w39374;
assign w39376 = w38318 & w38321;
assign w39377 = w39376 & w52298;
assign w39378 = ~w38210 & ~w39377;
assign w39379 = ~w38222 & w39378;
assign w39380 = ~w38221 & w38248;
assign w39381 = w37107 & ~w38236;
assign w39382 = w39380 & ~w39381;
assign w39383 = ~w39379 & w39382;
assign w39384 = ~w1 & w38220;
assign w39385 = w39383 & ~w39384;
assign w39386 = ~w38222 & ~w38248;
assign w39387 = ~w39380 & ~w39386;
assign w39388 = ~w39378 & w39387;
assign w39389 = w42 & ~w39388;
assign w39390 = w39379 & w39380;
assign w39391 = w39389 & ~w39390;
assign w39392 = ~w42 & ~w38249;
assign w39393 = w38221 & ~w38248;
assign w39394 = w39392 & ~w39393;
assign w39395 = w39378 & w39386;
assign w39396 = w39394 & ~w39395;
assign w39397 = ~w39385 & w39391;
assign w39398 = ~w39383 & w39396;
assign w39399 = ~w39397 & ~w39398;
assign w39400 = ~w38305 & ~w38339;
assign w39401 = ~w39353 & w39400;
assign w39402 = w80 & w38339;
assign w39403 = ~w39401 & ~w39402;
assign w39404 = w3 & ~w38209;
assign w39405 = ~w39403 & w39404;
assign w39406 = w3 & w38209;
assign w39407 = w39403 & w39406;
assign w39408 = ~w39405 & ~w39407;
assign w39409 = ~w80 & ~w39358;
assign w39410 = w39408 & ~w39409;
assign w39411 = w39399 & w39410;
assign w39412 = w39361 & ~w39375;
assign w39413 = w39411 & ~w39412;
assign w39414 = (w38189 & w38176) | (w38189 & w43229) | (w38176 & w43229);
assign w39415 = (w37286 & w38142) | (w37286 & w43230) | (w38142 & w43230);
assign w39416 = (~w37205 & w39415) | (~w37205 & w46371) | (w39415 & w46371);
assign w39417 = ~w1120 & w39416;
assign w39418 = w1120 & ~w39416;
assign w39419 = ~w39417 & ~w39418;
assign w39420 = ~w38339 & w39419;
assign w39421 = ~w38142 & w43231;
assign w39422 = w37288 & w39421;
assign w39423 = ~w37287 & w37288;
assign w39424 = w754 & ~w39423;
assign w39425 = (w39424 & ~w39421) | (w39424 & w46372) | (~w39421 & w46372);
assign w39426 = w612 & ~w37149;
assign w39427 = (~w39426 & w38336) | (~w39426 & w46373) | (w38336 & w46373);
assign w39428 = ~w39425 & w39427;
assign w39429 = ~w38192 & w46374;
assign w39430 = ~w37288 & ~w39429;
assign w39431 = w37287 & ~w37288;
assign w39432 = ~w39430 & w52299;
assign w39433 = w37192 & w37287;
assign w39434 = ~w39421 & w39433;
assign w39435 = ~w39432 & ~w39434;
assign w39436 = (w754 & w38336) | (w754 & w46375) | (w38336 & w46375);
assign w39437 = w39435 & w39436;
assign w39438 = ~w39428 & ~w39437;
assign w39439 = ~w754 & ~w37191;
assign w39440 = ~w754 & w39432;
assign w39441 = ~w38339 & w39440;
assign w39442 = ~w39439 & ~w39441;
assign w39443 = w39438 & w39442;
assign w39444 = w37222 & ~w39420;
assign w39445 = ~w37222 & w39419;
assign w39446 = ~w39443 & w39445;
assign w39447 = ~w39444 & ~w39446;
assign w39448 = w612 & w37149;
assign w39449 = w39428 & ~w39440;
assign w39450 = w39448 & ~w39449;
assign w39451 = w754 & w37191;
assign w39452 = ~w38339 & ~w39440;
assign w39453 = ~w39451 & ~w39452;
assign w39454 = w39438 & ~w39453;
assign w39455 = (w37287 & w38142) | (w37287 & w43233) | (w38142 & w43233);
assign w39456 = w39429 & ~w39455;
assign w39457 = w37290 & ~w39456;
assign w39458 = ~w37150 & ~w39457;
assign w39459 = w612 & ~w39458;
assign w39460 = ~w493 & w37294;
assign w39461 = w39459 & ~w39460;
assign w39462 = ~w612 & ~w37150;
assign w39463 = w37289 & ~w39460;
assign w39464 = w39462 & ~w39463;
assign w39465 = ~w612 & ~w37149;
assign w39466 = ~w39460 & ~w39465;
assign w39467 = ~w493 & w39466;
assign w39468 = ~w39464 & ~w39467;
assign w39469 = ~w612 & w39432;
assign w39470 = w39468 & ~w39469;
assign w39471 = w39439 & ~w39448;
assign w39472 = w39466 & ~w39471;
assign w39473 = w38339 & w39472;
assign w39474 = ~w39460 & w39464;
assign w39475 = w39432 & w39474;
assign w39476 = ~w39473 & ~w39475;
assign w39477 = ~w39459 & w39470;
assign w39478 = w39476 & ~w39477;
assign w39479 = ~w39422 & ~w39423;
assign w39480 = ~w39448 & ~w39479;
assign w39481 = ~w39426 & w39435;
assign w39482 = ~w38339 & ~w39481;
assign w39483 = ~w39436 & ~w39473;
assign w39484 = ~w39480 & w39482;
assign w39485 = w39483 & ~w39484;
assign w39486 = ~w39461 & w39478;
assign w39487 = ~w39485 & ~w39486;
assign w39488 = ~w39454 & w46376;
assign w39489 = ~w39447 & w39488;
assign w39490 = w39487 & ~w39489;
assign w39491 = (w38336 & w39168) | (w38336 & w46377) | (w39168 & w46377);
assign w39492 = w39167 & ~w39159;
assign w39493 = ~w39491 & ~w39492;
assign w39494 = (w38336 & w46378) | (w38336 & w46379) | (w46378 & w46379);
assign w39495 = (~w38336 & w46380) | (~w38336 & w46381) | (w46380 & w46381);
assign w39496 = ~w39494 & ~w39495;
assign w39497 = ~w2006 & w39158;
assign w39498 = ~w39493 & w39497;
assign w39499 = ~w2006 & ~w39158;
assign w39500 = ~w39496 & w39499;
assign w39501 = ~w39498 & ~w39500;
assign w39502 = ~w2285 & ~w38010;
assign w39503 = ~w39194 & w39502;
assign w39504 = w39501 & ~w39503;
assign w39505 = ~w2285 & w38010;
assign w39506 = w39194 & w39505;
assign w39507 = w39504 & ~w39506;
assign w39508 = w37239 & w37285;
assign w39509 = (w37279 & w38142) | (w37279 & w43235) | (w38142 & w43235);
assign w39510 = ~w38339 & w39509;
assign w39511 = ~w39510 & w43236;
assign w39512 = (~w39508 & w39510) | (~w39508 & w43237) | (w39510 & w43237);
assign w39513 = ~w39511 & ~w39512;
assign w39514 = ~w37205 & w37246;
assign w39515 = ~w38336 & w46382;
assign w39516 = ~w38339 & w43238;
assign w39517 = (w39514 & w39516) | (w39514 & w46383) | (w39516 & w46383);
assign w39518 = ~w39516 & w46384;
assign w39519 = ~w39517 & ~w39518;
assign w39520 = ~w1320 & w39513;
assign w39521 = w1120 & w39519;
assign w39522 = ~w39520 & ~w39521;
assign w39523 = w37165 & w39429;
assign w39524 = w37298 & ~w39523;
assign w39525 = ~w37123 & ~w39524;
assign w39526 = (w400 & w39364) | (w400 & w46385) | (w39364 & w46385);
assign w39527 = ~w37291 & ~w37296;
assign w39528 = (w39527 & w39455) | (w39527 & w46386) | (w39455 & w46386);
assign w39529 = w400 & ~w37122;
assign w39530 = ~w493 & w39529;
assign w39531 = ~w39528 & w39530;
assign w39532 = ~w39526 & ~w39531;
assign w39533 = w37122 & w38339;
assign w39534 = w37123 & w39528;
assign w39535 = ~w39533 & ~w39534;
assign w39536 = ~w400 & w39525;
assign w39537 = ~w39364 & w39536;
assign w39538 = ~w39526 & ~w39537;
assign w39539 = ~w351 & w37137;
assign w39540 = ~w38339 & w39539;
assign w39541 = ~w39538 & w39540;
assign w39542 = ~w351 & ~w37137;
assign w39543 = ~w39529 & ~w39542;
assign w39544 = w38339 & ~w39543;
assign w39545 = w400 & w37122;
assign w39546 = w39527 & w39545;
assign w39547 = (w39546 & w39455) | (w39546 & w46387) | (w39455 & w46387);
assign w39548 = (w39542 & w39364) | (w39542 & w48081) | (w39364 & w48081);
assign w39549 = ~w39547 & w39548;
assign w39550 = ~w39544 & ~w39549;
assign w39551 = ~w39541 & w39550;
assign w39552 = ~w39532 & w39535;
assign w39553 = w39551 & ~w39552;
assign w39554 = ~w38336 & w43239;
assign w39555 = ~w38339 & ~w39176;
assign w39556 = ~w39554 & ~w39555;
assign w39557 = w37254 & ~w37276;
assign w39558 = ~w1541 & ~w39557;
assign w39559 = (~w39558 & w38339) | (~w39558 & w46388) | (w38339 & w46388);
assign w39560 = ~w1541 & w39557;
assign w39561 = ~w38339 & w46389;
assign w39562 = (~w39560 & w38336) | (~w39560 & w46390) | (w38336 & w46390);
assign w39563 = ~w39555 & w39562;
assign w39564 = ~w39561 & ~w39563;
assign w39565 = ~w39556 & w39559;
assign w39566 = w39564 & ~w39565;
assign w39567 = ~w38339 & w46391;
assign w39568 = (~w1738 & w39178) | (~w1738 & w46392) | (w39178 & w46392);
assign w39569 = ~w39566 & ~w39568;
assign w39570 = w39553 & w39569;
assign w39571 = w39522 & w39570;
assign w39572 = w39186 & ~w39507;
assign w39573 = w39571 & ~w39572;
assign w39574 = w39490 & w39573;
assign w39575 = w39413 & w39574;
assign w39576 = ~w39341 & w39575;
assign w39577 = ~w39172 & ~w39556;
assign w39578 = w1320 & ~w39513;
assign w39579 = w1541 & w39557;
assign w39580 = w39577 & w39579;
assign w39581 = w1541 & ~w39557;
assign w39582 = (w39581 & w39556) | (w39581 & w43240) | (w39556 & w43240);
assign w39583 = ~w39578 & ~w39582;
assign w39584 = ~w39580 & w39583;
assign w39585 = w39522 & ~w39584;
assign w39586 = ~w945 & w37222;
assign w39587 = w39419 & w43241;
assign w39588 = ~w39454 & w46393;
assign w39589 = ~w945 & ~w37222;
assign w39590 = (w39589 & ~w39419) | (w39589 & w43242) | (~w39419 & w43242);
assign w39591 = ~w1120 & ~w39519;
assign w39592 = ~w39590 & ~w39591;
assign w39593 = w39588 & w39592;
assign w39594 = ~w39585 & w39593;
assign w39595 = w39490 & ~w39594;
assign w39596 = (~w38339 & w39458) | (~w38339 & w43243) | (w39458 & w43243);
assign w39597 = ~w612 & w39458;
assign w39598 = w39596 & ~w39597;
assign w39599 = ~w37294 & w39598;
assign w39600 = w493 & ~w39599;
assign w39601 = w37294 & ~w39598;
assign w39602 = w39600 & ~w39601;
assign w39603 = ~w493 & ~w39528;
assign w39604 = ~w38339 & ~w39603;
assign w39605 = w493 & w39528;
assign w39606 = w39604 & ~w39605;
assign w39607 = ~w37122 & ~w39606;
assign w39608 = ~w400 & ~w39607;
assign w39609 = w37122 & w39606;
assign w39610 = w39608 & ~w39609;
assign w39611 = ~w39602 & ~w39610;
assign w39612 = ~w39595 & w39611;
assign w39613 = ~w38209 & ~w39403;
assign w39614 = ~w3 & ~w39613;
assign w39615 = w38209 & w39403;
assign w39616 = w39614 & ~w39615;
assign w39617 = ~w38221 & ~w38222;
assign w39618 = w39378 & ~w39617;
assign w39619 = w39392 & ~w39618;
assign w39620 = ~w39378 & w39617;
assign w39621 = w39619 & ~w39620;
assign w39622 = ~w38220 & w38237;
assign w39623 = ~w39621 & ~w39622;
assign w39624 = ~w39616 & w39623;
assign w39625 = ~w38339 & ~w39538;
assign w39626 = w37137 & w39625;
assign w39627 = w351 & ~w39626;
assign w39628 = ~w37137 & ~w39625;
assign w39629 = w39627 & ~w39628;
assign w39630 = ~w252 & w39372;
assign w39631 = ~w39629 & ~w39630;
assign w39632 = w39361 & w39631;
assign w39633 = w39413 & ~w39632;
assign w39634 = w39399 & ~w39624;
assign w39635 = ~w39633 & ~w39634;
assign w39636 = w39413 & w39553;
assign w39637 = ~w39612 & w39636;
assign w39638 = w39635 & ~w39637;
assign w39639 = ~w39318 & w39576;
assign w39640 = w39638 & ~w39639;
assign w39641 = w5 & ~w9;
assign w39642 = a[126] & ~w1;
assign w39643 = w45 & a[122];
assign w39644 = a[120] & a[121];
assign w39645 = w83 & ~w85;
assign w39646 = ~w83 & ~w81;
assign w39647 = ~w100 & w50670;
assign w39648 = ~w55 & ~w107;
assign w39649 = (~w3 & w102) | (~w3 & w50671) | (w102 & w50671);
assign w39650 = w11 & a[123];
assign w39651 = a[122] & ~w1;
assign w39652 = a[122] & a[123];
assign w39653 = w24 & ~w35;
assign w39654 = w36 & w47;
assign w39655 = w36 & ~a[124];
assign w39656 = w157 & w159;
assign w39657 = w172 & a[122];
assign w39658 = w186 & w43244;
assign w39659 = ~w86 & ~w3;
assign w39660 = w90 & ~w3;
assign w39661 = w157 & ~w205;
assign w39662 = ~w223 & ~w224;
assign w39663 = ~w236 & a[119];
assign w39664 = ~w214 & w43245;
assign w39665 = (~w80 & w214) | (~w80 & w43246) | (w214 & w43246);
assign w39666 = ~w160 & ~w229;
assign w39667 = ~w251 & w259;
assign w39668 = ~w270 & ~w3;
assign w39669 = ~w199 & w3;
assign w39670 = ~w281 & ~w280;
assign w39671 = ~w293 & ~w292;
assign w39672 = ~w228 & ~w268;
assign w39673 = ~w312 & ~w313;
assign w39674 = w234 & w354;
assign w39675 = ~w234 & w358;
assign w39676 = w234 & w367;
assign w39677 = ~w368 & ~w80;
assign w39678 = w303 & ~w213;
assign w39679 = w290 & w219;
assign w39680 = (w43247 & w374) | (w43247 & w50672) | (w374 & w50672);
assign w39681 = (~a[119] & w43248) | (~a[119] & w52300) | (w43248 & w52300);
assign w39682 = w234 & w389;
assign w39683 = ~w234 & w391;
assign w39684 = w368 & w80;
assign w39685 = ~w332 & ~w330;
assign w39686 = (~w39685 & w50673) | (~w39685 & w50674) | (w50673 & w50674);
assign w39687 = ~w330 & w52301;
assign w39688 = ~w330 & w52302;
assign w39689 = ~w330 & w52303;
assign w39690 = (w39685 & w50678) | (w39685 & w50679) | (w50678 & w50679);
assign w39691 = (~w39685 & w50680) | (~w39685 & w50681) | (w50680 & w50681);
assign w39692 = ~w369 & ~w331;
assign w39693 = ~w467 & ~w274;
assign w39694 = (w273 & w370) | (w273 & w50682) | (w370 & w50682);
assign w39695 = (~w3 & w370) | (~w3 & w43249) | (w370 & w43249);
assign w39696 = ~w370 & w43250;
assign w39697 = w459 & w494;
assign w39698 = ~w511 & ~w510;
assign w39699 = ~w515 & w516;
assign w39700 = w515 & w518;
assign w39701 = w459 & ~w456;
assign w39702 = ~w526 & ~w527;
assign w39703 = w492 & w524;
assign w39704 = ~w515 & w537;
assign w39705 = w515 & w539;
assign w39706 = ~w441 & w506;
assign w39707 = (w419 & ~w548) | (w419 & w46394) | (~w548 & w46394);
assign w39708 = w548 & w46395;
assign w39709 = w515 & w553;
assign w39710 = ~w515 & w555;
assign w39711 = ~w492 & w570;
assign w39712 = w492 & w572;
assign w39713 = w492 & ~w577;
assign w39714 = ~w492 & w580;
assign w39715 = ~w492 & w584;
assign w39716 = w492 & w586;
assign w39717 = ~w492 & w597;
assign w39718 = w492 & w599;
assign w39719 = ~w492 & w595;
assign w39720 = w492 & w596;
assign w39721 = w613 & w619;
assign w39722 = w624 & w351;
assign w39723 = ~w628 & w630;
assign w39724 = w628 & w632;
assign w39725 = w588 & ~w252;
assign w39726 = ~w588 & w252;
assign w39727 = ~w628 & w644;
assign w39728 = w628 & w646;
assign w39729 = ~w660 & ~w661;
assign w39730 = ~w652 & w678;
assign w39731 = ~w624 & ~w351;
assign w39732 = w613 & w682;
assign w39733 = (~w57 & ~w606) | (~w57 & w50739) | (~w606 & w50739);
assign w39734 = w606 & w50740;
assign w39735 = w693 & ~w551;
assign w39736 = ~w693 & w50741;
assign w39737 = (w700 & w542) | (w700 & w50780) | (w542 & w50780);
assign w39738 = w543 & w545;
assign w39739 = w512 & w80;
assign w39740 = ~w552 & w50742;
assign w39741 = ~w512 & w727;
assign w39742 = ~w651 & w733;
assign w39743 = w716 & ~w711;
assign w39744 = w738 & ~w703;
assign w39745 = ~w711 & w52304;
assign w39746 = w551 & ~w693;
assign w39747 = (~w750 & ~w746) | (~w750 & w50744) | (~w746 & w50744);
assign w39748 = ~w651 & w760;
assign w39749 = ~w740 & w751;
assign w39750 = ~w773 & w720;
assign w39751 = ~w751 & ~w798;
assign w39752 = w672 & ~w627;
assign w39753 = (w748 & w50745) | (w748 & w50746) | (w50745 & w50746);
assign w39754 = w771 & ~w807;
assign w39755 = (~w869 & w753) | (~w869 & w43252) | (w753 & w43252);
assign w39756 = ~w885 & ~w886;
assign w39757 = w884 & w493;
assign w39758 = (w895 & ~w746) | (w895 & w50747) | (~w746 & w50747);
assign w39759 = ~w933 & ~w932;
assign w39760 = w878 & ~w931;
assign w39761 = w942 & w3;
assign w39762 = ~w877 & w43253;
assign w39763 = (~w351 & w877) | (~w351 & w43254) | (w877 & w43254);
assign w39764 = w1037 & ~w400;
assign w39765 = ~w856 & w252;
assign w39766 = ~w942 & ~w847;
assign w39767 = w1079 & w847;
assign w39768 = ~w1079 & w1083;
assign w39769 = w935 & w1092;
assign w39770 = ~w935 & ~w1092;
assign w39771 = w1079 & w1104;
assign w39772 = w1087 & ~w1097;
assign w39773 = (~w3 & ~w945) | (~w3 & w43255) | (~w945 & w43255);
assign w39774 = ~w1114 & ~w1117;
assign w39775 = ~w1112 & w1118;
assign w39776 = ~w1119 & w46396;
assign w39777 = w1078 & w1102;
assign w39778 = w1143 & ~w1140;
assign w39779 = ~w1143 & w1140;
assign w39780 = w1118 & ~w1157;
assign w39781 = ~w1119 & w46397;
assign w39782 = (w1164 & w1119) | (w1164 & w46398) | (w1119 & w46398);
assign w39783 = ~w1112 & w1169;
assign w39784 = w1170 & ~w1176;
assign w39785 = ~w1112 & ~w1117;
assign w39786 = ~w1114 & ~w978;
assign w39787 = w1118 & w1230;
assign w39788 = w1118 & ~w1245;
assign w39789 = w1118 & ~w1263;
assign w39790 = w1118 & w1268;
assign w39791 = w1118 & w1280;
assign w39792 = w1281 & w1284;
assign w39793 = ~w1281 & ~w1284;
assign w39794 = ~w1158 & w1022;
assign w39795 = w1118 & w1296;
assign w39796 = (~w1161 & w1119) | (~w1161 & w46399) | (w1119 & w46399);
assign w39797 = ~w1119 & w46400;
assign w39798 = (w400 & w1119) | (w400 & w48082) | (w1119 & w48082);
assign w39799 = (~w1314 & w1306) | (~w1314 & w43256) | (w1306 & w43256);
assign w39800 = ~w1307 & w1316;
assign w39801 = (~w1329 & w1215) | (~w1329 & w43257) | (w1215 & w43257);
assign w39802 = ~w1215 & w43258;
assign w39803 = (w1347 & w1215) | (w1347 & w43259) | (w1215 & w43259);
assign w39804 = (w1359 & w1215) | (w1359 & w43260) | (w1215 & w43260);
assign w39805 = ~w1215 & w43261;
assign w39806 = ~w1215 & w43262;
assign w39807 = (w1366 & w1215) | (w1366 & w43263) | (w1215 & w43263);
assign w39808 = ~w1215 & w43264;
assign w39809 = (w1374 & w1215) | (w1374 & w43265) | (w1215 & w43265);
assign w39810 = (w1384 & w1215) | (w1384 & w43266) | (w1215 & w43266);
assign w39811 = ~w1215 & w43267;
assign w39812 = (w493 & ~w1275) | (w493 & w43268) | (~w1275 & w43268);
assign w39813 = w1400 & ~w1401;
assign w39814 = (~w1407 & w1403) | (~w1407 & w43269) | (w1403 & w43269);
assign w39815 = ~w1317 & w1410;
assign w39816 = ~w1398 & w43270;
assign w39817 = (w1421 & w1398) | (w1421 & w43271) | (w1398 & w43271);
assign w39818 = ~w1398 & w43272;
assign w39819 = (~w1287 & w1398) | (~w1287 & w43273) | (w1398 & w43273);
assign w39820 = ~w1457 & ~w1458;
assign w39821 = (~w1466 & w1215) | (~w1466 & w43274) | (w1215 & w43274);
assign w39822 = (w1466 & w1215) | (w1466 & w43275) | (w1215 & w43275);
assign w39823 = (~w1202 & w1215) | (~w1202 & w46401) | (w1215 & w46401);
assign w39824 = ~w1215 & w46402;
assign w39825 = (w1319 & w46403) | (w1319 & w46404) | (w46403 & w46404);
assign w39826 = ~w1499 & w52305;
assign w39827 = w1476 & ~w1513;
assign w39828 = w1530 & ~w80;
assign w39829 = ~w1544 & w1545;
assign w39830 = w1544 & w1547;
assign w39831 = (w1554 & ~w1483) | (w1554 & w51385) | (~w1483 & w51385);
assign w39832 = (~w1555 & ~w1483) | (~w1555 & w51386) | (~w1483 & w51386);
assign w39833 = (w1477 & w46405) | (w1477 & w46406) | (w46405 & w46406);
assign w39834 = (~w1477 & w46407) | (~w1477 & w46408) | (w46407 & w46408);
assign w39835 = ~w1477 & w43276;
assign w39836 = (w1567 & w1477) | (w1567 & w43277) | (w1477 & w43277);
assign w39837 = w1120 & w52306;
assign w39838 = ~w1509 & w1584;
assign w39839 = w1509 & w1586;
assign w39840 = (w1590 & ~w1483) | (w1590 & w51387) | (~w1483 & w51387);
assign w39841 = ~w1570 & ~w1594;
assign w39842 = ~w1477 & w43278;
assign w39843 = (w1583 & w1477) | (w1583 & w43279) | (w1477 & w43279);
assign w39844 = (w1602 & ~w1483) | (w1602 & w51388) | (~w1483 & w51388);
assign w39845 = (~w1477 & w46411) | (~w1477 & w46412) | (w46411 & w46412);
assign w39846 = (w1477 & w46413) | (w1477 & w46414) | (w46413 & w46414);
assign w39847 = (~w1477 & w46415) | (~w1477 & w46416) | (w46415 & w46416);
assign w39848 = (w1477 & w46417) | (w1477 & w46418) | (w46417 & w46418);
assign w39849 = ~w1477 & w43280;
assign w39850 = (w1619 & w1477) | (w1619 & w43281) | (w1477 & w43281);
assign w39851 = ~w1477 & w43282;
assign w39852 = (w1616 & w1477) | (w1616 & w43283) | (w1477 & w43283);
assign w39853 = (~w1477 & w46419) | (~w1477 & w46420) | (w46419 & w46420);
assign w39854 = (w1477 & w46421) | (w1477 & w46422) | (w46421 & w46422);
assign w39855 = ~w1508 & w1652;
assign w39856 = ~w1653 & w1655;
assign w39857 = w1653 & w1657;
assign w39858 = w1509 & w1665;
assign w39859 = ~w1653 & w1692;
assign w39860 = w1653 & w1694;
assign w39861 = ~w1544 & w1700;
assign w39862 = w1544 & w1702;
assign w39863 = ~w1476 & w1483;
assign w39864 = w1529 & w46423;
assign w39865 = ~w1716 & w1729;
assign w39866 = (~w3 & ~w1649) | (~w3 & w46424) | (~w1649 & w46424);
assign w39867 = (w3 & ~w1649) | (w3 & w46425) | (~w1649 & w46425);
assign w39868 = ~w1722 & w1758;
assign w39869 = w1649 & w46426;
assign w39870 = (w1764 & ~w1649) | (w1764 & w46427) | (~w1649 & w46427);
assign w39871 = w1649 & w46428;
assign w39872 = (w1778 & ~w1649) | (w1778 & w46429) | (~w1649 & w46429);
assign w39873 = w1649 & w46430;
assign w39874 = (w1784 & ~w1649) | (w1784 & w46431) | (~w1649 & w46431);
assign w39875 = w1649 & w46432;
assign w39876 = ~w1737 & w1794;
assign w39877 = w1649 & w46433;
assign w39878 = (w1775 & ~w1649) | (w1775 & w46434) | (~w1649 & w46434);
assign w39879 = ~w1722 & w1807;
assign w39880 = w1649 & w46435;
assign w39881 = w1649 & w46436;
assign w39882 = (w1814 & ~w1649) | (w1814 & w46437) | (~w1649 & w46437);
assign w39883 = ~w1696 & w1659;
assign w39884 = ~w1856 & ~w1857;
assign w39885 = w1874 & w43284;
assign w39886 = (w1879 & ~w1874) | (w1879 & w43285) | (~w1874 & w43285);
assign w39887 = w1888 & w43286;
assign w39888 = (w1894 & ~w1888) | (w1894 & w43287) | (~w1888 & w43287);
assign w39889 = (w43288 & w1903) | (w43288 & w46438) | (w1903 & w46438);
assign w39890 = (w1913 & w43289) | (w1913 & w1904) | (w43289 & w1904);
assign w39891 = ~w1918 & w43290;
assign w39892 = w1649 & w46439;
assign w39893 = (w1934 & ~w1649) | (w1934 & w46440) | (~w1649 & w46440);
assign w39894 = w1649 & w46441;
assign w39895 = (w1943 & ~w1649) | (w1943 & w46442) | (~w1649 & w46442);
assign w39896 = ~w1896 & ~w1930;
assign w39897 = ~w1904 & w43291;
assign w39898 = (w1959 & w1904) | (w1959 & w43292) | (w1904 & w43292);
assign w39899 = ~w1896 & w1798;
assign w39900 = w2005 & w2043;
assign w39901 = w1861 & ~w2025;
assign w39902 = ~w1861 & w2025;
assign w39903 = w2005 & w2054;
assign w39904 = ~w2004 & ~w57;
assign w39905 = ~w2061 & ~w2060;
assign w39906 = w2005 & w2064;
assign w39907 = w1956 & w1915;
assign w39908 = ~w1961 & ~w2072;
assign w39909 = w2005 & ~w1843;
assign w39910 = w1961 & w2072;
assign w39911 = ~w2081 & w3;
assign w39912 = w2005 & ~w2094;
assign w39913 = w2082 & ~w3;
assign w39914 = ~w1881 & w2117;
assign w39915 = w1881 & ~w2117;
assign w39916 = ~w2002 & w43293;
assign w39917 = ~w2005 & ~w2123;
assign w39918 = ~w2002 & w43294;
assign w39919 = (w2000 & w43295) | (w2000 & w43296) | (w43295 & w43296);
assign w39920 = w2112 & w2021;
assign w39921 = w2005 & w2140;
assign w39922 = ~w2005 & w2142;
assign w39923 = ~w2004 & ~a[97];
assign w39924 = ~w2004 & w2163;
assign w39925 = ~w2164 & ~w2162;
assign w39926 = ~w2165 & w1541;
assign w39927 = ~w2164 & w2167;
assign w39928 = w2005 & w2173;
assign w39929 = ~w2005 & ~w2172;
assign w39930 = ~w1798 & w48083;
assign w39931 = (~w612 & w1798) | (~w612 & w48084) | (w1798 & w48084);
assign w39932 = w2005 & w2201;
assign w39933 = ~w2205 & ~w1802;
assign w39934 = w2005 & w2227;
assign w39935 = w2005 & w2235;
assign w39936 = ~w2005 & w2237;
assign w39937 = ~w2004 & w2240;
assign w39938 = w2241 & ~w1826;
assign w39939 = ~w2241 & w2250;
assign w39940 = w2241 & w2252;
assign w39941 = w2005 & w2260;
assign w39942 = ~w2005 & w2262;
assign w39943 = w2005 & w2273;
assign w39944 = ~w2279 & w2289;
assign w39945 = ~w2290 & w2059;
assign w39946 = ~w2290 & w2047;
assign w39947 = ~w2311 & w1541;
assign w39948 = ~w2330 & w2176;
assign w39949 = w2330 & ~w2176;
assign w39950 = (w2133 & w2281) | (w2133 & w43297) | (w2281 & w43297);
assign w39951 = ~w2344 & ~a[97];
assign w39952 = w2334 & ~w2360;
assign w39953 = ~w2185 & ~w2374;
assign w39954 = w2147 & ~w2376;
assign w39955 = ~w2148 & w2254;
assign w39956 = ~w2385 & ~w2386;
assign w39957 = w2378 & w40834;
assign w39958 = w2148 & w2247;
assign w39959 = w2134 & ~w493;
assign w39960 = ~w2148 & w2426;
assign w39961 = w2134 & ~w754;
assign w39962 = ~w2290 & w351;
assign w39963 = ~w2491 & ~w2494;
assign w39964 = ~w2491 & w2497;
assign w39965 = ~w2285 & w48085;
assign w39966 = (~w80 & w2285) | (~w80 & w48086) | (w2285 & w48086);
assign w39967 = (~w57 & w2554) | (~w57 & w43298) | (w2554 & w43298);
assign w39968 = ~w2491 & w2553;
assign w39969 = (w2542 & w2554) | (w2542 & w43299) | (w2554 & w43299);
assign w39970 = ~w2554 & w43300;
assign w39971 = (w2620 & w2554) | (w2620 & w43301) | (w2554 & w43301);
assign w39972 = ~w2578 & w42;
assign w39973 = w2635 & ~w2633;
assign w39974 = (~w400 & w2652) | (~w400 & w43302) | (w2652 & w43302);
assign w39975 = ~w2652 & w43303;
assign w39976 = ~w2661 & ~w2662;
assign w39977 = w2558 & w43304;
assign w39978 = ~w2654 & ~w2655;
assign w39979 = w2558 & w43305;
assign w39980 = (w2674 & ~w2558) | (w2674 & w43306) | (~w2558 & w43306);
assign w39981 = w2383 & ~w2688;
assign w39982 = ~w2383 & w2474;
assign w39983 = w2383 & w2693;
assign w39984 = w2555 & w2372;
assign w39985 = ~w2704 & w754;
assign w39986 = ~w2396 & w2712;
assign w39987 = w2555 & ~w2472;
assign w39988 = ~w2717 & ~w493;
assign w39989 = ~w2395 & w2456;
assign w39990 = ~w2728 & ~w2729;
assign w39991 = ~w2730 & ~w2731;
assign w39992 = w2555 & w2743;
assign w39993 = w2555 & w2753;
assign w39994 = ~w2555 & w2755;
assign w39995 = w2555 & w2759;
assign w39996 = (w2765 & w2554) | (w2765 & w43307) | (w2554 & w43307);
assign w39997 = (~w2767 & w2554) | (~w2767 & w43308) | (w2554 & w43308);
assign w39998 = ~w2554 & w51389;
assign w39999 = ~w2555 & w2774;
assign w40000 = w2704 & ~w754;
assign w40001 = ~w2554 & w43310;
assign w40002 = (w2802 & w2554) | (w2802 & w43311) | (w2554 & w43311);
assign w40003 = ~w2554 & w43313;
assign w40004 = ~w2554 & w43314;
assign w40005 = (w2820 & w2554) | (w2820 & w43315) | (w2554 & w43315);
assign w40006 = (w2818 & w2554) | (w2818 & w43316) | (w2554 & w43316);
assign w40007 = (w2830 & w2554) | (w2830 & w43317) | (w2554 & w43317);
assign w40008 = ~w2554 & w43318;
assign w40009 = (~w2006 & w2554) | (~w2006 & w43319) | (w2554 & w43319);
assign w40010 = ~w2866 & ~w2678;
assign w40011 = w2867 & ~w2641;
assign w40012 = w2867 & ~w57;
assign w40013 = ~w2867 & w57;
assign w40014 = ~w2867 & w2645;
assign w40015 = w3002 & w3175;
assign w40016 = ~w2707 & ~w3192;
assign w40017 = ~w3195 & ~w3194;
assign w40018 = ~w3197 & w2700;
assign w40019 = ~w3193 & w3201;
assign w40020 = w3198 & ~w493;
assign w40021 = w2723 & ~w2720;
assign w40022 = ~w2680 & w46443;
assign w40023 = ~w2680 & ~w2734;
assign w40024 = w3214 & w351;
assign w40025 = (w3226 & w2864) | (w3226 & w46444) | (w2864 & w46444);
assign w40026 = ~w3198 & w493;
assign w40027 = w3236 & w3229;
assign w40028 = ~w2891 & w46445;
assign w40029 = ~w3249 & ~w3247;
assign w40030 = (w3258 & w2966) | (w3258 & w43320) | (w2966 & w43320);
assign w40031 = ~w2966 & w43321;
assign w40032 = w3262 & w2285;
assign w40033 = w2967 & w3267;
assign w40034 = ~w2891 & w46446;
assign w40035 = ~w3271 & ~w3270;
assign w40036 = (~w3276 & w2966) | (~w3276 & w43322) | (w2966 & w43322);
assign w40037 = ~w2966 & w43323;
assign w40038 = ~w2966 & w43324;
assign w40039 = (w3291 & w2966) | (w3291 & w43325) | (w2966 & w43325);
assign w40040 = ~w2967 & w3295;
assign w40041 = w2967 & w3297;
assign w40042 = w2967 & w3265;
assign w40043 = w3138 & ~w2006;
assign w40044 = ~w3138 & w2006;
assign w40045 = ~w2967 & w3322;
assign w40046 = w3118 & ~w1541;
assign w40047 = ~w2891 & w46447;
assign w40048 = ~w3337 & ~w3336;
assign w40049 = w3343 & w3348;
assign w40050 = ~w3343 & w3350;
assign w40051 = ~w3308 & w3353;
assign w40052 = (w1320 & w2966) | (w1320 & w43326) | (w2966 & w43326);
assign w40053 = w2967 & w3341;
assign w40054 = w3343 & ~w3347;
assign w40055 = ~w2967 & ~w3161;
assign w40056 = w2967 & w3367;
assign w40057 = w2967 & ~w3372;
assign w40058 = ~w3049 & ~w3387;
assign w40059 = ~w3056 & w46448;
assign w40060 = (~w3385 & w3056) | (~w3385 & w46449) | (w3056 & w46449);
assign w40061 = (w3394 & w2966) | (w3394 & w43327) | (w2966 & w43327);
assign w40062 = (w3403 & w3241) | (w3403 & w43328) | (w3241 & w43328);
assign w40063 = (w3406 & w3241) | (w3406 & w43329) | (w3241 & w43329);
assign w40064 = ~w2999 & w3414;
assign w40065 = ~w2891 & w46450;
assign w40066 = ~w3241 & w46451;
assign w40067 = ~w2891 & w46452;
assign w40068 = ~w3434 & w400;
assign w40069 = w2998 & w3438;
assign w40070 = ~w2998 & ~w3438;
assign w40071 = ~w2891 & w46453;
assign w40072 = ~w3443 & ~w612;
assign w40073 = ~w2967 & ~w3077;
assign w40074 = w2967 & w3393;
assign w40075 = ~w3171 & ~w3078;
assign w40076 = ~w2967 & w2997;
assign w40077 = ~w3241 & w46454;
assign w40078 = w3354 & w3463;
assign w40079 = ~w3241 & w46455;
assign w40080 = (w754 & w3241) | (w754 & w46456) | (w3241 & w46456);
assign w40081 = w3435 & ~w400;
assign w40082 = ~w3429 & ~w3235;
assign w40083 = ~w2891 & w46457;
assign w40084 = ~w3481 & w3479;
assign w40085 = w3480 & ~w3189;
assign w40086 = ~w3480 & ~w3479;
assign w40087 = ~w3237 & w2955;
assign w40088 = ~w2966 & w43330;
assign w40089 = (~w80 & w2966) | (~w80 & w43331) | (w2966 & w43331);
assign w40090 = (w3 & w2966) | (w3 & w43332) | (w2966 & w43332);
assign w40091 = (~w3513 & w3510) | (~w3513 & w46458) | (w3510 & w46458);
assign w40092 = (~w3516 & w3241) | (~w3516 & w43333) | (w3241 & w43333);
assign w40093 = ~w3241 & w43334;
assign w40094 = w2967 & ~w3525;
assign w40095 = w3526 & w50228;
assign w40096 = ~w3535 & ~w2890;
assign w40097 = w3535 & w3540;
assign w40098 = (w57 & w2966) | (w57 & w43335) | (w2966 & w43335);
assign w40099 = ~w3241 & w43336;
assign w40100 = (w3551 & w3241) | (w3551 & w43337) | (w3241 & w43337);
assign w40101 = ~w2967 & w3555;
assign w40102 = (w3554 & w3237) | (w3554 & w46459) | (w3237 & w46459);
assign w40103 = ~w3237 & w46460;
assign w40104 = ~w2967 & w3562;
assign w40105 = (w2953 & w2966) | (w2953 & w43338) | (w2966 & w43338);
assign w40106 = w3236 & ~w3224;
assign w40107 = ~w3241 & w43339;
assign w40108 = ~w3481 & ~w3591;
assign w40109 = w3481 & w3591;
assign w40110 = (~w351 & w3521) | (~w351 & w43340) | (w3521 & w43340);
assign w40111 = (w351 & w3521) | (w351 & w43341) | (w3521 & w43341);
assign w40112 = (w3621 & w3521) | (w3621 & w43342) | (w3521 & w43342);
assign w40113 = (w3623 & w3521) | (w3623 & w43343) | (w3521 & w43343);
assign w40114 = w3553 & w3588;
assign w40115 = ~w3652 & w3654;
assign w40116 = w3354 & w3649;
assign w40117 = w3354 & w3664;
assign w40118 = w3354 & w3647;
assign w40119 = w3354 & w3676;
assign w40120 = ~w3521 & w43344;
assign w40121 = (w3759 & ~w3639) | (w3759 & w46461) | (~w3639 & w46461);
assign w40122 = (w3765 & ~w3639) | (w3765 & w46462) | (~w3639 & w46462);
assign w40123 = ~w3521 & w43345;
assign w40124 = (~a[89] & ~w3639) | (~a[89] & w46463) | (~w3639 & w46463);
assign w40125 = ~w3521 & w43346;
assign w40126 = (w3786 & ~w3639) | (w3786 & w46464) | (~w3639 & w46464);
assign w40127 = (w3792 & ~w3639) | (w3792 & w46465) | (~w3639 & w46465);
assign w40128 = ~w3521 & w43347;
assign w40129 = ~w3643 & ~w3813;
assign w40130 = (w2558 & ~w3639) | (w2558 & w46466) | (~w3639 & w46466);
assign w40131 = ~w3308 & w1738;
assign w40132 = w3615 & ~w3598;
assign w40133 = ~w3935 & w3937;
assign w40134 = (w3579 & ~w3639) | (w3579 & w46467) | (~w3639 & w46467);
assign w40135 = (~w3952 & ~w3937) | (~w3952 & ~w3506) | (~w3937 & ~w3506);
assign w40136 = (w3519 & ~w3639) | (w3519 & w46468) | (~w3639 & w46468);
assign w40137 = w3971 & ~w3934;
assign w40138 = ~w3615 & w3971;
assign w40139 = ~w3975 & ~w3974;
assign w40140 = (w3986 & w43348) | (w3986 & ~w3976) | (w43348 & ~w3976);
assign w40141 = ~w3972 & w3976;
assign w40142 = (~w80 & w43349) | (~w80 & ~w3646) | (w43349 & ~w3646);
assign w40143 = ~w4006 & ~w4005;
assign w40144 = ~w3521 & w43350;
assign w40145 = (w4033 & w43351) | (w4033 & ~w3976) | (w43351 & ~w3976);
assign w40146 = (~w57 & w4053) | (~w57 & w46469) | (w4053 & w46469);
assign w40147 = ~w4068 & ~w4072;
assign w40148 = w4018 & ~w3888;
assign w40149 = (~w4003 & w4053) | (~w4003 & w46470) | (w4053 & w46470);
assign w40150 = ~w4055 & w4003;
assign w40151 = (~w3 & w4081) | (~w3 & w51390) | (w4081 & w51390);
assign w40152 = ~w4055 & w3636;
assign w40153 = ~w4073 & w46471;
assign w40154 = ~w4117 & w4115;
assign w40155 = ~w4056 & w43352;
assign w40156 = (w42 & w4056) | (w42 & w43353) | (w4056 & w43353);
assign w40157 = (~w4029 & w50394) | (~w4029 & w50395) | (w50394 & w50395);
assign w40158 = w44098 & w48087;
assign w40159 = ~w4152 & w4155;
assign w40160 = (w400 & w4053) | (w400 & w46472) | (w4053 & w46472);
assign w40161 = (w4029 & w49274) | (w4029 & w49275) | (w49274 & w49275);
assign w40162 = (~w4029 & w50396) | (~w4029 & w50397) | (w50396 & w50397);
assign w40163 = (w4029 & w49276) | (w4029 & w49277) | (w49276 & w49277);
assign w40164 = (~w4029 & w50398) | (~w4029 & w50399) | (w50398 & w50399);
assign w40165 = ~w4152 & w4154;
assign w40166 = ~w4176 & ~w4178;
assign w40167 = (~w3904 & w43355) | (~w3904 & w43356) | (w43355 & w43356);
assign w40168 = (~w4186 & ~w4189) | (~w4186 & w46473) | (~w4189 & w46473);
assign w40169 = ~w4190 & ~w4200;
assign w40170 = (w4215 & w4053) | (w4215 & w46474) | (w4053 & w46474);
assign w40171 = w4216 & ~w3242;
assign w40172 = (w4233 & w4053) | (w4233 & w46475) | (w4053 & w46475);
assign w40173 = ~w4053 & w46476;
assign w40174 = ~w4053 & w46477;
assign w40175 = (~w4246 & w4053) | (~w4246 & w46478) | (w4053 & w46478);
assign w40176 = ~w4053 & w46479;
assign w40177 = (w4271 & w4053) | (w4271 & w46480) | (w4053 & w46480);
assign w40178 = ~w4053 & w46481;
assign w40179 = ~w4053 & w46482;
assign w40180 = w3867 & w1738;
assign w40181 = ~w3867 & ~w1738;
assign w40182 = w4055 & ~w4309;
assign w40183 = (~w1541 & w4309) | (~w1541 & w46483) | (w4309 & w46483);
assign w40184 = w4055 & ~w4314;
assign w40185 = ~w4336 & w3836;
assign w40186 = w4336 & ~w3836;
assign w40187 = ~w3931 & w51391;
assign w40188 = (w945 & w4053) | (w945 & w46484) | (w4053 & w46484);
assign w40189 = w4055 & w4353;
assign w40190 = ~w4309 & w46485;
assign w40191 = ~w4336 & w4366;
assign w40192 = w4336 & w4368;
assign w40193 = (w3901 & w4053) | (w3901 & w46486) | (w4053 & w46486);
assign w40194 = ~w3880 & w3896;
assign w40195 = (~w3901 & w4053) | (~w3901 & w46487) | (w4053 & w46487);
assign w40196 = w43357 & w52178;
assign w40197 = w4389 & w4361;
assign w40198 = (w4080 & w51477) | (w4080 & w51478) | (w51477 & w51478);
assign w40199 = ~w4390 & w4404;
assign w40200 = (~w4407 & w4139) | (~w4407 & w46488) | (w4139 & w46488);
assign w40201 = ~w4413 & ~w4407;
assign w40202 = (w4414 & w4443) | (w4414 & w4432) | (w4443 & w4432);
assign w40203 = w4411 & ~w4114;
assign w40204 = (w1738 & w4305) | (w1738 & w48088) | (w4305 & w48088);
assign w40205 = w4275 & w4292;
assign w40206 = ~w4388 & w49278;
assign w40207 = ~w4626 & ~w4625;
assign w40208 = w4389 & ~w4651;
assign w40209 = ~w4653 & ~w4652;
assign w40210 = ~w4372 & w43359;
assign w40211 = (w1120 & w4372) | (w1120 & w43360) | (w4372 & w43360);
assign w40212 = (w4395 & w46489) | (w4395 & w46490) | (w46489 & w46490);
assign w40213 = (~w4715 & w46491) | (~w4715 & w4693) | (w46491 & w4693);
assign w40214 = ~w4443 & w43362;
assign w40215 = ~w4444 & w4756;
assign w40216 = (~w4413 & w4443) | (~w4413 & w48089) | (w4443 & w48089);
assign w40217 = (w4168 & w4693) | (w4168 & w43364) | (w4693 & w43364);
assign w40218 = w4444 & ~w4418;
assign w40219 = w4418 & ~w4150;
assign w40220 = ~w4785 & w3;
assign w40221 = ~w4780 & w3;
assign w40222 = (~w4851 & w4606) | (~w4851 & w43365) | (w4606 & w43365);
assign w40223 = ~w4833 & w4891;
assign w40224 = w4892 & w4899;
assign w40225 = ~w4892 & w4901;
assign w40226 = w4920 & w4921;
assign w40227 = ~w4920 & w4923;
assign w40228 = w4920 & w4927;
assign w40229 = ~w4920 & w4929;
assign w40230 = w4935 & w4938;
assign w40231 = ~w4935 & w4940;
assign w40232 = ~w4892 & w4949;
assign w40233 = w4892 & w4951;
assign w40234 = w4956 & a[83];
assign w40235 = ~w4833 & w4991;
assign w40236 = w4935 & w5041;
assign w40237 = ~w4935 & w5043;
assign w40238 = ~w5048 & w4889;
assign w40239 = ~w4566 & w5053;
assign w40240 = w4566 & ~w4742;
assign w40241 = ~w5054 & w43366;
assign w40242 = (w5052 & w5054) | (w5052 & w43367) | (w5054 & w43367);
assign w40243 = ~w4833 & w5061;
assign w40244 = ~w4833 & w5065;
assign w40245 = ~w4566 & ~w4724;
assign w40246 = w4566 & ~w5067;
assign w40247 = ~w4833 & w5098;
assign w40248 = ~w4833 & w5108;
assign w40249 = w5118 & w5116;
assign w40250 = ~w5118 & ~w5116;
assign w40251 = (~w4663 & w5053) | (~w4663 & w43368) | (w5053 & w43368);
assign w40252 = (w5134 & w5136) | (w5134 & w46492) | (w5136 & w46492);
assign w40253 = ~w5136 & w43369;
assign w40254 = ~w5079 & w5146;
assign w40255 = w4962 & w4746;
assign w40256 = w4962 & w5175;
assign w40257 = w5199 & w5202;
assign w40258 = ~w5199 & w5204;
assign w40259 = w5199 & w5208;
assign w40260 = ~w5199 & w5210;
assign w40261 = w4962 & w5213;
assign w40262 = ~w4814 & w4813;
assign w40263 = (w5226 & w4750) | (w5226 & w43370) | (w4750 & w43370);
assign w40264 = ~w4814 & ~w4802;
assign w40265 = (~w4818 & w4750) | (~w4818 & w43371) | (w4750 & w43371);
assign w40266 = w5252 & ~w5258;
assign w40267 = (w4835 & w4750) | (w4835 & w43372) | (w4750 & w43372);
assign w40268 = ~w4987 & w5047;
assign w40269 = ~w4987 & w5427;
assign w40270 = (~w4877 & w4955) | (~w4877 & w43373) | (w4955 & w43373);
assign w40271 = ~w5048 & w5485;
assign w40272 = ~w5048 & w4888;
assign w40273 = (w5102 & w5551) | (w5102 & w43374) | (w5551 & w43374);
assign w40274 = ~w5282 & w5224;
assign w40275 = w5329 & w5673;
assign w40276 = w5667 & w80;
assign w40277 = ~w5282 & w5223;
assign w40278 = w5682 & w5679;
assign w40279 = ~w5682 & ~w5679;
assign w40280 = w5329 & ~w5181;
assign w40281 = ~w5695 & w3;
assign w40282 = w5653 & w5724;
assign w40283 = ~w5653 & w5726;
assign w40284 = (w5746 & w5752) | (w5746 & w43375) | (w5752 & w43375);
assign w40285 = ~w5752 & w43376;
assign w40286 = ~w5732 & w49279;
assign w40287 = ~w5744 & w5756;
assign w40288 = ~w5574 & ~w5628;
assign w40289 = w5762 & w52307;
assign w40290 = w5767 & w5769;
assign w40291 = ~w5771 & w5768;
assign w40292 = ~w5574 & w5779;
assign w40293 = ~w5780 & w5627;
assign w40294 = (~w5640 & ~w5743) | (~w5640 & w46493) | (~w5743 & w46493);
assign w40295 = w5777 & w46494;
assign w40296 = (w5732 & w46495) | (w5732 & w46496) | (w46495 & w46496);
assign w40297 = w612 & w52307;
assign w40298 = w5767 & w5793;
assign w40299 = w5743 & ~w493;
assign w40300 = (w5798 & w5732) | (w5798 & w46497) | (w5732 & w46497);
assign w40301 = w5743 & w493;
assign w40302 = (w5802 & w5732) | (w5802 & w46498) | (w5732 & w46498);
assign w40303 = (w351 & ~w5777) | (w351 & w46499) | (~w5777 & w46499);
assign w40304 = (w5811 & w5732) | (w5811 & w48090) | (w5732 & w48090);
assign w40305 = (w5814 & w5732) | (w5814 & w46500) | (w5732 & w46500);
assign w40306 = w5821 & w5824;
assign w40307 = (~w5791 & w5825) | (~w5791 & w46501) | (w5825 & w46501);
assign w40308 = w5835 & ~w5834;
assign w40309 = (~w57 & ~w5745) | (~w57 & w43377) | (~w5745 & w43377);
assign w40310 = ~w5732 & w43378;
assign w40311 = w5845 & w5849;
assign w40312 = ~w5845 & w5851;
assign w40313 = ~w5732 & w46502;
assign w40314 = ~w5744 & w5860;
assign w40315 = ~w5732 & w46503;
assign w40316 = ~w5743 & w5875;
assign w40317 = w5743 & w5879;
assign w40318 = (w5732 & w49812) | (w5732 & w49813) | (w49812 & w49813);
assign w40319 = w5743 & ~w2896;
assign w40320 = ~w5900 & ~w5529;
assign w40321 = ~w5437 & ~w5586;
assign w40322 = ~w5923 & ~w5926;
assign w40323 = ~w5732 & w46504;
assign w40324 = ~w5744 & w5930;
assign w40325 = w5923 & ~w5935;
assign w40326 = ~w5923 & ~w5939;
assign w40327 = ~w5744 & w5941;
assign w40328 = w5743 & ~w5945;
assign w40329 = (~w1738 & w5732) | (~w1738 & w46505) | (w5732 & w46505);
assign w40330 = ~w5422 & w5948;
assign w40331 = ~w5732 & w46506;
assign w40332 = ~w5422 & w5967;
assign w40333 = ~w5732 & w43379;
assign w40334 = ~w5721 & w43380;
assign w40335 = (~w5981 & ~w5743) | (~w5981 & w43381) | (~w5743 & w43381);
assign w40336 = ~w5985 & ~w5986;
assign w40337 = ~w5991 & ~w4838;
assign w40338 = (w5732 & w49814) | (w5732 & w49815) | (w49814 & w49815);
assign w40339 = w5743 & w6002;
assign w40340 = ~w5743 & w6006;
assign w40341 = (~w5732 & w43382) | (~w5732 & w43383) | (w43382 & w43383);
assign w40342 = (w4430 & w5983) | (w4430 & w43384) | (w5983 & w43384);
assign w40343 = ~w6016 & ~w6033;
assign w40344 = w5373 & w52308;
assign w40345 = ~w5743 & w6039;
assign w40346 = (w5732 & w49816) | (w5732 & w49817) | (w49816 & w49817);
assign w40347 = w5388 & ~w6040;
assign w40348 = w6040 & w5361;
assign w40349 = ~w6040 & ~w5361;
assign w40350 = (w5732 & w46507) | (w5732 & w46508) | (w46507 & w46508);
assign w40351 = ~w5385 & ~w5876;
assign w40352 = w5480 & ~w5483;
assign w40353 = w6062 & ~w6066;
assign w40354 = ~w6062 & w6066;
assign w40355 = w5743 & ~w5523;
assign w40356 = ~w5744 & ~w6069;
assign w40357 = (w1320 & w5721) | (w1320 & w43385) | (w5721 & w43385);
assign w40358 = ~w5732 & w46509;
assign w40359 = (w6079 & w5732) | (w6079 & w46510) | (w5732 & w46510);
assign w40360 = ~w5732 & w46511;
assign w40361 = ~w5732 & w46512;
assign w40362 = ~w5732 & w48091;
assign w40363 = ~w6116 & w5659;
assign w40364 = ~w6116 & w6118;
assign w40365 = (~w80 & ~w5745) | (~w80 & w49818) | (~w5745 & w49818);
assign w40366 = (w6125 & ~w6116) | (w6125 & w46513) | (~w6116 & w46513);
assign w40367 = ~w6116 & w5691;
assign w40368 = ~w5821 & ~w5824;
assign w40369 = ~w5732 & w46514;
assign w40370 = w6176 & w612;
assign w40371 = (~w5502 & w6182) | (~w5502 & w46515) | (w6182 & w46515);
assign w40372 = w5744 & w6186;
assign w40373 = w5744 & w6194;
assign w40374 = ~w6176 & ~w612;
assign w40375 = w6198 & ~w6179;
assign w40376 = ~w5422 & w5820;
assign w40377 = ~w6182 & w46516;
assign w40378 = w5743 & ~w5501;
assign w40379 = w6210 & ~w945;
assign w40380 = ~w5732 & w46517;
assign w40381 = ~w5732 & w46518;
assign w40382 = ~w6212 & ~w6179;
assign w40383 = ~w5732 & w46519;
assign w40384 = (w945 & w5732) | (w945 & w46520) | (w5732 & w46520);
assign w40385 = w6160 & w6134;
assign w40386 = (w5855 & w6061) | (w5855 & w46521) | (w6061 & w46521);
assign w40387 = ~w6160 & ~w6248;
assign w40388 = ~w5721 & w43386;
assign w40389 = (w6252 & w5721) | (w6252 & w43387) | (w5721 & w43387);
assign w40390 = (w6269 & w5917) | (w6269 & w46522) | (w5917 & w46522);
assign w40391 = w5854 & w6228;
assign w40392 = w6326 & ~w6323;
assign w40393 = w6249 & w6342;
assign w40394 = (w5330 & w6344) | (w5330 & w43388) | (w6344 & w43388);
assign w40395 = w6243 & ~w4838;
assign w40396 = ~w6346 & w6376;
assign w40397 = w6243 & w6011;
assign w40398 = ~w6243 & ~w6011;
assign w40399 = w6249 & w6384;
assign w40400 = w6243 & w6402;
assign w40401 = ~w6243 & w6404;
assign w40402 = w6243 & w6033;
assign w40403 = w6243 & ~w4056;
assign w40404 = w3646 & ~w6056;
assign w40405 = ~w6114 & w6469;
assign w40406 = ~w6114 & w6484;
assign w40407 = (w6503 & w5917) | (w6503 & w46523) | (w5917 & w46523);
assign w40408 = ~w6114 & w6507;
assign w40409 = ~w6114 & w6526;
assign w40410 = (w2558 & w6454) | (w2558 & w3278) | (w6454 & w3278);
assign w40411 = w6536 & w6520;
assign w40412 = ~w6077 & w6234;
assign w40413 = w6569 & ~w945;
assign w40414 = w6570 & w43389;
assign w40415 = (~w6572 & w43390) | (~w6572 & w43391) | (w43390 & w43391);
assign w40416 = w6234 & ~w6074;
assign w40417 = ~w6110 & w5974;
assign w40418 = (w945 & w6580) | (w945 & w43392) | (w6580 & w43392);
assign w40419 = ~w6114 & w6597;
assign w40420 = ~w6264 & w49819;
assign w40421 = ~w6200 & w5831;
assign w40422 = ~w6114 & w6633;
assign w40423 = (w57 & w6264) | (w57 & w49820) | (w6264 & w49820);
assign w40424 = (~w80 & w6646) | (~w80 & w46524) | (w6646 & w46524);
assign w40425 = w6243 & ~w6667;
assign w40426 = ~w6702 & w6226;
assign w40427 = ~w6703 & w6197;
assign w40428 = ~w6212 & ~w6702;
assign w40429 = (w6112 & w49821) | (w6112 & w49822) | (w49821 & w49822);
assign w40430 = (~w6112 & w49823) | (~w6112 & w49824) | (w49823 & w49824);
assign w40431 = (w6735 & ~w6718) | (w6735 & w46525) | (~w6718 & w46525);
assign w40432 = w6584 & ~w945;
assign w40433 = ~w6593 & ~w6738;
assign w40434 = (w6318 & ~w6762) | (w6318 & w43393) | (~w6762 & w43393);
assign w40435 = w6536 & w6518;
assign w40436 = ~w6499 & w6466;
assign w40437 = w6766 & w43394;
assign w40438 = (~w6822 & ~w6762) | (~w6822 & w48092) | (~w6762 & w48092);
assign w40439 = (w6824 & ~w6762) | (w6824 & w52088) | (~w6762 & w52088);
assign w40440 = ~w6768 & w6832;
assign w40441 = (w6840 & ~w6762) | (w6840 & w48093) | (~w6762 & w48093);
assign w40442 = ~w6768 & w6853;
assign w40443 = w6766 & w43395;
assign w40444 = ~w6869 & ~w6868;
assign w40445 = ~w6768 & w6871;
assign w40446 = w6767 & ~w6877;
assign w40447 = ~w6879 & ~w6878;
assign w40448 = ~w6879 & w6883;
assign w40449 = ~w6392 & w43396;
assign w40450 = (w6969 & ~w6762) | (w6969 & w48094) | (~w6762 & w48094);
assign w40451 = w6767 & w7012;
assign w40452 = (~w7013 & ~w6762) | (~w7013 & w48095) | (~w6762 & w48095);
assign w40453 = ~w6607 & ~w7103;
assign w40454 = ~w6608 & w6746;
assign w40455 = (w7140 & ~w6762) | (w7140 & w48096) | (~w6762 & w48096);
assign w40456 = ~w6608 & w7180;
assign w40457 = w7150 & w43397;
assign w40458 = (w7224 & ~w7150) | (w7224 & w43398) | (~w7150 & w43398);
assign w40459 = ~w6768 & w7229;
assign w40460 = ~w7221 & w7234;
assign w40461 = w7221 & w7236;
assign w40462 = (~w6316 & ~w6762) | (~w6316 & w43399) | (~w6762 & w43399);
assign w40463 = (w7252 & ~w6762) | (w7252 & w43400) | (~w6762 & w43400);
assign w40464 = w6765 & ~w7260;
assign w40465 = ~w6765 & w7260;
assign w40466 = w7121 & ~w612;
assign w40467 = ~w6735 & w7296;
assign w40468 = ~w7299 & ~w400;
assign w40469 = w7192 & w351;
assign w40470 = ~w7304 & ~w7314;
assign w40471 = ~w6821 & w6796;
assign w40472 = w7331 & ~w1541;
assign w40473 = ~w7338 & ~w7009;
assign w40474 = w7333 & w7010;
assign w40475 = ~w6986 & w48097;
assign w40476 = ~w7270 & w50140;
assign w40477 = ~w7101 & w7280;
assign w40478 = ~w7101 & w7394;
assign w40479 = (w7082 & w43401) | (w7082 & w43402) | (w43401 & w43402);
assign w40480 = (~w7082 & w43403) | (~w7082 & w43404) | (w43403 & w43404);
assign w40481 = ~w7395 & w7403;
assign w40482 = w7395 & w7115;
assign w40483 = (~w612 & ~w7315) | (~w612 & w49825) | (~w7315 & w49825);
assign w40484 = (w7269 & w7082) | (w7269 & w43406) | (w7082 & w43406);
assign w40485 = w7315 & w49280;
assign w40486 = ~w7378 & w7124;
assign w40487 = w7436 & w49281;
assign w40488 = w7388 & w493;
assign w40489 = w7458 & w7455;
assign w40490 = (~w1541 & ~w7314) | (~w1541 & w49282) | (~w7314 & w49282);
assign w40491 = ~w7456 & w7021;
assign w40492 = w7458 & ~w7509;
assign w40493 = ~w7458 & w7509;
assign w40494 = ~w7526 & ~w7468;
assign w40495 = w7601 & w7603;
assign w40496 = ~w7601 & w7606;
assign w40497 = w7601 & w7614;
assign w40498 = ~w7601 & w7617;
assign w40499 = ~w7625 & w7627;
assign w40500 = w7625 & w7630;
assign w40501 = ~w6862 & ~w7637;
assign w40502 = (w7642 & w7314) | (w7642 & w49283) | (w7314 & w49283);
assign w40503 = ~w7314 & w49284;
assign w40504 = ~w7625 & w7649;
assign w40505 = w7625 & w7652;
assign w40506 = w7640 & ~w7658;
assign w40507 = ~w7640 & ~w7660;
assign w40508 = ~w7314 & w49285;
assign w40509 = (w7680 & w7314) | (w7680 & w49286) | (w7314 & w49286);
assign w40510 = ~w5330 & ~w6874;
assign w40511 = ~w7684 & w7683;
assign w40512 = w7684 & ~w7683;
assign w40513 = (w3242 & w6957) | (w3242 & w49287) | (w6957 & w49287);
assign w40514 = ~w7698 & w6982;
assign w40515 = ~w6960 & ~w3242;
assign w40516 = w6960 & w3242;
assign w40517 = ~w7709 & ~w7700;
assign w40518 = ~w7710 & w6982;
assign w40519 = w7710 & ~w6982;
assign w40520 = w7675 & w7725;
assign w40521 = ~w7675 & w7728;
assign w40522 = ~w7710 & w7750;
assign w40523 = w7710 & w7752;
assign w40524 = ~w3242 & w7754;
assign w40525 = ~w7306 & ~w7194;
assign w40526 = w7789 & w7194;
assign w40527 = (w43408 & w43407) | (w43408 & ~w7304) | (w43407 & ~w7304);
assign w40528 = ~w7805 & w252;
assign w40529 = w7301 & w7308;
assign w40530 = (w40470 & w49288) | (w40470 & w49289) | (w49288 & w49289);
assign w40531 = w43410 & ~w7315;
assign w40532 = w7805 & ~w252;
assign w40533 = ~w7828 & w7315;
assign w40534 = w7828 & ~w7315;
assign w40535 = w46526 & ~w7315;
assign w40536 = (w40470 & w49290) | (w40470 & w49291) | (w49290 & w49291);
assign w40537 = ~w7843 & w7844;
assign w40538 = w7844 & w49292;
assign w40539 = (w7886 & ~w7852) | (w7886 & w52089) | (~w7852 & w52089);
assign w40540 = ~w7843 & w7888;
assign w40541 = w7914 & ~w7910;
assign w40542 = (w7519 & w43411) | (w7519 & w43412) | (w43411 & w43412);
assign w40543 = (~w7933 & ~w7526) | (~w7933 & w49293) | (~w7526 & w49293);
assign w40544 = w7934 & ~w7932;
assign w40545 = w7923 & w7927;
assign w40546 = ~w7527 & w7946;
assign w40547 = (~w7923 & w7950) | (~w7923 & w43413) | (w7950 & w43413);
assign w40548 = w7841 & ~w493;
assign w40549 = ~w7953 & ~w7952;
assign w40550 = w7967 & w7412;
assign w40551 = ~w7967 & ~w7412;
assign w40552 = ~w7983 & w7984;
assign w40553 = w7983 & w7986;
assign w40554 = ~w7527 & ~w7989;
assign w40555 = ~w7840 & w43416;
assign w40556 = ~w7995 & ~w7996;
assign w40557 = ~w7997 & w8001;
assign w40558 = w7997 & w8003;
assign w40559 = w945 & ~w7943;
assign w40560 = ~w7983 & w8008;
assign w40561 = w7983 & w8010;
assign w40562 = (~w7932 & ~w8015) | (~w7932 & w43417) | (~w8015 & w43417);
assign w40563 = w8015 & w43418;
assign w40564 = (w7904 & w43419) | (w7904 & w43420) | (w43419 & w43420);
assign w40565 = w7997 & w8023;
assign w40566 = ~w7997 & w8025;
assign w40567 = w7967 & w8029;
assign w40568 = ~w7967 & w8031;
assign w40569 = w7427 & ~w7442;
assign w40570 = (~w400 & w8041) | (~w400 & w48098) | (w8041 & w48098);
assign w40571 = ~w8041 & w48099;
assign w40572 = ~w7903 & w8048;
assign w40573 = ~w8041 & w48100;
assign w40574 = w7783 & w351;
assign w40575 = ~w7783 & ~w351;
assign w40576 = (~w7911 & w7991) | (~w7911 & w52090) | (w7991 & w52090);
assign w40577 = ~w8078 & ~w7832;
assign w40578 = w8081 & ~w8078;
assign w40579 = w7923 & w7807;
assign w40580 = w8080 & ~w8085;
assign w40581 = w7841 & w57;
assign w40582 = ~w8089 & ~w8088;
assign w40583 = ~w7903 & w8091;
assign w40584 = w7781 & w8102;
assign w40585 = w8107 & ~w7923;
assign w40586 = ~w8107 & ~w7923;
assign w40587 = w7783 & w7832;
assign w40588 = ~w7783 & w8160;
assign w40589 = ~w7923 & w7831;
assign w40590 = w7923 & ~w7831;
assign w40591 = w7841 & ~w8210;
assign w40592 = ~w7923 & ~w8203;
assign w40593 = ~w7840 & w43421;
assign w40594 = ~w8229 & ~w8228;
assign w40595 = ~w7903 & w8231;
assign w40596 = ~w7840 & w43422;
assign w40597 = ~w8237 & ~w8236;
assign w40598 = ~w7903 & w8241;
assign w40599 = w7923 & w8246;
assign w40600 = ~w7903 & w8250;
assign w40601 = ~w7903 & w8255;
assign w40602 = ~w7903 & w8260;
assign w40603 = ~w7903 & w8270;
assign w40604 = ~w7903 & w8287;
assign w40605 = ~w7903 & w8297;
assign w40606 = ~w7840 & w43423;
assign w40607 = ~w8306 & ~w8307;
assign w40608 = ~w7903 & w8309;
assign w40609 = w7923 & w3646;
assign w40610 = ~w7923 & w8318;
assign w40611 = ~w7903 & w8344;
assign w40612 = ~w7903 & w8356;
assign w40613 = ~w7840 & w43424;
assign w40614 = ~w8375 & ~w8374;
assign w40615 = ~w7903 & w8377;
assign w40616 = ~w8389 & ~w8404;
assign w40617 = w7668 & w8409;
assign w40618 = ~w8419 & ~w8420;
assign w40619 = (w7782 & w52091) | (w7782 & w52092) | (w52091 & w52092);
assign w40620 = (~w7782 & w52093) | (~w7782 & w52094) | (w52093 & w52094);
assign w40621 = ~w7840 & w43425;
assign w40622 = ~w8432 & ~w8431;
assign w40623 = ~w7903 & w8434;
assign w40624 = (~w7782 & w52095) | (~w7782 & w52096) | (w52095 & w52096);
assign w40625 = (w7782 & w52097) | (w7782 & w52098) | (w52097 & w52098);
assign w40626 = w7668 & w7734;
assign w40627 = w7841 & ~w7762;
assign w40628 = w7841 & w8464;
assign w40629 = w7841 & w8474;
assign w40630 = w7841 & w8486;
assign w40631 = (w7482 & w7765) | (w7482 & w48101) | (w7765 & w48101);
assign w40632 = ~w7840 & w43426;
assign w40633 = ~w8506 & ~w8507;
assign w40634 = ~w8508 & w1738;
assign w40635 = w8508 & ~w1738;
assign w40636 = ~w8523 & ~w8524;
assign w40637 = w8429 & w8521;
assign w40638 = ~w8523 & w8547;
assign w40639 = ~w7527 & ~w7468;
assign w40640 = w7841 & w7524;
assign w40641 = w8448 & ~w8543;
assign w40642 = ~w8555 & ~w8556;
assign w40643 = ~w8583 & ~w1320;
assign w40644 = (w8586 & ~w8015) | (w8586 & w46528) | (~w8015 & w46528);
assign w40645 = w8015 & w46529;
assign w40646 = w8582 & w48102;
assign w40647 = (~w7945 & ~w8582) | (~w7945 & w46530) | (~w8582 & w46530);
assign w40648 = ~w8443 & w8518;
assign w40649 = ~w8157 & ~w8623;
assign w40650 = w8645 & w8647;
assign w40651 = w8157 & ~w1541;
assign w40652 = w8645 & w8497;
assign w40653 = (w8682 & w8404) | (w8682 & w46531) | (w8404 & w46531);
assign w40654 = (~w2896 & w8404) | (~w2896 & w43427) | (w8404 & w43427);
assign w40655 = (~w8458 & w8404) | (~w8458 & w46532) | (w8404 & w46532);
assign w40656 = w8157 & ~w8698;
assign w40657 = ~w8645 & w8709;
assign w40658 = w8157 & w8726;
assign w40659 = ~w8274 & w8295;
assign w40660 = w8157 & w8799;
assign w40661 = w8157 & ~w3242;
assign w40662 = w8582 & w46533;
assign w40663 = (w8979 & ~w8582) | (w8979 & w46534) | (~w8582 & w46534);
assign w40664 = w8570 & w8021;
assign w40665 = w8157 & w8997;
assign w40666 = w8157 & ~w252;
assign w40667 = w8157 & ~w7970;
assign w40668 = w8983 & ~w9090;
assign w40669 = w9092 & w52309;
assign w40670 = w8983 & w9094;
assign w40671 = ~w9095 & w52310;
assign w40672 = w8188 & w493;
assign w40673 = (~w9102 & ~w40672) | (~w9102 & w46535) | (~w40672 & w46535);
assign w40674 = ~w8188 & w8086;
assign w40675 = ~w8101 & w8086;
assign w40676 = ~w9014 & ~w8142;
assign w40677 = w9014 & w8142;
assign w40678 = w9044 & ~w8170;
assign w40679 = w9117 & w80;
assign w40680 = w8999 & ~w612;
assign w40681 = w9086 & w400;
assign w40682 = w9043 & w46536;
assign w40683 = (~w8158 & ~w9043) | (~w8158 & w46537) | (~w9043 & w46537);
assign w40684 = ~w9044 & w9160;
assign w40685 = w9120 & w3;
assign w40686 = ~w9020 & w42;
assign w40687 = w8125 & ~w9184;
assign w40688 = ~w8178 & w42;
assign w40689 = w8763 & ~w9198;
assign w40690 = ~w9210 & w9214;
assign w40691 = ~w8971 & w9252;
assign w40692 = ~w9259 & ~w9258;
assign w40693 = ~w8973 & w9229;
assign w40694 = ~w9227 & ~w9230;
assign w40695 = w9285 & w9289;
assign w40696 = ~w9285 & ~w9289;
assign w40697 = ~w8674 & ~w1320;
assign w40698 = w8674 & w1320;
assign w40699 = ~w8972 & ~w8747;
assign w40700 = ~w8971 & w8745;
assign w40701 = ~w8971 & w9339;
assign w40702 = w9342 & ~w2006;
assign w40703 = ~w7924 & ~w7315;
assign w40704 = ~w9381 & a[67];
assign w40705 = w9381 & ~a[67];
assign w40706 = w7924 & w7315;
assign w40707 = ~w9406 & w9408;
assign w40708 = w9406 & w9410;
assign w40709 = ~w9406 & w9414;
assign w40710 = w9406 & w9416;
assign w40711 = ~w9174 & ~w9178;
assign w40712 = ~w9422 & w9424;
assign w40713 = w9422 & w9426;
assign w40714 = ~w9422 & w9433;
assign w40715 = w9422 & w9435;
assign w40716 = ~w8948 & w9452;
assign w40717 = ~w8948 & w9481;
assign w40718 = w8935 & w8906;
assign w40719 = ~w9487 & ~w9488;
assign w40720 = ~w9461 & w9494;
assign w40721 = ~w9514 & w9508;
assign w40722 = w9514 & ~w9508;
assign w40723 = ~w9525 & w9528;
assign w40724 = w9535 & w9537;
assign w40725 = ~w9525 & ~w9528;
assign w40726 = w9525 & w9528;
assign w40727 = ~w9535 & w9557;
assign w40728 = w9535 & w9559;
assign w40729 = w8966 & w9574;
assign w40730 = ~w8966 & ~w9574;
assign w40731 = ~w9573 & ~w2285;
assign w40732 = w9005 & ~w9145;
assign w40733 = w9145 & w9588;
assign w40734 = ~w9589 & w9042;
assign w40735 = w9592 & w57;
assign w40736 = w9145 & ~w9587;
assign w40737 = ~w9619 & ~w9620;
assign w40738 = w9619 & w9620;
assign w40739 = w9643 & w9648;
assign w40740 = ~w80 & w9650;
assign w40741 = ~w9679 & ~w9104;
assign w40742 = ~w9694 & w9693;
assign w40743 = w9694 & ~w9693;
assign w40744 = ~w9707 & w9711;
assign w40745 = w9715 & ~w493;
assign w40746 = w9687 & w351;
assign w40747 = ~w9715 & w493;
assign w40748 = ~w9592 & ~w57;
assign w40749 = w9619 & w9747;
assign w40750 = ~w9619 & w9749;
assign w40751 = ~w9643 & ~w9647;
assign w40752 = ~w8969 & w2285;
assign w40753 = ~w8734 & w2006;
assign w40754 = w9247 & ~w9209;
assign w40755 = w9582 & w9798;
assign w40756 = w9799 & ~w9805;
assign w40757 = ~w9799 & w9805;
assign w40758 = ~w9814 & ~w9815;
assign w40759 = ~w9838 & w9553;
assign w40760 = ~w9838 & w9844;
assign w40761 = ~w9895 & w9373;
assign w40762 = w9895 & ~w9373;
assign w40763 = ~w9901 & w9903;
assign w40764 = w9901 & w9905;
assign w40765 = ~w9895 & w9908;
assign w40766 = w9895 & w9910;
assign w40767 = w9195 & w9915;
assign w40768 = w9352 & ~w9919;
assign w40769 = w9899 & w9913;
assign w40770 = ~w9395 & w9428;
assign w40771 = ~w9934 & w9437;
assign w40772 = w9935 & ~w9963;
assign w40773 = w9956 & w9965;
assign w40774 = ~w9976 & w9977;
assign w40775 = w9976 & w9979;
assign w40776 = ~w10001 & ~w4838;
assign w40777 = ~w9976 & w10015;
assign w40778 = w9976 & w10017;
assign w40779 = ~w9473 & w9495;
assign w40780 = w10031 & w10032;
assign w40781 = ~w10031 & w10034;
assign w40782 = ~w9473 & ~w9479;
assign w40783 = w9940 & ~w9470;
assign w40784 = w10047 & ~w9459;
assign w40785 = ~w10001 & w4838;
assign w40786 = ~w10061 & ~w10070;
assign w40787 = ~w9838 & ~w9551;
assign w40788 = w10031 & w10087;
assign w40789 = ~w10031 & w10089;
assign w40790 = ~w10044 & w4056;
assign w40791 = w10047 & w10097;
assign w40792 = w10100 & ~w10094;
assign w40793 = w9248 & w9769;
assign w40794 = w10111 & w43428;
assign w40795 = ~w10113 & ~w10114;
assign w40796 = w80 & w10119;
assign w40797 = ~w80 & w10122;
assign w40798 = (w9349 & w43429) | (w9349 & w43430) | (w43429 & w43430);
assign w40799 = w3 & w10136;
assign w40800 = ~w3 & w10139;
assign w40801 = ~w10107 & w10111;
assign w40802 = ~w10147 & w9738;
assign w40803 = w57 & w10153;
assign w40804 = ~w57 & w10156;
assign w40805 = ~w252 & w10166;
assign w40806 = ~w10147 & w10169;
assign w40807 = w252 & w10169;
assign w40808 = w57 & w10176;
assign w40809 = ~w57 & w10179;
assign w40810 = w80 & w10186;
assign w40811 = ~w80 & w10189;
assign w40812 = ~w9781 & w43431;
assign w40813 = (w10213 & w9781) | (w10213 & w43432) | (w9781 & w43432);
assign w40814 = ~w10146 & w10217;
assign w40815 = ~w10107 & w10219;
assign w40816 = ~w9777 & w10253;
assign w40817 = w10252 & ~w400;
assign w40818 = ~w9583 & w10106;
assign w40819 = w9777 & ~w9705;
assign w40820 = ~w9208 & w493;
assign w40821 = w9306 & w9311;
assign w40822 = ~w10281 & ~w10284;
assign w40823 = w10281 & w10284;
assign w40824 = w10290 & w612;
assign w40825 = w9208 & ~w493;
assign w40826 = w9306 & ~w10306;
assign w40827 = ~w9306 & w10306;
assign w40828 = ~w10290 & ~w612;
assign w40829 = w9769 & ~w9268;
assign w40830 = ~w1120 & ~w945;
assign w40831 = ~w10353 & ~w10354;
assign w40832 = (~w9295 & w10340) | (~w9295 & w43433) | (w10340 & w43433);
assign w40833 = (w10358 & w10340) | (w10358 & w43434) | (w10340 & w43434);
assign w40834 = w1120 & w945;
assign w40835 = ~w9781 & w43435;
assign w40836 = (w10407 & w9781) | (w10407 & w43436) | (w9781 & w43436);
assign w40837 = ~w10416 & w10218;
assign w40838 = w9863 & w10423;
assign w40839 = w10434 & ~w10369;
assign w40840 = ~w10394 & w10417;
assign w40841 = ~w10103 & w10393;
assign w40842 = w10444 & w10459;
assign w40843 = w10434 & w10352;
assign w40844 = w10388 & w10469;
assign w40845 = ~w10470 & ~w10400;
assign w40846 = w10418 & ~w754;
assign w40847 = ~w10484 & ~w10452;
assign w40848 = ~w10486 & ~w10487;
assign w40849 = ~w10494 & ~w10492;
assign w40850 = ~w10498 & w493;
assign w40851 = ~w10433 & w43437;
assign w40852 = w10510 & w10512;
assign w40853 = ~w10510 & w10514;
assign w40854 = w10388 & w10446;
assign w40855 = ~w10519 & w10453;
assign w40856 = w10418 & ~w400;
assign w40857 = ~w10524 & w10526;
assign w40858 = w10524 & w10528;
assign w40859 = ~w10532 & w10533;
assign w40860 = w10498 & ~w493;
assign w40861 = ~w10519 & w10547;
assign w40862 = w10524 & w10560;
assign w40863 = ~w10524 & w10562;
assign w40864 = w10418 & w57;
assign w40865 = ~w10246 & ~w10414;
assign w40866 = ~w10367 & ~w10402;
assign w40867 = ~w10576 & w10579;
assign w40868 = w10418 & w10583;
assign w40869 = w10576 & w10582;
assign w40870 = ~w10394 & w10597;
assign w40871 = ~w10600 & w10195;
assign w40872 = w10418 & w10603;
assign w40873 = ~w10394 & w10614;
assign w40874 = ~w10394 & w10633;
assign w40875 = w10418 & w80;
assign w40876 = w10636 & w10639;
assign w40877 = ~w10636 & w10641;
assign w40878 = (~w10578 & w10418) | (~w10578 & w43438) | (w10418 & w43438);
assign w40879 = w10654 & ~w10636;
assign w40880 = (w10396 & w43439) | (w10396 & w43440) | (w43439 & w43440);
assign w40881 = w10418 & w1120;
assign w40882 = (w10396 & w43441) | (w10396 & w43442) | (w43441 & w43442);
assign w40883 = ~w10674 & w52311;
assign w40884 = w10510 & w10362;
assign w40885 = w10431 & w10376;
assign w40886 = (~w9823 & w10689) | (~w9823 & w43443) | (w10689 & w43443);
assign w40887 = (w9836 & w10689) | (w9836 & w43444) | (w10689 & w43444);
assign w40888 = w10431 & w10734;
assign w40889 = w10418 & w10744;
assign w40890 = ~w2006 & ~w10746;
assign w40891 = ~w10753 & ~w10752;
assign w40892 = ~w10102 & ~w10389;
assign w40893 = w10418 & ~w9850;
assign w40894 = ~w10773 & w10772;
assign w40895 = w10773 & ~w10772;
assign w40896 = w10418 & w10085;
assign w40897 = (w10396 & w43445) | (w10396 & w43446) | (w43445 & w43446);
assign w40898 = w10781 & ~w10748;
assign w40899 = ~w10100 & w10785;
assign w40900 = w10418 & ~w10057;
assign w40901 = w10095 & w4056;
assign w40902 = ~w10095 & ~w4056;
assign w40903 = ~w10794 & w10795;
assign w40904 = w10794 & w10797;
assign w40905 = w10802 & w10804;
assign w40906 = ~w10802 & w10806;
assign w40907 = ~w3242 & ~w10788;
assign w40908 = ~w10794 & w10811;
assign w40909 = w10794 & w10813;
assign w40910 = ~w2558 & ~w10777;
assign w40911 = w10418 & w9850;
assign w40912 = ~w9930 & ~w10000;
assign w40913 = ~w10874 & ~w10873;
assign w40914 = ~w9930 & w10888;
assign w40915 = ~w10418 & ~w10899;
assign w40916 = w10418 & w10904;
assign w40917 = w10418 & w10914;
assign w40918 = w10802 & w10922;
assign w40919 = ~w10802 & w10924;
assign w40920 = w10394 & w10937;
assign w40921 = ~w10941 & w10944;
assign w40922 = w10418 & w10971;
assign w40923 = ~w10418 & w10965;
assign w40924 = w10418 & w11002;
assign w40925 = ~w10418 & w11004;
assign w40926 = ~w10974 & w8666;
assign w40927 = ~w10418 & w11018;
assign w40928 = ~w10956 & w11022;
assign w40929 = ~w11031 & w11033;
assign w40930 = w11031 & w11035;
assign w40931 = ~w11043 & w11045;
assign w40932 = w11043 & w11047;
assign w40933 = ~w11031 & w11066;
assign w40934 = w11031 & w11068;
assign w40935 = ~w11054 & w11071;
assign w40936 = w11054 & w11073;
assign w40937 = ~w9900 & w9912;
assign w40938 = ~w11043 & w11106;
assign w40939 = w11043 & w11108;
assign w40940 = w10418 & w11122;
assign w40941 = (w11140 & w10862) | (w11140 & w48103) | (w10862 & w48103);
assign w40942 = (~w10592 & w10570) | (~w10592 & w43447) | (w10570 & w43447);
assign w40943 = (w10683 & w10862) | (w10683 & w43448) | (w10862 & w43448);
assign w40944 = (w10684 & w10862) | (w10684 & w43449) | (w10862 & w43449);
assign w40945 = ~w11077 & ~w5330;
assign w40946 = w5330 & ~w11238;
assign w40947 = ~w5330 & ~w10903;
assign w40948 = ~w11077 & ~w10903;
assign w40949 = ~w11281 & ~w4430;
assign w40950 = ~w11280 & w50561;
assign w40951 = w11250 & ~w11255;
assign w40952 = w10932 & w10926;
assign w40953 = (w10808 & w11223) | (w10808 & w43450) | (w11223 & w43450);
assign w40954 = ~w10870 & ~w11335;
assign w40955 = w11232 & ~w11343;
assign w40956 = (w11346 & w11223) | (w11346 & w43451) | (w11223 & w43451);
assign w40957 = ~w11360 & w10764;
assign w40958 = ~w11360 & w10782;
assign w40959 = ~w11390 & w11394;
assign w40960 = w11390 & w11397;
assign w40961 = ~w11360 & w10783;
assign w40962 = w10935 & w11134;
assign w40963 = (w6264 & ~w10685) | (w6264 & w43452) | (~w10685 & w43452);
assign w40964 = w10935 & w10784;
assign w40965 = w11011 & w11026;
assign w40966 = ~w11528 & ~w11527;
assign w40967 = ~w10869 & w11536;
assign w40968 = (~w11232 & ~w11579) | (~w11232 & w43453) | (~w11579 & w43453);
assign w40969 = (~w11591 & ~w11134) | (~w11591 & w43454) | (~w11134 & w43454);
assign w40970 = ~w10869 & w11599;
assign w40971 = ~w10672 & ~a[59];
assign w40972 = (w11611 & ~w11134) | (w11611 & w43455) | (~w11134 & w43455);
assign w40973 = (~w11626 & ~w11134) | (~w11626 & w43456) | (~w11134 & w43456);
assign w40974 = w10571 & w10661;
assign w40975 = ~w10869 & w11655;
assign w40976 = ~w11598 & ~w11693;
assign w40977 = ~w11390 & w11718;
assign w40978 = w11390 & w11721;
assign w40979 = ~w10869 & w11822;
assign w40980 = ~w10869 & w11832;
assign w40981 = (w11835 & ~w11134) | (w11835 & w43457) | (~w11134 & w43457);
assign w40982 = w11138 & w42;
assign w40983 = w11862 & ~w11855;
assign w40984 = (~w11869 & w11815) | (~w11869 & w43458) | (w11815 & w43458);
assign w40985 = w11149 & ~w11874;
assign w40986 = w11864 & w7315;
assign w40987 = ~w11893 & ~w11894;
assign w40988 = ~w11865 & w11896;
assign w40989 = (w11905 & w11815) | (w11905 & w43459) | (w11815 & w43459);
assign w40990 = w11864 & w11597;
assign w40991 = ~w11865 & w11918;
assign w40992 = ~w11917 & ~w11920;
assign w40993 = w11864 & ~w11699;
assign w40994 = ~w11925 & ~w11926;
assign w40995 = ~w7315 & ~w11927;
assign w40996 = w11927 & w7315;
assign w40997 = w11864 & a[57];
assign w40998 = ~w11943 & ~w11944;
assign w40999 = (w11946 & w11815) | (w11946 & w43460) | (w11815 & w43460);
assign w41000 = (w11949 & w11815) | (w11949 & w43461) | (w11815 & w43461);
assign w41001 = (w11954 & w11815) | (w11954 & w43462) | (w11815 & w43462);
assign w41002 = (w11962 & w11815) | (w11962 & w43463) | (w11815 & w43463);
assign w41003 = w11862 & w11967;
assign w41004 = w11968 & ~w11964;
assign w41005 = ~w11970 & ~w11969;
assign w41006 = (w11981 & w11815) | (w11981 & w43464) | (w11815 & w43464);
assign w41007 = (w11983 & w11815) | (w11983 & w43465) | (w11815 & w43465);
assign w41008 = (~w11966 & w11815) | (~w11966 & w43466) | (w11815 & w43466);
assign w41009 = w11863 & w11999;
assign w41010 = ~w12001 & ~w12000;
assign w41011 = ~w12003 & ~w12007;
assign w41012 = (w12023 & w11815) | (w12023 & w43467) | (w11815 & w43467);
assign w41013 = ~w11988 & ~w12002;
assign w41014 = ~w11703 & ~w11573;
assign w41015 = ~w12068 & ~w12073;
assign w41016 = ~w11705 & w12077;
assign w41017 = w11705 & w12079;
assign w41018 = w40983 & w50562;
assign w41019 = w11705 & w12098;
assign w41020 = w12104 & ~w12099;
assign w41021 = w12107 & w12099;
assign w41022 = w40983 & w50563;
assign w41023 = w5330 & w11302;
assign w41024 = w40983 & w50564;
assign w41025 = w12144 & ~w12099;
assign w41026 = w12147 & w12099;
assign w41027 = w40983 & w49294;
assign w41028 = (w12123 & w12137) | (w12123 & w48104) | (w12137 & w48104);
assign w41029 = w11864 & w5745;
assign w41030 = ~w12177 & ~w12176;
assign w41031 = w12180 & w50230;
assign w41032 = (w11814 & w48105) | (w11814 & w48106) | (w48105 & w48106);
assign w41033 = w40983 & w49295;
assign w41034 = ~w11865 & ~w12204;
assign w41035 = ~w11869 & ~w12164;
assign w41036 = w11414 & w43468;
assign w41037 = w11414 & w49296;
assign w41038 = ~w11742 & ~w11758;
assign w41039 = ~w12218 & w12221;
assign w41040 = ~w12218 & w12232;
assign w41041 = (~w12237 & ~w12232) | (~w12237 & w43469) | (~w12232 & w43469);
assign w41042 = ~w11344 & w12249;
assign w41043 = w40983 & w50565;
assign w41044 = ~w12251 & ~w12252;
assign w41045 = (w46538 & w46539) | (w46538 & ~w11814) | (w46539 & ~w11814);
assign w41046 = (w11709 & w50566) | (w11709 & w50567) | (w50566 & w50567);
assign w41047 = ~w11344 & w12263;
assign w41048 = w11864 & w1320;
assign w41049 = ~w12265 & ~w12266;
assign w41050 = (~w11814 & w46542) | (~w11814 & w46543) | (w46542 & w46543);
assign w41051 = (w11814 & w46544) | (w11814 & w46545) | (w46544 & w46545);
assign w41052 = w12277 & w11343;
assign w41053 = w12277 & ~w40955;
assign w41054 = (w11332 & w43470) | (w11332 & w43471) | (w43470 & w43471);
assign w41055 = (w11332 & w43472) | (w11332 & w43473) | (w43472 & w43473);
assign w41056 = ~w12306 & ~w11343;
assign w41057 = ~w12306 & w40955;
assign w41058 = ~w11344 & w12320;
assign w41059 = w11864 & ~w2558;
assign w41060 = ~w12323 & ~w12324;
assign w41061 = w12318 & ~w12325;
assign w41062 = (w11814 & w48107) | (w11814 & w48108) | (w48107 & w48108);
assign w41063 = w11358 & ~w11344;
assign w41064 = w12349 & ~w12325;
assign w41065 = ~w12246 & w49297;
assign w41066 = w11864 & w3242;
assign w41067 = ~w12358 & ~w12357;
assign w41068 = w11705 & w12385;
assign w41069 = (w11814 & w46546) | (w11814 & w46547) | (w46546 & w46547);
assign w41070 = w12179 & w50230;
assign w41071 = ~w12169 & ~w12213;
assign w41072 = w11864 & w11712;
assign w41073 = ~w12424 & ~w12425;
assign w41074 = ~w12218 & w12430;
assign w41075 = (~w493 & w12431) | (~w493 & w50568) | (w12431 & w50568);
assign w41076 = ~w12431 & w50569;
assign w41077 = ~w11807 & ~w11869;
assign w41078 = ~w12457 & w12460;
assign w41079 = ~w12431 & w50570;
assign w41080 = (w493 & w12431) | (w493 & w50571) | (w12431 & w50571);
assign w41081 = w11491 & ~w11207;
assign w41082 = w11864 & w351;
assign w41083 = ~w12490 & ~w12491;
assign w41084 = w12495 & ~w12492;
assign w41085 = (w11814 & w50572) | (w11814 & w50573) | (w50572 & w50573);
assign w41086 = ~w12500 & ~w12502;
assign w41087 = ~w11344 & w12501;
assign w41088 = w12500 & w12502;
assign w41089 = w12510 & ~w57;
assign w41090 = w12525 & w351;
assign w41091 = ~w12510 & w57;
assign w41092 = ~w11870 & w11780;
assign w41093 = ~w11870 & ~w80;
assign w41094 = ~w11865 & w12544;
assign w41095 = (~w351 & w11870) | (~w351 & w43476) | (w11870 & w43476);
assign w41096 = (w11814 & w46548) | (w11814 & w46549) | (w46548 & w46549);
assign w41097 = w12562 & ~w12492;
assign w41098 = w12592 & w12565;
assign w41099 = (w11814 & w46550) | (w11814 & w46551) | (w46550 & w46551);
assign w41100 = (~w11814 & w46552) | (~w11814 & w46553) | (w46552 & w46553);
assign w41101 = (w11814 & w50574) | (w11814 & w50575) | (w50574 & w50575);
assign w41102 = w12268 & w52312;
assign w41103 = w12615 & ~w11888;
assign w41104 = w12421 & w12620;
assign w41105 = ~w12622 & w48109;
assign w41106 = ~w12581 & w49298;
assign w41107 = w12421 & w12649;
assign w41108 = w12653 & ~w12654;
assign w41109 = (w12027 & w12581) | (w12027 & w48110) | (w12581 & w48110);
assign w41110 = ~w12581 & w48111;
assign w41111 = w12421 & ~w11909;
assign w41112 = ~w12717 & w48112;
assign w41113 = (~w7924 & ~w12726) | (~w7924 & w50576) | (~w12726 & w50576);
assign w41114 = ~w12581 & w48113;
assign w41115 = (~w12034 & w12051) | (~w12034 & w50577) | (w12051 & w50577);
assign w41116 = (w12747 & w12051) | (w12747 & w50578) | (w12051 & w50578);
assign w41117 = w12615 & ~w12753;
assign w41118 = w12772 & w12613;
assign w41119 = w12615 & w12785;
assign w41120 = w12615 & w12797;
assign w41121 = (w12159 & ~w12836) | (w12159 & w43477) | (~w12836 & w43477);
assign w41122 = w12615 & w12212;
assign w41123 = ~w12836 & w43478;
assign w41124 = (~w4056 & w12836) | (~w4056 & w43479) | (w12836 & w43479);
assign w41125 = w12867 & w12157;
assign w41126 = ~w12615 & w12880;
assign w41127 = w12421 & w12402;
assign w41128 = (w12915 & w12581) | (w12915 & w48114) | (w12581 & w48114);
assign w41129 = (~w12835 & w12045) | (~w12835 & w46554) | (w12045 & w46554);
assign w41130 = w12421 & w12926;
assign w41131 = ~w12421 & ~w12192;
assign w41132 = ~w12945 & ~w12944;
assign w41133 = (~w12401 & w12581) | (~w12401 & w48115) | (w12581 & w48115);
assign w41134 = ~w12951 & w43480;
assign w41135 = ~w12958 & ~w12961;
assign w41136 = ~w12772 & ~w12581;
assign w41137 = w12940 & w12943;
assign w41138 = ~w12978 & w46555;
assign w41139 = w12615 & ~w945;
assign w41140 = ~w12214 & w12998;
assign w41141 = ~w13002 & ~w13001;
assign w41142 = w13003 & w13007;
assign w41143 = w12615 & w945;
assign w41144 = w13003 & w13023;
assign w41145 = w13003 & ~w13006;
assign w41146 = w13003 & w13037;
assign w41147 = ~w13035 & w12606;
assign w41148 = ~w13035 & w43481;
assign w41149 = ~w12999 & w13054;
assign w41150 = ~w12075 & w13092;
assign w41151 = ~w12075 & w13098;
assign w41152 = ~w13097 & w13103;
assign w41153 = ~w12075 & w12592;
assign w41154 = ~w12581 & w48116;
assign w41155 = ~w12075 & w12594;
assign w41156 = ~w12581 & w48117;
assign w41157 = ~w12581 & w48118;
assign w41158 = ~w12581 & w48119;
assign w41159 = (w13238 & w12581) | (w13238 & w48120) | (w12581 & w48120);
assign w41160 = (~w2006 & w12581) | (~w2006 & w48121) | (w12581 & w48121);
assign w41161 = ~w12583 & w50579;
assign w41162 = (~w13258 & w12583) | (~w13258 & w50580) | (w12583 & w50580);
assign w41163 = w13281 & w13287;
assign w41164 = ~w12615 & w12330;
assign w41165 = w13281 & w12331;
assign w41166 = (w2558 & w12581) | (w2558 & w48122) | (w12581 & w48122);
assign w41167 = ~w12583 & w50581;
assign w41168 = (w13314 & w12583) | (w13314 & w50582) | (w12583 & w50582);
assign w41169 = ~w12583 & w50583;
assign w41170 = (w13321 & w12583) | (w13321 & w50584) | (w12583 & w50584);
assign w41171 = ~w12583 & w50620;
assign w41172 = (w13329 & w12583) | (w13329 & w50585) | (w12583 & w50585);
assign w41173 = w12986 & ~w13349;
assign w41174 = w12974 & ~w12991;
assign w41175 = ~w13334 & w43482;
assign w41176 = ~w13334 & w43483;
assign w41177 = w12986 & ~w13774;
assign w41178 = (w13333 & w12893) | (w13333 & w48123) | (w12893 & w48123);
assign w41179 = ~w13349 & w43484;
assign w41180 = (~w13876 & w13349) | (~w13876 & w43485) | (w13349 & w43485);
assign w41181 = (w13131 & w13774) | (w13131 & w43486) | (w13774 & w43486);
assign w41182 = ~w12894 & ~w13326;
assign w41183 = ~w13957 & ~w13956;
assign w41184 = ~w13988 & w13991;
assign w41185 = w13988 & w13993;
assign w41186 = w14016 & w13818;
assign w41187 = w14035 & ~w13881;
assign w41188 = ~w14082 & w14087;
assign w41189 = w14082 & w14089;
assign w41190 = w14082 & w14098;
assign w41191 = ~w14082 & w14100;
assign w41192 = ~w14102 & w14091;
assign w41193 = ~w14075 & w14114;
assign w41194 = ~w13404 & w6769;
assign w41195 = w14143 & w14144;
assign w41196 = ~w14143 & w14146;
assign w41197 = ~w14150 & ~w14149;
assign w41198 = ~w14154 & w14156;
assign w41199 = w14154 & w14141;
assign w41200 = ~w13481 & w13406;
assign w41201 = ~w14192 & w13590;
assign w41202 = ~w14154 & w14206;
assign w41203 = w14154 & w14142;
assign w41204 = ~w14204 & ~w14200;
assign w41205 = ~w14216 & ~w14215;
assign w41206 = ~w14218 & w14230;
assign w41207 = ~w14250 & w14253;
assign w41208 = ~w13614 & ~w14266;
assign w41209 = ~w13622 & w2896;
assign w41210 = w14285 & w14284;
assign w41211 = ~w14285 & ~w14284;
assign w41212 = w14035 & ~w14308;
assign w41213 = a[51] & ~w14304;
assign w41214 = w14035 & ~w14326;
assign w41215 = w14035 & w14330;
assign w41216 = w14035 & w14359;
assign w41217 = ~w14384 & w14391;
assign w41218 = w14384 & w14393;
assign w41219 = w13668 & w9781;
assign w41220 = ~w13668 & ~w9781;
assign w41221 = w14389 & w14416;
assign w41222 = ~w14213 & w14300;
assign w41223 = (w14441 & w13738) | (w14441 & w48124) | (w13738 & w48124);
assign w41224 = w14035 & ~w1541;
assign w41225 = w14035 & w13955;
assign w41226 = ~w13738 & ~w13980;
assign w41227 = ~w14440 & w14003;
assign w41228 = (w1120 & ~w14039) | (w1120 & w49299) | (~w14039 & w49299);
assign w41229 = w14039 & w49300;
assign w41230 = w14016 & ~w14021;
assign w41231 = (w14018 & w50586) | (w14018 & w50587) | (w50586 & w50587);
assign w41232 = w14490 & w13758;
assign w41233 = ~w14490 & w14494;
assign w41234 = ~w14492 & ~w14489;
assign w41235 = (~w612 & ~w14039) | (~w612 & w49826) | (~w14039 & w49826);
assign w41236 = ~w14485 & w43488;
assign w41237 = w13738 & w14505;
assign w41238 = ~w14501 & ~w14513;
assign w41239 = w14467 & ~w14465;
assign w41240 = w13738 & w14529;
assign w41241 = w13969 & ~w1541;
assign w41242 = ~w13738 & ~w14529;
assign w41243 = w14226 & ~w14552;
assign w41244 = ~w14226 & ~w14556;
assign w41245 = ~w14267 & ~w14269;
assign w41246 = ~w14514 & w14527;
assign w41247 = w14527 & ~w14588;
assign w41248 = ~w14589 & ~w14584;
assign w41249 = w14599 & ~w80;
assign w41250 = w14596 & w80;
assign w41251 = w13815 & w14618;
assign w41252 = w13852 & w14618;
assign w41253 = w14035 & ~w14635;
assign w41254 = w14035 & w14635;
assign w41255 = w14638 & w49827;
assign w41256 = (w351 & w14039) | (w351 & w46556) | (w14039 & w46556);
assign w41257 = ~w14039 & w46557;
assign w41258 = ~w14660 & ~w13770;
assign w41259 = ~w14488 & ~w13758;
assign w41260 = ~w14658 & ~w14694;
assign w41261 = (w14696 & w48125) | (w14696 & w48126) | (w48125 & w48126);
assign w41262 = ~w14713 & ~w13932;
assign w41263 = w14035 & w13895;
assign w41264 = ~w14574 & w14588;
assign w41265 = ~w14436 & w14762;
assign w41266 = (~w14767 & ~w14696) | (~w14767 & w46559) | (~w14696 & w46559);
assign w41267 = w14696 & w46560;
assign w41268 = w14780 & ~w57;
assign w41269 = (w14778 & w48127) | (w14778 & w48128) | (w48127 & w48128);
assign w41270 = (w14671 & w14765) | (w14671 & w43489) | (w14765 & w43489);
assign w41271 = ~w14705 & w14670;
assign w41272 = ~w14833 & ~w14834;
assign w41273 = ~w14704 & ~w14843;
assign w41274 = w14844 & w48129;
assign w41275 = ~w14884 & w14885;
assign w41276 = ~w14876 & ~w14455;
assign w41277 = ~w14757 & w43490;
assign w41278 = ~w14454 & w1120;
assign w41279 = w14876 & w14517;
assign w41280 = w14759 & ~w14938;
assign w41281 = (w15020 & ~w15021) | (w15020 & w43491) | (~w15021 & w43491);
assign w41282 = w15021 & w43492;
assign w41283 = ~w14436 & w15021;
assign w41284 = ~w14213 & w15059;
assign w41285 = ~w15060 & w15066;
assign w41286 = w15064 & ~w15060;
assign w41287 = ~w14213 & ~w14297;
assign w41288 = (w14189 & w46561) | (w14189 & w46562) | (w46561 & w46562);
assign w41289 = w14759 & ~w15093;
assign w41290 = ~w15088 & w15130;
assign w41291 = (w14189 & w46563) | (w14189 & w46564) | (w46563 & w46564);
assign w41292 = (~w14189 & w46565) | (~w14189 & w46566) | (w46565 & w46566);
assign w41293 = ~w15236 & ~w15235;
assign w41294 = (~w6769 & w14761) | (~w6769 & w43493) | (w14761 & w43493);
assign w41295 = ~w14765 & w46567;
assign w41296 = (w15268 & w14765) | (w15268 & w46568) | (w14765 & w46568);
assign w41297 = (~w7315 & w15289) | (~w7315 & w43494) | (w15289 & w43494);
assign w41298 = ~w15289 & w43495;
assign w41299 = w14389 & w14395;
assign w41300 = (~w15319 & w14761) | (~w15319 & w43496) | (w14761 & w43496);
assign w41301 = ~w14761 & w43497;
assign w41302 = ~w14761 & w43498;
assign w41303 = (w15338 & w14761) | (w15338 & w43499) | (w14761 & w43499);
assign w41304 = w14759 & w14383;
assign w41305 = ~w14765 & w46569;
assign w41306 = (w15358 & w14765) | (w15358 & w46570) | (w14765 & w46570);
assign w41307 = ~w15395 & ~w15408;
assign w41308 = w14759 & ~w15425;
assign w41309 = ~w15423 & w14565;
assign w41310 = w15442 & w15444;
assign w41311 = ~w15404 & w15409;
assign w41312 = ~w14763 & w15459;
assign w41313 = w14759 & w15473;
assign w41314 = w15460 & w13384;
assign w41315 = w14759 & ~w15492;
assign w41316 = (w14761 & w43500) | (w14761 & w43501) | (w43500 & w43501);
assign w41317 = ~w15502 & ~w15412;
assign w41318 = ~w15450 & w15388;
assign w41319 = ~w15212 & ~w4838;
assign w41320 = w15172 & w4430;
assign w41321 = w15606 & w15608;
assign w41322 = w15603 & w15605;
assign w41323 = ~w15574 & ~w15620;
assign w41324 = ~w15535 & w15826;
assign w41325 = ~w15535 & w15378;
assign w41326 = ~w15537 & w15572;
assign w41327 = (w15571 & w46571) | (w15571 & w46572) | (w46571 & w46572);
assign w41328 = ~w15571 & w46573;
assign w41329 = ~w16261 & w16262;
assign w41330 = (w16273 & ~w15572) | (w16273 & w43504) | (~w15572 & w43504);
assign w41331 = (w16303 & w15620) | (w16303 & w43505) | (w15620 & w43505);
assign w41332 = (~w14969 & w43506) | (~w14969 & w15620) | (w43506 & w15620);
assign w41333 = ~w16302 & w16389;
assign w41334 = ~w16302 & w16394;
assign w41335 = ~w16422 & ~w16423;
assign w41336 = ~w15620 & w43507;
assign w41337 = ~w16455 & ~w16456;
assign w41338 = w16455 & w16456;
assign w41339 = w16400 & w16464;
assign w41340 = ~w16400 & w16466;
assign w41341 = (w14806 & w15677) | (w14806 & w46574) | (w15677 & w46574);
assign w41342 = ~w16476 & w14994;
assign w41343 = w15680 & w16481;
assign w41344 = ~w15800 & w16488;
assign w41345 = ~w16476 & w14993;
assign w41346 = w16245 & w16515;
assign w41347 = ~w16299 & w16524;
assign w41348 = w16363 & w754;
assign w41349 = w16357 & w754;
assign w41350 = ~w16515 & ~w16529;
assign w41351 = (w15640 & ~w15714) | (w15640 & w48130) | (~w15714 & w48130);
assign w41352 = w16547 & ~w15736;
assign w41353 = ~w16547 & w15736;
assign w41354 = (w41346 & w49301) | (w41346 & w49302) | (w49301 & w49302);
assign w41355 = ~w16299 & w16551;
assign w41356 = (w16565 & w16299) | (w16565 & w43508) | (w16299 & w43508);
assign w41357 = (w16537 & w16299) | (w16537 & w43509) | (w16299 & w43509);
assign w41358 = w16559 & w43510;
assign w41359 = ~w15939 & w16518;
assign w41360 = (w16518 & w16296) | (w16518 & w43511) | (w16296 & w43511);
assign w41361 = (~w16621 & w16619) | (~w16621 & w43512) | (w16619 & w43512);
assign w41362 = ~w16299 & w16550;
assign w41363 = w16541 & w945;
assign w41364 = ~w16627 & ~w16626;
assign w41365 = w16541 & ~w945;
assign w41366 = ~w16561 & w16630;
assign w41367 = ~w16617 & ~w16619;
assign w41368 = w16541 & ~w16226;
assign w41369 = w16642 & w48131;
assign w41370 = w16556 & w16672;
assign w41371 = (w945 & ~w16642) | (w945 & w48132) | (~w16642 & w48132);
assign w41372 = w16556 & w16684;
assign w41373 = ~w16694 & ~w16695;
assign w41374 = (~w16516 & ~w16704) | (~w16516 & w43513) | (~w16704 & w43513);
assign w41375 = ~w16521 & w46575;
assign w41376 = w16725 & ~w41382;
assign w41377 = ~w16726 & w16417;
assign w41378 = (w16737 & w16299) | (w16737 & w43514) | (w16299 & w43514);
assign w41379 = w16556 & w16526;
assign w41380 = ~w16556 & w16462;
assign w41381 = w16556 & w16463;
assign w41382 = (w16538 & w16299) | (w16538 & w41375) | (w16299 & w41375);
assign w41383 = ~w16556 & w16761;
assign w41384 = w16556 & w16769;
assign w41385 = (w16540 & w16299) | (w16540 & w43515) | (w16299 & w43515);
assign w41386 = w16556 & w3;
assign w41387 = w16556 & ~w16432;
assign w41388 = ~w16556 & w5330;
assign w41389 = w16556 & w16832;
assign w41390 = ~w16841 & w16842;
assign w41391 = ~w16556 & w5745;
assign w41392 = w16556 & ~w4838;
assign w41393 = ~w15939 & w16038;
assign w41394 = (~w16040 & w43516) | (~w16040 & w16867) | (w43516 & w16867);
assign w41395 = ~w16116 & w16704;
assign w41396 = ~w16893 & ~w16894;
assign w41397 = w15939 & w16901;
assign w41398 = w16907 & ~w16109;
assign w41399 = (~w16916 & ~w16915) | (~w16916 & w48133) | (~w16915 & w48133);
assign w41400 = w16556 & w16110;
assign w41401 = w16917 & ~w2006;
assign w41402 = ~w16914 & w16096;
assign w41403 = w16933 & ~w2285;
assign w41404 = ~w16909 & w16915;
assign w41405 = w16983 & ~w16988;
assign w41406 = ~w16983 & w16988;
assign w41407 = ~w16556 & ~w16994;
assign w41408 = ~w16996 & w3646;
assign w41409 = ~w17000 & ~w16999;
assign w41410 = ~w16556 & ~w16108;
assign w41411 = w17026 & ~w2896;
assign w41412 = (~w15886 & w16842) | (~w15886 & w43517) | (w16842 & w43517);
assign w41413 = ~w17065 & w43518;
assign w41414 = (w7315 & w17065) | (w7315 & w43519) | (w17065 & w43519);
assign w41415 = w16556 & ~w17081;
assign w41416 = ~w17114 & ~w17113;
assign w41417 = ~w17116 & ~w17117;
assign w41418 = ~w15727 & w15739;
assign w41419 = w16556 & w10419;
assign w41420 = w16556 & ~w17142;
assign w41421 = ~w17155 & w43520;
assign w41422 = ~w16556 & ~w15807;
assign w41423 = ~w17170 & w8666;
assign w41424 = ~w16556 & w15808;
assign w41425 = w17168 & w9195;
assign w41426 = w17170 & ~w8666;
assign w41427 = (~w17123 & w17184) | (~w17123 & w48134) | (w17184 & w48134);
assign w41428 = w16556 & w17205;
assign w41429 = ~w16556 & w17207;
assign w41430 = ~w16556 & w17214;
assign w41431 = w16556 & w17213;
assign w41432 = w16556 & w17219;
assign w41433 = ~w16556 & w17221;
assign w41434 = ~w16299 & w17259;
assign w41435 = w16556 & w17270;
assign w41436 = w16556 & w17280;
assign w41437 = ~w17286 & w10419;
assign w41438 = w16541 & w17302;
assign w41439 = ~w16299 & w17305;
assign w41440 = ~w16556 & ~w15639;
assign w41441 = w16556 & w17318;
assign w41442 = w17292 & ~w17275;
assign w41443 = ~w16979 & w17351;
assign w41444 = ~w17352 & w16830;
assign w41445 = w17224 & ~w17328;
assign w41446 = ~w17396 & ~w17140;
assign w41447 = (~w9195 & w17356) | (~w9195 & w48135) | (w17356 & w48135);
assign w41448 = ~w17396 & w17430;
assign w41449 = ~w17343 & ~w17189;
assign w41450 = (w17351 & w17194) | (w17351 & w48136) | (w17194 & w48136);
assign w41451 = ~w17443 & ~w6769;
assign w41452 = w17450 & w43521;
assign w41453 = w17507 & ~w17514;
assign w41454 = (~w17350 & w17194) | (~w17350 & w48137) | (w17194 & w48137);
assign w41455 = (~w17531 & w17194) | (~w17531 & w48138) | (w17194 & w48138);
assign w41456 = ~w17194 & w48139;
assign w41457 = ~w17356 & w48140;
assign w41458 = ~w17343 & w17541;
assign w41459 = (w17570 & w17194) | (w17570 & w48141) | (w17194 & w48141);
assign w41460 = ~w17195 & w17737;
assign w41461 = (w16949 & w17747) | (w16949 & w43522) | (w17747 & w43522);
assign w41462 = ~w17747 & w43523;
assign w41463 = ~w17745 & ~w17747;
assign w41464 = ~w17791 & ~w2558;
assign w41465 = (w17804 & w17448) | (w17804 & w43524) | (w17448 & w43524);
assign w41466 = ~w17051 & w48142;
assign w41467 = ~w17375 & w43525;
assign w41468 = ~w17051 & w48143;
assign w41469 = ~w16979 & w17363;
assign w41470 = ~w18079 & ~w16636;
assign w41471 = ~w17051 & w48144;
assign w41472 = w16723 & w18108;
assign w41473 = w17753 & w18116;
assign w41474 = ~w17380 & ~w17846;
assign w41475 = ~w18089 & ~w18126;
assign w41476 = w17379 & w612;
assign w41477 = w18128 & w18132;
assign w41478 = ~w18128 & w18134;
assign w41479 = ~w18139 & ~w18138;
assign w41480 = ~w18139 & w18142;
assign w41481 = w18141 & w18148;
assign w41482 = w18141 & w18159;
assign w41483 = ~w18020 & ~w351;
assign w41484 = w18163 & ~w18165;
assign w41485 = ~w18128 & w18167;
assign w41486 = w18128 & w18169;
assign w41487 = ~w18173 & ~w18166;
assign w41488 = ~w18182 & ~w17395;
assign w41489 = w18182 & w18189;
assign w41490 = ~w18194 & ~w17697;
assign w41491 = ~w18182 & ~w17688;
assign w41492 = w18207 & w10419;
assign w41493 = ~w18182 & w17680;
assign w41494 = w18216 & w11138;
assign w41495 = ~w18207 & ~w10419;
assign w41496 = ~w18182 & w18231;
assign w41497 = ~w18238 & ~w17416;
assign w41498 = ~w18182 & w18243;
assign w41499 = ~w18184 & ~w17720;
assign w41500 = ~w18182 & w18254;
assign w41501 = ~w18182 & w18259;
assign w41502 = ~w18182 & ~w17405;
assign w41503 = ~w17731 & ~w17423;
assign w41504 = ~w18182 & ~w17475;
assign w41505 = ~w18182 & ~w7924;
assign w41506 = w18182 & w18269;
assign w41507 = ~w18276 & w18286;
assign w41508 = ~w18297 & w18300;
assign w41509 = ~w18182 & w17523;
assign w41510 = w18305 & w4056;
assign w41511 = ~w17582 & w18298;
assign w41512 = ~w18182 & w18316;
assign w41513 = ~w18309 & w18323;
assign w41514 = ~w18182 & w18326;
assign w41515 = ~w18337 & ~w17581;
assign w41516 = ~w18182 & w18356;
assign w41517 = ~w17731 & w18368;
assign w41518 = ~w18182 & w18379;
assign w41519 = w18182 & w18402;
assign w41520 = w18403 & ~w16559;
assign w41521 = ~w18182 & w18415;
assign w41522 = w18182 & w18414;
assign w41523 = ~w18408 & w15681;
assign w41524 = w18182 & ~w18430;
assign w41525 = ~w18182 & ~w17595;
assign w41526 = w18182 & w18470;
assign w41527 = w18182 & ~w18487;
assign w41528 = w18182 & w18499;
assign w41529 = ~w18182 & ~w17696;
assign w41530 = w18182 & w18508;
assign w41531 = w18482 & w18515;
assign w41532 = ~w18216 & ~w11138;
assign w41533 = ~w18053 & w18538;
assign w41534 = ~w18543 & ~w17814;
assign w41535 = ~w18053 & w18553;
assign w41536 = ~w18051 & ~w18556;
assign w41537 = w18051 & w18556;
assign w41538 = ~w18182 & w17812;
assign w41539 = ~w18543 & ~w18567;
assign w41540 = ~w18570 & w18566;
assign w41541 = w18570 & w18571;
assign w41542 = ~w18053 & w18575;
assign w41543 = ~w18578 & w18581;
assign w41544 = ~w18583 & w18584;
assign w41545 = w18583 & w18586;
assign w41546 = ~w18570 & w17814;
assign w41547 = w18570 & ~w17814;
assign w41548 = ~w18606 & ~w18612;
assign w41549 = w18621 & ~w18623;
assign w41550 = w17912 & w18641;
assign w41551 = ~w18182 & w18648;
assign w41552 = ~w18611 & w18653;
assign w41553 = ~w18583 & w17773;
assign w41554 = w18583 & ~w17773;
assign w41555 = ~w18053 & w18671;
assign w41556 = ~w18182 & ~w2006;
assign w41557 = w18674 & w18677;
assign w41558 = ~w18674 & w18679;
assign w41559 = w17582 & w17556;
assign w41560 = ~w18686 & w18690;
assign w41561 = ~w18182 & w17566;
assign w41562 = ~w18698 & w3242;
assign w41563 = ~w17584 & w18702;
assign w41564 = ~w18706 & w18708;
assign w41565 = w18706 & w18710;
assign w41566 = w18698 & ~w3242;
assign w41567 = ~w18686 & w17895;
assign w41568 = ~w18182 & w18719;
assign w41569 = ~w18182 & w18726;
assign w41570 = ~w18706 & w18733;
assign w41571 = w18706 & w18735;
assign w41572 = w18182 & ~w18743;
assign w41573 = w18182 & w18743;
assign w41574 = ~w18754 & w18756;
assign w41575 = ~w18759 & ~w18758;
assign w41576 = ~w18757 & ~w18763;
assign w41577 = w18077 & w612;
assign w41578 = ~w18124 & ~w18768;
assign w41579 = w18124 & ~w18174;
assign w41580 = ~w18124 & ~w18776;
assign w41581 = w18124 & ~w18121;
assign w41582 = ~w18182 & w18802;
assign w41583 = ~w18182 & w18808;
assign w41584 = ~w18182 & ~w17537;
assign w41585 = ~w18831 & ~w18832;
assign w41586 = w17577 & ~w3646;
assign w41587 = w18674 & ~w18676;
assign w41588 = ~w18674 & w18676;
assign w41589 = w18633 & w1541;
assign w41590 = ~w18179 & w18006;
assign w41591 = ~w18863 & w18866;
assign w41592 = w18182 & ~w18044;
assign w41593 = ~w18182 & w17974;
assign w41594 = ~w18887 & w42;
assign w41595 = ~w18913 & ~w18914;
assign w41596 = w18913 & w18914;
assign w41597 = w18179 & ~w18023;
assign w41598 = w18922 & ~w18921;
assign w41599 = ~w18930 & w57;
assign w41600 = w18910 & w18936;
assign w41601 = ~w18910 & w18938;
assign w41602 = (w18942 & w18457) | (w18942 & w48145) | (w18457 & w48145);
assign w41603 = ~w18457 & w48146;
assign w41604 = (w18945 & w18457) | (w18945 & w48147) | (w18457 & w48147);
assign w41605 = ~w18182 & w18022;
assign w41606 = ~w18457 & w48148;
assign w41607 = ~w18959 & ~w18178;
assign w41608 = w18964 & ~w18960;
assign w41609 = ~w18965 & w18171;
assign w41610 = ~w18182 & ~w400;
assign w41611 = ~w18965 & w18974;
assign w41612 = ~w18182 & w612;
assign w41613 = w18760 & ~w18175;
assign w41614 = ~w18981 & w18985;
assign w41615 = w18981 & w18987;
assign w41616 = ~w18995 & ~w18997;
assign w41617 = w18981 & w19001;
assign w41618 = ~w18981 & w19003;
assign w41619 = ~w18965 & w19010;
assign w41620 = ~w19026 & w18920;
assign w41621 = ~w18981 & ~w18984;
assign w41622 = w18981 & w18984;
assign w41623 = w19026 & ~w19037;
assign w41624 = ~w19039 & ~w18789;
assign w41625 = w18730 & ~w18838;
assign w41626 = ~w19063 & w2285;
assign w41627 = w18730 & ~w18701;
assign w41628 = ~w19100 & ~w2558;
assign w41629 = w18534 & w19106;
assign w41630 = ~w18730 & ~w18835;
assign w41631 = w19039 & ~w18700;
assign w41632 = (~w2896 & w19030) | (~w2896 & w43526) | (w19030 & w43526);
assign w41633 = ~w19030 & w43527;
assign w41634 = w18730 & w19130;
assign w41635 = ~w19139 & w19140;
assign w41636 = w19139 & w19142;
assign w41637 = (w18668 & w19150) | (w18668 & w43528) | (w19150 & w43528);
assign w41638 = ~w19139 & w19165;
assign w41639 = w19139 & w19167;
assign w41640 = w19116 & w2896;
assign w41641 = ~w19139 & w19203;
assign w41642 = w19139 & w19205;
assign w41643 = ~w2006 & ~w19161;
assign w41644 = ~w19139 & w18594;
assign w41645 = w19139 & ~w18594;
assign w41646 = ~w19223 & w18800;
assign w41647 = ~w19238 & w43529;
assign w41648 = (w19221 & w19238) | (w19221 & w43530) | (w19238 & w43530);
assign w41649 = w19039 & ~w4430;
assign w41650 = ~w19030 & w43531;
assign w41651 = (w19255 & w19030) | (w19255 & w43532) | (w19030 & w43532);
assign w41652 = ~w19266 & ~w19267;
assign w41653 = ~w18597 & w18682;
assign w41654 = ~w19278 & ~w18844;
assign w41655 = ~w19283 & ~w19284;
assign w41656 = ~w19217 & w19289;
assign w41657 = w19294 & ~w8666;
assign w41658 = ~w19313 & ~w18221;
assign w41659 = w19039 & w19319;
assign w41660 = ~w19298 & w18258;
assign w41661 = ~w19039 & w19329;
assign w41662 = ~w19334 & w7924;
assign w41663 = ~w19294 & w19339;
assign w41664 = ~w19039 & w19341;
assign w41665 = ~w19298 & w19348;
assign w41666 = ~w19039 & w19351;
assign w41667 = ~w19353 & w19356;
assign w41668 = w19353 & w19359;
assign w41669 = w19334 & ~w7924;
assign w41670 = ~w19298 & w18264;
assign w41671 = w19353 & w19380;
assign w41672 = ~w19017 & ~w19024;
assign w41673 = w19039 & w19442;
assign w41674 = ~w19039 & ~w19444;
assign w41675 = w18862 & w19450;
assign w41676 = ~w19039 & w19475;
assign w41677 = w19039 & w19484;
assign w41678 = w19039 & w18477;
assign w41679 = ~w19039 & w19496;
assign w41680 = ~w19039 & w19501;
assign w41681 = ~w19039 & w19510;
assign w41682 = w18482 & w18514;
assign w41683 = ~w19537 & ~w19536;
assign w41684 = w19555 & w10419;
assign w41685 = w19569 & w11870;
assign w41686 = ~w19039 & w19575;
assign w41687 = w19039 & w19583;
assign w41688 = ~w19039 & w19585;
assign w41689 = w19039 & w19598;
assign w41690 = ~w19039 & w19600;
assign w41691 = w19039 & w19603;
assign w41692 = ~w19039 & w19605;
assign w41693 = ~w19569 & ~w11870;
assign w41694 = w19616 & w19565;
assign w41695 = ~w19554 & ~w10419;
assign w41696 = w19564 & ~w19620;
assign w41697 = w19223 & w18533;
assign w41698 = w18288 & ~w18799;
assign w41699 = w19039 & w19641;
assign w41700 = w19039 & w19653;
assign w41701 = ~w19039 & ~w19663;
assign w41702 = w19217 & ~w19678;
assign w41703 = w19660 & w18797;
assign w41704 = w19039 & w19690;
assign w41705 = ~w19701 & w19671;
assign w41706 = w19039 & w19747;
assign w41707 = ~w19742 & w19751;
assign w41708 = w19039 & w18752;
assign w41709 = ~w19754 & ~w19052;
assign w41710 = ~w19764 & w19767;
assign w41711 = w19764 & w19770;
assign w41712 = w19039 & w19780;
assign w41713 = ~w19742 & w19784;
assign w41714 = w19039 & ~w945;
assign w41715 = ~w19039 & w19050;
assign w41716 = w19793 & w43533;
assign w41717 = ~w19808 & ~w19812;
assign w41718 = ~w19039 & ~w18934;
assign w41719 = w18861 & w19016;
assign w41720 = w19819 & w50231;
assign w41721 = (~w18827 & w43534) | (~w18827 & w43535) | (w43534 & w43535);
assign w41722 = ~w19036 & ~w19024;
assign w41723 = ~w18861 & w19037;
assign w41724 = (~w42 & ~w19040) | (~w42 & w43536) | (~w19040 & w43536);
assign w41725 = ~w18955 & w52313;
assign w41726 = ~w19039 & w19846;
assign w41727 = (~w80 & w19841) | (~w80 & w43537) | (w19841 & w43537);
assign w41728 = ~w19818 & w50231;
assign w41729 = w19856 & w18978;
assign w41730 = w19039 & ~w252;
assign w41731 = (w18827 & w48149) | (w18827 & w48150) | (w48149 & w48150);
assign w41732 = ~w19039 & w19879;
assign w41733 = w18861 & w19881;
assign w41734 = ~w18861 & w19884;
assign w41735 = w19039 & ~w19893;
assign w41736 = ~w18861 & ~w19034;
assign w41737 = ~w19899 & w19905;
assign w41738 = ~w19908 & w19909;
assign w41739 = w19908 & w19911;
assign w41740 = w19040 & w43538;
assign w41741 = ~w19854 & w19942;
assign w41742 = (w19949 & w19030) | (w19949 & w48151) | (w19030 & w48151);
assign w41743 = ~w19030 & w48152;
assign w41744 = ~w19908 & w19959;
assign w41745 = w19908 & w19961;
assign w41746 = ~w19854 & w19973;
assign w41747 = w19814 & ~w19974;
assign w41748 = ~w19708 & ~w19999;
assign w41749 = ~w19734 & ~w20001;
assign w41750 = ~w19671 & ~w19659;
assign w41751 = ~w19416 & w20035;
assign w41752 = w20044 & ~w19171;
assign w41753 = ~w20044 & w20064;
assign w41754 = (w19986 & w19736) | (w19986 & w19999) | (w19736 & w19999);
assign w41755 = ~w20033 & w20077;
assign w41756 = ~w20000 & ~w20070;
assign w41757 = w20122 & ~w20128;
assign w41758 = ~w20122 & w20128;
assign w41759 = ~w20044 & w20141;
assign w41760 = w20000 & w20145;
assign w41761 = ~w20000 & w20147;
assign w41762 = w20172 & ~w2285;
assign w41763 = ~w20171 & w2285;
assign w41764 = ~w20174 & w20191;
assign w41765 = ~w20196 & w2558;
assign w41766 = w20197 & ~w2558;
assign w41767 = ~w20121 & w20228;
assign w41768 = ~w20233 & ~w20232;
assign w41769 = ~w19631 & w43539;
assign w41770 = (~w20301 & w19631) | (~w20301 & w43540) | (w19631 & w43540);
assign w41771 = (~w20318 & w19999) | (~w20318 & w43541) | (w19999 & w43541);
assign w41772 = ~w19999 & w43542;
assign w41773 = (w20334 & w19999) | (w20334 & w43543) | (w19999 & w43543);
assign w41774 = ~w19999 & w43544;
assign w41775 = (w20361 & w19999) | (w20361 & w43545) | (w19999 & w43545);
assign w41776 = ~w19999 & w43546;
assign w41777 = w20206 & w20150;
assign w41778 = ~w20456 & ~w20460;
assign w41779 = w20456 & w20471;
assign w41780 = ~w20456 & w20473;
assign w41781 = w20479 & w20483;
assign w41782 = ~w20479 & w20485;
assign w41783 = ~w20479 & ~w20482;
assign w41784 = w20479 & w20482;
assign w41785 = (~w20637 & w19999) | (~w20637 & w43547) | (w19999 & w43547);
assign w41786 = (~w20639 & w19999) | (~w20639 & w46576) | (w19999 & w46576);
assign w41787 = (w20668 & w19999) | (w20668 & w43548) | (w19999 & w43548);
assign w41788 = ~w19999 & w43549;
assign w41789 = (w10419 & w19999) | (w10419 & w43550) | (w19999 & w43550);
assign w41790 = (w20736 & w19999) | (w20736 & w43551) | (w19999 & w43551);
assign w41791 = ~w19999 & w43552;
assign w41792 = ~w20716 & ~w20752;
assign w41793 = (~w20226 & w20108) | (~w20226 & w46577) | (w20108 & w46577);
assign w41794 = ~w20716 & w20775;
assign w41795 = ~w19734 & w19982;
assign w41796 = ~w20542 & ~w20621;
assign w41797 = ~w20542 & w20938;
assign w41798 = ~w20624 & w43553;
assign w41799 = ~w20624 & w43554;
assign w41800 = w20715 & w20760;
assign w41801 = ~w21255 & w21261;
assign w41802 = (~w21324 & ~w21322) | (~w21324 & w43555) | (~w21322 & w43555);
assign w41803 = ~w20170 & ~w20221;
assign w41804 = (w21442 & w20781) | (w21442 & w43556) | (w20781 & w43556);
assign w41805 = (w20201 & w20781) | (w20201 & w43557) | (w20781 & w43557);
assign w41806 = (w21473 & w20781) | (w21473 & w43558) | (w20781 & w43558);
assign w41807 = ~w21494 & w21497;
assign w41808 = ~w21494 & ~w21491;
assign w41809 = (w21566 & w20910) | (w21566 & w43559) | (w20910 & w43559);
assign w41810 = ~w20910 & w43560;
assign w41811 = (w20384 & w20910) | (w20384 & w43561) | (w20910 & w43561);
assign w41812 = ~w20910 & w43562;
assign w41813 = w21708 & w48153;
assign w41814 = ~w21794 & ~w21806;
assign w41815 = w21815 & ~w21812;
assign w41816 = ~w21705 & w21827;
assign w41817 = w21709 & w21838;
assign w41818 = w21709 & ~w21838;
assign w41819 = (w493 & ~w21708) | (w493 & w48154) | (~w21708 & w48154);
assign w41820 = w21702 & ~w21697;
assign w41821 = w21708 & w48155;
assign w41822 = w21708 & w48156;
assign w41823 = w21708 & w48157;
assign w41824 = w21873 & w48158;
assign w41825 = (~w21792 & w21490) | (~w21792 & w48159) | (w21490 & w48159);
assign w41826 = (w21380 & ~w21879) | (w21380 & w48160) | (~w21879 & w48160);
assign w41827 = ~w21880 & w21881;
assign w41828 = ~w21709 & ~w252;
assign w41829 = w21708 & w48161;
assign w41830 = ~w21794 & w21825;
assign w41831 = (w57 & ~w21708) | (w57 & w48162) | (~w21708 & w48162);
assign w41832 = ~w21800 & w48163;
assign w41833 = (~w21904 & w21800) | (~w21904 & w48164) | (w21800 & w48164);
assign w41834 = ~w21703 & w21925;
assign w41835 = w21909 & ~w21651;
assign w41836 = w21709 & ~w21940;
assign w41837 = w21911 & w21947;
assign w41838 = ~w21911 & w21949;
assign w41839 = ~w21971 & w21972;
assign w41840 = ~w21709 & w21975;
assign w41841 = ~w21709 & w21978;
assign w41842 = w21971 & ~w21972;
assign w41843 = w21706 & ~w21881;
assign w41844 = ~w21709 & w21994;
assign w41845 = w21880 & w21881;
assign w41846 = ~w21998 & ~w612;
assign w41847 = w21708 & w46578;
assign w41848 = w21761 & w21507;
assign w41849 = ~w22016 & ~w22015;
assign w41850 = ~w22036 & ~w22035;
assign w41851 = ~w22037 & w21792;
assign w41852 = ~w22027 & w945;
assign w41853 = ~w21709 & w21434;
assign w41854 = w21708 & w46579;
assign w41855 = ~w21756 & w22009;
assign w41856 = w22072 & w2285;
assign w41857 = w22076 & w21785;
assign w41858 = ~w22076 & ~w21785;
assign w41859 = w21761 & w22081;
assign w41860 = ~w22092 & ~w22091;
assign w41861 = w22103 & ~w21778;
assign w41862 = ~w21709 & w22109;
assign w41863 = w22093 & w21779;
assign w41864 = w22105 & ~w1738;
assign w41865 = ~w21709 & ~w1738;
assign w41866 = ~w22103 & w22126;
assign w41867 = w22111 & ~w1738;
assign w41868 = w22121 & w22138;
assign w41869 = ~w22121 & w22140;
assign w41870 = w21780 & w22100;
assign w41871 = ~w21709 & w1541;
assign w41872 = w21709 & w21485;
assign w41873 = ~w21709 & w22160;
assign w41874 = w21709 & w22162;
assign w41875 = ~w21709 & w22166;
assign w41876 = w21709 & w22168;
assign w41877 = ~w22019 & w22007;
assign w41878 = w22003 & w22178;
assign w41879 = ~w22003 & w22180;
assign w41880 = ~w22111 & w1738;
assign w41881 = w22076 & w22192;
assign w41882 = ~w22076 & w22194;
assign w41883 = (w22216 & ~w21708) | (w22216 & w48165) | (~w21708 & w48165);
assign w41884 = w21708 & w48166;
assign w41885 = (w22225 & ~w21708) | (w22225 & w48167) | (~w21708 & w48167);
assign w41886 = w21708 & w48168;
assign w41887 = w21708 & w48169;
assign w41888 = (w22221 & ~w21708) | (w22221 & w48170) | (~w21708 & w48170);
assign w41889 = w21708 & w48171;
assign w41890 = w21708 & w48172;
assign w41891 = (w21120 & ~w21708) | (w21120 & w48173) | (~w21708 & w48173);
assign w41892 = w21708 & w48174;
assign w41893 = w21708 & w48175;
assign w41894 = ~w22308 & w22310;
assign w41895 = w22308 & w22312;
assign w41896 = ~w21005 & w21248;
assign w41897 = ~w22320 & w22321;
assign w41898 = w22320 & w22323;
assign w41899 = w21134 & ~w20998;
assign w41900 = w21709 & ~w22339;
assign w41901 = w21709 & w22350;
assign w41902 = ~w21709 & w22330;
assign w41903 = w21709 & ~w22348;
assign w41904 = ~w21127 & ~w21131;
assign w41905 = ~w22380 & w22382;
assign w41906 = w22380 & w22384;
assign w41907 = ~w22392 & ~w22393;
assign w41908 = ~w21709 & w22407;
assign w41909 = ~w21134 & w22417;
assign w41910 = ~w21709 & w20947;
assign w41911 = w21709 & ~w22429;
assign w41912 = ~w21709 & w22447;
assign w41913 = w21708 & w48176;
assign w41914 = w21708 & w48177;
assign w41915 = w22474 & w22326;
assign w41916 = w21709 & ~w22438;
assign w41917 = ~w22380 & w22487;
assign w41918 = w22380 & w22489;
assign w41919 = w22308 & ~w22309;
assign w41920 = ~w22308 & w22309;
assign w41921 = ~w22315 & w21237;
assign w41922 = ~w22512 & w22508;
assign w41923 = w22512 & ~w22508;
assign w41924 = ~w22320 & w21221;
assign w41925 = w22320 & ~w21221;
assign w41926 = ~w22315 & w22525;
assign w41927 = (~w21214 & ~w21708) | (~w21214 & w46580) | (~w21708 & w46580);
assign w41928 = (~w7315 & w21800) | (~w7315 & w46581) | (w21800 & w46581);
assign w41929 = w21170 & ~w22535;
assign w41930 = (~w21298 & ~w21708) | (~w21298 & w46582) | (~w21708 & w46582);
assign w41931 = (~w5745 & w21800) | (~w5745 & w46583) | (w21800 & w46583);
assign w41932 = ~w22535 & ~w21299;
assign w41933 = w21170 & ~w21299;
assign w41934 = ~w22548 & ~w22547;
assign w41935 = w22548 & w22547;
assign w41936 = ~w22315 & w21238;
assign w41937 = ~w21800 & w46584;
assign w41938 = ~w22315 & w22571;
assign w41939 = ~w21709 & w22581;
assign w41940 = ~w21709 & w22590;
assign w41941 = ~w21709 & w22595;
assign w41942 = (~w5330 & ~w21708) | (~w5330 & w46585) | (~w21708 & w46585);
assign w41943 = w22604 & w22611;
assign w41944 = w22586 & w22534;
assign w41945 = ~w22617 & w22522;
assign w41946 = ~w22623 & ~w21768;
assign w41947 = w21708 & w46586;
assign w41948 = w21708 & w46587;
assign w41949 = (~w22659 & ~w21708) | (~w22659 & w48178) | (~w21708 & w48178);
assign w41950 = ~w21757 & w48179;
assign w41951 = ~w22623 & ~w22661;
assign w41952 = w21170 & w21749;
assign w41953 = w21357 & ~w21752;
assign w41954 = ~w21800 & w48180;
assign w41955 = (w22683 & w21800) | (w22683 & w48181) | (w21800 & w48181);
assign w41956 = ~w21800 & w48182;
assign w41957 = (w22693 & w21800) | (w22693 & w48183) | (w21800 & w48183);
assign w41958 = (~w21350 & ~w21708) | (~w21350 & w48184) | (~w21708 & w48184);
assign w41959 = ~w21800 & w48185;
assign w41960 = (w22712 & w21254) | (w22712 & w43563) | (w21254 & w43563);
assign w41961 = (~w4838 & ~w21708) | (~w4838 & w46588) | (~w21708 & w46588);
assign w41962 = ~w21800 & w46589;
assign w41963 = (~w22734 & w21800) | (~w22734 & w46590) | (w21800 & w46590);
assign w41964 = w22727 & ~w22743;
assign w41965 = ~w22512 & w22746;
assign w41966 = w22512 & w22748;
assign w41967 = ~w22207 & ~w22204;
assign w41968 = w22498 & w22486;
assign w41969 = (w22791 & ~w22781) | (w22791 & w48186) | (~w22781 & w48186);
assign w41970 = ~w22829 & w48187;
assign w41971 = ~w22789 & w22602;
assign w41972 = w21970 & w22545;
assign w41973 = ~w22872 & w22545;
assign w41974 = w22498 & w22485;
assign w41975 = w22473 & w22446;
assign w41976 = w22366 & w48188;
assign w41977 = ~w22929 & w49303;
assign w41978 = ~w22929 & w49304;
assign w41979 = ~w22499 & w22991;
assign w41980 = ~w22997 & w22998;
assign w41981 = w22997 & w23000;
assign w41982 = ~w23021 & w22505;
assign w41983 = w23021 & ~w22505;
assign w41984 = ~w23021 & w23028;
assign w41985 = w23021 & w23030;
assign w41986 = w22767 & w48189;
assign w41987 = ~w22997 & w23043;
assign w41988 = w22997 & w23045;
assign w41989 = w23050 & w5745;
assign w41990 = (~w5745 & w22829) | (~w5745 & w9992) | (w22829 & w9992);
assign w41991 = ~w22207 & w48190;
assign w41992 = (w22291 & w22207) | (w22291 & w48191) | (w22207 & w48191);
assign w41993 = ~w22207 & w43564;
assign w41994 = (w23077 & w22207) | (w23077 & w43565) | (w22207 & w43565);
assign w41995 = ~w21955 & w48192;
assign w41996 = ~w22764 & w23100;
assign w41997 = (w22228 & w22204) | (w22228 & w48193) | (w22204 & w48193);
assign w41998 = ~w22204 & w48194;
assign w41999 = w23163 & w23167;
assign w42000 = (w23169 & w22207) | (w23169 & w48195) | (w22207 & w48195);
assign w42001 = (~w23166 & w22207) | (~w23166 & w43566) | (w22207 & w43566);
assign w42002 = ~w22207 & w43567;
assign w42003 = ~w22204 & w46591;
assign w42004 = (w23219 & w22204) | (w23219 & w46592) | (w22204 & w46592);
assign w42005 = w22767 & w43568;
assign w42006 = (~w23265 & w22204) | (~w23265 & w43569) | (w22204 & w43569);
assign w42007 = (w22766 & w46593) | (w22766 & w46594) | (w46593 & w46594);
assign w42008 = (~w11870 & ~w22767) | (~w11870 & w43570) | (~w22767 & w43570);
assign w42009 = w12666 & ~w23266;
assign w42010 = ~w22204 & w46595;
assign w42011 = (~w23304 & w22204) | (~w23304 & w46596) | (w22204 & w46596);
assign w42012 = (w23316 & w22204) | (w23316 & w46597) | (w22204 & w46597);
assign w42013 = ~w22204 & w46598;
assign w42014 = ~w23348 & w23368;
assign w42015 = (w23051 & ~w23338) | (w23051 & w48196) | (~w23338 & w48196);
assign w42016 = ~w21955 & w43571;
assign w42017 = ~w22477 & ~w23375;
assign w42018 = ~w22761 & w22742;
assign w42019 = ~w22206 & w43572;
assign w42020 = ~w22705 & w52314;
assign w42021 = w22477 & w22762;
assign w42022 = (~w22705 & w22204) | (~w22705 & w49305) | (w22204 & w49305);
assign w42023 = w23450 & w23404;
assign w42024 = ~w4838 & w5330;
assign w42025 = ~w23498 & ~w23499;
assign w42026 = (w22137 & w22730) | (w22137 & w46599) | (w22730 & w46599);
assign w42027 = ~w22764 & ~w22118;
assign w42028 = ~w23532 & w22175;
assign w42029 = ~w23532 & w23536;
assign w42030 = ~w23532 & w22183;
assign w42031 = (w43573 & w22203) | (w43573 & w48197) | (w22203 & w48197);
assign w42032 = (w43574 & w22203) | (w43574 & w48198) | (w22203 & w48198);
assign w42033 = (w23556 & w43575) | (w23556 & w22204) | (w43575 & w22204);
assign w42034 = (w23556 & w43576) | (w23556 & w22204) | (w43576 & w22204);
assign w42035 = (w43577 & w22203) | (w43577 & w48199) | (w22203 & w48199);
assign w42036 = (w43578 & w22203) | (w43578 & w48200) | (w22203 & w48200);
assign w42037 = (w23570 & w43579) | (w23570 & w22204) | (w43579 & w22204);
assign w42038 = (w23570 & w43580) | (w23570 & w22204) | (w43580 & w22204);
assign w42039 = ~w23621 & w23637;
assign w42040 = ~w23504 & w23593;
assign w42041 = ~w23532 & w23685;
assign w42042 = ~w23504 & w23752;
assign w42043 = w23504 & w23759;
assign w42044 = ~w23835 & ~w23834;
assign w42045 = ~w23504 & w23837;
assign w42046 = ~w23851 & w23853;
assign w42047 = (~w14766 & w23204) | (~w14766 & w43581) | (w23204 & w43581);
assign w42048 = ~w23504 & w23849;
assign w42049 = ~w23348 & w24264;
assign w42050 = (~w24267 & w24265) | (~w24267 & w43582) | (w24265 & w43582);
assign w42051 = ~w23504 & w23530;
assign w42052 = ~w24606 & ~w23543;
assign w42053 = ~w24609 & w24615;
assign w42054 = ~w23842 & w24613;
assign w42055 = w23806 & w1120;
assign w42056 = w23806 & ~w945;
assign w42057 = ~w23842 & w23588;
assign w42058 = w23842 & ~w24628;
assign w42059 = ~w23630 & w24682;
assign w42060 = (~w24678 & ~w24688) | (~w24678 & w48201) | (~w24688 & w48201);
assign w42061 = w24688 & w24736;
assign w42062 = ~w24633 & w24697;
assign w42063 = ~w23845 & ~w23768;
assign w42064 = w23741 & ~w23768;
assign w42065 = w23806 & w252;
assign w42066 = ~w24728 & w24725;
assign w42067 = w24728 & ~w24725;
assign w42068 = ~w23842 & w23729;
assign w42069 = w24732 & ~w252;
assign w42070 = ~w24764 & ~w24748;
assign w42071 = ~w24732 & w252;
assign w42072 = ~w24785 & ~w23863;
assign w42073 = ~w23763 & w23745;
assign w42074 = ~w23842 & ~w80;
assign w42075 = ~w23856 & ~w23682;
assign w42076 = w24822 & w24827;
assign w42077 = ~w24822 & w24829;
assign w42078 = w23802 & ~w23821;
assign w42079 = ~w24794 & w23665;
assign w42080 = ~w24794 & ~w23665;
assign w42081 = w24794 & ~w23665;
assign w42082 = w24794 & w23665;
assign w42083 = w24822 & w24853;
assign w42084 = ~w24822 & w24855;
assign w42085 = ~w24833 & ~w24859;
assign w42086 = w24865 & w24016;
assign w42087 = ~w24865 & w24891;
assign w42088 = ~w24902 & w24903;
assign w42089 = w24865 & ~w24907;
assign w42090 = ~w24038 & w24909;
assign w42091 = (w24787 & w46600) | (w24787 & w46601) | (w46600 & w46601);
assign w42092 = ~w24918 & w24920;
assign w42093 = (w10419 & ~w24914) | (w10419 & w46602) | (~w24914 & w46602);
assign w42094 = ~w24931 & w23997;
assign w42095 = ~w24865 & w24939;
assign w42096 = (w11870 & ~w24939) | (w11870 & w43583) | (~w24939 & w43583);
assign w42097 = ~w24931 & ~w23996;
assign w42098 = ~w24865 & w24951;
assign w42099 = ~w24871 & ~w23995;
assign w42100 = w24871 & w24960;
assign w42101 = (~w12666 & w24873) | (~w12666 & w46603) | (w24873 & w46603);
assign w42102 = (w7315 & w24862) | (w7315 & w46604) | (w24862 & w46604);
assign w42103 = w24871 & w24984;
assign w42104 = w24990 & w24539;
assign w42105 = ~w24990 & w24979;
assign w42106 = w24038 & w23976;
assign w42107 = ~w25001 & w24025;
assign w42108 = w25001 & ~w24025;
assign w42109 = (w24556 & w24862) | (w24556 & w46605) | (w24862 & w46605);
assign w42110 = ~w25034 & ~w25035;
assign w42111 = ~w24871 & ~w23960;
assign w42112 = w24865 & w23941;
assign w42113 = (~w9781 & w25041) | (~w9781 & w43584) | (w25041 & w43584);
assign w42114 = ~w25041 & w43585;
assign w42115 = w25065 & ~w6769;
assign w42116 = ~w25065 & w25068;
assign w42117 = w25071 & w24516;
assign w42118 = ~w25071 & ~w24516;
assign w42119 = ~w24865 & w25089;
assign w42120 = ~w25088 & ~w25091;
assign w42121 = (w24158 & w24865) | (w24158 & w46606) | (w24865 & w46606);
assign w42122 = ~w24865 & w46607;
assign w42123 = ~w25150 & ~w25149;
assign w42124 = ~w24865 & w25182;
assign w42125 = ~w25189 & ~w25188;
assign w42126 = (~w25204 & w24871) | (~w25204 & w46608) | (w24871 & w46608);
assign w42127 = w25202 & w25207;
assign w42128 = w24868 & w46609;
assign w42129 = (~w20000 & ~w24868) | (~w20000 & w46610) | (~w24868 & w46610);
assign w42130 = (~w25299 & w24871) | (~w25299 & w46611) | (w24871 & w46611);
assign w42131 = ~w24865 & w25304;
assign w42132 = (w43586 & w24873) | (w43586 & w46612) | (w24873 & w46612);
assign w42133 = ~w25311 & w25315;
assign w42134 = ~w25339 & w25341;
assign w42135 = ~w24871 & ~w2558;
assign w42136 = ~w24356 & w52315;
assign w42137 = w24865 & ~w24342;
assign w42138 = ~w25349 & w43587;
assign w42139 = (~w24288 & ~w25341) | (~w24288 & w43588) | (~w25341 & w43588);
assign w42140 = w24871 & ~w24326;
assign w42141 = (w25387 & ~w25386) | (w25387 & w48202) | (~w25386 & w48202);
assign w42142 = ~w25385 & ~w24298;
assign w42143 = ~w24871 & ~w24586;
assign w42144 = (~w24585 & ~w25386) | (~w24585 & w43589) | (~w25386 & w43589);
assign w42145 = ~w25392 & w46613;
assign w42146 = ~w24862 & w48203;
assign w42147 = (w24873 & w43590) | (w24873 & w43591) | (w43590 & w43591);
assign w42148 = (~w24873 & w43592) | (~w24873 & w43593) | (w43592 & w43593);
assign w42149 = ~w24862 & w48204;
assign w42150 = (~w24873 & w43594) | (~w24873 & w43595) | (w43594 & w43595);
assign w42151 = (w24873 & w43596) | (w24873 & w43597) | (w43596 & w43597);
assign w42152 = (~w24873 & w43598) | (~w24873 & w43599) | (w43598 & w43599);
assign w42153 = (w24873 & w43600) | (w24873 & w43601) | (w43600 & w43601);
assign w42154 = ~w24867 & w25439;
assign w42155 = ~w25458 & w25461;
assign w42156 = ~w25460 & ~w25463;
assign w42157 = w24865 & w25469;
assign w42158 = w25471 & w4838;
assign w42159 = ~w25475 & ~w24563;
assign w42160 = ~w25481 & ~w25480;
assign w42161 = w24865 & w25486;
assign w42162 = ~w25492 & w46614;
assign w42163 = ~w25457 & ~w25494;
assign w42164 = w25458 & ~w24562;
assign w42165 = w25497 & ~w5330;
assign w42166 = ~w24034 & w25501;
assign w42167 = (~w25502 & w24022) | (~w25502 & w46615) | (w24022 & w46615);
assign w42168 = w24871 & w25504;
assign w42169 = (w24787 & w46616) | (w24787 & w46617) | (w46616 & w46617);
assign w42170 = ~w25507 & w25508;
assign w42171 = (w25512 & w25507) | (w25512 & w48205) | (w25507 & w48205);
assign w42172 = ~w25492 & w46618;
assign w42173 = ~w4838 & ~w25471;
assign w42174 = ~w24871 & ~w24355;
assign w42175 = ~w24573 & w25533;
assign w42176 = w24865 & w24355;
assign w42177 = ~w25530 & w46619;
assign w42178 = ~w24573 & ~w24387;
assign w42179 = ~w24573 & w3646;
assign w42180 = ~w25552 & w25553;
assign w42181 = w24865 & ~w25557;
assign w42182 = (w25559 & ~w24573) | (w25559 & w46620) | (~w24573 & w46620);
assign w42183 = w24865 & ~w4838;
assign w42184 = (w24873 & w43602) | (w24873 & w43603) | (w43602 & w43603);
assign w42185 = w25571 & ~w25567;
assign w42186 = w25577 & ~w25582;
assign w42187 = ~w25577 & w25582;
assign w42188 = w24865 & w24417;
assign w42189 = ~w3646 & ~w25586;
assign w42190 = ~w25592 & ~w25591;
assign w42191 = ~w25595 & w25593;
assign w42192 = w24865 & w24423;
assign w42193 = (w24873 & w46621) | (w24873 & w46622) | (w46621 & w46622);
assign w42194 = ~w25552 & ~w24386;
assign w42195 = w25552 & w24386;
assign w42196 = w24865 & w3242;
assign w42197 = w25623 & w52316;
assign w42198 = (w24873 & w43604) | (w24873 & w43605) | (w43604 & w43605);
assign w42199 = (~w2285 & w25349) | (~w2285 & w46623) | (w25349 & w46623);
assign w42200 = w24868 & w48206;
assign w42201 = (w80 & w24862) | (w80 & w48207) | (w24862 & w48207);
assign w42202 = ~w25660 & w25662;
assign w42203 = ~w24871 & ~w57;
assign w42204 = ~w24865 & ~w25661;
assign w42205 = ~w25660 & ~w24734;
assign w42206 = w24865 & ~w24747;
assign w42207 = w24865 & ~w252;
assign w42208 = w25686 & w52317;
assign w42209 = (w24873 & w43606) | (w24873 & w43607) | (w43606 & w43607);
assign w42210 = ~w25684 & ~w57;
assign w42211 = ~w25683 & w377;
assign w42212 = w24573 & w24895;
assign w42213 = ~w25711 & w24761;
assign w42214 = w24871 & ~w24667;
assign w42215 = w24555 & w25722;
assign w42216 = w24706 & w46624;
assign w42217 = w24871 & ~w25729;
assign w42218 = (w24632 & w24871) | (w24632 & w43608) | (w24871 & w43608);
assign w42219 = w25756 & ~w25754;
assign w42220 = w25756 & w25760;
assign w42221 = w25759 & ~w25764;
assign w42222 = ~w25511 & ~w24497;
assign w42223 = ~w25790 & w5745;
assign w42224 = w25616 & ~w25798;
assign w42225 = w25311 & w25326;
assign w42226 = ~w25616 & ~w25631;
assign w42227 = (w25313 & w25264) | (w25313 & w43609) | (w25264 & w43609);
assign w42228 = (~w25589 & w25852) | (~w25589 & w25613) | (w25852 & w25613);
assign w42229 = (~w25312 & w25264) | (~w25312 & w43610) | (w25264 & w43610);
assign w42230 = w25616 & w26803;
assign w42231 = ~w26807 & w26803;
assign w42232 = w26051 & w26815;
assign w42233 = w26816 & w26818;
assign w42234 = ~w26816 & w26820;
assign w42235 = ~w26439 & w26826;
assign w42236 = w26816 & w26828;
assign w42237 = ~w26816 & w26830;
assign w42238 = ~w26822 & w26832;
assign w42239 = w25850 & w26845;
assign w42240 = w25850 & w25359;
assign w42241 = w26747 & ~w1120;
assign w42242 = w26738 & w26863;
assign w42243 = ~w26738 & w26865;
assign w42244 = ~w26752 & ~w26755;
assign w42245 = w26752 & w26755;
assign w42246 = ~w26070 & ~w26076;
assign w42247 = ~w26890 & ~w26894;
assign w42248 = w26003 & ~w26884;
assign w42249 = (w26065 & w26826) | (w26065 & w43611) | (w26826 & w43611);
assign w42250 = ~w26439 & w26942;
assign w42251 = w26437 & w46625;
assign w42252 = ~w26960 & w46626;
assign w42253 = w26077 & w26750;
assign w42254 = (~w1120 & w26893) | (~w1120 & w49828) | (w26893 & w49828);
assign w42255 = (w754 & w26960) | (w754 & w46627) | (w26960 & w46627);
assign w42256 = ~w26794 & w27027;
assign w42257 = w26794 & ~w26802;
assign w42258 = ~w26824 & ~w27054;
assign w42259 = ~w27072 & w27076;
assign w42260 = w27072 & w2285;
assign w42261 = (w27089 & w26287) | (w27089 & w43612) | (w26287 & w43612);
assign w42262 = (w26720 & w26287) | (w26720 & w43613) | (w26287 & w43613);
assign w42263 = ~w26893 & w46628;
assign w42264 = (w26718 & w26287) | (w26718 & w43614) | (w26287 & w43614);
assign w42265 = (w27143 & w26317) | (w27143 & w48208) | (w26317 & w48208);
assign w42266 = w26430 & ~w27144;
assign w42267 = w27150 & ~w27144;
assign w42268 = ~w26317 & w48209;
assign w42269 = (w27163 & w26287) | (w27163 & w48210) | (w26287 & w48210);
assign w42270 = w26318 & w27183;
assign w42271 = (~w27184 & w26287) | (~w27184 & w50141) | (w26287 & w50141);
assign w42272 = w26851 & w27021;
assign w42273 = w26978 & ~w27259;
assign w42274 = (~w27265 & w26074) | (~w27265 & w46629) | (w26074 & w46629);
assign w42275 = ~w26861 & w46630;
assign w42276 = ~w26893 & w46631;
assign w42277 = (~w27276 & w26894) | (~w27276 & w46632) | (w26894 & w46632);
assign w42278 = ~w26893 & w49829;
assign w42279 = ~w26075 & w26484;
assign w42280 = ~w26893 & w46633;
assign w42281 = (w27314 & w26074) | (w27314 & w46634) | (w26074 & w46634);
assign w42282 = (w27322 & w26074) | (w27322 & w46635) | (w26074 & w46635);
assign w42283 = ~w27310 & ~w23843;
assign w42284 = ~w26861 & w46636;
assign w42285 = (w27374 & w26074) | (w27374 & w46637) | (w26074 & w46637);
assign w42286 = ~w26565 & w27389;
assign w42287 = ~w26077 & ~w27392;
assign w42288 = ~w27392 & w26615;
assign w42289 = ~w26077 & ~w27403;
assign w42290 = (~w27447 & w26894) | (~w27447 & w46638) | (w26894 & w46638);
assign w42291 = ~w26565 & w26622;
assign w42292 = ~w26077 & w27474;
assign w42293 = ~w26698 & w43615;
assign w42294 = (w27488 & w26698) | (w27488 & w43616) | (w26698 & w43616);
assign w42295 = (w26282 & w26698) | (w26282 & w43617) | (w26698 & w43617);
assign w42296 = ~w27510 & ~w27509;
assign w42297 = w27524 & w27527;
assign w42298 = ~w27524 & w27529;
assign w42299 = ~w27541 & ~w14039;
assign w42300 = w27541 & w14039;
assign w42301 = ~w27547 & w27538;
assign w42302 = w27547 & w27551;
assign w42303 = ~w27547 & w27559;
assign w42304 = w27547 & w27566;
assign w42305 = w27524 & w27588;
assign w42306 = ~w27524 & w27590;
assign w42307 = ~w27604 & ~w27603;
assign w42308 = ~w27628 & w46639;
assign w42309 = (~w26127 & w27628) | (~w26127 & w46640) | (w27628 & w46640);
assign w42310 = w27641 & ~w27634;
assign w42311 = ~w26077 & ~w10419;
assign w42312 = ~w27677 & ~w27679;
assign w42313 = ~w26965 & w27685;
assign w42314 = ~w26087 & w26248;
assign w42315 = ~w26965 & w27727;
assign w42316 = w26158 & w27729;
assign w42317 = w26158 & w27733;
assign w42318 = (w10419 & ~w26880) | (w10419 & w43618) | (~w26880 & w43618);
assign w42319 = ~w27717 & w27748;
assign w42320 = ~w27717 & w27754;
assign w42321 = ~w27717 & w27765;
assign w42322 = w27717 & w27767;
assign w42323 = (~w27752 & w27778) | (~w27752 & w49830) | (w27778 & w49830);
assign w42324 = ~w27790 & ~w27789;
assign w42325 = ~w26077 & w6264;
assign w42326 = ~w26965 & w27827;
assign w42327 = ~w27832 & ~w27848;
assign w42328 = w26880 & w43619;
assign w42329 = ~w27762 & ~w27752;
assign w42330 = w27905 & ~w27260;
assign w42331 = ~w26889 & w27910;
assign w42332 = (w26882 & w48211) | (w26882 & w48212) | (w48211 & w48212);
assign w42333 = w27951 & ~w26884;
assign w42334 = ~w26074 & w49306;
assign w42335 = ~w27639 & ~w27651;
assign w42336 = ~w28037 & ~w28039;
assign w42337 = ~w28036 & w49307;
assign w42338 = (w28099 & w28049) | (w28099 & w43621) | (w28049 & w43621);
assign w42339 = (w43622 & w27260) | (w43622 & w50142) | (w27260 & w50142);
assign w42340 = w42337 & w46641;
assign w42341 = (w28183 & w28049) | (w28183 & w43623) | (w28049 & w43623);
assign w42342 = ~w28192 & w43624;
assign w42343 = ~w28050 & ~w28237;
assign w42344 = ~w28050 & w28244;
assign w42345 = w26978 & w27216;
assign w42346 = w28272 & ~w28251;
assign w42347 = ~w28049 & w43625;
assign w42348 = (w28275 & w28049) | (w28275 & w43626) | (w28049 & w43626);
assign w42349 = w28050 & w27515;
assign w42350 = (w11138 & w28324) | (w11138 & w43627) | (w28324 & w43627);
assign w42351 = ~w28050 & w28347;
assign w42352 = ~w28049 & w43628;
assign w42353 = ~w28409 & w46642;
assign w42354 = (~w14039 & w28421) | (~w14039 & w43629) | (w28421 & w43629);
assign w42355 = ~w28295 & ~w15681;
assign w42356 = w28295 & w15681;
assign w42357 = ~w28435 & w43630;
assign w42358 = (~w27616 & w28435) | (~w27616 & w43631) | (w28435 & w43631);
assign w42359 = ~w28421 & w50143;
assign w42360 = ~w28446 & w43632;
assign w42361 = ~w28455 & w46643;
assign w42362 = ~w28049 & w43633;
assign w42363 = ~w28050 & w28469;
assign w42364 = ~w28049 & w43634;
assign w42365 = ~w28050 & w28490;
assign w42366 = ~w27746 & ~w27874;
assign w42367 = (~w27260 & w50144) | (~w27260 & w50145) | (w50144 & w50145);
assign w42368 = (w28076 & w43638) | (w28076 & w43639) | (w43638 & w43639);
assign w42369 = (~w28076 & w43640) | (~w28076 & w43641) | (w43640 & w43641);
assign w42370 = (~w28076 & w43642) | (~w28076 & w43643) | (w43642 & w43643);
assign w42371 = (w28076 & w43644) | (w28076 & w43645) | (w43644 & w43645);
assign w42372 = w28050 & ~w5745;
assign w42373 = ~w28050 & w28548;
assign w42374 = ~w28564 & w28565;
assign w42375 = (w28507 & w28049) | (w28507 & w43646) | (w28049 & w43646);
assign w42376 = (w7315 & w28049) | (w7315 & w43647) | (w28049 & w43647);
assign w42377 = ~w28583 & ~w28584;
assign w42378 = (w43648 & w27260) | (w43648 & w50146) | (w27260 & w50146);
assign w42379 = ~w28564 & w28610;
assign w42380 = (w27216 & ~w27904) | (w27216 & w43649) | (~w27904 & w43649);
assign w42381 = ~w28050 & ~w28636;
assign w42382 = ~w28049 & w43650;
assign w42383 = (~w28076 & w43651) | (~w28076 & w43652) | (w43651 & w43652);
assign w42384 = ~w28049 & w43653;
assign w42385 = w28050 & ~w28711;
assign w42386 = ~w27907 & w46644;
assign w42387 = w42386 & w49831;
assign w42388 = ~w28719 & ~w28718;
assign w42389 = w27006 & w26994;
assign w42390 = (~w26975 & w28717) | (~w26975 & w48213) | (w28717 & w48213);
assign w42391 = ~w28049 & w43654;
assign w42392 = (w28076 & w43655) | (w28076 & w43656) | (w43655 & w43656);
assign w42393 = w28761 & ~w28755;
assign w42394 = (w28076 & w43657) | (w28076 & w43658) | (w43657 & w43658);
assign w42395 = w28050 & w26991;
assign w42396 = ~w28773 & w27248;
assign w42397 = ~w28777 & ~w28778;
assign w42398 = ~w27905 & w28783;
assign w42399 = w28050 & ~w28792;
assign w42400 = ~w28809 & ~w28810;
assign w42401 = ~w28815 & w46645;
assign w42402 = w28816 & w612;
assign w42403 = ~w28816 & ~w612;
assign w42404 = ~w28859 & ~w28858;
assign w42405 = ~w28050 & w28862;
assign w42406 = (w28689 & w43660) | (w28689 & w43661) | (w43660 & w43661);
assign w42407 = (~w27260 & w50147) | (~w27260 & w50148) | (w50147 & w50148);
assign w42408 = ~w28077 & w43663;
assign w42409 = (w28880 & w28077) | (w28880 & w43664) | (w28077 & w43664);
assign w42410 = ~w28076 & w50149;
assign w42411 = ~w28923 & w28922;
assign w42412 = ~w28770 & ~w28936;
assign w42413 = (w28943 & w28049) | (w28943 & w43665) | (w28049 & w43665);
assign w42414 = ~w28049 & w43666;
assign w42415 = (w1541 & w28049) | (w1541 & w43667) | (w28049 & w43667);
assign w42416 = ~w28049 & w43668;
assign w42417 = (w28076 & w43669) | (w28076 & w43670) | (w43669 & w43670);
assign w42418 = ~w29041 & w29043;
assign w42419 = w28050 & w27158;
assign w42420 = (w29053 & w48214) | (w29053 & w48215) | (w48214 & w48215);
assign w42421 = w28077 & w46646;
assign w42422 = (w2558 & ~w28077) | (w2558 & w43672) | (~w28077 & w43672);
assign w42423 = (~w29078 & w28049) | (~w29078 & w43673) | (w28049 & w43673);
assign w42424 = ~w29079 & w43674;
assign w42425 = ~w28050 & ~w29039;
assign w42426 = (~w29092 & w28049) | (~w29092 & w43675) | (w28049 & w43675);
assign w42427 = w29092 & w52318;
assign w42428 = w29099 & w4056;
assign w42429 = ~w29108 & ~w29109;
assign w42430 = (w28076 & w43677) | (w28076 & w43678) | (w43677 & w43678);
assign w42431 = (~w28076 & w43679) | (~w28076 & w43680) | (w43679 & w43680);
assign w42432 = (~w28076 & w43681) | (~w28076 & w43682) | (w43681 & w43682);
assign w42433 = (w28076 & w43683) | (w28076 & w43684) | (w43683 & w43684);
assign w42434 = (w2896 & w29079) | (w2896 & w46647) | (w29079 & w46647);
assign w42435 = w28930 & ~w29208;
assign w42436 = w29157 & w43685;
assign w42437 = w28919 & w43686;
assign w42438 = w29157 & w43687;
assign w42439 = (w29645 & ~w29157) | (w29645 & w43688) | (~w29157 & w43688);
assign w42440 = ~w28938 & w945;
assign w42441 = w28919 & w46648;
assign w42442 = ~w28770 & w28882;
assign w42443 = ~w28936 & w46649;
assign w42444 = (w30058 & w28936) | (w30058 & w46650) | (w28936 & w46650);
assign w42445 = w28681 & w30073;
assign w42446 = ~w29157 & w252;
assign w42447 = w29157 & w28743;
assign w42448 = w28738 & w30107;
assign w42449 = ~w42 & ~w30043;
assign w42450 = w30120 & w30122;
assign w42451 = ~w29722 & w30151;
assign w42452 = w29722 & w30153;
assign w42453 = ~w29722 & w30162;
assign w42454 = w29722 & w30164;
assign w42455 = w30161 & ~w4838;
assign w42456 = ~w29157 & ~w4838;
assign w42457 = w29157 & w29687;
assign w42458 = w28546 & w30189;
assign w42459 = ~w29113 & w3242;
assign w42460 = ~w29157 & ~w29132;
assign w42461 = ~w30236 & ~w30148;
assign w42462 = ~w30149 & ~w30238;
assign w42463 = w30032 & w29997;
assign w42464 = (w30241 & w43689) | (w30241 & w52319) | (w43689 & w52319);
assign w42465 = (w43690 & w30250) | (w43690 & w46651) | (w30250 & w46651);
assign w42466 = ~w30249 & w49308;
assign w42467 = (~w29977 & w30147) | (~w29977 & w46652) | (w30147 & w46652);
assign w42468 = w30273 & w30284;
assign w42469 = (w30289 & w30286) | (w30289 & w46653) | (w30286 & w46653);
assign w42470 = ~w30286 & w46654;
assign w42471 = (w30294 & w30238) | (w30294 & w46655) | (w30238 & w46655);
assign w42472 = (~w29926 & w30147) | (~w29926 & w46656) | (w30147 & w46656);
assign w42473 = ~w30307 & w30303;
assign w42474 = w30313 & w30315;
assign w42475 = (w30317 & w30286) | (w30317 & w46657) | (w30286 & w46657);
assign w42476 = ~w30286 & w46658;
assign w42477 = ~w30312 & w30322;
assign w42478 = ~w30273 & ~w30283;
assign w42479 = ~w30313 & w30333;
assign w42480 = w30313 & w30335;
assign w42481 = ~w30308 & w43691;
assign w42482 = ~w30361 & ~w30360;
assign w42483 = (w30030 & w30242) | (w30030 & w30035) | (w30242 & w30035);
assign w42484 = ~w29963 & w30446;
assign w42485 = (~w30525 & w30147) | (~w30525 & w46659) | (w30147 & w46659);
assign w42486 = (w28077 & ~w30148) | (w28077 & w46660) | (~w30148 & w46660);
assign w42487 = (w30547 & w30147) | (w30547 & w48216) | (w30147 & w48216);
assign w42488 = ~w30238 & w46661;
assign w42489 = ~w30564 & w46662;
assign w42490 = ~w30148 & ~w30596;
assign w42491 = w29474 & w24874;
assign w42492 = ~w29474 & ~w24874;
assign w42493 = ~w30606 & w30609;
assign w42494 = w30606 & w30612;
assign w42495 = ~w30145 & w30628;
assign w42496 = ~w30236 & w30629;
assign w42497 = ~w30148 & ~w30648;
assign w42498 = w30629 & w30658;
assign w42499 = ~w30237 & w46663;
assign w42500 = (~w29484 & w30237) | (~w29484 & w46664) | (w30237 & w46664);
assign w42501 = (~w29489 & w29474) | (~w29489 & w43692) | (w29474 & w43692);
assign w42502 = ~w30669 & ~w30682;
assign w42503 = w29516 & ~w29264;
assign w42504 = ~w29516 & w29358;
assign w42505 = ~w29654 & w29338;
assign w42506 = ~w29277 & w30787;
assign w42507 = ~w29963 & w30237;
assign w42508 = ~w12666 & w30787;
assign w42509 = ~w30800 & w46665;
assign w42510 = (~w29336 & ~w30785) | (~w29336 & w43693) | (~w30785 & w43693);
assign w42511 = (w11870 & w30800) | (w11870 & w46666) | (w30800 & w46666);
assign w42512 = w29647 & ~w14766;
assign w42513 = ~w29647 & w14766;
assign w42514 = (w30785 & w46667) | (w30785 & w46668) | (w46667 & w46668);
assign w42515 = ~w30862 & w30865;
assign w42516 = ~w30145 & w29343;
assign w42517 = ~w29517 & w29266;
assign w42518 = w30238 & w46669;
assign w42519 = (w30836 & ~w30238) | (w30836 & w46670) | (~w30238 & w46670);
assign w42520 = ~w30800 & w48217;
assign w42521 = (w15681 & w30800) | (w15681 & w46671) | (w30800 & w46671);
assign w42522 = ~w29664 & w29633;
assign w42523 = ~w29664 & w30957;
assign w42524 = w29662 & w30987;
assign w42525 = w29662 & w29617;
assign w42526 = ~w30148 & w31002;
assign w42527 = w30148 & w31005;
assign w42528 = w31011 & ~w31012;
assign w42529 = ~w31011 & w31015;
assign w42530 = ~w31023 & w31029;
assign w42531 = ~w30942 & ~w31048;
assign w42532 = ~w30148 & w31050;
assign w42533 = w30148 & w31053;
assign w42534 = ~w31029 & w31023;
assign w42535 = ~w29546 & ~w31069;
assign w42536 = ~w31076 & w31079;
assign w42537 = ~w31083 & ~w31082;
assign w42538 = ~w29546 & w31089;
assign w42539 = w30239 & w46672;
assign w42540 = ~w29546 & ~w31107;
assign w42541 = w31116 & w30239;
assign w42542 = w31118 & ~w30239;
assign w42543 = ~w29546 & ~w30174;
assign w42544 = w31137 & w30239;
assign w42545 = w31139 & ~w30239;
assign w42546 = w29546 & ~w31146;
assign w42547 = ~w30238 & w46673;
assign w42548 = (~w5330 & w30238) | (~w5330 & w46674) | (w30238 & w46674);
assign w42549 = (~w5745 & w30238) | (~w5745 & w46675) | (w30238 & w46675);
assign w42550 = ~w29593 & ~w29537;
assign w42551 = w31167 & w5330;
assign w42552 = w31195 & w30239;
assign w42553 = w31197 & ~w30239;
assign w42554 = (w4056 & ~w30239) | (w4056 & w46676) | (~w30239 & w46676);
assign w42555 = w31206 & w30239;
assign w42556 = w31208 & ~w30239;
assign w42557 = w30246 & w46677;
assign w42558 = ~w30308 & w43694;
assign w42559 = ~w31248 & w31251;
assign w42560 = (~w31250 & w30147) | (~w31250 & w46678) | (w30147 & w46678);
assign w42561 = (w31271 & w30238) | (w31271 & w46679) | (w30238 & w46679);
assign w42562 = ~w31248 & w31274;
assign w42563 = ~w30238 & w46680;
assign w42564 = ~w31248 & w31280;
assign w42565 = ~w30238 & w46681;
assign w42566 = (w31285 & w30238) | (w31285 & w46682) | (w30238 & w46682);
assign w42567 = ~w29675 & ~w30216;
assign w42568 = (w31298 & w31289) | (w31298 & w46683) | (w31289 & w46683);
assign w42569 = ~w30238 & w46684;
assign w42570 = (w31304 & w30238) | (w31304 & w46685) | (w30238 & w46685);
assign w42571 = (w31310 & w30238) | (w31310 & w46686) | (w30238 & w46686);
assign w42572 = ~w30238 & w46687;
assign w42573 = w31322 & ~w3242;
assign w42574 = ~w31322 & ~w31325;
assign w42575 = ~w30148 & ~w31337;
assign w42576 = ~w31076 & w31342;
assign w42577 = w31345 & ~w31349;
assign w42578 = ~w31322 & ~w31246;
assign w42579 = ~w31247 & w46688;
assign w42580 = ~w31416 & w30516;
assign w42581 = ~w31430 & w31435;
assign w42582 = ~w31437 & ~w31429;
assign w42583 = w31213 & w31428;
assign w42584 = w30779 & w31448;
assign w42585 = ~w31465 & w31468;
assign w42586 = w31367 & ~w30468;
assign w42587 = ~w31475 & ~w31421;
assign w42588 = w31416 & ~w1320;
assign w42589 = ~w31464 & w43695;
assign w42590 = ~w31464 & w43696;
assign w42591 = w31446 & ~w31455;
assign w42592 = ~w31464 & w43697;
assign w42593 = (w31534 & w31421) | (w31534 & w43698) | (w31421 & w43698);
assign w42594 = (w31580 & w31421) | (w31580 & w43699) | (w31421 & w43699);
assign w42595 = ~w31421 & w43700;
assign w42596 = w31421 & w46689;
assign w42597 = (~w30877 & ~w31421) | (~w30877 & w43701) | (~w31421 & w43701);
assign w42598 = w31421 & w43702;
assign w42599 = (w31671 & ~w31421) | (w31671 & w43703) | (~w31421 & w43703);
assign w42600 = ~w30683 & ~w30730;
assign w42601 = w31421 & w43704;
assign w42602 = (w31692 & ~w31421) | (w31692 & w43705) | (~w31421 & w43705);
assign w42603 = w31421 & w43706;
assign w42604 = (w31700 & ~w31421) | (w31700 & w43707) | (~w31421 & w43707);
assign w42605 = (~w31762 & w31421) | (~w31762 & ~w31761) | (w31421 & ~w31761);
assign w42606 = (~w31773 & w31421) | (~w31773 & w46690) | (w31421 & w46690);
assign w42607 = (~w31785 & w31421) | (~w31785 & w43708) | (w31421 & w43708);
assign w42608 = (~w31794 & w31421) | (~w31794 & w46691) | (w31421 & w46691);
assign w42609 = ~w31464 & w43709;
assign w42610 = (~w31819 & w31421) | (~w31819 & w43710) | (w31421 & w43710);
assign w42611 = (w31824 & w31421) | (w31824 & w46692) | (w31421 & w46692);
assign w42612 = w31367 & w31839;
assign w42613 = w31494 & w31846;
assign w42614 = (w31852 & ~w31421) | (w31852 & w43711) | (~w31421 & w43711);
assign w42615 = (~w31873 & w31421) | (~w31873 & w43712) | (w31421 & w43712);
assign w42616 = (~w31877 & w31421) | (~w31877 & w46693) | (w31421 & w46693);
assign w42617 = ~w31901 & ~w31902;
assign w42618 = ~w31955 & w31954;
assign w42619 = (~w31967 & w31421) | (~w31967 & w43713) | (w31421 & w43713);
assign w42620 = ~w31978 & w31977;
assign w42621 = w31367 & w31997;
assign w42622 = w31421 & w43714;
assign w42623 = (w32004 & ~w31421) | (w32004 & w43715) | (~w31421 & w43715);
assign w42624 = w31421 & w43716;
assign w42625 = (w30588 & ~w31421) | (w30588 & w43717) | (~w31421 & w43717);
assign w42626 = ~w32079 & ~w32080;
assign w42627 = ~w32074 & w43718;
assign w42628 = (~w4838 & w31421) | (~w4838 & w43719) | (w31421 & w43719);
assign w42629 = ~w32269 & ~w32268;
assign w42630 = w32284 & ~w32285;
assign w42631 = ~w32330 & ~w32331;
assign w42632 = w31367 & w32434;
assign w42633 = w31367 & w32446;
assign w42634 = ~w32456 & w30508;
assign w42635 = w31477 & w43720;
assign w42636 = (~w32445 & ~w31477) | (~w32445 & w43721) | (~w31477 & w43721);
assign w42637 = w31367 & w32466;
assign w42638 = w31421 & w43722;
assign w42639 = w31421 & w43723;
assign w42640 = (~w30507 & w32455) | (~w30507 & w43724) | (w32455 & w43724);
assign w42641 = w32576 & ~w32581;
assign w42642 = w32379 & ~w32697;
assign w42643 = (~w32721 & w32697) | (~w32721 & w43725) | (w32697 & w43725);
assign w42644 = ~w32428 & w32724;
assign w42645 = (~w32579 & w32697) | (~w32579 & w43726) | (w32697 & w43726);
assign w42646 = w32711 & w46694;
assign w42647 = ~w32428 & w32574;
assign w42648 = ~w32428 & w32760;
assign w42649 = (w32444 & w32697) | (w32444 & w43727) | (w32697 & w43727);
assign w42650 = ~w32697 & w43728;
assign w42651 = (w32444 & w32697) | (w32444 & w46695) | (w32697 & w46695);
assign w42652 = ~w32697 & w43729;
assign w42653 = (w32554 & w32235) | (w32554 & w43730) | (w32235 & w43730);
assign w42654 = ~w32698 & w43731;
assign w42655 = (w32828 & w32698) | (w32828 & w43732) | (w32698 & w43732);
assign w42656 = ~w32698 & w43733;
assign w42657 = (w32852 & w32698) | (w32852 & w43734) | (w32698 & w43734);
assign w42658 = ~w32259 & w43735;
assign w42659 = (~w32236 & w32419) | (~w32236 & w43736) | (w32419 & w43736);
assign w42660 = (~w32825 & w32698) | (~w32825 & w43737) | (w32698 & w43737);
assign w42661 = ~w32698 & w43738;
assign w42662 = (w31971 & w32697) | (w31971 & w46696) | (w32697 & w46696);
assign w42663 = ~w32697 & w43739;
assign w42664 = (w33020 & w32697) | (w33020 & w43740) | (w32697 & w43740);
assign w42665 = ~w32697 & w43741;
assign w42666 = (w33030 & w32697) | (w33030 & w43742) | (w32697 & w43742);
assign w42667 = ~w32697 & w43743;
assign w42668 = (w33072 & w32697) | (w33072 & w43744) | (w32697 & w43744);
assign w42669 = ~w32697 & w43745;
assign w42670 = (~w31668 & w32697) | (~w31668 & w46697) | (w32697 & w46697);
assign w42671 = w33519 & ~w9195;
assign w42672 = (~w33632 & w32697) | (~w33632 & w43746) | (w32697 & w43746);
assign w42673 = ~w33519 & w9195;
assign w42674 = (~w6264 & w32698) | (~w6264 & w46698) | (w32698 & w46698);
assign w42675 = w33677 & w33679;
assign w42676 = w5330 & ~w33689;
assign w42677 = w32129 & w4430;
assign w42678 = w33591 & w33707;
assign w42679 = ~w33591 & w33709;
assign w42680 = ~w32997 & w46699;
assign w42681 = w33631 & w32968;
assign w42682 = w33737 & ~w33741;
assign w42683 = w33744 & ~w33735;
assign w42684 = ~w33696 & w33728;
assign w42685 = (~w32717 & w32997) | (~w32717 & w43747) | (w32997 & w43747);
assign w42686 = (w33788 & w33736) | (w33788 & w43748) | (w33736 & w43748);
assign w42687 = (w32872 & w33736) | (w32872 & w43749) | (w33736 & w43749);
assign w42688 = ~w32998 & w33812;
assign w42689 = (w33861 & w32997) | (w33861 & w43750) | (w32997 & w43750);
assign w42690 = ~w32997 & w43751;
assign w42691 = (~w33872 & w32997) | (~w33872 & w43753) | (w32997 & w43753);
assign w42692 = ~w32997 & w46700;
assign w42693 = (w33879 & w32997) | (w33879 & w43754) | (w32997 & w43754);
assign w42694 = ~w32997 & w43755;
assign w42695 = ~w32997 & w43756;
assign w42696 = ~w32997 & w43757;
assign w42697 = (~w33896 & w32997) | (~w33896 & w43758) | (w32997 & w43758);
assign w42698 = ~w33729 & ~w32997;
assign w42699 = (w33911 & w32997) | (w33911 & w43759) | (w32997 & w43759);
assign w42700 = ~w32997 & w43760;
assign w42701 = (w33878 & w32997) | (w33878 & w43761) | (w32997 & w43761);
assign w42702 = ~w32997 & w43762;
assign w42703 = (~w33931 & w32997) | (~w33931 & w43763) | (w32997 & w43763);
assign w42704 = (~w33937 & w32789) | (~w33937 & w46701) | (w32789 & w46701);
assign w42705 = ~w32789 & w46702;
assign w42706 = ~w32789 & w46703;
assign w42707 = (~w33080 & w32789) | (~w33080 & w46704) | (w32789 & w46704);
assign w42708 = w33936 & ~w33935;
assign w42709 = w32790 & w33972;
assign w42710 = (w33098 & w32789) | (w33098 & w46705) | (w32789 & w46705);
assign w42711 = ~w32997 & w46706;
assign w42712 = (w33987 & w32997) | (w33987 & w46707) | (w32997 & w46707);
assign w42713 = ~w33100 & ~w33144;
assign w42714 = (w34000 & w32789) | (w34000 & w46708) | (w32789 & w46708);
assign w42715 = ~w34005 & ~w34004;
assign w42716 = ~w32998 & w34010;
assign w42717 = w32790 & ~w34016;
assign w42718 = w32790 & w34019;
assign w42719 = (~w32997 & w48218) | (~w32997 & w48219) | (w48218 & w48219);
assign w42720 = w33109 & w52320;
assign w42721 = w32790 & w34031;
assign w42722 = (w32997 & w48220) | (w32997 & w48221) | (w48220 & w48221);
assign w42723 = (~w32997 & w48222) | (~w32997 & w48223) | (w48222 & w48223);
assign w42724 = ~w34055 & ~w34056;
assign w42725 = ~w33177 & w19040;
assign w42726 = ~w32789 & w46709;
assign w42727 = ~w32789 & w46710;
assign w42728 = (w32997 & w48224) | (w32997 & w48225) | (w48224 & w48225);
assign w42729 = (~w32997 & w48226) | (~w32997 & w48227) | (w48226 & w48227);
assign w42730 = ~w34006 & ~w34011;
assign w42731 = (w32997 & w48228) | (w32997 & w48229) | (w48228 & w48229);
assign w42732 = w34123 & w52320;
assign w42733 = ~w32997 & w46711;
assign w42734 = (w34128 & w32997) | (w34128 & w46712) | (w32997 & w46712);
assign w42735 = ~w32997 & w46713;
assign w42736 = ~w32998 & w34146;
assign w42737 = ~w32997 & w46714;
assign w42738 = ~w32998 & w34155;
assign w42739 = ~w33247 & w34170;
assign w42740 = w32998 & w34176;
assign w42741 = w32998 & w34183;
assign w42742 = ~w34200 & ~w11870;
assign w42743 = w33306 & w14766;
assign w42744 = ~w33306 & ~w14766;
assign w42745 = (w34209 & w34208) | (w34209 & w43764) | (w34208 & w43764);
assign w42746 = ~w32998 & w33335;
assign w42747 = ~w33731 & w43765;
assign w42748 = (~w34202 & w33731) | (~w34202 & w43766) | (w33731 & w43766);
assign w42749 = ~w34208 & w46715;
assign w42750 = ~w34229 & ~w34233;
assign w42751 = w33306 & w33459;
assign w42752 = ~w33731 & w43767;
assign w42753 = (w34252 & w33731) | (w34252 & w43768) | (w33731 & w43768);
assign w42754 = w32998 & w33274;
assign w42755 = ~w34264 & ~w14766;
assign w42756 = ~w32998 & w34269;
assign w42757 = ~w32998 & w34272;
assign w42758 = w34264 & w14766;
assign w42759 = ~w34288 & ~w34289;
assign w42760 = w32998 & w34294;
assign w42761 = w32998 & w34181;
assign w42762 = ~w34180 & ~w34267;
assign w42763 = (w34584 & ~w34217) | (w34584 & w46716) | (~w34217 & w46716);
assign w42764 = (~w33450 & w33656) | (~w33450 & w46717) | (w33656 & w46717);
assign w42765 = w34320 & w52321;
assign w42766 = (w33555 & w46718) | (w33555 & w46719) | (w46718 & w46719);
assign w42767 = ~w32997 & w46720;
assign w42768 = ~w33555 & w46721;
assign w42769 = (~w34331 & w33555) | (~w34331 & w46722) | (w33555 & w46722);
assign w42770 = w32998 & w34338;
assign w42771 = w33552 & w33471;
assign w42772 = ~w34352 & ~w34349;
assign w42773 = (~w33659 & w34353) | (~w33659 & w46723) | (w34353 & w46723);
assign w42774 = w32998 & ~w34348;
assign w42775 = ~w32997 & w46724;
assign w42776 = (w33555 & w33451) | (w33555 & w46725) | (w33451 & w46725);
assign w42777 = ~w34370 & ~w34371;
assign w42778 = ~w33428 & ~w5330;
assign w42779 = ~w32997 & w46726;
assign w42780 = ~w32997 & w46727;
assign w42781 = ~w32998 & w34354;
assign w42782 = ~w33669 & w33452;
assign w42783 = ~w34391 & ~w33676;
assign w42784 = ~w32997 & w46728;
assign w42785 = ~w34395 & w34398;
assign w42786 = w34395 & w34400;
assign w42787 = w34395 & w34410;
assign w42788 = ~w34395 & w34412;
assign w42789 = (~w34423 & ~w33695) | (~w34423 & w46729) | (~w33695 & w46729);
assign w42790 = ~w34428 & ~w34427;
assign w42791 = ~w32997 & w46730;
assign w42792 = w33453 & ~w33699;
assign w42793 = (w33702 & w33695) | (w33702 & w46731) | (w33695 & w46731);
assign w42794 = (w34444 & w32789) | (w34444 & w46732) | (w32789 & w46732);
assign w42795 = (~w34469 & ~w34463) | (~w34469 & w46733) | (~w34463 & w46733);
assign w42796 = w34463 & w46734;
assign w42797 = w32998 & ~w34474;
assign w42798 = ~w33507 & ~w33551;
assign w42799 = w34482 & w34489;
assign w42800 = ~w34482 & w34491;
assign w42801 = ~w34494 & ~w33536;
assign w42802 = w34494 & w34502;
assign w42803 = ~w32790 & ~w34512;
assign w42804 = ~w34494 & ~w33639;
assign w42805 = w34482 & w34485;
assign w42806 = ~w34482 & w34488;
assign w42807 = w32998 & w34524;
assign w42808 = ~w32997 & w46735;
assign w42809 = w34479 & w34535;
assign w42810 = ~w34540 & w34537;
assign w42811 = w34540 & ~w34537;
assign w42812 = ~w34480 & w46736;
assign w42813 = (~w9781 & w34480) | (~w9781 & w46737) | (w34480 & w46737);
assign w42814 = ~w32997 & w46738;
assign w42815 = ~w33405 & w34463;
assign w42816 = ~w32997 & w46739;
assign w42817 = w34379 & ~w34572;
assign w42818 = (w34593 & w33739) | (w34593 & w46740) | (w33739 & w46740);
assign w42819 = (w32807 & w32997) | (w32807 & w46741) | (w32997 & w46741);
assign w42820 = (~w34610 & w32997) | (~w34610 & w46742) | (w32997 & w46742);
assign w42821 = (w34610 & w32997) | (w34610 & w46743) | (w32997 & w46743);
assign w42822 = (w32842 & w32997) | (w32842 & w43770) | (w32997 & w43770);
assign w42823 = (w34642 & w33739) | (w34642 & w43771) | (w33739 & w43771);
assign w42824 = (w2896 & w32789) | (w2896 & w46744) | (w32789 & w46744);
assign w42825 = ~w34668 & ~w34669;
assign w42826 = (w34671 & ~w33695) | (w34671 & w46745) | (~w33695 & w46745);
assign w42827 = w34667 & w34676;
assign w42828 = ~w34667 & w34678;
assign w42829 = w33453 & w33705;
assign w42830 = w34668 & w33705;
assign w42831 = ~w34683 & ~w33590;
assign w42832 = w32790 & w34687;
assign w42833 = ~w32997 & w46746;
assign w42834 = w34692 & w34696;
assign w42835 = ~w34692 & w34698;
assign w42836 = ~w34683 & w34703;
assign w42837 = ~w34668 & ~w34705;
assign w42838 = ~w34706 & w34707;
assign w42839 = ~w32997 & w46747;
assign w42840 = w34712 & ~w2896;
assign w42841 = (w34717 & w32997) | (w34717 & w46748) | (w32997 & w46748);
assign w42842 = ~w32997 & w46749;
assign w42843 = ~w34712 & w2896;
assign w42844 = ~w33610 & w50232;
assign w42845 = (w33695 & w46750) | (w33695 & w46751) | (w46750 & w46751);
assign w42846 = w3646 & w52322;
assign w42847 = ~w34734 & w34736;
assign w42848 = w34734 & w34738;
assign w42849 = ~w32997 & w43772;
assign w42850 = w34747 & w34753;
assign w42851 = w34757 & ~w34746;
assign w42852 = ~w33723 & ~w34769;
assign w42853 = (~w1738 & ~w33731) | (~w1738 & w43773) | (~w33731 & w43773);
assign w42854 = ~w34692 & w34776;
assign w42855 = w34692 & w34778;
assign w42856 = ~w32997 & w43774;
assign w42857 = ~w33730 & w43775;
assign w42858 = w34786 & w34795;
assign w42859 = ~w32997 & w46752;
assign w42860 = ~w32996 & w33722;
assign w42861 = ~w32997 & w46753;
assign w42862 = w34786 & ~w32964;
assign w42863 = w33731 & w43776;
assign w42864 = w34813 & w46754;
assign w42865 = w34834 & w34839;
assign w42866 = ~w34734 & w34846;
assign w42867 = w34734 & w34848;
assign w42868 = ~w34833 & w34819;
assign w42869 = ~w34861 & ~w34860;
assign w42870 = ~w34536 & ~w34544;
assign w42871 = w34701 & w34628;
assign w42872 = w34589 & w34821;
assign w42873 = w34856 & w50233;
assign w42874 = (~w34895 & w34871) | (~w34895 & w48230) | (w34871 & w48230);
assign w42875 = w33855 & w34925;
assign w42876 = ~w33855 & w34939;
assign w42877 = w33855 & w34941;
assign w42878 = w33855 & w34949;
assign w42879 = ~w33855 & ~w33934;
assign w42880 = w33855 & w34938;
assign w42881 = (w33855 & w34964) | (w33855 & w43778) | (w34964 & w43778);
assign w42882 = (w34995 & w49309) | (w34995 & w49310) | (w49309 & w49310);
assign w42883 = (~w35002 & w34871) | (~w35002 & w48231) | (w34871 & w48231);
assign w42884 = (~a[9] & w33855) | (~a[9] & w49311) | (w33855 & w49311);
assign w42885 = w34871 & w35036;
assign w42886 = ~w34871 & w49312;
assign w42887 = ~w33855 & w33915;
assign w42888 = (w43780 & w34995) | (w43780 & w49313) | (w34995 & w49313);
assign w42889 = w33924 & w33992;
assign w42890 = ~w35168 & ~w35167;
assign w42891 = w33855 & ~w35180;
assign w42892 = (~w19040 & w35180) | (~w19040 & w43781) | (w35180 & w43781);
assign w42893 = (~w20906 & w34919) | (~w20906 & w49314) | (w34919 & w49314);
assign w42894 = w33855 & w35224;
assign w42895 = ~w33855 & ~w35144;
assign w42896 = w33855 & w35233;
assign w42897 = ~w33855 & w34149;
assign w42898 = (w16559 & w43782) | (w16559 & w34899) | (w43782 & w34899);
assign w42899 = ~w34919 & w49315;
assign w42900 = ~w33855 & w34097;
assign w42901 = w33855 & w35254;
assign w42902 = (w43783 & w34898) | (w43783 & w49316) | (w34898 & w49316);
assign w42903 = (~w34588 & w34316) | (~w34588 & w43784) | (w34316 & w43784);
assign w42904 = ~w34590 & ~w34881;
assign w42905 = ~w33855 & ~w7315;
assign w42906 = ~w35411 & w43785;
assign w42907 = ~w34314 & w43786;
assign w42908 = ~w35420 & w35423;
assign w42909 = ~w34314 & w43787;
assign w42910 = (w42908 & w46755) | (w42908 & w46756) | (w46755 & w46756);
assign w42911 = (~w35435 & w49832) | (~w35435 & w49833) | (w49832 & w49833);
assign w42912 = (~w42908 & w46757) | (~w42908 & w46758) | (w46757 & w46758);
assign w42913 = ~w35427 & ~w35433;
assign w42914 = w35454 & w43788;
assign w42915 = ~w34899 & w43789;
assign w42916 = ~w35464 & w35468;
assign w42917 = ~w35464 & w35441;
assign w42918 = ~w33855 & ~w34292;
assign w42919 = (~w9781 & w34899) | (~w9781 & w43790) | (w34899 & w43790);
assign w42920 = w33855 & ~w35494;
assign w42921 = ~w34899 & w43791;
assign w42922 = ~w34279 & w34311;
assign w42923 = ~w34220 & w34313;
assign w42924 = ~w33855 & ~w34248;
assign w42925 = ~w34899 & w43792;
assign w42926 = (w8666 & w34899) | (w8666 & w43793) | (w34899 & w43793);
assign w42927 = ~w33855 & ~w6769;
assign w42928 = ~w35331 & w43794;
assign w42929 = (w10419 & w34899) | (w10419 & w43795) | (w34899 & w43795);
assign w42930 = ~w33855 & w5745;
assign w42931 = (w35580 & w43796) | (w35580 & w34899) | (w43796 & w34899);
assign w42932 = (w43797 & w34898) | (w43797 & w49317) | (w34898 & w49317);
assign w42933 = (~w35641 & w46759) | (~w35641 & w50234) | (w46759 & w50234);
assign w42934 = (w43798 & w35582) | (w43798 & w49318) | (w35582 & w49318);
assign w42935 = (~w35693 & w34881) | (~w35693 & w43799) | (w34881 & w43799);
assign w42936 = w35699 & w34835;
assign w42937 = (~w34835 & w35694) | (~w34835 & w43800) | (w35694 & w43800);
assign w42938 = ~w35706 & ~w35707;
assign w42939 = ~w33855 & w35722;
assign w42940 = (~w35717 & w35716) | (~w35717 & w43801) | (w35716 & w43801);
assign w42941 = ~w35726 & ~w2285;
assign w42942 = ~w34900 & w43802;
assign w42943 = w33855 & ~w34833;
assign w42944 = ~w33855 & w1320;
assign w42945 = (w33850 & w34870) | (w33850 & w49319) | (w34870 & w49319);
assign w42946 = (~w33845 & w34870) | (~w33845 & w49320) | (w34870 & w49320);
assign w42947 = ~w33855 & w252;
assign w42948 = (w35850 & w43803) | (w35850 & w34899) | (w43803 & w34899);
assign w42949 = (w43804 & w34898) | (w43804 & w49321) | (w34898 & w49321);
assign w42950 = ~w34859 & w35863;
assign w42951 = ~w35867 & w35875;
assign w42952 = ~w35867 & w35879;
assign w42953 = ~w35877 & ~w35880;
assign w42954 = w33855 & w35882;
assign w42955 = ~w33855 & ~w34617;
assign w42956 = ~w33855 & w351;
assign w42957 = (w35903 & w43805) | (w35903 & w34899) | (w43805 & w34899);
assign w42958 = (w43806 & w34898) | (w43806 & w49322) | (w34898 & w49322);
assign w42959 = w33855 & ~w34650;
assign w42960 = w35924 & ~w35925;
assign w42961 = ~w35924 & w35925;
assign w42962 = ~w35872 & ~w400;
assign w42963 = w35872 & ~w400;
assign w42964 = ~w35898 & ~w35902;
assign w42965 = w35916 & w612;
assign w42966 = ~w35794 & ~w35961;
assign w42967 = w35409 & w35936;
assign w42968 = ~w35979 & ~w35978;
assign w42969 = w35804 & ~w35794;
assign w42970 = w35980 & ~w35998;
assign w42971 = w35811 & w36001;
assign w42972 = ~w35811 & w36003;
assign w42973 = w35811 & w36006;
assign w42974 = ~w35811 & w36008;
assign w42975 = (~w42968 & w48232) | (~w42968 & w48233) | (w48232 & w48233);
assign w42976 = (w48234 & w50401) | (w48234 & w42968) | (w50401 & w42968);
assign w42977 = w35983 & w46760;
assign w42978 = w35634 & w36025;
assign w42979 = w35328 & w35668;
assign w42980 = (w48235 & w50402) | (w48235 & w42968) | (w50402 & w42968);
assign w42981 = (w48236 & w50403) | (w48236 & w42968) | (w50403 & w42968);
assign w42982 = (~w42968 & w48237) | (~w42968 & w48238) | (w48237 & w48238);
assign w42983 = (w48239 & w50404) | (w48239 & w42968) | (w50404 & w42968);
assign w42984 = w35980 & w29158;
assign w42985 = (w48240 & w50405) | (w48240 & w42968) | (w50405 & w42968);
assign w42986 = (w48241 & w50406) | (w48241 & w42968) | (w50406 & w42968);
assign w42987 = (~w42968 & w48242) | (~w42968 & w48243) | (w48242 & w48243);
assign w42988 = (w48244 & w50407) | (w48244 & w42968) | (w50407 & w42968);
assign w42989 = (w48245 & w50408) | (w48245 & w42968) | (w50408 & w42968);
assign w42990 = (~w42968 & w48246) | (~w42968 & w48247) | (w48246 & w48247);
assign w42991 = (w48248 & w50409) | (w48248 & w42968) | (w50409 & w42968);
assign w42992 = (~w42968 & w48249) | (~w42968 & w48250) | (w48249 & w48250);
assign w42993 = w35980 & ~w36169;
assign w42994 = (~w42968 & w48251) | (~w42968 & w48252) | (w48251 & w48252);
assign w42995 = (w42968 & w48253) | (w42968 & w48254) | (w48253 & w48254);
assign w42996 = (w48255 & w50410) | (w48255 & w42968) | (w50410 & w42968);
assign w42997 = w36228 & w36243;
assign w42998 = ~w35980 & w35228;
assign w42999 = w35980 & w36255;
assign w43000 = ~w35139 & w35279;
assign w43001 = ~w35980 & w36273;
assign w43002 = ~w35980 & w36283;
assign w43003 = ~w35980 & ~w35213;
assign w43004 = w35980 & w36292;
assign w43005 = ~w35980 & w36297;
assign w43006 = w36228 & w36304;
assign w43007 = ~w35980 & w36310;
assign w43008 = ~w35980 & w36317;
assign w43009 = w36228 & ~w35250;
assign w43010 = ~w35980 & w36328;
assign w43011 = ~w35980 & w36338;
assign w43012 = ~w35980 & w36343;
assign w43013 = ~w35980 & ~w35236;
assign w43014 = w35980 & w36272;
assign w43015 = w35980 & ~w36359;
assign w43016 = ~w36372 & w35308;
assign w43017 = w36372 & ~w35308;
assign w43018 = w36389 & w35543;
assign w43019 = w35980 & w35480;
assign w43020 = (w36401 & w36393) | (w36401 & w43807) | (w36393 & w43807);
assign w43021 = w36389 & w36413;
assign w43022 = ~w36414 & w43808;
assign w43023 = ~w7924 & w36411;
assign w43024 = ~w35978 & w50235;
assign w43025 = (w36431 & w36393) | (w36431 & w43809) | (w36393 & w43809);
assign w43026 = ~w36455 & w36457;
assign w43027 = ~w36455 & ~w35542;
assign w43028 = ~w36469 & ~w36458;
assign w43029 = w36478 & w36476;
assign w43030 = ~w36478 & ~w36476;
assign w43031 = ~w35980 & ~w35553;
assign w43032 = w36484 & ~w10419;
assign w43033 = ~w36389 & ~w36488;
assign w43034 = w36389 & w36488;
assign w43035 = w35328 & ~w35618;
assign w43036 = w36504 & w35616;
assign w43037 = ~w36504 & w36506;
assign w43038 = ~w35980 & w36510;
assign w43039 = ~w36502 & w36517;
assign w43040 = w35980 & ~w36528;
assign w43041 = ~w36484 & w10419;
assign w43042 = ~w36502 & w36540;
assign w43043 = w36502 & w36542;
assign w43044 = w36550 & w36475;
assign w43045 = ~w36475 & ~w36464;
assign w43046 = w36571 & ~w36575;
assign w43047 = ~w35775 & ~w35799;
assign w43048 = w35980 & ~w36578;
assign w43049 = ~w35980 & w35791;
assign w43050 = ~w35980 & ~w35791;
assign w43051 = ~w35775 & ~w35807;
assign w43052 = ~w35760 & w35747;
assign w43053 = w35980 & w36606;
assign w43054 = ~w35980 & ~w1320;
assign w43055 = ~w35980 & w1320;
assign w43056 = w35980 & w36631;
assign w43057 = w35634 & w35743;
assign w43058 = ~w35980 & w1541;
assign w43059 = ~w36642 & w36651;
assign w43060 = w35980 & ~w36673;
assign w43061 = ~w35760 & w36675;
assign w43062 = w35980 & ~w2285;
assign w43063 = (~w42968 & w48257) | (~w42968 & w48258) | (w48257 & w48258);
assign w43064 = ~w35993 & w48259;
assign w43065 = (~w36692 & w35993) | (~w36692 & w48260) | (w35993 & w48260);
assign w43066 = ~w36603 & w36665;
assign w43067 = ~w36642 & w36720;
assign w43068 = ~w36630 & ~w36716;
assign w43069 = ~w36740 & ~w36741;
assign w43070 = w36740 & w36741;
assign w43071 = ~w36748 & ~w35932;
assign w43072 = (w48261 & w50411) | (w48261 & w42968) | (w50411 & w42968);
assign w43073 = (~w42968 & w48262) | (~w42968 & w48263) | (w48262 & w48263);
assign w43074 = (~w42968 & w48264) | (~w42968 & w48265) | (w48264 & w48265);
assign w43075 = ~w36765 & ~w36764;
assign w43076 = ~w35980 & w612;
assign w43077 = w36795 & w36783;
assign w43078 = ~w35635 & w35665;
assign w43079 = w3646 & w35392;
assign w43080 = (~w36834 & ~w35994) | (~w36834 & w43810) | (~w35994 & w43810);
assign w43081 = w35994 & w43811;
assign w43082 = ~w36828 & w36834;
assign w43083 = w35980 & ~w36842;
assign w43084 = w36867 & ~w36864;
assign w43085 = ~w36867 & w36864;
assign w43086 = w36883 & ~w36878;
assign w43087 = ~w36883 & w36878;
assign w43088 = w35328 & w36881;
assign w43089 = ~w35980 & w36899;
assign w43090 = ~w35980 & w36903;
assign w43091 = ~w35980 & w35646;
assign w43092 = w36916 & ~w36921;
assign w43093 = ~w35669 & w4056;
assign w43094 = ~w36929 & w35579;
assign w43095 = w36929 & ~w36932;
assign w43096 = w35328 & w36940;
assign w43097 = w35328 & w36952;
assign w43098 = ~w35980 & w35660;
assign w43099 = ~w36955 & ~w4056;
assign w43100 = ~w36929 & w36960;
assign w43101 = w36929 & w36962;
assign w43102 = w35980 & w35946;
assign w43103 = ~w36975 & ~w35859;
assign w43104 = (w48266 & w50412) | (w48266 & w42968) | (w50412 & w42968);
assign w43105 = w35980 & w37003;
assign w43106 = w35994 & w43812;
assign w43107 = (w37011 & ~w35994) | (w37011 & w43813) | (~w35994 & w43813);
assign w43108 = w36975 & w35947;
assign w43109 = ~w35980 & w37074;
assign w43110 = ~w35980 & w37082;
assign w43111 = w36955 & w4056;
assign w43112 = ~w36850 & w46761;
assign w43113 = ~w37102 & w37057;
assign w43114 = ~w37110 & ~w37109;
assign w43115 = ~w37110 & w37141;
assign w43116 = (w37172 & ~w37168) | (w37172 & w43814) | (~w37168 & w43814);
assign w43117 = ~w37110 & w37168;
assign w43118 = (~w37171 & ~w37168) | (~w37171 & w43815) | (~w37168 & w43815);
assign w43119 = ~w37169 & w37207;
assign w43120 = (~w37064 & ~w37225) | (~w37064 & w43816) | (~w37225 & w43816);
assign w43121 = ~w37110 & w37225;
assign w43122 = ~w37110 & w37256;
assign w43123 = w37057 & w46762;
assign w43124 = w37057 & w46763;
assign w43125 = w37057 & w46764;
assign w43126 = w37057 & w46765;
assign w43127 = w37057 & w46766;
assign w43128 = w37057 & w46767;
assign w43129 = w37057 & w46768;
assign w43130 = ~w37698 & ~w36549;
assign w43131 = ~w36552 & w36573;
assign w43132 = ~w37698 & w37907;
assign w43133 = w37057 & w46769;
assign w43134 = w36571 & ~w37997;
assign w43135 = w37057 & w46770;
assign w43136 = ~w38040 & ~w38041;
assign w43137 = w37057 & w46771;
assign w43138 = w37057 & w46772;
assign w43139 = (w38094 & w36575) | (w38094 & w43817) | (w36575 & w43817);
assign w43140 = (w38100 & w36575) | (w38100 & w43818) | (w36575 & w43818);
assign w43141 = w37106 & ~w4430;
assign w43142 = ~w38109 & w38108;
assign w43143 = w38109 & ~w38108;
assign w43144 = ~w38104 & w4056;
assign w43145 = (w38130 & w37107) | (w38130 & w43819) | (w37107 & w43819);
assign w43146 = ~w37107 & w43820;
assign w43147 = ~w38136 & w38138;
assign w43148 = w37106 & w38152;
assign w43149 = w2558 & w38178;
assign w43150 = ~w2558 & w38183;
assign w43151 = ~w38198 & w38199;
assign w43152 = w37106 & ~w57;
assign w43153 = ~w38198 & w38211;
assign w43154 = ~w37106 & w37013;
assign w43155 = w37106 & ~w3;
assign w43156 = ~w37309 & w351;
assign w43157 = ~w37301 & w38257;
assign w43158 = w37106 & ~w36761;
assign w43159 = ~w37114 & w38275;
assign w43160 = ~w37106 & ~w252;
assign w43161 = ~w37106 & w252;
assign w43162 = ~w37316 & w38328;
assign w43163 = w37315 & w38292;
assign w43164 = ~w38337 & w43821;
assign w43165 = (w38380 & w38337) | (w38380 & w43822) | (w38337 & w43822);
assign w43166 = (~w38403 & w38337) | (~w38403 & w43823) | (w38337 & w43823);
assign w43167 = (~w38433 & w38337) | (~w38433 & w43824) | (w38337 & w43824);
assign w43168 = (w38452 & w38337) | (w38452 & w43825) | (w38337 & w43825);
assign w43169 = ~w38337 & w43826;
assign w43170 = (w38448 & w38337) | (w38448 & w43827) | (w38337 & w43827);
assign w43171 = (w38469 & w38337) | (w38469 & w43828) | (w38337 & w43828);
assign w43172 = ~w37494 & w37369;
assign w43173 = (w38485 & w38337) | (w38485 & w43829) | (w38337 & w43829);
assign w43174 = (w38336 & w43830) | (w38336 & w43831) | (w43830 & w43831);
assign w43175 = ~w38338 & w38501;
assign w43176 = ~w38338 & w38509;
assign w43177 = w37694 & w43832;
assign w43178 = (~w38525 & w37678) | (~w38525 & w43833) | (w37678 & w43833);
assign w43179 = w38533 & ~w38536;
assign w43180 = ~w38533 & w38536;
assign w43181 = (w38526 & w38337) | (w38526 & w43834) | (w38337 & w43834);
assign w43182 = (~w37829 & w37678) | (~w37829 & w43835) | (w37678 & w43835);
assign w43183 = ~w38337 & w43836;
assign w43184 = ~w38338 & w38544;
assign w43185 = ~w38338 & ~w38555;
assign w43186 = w38338 & w38564;
assign w43187 = w38554 & ~w38540;
assign w43188 = ~w38578 & ~w37823;
assign w43189 = ~w38583 & w37753;
assign w43190 = ~w38578 & w38585;
assign w43191 = ~w38337 & w43837;
assign w43192 = ~w38592 & w38597;
assign w43193 = ~w38336 & w43838;
assign w43194 = w37667 & w22767;
assign w43195 = ~w37667 & ~w22767;
assign w43196 = (w38681 & w37678) | (w38681 & w43839) | (w37678 & w43839);
assign w43197 = ~w37678 & w43840;
assign w43198 = ~w38338 & ~w38685;
assign w43199 = ~w37677 & ~w37639;
assign w43200 = (w38336 & w43841) | (w38336 & w43842) | (w43841 & w43842);
assign w43201 = ~w38338 & ~w38875;
assign w43202 = (w38590 & w38336) | (w38590 & w43843) | (w38336 & w43843);
assign w43203 = (~w37775 & w38337) | (~w37775 & w43844) | (w38337 & w43844);
assign w43204 = ~w37985 & w38162;
assign w43205 = w10419 & ~w37954;
assign w43206 = ~w10419 & ~w38159;
assign w43207 = w37939 & ~w37987;
assign w43208 = ~w38959 & w38962;
assign w43209 = (w39026 & w39031) | (w39026 & w43845) | (w39031 & w43845);
assign w43210 = ~w39031 & w43846;
assign w43211 = ~w39028 & w39051;
assign w43212 = (~w38136 & ~w39093) | (~w38136 & w43847) | (~w39093 & w43847);
assign w43213 = (~w39095 & ~w39093) | (~w39095 & w43848) | (~w39093 & w43848);
assign w43214 = ~w38338 & ~w2285;
assign w43215 = (w39152 & ~w39093) | (w39152 & w43849) | (~w39093 & w43849);
assign w43216 = (w2285 & w38337) | (w2285 & w43850) | (w38337 & w43850);
assign w43217 = (w39169 & w38176) | (w39169 & w43851) | (w38176 & w43851);
assign w43218 = (w37272 & w38142) | (w37272 & w43852) | (w38142 & w43852);
assign w43219 = (~w39168 & w38176) | (~w39168 & w43853) | (w38176 & w43853);
assign w43220 = ~w39175 & w43854;
assign w43221 = (w39151 & ~w39093) | (w39151 & w43855) | (~w39093 & w43855);
assign w43222 = ~w39032 & ~w37867;
assign w43223 = ~w38337 & w43856;
assign w43224 = (w39300 & w38336) | (w39300 & w43857) | (w38336 & w43857);
assign w43225 = ~w38336 & w43858;
assign w43226 = ~w37316 & w38271;
assign w43227 = ~w38176 & w46773;
assign w43228 = ~w37316 & w38291;
assign w43229 = w38140 & w38189;
assign w43230 = ~w39414 & w37286;
assign w43231 = w39414 & w37248;
assign w43232 = ~w38176 & w43859;
assign w43233 = ~w38176 & w43860;
assign w43234 = ~w38337 & w43861;
assign w43235 = ~w39414 & w37279;
assign w43236 = (w39508 & w38336) | (w39508 & w43862) | (w38336 & w43862);
assign w43237 = ~w38336 & w43863;
assign w43238 = ~w39415 & w37239;
assign w43239 = ~w38337 & w43864;
assign w43240 = w39172 & w39581;
assign w43241 = ~w38339 & w39586;
assign w43242 = w38339 & w39589;
assign w43243 = ~w612 & ~w38339;
assign w43244 = ~w187 & w42;
assign w43245 = w239 & w80;
assign w43246 = ~w239 & ~w80;
assign w43247 = w379 & a[119];
assign w43248 = ~w379 & ~a[119];
assign w43249 = ~w369 & ~w3;
assign w43250 = w369 & w3;
assign w43251 = ~w642 & w80;
assign w43252 = ~w870 & ~w869;
assign w43253 = w400 & w351;
assign w43254 = ~w400 & ~w351;
assign w43255 = w819 & ~w3;
assign w43256 = w1292 & ~w1314;
assign w43257 = ~w1224 & ~w1329;
assign w43258 = w1224 & ~w1340;
assign w43259 = ~w1224 & w1347;
assign w43260 = ~w1224 & w1359;
assign w43261 = w1224 & w1361;
assign w43262 = w1224 & w1367;
assign w43263 = ~w1224 & w1366;
assign w43264 = w1224 & w1372;
assign w43265 = ~w1224 & w1374;
assign w43266 = ~w1224 & w1384;
assign w43267 = w1224 & ~w1387;
assign w43268 = ~w612 & w493;
assign w43269 = w1406 & ~w1407;
assign w43270 = ~w1397 & w1419;
assign w43271 = w1397 & w1421;
assign w43272 = ~w1397 & w1287;
assign w43273 = w1397 & ~w1287;
assign w43274 = ~w1224 & ~w1466;
assign w43275 = ~w1224 & w1466;
assign w43276 = w1508 & w1565;
assign w43277 = ~w1508 & w1567;
assign w43278 = w1508 & ~w1576;
assign w43279 = ~w1508 & w1583;
assign w43280 = w1508 & w1617;
assign w43281 = ~w1508 & w1619;
assign w43282 = w1508 & w1390;
assign w43283 = ~w1508 & w1616;
assign w43284 = (w1877 & ~w1649) | (w1877 & w46774) | (~w1649 & w46774);
assign w43285 = w1649 & w46775;
assign w43286 = (w1892 & ~w1649) | (w1892 & w46776) | (~w1649 & w46776);
assign w43287 = w1649 & w46777;
assign w43288 = w252 & w1911;
assign w43289 = ~w252 & w1913;
assign w43290 = ~w1901 & w1924;
assign w43291 = w252 & w1957;
assign w43292 = ~w252 & w1959;
assign w43293 = w2004 & w2116;
assign w43294 = w2004 & w1860;
assign w43295 = w351 & w1860;
assign w43296 = w351 & w39918;
assign w43297 = ~w2279 & w2133;
assign w43298 = ~w2517 & ~w57;
assign w43299 = ~w2586 & w2542;
assign w43300 = w2517 & ~w80;
assign w43301 = ~w2586 & w2620;
assign w43302 = ~w2438 & ~w400;
assign w43303 = w2438 & w400;
assign w43304 = ~w351 & w2662;
assign w43305 = ~w351 & w2672;
assign w43306 = w351 & w2674;
assign w43307 = ~w2517 & w2765;
assign w43308 = ~w2517 & ~w2767;
assign w43309 = ~w2517 & w2789;
assign w43310 = w2517 & w2800;
assign w43311 = ~w2517 & w2802;
assign w43312 = ~w2517 & w2806;
assign w43313 = w2517 & ~w2285;
assign w43314 = w2814 & w2006;
assign w43315 = ~w2517 & w2820;
assign w43316 = ~w2517 & w2818;
assign w43317 = ~w2517 & w2830;
assign w43318 = w2517 & w2832;
assign w43319 = ~w2814 & ~w2006;
assign w43320 = w2964 & w3258;
assign w43321 = ~w2964 & w3260;
assign w43322 = w2964 & ~w3276;
assign w43323 = ~w2964 & w3284;
assign w43324 = ~w2964 & w3289;
assign w43325 = w2964 & w3291;
assign w43326 = w2964 & w1320;
assign w43327 = w2964 & w3394;
assign w43328 = ~w40061 & w3403;
assign w43329 = ~w40061 & w3406;
assign w43330 = ~w2964 & ~w2936;
assign w43331 = w2964 & ~w80;
assign w43332 = w2964 & w3;
assign w43333 = ~w40090 & ~w3516;
assign w43334 = w40090 & w3516;
assign w43335 = w2964 & w57;
assign w43336 = w40098 & w3549;
assign w43337 = ~w40098 & w3551;
assign w43338 = w2964 & w2953;
assign w43339 = w40105 & w57;
assign w43340 = w3545 & ~w351;
assign w43341 = w3545 & w351;
assign w43342 = w3545 & w3621;
assign w43343 = w3545 & w3623;
assign w43344 = ~w3545 & w3754;
assign w43345 = ~w3545 & w3771;
assign w43346 = ~w3545 & ~w3247;
assign w43347 = ~w3545 & w3797;
assign w43348 = w3605 & w3986;
assign w43349 = ~w3995 & ~w80;
assign w43350 = ~w3545 & ~w3597;
assign w43351 = w3605 & w4033;
assign w43352 = w4123 & ~w42;
assign w43353 = ~w4123 & w42;
assign w43354 = w3661 & w252;
assign w43355 = ~w3737 & w4188;
assign w43356 = (~w3737 & ~w3888) | (~w3737 & w43355) | (~w3888 & w43355);
assign w43357 = ~w4380 & w46778;
assign w43358 = ~w4385 & w1120;
assign w43359 = w4377 & ~w1120;
assign w43360 = ~w4377 & w1120;
assign w43361 = w4396 & ~w4204;
assign w43362 = ~w4431 & w4112;
assign w43363 = (~w4111 & w4184) | (~w4111 & w48267) | (w4184 & w48267);
assign w43364 = ~w4717 & w4168;
assign w43365 = w4611 & ~w4851;
assign w43366 = ~w4742 & ~w5052;
assign w43367 = w4742 & w5052;
assign w43368 = (~w4663 & w4742) | (~w4663 & w48268) | (w4742 & w48268);
assign w43369 = w40251 & ~w5134;
assign w43370 = ~w40262 & w5226;
assign w43371 = ~w40264 & ~w4818;
assign w43372 = ~w40262 & w4835;
assign w43373 = ~w4904 & ~w4877;
assign w43374 = ~w5290 & w5102;
assign w43375 = w5747 & w5746;
assign w43376 = ~w5747 & ~w5746;
assign w43377 = ~w5839 & ~w57;
assign w43378 = w5743 & ~w351;
assign w43379 = w5743 & w5482;
assign w43380 = w40333 & ~w1320;
assign w43381 = w5979 & ~w5981;
assign w43382 = w4838 & w5981;
assign w43383 = (w5743 & w43382) | (w5743 & w49323) | (w43382 & w49323);
assign w43384 = (w5732 & w49324) | (w5732 & w49325) | (w49324 & w49325);
assign w43385 = (w1320 & w5732) | (w1320 & w48269) | (w5732 & w48269);
assign w43386 = ~w5732 & w48270;
assign w43387 = (w6252 & w5732) | (w6252 & w48271) | (w5732 & w48271);
assign w43388 = w6345 & w5330;
assign w43389 = w945 & w6211;
assign w43390 = ~w754 & w6211;
assign w43391 = w6570 & w48272;
assign w43392 = w6583 & w945;
assign w43393 = ~w6767 & w6318;
assign w43394 = ~w6764 & w6319;
assign w43395 = ~w6764 & w6867;
assign w43396 = ~w6427 & ~w6426;
assign w43397 = w7151 & w80;
assign w43398 = ~w7151 & w7224;
assign w43399 = w6764 & ~w6316;
assign w43400 = ~w6767 & w7252;
assign w43401 = ~w7270 & w49326;
assign w43402 = w7394 & w48273;
assign w43403 = (w7399 & w7270) | (w7399 & w49327) | (w7270 & w49327);
assign w43404 = (w7399 & ~w7394) | (w7399 & w48274) | (~w7394 & w48274);
assign w43405 = w7086 & w7417;
assign w43406 = w7086 & w7269;
assign w43407 = ~w7802 & ~w7194;
assign w43408 = ~w7802 & ~w7801;
assign w43409 = w252 & w7814;
assign w43410 = ~w252 & w7816;
assign w43411 = w1320 & ~w7468;
assign w43412 = w1320 & w40494;
assign w43413 = ~w7949 & ~w7923;
assign w43414 = w7979 & w7468;
assign w43415 = w7979 & ~w40494;
assign w43416 = ~w7783 & w754;
assign w43417 = w7935 & ~w7932;
assign w43418 = ~w7935 & w7932;
assign w43419 = ~w945 & w7927;
assign w43420 = ~w945 & w40545;
assign w43421 = ~w7783 & ~w8227;
assign w43422 = ~w7783 & ~w8235;
assign w43423 = ~w7783 & w4056;
assign w43424 = ~w7783 & ~w8373;
assign w43425 = ~w7783 & ~w2285;
assign w43426 = ~w7783 & w8505;
assign w43427 = w8539 & ~w2896;
assign w43428 = w9609 & ~w10107;
assign w43429 = w10129 & ~w40794;
assign w43430 = w10129 & ~w10112;
assign w43431 = ~w3 & w10211;
assign w43432 = w3 & w10213;
assign w43433 = ~w10339 & ~w9295;
assign w43434 = ~w10339 & w10358;
assign w43435 = w252 & w10405;
assign w43436 = ~w252 & w10407;
assign w43437 = w10388 & ~w10351;
assign w43438 = ~w10575 & ~w10578;
assign w43439 = w10656 & w80;
assign w43440 = w10656 & w40875;
assign w43441 = w10674 & w1120;
assign w43442 = w10674 & w40881;
assign w43443 = ~w10376 & ~w9823;
assign w43444 = ~w10376 & w9836;
assign w43445 = w2558 & w10085;
assign w43446 = w2558 & w40896;
assign w43447 = ~w10545 & ~w10592;
assign w43448 = ~w10868 & w10683;
assign w43449 = ~w10868 & w10684;
assign w43450 = ~w40952 & w10808;
assign w43451 = ~w10933 & w11346;
assign w43452 = ~w10645 & w6264;
assign w43453 = w11580 & ~w11232;
assign w43454 = w10863 & ~w11591;
assign w43455 = w10863 & w11611;
assign w43456 = w10863 & ~w11626;
assign w43457 = w10863 & w11835;
assign w43458 = ~w11864 & ~w11869;
assign w43459 = ~w11864 & w11905;
assign w43460 = ~w11864 & w11946;
assign w43461 = ~w11864 & w11949;
assign w43462 = ~w11864 & w11954;
assign w43463 = ~w11864 & w11962;
assign w43464 = ~w11864 & w11981;
assign w43465 = ~w11968 & w11983;
assign w43466 = ~w11968 & ~w11966;
assign w43467 = ~w11864 & w12023;
assign w43468 = w11435 & w11343;
assign w43469 = ~w12234 & ~w12237;
assign w43470 = w12280 & ~w41053;
assign w43471 = w12280 & ~w41052;
assign w43472 = w12293 & ~w41053;
assign w43473 = w12293 & ~w41052;
assign w43474 = w12307 & ~w41056;
assign w43475 = w12307 & ~w41057;
assign w43476 = w12523 & ~w351;
assign w43477 = ~w12143 & w12159;
assign w43478 = ~w12858 & w4056;
assign w43479 = w12858 & ~w4056;
assign w43480 = ~w12912 & w48275;
assign w43481 = w1120 & w13051;
assign w43482 = w13280 & ~w13740;
assign w43483 = w13280 & ~w13089;
assign w43484 = w13859 & ~w13358;
assign w43485 = ~w13859 & ~w13876;
assign w43486 = ~w13885 & w13131;
assign w43487 = w13840 & ~w14491;
assign w43488 = w14490 & ~w13937;
assign w43489 = ~w14761 & w14671;
assign w43490 = ~w14753 & w14516;
assign w43491 = ~w15024 & w15020;
assign w43492 = w15024 & ~w15020;
assign w43493 = ~w15247 & ~w6769;
assign w43494 = ~w15288 & ~w7315;
assign w43495 = w15288 & w7315;
assign w43496 = w15314 & ~w15319;
assign w43497 = ~w15314 & w15319;
assign w43498 = ~w15314 & w15336;
assign w43499 = w15314 & w15338;
assign w43500 = ~a[51] & ~w14039;
assign w43501 = ~a[51] & w15423;
assign w43502 = ~w16086 & w16085;
assign w43503 = w16086 & ~w16085;
assign w43504 = ~w16130 & w16273;
assign w43505 = ~w14972 & w46779;
assign w43506 = ~w14925 & ~w14969;
assign w43507 = w14966 & w14982;
assign w43508 = ~w16521 & w48276;
assign w43509 = w16522 & w16537;
assign w43510 = w16610 & ~w612;
assign w43511 = ~w16270 & w50236;
assign w43512 = ~w16620 & ~w16621;
assign w43513 = w16281 & ~w16516;
assign w43514 = w16522 & w16737;
assign w43515 = w16522 & w16540;
assign w43516 = ~w16868 & ~w16040;
assign w43517 = w15871 & ~w15886;
assign w43518 = w41412 & ~w7315;
assign w43519 = ~w41412 & w7315;
assign w43520 = ~w17153 & ~w9195;
assign w43521 = w17443 & w6769;
assign w43522 = w17045 & w16949;
assign w43523 = ~w17045 & w16951;
assign w43524 = ~w3242 & w17804;
assign w43525 = w17357 & ~w2006;
assign w43526 = ~w41631 & ~w2896;
assign w43527 = w19100 & w2558;
assign w43528 = w19147 & w18668;
assign w43529 = ~w19236 & ~w19221;
assign w43530 = w19236 & w19221;
assign w43531 = w41649 & w19253;
assign w43532 = ~w41649 & w19255;
assign w43533 = ~w19794 & ~w612;
assign w43534 = w18957 & ~w19819;
assign w43535 = w18957 & ~w41720;
assign w43536 = w18917 & ~w42;
assign w43537 = ~w41724 & ~w80;
assign w43538 = ~w18917 & w42;
assign w43539 = w20035 & w20301;
assign w43540 = ~w20035 & ~w20301;
assign w43541 = w5330 & ~w20318;
assign w43542 = ~w5330 & ~w20320;
assign w43543 = ~w5745 & w20334;
assign w43544 = w5745 & w20337;
assign w43545 = w5330 & w20361;
assign w43546 = ~w5330 & w20364;
assign w43547 = ~w19626 & ~w20637;
assign w43548 = w10419 & w20668;
assign w43549 = ~w10419 & w20671;
assign w43550 = ~w20705 & w10419;
assign w43551 = w10419 & w20736;
assign w43552 = ~w10419 & w20739;
assign w43553 = w20713 & w20678;
assign w43554 = w20713 & w20676;
assign w43555 = w20326 & ~w21324;
assign w43556 = ~w20210 & w21442;
assign w43557 = ~w20210 & w20201;
assign w43558 = ~w20210 & w21473;
assign w43559 = ~w20904 & w21566;
assign w43560 = w20904 & w21568;
assign w43561 = ~w20904 & w20384;
assign w43562 = w20904 & ~w20384;
assign w43563 = ~w21341 & w22712;
assign w43564 = w23066 & w23075;
assign w43565 = ~w23066 & w23077;
assign w43566 = w23160 & ~w23166;
assign w43567 = ~w23160 & w23166;
assign w43568 = w23242 & w11870;
assign w43569 = ~w23264 & ~w23265;
assign w43570 = ~w23242 & ~w11870;
assign w43571 = ~w21969 & w22647;
assign w43572 = w21970 & w22647;
assign w43573 = w945 & w23546;
assign w43574 = ~w945 & w23546;
assign w43575 = w945 & w23556;
assign w43576 = ~w945 & w23556;
assign w43577 = w945 & w23564;
assign w43578 = ~w945 & w23564;
assign w43579 = w945 & w23570;
assign w43580 = ~w945 & w23570;
assign w43581 = ~w23205 & ~w14766;
assign w43582 = ~w24266 & ~w24267;
assign w43583 = w24010 & w11870;
assign w43584 = ~w25048 & ~w9781;
assign w43585 = w25048 & w9781;
assign w43586 = ~w25303 & ~w16559;
assign w43587 = w25351 & w48277;
assign w43588 = w24331 & ~w24288;
assign w43589 = w24313 & ~w24585;
assign w43590 = w25402 & w1120;
assign w43591 = w25402 & w42146;
assign w43592 = w25404 & ~w1120;
assign w43593 = w25404 & ~w42146;
assign w43594 = w25419 & ~w1541;
assign w43595 = w25419 & ~w42149;
assign w43596 = w25421 & w1541;
assign w43597 = w25421 & w42149;
assign w43598 = ~w25418 & ~w1541;
assign w43599 = ~w25418 & ~w42149;
assign w43600 = w25418 & w1541;
assign w43601 = w25418 & w42149;
assign w43602 = w25569 & ~w4838;
assign w43603 = w25569 & w42183;
assign w43604 = w25625 & w3242;
assign w43605 = w25625 & w42196;
assign w43606 = ~w25686 & ~w252;
assign w43607 = ~w25686 & w42207;
assign w43608 = ~w493 & w24632;
assign w43609 = w25307 & w25313;
assign w43610 = w25307 & ~w25312;
assign w43611 = (w26065 & w26861) | (w26065 & w48278) | (w26861 & w48278);
assign w43612 = ~w26318 & w27089;
assign w43613 = (w26720 & w26317) | (w26720 & w46780) | (w26317 & w46780);
assign w43614 = (w26718 & w26317) | (w26718 & w46781) | (w26317 & w46781);
assign w43615 = ~w26688 & ~w27488;
assign w43616 = w26688 & w27488;
assign w43617 = ~w26944 & w26282;
assign w43618 = ~w27726 & w10419;
assign w43619 = w27726 & ~w10419;
assign w43620 = (w28080 & w28036) | (w28080 & w49834) | (w28036 & w49834);
assign w43621 = ~w28037 & w28099;
assign w43622 = (~w28036 & w49835) | (~w28036 & w49836) | (w49835 & w49836);
assign w43623 = ~w28037 & w28183;
assign w43624 = (~w28193 & w46783) | (~w28193 & w28037) | (w46783 & w28037);
assign w43625 = w28037 & w20000;
assign w43626 = ~w28037 & w28275;
assign w43627 = ~w28321 & w46784;
assign w43628 = ~w28036 & w49837;
assign w43629 = w28419 & ~w14039;
assign w43630 = (w27616 & w28433) | (w27616 & w48279) | (w28433 & w48279);
assign w43631 = ~w28433 & w48280;
assign w43632 = (~w27482 & w28037) | (~w27482 & w49838) | (w28037 & w49838);
assign w43633 = w28037 & ~w27401;
assign w43634 = w28037 & w9781;
assign w43635 = (~w28512 & w28036) | (~w28512 & w49839) | (w28036 & w49839);
assign w43636 = ~w28036 & w49840;
assign w43637 = ~w28036 & w49841;
assign w43638 = w28528 & ~w5330;
assign w43639 = ~w28049 & w46785;
assign w43640 = w28530 & w5330;
assign w43641 = (w28530 & w28049) | (w28530 & w46786) | (w28049 & w46786);
assign w43642 = ~w28527 & w5330;
assign w43643 = (~w28527 & w28049) | (~w28527 & w46787) | (w28049 & w46787);
assign w43644 = w28527 & ~w5330;
assign w43645 = ~w28049 & w46788;
assign w43646 = (w42366 & w50150) | (w42366 & w50151) | (w50150 & w50151);
assign w43647 = (w7315 & w28036) | (w7315 & w49842) | (w28036 & w49842);
assign w43648 = ~w28036 & w49843;
assign w43649 = w27881 & w27216;
assign w43650 = w28037 & w28646;
assign w43651 = w8666 & ~w28646;
assign w43652 = (w8666 & w28049) | (w8666 & w46789) | (w28049 & w46789);
assign w43653 = ~w28036 & w49844;
assign w43654 = w28037 & w493;
assign w43655 = w28759 & w493;
assign w43656 = w28759 & w42391;
assign w43657 = ~w28696 & w252;
assign w43658 = ~w28049 & w46790;
assign w43659 = (~w80 & w28036) | (~w80 & w49845) | (w28036 & w49845);
assign w43660 = w3 & w28858;
assign w43661 = w3 & ~w42404;
assign w43662 = (w28001 & w28036) | (w28001 & w49846) | (w28036 & w49846);
assign w43663 = w57 & w28878;
assign w43664 = ~w57 & w28880;
assign w43665 = ~w28037 & w28943;
assign w43666 = w28037 & w28954;
assign w43667 = ~w28037 & w1541;
assign w43668 = ~w28036 & w49847;
assign w43669 = w2006 & w27196;
assign w43670 = ~w28049 & w46791;
assign w43671 = w27202 & w29054;
assign w43672 = ~w42420 & w2558;
assign w43673 = ~w28037 & ~w29078;
assign w43674 = w27177 & ~w2896;
assign w43675 = (~w29092 & ~w45723) | (~w29092 & w48281) | (~w45723 & w48281);
assign w43676 = ~w28036 & w49848;
assign w43677 = w29123 & w3646;
assign w43678 = ~w28049 & w46792;
assign w43679 = w29125 & ~w3646;
assign w43680 = (w29125 & w28049) | (w29125 & w46793) | (w28049 & w46793);
assign w43681 = ~w29122 & ~w3646;
assign w43682 = (~w29122 & w28049) | (~w29122 & w46794) | (w28049 & w46794);
assign w43683 = w29122 & w3646;
assign w43684 = ~w28049 & w46795;
assign w43685 = ~w29350 & w28472;
assign w43686 = ~w28929 & w29416;
assign w43687 = ~w29350 & w29643;
assign w43688 = w29350 & w29645;
assign w43689 = w30026 & w30241;
assign w43690 = ~w30026 & ~w30241;
assign w43691 = w30339 & ~w30246;
assign w43692 = w29485 & ~w29489;
assign w43693 = ~w29653 & ~w29336;
assign w43694 = (~w2006 & w30205) | (~w2006 & w46796) | (w30205 & w46796);
assign w43695 = w31469 & w31500;
assign w43696 = w31469 & ~w30509;
assign w43697 = w31469 & w31541;
assign w43698 = w57 & w31534;
assign w43699 = ~w14766 & w31580;
assign w43700 = w14766 & w31584;
assign w43701 = w31662 & ~w30877;
assign w43702 = ~w31662 & w31669;
assign w43703 = w31662 & w31671;
assign w43704 = w31684 & w31690;
assign w43705 = ~w31684 & w31692;
assign w43706 = w31684 & w31698;
assign w43707 = ~w31684 & w31700;
assign w43708 = ~w31784 & ~w31785;
assign w43709 = w31469 & w30517;
assign w43710 = ~w31818 & ~w31819;
assign w43711 = ~w31810 & w31852;
assign w43712 = ~w31872 & ~w31873;
assign w43713 = (~w31966 & ~w31964) | (~w31966 & w46797) | (~w31964 & w46797);
assign w43714 = w31996 & w32002;
assign w43715 = ~w31996 & w32004;
assign w43716 = w31996 & w32033;
assign w43717 = ~w31996 & w30588;
assign w43718 = ~w30468 & w46798;
assign w43719 = ~w31193 & ~w4838;
assign w43720 = ~w754 & w32445;
assign w43721 = w754 & ~w32445;
assign w43722 = ~w30511 & w32483;
assign w43723 = ~w31492 & w32492;
assign w43724 = ~w32454 & ~w30507;
assign w43725 = ~w32722 & ~w32721;
assign w43726 = ~w32510 & ~w32579;
assign w43727 = ~w400 & w32444;
assign w43728 = w400 & ~w32444;
assign w43729 = ~w400 & ~w32444;
assign w43730 = ~w32375 & w32554;
assign w43731 = w754 & w32826;
assign w43732 = ~w754 & w32828;
assign w43733 = w945 & w32850;
assign w43734 = ~w945 & w32852;
assign w43735 = ~w32250 & ~w32236;
assign w43736 = w32422 & w46799;
assign w43737 = ~w754 & ~w32825;
assign w43738 = w754 & w32825;
assign w43739 = ~w33001 & ~w31971;
assign w43740 = ~w33019 & w33020;
assign w43741 = w33019 & w33023;
assign w43742 = w33001 & w33030;
assign w43743 = ~w33001 & w33032;
assign w43744 = ~w33019 & w33072;
assign w43745 = w33019 & w33075;
assign w43746 = w10419 & ~w33632;
assign w43747 = ~w32789 & w46800;
assign w43748 = ~w32968 & w33788;
assign w43749 = (w32872 & w32967) | (w32872 & w49328) | (w32967 & w49328);
assign w43750 = w32790 & w33861;
assign w43751 = ~w32790 & w33863;
assign w43752 = w32710 & ~w33869;
assign w43753 = ~w33872 & w50238;
assign w43754 = w32790 & w33879;
assign w43755 = ~w32790 & w33881;
assign w43756 = ~w32790 & w33892;
assign w43757 = ~w32790 & ~w33858;
assign w43758 = w32790 & ~w33896;
assign w43759 = w32790 & w33911;
assign w43760 = ~w32790 & w33877;
assign w43761 = w32790 & w33878;
assign w43762 = ~w32790 & ~w33004;
assign w43763 = w32790 & ~w33931;
assign w43764 = ~w33361 & w34209;
assign w43765 = w42745 & w34202;
assign w43766 = ~w42745 & ~w34202;
assign w43767 = w42745 & w34250;
assign w43768 = ~w42745 & w34252;
assign w43769 = ~w32968 & w32870;
assign w43770 = ~w32789 & w46801;
assign w43771 = w34642 & w50239;
assign w43772 = (w34745 & w32789) | (w34745 & w46802) | (w32789 & w46802);
assign w43773 = ~w32931 & ~w1738;
assign w43774 = (~w1541 & w32789) | (~w1541 & w46803) | (w32789 & w46803);
assign w43775 = ~w32997 & w46804;
assign w43776 = w32931 & w1738;
assign w43777 = w34856 & w49329;
assign w43778 = ~w24874 & w33855;
assign w43779 = ~w33852 & w34892;
assign w43780 = ~w34895 & w35085;
assign w43781 = ~w34114 & ~w19040;
assign w43782 = ~w42897 & w16559;
assign w43783 = w42897 & ~w16559;
assign w43784 = ~w42763 & ~w34588;
assign w43785 = w34877 & w33855;
assign w43786 = ~w34312 & w35419;
assign w43787 = ~w34312 & w35426;
assign w43788 = ~w33855 & ~w35432;
assign w43789 = w42914 & ~w8666;
assign w43790 = ~w42918 & ~w9781;
assign w43791 = w42918 & w9781;
assign w43792 = w42924 & ~w10419;
assign w43793 = (w8666 & ~w35454) | (w8666 & w46805) | (~w35454 & w46805);
assign w43794 = w35530 & w33855;
assign w43795 = ~w42924 & w10419;
assign w43796 = ~w42930 & w35580;
assign w43797 = w42930 & ~w35580;
assign w43798 = ~w35639 & w35641;
assign w43799 = ~w35692 & ~w35693;
assign w43800 = ~w35698 & ~w34835;
assign w43801 = w35679 & ~w35717;
assign w43802 = w42940 & w2285;
assign w43803 = ~w42947 & w35850;
assign w43804 = w42947 & ~w35850;
assign w43805 = ~w42956 & w35903;
assign w43806 = w42956 & w35905;
assign w43807 = ~w36392 & w36401;
assign w43808 = ~w36412 & ~w35463;
assign w43809 = ~w35518 & w36431;
assign w43810 = w3242 & ~w36834;
assign w43811 = ~w3242 & w36834;
assign w43812 = ~w252 & w37009;
assign w43813 = w252 & w37011;
assign w43814 = ~w37166 & w37172;
assign w43815 = ~w37166 & ~w37171;
assign w43816 = ~w37063 & ~w37064;
assign w43817 = ~w37086 & w38094;
assign w43818 = ~w37086 & w38100;
assign w43819 = ~w5330 & w38130;
assign w43820 = w5330 & w38132;
assign w43821 = w38325 & w38361;
assign w43822 = ~w38325 & w38380;
assign w43823 = ~w38325 & ~w38403;
assign w43824 = ~w38325 & ~w38433;
assign w43825 = ~w38325 & w38452;
assign w43826 = w38325 & ~w37472;
assign w43827 = ~w38325 & w38448;
assign w43828 = ~w38325 & w38469;
assign w43829 = ~w38325 & w38485;
assign w43830 = ~w38484 & w38485;
assign w43831 = ~w38484 & w43173;
assign w43832 = ~w37691 & ~w37810;
assign w43833 = ~w43177 & ~w38525;
assign w43834 = ~w38325 & w38526;
assign w43835 = ~w37695 & ~w37829;
assign w43836 = w38325 & w37809;
assign w43837 = w38325 & ~w12666;
assign w43838 = w43191 & w38599;
assign w43839 = ~w37694 & w38681;
assign w43840 = w37694 & ~w38681;
assign w43841 = w38771 & w38485;
assign w43842 = w38771 & w43173;
assign w43843 = ~w43191 & w38590;
assign w43844 = ~w38325 & ~w37775;
assign w43845 = w37878 & w39026;
assign w43846 = ~w37878 & ~w39026;
assign w43847 = w38120 & ~w38136;
assign w43848 = w4430 & ~w39095;
assign w43849 = w38120 & w39152;
assign w43850 = ~w38325 & w2285;
assign w43851 = w38140 & w39169;
assign w43852 = ~w43217 & w37272;
assign w43853 = w38140 & ~w39168;
assign w43854 = w2006 & ~w37272;
assign w43855 = w38120 & w39151;
assign w43856 = w38325 & w4838;
assign w43857 = ~w43223 & w39300;
assign w43858 = w43223 & ~w39300;
assign w43859 = ~w38140 & w39431;
assign w43860 = ~w38140 & w37287;
assign w43861 = w38325 & w1541;
assign w43862 = ~w43234 & w39508;
assign w43863 = w43234 & ~w39508;
assign w43864 = w38325 & ~w1738;
assign w43865 = w41 & ~w35;
assign w43866 = w105 & w50683;
assign w43867 = ~w160 & w230;
assign w43868 = w309 & ~w267;
assign w43869 = ~w228 & ~w212;
assign w43870 = w270 & w3;
assign w43871 = ~w233 & ~w337;
assign w43872 = w233 & ~w339;
assign w43873 = ~w233 & ~a[117];
assign w43874 = (w346 & ~w43873) | (w346 & w50684) | (~w43873 & w50684);
assign w43875 = w233 & ~w357;
assign w43876 = ~w233 & w378;
assign w43877 = (a[118] & ~w43876) | (a[118] & w50685) | (~w43876 & w50685);
assign w43878 = ~w397 & w416;
assign w43879 = w397 & w415;
assign w43880 = ~w396 & ~w388;
assign w43881 = ~w438 & ~w3;
assign w43882 = w438 & w3;
assign w43883 = w329 & w273;
assign w43884 = w488 & ~w42;
assign w43885 = ~w525 & ~w456;
assign w43886 = ~w525 & w39701;
assign w43887 = w530 & ~w456;
assign w43888 = w530 & w39701;
assign w43889 = ~w397 & ~w564;
assign w43890 = ~w330 & w52323;
assign w43891 = ~a[115] & ~w397;
assign w43892 = w515 & w455;
assign w43893 = ~w515 & ~w455;
assign w43894 = ~w512 & w535;
assign w43895 = ~w543 & w510;
assign w43896 = w543 & w544;
assign w43897 = ~w694 & w80;
assign w43898 = ~w697 & ~w643;
assign w43899 = w770 & w3;
assign w43900 = w778 & ~w771;
assign w43901 = ~w39751 & ~w799;
assign w43902 = ~w703 & ~w720;
assign w43903 = ~w703 & ~w39750;
assign w43904 = w825 & ~w57;
assign w43905 = ~w769 & ~w3;
assign w43906 = w748 & w894;
assign w43907 = w876 & w400;
assign w43908 = w893 & ~w878;
assign w43909 = (w936 & ~w748) | (w936 & w50748) | (~w748 & w50748);
assign w43910 = w828 & w940;
assign w43911 = ~w948 & ~w946;
assign w43912 = ~w958 & w834;
assign w43913 = ~w980 & w42;
assign w43914 = w943 & w57;
assign w43915 = w42 & ~w1114;
assign w43916 = ~w983 & w1133;
assign w43917 = w984 & w1152;
assign w43918 = ~w1135 & ~w252;
assign w43919 = ~w983 & w400;
assign w43920 = ~w983 & ~w1096;
assign w43921 = ~w983 & w1086;
assign w43922 = ~w1199 & ~w80;
assign w43923 = ~w983 & ~w1301;
assign w43924 = ~w1312 & ~w1314;
assign w43925 = ~w1312 & w39799;
assign w43926 = ~w1168 & w1327;
assign w43927 = ~w1399 & w1414;
assign w43928 = ~w1415 & w493;
assign w43929 = ~w400 & w351;
assign w43930 = w351 & ~w1314;
assign w43931 = w351 & w39799;
assign w43932 = ~w39820 & w1311;
assign w43933 = w39820 & ~w1311;
assign w43934 = ~w1441 & ~w1462;
assign w43935 = ~w1320 & w46806;
assign w43936 = (w80 & w1320) | (w80 & w46807) | (w1320 & w46807);
assign w43937 = (w57 & w1320) | (w57 & w46808) | (w1320 & w46808);
assign w43938 = ~w1168 & ~w1326;
assign w43939 = (w1486 & w1215) | (w1486 & w46809) | (w1215 & w46809);
assign w43940 = (~w80 & w1215) | (~w80 & w46810) | (w1215 & w46810);
assign w43941 = (~w1212 & w1167) | (~w1212 & w51392) | (w1167 & w51392);
assign w43942 = w1483 & w48282;
assign w43943 = ~w1512 & w1527;
assign w43944 = ~w1530 & ~w1533;
assign w43945 = ~w1536 & ~w1336;
assign w43946 = w1536 & w1538;
assign w43947 = w1528 & ~w1509;
assign w43948 = w1557 & w52324;
assign w43949 = w1591 & w1370;
assign w43950 = ~w1675 & w1676;
assign w43951 = w1675 & w1678;
assign w43952 = ~w1648 & w1681;
assign w43953 = (w1687 & w1509) | (w1687 & w48283) | (w1509 & w48283);
assign w43954 = ~w1509 & w48284;
assign w43955 = ~w1810 & w1320;
assign w43956 = ~w1803 & w1798;
assign w43957 = w1835 & ~w1837;
assign w43958 = ~w1835 & w1837;
assign w43959 = ~w1607 & w1645;
assign w43960 = (~w1671 & ~w1647) | (~w1671 & w46811) | (~w1647 & w46811);
assign w43961 = ~w2014 & w2016;
assign w43962 = w2014 & w2018;
assign w43963 = ~w2036 & ~w2039;
assign w43964 = w2036 & w2039;
assign w43965 = ~w2005 & w2084;
assign w43966 = ~w2005 & ~w2092;
assign w43967 = w1867 & w1948;
assign w43968 = w39914 & w2117;
assign w43969 = (w2117 & w39914) | (w2117 & w2120) | (w39914 & w2120);
assign w43970 = ~w2120 & w39915;
assign w43971 = ~w2005 & w2042;
assign w43972 = w2101 & ~w2133;
assign w43973 = ~w2005 & w2199;
assign w43974 = ~w2135 & w46812;
assign w43975 = ~w2135 & w46813;
assign w43976 = (w1120 & w2135) | (w1120 & w46814) | (w2135 & w46814);
assign w43977 = w2136 & ~w2409;
assign w43978 = ~w2088 & w51393;
assign w43979 = (w2420 & ~w43977) | (w2420 & w46815) | (~w43977 & w46815);
assign w43980 = w43977 & w46816;
assign w43981 = (w612 & w2135) | (w612 & w46817) | (w2135 & w46817);
assign w43982 = ~w2431 & w2434;
assign w43983 = w2431 & w2436;
assign w43984 = w43977 & w46818;
assign w43985 = (w2441 & ~w43977) | (w2441 & w46819) | (~w43977 & w46819);
assign w43986 = w2136 & w2450;
assign w43987 = w43986 & w46820;
assign w43988 = (w2454 & ~w43986) | (w2454 & w46821) | (~w43986 & w46821);
assign w43989 = (~w2451 & ~w43986) | (~w2451 & w46822) | (~w43986 & w46822);
assign w43990 = w43986 & w46823;
assign w43991 = ~w2282 & ~w2127;
assign w43992 = w2484 & w252;
assign w43993 = ~w2285 & w48285;
assign w43994 = ~w2135 & w46824;
assign w43995 = ~w2135 & w46825;
assign w43996 = ~w2135 & w46826;
assign w43997 = (w80 & w2135) | (w80 & w46827) | (w2135 & w46827);
assign w43998 = ~w2528 & w2531;
assign w43999 = w2528 & w2533;
assign w44000 = ~w2528 & w2538;
assign w44001 = w2528 & w2540;
assign w44002 = ~w2517 & w57;
assign w44003 = ~w2496 & w80;
assign w44004 = w2542 & w2535;
assign w44005 = ~w2576 & ~w2578;
assign w44006 = (~w2492 & w51394) | (~w2492 & w51395) | (w51394 & w51395);
assign w44007 = w2591 & ~w2603;
assign w44008 = ~w2591 & w2608;
assign w44009 = ~w2635 & w2633;
assign w44010 = w2638 & ~w2639;
assign w44011 = w2555 & ~w351;
assign w44012 = ~w2686 & w39982;
assign w44013 = w2362 & w2748;
assign w44014 = ~w2362 & ~w2748;
assign w44015 = w2792 & w2789;
assign w44016 = (w2554 & w44015) | (w2554 & w46828) | (w44015 & w46828);
assign w44017 = ~w2792 & ~w2789;
assign w44018 = ~w2792 & w50240;
assign w44019 = ~w2805 & ~w2806;
assign w44020 = (~w2554 & w44019) | (~w2554 & w46829) | (w44019 & w46829);
assign w44021 = (w2808 & w2554) | (w2808 & w48286) | (w2554 & w48286);
assign w44022 = (w2557 & w46830) | (w2557 & w46831) | (w46830 & w46831);
assign w44023 = (~w2557 & w48287) | (~w2557 & w48288) | (w48287 & w48288);
assign w44024 = ~w2822 & w1738;
assign w44025 = w2357 & w2767;
assign w44026 = w2357 & ~w39997;
assign w44027 = ~w1320 & ~w2765;
assign w44028 = ~w1320 & ~w39996;
assign w44029 = w2869 & ~w2646;
assign w44030 = (w2878 & ~w2861) | (w2878 & w48289) | (~w2861 & w48289);
assign w44031 = ~w2626 & w46832;
assign w44032 = w2862 & ~w2671;
assign w44033 = ~w2842 & ~w2848;
assign w44034 = (~w945 & w2987) | (~w945 & w46833) | (w2987 & w46833);
assign w44035 = w2897 & ~w3020;
assign w44036 = (w3032 & w2898) | (w3032 & w46834) | (w2898 & w46834);
assign w44037 = ~w2898 & w46835;
assign w44038 = w3039 & w2795;
assign w44039 = w3044 & ~w1320;
assign w44040 = ~w3030 & w3052;
assign w44041 = (~w3058 & w2898) | (~w3058 & w46836) | (w2898 & w46836);
assign w44042 = (w3060 & ~w2680) | (w3060 & w48290) | (~w2680 & w48290);
assign w44043 = w2897 & w3062;
assign w44044 = ~w3039 & w1320;
assign w44045 = w3055 & w3074;
assign w44046 = ~w2987 & w46837;
assign w44047 = w2862 & w3092;
assign w44048 = (~w3100 & ~w2680) | (~w3100 & w46838) | (~w2680 & w46838);
assign w44049 = w2627 & w3102;
assign w44050 = w2627 & ~w3110;
assign w44051 = ~w3112 & w3113;
assign w44052 = ~w3121 & ~w3125;
assign w44053 = (~w2897 & w46839) | (~w2897 & w46840) | (w46839 & w46840);
assign w44054 = ~w2558 & a[92];
assign w44055 = w2908 & ~w2824;
assign w44056 = w2908 & w3147;
assign w44057 = w2558 & ~a[92];
assign w44058 = w3139 & ~w3138;
assign w44059 = ~w3115 & w3158;
assign w44060 = ~w3115 & ~w3118;
assign w44061 = w3024 & w1738;
assign w44062 = w3190 & ~w3220;
assign w44063 = w3163 & w3221;
assign w44064 = w3223 & ~w2967;
assign w44065 = ~w3334 & ~w3333;
assign w44066 = (w3234 & w3160) | (w3234 & w51396) | (w3160 & w51396);
assign w44067 = ~w3425 & w493;
assign w44068 = w2945 & w48291;
assign w44069 = ~w3532 & w3531;
assign w44070 = ~w40089 & w3580;
assign w44071 = w40090 & w2957;
assign w44072 = ~w3644 & ~w3620;
assign w44073 = w3461 & ~w3648;
assign w44074 = w3461 & w3650;
assign w44075 = ~w3663 & ~w3664;
assign w44076 = w3399 & w48292;
assign w44077 = w3666 & ~w3649;
assign w44078 = w3399 & w48293;
assign w44079 = w3461 & ~w3674;
assign w44080 = ~w3675 & ~w3676;
assign w44081 = w3399 & w48294;
assign w44082 = (w3704 & w3620) | (w3704 & w48295) | (w3620 & w48295);
assign w44083 = w3716 & w3722;
assign w44084 = w3716 & w3718;
assign w44085 = ~w3716 & w3721;
assign w44086 = (w2896 & w3768) | (w2896 & w46841) | (w3768 & w46841);
assign w44087 = ~w3644 & w3798;
assign w44088 = (~w2896 & ~w3620) | (~w2896 & w46842) | (~w3620 & w46842);
assign w44089 = (~w2558 & w3768) | (~w2558 & w46843) | (w3768 & w46843);
assign w44090 = ~w3768 & w46844;
assign w44091 = (w3818 & ~w3620) | (w3818 & w48296) | (~w3620 & w48296);
assign w44092 = w3620 & w48297;
assign w44093 = (~w3369 & w3301) | (~w3369 & w51397) | (w3301 & w51397);
assign w44094 = ~w3620 & w48298;
assign w44095 = ~w3645 & w51398;
assign w44096 = (w3907 & w3620) | (w3907 & w46845) | (w3620 & w46845);
assign w44097 = ~w3620 & w46846;
assign w44098 = ~w3703 & ~w3922;
assign w44099 = w3920 & w3915;
assign w44100 = w3662 & w3638;
assign w44101 = w3810 & w3881;
assign w44102 = w3939 & ~w3938;
assign w44103 = (~w3944 & w3620) | (~w3944 & w48299) | (w3620 & w48299);
assign w44104 = ~w3620 & w48300;
assign w44105 = (w3936 & w46847) | (w3936 & w46848) | (w46847 & w46848);
assign w44106 = ~w3960 & ~w3968;
assign w44107 = (w3983 & w3620) | (w3983 & w46849) | (w3620 & w46849);
assign w44108 = ~w3620 & w46850;
assign w44109 = ~w3968 & ~w3991;
assign w44110 = (w57 & w3620) | (w57 & w46851) | (w3620 & w46851);
assign w44111 = (w4030 & w3620) | (w4030 & w46852) | (w3620 & w46852);
assign w44112 = ~w3620 & w46853;
assign w44113 = ~w3968 & w4038;
assign w44114 = ~w3920 & w4019;
assign w44115 = w40148 & w51399;
assign w44116 = ~w4078 & ~w4077;
assign w44117 = (w4083 & w4051) | (w4083 & w48301) | (w4051 & w48301);
assign w44118 = (w3638 & w4051) | (w3638 & w48302) | (w4051 & w48302);
assign w44119 = (w57 & w4105) | (w57 & w48303) | (w4105 & w48303);
assign w44120 = w4146 & w40157;
assign w44121 = ~w3889 & w4152;
assign w44122 = (~w3904 & w51400) | (~w3904 & w51401) | (w51400 & w51401);
assign w44123 = (~w3737 & w40167) | (~w3737 & w3889) | (w40167 & w3889);
assign w44124 = w3810 & w3880;
assign w44125 = ~w4051 & w48304;
assign w44126 = ~w3889 & ~w3905;
assign w44127 = (w4373 & w4318) | (w4373 & w48305) | (w4318 & w48305);
assign w44128 = ~w4318 & w48306;
assign w44129 = w4211 & ~w4404;
assign w44130 = (w4211 & w4295) | (w4211 & w49330) | (w4295 & w49330);
assign w44131 = ~w4105 & w48307;
assign w44132 = ~w4141 & ~w4407;
assign w44133 = (w3646 & w4406) | (w3646 & w46854) | (w4406 & w46854);
assign w44134 = (w1738 & w4585) | (w1738 & w46855) | (w4585 & w46855);
assign w44135 = w4267 & w2285;
assign w44136 = w4506 & ~w4595;
assign w44137 = ~w4506 & ~w4597;
assign w44138 = ~w4585 & w46856;
assign w44139 = ~w4659 & w46857;
assign w44140 = (w754 & w4659) | (w754 & w46858) | (w4659 & w46858);
assign w44141 = ~w4343 & w46859;
assign w44142 = (w46860 & w46861) | (w46860 & w4343) | (w46861 & w4343);
assign w44143 = (~w42 & w4391) | (~w42 & w48308) | (w4391 & w48308);
assign w44144 = w4446 & w4759;
assign w44145 = (w4808 & w4804) | (w4808 & w46862) | (w4804 & w46862);
assign w44146 = ~w4804 & w46863;
assign w44147 = ~w4804 & w46864;
assign w44148 = (w4826 & w4804) | (w4826 & w46865) | (w4804 & w46865);
assign w44149 = ~w4590 & w40222;
assign w44150 = ~w4590 & ~w4850;
assign w44151 = ~w4860 & w40222;
assign w44152 = ~w4860 & ~w4850;
assign w44153 = ~w4833 & w4978;
assign w44154 = w5062 & w612;
assign w44155 = ~w5154 & w1738;
assign w44156 = ~w5275 & w400;
assign w44157 = ~w5271 & ~w351;
assign w44158 = ~w4955 & w4903;
assign w44159 = w5329 & w4849;
assign w44160 = ~w5329 & ~w5336;
assign w44161 = w5329 & a[79];
assign w44162 = (w5346 & w5329) | (w5346 & w46866) | (w5329 & w46866);
assign w44163 = ~w5329 & w46867;
assign w44164 = w5329 & w5358;
assign w44165 = ~w5329 & w5357;
assign w44166 = (w5362 & w5329) | (w5362 & w46868) | (w5329 & w46868);
assign w44167 = ~w5329 & w46869;
assign w44168 = ~w5329 & ~w4430;
assign w44169 = ~w5329 & ~w5375;
assign w44170 = w5329 & ~w4056;
assign w44171 = ~w5329 & w5004;
assign w44172 = w5329 & w5403;
assign w44173 = ~w5329 & w5407;
assign w44174 = w5329 & w4986;
assign w44175 = ~w5329 & w5416;
assign w44176 = ~w5426 & w4931;
assign w44177 = ~w5426 & w5431;
assign w44178 = w5329 & ~w4947;
assign w44179 = w5329 & w5446;
assign w44180 = w5329 & w5452;
assign w44181 = w5329 & w5457;
assign w44182 = w5329 & w5467;
assign w44183 = ~w5329 & w5469;
assign w44184 = w5329 & w5157;
assign w44185 = ~w4877 & w4868;
assign w44186 = w5484 & ~w5489;
assign w44187 = w5329 & ~w5161;
assign w44188 = (w5328 & w46870) | (w5328 & w46871) | (w46870 & w46871);
assign w44189 = w5164 & w5503;
assign w44190 = w5329 & w5509;
assign w44191 = w1120 & ~w5500;
assign w44192 = ~w5157 & ~w5517;
assign w44193 = w5157 & w5517;
assign w44194 = w5329 & w5150;
assign w44195 = w1320 & ~w5521;
assign w44196 = ~w5329 & w5534;
assign w44197 = w5329 & ~w5537;
assign w44198 = (w5328 & w46872) | (w5328 & w46873) | (w46872 & w46873);
assign w44199 = w5552 & w5102;
assign w44200 = (~w754 & w5330) | (~w754 & w46874) | (w5330 & w46874);
assign w44201 = w5329 & w1120;
assign w44202 = ~w5329 & w5504;
assign w44203 = w5329 & w2558;
assign w44204 = ~w5329 & ~w5430;
assign w44205 = (~w5133 & w5329) | (~w5133 & w49331) | (w5329 & w49331);
assign w44206 = w5128 & ~w5593;
assign w44207 = ~w5596 & w5595;
assign w44208 = w5329 & ~w5132;
assign w44209 = ~w5592 & w49332;
assign w44210 = ~w5607 & ~w5606;
assign w44211 = w40273 & ~w5610;
assign w44212 = w5329 & w5615;
assign w44213 = w5329 & ~w493;
assign w44214 = ~w5622 & w52325;
assign w44215 = (w5328 & w49333) | (w5328 & w49334) | (w49333 & w49334);
assign w44216 = w5329 & w400;
assign w44217 = (w5328 & w49335) | (w5328 & w49336) | (w49335 & w49336);
assign w44218 = ~w5632 & w52326;
assign w44219 = ~w5633 & ~w5631;
assign w44220 = ~w5652 & ~w5278;
assign w44221 = ~w5666 & ~w80;
assign w44222 = ~w5683 & ~w5685;
assign w44223 = ~w5577 & w5720;
assign w44224 = ~w5743 & ~w5886;
assign w44225 = ~w5743 & ~w5901;
assign w44226 = ~w5721 & w52099;
assign w44227 = (w5909 & w5721) | (w5909 & w52100) | (w5721 & w52100);
assign w44228 = (~w4430 & w5721) | (~w4430 & w52101) | (w5721 & w52101);
assign w44229 = ~w5881 & ~w3646;
assign w44230 = ~w6071 & ~w1120;
assign w44231 = w5899 & w6084;
assign w44232 = (w6286 & w48309) | (w6286 & w48310) | (w48309 & w48310);
assign w44233 = (w6297 & ~w6287) | (w6297 & w46876) | (~w6287 & w46876);
assign w44234 = (~w6228 & w6112) | (~w6228 & w48311) | (w6112 & w48311);
assign w44235 = (~w6361 & w6261) | (~w6361 & w49337) | (w6261 & w49337);
assign w44236 = w6263 & ~w6363;
assign w44237 = (w6413 & w6261) | (w6413 & w49338) | (w6261 & w49338);
assign w44238 = ~w6261 & w49339;
assign w44239 = w6420 & w48312;
assign w44240 = (w6436 & w6261) | (w6436 & w49340) | (w6261 & w49340);
assign w44241 = ~w6261 & w49341;
assign w44242 = ~w6433 & ~w6455;
assign w44243 = ~w6429 & w6456;
assign w44244 = w6461 & w6462;
assign w44245 = ~w6461 & w6464;
assign w44246 = w6461 & w6495;
assign w44247 = ~w6461 & w6497;
assign w44248 = ~w6113 & w6687;
assign w44249 = (~w6694 & w6261) | (~w6694 & w49342) | (w6261 & w49342);
assign w44250 = w400 & ~w6695;
assign w44251 = w5962 & w49849;
assign w44252 = ~w6076 & w6237;
assign w44253 = (w6178 & w6261) | (w6178 & w50413) | (w6261 & w50413);
assign w44254 = ~w493 & w52327;
assign w44255 = (w6726 & w6261) | (w6726 & w49343) | (w6261 & w49343);
assign w44256 = w6263 & w6730;
assign w44257 = w493 & ~w6708;
assign w44258 = (w6562 & w6456) | (w6562 & w46877) | (w6456 & w46877);
assign w44259 = ~w6812 & ~w6811;
assign w44260 = ~w6429 & w6443;
assign w44261 = (w6556 & w6456) | (w6556 & w46878) | (w6456 & w46878);
assign w44262 = w7049 & w6318;
assign w44263 = w7049 & w40434;
assign w44264 = ~w6432 & w6318;
assign w44265 = ~w6432 & w40434;
assign w44266 = w7058 & w6318;
assign w44267 = w7058 & w40434;
assign w44268 = ~w7053 & ~w2896;
assign w44269 = (w1541 & w48313) | (w1541 & ~w6769) | (w48313 & ~w6769);
assign w44270 = w7072 & w6318;
assign w44271 = w7072 & w40434;
assign w44272 = w6998 & ~w7069;
assign w44273 = ~w7087 & w6821;
assign w44274 = w7097 & w6318;
assign w44275 = w7097 & w40434;
assign w44276 = w6591 & w6318;
assign w44277 = w6591 & w40434;
assign w44278 = ~w7111 & w754;
assign w44279 = ~w7108 & ~w6592;
assign w44280 = ~w7108 & w7118;
assign w44281 = ~w6578 & w6318;
assign w44282 = ~w6578 & w40434;
assign w44283 = ~w6680 & w6642;
assign w44284 = w252 & w6318;
assign w44285 = w252 & w40434;
assign w44286 = ~w7166 & ~w7165;
assign w44287 = ~w7169 & ~w7168;
assign w44288 = w7170 & w7167;
assign w44289 = w6735 & ~w6711;
assign w44290 = ~w7189 & ~w7190;
assign w44291 = (~w351 & ~w6769) | (~w351 & w49344) | (~w6769 & w49344);
assign w44292 = ~w7196 & w48315;
assign w44293 = (w7199 & w7196) | (w7199 & w48316) | (w7196 & w48316);
assign w44294 = ~w7196 & w48317;
assign w44295 = (w7214 & w7196) | (w7214 & w48318) | (w7196 & w48318);
assign w44296 = (w7142 & w49345) | (w7142 & w49346) | (w49345 & w49346);
assign w44297 = ~w7244 & w7153;
assign w44298 = w6762 & w48319;
assign w44299 = (~w42 & w7249) | (~w42 & w48320) | (w7249 & w48320);
assign w44300 = ~w7179 & w7267;
assign w44301 = ~w6605 & w6318;
assign w44302 = (~w6762 & w44301) | (~w6762 & w48321) | (w44301 & w48321);
assign w44303 = (~w6737 & w50152) | (~w6737 & w50153) | (w50152 & w50153);
assign w44304 = w7111 & ~w754;
assign w44305 = ~w7249 & w48322;
assign w44306 = w7293 & ~w7301;
assign w44307 = w40471 & w6796;
assign w44308 = (~w7082 & w44307) | (~w7082 & w48323) | (w44307 & w48323);
assign w44309 = w7325 & ~w945;
assign w44310 = w7085 & ~w1120;
assign w44311 = ~w7067 & ~w7082;
assign w44312 = (w48324 & w50415) | (w48324 & w44300) | (w50415 & w44300);
assign w44313 = (~w44300 & w48325) | (~w44300 & w48326) | (w48325 & w48326);
assign w44314 = ~w7270 & w50154;
assign w44315 = (~w44300 & w48327) | (~w44300 & w48328) | (w48327 & w48328);
assign w44316 = ~w7416 & ~w7417;
assign w44317 = (~w7082 & w44316) | (~w7082 & w48329) | (w44316 & w48329);
assign w44318 = w7420 & ~w7269;
assign w44319 = w7420 & ~w40484;
assign w44320 = ~w7315 & w49347;
assign w44321 = (~w44300 & w48330) | (~w44300 & w48331) | (w48330 & w48331);
assign w44322 = (~w44300 & w48332) | (~w44300 & w48333) | (w48332 & w48333);
assign w44323 = (~w44300 & w48334) | (~w44300 & w48335) | (w48334 & w48335);
assign w44324 = (~w44300 & w48336) | (~w44300 & w48337) | (w48336 & w48337);
assign w44325 = (~w44300 & w48338) | (~w44300 & w48339) | (w48338 & w48339);
assign w44326 = (~w44300 & w48340) | (~w44300 & w48341) | (w48340 & w48341);
assign w44327 = (~w44300 & w48342) | (~w44300 & w48343) | (w48342 & w48343);
assign w44328 = (~w44300 & w48344) | (~w44300 & w48345) | (w48344 & w48345);
assign w44329 = (~w44300 & w48346) | (~w44300 & w48347) | (w48346 & w48347);
assign w44330 = (~w44300 & w48348) | (~w44300 & w48349) | (w48348 & w48349);
assign w44331 = (~w44300 & w48350) | (~w44300 & w48351) | (w48350 & w48351);
assign w44332 = (~w44300 & w48352) | (~w44300 & w48353) | (w48352 & w48353);
assign w44333 = (w44300 & w48354) | (w44300 & w48355) | (w48354 & w48355);
assign w44334 = w40526 & w7194;
assign w44335 = (~w44300 & w48356) | (~w44300 & w48357) | (w48356 & w48357);
assign w44336 = ~w7839 & ~w7783;
assign w44337 = w7178 & ~w7844;
assign w44338 = w7178 & ~w40537;
assign w44339 = w3 & w52328;
assign w44340 = (~w44300 & w48358) | (~w44300 & w48359) | (w48358 & w48359);
assign w44341 = w7874 & ~w7855;
assign w44342 = w7874 & ~w40538;
assign w44343 = w7901 & w7841;
assign w44344 = w7781 & w7903;
assign w44345 = ~w42 & ~w7908;
assign w44346 = ~w7948 & w46879;
assign w44347 = (~w612 & w7948) | (~w612 & w46880) | (w7948 & w46880);
assign w44348 = w7978 & w50241;
assign w44349 = ~w8035 & w7976;
assign w44350 = ~w8055 & ~w8058;
assign w44351 = w8062 & ~w8064;
assign w44352 = (w252 & w7904) | (w252 & w46881) | (w7904 & w46881);
assign w44353 = (~w7783 & w7452) | (~w7783 & w48360) | (w7452 & w48360);
assign w44354 = ~w7887 & w48361;
assign w44355 = ~w7820 & w7922;
assign w44356 = ~w8090 & w8095;
assign w44357 = w8090 & w8097;
assign w44358 = w7900 & w8105;
assign w44359 = w7900 & w8120;
assign w44360 = w7900 & w8127;
assign w44361 = w7900 & w8134;
assign w44362 = w8050 & w351;
assign w44363 = ~w8291 & ~w8287;
assign w44364 = ~w8291 & ~w40604;
assign w44365 = ~w7887 & w46882;
assign w44366 = w8296 & w7922;
assign w44367 = w8300 & w8297;
assign w44368 = w8300 & w40605;
assign w44369 = ~w8294 & w8302;
assign w44370 = ~w8274 & w8303;
assign w44371 = ~w7562 & w8297;
assign w44372 = ~w7562 & w40605;
assign w44373 = w8333 & ~w8287;
assign w44374 = w8333 & ~w40604;
assign w44375 = w8335 & w8287;
assign w44376 = w8335 & w40604;
assign w44377 = w8360 & ~w8356;
assign w44378 = w8360 & ~w40612;
assign w44379 = w8362 & w8356;
assign w44380 = w8362 & w40612;
assign w44381 = w8381 & w8356;
assign w44382 = w8381 & w40612;
assign w44383 = w8383 & ~w8356;
assign w44384 = w8383 & ~w40612;
assign w44385 = w8347 & ~w4056;
assign w44386 = (~w2896 & ~w8472) | (~w2896 & w48362) | (~w8472 & w48362);
assign w44387 = ~w8617 & w46883;
assign w44388 = ~w8541 & w8577;
assign w44389 = ~w8617 & w46884;
assign w44390 = (w8612 & w8617) | (w8612 & w46885) | (w8617 & w46885);
assign w44391 = w8443 & ~w8520;
assign w44392 = w8650 & w8655;
assign w44393 = ~w8650 & w8657;
assign w44394 = w8650 & w8661;
assign w44395 = ~w8650 & w8663;
assign w44396 = w8390 & ~w8616;
assign w44397 = w8448 & w8479;
assign w44398 = ~w8448 & w8428;
assign w44399 = w8710 & w8709;
assign w44400 = w8710 & w8390;
assign w44401 = ~w8713 & ~w8709;
assign w44402 = ~w8713 & ~w8390;
assign w44403 = ~w8686 & ~w8729;
assign w44404 = w8686 & w8729;
assign w44405 = (~w8391 & ~w8339) | (~w8391 & w50416) | (~w8339 & w50416);
assign w44406 = (~w8391 & ~w8792) | (~w8391 & w50417) | (~w8792 & w50417);
assign w44407 = ~w8388 & ~w8833;
assign w44408 = ~w8184 & w49850;
assign w44409 = ~w8983 & ~w8007;
assign w44410 = w8987 & ~w8007;
assign w44411 = ~w8985 & w46886;
assign w44412 = (~w8982 & w8985) | (~w8982 & w46887) | (w8985 & w46887);
assign w44413 = ~w754 & ~w9001;
assign w44414 = ~w9015 & w8099;
assign w44415 = ~w9015 & w8183;
assign w44416 = ~w8983 & w9029;
assign w44417 = w8987 & w9029;
assign w44418 = (w9033 & w8985) | (w9033 & w46888) | (w8985 & w46888);
assign w44419 = ~w9009 & w9044;
assign w44420 = w9009 & ~w9065;
assign w44421 = (w8983 & ~w9032) | (w8983 & w46889) | (~w9032 & w46889);
assign w44422 = (~w8985 & w52102) | (~w8985 & w52103) | (w52102 & w52103);
assign w44423 = (w9081 & w8985) | (w9081 & w46890) | (w8985 & w46890);
assign w44424 = w9001 & ~w9137;
assign w44425 = ~w8189 & ~w9101;
assign w44426 = w9140 & ~w493;
assign w44427 = ~w9116 & ~w80;
assign w44428 = w9005 & ~w9104;
assign w44429 = w9582 & w9765;
assign w44430 = w9817 & w9826;
assign w44431 = ~w9817 & ~w9826;
assign w44432 = ~w9829 & w9831;
assign w44433 = w9829 & w9833;
assign w44434 = w10007 & ~w10001;
assign w44435 = ~w9829 & w10379;
assign w44436 = w9829 & w10381;
assign w44437 = ~w10414 & w10230;
assign w44438 = ~w10324 & w10294;
assign w44439 = ~w10467 & w10471;
assign w44440 = ~w40851 & w10399;
assign w44441 = w10418 & w493;
assign w44442 = ~w10549 & w10552;
assign w44443 = w10549 & w10554;
assign w44444 = w10549 & w10565;
assign w44445 = ~w10549 & w10567;
assign w44446 = ~w10663 & w10627;
assign w44447 = ~w42 & ~w10669;
assign w44448 = w754 & ~w10362;
assign w44449 = w754 & ~w40884;
assign w44450 = ~w40886 & ~w10687;
assign w44451 = w10418 & w10700;
assign w44452 = w10696 & ~w10701;
assign w44453 = ~w40887 & w10704;
assign w44454 = ~w40887 & w10383;
assign w44455 = w10418 & w10717;
assign w44456 = w10418 & w9822;
assign w44457 = ~w10375 & w10722;
assign w44458 = w10375 & ~w10722;
assign w44459 = w10418 & ~w3242;
assign w44460 = ~w10755 & w10760;
assign w44461 = w10755 & w10762;
assign w44462 = ~w10765 & ~w10389;
assign w44463 = ~w10765 & w40892;
assign w44464 = ~w10755 & ~w10759;
assign w44465 = ~w10725 & ~w10727;
assign w44466 = w10746 & w2006;
assign w44467 = ~w40887 & w10838;
assign w44468 = ~w10705 & ~w9812;
assign w44469 = ~w10023 & ~w9996;
assign w44470 = w10570 & ~w10592;
assign w44471 = w10673 & ~w57;
assign w44472 = ~w11137 & w48363;
assign w44473 = (~w10464 & w11137) | (~w10464 & w48364) | (w11137 & w48364);
assign w44474 = w11152 & ~w40943;
assign w44475 = ~w10673 & w10569;
assign w44476 = ~w40944 & w11161;
assign w44477 = ~w40943 & w10517;
assign w44478 = w10673 & ~w493;
assign w44479 = w11176 & w11179;
assign w44480 = ~w11176 & w11181;
assign w44481 = w11176 & w11190;
assign w44482 = ~w11176 & w11192;
assign w44483 = ~w40943 & w10516;
assign w44484 = ~w40943 & w11198;
assign w44485 = w11345 & ~w11346;
assign w44486 = w11345 & ~w40956;
assign w44487 = w10673 & ~w10790;
assign w44488 = ~w10673 & ~w11349;
assign w44489 = w10824 & w11363;
assign w44490 = w10780 & w11365;
assign w44491 = ~w11370 & ~w2006;
assign w44492 = w11375 & w11374;
assign w44493 = ~w11375 & ~w11374;
assign w44494 = ~w11381 & ~w1738;
assign w44495 = w10672 & ~w2896;
assign w44496 = w10673 & w11407;
assign w44497 = ~w11418 & ~w11419;
assign w44498 = w10673 & ~w11421;
assign w44499 = ~w11137 & w46891;
assign w44500 = w11416 & w11425;
assign w44501 = ~w11416 & ~w11428;
assign w44502 = w10673 & ~w10702;
assign w44503 = ~w11137 & w46892;
assign w44504 = w10686 & ~w10679;
assign w44505 = w11447 & ~w754;
assign w44506 = w10673 & w11461;
assign w44507 = ~w11416 & w11466;
assign w44508 = ~w11416 & w11464;
assign w44509 = ~w11478 & ~w11477;
assign w44510 = w10686 & ~w11480;
assign w44511 = w10686 & w11480;
assign w44512 = ~w10673 & w11305;
assign w44513 = w11504 & w11507;
assign w44514 = ~w11504 & w11509;
assign w44515 = ~w11515 & w11518;
assign w44516 = ~w11547 & ~w11533;
assign w44517 = w10673 & ~w11061;
assign w44518 = ~w10673 & w11558;
assign w44519 = ~w10673 & w11565;
assign w44520 = w11592 & w10993;
assign w44521 = ~w11592 & ~w10993;
assign w44522 = w10645 & ~a[59];
assign w44523 = ~w11604 & w9781;
assign w44524 = ~w9195 & ~w11598;
assign w44525 = (w1541 & w11137) | (w1541 & w46893) | (w11137 & w46893);
assign w44526 = ~w11137 & w48365;
assign w44527 = w10673 & w11727;
assign w44528 = w11371 & w2006;
assign w44529 = w10673 & ~w10779;
assign w44530 = ~w11736 & w2285;
assign w44531 = ~w11743 & ~w11742;
assign w44532 = ~w11447 & w754;
assign w44533 = w11468 & ~w11472;
assign w44534 = ~w11432 & w1320;
assign w44535 = w11204 & w493;
assign w44536 = ~w11765 & ~w11713;
assign w44537 = ~w11748 & w11212;
assign w44538 = ~w11770 & ~w11213;
assign w44539 = ~w11781 & w11785;
assign w44540 = ~w11771 & ~w11148;
assign w44541 = ~w40942 & ~w10463;
assign w44542 = ~w11797 & w11796;
assign w44543 = w11790 & w3;
assign w44544 = w11760 & ~w11713;
assign w44545 = ~w11813 & w11865;
assign w44546 = ~w11869 & w52329;
assign w44547 = (~w11869 & w40984) | (~w11869 & w11813) | (w40984 & w11813);
assign w44548 = ~w11694 & ~w11701;
assign w44549 = w40989 & w11905;
assign w44550 = (w11905 & w40989) | (w11905 & w11813) | (w40989 & w11813);
assign w44551 = w11646 & w8666;
assign w44552 = w40999 & w11946;
assign w44553 = (w11946 & w40999) | (w11946 & w11813) | (w40999 & w11813);
assign w44554 = w41000 & w11949;
assign w44555 = (w11949 & w41000) | (w11949 & w11813) | (w41000 & w11813);
assign w44556 = w41001 & w11954;
assign w44557 = (w11954 & w41001) | (w11954 & w11813) | (w41001 & w11813);
assign w44558 = ~w11947 & w11942;
assign w44559 = w41002 & w11962;
assign w44560 = (w11962 & w41002) | (w11962 & w11813) | (w41002 & w11813);
assign w44561 = w11828 & ~w11965;
assign w44562 = w41006 & w11981;
assign w44563 = (w11981 & w41006) | (w11981 & w11813) | (w41006 & w11813);
assign w44564 = w41008 & ~w11966;
assign w44565 = (~w11966 & w41008) | (~w11966 & w11813) | (w41008 & w11813);
assign w44566 = ~w11982 & ~w9781;
assign w44567 = ~w11963 & ~w10419;
assign w44568 = w41012 & w12023;
assign w44569 = (w12023 & w41012) | (w12023 & w11813) | (w41012 & w11813);
assign w44570 = ~w11985 & w9781;
assign w44571 = w11903 & w11939;
assign w44572 = w11928 & ~w6264;
assign w44573 = ~w11574 & ~w11581;
assign w44574 = ~w11813 & w12086;
assign w44575 = ~w11813 & w12109;
assign w44576 = ~w12076 & ~w12118;
assign w44577 = ~w12076 & ~w12126;
assign w44578 = ~w12120 & w12138;
assign w44579 = ~w11813 & w12140;
assign w44580 = ~w11813 & w12149;
assign w44581 = ~w11813 & w12186;
assign w44582 = ~w11870 & w48366;
assign w44583 = w41038 & ~w11757;
assign w44584 = w41041 | ~w12237;
assign w44585 = (~w12237 & w41041) | (~w12237 & w12218) | (w41041 & w12218);
assign w44586 = (w754 & w11870) | (w754 & w48367) | (w11870 & w48367);
assign w44587 = w41054 & ~w12281;
assign w44588 = ~w41054 & w12281;
assign w44589 = ~w41055 & ~w12292;
assign w44590 = ~w41054 & w12295;
assign w44591 = w2285 & ~w12307;
assign w44592 = (w11332 & w49348) | (w11332 & w49349) | (w49348 & w49349);
assign w44593 = ~w2285 & w12307;
assign w44594 = ~w2285 & w52330;
assign w44595 = w12334 & w12317;
assign w44596 = w12340 & w11358;
assign w44597 = w12340 & w41063;
assign w44598 = w11232 & ~w11869;
assign w44599 = w12364 & w11358;
assign w44600 = w12364 & w41063;
assign w44601 = w11322 & ~w11327;
assign w44602 = ~w12443 & ~w12444;
assign w44603 = ~w12484 & w12485;
assign w44604 = ~w12486 & w12487;
assign w44605 = ~w12484 & ~w11764;
assign w44606 = w12516 & ~w12517;
assign w44607 = ~w12516 & w12517;
assign w44608 = w12463 & ~w612;
assign w44609 = w12240 & ~w754;
assign w44610 = w12602 & w12243;
assign w44611 = w12640 & ~w12669;
assign w44612 = w12615 & w12683;
assign w44613 = ~w12421 & w11902;
assign w44614 = ~w12775 & w6264;
assign w44615 = w12777 & ~w6264;
assign w44616 = ~w12640 & w12202;
assign w44617 = w12640 & w12821;
assign w44618 = ~w12839 & ~w3242;
assign w44619 = w12839 & w12843;
assign w44620 = (~w12393 & w12724) | (~w12393 & w50588) | (w12724 & w50588);
assign w44621 = w12636 & w12584;
assign w44622 = w12839 & ~w12212;
assign w44623 = ~w12886 & ~w12889;
assign w44624 = (w2558 & ~w44623) | (w2558 & w50589) | (~w44623 & w50589);
assign w44625 = w11888 & ~w4430;
assign w44626 = ~w12963 & w12965;
assign w44627 = ~w12640 & w12970;
assign w44628 = ~w12336 & w12998;
assign w44629 = ~w12640 & w754;
assign w44630 = w13028 & w13022;
assign w44631 = ~w13028 & ~w13022;
assign w44632 = w12615 & ~w13038;
assign w44633 = w12640 & w12605;
assign w44634 = w12640 & w13048;
assign w44635 = w12317 & w52331;
assign w44636 = ~w13055 & ~w13057;
assign w44637 = ~w12640 & w12598;
assign w44638 = w12203 & w12412;
assign w44639 = ~w12640 & w12301;
assign w44640 = w13080 & w1320;
assign w44641 = ~w12640 & ~w12598;
assign w44642 = ~w12608 & ~w12591;
assign w44643 = ~w12608 & w13098;
assign w44644 = ~w12640 & w13118;
assign w44645 = ~w12465 & w12441;
assign w44646 = (w13118 & w12581) | (w13118 & w48368) | (w12581 & w48368);
assign w44647 = w12640 & ~w13132;
assign w44648 = ~w12640 & ~w13136;
assign w44649 = ~w13143 & w351;
assign w44650 = ~w12543 & ~w12575;
assign w44651 = w12615 & w3;
assign w44652 = w12534 & ~w12575;
assign w44653 = w13186 & ~w3;
assign w44654 = ~w12574 & ~w3;
assign w44655 = w12616 & ~w12513;
assign w44656 = ~w13221 & ~w13225;
assign w44657 = w12640 & w13231;
assign w44658 = ~w12640 & ~w13238;
assign w44659 = ~w13260 & w13269;
assign w44660 = ~w12640 & w1738;
assign w44661 = w13272 & w13275;
assign w44662 = ~w13272 & w13277;
assign w44663 = ~w13282 & w13285;
assign w44664 = ~w13288 & ~w13289;
assign w44665 = ~w13282 & w13295;
assign w44666 = ~w13297 & ~w13298;
assign w44667 = w44623 & w50591;
assign w44668 = ~w13272 & ~w13274;
assign w44669 = w13272 & w13274;
assign w44670 = ~w13045 & ~w13066;
assign w44671 = ~w13228 & ~w13233;
assign w44672 = w13143 & ~w351;
assign w44673 = ~w13380 & ~w13379;
assign w44674 = ~w13388 & w12805;
assign w44675 = w13388 & ~w12805;
assign w44676 = ~w12700 & w12742;
assign w44677 = w13401 & w13393;
assign w44678 = ~w13401 & ~w13393;
assign w44679 = ~w13432 & w13434;
assign w44680 = w13432 & w13436;
assign w44681 = ~w13442 & w13443;
assign w44682 = w13442 & w13445;
assign w44683 = ~w13432 & w13461;
assign w44684 = ~w13442 & w12708;
assign w44685 = w13442 & ~w12708;
assign w44686 = w13150 & w48369;
assign w44687 = w13256 & w13473;
assign w44688 = ~w12827 & ~w12950;
assign w44689 = w12806 & w13503;
assign w44690 = ~w13504 & w13508;
assign w44691 = w13523 & ~w12800;
assign w44692 = ~w13523 & w12800;
assign w44693 = ~w13538 & ~w12877;
assign w44694 = ~w13560 & w13559;
assign w44695 = w13560 & ~w13559;
assign w44696 = w13570 & w13569;
assign w44697 = ~w13570 & ~w13569;
assign w44698 = w13523 & w13586;
assign w44699 = ~w13523 & w13588;
assign w44700 = w13492 & w48370;
assign w44701 = ~w13599 & w13601;
assign w44702 = w13599 & w13603;
assign w44703 = ~w13493 & ~w12918;
assign w44704 = ~w12984 & w13535;
assign w44705 = a[52] & w13633;
assign w44706 = w13257 & w13636;
assign w44707 = ~w13638 & w48371;
assign w44708 = (w11870 & w13638) | (w11870 & w48372) | (w13638 & w48372);
assign w44709 = a[52] & w13654;
assign w44710 = w13672 & w13673;
assign w44711 = ~w13672 & w13675;
assign w44712 = w13691 & ~w13697;
assign w44713 = ~w13691 & w13699;
assign w44714 = ~w13672 & w12692;
assign w44715 = w13672 & ~w12692;
assign w44716 = ~w13599 & w13724;
assign w44717 = w13599 & w13726;
assign w44718 = (w13088 & w13343) | (w13088 & w48373) | (w13343 & w48373);
assign w44719 = ~w13741 & w13743;
assign w44720 = ~w13744 & w13044;
assign w44721 = ~w13746 & w13748;
assign w44722 = w13749 & ~w13045;
assign w44723 = ~w13755 & ~w13754;
assign w44724 = ~w13034 & ~w13147;
assign w44725 = w13777 & ~w13775;
assign w44726 = ~w13782 & ~w13780;
assign w44727 = w13788 & ~w13775;
assign w44728 = ~w13806 & ~w13805;
assign w44729 = w13810 & ~w493;
assign w44730 = w13861 & w48374;
assign w44731 = w13384 & w46894;
assign w44732 = (~w13896 & w46895) | (~w13896 & ~w13384) | (w46895 & ~w13384);
assign w44733 = ~w13475 & w48375;
assign w44734 = (~w13917 & w13475) | (~w13917 & w48376) | (w13475 & w48376);
assign w44735 = ~w13930 & ~w13933;
assign w44736 = ~w13944 & w13333;
assign w44737 = ~w13944 & w12994;
assign w44738 = ~w13947 & ~w13946;
assign w44739 = ~w13819 & w13949;
assign w44740 = w13958 & ~w13960;
assign w44741 = ~w13958 & w13964;
assign w44742 = ~w1320 & ~w14014;
assign w44743 = ~w14017 & ~w14016;
assign w44744 = w14033 & w14035;
assign w44745 = w14026 & w14037;
assign w44746 = ~w13855 & w13737;
assign w44747 = (~w14031 & w13854) | (~w14031 & w48377) | (w13854 & w48377);
assign w44748 = w13894 & ~w14052;
assign w44749 = ~w14038 & ~w80;
assign w44750 = w14061 & w14065;
assign w44751 = ~w14061 & w14067;
assign w44752 = w14061 & w14070;
assign w44753 = ~w14061 & w14072;
assign w44754 = (~w44745 & w49851) | (~w44745 & w49852) | (w49851 & w49852);
assign w44755 = w14038 & w14094;
assign w44756 = (~w44745 & w49853) | (~w44745 & w49854) | (w49853 & w49854);
assign w44757 = (~w44745 & w49855) | (~w44745 & w49856) | (w49855 & w49856);
assign w44758 = w14038 & ~w14122;
assign w44759 = (~w44745 & w49857) | (~w44745 & w49858) | (w49857 & w49858);
assign w44760 = ~w5745 & w52332;
assign w44761 = (w14025 & w49859) | (w14025 & w49860) | (w49859 & w49860);
assign w44762 = (~w44745 & w49861) | (~w44745 & w49862) | (w49861 & w49862);
assign w44763 = ~w14038 & w14178;
assign w44764 = (~w44745 & w49863) | (~w44745 & w49864) | (w49863 & w49864);
assign w44765 = w14143 & ~w13526;
assign w44766 = ~w14143 & w13526;
assign w44767 = (w14025 & w49865) | (w14025 & w49866) | (w49865 & w49866);
assign w44768 = w14188 & w14213;
assign w44769 = (~w44745 & w49867) | (~w44745 & w49868) | (w49867 & w49868);
assign w44770 = ~w2558 & ~w14221;
assign w44771 = (~w44745 & w49869) | (~w44745 & w49870) | (w49869 & w49870);
assign w44772 = w2285 & ~w14238;
assign w44773 = w13614 & w13728;
assign w44774 = (~w44745 & w49871) | (~w44745 & w49872) | (w49871 & w49872);
assign w44775 = (w14025 & w49873) | (w14025 & w49874) | (w49873 & w49874);
assign w44776 = ~w14038 & ~w13622;
assign w44777 = w14265 & w14266;
assign w44778 = w14265 & ~w41208;
assign w44779 = w14038 & ~w14267;
assign w44780 = ~w14265 & ~w14266;
assign w44781 = ~w14265 & w41208;
assign w44782 = (~w44745 & w49875) | (~w44745 & w49876) | (w49875 & w49876);
assign w44783 = (w14025 & w49877) | (w14025 & w49878) | (w49877 & w49878);
assign w44784 = (~w44745 & w49879) | (~w44745 & w49880) | (w49879 & w49880);
assign w44785 = (w14025 & w49881) | (w14025 & w49882) | (w49881 & w49882);
assign w44786 = ~w3646 & ~w14280;
assign w44787 = w4430 & ~w14197;
assign w44788 = w13855 & w14314;
assign w44789 = ~w14038 & w14344;
assign w44790 = w14038 & w14346;
assign w44791 = ~w14038 & w14353;
assign w44792 = w14038 & w14355;
assign w44793 = w14038 & w14367;
assign w44794 = ~w14038 & w14369;
assign w44795 = w14038 & w14384;
assign w44796 = ~w14038 & w14410;
assign w44797 = w14038 & w14412;
assign w44798 = ~w14038 & w14426;
assign w44799 = w14038 & w14428;
assign w44800 = ~w14421 & w14300;
assign w44801 = w14038 & ~w14442;
assign w44802 = ~w14038 & w1120;
assign w44803 = w14468 & w14472;
assign w44804 = ~w14468 & w14474;
assign w44805 = w14468 & w14479;
assign w44806 = ~w14468 & w14481;
assign w44807 = ~w14038 & w13841;
assign w44808 = w14508 & ~w14505;
assign w44809 = w14508 & ~w41237;
assign w44810 = w14509 & w13937;
assign w44811 = w14509 & ~w41236;
assign w44812 = ~w14038 & ~w13936;
assign w44813 = (~w44745 & w49883) | (~w44745 & w49884) | (w49883 & w49884);
assign w44814 = ~w14542 & ~w1738;
assign w44815 = (w14025 & w49885) | (w14025 & w49886) | (w49885 & w49886);
assign w44816 = (~w44745 & w49887) | (~w44745 & w49888) | (w49887 & w49888);
assign w44817 = w2006 & ~w14560;
assign w44818 = ~w14264 & ~w2896;
assign w44819 = w14221 & w2558;
assign w44820 = ~w14291 & ~w4056;
assign w44821 = ~w14261 & w3242;
assign w44822 = w14238 & ~w2285;
assign w44823 = w14560 & ~w2006;
assign w44824 = w14604 & w14612;
assign w44825 = ~w14604 & ~w14611;
assign w44826 = ~w14038 & ~w13848;
assign w44827 = (~w44745 & w49889) | (~w44745 & w49890) | (w49889 & w49890);
assign w44828 = w14666 & ~w14662;
assign w44829 = (w14025 & w49891) | (w14025 & w49892) | (w49891 & w49892);
assign w44830 = w14672 & ~w14662;
assign w44831 = (w14025 & w49893) | (w14025 & w49894) | (w49893 & w49894);
assign w44832 = (~w44745 & w49895) | (~w44745 & w49896) | (w49895 & w49896);
assign w44833 = (w14025 & w49897) | (w14025 & w49898) | (w49897 & w49898);
assign w44834 = w14684 & ~w14677;
assign w44835 = (w14025 & w49899) | (w14025 & w49900) | (w49899 & w49900);
assign w44836 = w14702 & ~w14677;
assign w44837 = (~w44745 & w49901) | (~w44745 & w49902) | (w49901 & w49902);
assign w44838 = w14720 & w14724;
assign w44839 = ~w14720 & w14726;
assign w44840 = ~w14716 & ~w14074;
assign w44841 = ~w14716 & ~w41261;
assign w44842 = (w14025 & w49903) | (w14025 & w49904) | (w49903 & w49904);
assign w44843 = ~w14743 & ~w14720;
assign w44844 = w14689 & ~w14753;
assign w44845 = w14566 & w14759;
assign w44846 = ~w14764 & w14761;
assign w44847 = w14568 & w41266;
assign w44848 = w41267 & w14767;
assign w44849 = (w14767 & w41267) | (w14767 & ~w14568) | (w41267 & ~w14568);
assign w44850 = w41268 & ~w57;
assign w44851 = (~w57 & w41268) | (~w57 & ~w14568) | (w41268 & ~w14568);
assign w44852 = w41269 & ~w14615;
assign w44853 = (w14439 & w48378) | (w14439 & w48379) | (w48378 & w48379);
assign w44854 = (~w14792 & ~w14761) | (~w14792 & w46896) | (~w14761 & w46896);
assign w44855 = ~w14439 & w48380;
assign w44856 = w41271 & w14670;
assign w44857 = (w14439 & w48381) | (w14439 & w48382) | (w48381 & w48382);
assign w44858 = (w14704 & w14439) | (w14704 & w48383) | (w14439 & w48383);
assign w44859 = w14836 & ~w14840;
assign w44860 = w41273 & ~w14843;
assign w44861 = (~w14843 & w41273) | (~w14843 & ~w14568) | (w41273 & ~w14568);
assign w44862 = w14759 & w14527;
assign w44863 = ~w14872 & ~w14876;
assign w44864 = w14880 & ~w14858;
assign w44865 = ~w14514 & ~w14526;
assign w44866 = w14519 & ~w14526;
assign w44867 = ~w14863 & w14866;
assign w44868 = (w493 & w14887) | (w493 & w46897) | (w14887 & w46897);
assign w44869 = ~w41276 & ~w14516;
assign w44870 = (w14905 & ~w14761) | (w14905 & w48384) | (~w14761 & w48384);
assign w44871 = w14761 & w48385;
assign w44872 = ~w41276 & w14910;
assign w44873 = (w14927 & ~w14761) | (w14927 & w48386) | (~w14761 & w48386);
assign w44874 = w14761 & w48387;
assign w44875 = ~w41276 & w14932;
assign w44876 = (w14947 & ~w14761) | (w14947 & w48388) | (~w14761 & w48388);
assign w44877 = w14950 & ~w14517;
assign w44878 = w14950 & ~w41279;
assign w44879 = w14761 & w48389;
assign w44880 = w14945 & w14960;
assign w44881 = ~w14945 & w14962;
assign w44882 = w14971 & w14900;
assign w44883 = ~w14887 & w46898;
assign w44884 = ~w14771 & w15001;
assign w44885 = w14761 & w46899;
assign w44886 = ~w14438 & ~w14586;
assign w44887 = w14438 & w15022;
assign w44888 = ~w14438 & ~w15022;
assign w44889 = (w1738 & ~w14761) | (w1738 & w48390) | (~w14761 & w48390);
assign w44890 = ~w14421 & w15059;
assign w44891 = w15062 & ~w15065;
assign w44892 = (w2285 & ~w14761) | (w2285 & w48391) | (~w14761 & w48391);
assign w44893 = ~w15062 & ~w2285;
assign w44894 = w15062 & ~w15078;
assign w44895 = ~w14421 & ~w14297;
assign w44896 = w14579 & ~w15091;
assign w44897 = w14579 & ~w15090;
assign w44898 = ~w15112 & ~w15119;
assign w44899 = w15090 & w15133;
assign w44900 = w14766 & w48392;
assign w44901 = (~w3242 & ~w14766) | (~w3242 & w48393) | (~w14766 & w48393);
assign w44902 = ~w15159 & w48394;
assign w44903 = ~w15160 & w15175;
assign w44904 = (~w4430 & ~w14761) | (~w4430 & w46900) | (~w14761 & w46900);
assign w44905 = (w15184 & ~w14761) | (w15184 & w46901) | (~w14761 & w46901);
assign w44906 = (w15204 & w15159) | (w15204 & w48395) | (w15159 & w48395);
assign w44907 = ~w15159 & w48396;
assign w44908 = ~w15159 & w48397;
assign w44909 = (w15224 & ~w14761) | (w15224 & w46902) | (~w14761 & w46902);
assign w44910 = w14761 & w46903;
assign w44911 = ~w14419 & ~w14103;
assign w44912 = ~w15240 & w15242;
assign w44913 = (~w14126 & ~w14761) | (~w14126 & w46904) | (~w14761 & w46904);
assign w44914 = (~w15305 & ~w14761) | (~w15305 & w48398) | (~w14761 & w48398);
assign w44915 = ~w15160 & w14113;
assign w44916 = ~w14765 & w46905;
assign w44917 = ~w15372 & ~w15374;
assign w44918 = w14764 & w15395;
assign w44919 = w14568 & w15404;
assign w44920 = w14763 & w41316;
assign w44921 = w41316 & w50242;
assign w44922 = ~w15377 & w15234;
assign w44923 = w14761 & w46906;
assign w44924 = (~w5745 & ~w14761) | (~w5745 & w48400) | (~w14761 & w48400);
assign w44925 = w14761 & w48401;
assign w44926 = w15102 & ~w15106;
assign w44927 = w41321 & w15608;
assign w44928 = (w14439 & w44927) | (w14439 & w48402) | (w44927 & w48402);
assign w44929 = w41322 & w15605;
assign w44930 = (w14439 & w44929) | (w14439 & w48403) | (w44929 & w48403);
assign w44931 = w15625 & w15538;
assign w44932 = ~w15581 & ~w15648;
assign w44933 = ~w15451 & w15650;
assign w44934 = ~w15511 & w15529;
assign w44935 = w15564 & ~w15551;
assign w44936 = ~w15335 & w15233;
assign w44937 = w15581 & ~w14777;
assign w44938 = (~w15718 & w15678) | (~w15718 & w46907) | (w15678 & w46907);
assign w44939 = (w15719 & w15678) | (w15719 & w46908) | (w15678 & w46908);
assign w44940 = (w15707 & w15678) | (w15707 & w46909) | (w15678 & w46909);
assign w44941 = (w15744 & w15678) | (w15744 & w46910) | (w15678 & w46910);
assign w44942 = ~w15679 & ~w15760;
assign w44943 = ~w15679 & w15762;
assign w44944 = (~w15514 & w15678) | (~w15514 & w46911) | (w15678 & w46911);
assign w44945 = ~w14974 & w15678;
assign w44946 = (~w15374 & w15323) | (~w15374 & w48404) | (w15323 & w48404);
assign w44947 = ~w15663 & w15549;
assign w44948 = ~w15533 & w15296;
assign w44949 = (w15233 & w15311) | (w15233 & w46912) | (w15311 & w46912);
assign w44950 = ~w15663 & w15951;
assign w44951 = (~w15195 & w15678) | (~w15195 & w46913) | (w15678 & w46913);
assign w44952 = (~w3646 & w15678) | (~w3646 & w46914) | (w15678 & w46914);
assign w44953 = ~w15533 & w15232;
assign w44954 = w15533 & w16009;
assign w44955 = (w16016 & w15678) | (w16016 & w46915) | (w15678 & w46915);
assign w44956 = w16056 & ~w15536;
assign w44957 = ~w15679 & ~w16065;
assign w44958 = ~w16086 & ~w15572;
assign w44959 = ~w16086 & w15536;
assign w44960 = ~w15124 & w15580;
assign w44961 = ~w15581 & w16124;
assign w44962 = w15660 & w1738;
assign w44963 = w16154 & ~w1738;
assign w44964 = w15660 & ~w16169;
assign w44965 = ~w15679 & w16152;
assign w44966 = ~w1120 & ~w15620;
assign w44967 = ~w1120 & w15538;
assign w44968 = w1120 & w15620;
assign w44969 = w1120 & ~w15538;
assign w44970 = ~w14925 & w15620;
assign w44971 = ~w14925 & ~w15538;
assign w44972 = w16194 & ~w15620;
assign w44973 = w16194 & w15538;
assign w44974 = ~w15679 & ~w14968;
assign w44975 = ~w16161 & w1541;
assign w44976 = ~w15551 & w16130;
assign w44977 = w15618 & w14966;
assign w44978 = ~w15619 & w46916;
assign w44979 = (w16310 & ~w15536) | (w16310 & w46917) | (~w15536 & w46917);
assign w44980 = w15793 & ~w16320;
assign w44981 = (w400 & w15678) | (w400 & w46918) | (w15678 & w46918);
assign w44982 = w15618 & w16421;
assign w44983 = w15666 & w49350;
assign w44984 = w16490 & w16488;
assign w44985 = w16490 & w15797;
assign w44986 = ~w14776 & w16488;
assign w44987 = ~w14776 & w15797;
assign w44988 = w16500 & ~w16488;
assign w44989 = w16500 & ~w15797;
assign w44990 = ~w16494 & ~w16503;
assign w44991 = w16512 & w48405;
assign w44992 = (~w3 & ~w16512) | (~w3 & w48406) | (~w16512 & w48406);
assign w44993 = ~w16234 & ~w945;
assign w44994 = (~w16234 & w16474) | (~w16234 & w48407) | (w16474 & w48407);
assign w44995 = w16550 & w16234;
assign w44996 = w16623 & ~w754;
assign w44997 = w16629 & w16623;
assign w44998 = w16623 & w754;
assign w44999 = ~w16609 & w16592;
assign w45000 = ~w17374 & w17357;
assign w45001 = ~w2558 & ~w17376;
assign w45002 = (~w45000 & w46920) | (~w45000 & w46921) | (w46920 & w46921);
assign w45003 = w41444 & w48408;
assign w45004 = ~w17778 & ~w17014;
assign w45005 = (~w17819 & w17051) | (~w17819 & w48409) | (w17051 & w48409);
assign w45006 = w17062 & w17829;
assign w45007 = ~w17380 & w17856;
assign w45008 = ~w16968 & ~w17862;
assign w45009 = w16829 & ~w2006;
assign w45010 = w16968 & w17862;
assign w45011 = ~w17872 & w1738;
assign w45012 = w17873 & ~w1738;
assign w45013 = w17379 & ~w17092;
assign w45014 = ~w5330 & ~w17889;
assign w45015 = ~w17921 & w17369;
assign w45016 = ~w17921 & w17942;
assign w45017 = ~w17921 & ~w17368;
assign w45018 = ~w17370 & ~w16825;
assign w45019 = ~w17379 & ~w16578;
assign w45020 = ~w16722 & ~w17643;
assign w45021 = w17984 & w57;
assign w45022 = w18020 & w351;
assign w45023 = w17370 & ~w17920;
assign w45024 = ~w17376 & ~w16680;
assign w45025 = ~w41502 & ~w7924;
assign w45026 = ~w41504 & ~w7315;
assign w45027 = (~w5330 & w18182) | (~w5330 & w48410) | (w18182 & w48410);
assign w45028 = ~w18362 & w5330;
assign w45029 = ~w18182 & w17510;
assign w45030 = ~w18391 & ~w6769;
assign w45031 = ~w18405 & ~w18406;
assign w45032 = ~w18405 & w18409;
assign w45033 = ~w41525 & a[43];
assign w45034 = ~w18461 & w18463;
assign w45035 = ~w17637 & w18470;
assign w45036 = ~w17637 & w41526;
assign w45037 = (~w1541 & w18182) | (~w1541 & w48411) | (w18182 & w48411);
assign w45038 = ~w18182 & ~w1320;
assign w45039 = w18655 & w18660;
assign w45040 = ~w18655 & w18662;
assign w45041 = w18930 & ~w57;
assign w45042 = w18533 & ~w18515;
assign w45043 = w18533 & w18480;
assign w45044 = w18753 & w19055;
assign w45045 = w18837 & ~w19125;
assign w45046 = w18837 & w19132;
assign w45047 = w19129 & w2285;
assign w45048 = ~w19129 & ~w2285;
assign w45049 = ~w18383 & w19222;
assign w45050 = ~w19227 & w19222;
assign w45051 = ~w19039 & w41647;
assign w45052 = ~w19039 & w41648;
assign w45053 = ~w19039 & w19249;
assign w45054 = w19039 & ~w19263;
assign w45055 = ~w19268 & ~w4430;
assign w45056 = ~w19039 & w19306;
assign w45057 = ~w19424 & w18183;
assign w45058 = w19424 & w18920;
assign w45059 = ~w19431 & ~w19432;
assign w45060 = w19020 & w19449;
assign w45061 = ~w41673 & w19458;
assign w45062 = w19503 & ~w19501;
assign w45063 = w19503 & ~w41680;
assign w45064 = w19505 & w19501;
assign w45065 = w19505 & w41680;
assign w45066 = w19511 & ~w19510;
assign w45067 = w19511 & ~w41681;
assign w45068 = w19513 & w19510;
assign w45069 = w19513 & w41681;
assign w45070 = w19520 & ~w19510;
assign w45071 = w19520 & ~w41681;
assign w45072 = w19522 & w19510;
assign w45073 = w19522 & w41681;
assign w45074 = w19525 & ~w19501;
assign w45075 = w19525 & ~w41680;
assign w45076 = w19527 & w19501;
assign w45077 = w19527 & w41680;
assign w45078 = w19530 & ~w19519;
assign w45079 = w19039 & ~w18473;
assign w45080 = ~w19039 & w19593;
assign w45081 = ~w19039 & w19573;
assign w45082 = ~w11138 & ~w19612;
assign w45083 = w19039 & w612;
assign w45084 = ~w19799 & w19801;
assign w45085 = w19799 & w19803;
assign w45086 = ~w19799 & ~w19800;
assign w45087 = w19799 & w19800;
assign w45088 = w19039 & w18933;
assign w45089 = ~w41724 & w3;
assign w45090 = ~w19834 & ~w18918;
assign w45091 = w19293 & ~w19958;
assign w45092 = w20004 & w20006;
assign w45093 = ~w20008 & ~w20011;
assign w45094 = w20008 & w20011;
assign w45095 = ~w20022 & ~w20021;
assign w45096 = ~w20060 & ~w20059;
assign w45097 = ~w1320 & w20071;
assign w45098 = w1320 & w20074;
assign w45099 = w19287 & ~w1120;
assign w45100 = w20073 & ~w20098;
assign w45101 = ~w20004 & ~w20006;
assign w45102 = ~w20136 & w20139;
assign w45103 = w20175 & ~w20180;
assign w45104 = ~w20175 & w20180;
assign w45105 = ~w20175 & w19986;
assign w45106 = ~w20237 & w2896;
assign w45107 = ~w20231 & w19257;
assign w45108 = ~w19625 & ~w19627;
assign w45109 = w20281 & w20284;
assign w45110 = ~w20281 & ~w20284;
assign w45111 = ~w20295 & w20296;
assign w45112 = w20295 & w20298;
assign w45113 = ~w19998 & w20313;
assign w45114 = ~w19998 & w20329;
assign w45115 = w20330 & w20349;
assign w45116 = ~w20330 & w20351;
assign w45117 = ~w20295 & w20356;
assign w45118 = w20295 & w20358;
assign w45119 = w20237 & ~w2896;
assign w45120 = ~w20387 & ~w20241;
assign w45121 = ~w19708 & ~w20493;
assign w45122 = ~w20495 & w20500;
assign w45123 = w20495 & w20501;
assign w45124 = ~w20495 & w20517;
assign w45125 = w20495 & w20519;
assign w45126 = w20495 & w20534;
assign w45127 = ~w20495 & w20536;
assign w45128 = ~w19531 & w20564;
assign w45129 = ~w19708 & ~w20608;
assign w45130 = ~w20610 & w20614;
assign w45131 = w20610 & w20616;
assign w45132 = w20634 & w9195;
assign w45133 = ~w20634 & ~w9195;
assign w45134 = ~w19998 & w20665;
assign w45135 = w20727 & w20729;
assign w45136 = ~w20727 & w20731;
assign w45137 = w20727 & w20755;
assign w45138 = ~w20727 & w20757;
assign w45139 = ~w20263 & w20760;
assign w45140 = ~w20769 & w20773;
assign w45141 = w20787 & ~w20789;
assign w45142 = w20786 & w19918;
assign w45143 = ~w20819 & ~w19970;
assign w45144 = ~w19998 & w20821;
assign w45145 = ~w20819 & w19971;
assign w45146 = w20833 & w20831;
assign w45147 = ~w20833 & ~w20831;
assign w45148 = w20852 & w20857;
assign w45149 = ~w20852 & w20859;
assign w45150 = ~w20787 & w19969;
assign w45151 = w20852 & w20884;
assign w45152 = ~w20852 & w20886;
assign w45153 = ~w20774 & w20765;
assign w45154 = ~w20879 & w20904;
assign w45155 = w20879 & ~w20753;
assign w45156 = ~w20917 & ~w20916;
assign w45157 = w20930 & w20590;
assign w45158 = ~w20930 & ~w20590;
assign w45159 = ~w20953 & ~w20956;
assign w45160 = w20976 & w20551;
assign w45161 = w20990 & w20993;
assign w45162 = w21008 & w21012;
assign w45163 = w21008 & w21027;
assign w45164 = ~w20903 & w21048;
assign w45165 = ~w21105 & w21106;
assign w45166 = w21105 & w21108;
assign w45167 = ~w21122 & w20407;
assign w45168 = w21122 & ~w20407;
assign w45169 = ~w21139 & w21007;
assign w45170 = ~w21186 & w21185;
assign w45171 = ~w21185 & ~w21190;
assign w45172 = w21204 & w20655;
assign w45173 = ~w21208 & ~w20655;
assign w45174 = w21225 & w20599;
assign w45175 = w21225 & w21244;
assign w45176 = w20879 & ~w20287;
assign w45177 = ~w20906 & w48412;
assign w45178 = w21276 & w20277;
assign w45179 = ~w5745 & w21277;
assign w45180 = w21291 & ~w21294;
assign w45181 = ~w21272 & ~w5330;
assign w45182 = w21303 & ~w21273;
assign w45183 = w21308 & ~w21311;
assign w45184 = ~w21325 & ~w21320;
assign w45185 = ~w21334 & ~w21333;
assign w45186 = w21325 & w20369;
assign w45187 = ~w20212 & w21360;
assign w45188 = ~w21362 & w21367;
assign w45189 = ~w21362 & w20107;
assign w45190 = w21376 & ~w945;
assign w45191 = w20781 & w21383;
assign w45192 = ~w20098 & ~w754;
assign w45193 = w21398 & w21404;
assign w45194 = ~w21405 & ~w21408;
assign w45195 = ~w20903 & w754;
assign w45196 = w754 & w20098;
assign w45197 = ~w20903 & ~w20151;
assign w45198 = w21448 & w1320;
assign w45199 = w21477 & ~w21478;
assign w45200 = ~w21479 & w1738;
assign w45201 = ~w20251 & ~w20385;
assign w45202 = w20240 & ~w2558;
assign w45203 = ~w20903 & ~w2285;
assign w45204 = w21536 & w20208;
assign w45205 = ~w20903 & w20209;
assign w45206 = ~w21550 & w21553;
assign w45207 = ~w20895 & ~w20830;
assign w45208 = ~w20903 & ~w20878;
assign w45209 = ~w21614 & ~w21615;
assign w45210 = ~w21613 & ~w20891;
assign w45211 = w21628 & w21631;
assign w45212 = ~w21628 & w21633;
assign w45213 = ~w21612 & w21639;
assign w45214 = ~w21612 & ~w20889;
assign w45215 = w21642 & ~w57;
assign w45216 = w57 & w21652;
assign w45217 = ~w20032 & ~w20770;
assign w45218 = ~w21651 & ~w21675;
assign w45219 = ~w21677 & ~w20225;
assign w45220 = ~w20903 & w21683;
assign w45221 = ~w21693 & ~w493;
assign w45222 = w21676 & w21636;
assign w45223 = w80 & w21710;
assign w45224 = ~w80 & w21713;
assign w45225 = ~w21642 & w57;
assign w45226 = w21741 & w21636;
assign w45227 = ~w21303 & w21338;
assign w45228 = ~w21762 & ~w21763;
assign w45229 = ~w21766 & w3242;
assign w45230 = w21479 & ~w1738;
assign w45231 = ~w21810 & ~w21809;
assign w45232 = w22011 & w21558;
assign w45233 = w21241 & ~w1541;
assign w45234 = ~w22143 & w21780;
assign w45235 = ~w21709 & w22231;
assign w45236 = ~w21709 & w22266;
assign w45237 = w21709 & w22265;
assign w45238 = w22283 & w21131;
assign w45239 = ~w22272 & w22303;
assign w45240 = w21241 & w22352;
assign w45241 = ~w22353 & ~w22354;
assign w45242 = w21241 & ~w22400;
assign w45243 = w21241 & w22442;
assign w45244 = (~w21283 & ~w21708) | (~w21283 & w46922) | (~w21708 & w46922);
assign w45245 = ~w21800 & w46923;
assign w45246 = w21241 & ~w21168;
assign w45247 = ~w22558 & w6769;
assign w45248 = ~w22553 & ~w5330;
assign w45249 = ~w22715 & ~w22717;
assign w45250 = w21709 & w22735;
assign w45251 = ~w21800 & w46924;
assign w45252 = (~w22603 & w21800) | (~w22603 & w46925) | (w21800 & w46925);
assign w45253 = w22754 & w22761;
assign w45254 = ~w22763 & ~w22768;
assign w45255 = w22205 & w22771;
assign w45256 = (w22771 & w45255) | (w22771 & w22769) | (w45255 & w22769);
assign w45257 = ~w22772 & w22773;
assign w45258 = w22473 & ~w10419;
assign w45259 = w22936 & w22937;
assign w45260 = w22936 & w22969;
assign w45261 = ~w22953 & w23209;
assign w45262 = ~w22272 & w23275;
assign w45263 = w23314 & ~w23281;
assign w45264 = ~w23314 & w23281;
assign w45265 = w23346 & w23026;
assign w45266 = ~w42016 & ~w23373;
assign w45267 = w22725 & ~w22726;
assign w45268 = ~w23379 & ~w22638;
assign w45269 = w23384 & ~w2006;
assign w45270 = ~w22764 & w2006;
assign w45271 = w23397 & w23399;
assign w45272 = ~w23397 & w23401;
assign w45273 = w23397 & w23405;
assign w45274 = ~w23397 & w23407;
assign w45275 = w22695 & w23412;
assign w45276 = w22695 & w42020;
assign w45277 = w23378 & ~w23421;
assign w45278 = ~w23378 & w23421;
assign w45279 = ~w23382 & w2006;
assign w45280 = ~w23397 & ~w22079;
assign w45281 = (~w2558 & w23427) | (~w2558 & w3095) | (w23427 & w3095);
assign w45282 = ~w23518 & w48413;
assign w45283 = ~w22763 & w22199;
assign w45284 = ~w23533 & w42028;
assign w45285 = ~w23533 & w42029;
assign w45286 = ~w22767 & w48414;
assign w45287 = ~w23533 & w42030;
assign w45288 = w23521 & w23606;
assign w45289 = ~w23521 & w23608;
assign w45290 = w80 & ~w21915;
assign w45291 = w22205 & w22770;
assign w45292 = (w22770 & w45291) | (w22770 & w22769) | (w45291 & w22769);
assign w45293 = ~w23533 & w42041;
assign w45294 = (w23712 & w22767) | (w23712 & w48415) | (w22767 & w48415);
assign w45295 = ~w22767 & w48416;
assign w45296 = ~w22767 & w48417;
assign w45297 = ~w22767 & w48418;
assign w45298 = (w23734 & w22767) | (w23734 & w48419) | (w22767 & w48419);
assign w45299 = w23741 & ~w23627;
assign w45300 = w23803 & ~w23751;
assign w45301 = ~w23804 & ~w23806;
assign w45302 = ~w23640 & ~w23807;
assign w45303 = ~w23874 & w23877;
assign w45304 = w23874 & w23879;
assign w45305 = w23874 & w23882;
assign w45306 = ~w23874 & w23884;
assign w45307 = w23892 & w23894;
assign w45308 = ~w23892 & w23896;
assign w45309 = w23206 & w14766;
assign w45310 = ~w42047 & w23333;
assign w45311 = ~w23924 & ~w23244;
assign w45312 = w23940 & ~w10419;
assign w45313 = w23966 & w23969;
assign w45314 = ~w23966 & w23971;
assign w45315 = ~w23980 & ~w23307;
assign w45316 = ~w23985 & ~w13384;
assign w45317 = w23985 & w13384;
assign w45318 = w23842 & w23990;
assign w45319 = ~w23741 & w23998;
assign w45320 = w23914 & w46926;
assign w45321 = ~w23892 & ~w23893;
assign w45322 = w23892 & w23893;
assign w45323 = ~w23966 & w24027;
assign w45324 = w23966 & w24029;
assign w45325 = w24021 & ~w24034;
assign w45326 = ~w23842 & w24062;
assign w45327 = w23845 & w24068;
assign w45328 = ~w24069 & w24073;
assign w45329 = w23771 & w24088;
assign w45330 = ~w24092 & ~w24091;
assign w45331 = w24133 & ~w24138;
assign w45332 = ~w24141 & ~w20000;
assign w45333 = w24152 & w23147;
assign w45334 = w24157 & ~w19040;
assign w45335 = w24169 & ~w23153;
assign w45336 = ~w24169 & w23153;
assign w45337 = (~w17380 & w23760) | (~w17380 & w48420) | (w23760 & w48420);
assign w45338 = ~w24190 & ~w24192;
assign w45339 = ~w23842 & w18183;
assign w45340 = (~w24161 & ~w23842) | (~w24161 & w46927) | (~w23842 & w46927);
assign w45341 = ~w24040 & w24035;
assign w45342 = w23050 & ~w23498;
assign w45343 = ~w23596 & ~w23499;
assign w45344 = ~w23370 & w24268;
assign w45345 = ~w23476 & ~w24269;
assign w45346 = (~w23476 & w24268) | (~w23476 & w45345) | (w24268 & w45345);
assign w45347 = w24271 & ~w24267;
assign w45348 = (w24265 & w45347) | (w24265 & w48421) | (w45347 & w48421);
assign w45349 = (~w23488 & w23807) | (~w23488 & w48422) | (w23807 & w48422);
assign w45350 = ~w24335 & w24333;
assign w45351 = ~w24365 & w24367;
assign w45352 = w24365 & w24369;
assign w45353 = w24365 & w24388;
assign w45354 = ~w24365 & w24390;
assign w45355 = ~w23058 & ~w22871;
assign w45356 = ~w24405 & ~w24406;
assign w45357 = w24427 & w24428;
assign w45358 = ~w24427 & w24431;
assign w45359 = ~w24439 & w24441;
assign w45360 = w24439 & w24444;
assign w45361 = w24427 & w24451;
assign w45362 = ~w24427 & w24454;
assign w45363 = ~w23348 & w23361;
assign w45364 = w24467 & w24469;
assign w45365 = ~w24467 & w23362;
assign w45366 = ~w24512 & ~w24513;
assign w45367 = w24512 & w24513;
assign w45368 = ~w24525 & w24528;
assign w45369 = w24525 & w24530;
assign w45370 = w24525 & w24541;
assign w45371 = ~w24525 & w24543;
assign w45372 = w24512 & w24546;
assign w45373 = ~w24512 & w24548;
assign w45374 = ~w24425 & ~w24492;
assign w45375 = w23808 & w24604;
assign w45376 = ~w23808 & w24621;
assign w45377 = w24641 & w24644;
assign w45378 = ~w24641 & w24646;
assign w45379 = w24655 & w24658;
assign w45380 = ~w24655 & w24660;
assign w45381 = ~w24655 & w24668;
assign w45382 = w24655 & w24670;
assign w45383 = ~w24397 & w24699;
assign w45384 = w24641 & w24749;
assign w45385 = ~w24641 & w24751;
assign w45386 = w24594 & w24754;
assign w45387 = ~w24594 & w24756;
assign w45388 = ~w24707 & w24767;
assign w45389 = w23863 & w24833;
assign w45390 = w24557 & ~w24865;
assign w45391 = w24256 & w24038;
assign w45392 = w24870 & ~w24016;
assign w45393 = w42090 | w24909;
assign w45394 = (w24909 & w42090) | (w24909 & ~w24256) | (w42090 & ~w24256);
assign w45395 = w24870 & ~w11138;
assign w45396 = w10419 & w24920;
assign w45397 = w10419 & w42092;
assign w45398 = w24904 & ~w11138;
assign w45399 = w42094 | w23997;
assign w45400 = (w23997 & w42094) | (w23997 & ~w24256) | (w42094 & ~w24256);
assign w45401 = ~w42095 & w24010;
assign w45402 = w24871 & w24942;
assign w45403 = w42097 | ~w23996;
assign w45404 = (w24255 & w45403) | (w24255 & w48423) | (w45403 & w48423);
assign w45405 = ~w24953 & ~w24952;
assign w45406 = ~w42102 & ~w24974;
assign w45407 = (~w24540 & w24034) | (~w24540 & w46928) | (w24034 & w46928);
assign w45408 = ~w24532 & ~w24976;
assign w45409 = ~w24983 & ~w24984;
assign w45410 = ~w24983 & ~w42103;
assign w45411 = w24256 & w42106;
assign w45412 = ~w24871 & w25008;
assign w45413 = (~w7924 & w24901) | (~w7924 & w46929) | (w24901 & w46929);
assign w45414 = ~w24871 & ~w25027;
assign w45415 = (~w9195 & w24901) | (~w9195 & w46930) | (w24901 & w46930);
assign w45416 = ~w24901 & w46931;
assign w45417 = ~w24901 & w46932;
assign w45418 = w24976 & w42115;
assign w45419 = ~w24895 & w24765;
assign w45420 = w24702 & w25197;
assign w45421 = w24702 & ~w25200;
assign w45422 = ~w25210 & ~w25207;
assign w45423 = w24871 & w25218;
assign w45424 = ~w24871 & ~w25220;
assign w45425 = w25240 & ~w25110;
assign w45426 = w25240 & ~w42128;
assign w45427 = ~w42129 & w25245;
assign w45428 = (w24142 & w24865) | (w24142 & w46933) | (w24865 & w46933);
assign w45429 = w25251 & ~w25110;
assign w45430 = w25251 & ~w42128;
assign w45431 = w25253 & w25110;
assign w45432 = w25253 & w42128;
assign w45433 = ~w24178 & w24247;
assign w45434 = ~w24871 & ~w24220;
assign w45435 = w24208 & ~w25279;
assign w45436 = (w24208 & ~w24871) | (w24208 & w45435) | (~w24871 & w45435);
assign w45437 = w24197 & w25289;
assign w45438 = (w24197 & ~w24871) | (w24197 & w45437) | (~w24871 & w45437);
assign w45439 = ~w24197 & ~w25289;
assign w45440 = w24871 & w45439;
assign w45441 = (w14039 & w24901) | (w14039 & w48424) | (w24901 & w48424);
assign w45442 = ~w25332 & w25339;
assign w45443 = w25330 & ~w25341;
assign w45444 = w25330 & ~w42134;
assign w45445 = ~w25330 & w25341;
assign w45446 = ~w25330 & w42134;
assign w45447 = ~w24703 & w25373;
assign w45448 = w1738 & ~w25372;
assign w45449 = (w1738 & w25373) | (w1738 & w45448) | (w25373 & w45448);
assign w45450 = ~w1738 & w25372;
assign w45451 = ~w25373 & w45450;
assign w45452 = w25385 & ~w25388;
assign w45453 = w25377 & ~w1541;
assign w45454 = w25473 & w25476;
assign w45455 = ~w24703 & w24573;
assign w45456 = ~w24575 & w24387;
assign w45457 = ~w24575 & ~w42178;
assign w45458 = ~w24261 & w46934;
assign w45459 = w24871 & w23863;
assign w45460 = ~w42201 & w23862;
assign w45461 = ~w24700 & w24766;
assign w45462 = w25668 & w48425;
assign w45463 = ~w24707 & w24765;
assign w45464 = w25669 & ~w80;
assign w45465 = w25438 & w25712;
assign w45466 = ~w24866 & w25722;
assign w45467 = ~w24871 & ~w24666;
assign w45468 = ~w25753 & w25754;
assign w45469 = ~w25753 & ~w42219;
assign w45470 = ~w24871 & ~w25752;
assign w45471 = ~w25717 & w25770;
assign w45472 = ~w25777 & ~w25720;
assign w45473 = w25072 & ~w6264;
assign w45474 = ~w25507 & w24497;
assign w45475 = ~w25789 & ~w25500;
assign w45476 = ~w25672 & ~w25816;
assign w45477 = ~w25856 & w25801;
assign w45478 = ~w25787 & ~w25779;
assign w45479 = ~w25850 & ~w25670;
assign w45480 = w25850 & w80;
assign w45481 = ~w25880 & w25883;
assign w45482 = w25880 & w25885;
assign w45483 = w25850 & ~w57;
assign w45484 = w25893 & w25894;
assign w45485 = ~w25893 & w25896;
assign w45486 = (~w25783 & w25436) | (~w25783 & w49351) | (w25436 & w49351);
assign w45487 = ~w25456 & w25786;
assign w45488 = ~w25844 & ~w25917;
assign w45489 = ~w25905 & w48426;
assign w45490 = w25893 & w25926;
assign w45491 = ~w25893 & w25928;
assign w45492 = w25880 & w25932;
assign w45493 = ~w25880 & w25934;
assign w45494 = ~w25850 & w612;
assign w45495 = (w45486 & w25785) | (w45486 & w48427) | (w25785 & w48427);
assign w45496 = ~w25850 & ~w25969;
assign w45497 = w25850 & ~w25735;
assign w45498 = (w400 & w25968) | (w400 & w48428) | (w25968 & w48428);
assign w45499 = w25850 & ~w25448;
assign w45500 = ~w25992 & w48429;
assign w45501 = ~w26000 & w612;
assign w45502 = w25850 & ~w26006;
assign w45503 = ~w25850 & w48430;
assign w45504 = (~w26006 & w25850) | (~w26006 & w48431) | (w25850 & w48431);
assign w45505 = w25980 & ~w400;
assign w45506 = (~w351 & w25973) | (~w351 & w49352) | (w25973 & w49352);
assign w45507 = ~w26030 & ~w25947;
assign w45508 = (~w26053 & ~w26051) | (~w26053 & w46935) | (~w26051 & w46935);
assign w45509 = (~w26056 & w25850) | (~w26056 & w48432) | (w25850 & w48432);
assign w45510 = ~w25850 & w25398;
assign w45511 = w26061 & w26049;
assign w45512 = ~w26061 & ~w26049;
assign w45513 = ~w26072 & ~w25945;
assign w45514 = w25315 & ~w24971;
assign w45515 = w26083 & w25050;
assign w45516 = ~w26083 & ~w25050;
assign w45517 = (~w26089 & w25850) | (~w26089 & w49905) | (w25850 & w49905);
assign w45518 = w25850 & w26111;
assign w45519 = w26131 & w26133;
assign w45520 = ~w26131 & w26135;
assign w45521 = w26131 & w26139;
assign w45522 = ~w26131 & w26141;
assign w45523 = ~w25849 & w49906;
assign w45524 = w10419 & ~w26146;
assign w45525 = ~w26150 & w26115;
assign w45526 = w26152 & ~w26087;
assign w45527 = ~w24971 & w50244;
assign w45528 = ~w25849 & w49908;
assign w45529 = w25059 & ~w26079;
assign w45530 = (~w26206 & w25843) | (~w26206 & w49909) | (w25843 & w49909);
assign w45531 = w26180 & ~w26079;
assign w45532 = w26178 & ~w26079;
assign w45533 = (w26217 & w25843) | (w26217 & w49910) | (w25843 & w49910);
assign w45534 = (w25842 & w49911) | (w25842 & w49912) | (w49911 & w49912);
assign w45535 = w26235 & ~w26079;
assign w45536 = w26242 & w26244;
assign w45537 = ~w26242 & w26246;
assign w45538 = w25850 & w14039;
assign w45539 = ~w25850 & w26273;
assign w45540 = ~w26242 & w26288;
assign w45541 = w26242 & w26290;
assign w45542 = ~w25849 & w49913;
assign w45543 = ~w25850 & ~w26299;
assign w45544 = ~w25079 & w25798;
assign w45545 = w42228 & w26320;
assign w45546 = ~w25079 & w25796;
assign w45547 = ~w26348 & ~w26349;
assign w45548 = w25850 & ~w26361;
assign w45549 = w26375 & ~w4056;
assign w45550 = (w26362 & w25843) | (w26362 & w49914) | (w25843 & w49914);
assign w45551 = ~w25079 & w25795;
assign w45552 = w25850 & w26397;
assign w45553 = ~w26375 & w4056;
assign w45554 = w25850 & w26442;
assign w45555 = w23843 & w26447;
assign w45556 = w25840 & a[26];
assign w45557 = w25850 & w24874;
assign w45558 = ~w26493 & ~w26495;
assign w45559 = (w26462 & w48433) | (w26462 & w48434) | (w48433 & w48434);
assign w45560 = ~w25850 & w26506;
assign w45561 = (w26527 & w25850) | (w26527 & w49915) | (w25850 & w49915);
assign w45562 = ~w25850 & w49916;
assign w45563 = (w26542 & w25850) | (w26542 & w49917) | (w25850 & w49917);
assign w45564 = ~w25850 & w49918;
assign w45565 = w25850 & w26553;
assign w45566 = ~w25850 & w26555;
assign w45567 = (w25306 & w25850) | (w25306 & w48435) | (w25850 & w48435);
assign w45568 = ~w25850 & w48436;
assign w45569 = ~w25849 & w49919;
assign w45570 = ~w25850 & w26577;
assign w45571 = w25850 & w26594;
assign w45572 = ~w25850 & w26596;
assign w45573 = (~w26541 & w25850) | (~w26541 & w49920) | (w25850 & w49920);
assign w45574 = ~w26628 & ~w26627;
assign w45575 = ~w26639 & w25101;
assign w45576 = ~w25850 & w26645;
assign w45577 = ~w25849 & w48437;
assign w45578 = (w25842 & w48438) | (w25842 & w48439) | (w48438 & w48439);
assign w45579 = w26665 & w26593;
assign w45580 = ~w26565 & w26667;
assign w45581 = w25850 & w26672;
assign w45582 = w25850 & w26676;
assign w45583 = ~w25850 & w26678;
assign w45584 = w26265 & ~w26704;
assign w45585 = ~w25856 & w26051;
assign w45586 = ~w25849 & w49921;
assign w45587 = (~w25842 & w46936) | (~w25842 & w46937) | (w46936 & w46937);
assign w45588 = (w25842 & w46938) | (w25842 & w46939) | (w46938 & w46939);
assign w45589 = (~w25426 & w25849) | (~w25426 & w49922) | (w25849 & w49922);
assign w45590 = (~w25434 & w25849) | (~w25434 & w49923) | (w25849 & w49923);
assign w45591 = w42228 & ~w26763;
assign w45592 = ~w25796 & ~w26763;
assign w45593 = ~w26766 & ~w26765;
assign w45594 = w26776 & ~w2285;
assign w45595 = ~w25849 & w49924;
assign w45596 = (~w25621 & w25843) | (~w25621 & w49925) | (w25843 & w49925);
assign w45597 = w26722 & w26825;
assign w45598 = w26728 & w26834;
assign w45599 = ~w26728 & w26836;
assign w45600 = ~w26878 & ~w26078;
assign w45601 = ~w26876 & w26066;
assign w45602 = w26707 & w26884;
assign w45603 = w26439 & w48440;
assign w45604 = (w493 & ~w26886) | (w493 & w48441) | (~w26886 & w48441);
assign w45605 = w26707 & ~w26930;
assign w45606 = w26722 & w26824;
assign w45607 = (~w26958 & w26078) | (~w26958 & w49926) | (w26078 & w49926);
assign w45608 = (w26070 & w50155) | (w26070 & w50156) | (w50155 & w50156);
assign w45609 = w26977 & ~w26906;
assign w45610 = (w26827 & w48442) | (w26827 & w48443) | (w48442 & w48443);
assign w45611 = (w26957 & w48444) | (w26957 & w48445) | (w48444 & w48445);
assign w45612 = (~w26827 & w48446) | (~w26827 & w48447) | (w48446 & w48447);
assign w45613 = w26707 & ~w27062;
assign w45614 = (~w27063 & w48448) | (~w27063 & w48449) | (w48448 & w48449);
assign w45615 = (w3646 & w26078) | (w3646 & w46940) | (w26078 & w46940);
assign w45616 = (~w4056 & ~w27111) | (~w4056 & w46941) | (~w27111 & w46941);
assign w45617 = w27111 & w46942;
assign w45618 = (w4056 & w26078) | (w4056 & w46943) | (w26078 & w46943);
assign w45619 = w27145 & w48450;
assign w45620 = w27145 & w48451;
assign w45621 = ~w26429 & w26357;
assign w45622 = w27180 & w27184;
assign w45623 = (w27180 & ~w26700) | (w27180 & w49927) | (~w26700 & w49927);
assign w45624 = ~w27180 & ~w27184;
assign w45625 = w26700 & w49928;
assign w45626 = (~w26827 & w48452) | (~w26827 & w48453) | (w48452 & w48453);
assign w45627 = w27246 & w27251;
assign w45628 = (w26070 & w46944) | (w26070 & w46945) | (w46944 & w46945);
assign w45629 = ~w26521 & w27364;
assign w45630 = (~w26070 & w49929) | (~w26070 & w49930) | (w49929 & w49930);
assign w45631 = ~w27448 & ~w19040;
assign w45632 = ~w26708 & w48454;
assign w45633 = ~w27511 & ~w11870;
assign w45634 = ~w26151 & w26115;
assign w45635 = w27657 & w27665;
assign w45636 = (w8666 & w27661) | (w8666 & w49931) | (w27661 & w49931);
assign w45637 = ~w26073 & ~w26148;
assign w45638 = w27677 & w27672;
assign w45639 = w26964 & ~w27686;
assign w45640 = (~w45639 & w48455) | (~w45639 & w48456) | (w48455 & w48456);
assign w45641 = w26177 & ~w27693;
assign w45642 = ~w26177 & w27693;
assign w45643 = ~w26151 & w26114;
assign w45644 = (~w9195 & w26078) | (~w9195 & w49932) | (w26078 & w49932);
assign w45645 = w26152 & w42314;
assign w45646 = ~w27717 & w26292;
assign w45647 = w26138 & w27726;
assign w45648 = ~w26861 & w48457;
assign w45649 = w27808 & ~w27792;
assign w45650 = ~w26073 & w26263;
assign w45651 = w26264 & w27789;
assign w45652 = w26264 & ~w42324;
assign w45653 = w26964 & ~w27826;
assign w45654 = ~w27824 & ~w5745;
assign w45655 = ~w27812 & w27838;
assign w45656 = w27812 & w27841;
assign w45657 = (~w7315 & w26078) | (~w7315 & w49933) | (w26078 & w49933);
assign w45658 = ~w27659 & ~w8666;
assign w45659 = w27662 & w27701;
assign w45660 = ~w27859 & w27857;
assign w45661 = w27687 & ~w9781;
assign w45662 = (w25899 & w26892) | (w25899 & w49934) | (w26892 & w49934);
assign w45663 = (w25899 & ~w26439) | (w25899 & w48458) | (~w26439 & w48458);
assign w45664 = (w25898 & w26892) | (w25898 & w49935) | (w26892 & w49935);
assign w45665 = (w25898 & ~w26439) | (w25898 & w48459) | (~w26439 & w48459);
assign w45666 = w26877 & ~w25947;
assign w45667 = ~w42332 & w27930;
assign w45668 = (w26070 & w49936) | (w26070 & w49937) | (w49936 & w49937);
assign w45669 = ~w26861 & w48460;
assign w45670 = ~w26861 & w48461;
assign w45671 = ~w27956 & ~w26021;
assign w45672 = w27978 & ~w252;
assign w45673 = ~w27956 & w27981;
assign w45674 = ~w27987 & w27990;
assign w45675 = w27987 & w27993;
assign w45676 = ~w27929 & ~w42332;
assign w45677 = w28004 & ~w42332;
assign w45678 = (~w26885 & w48462) | (~w26885 & w48463) | (w48462 & w48463);
assign w45679 = w26880 & w49938;
assign w45680 = (w28022 & ~w26880) | (w28022 & w48464) | (~w26880 & w48464);
assign w45681 = ~w28017 & w28026;
assign w45682 = ~w28036 & w28039;
assign w45683 = w27873 & w27651;
assign w45684 = w27873 & ~w27487;
assign w45685 = w27837 & ~w27880;
assign w45686 = w27868 & ~w27723;
assign w45687 = w28065 & ~w28050;
assign w45688 = w28113 & w28039;
assign w45689 = w26978 & w50245;
assign w45690 = ~w28050 & w46946;
assign w45691 = ~w28050 & w46947;
assign w45692 = (w28076 & w50157) | (w28076 & w50158) | (w50157 & w50158);
assign w45693 = (~w24874 & w28050) | (~w24874 & w46948) | (w28050 & w46948);
assign w45694 = ~w28171 & w28170;
assign w45695 = (~w28049 & w50159) | (~w28049 & w50160) | (w50159 & w50160);
assign w45696 = (~w28076 & w50161) | (~w28076 & w50162) | (w50161 & w50162);
assign w45697 = (w28049 & w50163) | (w28049 & w50164) | (w50163 & w50164);
assign w45698 = (~w27636 & w27483) | (~w27636 & w46949) | (w27483 & w46949);
assign w45699 = ~w15681 & ~w28457;
assign w45700 = w15681 & ~w28456;
assign w45701 = w15681 & w28076;
assign w45702 = w28479 & w28426;
assign w45703 = ~w27873 & w48465;
assign w45704 = (w28508 & w27487) | (w28508 & w48466) | (w27487 & w48466);
assign w45705 = ~w27873 & w48467;
assign w45706 = (~w27880 & w27487) | (~w27880 & w48468) | (w27487 & w48468);
assign w45707 = w27006 & w48469;
assign w45708 = w28716 & w351;
assign w45709 = (w28701 & w28766) | (w28701 & w49940) | (w28766 & w49940);
assign w45710 = ~w27252 & w46950;
assign w45711 = w27084 & w28958;
assign w45712 = w28050 & w27211;
assign w45713 = w28979 & ~w1738;
assign w45714 = w27084 & w27026;
assign w45715 = ~w28979 & w1738;
assign w45716 = ~w27178 & w27206;
assign w45717 = w29019 & ~w29011;
assign w45718 = (~w27191 & ~w29020) | (~w27191 & w48470) | (~w29020 & w48470);
assign w45719 = w29022 & w48471;
assign w45720 = ~w29036 & ~w2006;
assign w45721 = ~w29010 & ~w29018;
assign w45722 = ~w29021 & ~w29042;
assign w45723 = w27949 & ~w4430;
assign w45724 = ~w28050 & w29096;
assign w45725 = w29105 & w29104;
assign w45726 = ~w29105 & ~w29104;
assign w45727 = w28050 & w29111;
assign w45728 = ~w29112 & ~w3646;
assign w45729 = w29112 & w3646;
assign w45730 = w28935 & w28852;
assign w45731 = ~w28763 & ~w29161;
assign w45732 = ~w29157 & w29171;
assign w45733 = ~w29166 & w29170;
assign w45734 = ~w29157 & ~w28743;
assign w45735 = w29166 & ~w29170;
assign w45736 = w29157 & ~w29196;
assign w45737 = w28218 & ~w29205;
assign w45738 = ~w28218 & w29205;
assign w45739 = ~w29157 & w29217;
assign w45740 = w29157 & w29219;
assign w45741 = w29226 & ~w28150;
assign w45742 = ~w29226 & ~w28190;
assign w45743 = ~w29157 & w29243;
assign w45744 = ~w29157 & ~w28281;
assign w45745 = w29157 & w29272;
assign w45746 = ~w29157 & w12666;
assign w45747 = w29157 & w29280;
assign w45748 = w28291 & ~w28473;
assign w45749 = ~w29157 & w29309;
assign w45750 = ~w29157 & w29317;
assign w45751 = w29188 & w29339;
assign w45752 = ~w29188 & w29341;
assign w45753 = w28284 & w16559;
assign w45754 = w29157 & w29385;
assign w45755 = ~w29157 & ~w29394;
assign w45756 = w29157 & w29396;
assign w45757 = ~w29163 & w29142;
assign w45758 = ~w29411 & w26880;
assign w45759 = w28681 & ~w29142;
assign w45760 = w29157 & w29441;
assign w45761 = w29157 & ~w29450;
assign w45762 = w29157 & w29459;
assign w45763 = w29157 & w29505;
assign w45764 = w28498 & ~w29522;
assign w45765 = ~w29529 & ~w29528;
assign w45766 = ~w29157 & ~w28629;
assign w45767 = (w28677 & w28499) | (w28677 & w46951) | (w28499 & w46951);
assign w45768 = ~w29540 & ~w29541;
assign w45769 = ~w28500 & w28675;
assign w45770 = ~w29157 & ~w28645;
assign w45771 = w29552 & w7924;
assign w45772 = w29157 & ~w29557;
assign w45773 = ~w29157 & w28384;
assign w45774 = ~w29586 & w9195;
assign w45775 = w29534 & ~w7315;
assign w45776 = ~w29552 & ~w7924;
assign w45777 = ~w29595 & w29598;
assign w45778 = ~w29602 & w28326;
assign w45779 = w29602 & ~w28326;
assign w45780 = ~w29157 & ~w11870;
assign w45781 = w29157 & w29608;
assign w45782 = ~w29630 & ~w29631;
assign w45783 = w29368 & w29635;
assign w45784 = ~w29157 & w29648;
assign w45785 = (w29363 & w29287) | (w29363 & w46952) | (w29287 & w46952);
assign w45786 = ~w29540 & ~w28623;
assign w45787 = w29665 & ~w29675;
assign w45788 = w28667 & w28556;
assign w45789 = w29682 & ~w28546;
assign w45790 = w29679 & w29693;
assign w45791 = ~w29679 & w29695;
assign w45792 = ~w29682 & w29707;
assign w45793 = w29727 & ~w29742;
assign w45794 = ~w29727 & w29742;
assign w45795 = ~w29157 & w28587;
assign w45796 = w28500 & ~w29683;
assign w45797 = w28668 & w29148;
assign w45798 = w29773 & w29766;
assign w45799 = ~w29775 & w29772;
assign w45800 = w29775 & ~w29772;
assign w45801 = ~w29774 & w29786;
assign w45802 = ~w29157 & w29790;
assign w45803 = ~w28681 & ~w29103;
assign w45804 = w29806 & ~w3242;
assign w45805 = ~w29810 & ~w29811;
assign w45806 = ~w29157 & w29132;
assign w45807 = w29773 & w29090;
assign w45808 = ~w29825 & w29827;
assign w45809 = ~w29157 & w1541;
assign w45810 = w29829 & w29824;
assign w45811 = ~w29829 & ~w29824;
assign w45812 = ~w29825 & w29837;
assign w45813 = ~w29157 & w1320;
assign w45814 = w29840 & w29836;
assign w45815 = w29848 & ~w29850;
assign w45816 = ~w29848 & w29850;
assign w45817 = ~w29157 & ~w28981;
assign w45818 = w29829 & w29858;
assign w45819 = ~w29829 & w29860;
assign w45820 = w29773 & w29084;
assign w45821 = w29865 & w1738;
assign w45822 = w29884 & ~w29887;
assign w45823 = ~w29884 & w29887;
assign w45824 = ~w29890 & w29046;
assign w45825 = w29890 & ~w29046;
assign w45826 = ~w29157 & w28780;
assign w45827 = ~w29006 & ~w28795;
assign w45828 = ~w29904 & ~w29908;
assign w45829 = w29911 & ~w29902;
assign w45830 = w28930 & ~w945;
assign w45831 = ~w29922 & ~w754;
assign w45832 = ~w29825 & w29932;
assign w45833 = ~w29157 & ~w1120;
assign w45834 = ~w29936 & w29939;
assign w45835 = w29936 & w29941;
assign w45836 = ~w29936 & ~w29938;
assign w45837 = w29936 & w29938;
assign w45838 = ~w29967 & w29970;
assign w45839 = w29971 & ~w29972;
assign w45840 = ~w29157 & w29974;
assign w45841 = w29006 & w29965;
assign w45842 = w29982 & w29991;
assign w45843 = ~w29998 & w30004;
assign w45844 = ~w29157 & ~w30011;
assign w45845 = w29982 & w30018;
assign w45846 = w30007 & ~w30012;
assign w45847 = ~w29890 & w30208;
assign w45848 = ~w30222 & w2558;
assign w45849 = w42463 | w29997;
assign w45850 = (w29997 & w42463) | (w29997 & w29960) | (w42463 & w29960);
assign w45851 = w30239 & w46953;
assign w45852 = (w30265 & ~w30239) | (w30265 & w46954) | (~w30239 & w46954);
assign w45853 = (~w30262 & ~w30239) | (~w30262 & w46955) | (~w30239 & w46955);
assign w45854 = w30239 & w46956;
assign w45855 = (w28077 & w30147) | (w28077 & w48472) | (w30147 & w48472);
assign w45856 = w30703 & w20906;
assign w45857 = ~w30703 & ~w20906;
assign w45858 = ~w30764 & ~w17380;
assign w45859 = w30796 & w11138;
assign w45860 = w30821 & ~w12666;
assign w45861 = w30933 & w30917;
assign w45862 = ~w29588 & ~w30957;
assign w45863 = ~w29588 & ~w42523;
assign w45864 = ~w30959 & w29569;
assign w45865 = ~w30959 & ~w30971;
assign w45866 = w9195 & ~w30238;
assign w45867 = w9195 & w29677;
assign w45868 = w30978 & w30981;
assign w45869 = ~w30978 & w30983;
assign w45870 = ~w30988 & ~w30987;
assign w45871 = ~w30988 & ~w42524;
assign w45872 = w30990 & ~w29617;
assign w45873 = w30990 & ~w42525;
assign w45874 = ~w30992 & w29626;
assign w45875 = w30976 & w30994;
assign w45876 = w30978 & w31033;
assign w45877 = ~w30978 & w31035;
assign w45878 = ~w31038 & w30986;
assign w45879 = w29368 & w31147;
assign w45880 = w29665 & w31146;
assign w45881 = ~w29665 & ~w31146;
assign w45882 = w29665 & w31158;
assign w45883 = w31177 & w46957;
assign w45884 = ~w31178 & ~w31182;
assign w45885 = ~w31222 & ~w31225;
assign w45886 = w30239 & w46958;
assign w45887 = (w31236 & ~w30239) | (w31236 & w46959) | (~w30239 & w46959);
assign w45888 = w30239 & w46960;
assign w45889 = (w31370 & ~w30239) | (w31370 & w46961) | (~w30239 & w46961);
assign w45890 = ~w42579 & w31376;
assign w45891 = (~w31233 & ~w30239) | (~w31233 & w46962) | (~w30239 & w46962);
assign w45892 = w30239 & w46963;
assign w45893 = w31253 & w31389;
assign w45894 = (w31391 & ~w30239) | (w31391 & w46964) | (~w30239 & w46964);
assign w45895 = w31039 & w30968;
assign w45896 = w31443 & w31436;
assign w45897 = ~w31403 & w31191;
assign w45898 = ~w32135 & w32138;
assign w45899 = ~w32135 & w32137;
assign w45900 = ~w32183 & w32137;
assign w45901 = ~w32183 & w45899;
assign w45902 = w32186 & w3646;
assign w45903 = ~w32164 & w31334;
assign w45904 = ~w32206 & ~w32207;
assign w45905 = w32212 & ~w2285;
assign w45906 = ~w32206 & w31307;
assign w45907 = w32181 & ~w32236;
assign w45908 = w30997 & ~w31032;
assign w45909 = ~w31217 & w31415;
assign w45910 = w32260 & w32375;
assign w45911 = w31539 & w31518;
assign w45912 = ~w32465 & w32473;
assign w45913 = w32465 & w32475;
assign w45914 = ~w612 & w32480;
assign w45915 = w612 & w32483;
assign w45916 = ~w493 & w32489;
assign w45917 = w493 & w32492;
assign w45918 = w32465 & w32511;
assign w45919 = ~w32465 & w32513;
assign w45920 = w32538 & w945;
assign w45921 = ~w32545 & ~w31494;
assign w45922 = ~w32549 & w31229;
assign w45923 = w32556 & w32559;
assign w45924 = ~w32556 & w32561;
assign w45925 = w32556 & w32591;
assign w45926 = ~w32556 & w32593;
assign w45927 = ~w32610 & w46965;
assign w45928 = ~w32610 & w46966;
assign w45929 = ~w31491 & ~w32644;
assign w45930 = ~w32645 & ~w32646;
assign w45931 = ~w3 & w32667;
assign w45932 = ~w32698 & w46967;
assign w45933 = (~w32621 & w32698) | (~w32621 & w46968) | (w32698 & w46968);
assign w45934 = w32573 & ~w32479;
assign w45935 = ~w32488 & w32515;
assign w45936 = ~w32749 & ~w57;
assign w45937 = w32762 & w32462;
assign w45938 = ~w32762 & w32804;
assign w45939 = w32762 & w32809;
assign w45940 = ~w32762 & w32811;
assign w45941 = w32376 & w32589;
assign w45942 = ~w42653 & w32589;
assign w45943 = ~w32817 & w32571;
assign w45944 = ~w32814 & ~w32583;
assign w45945 = ~w32192 & w32202;
assign w45946 = ~w32424 & w32239;
assign w45947 = w32887 & ~w2006;
assign w45948 = ~w32887 & w2006;
assign w45949 = ~w32428 & ~w32544;
assign w45950 = ~w32901 & ~w1541;
assign w45951 = w32905 & w32907;
assign w45952 = ~w32905 & w32909;
assign w45953 = ~w32888 & ~w32890;
assign w45954 = w32891 & w1738;
assign w45955 = ~w32923 & ~w32922;
assign w45956 = ~w32372 & ~w2285;
assign w45957 = w32921 & w32237;
assign w45958 = ~w2558 & w32940;
assign w45959 = ~w1541 & w32911;
assign w45960 = ~w32698 & w49353;
assign w45961 = w612 & w32813;
assign w45962 = ~w32720 & ~w32710;
assign w45963 = ~w32688 & w33009;
assign w45964 = ~w33010 & w33014;
assign w45965 = ~w33050 & ~w30239;
assign w45966 = ~w32025 & ~w26880;
assign w45967 = w33106 & w32031;
assign w45968 = ~w33106 & ~w32031;
assign w45969 = ~w33135 & w33137;
assign w45970 = w33135 & w33139;
assign w45971 = w33135 & w33194;
assign w45972 = ~w33135 & w33196;
assign w45973 = ~w33168 & w33232;
assign w45974 = w33275 & ~w33290;
assign w45975 = w33268 & w15681;
assign w45976 = ~w33268 & ~w33339;
assign w45977 = ~w32688 & w31668;
assign w45978 = ~w33346 & ~w33349;
assign w45979 = ~w31703 & w31697;
assign w45980 = ~w33313 & w33380;
assign w45981 = ~w33385 & ~w33388;
assign w45982 = w33385 & w33388;
assign w45983 = ~w33313 & w31601;
assign w45984 = ~w32409 & w33412;
assign w45985 = ~w5745 & w32422;
assign w45986 = w5745 & ~w32422;
assign w45987 = (w32323 & w33414) | (w32323 & w46969) | (w33414 & w46969);
assign w45988 = ~w32409 & w33411;
assign w45989 = ~w33432 & ~w33433;
assign w45990 = ~w33441 & ~w33440;
assign w45991 = ~w33443 & ~w33444;
assign w45992 = ~w32404 & ~w33472;
assign w45993 = w32404 & w32279;
assign w45994 = ~w32404 & ~w8666;
assign w45995 = w33475 & w7924;
assign w45996 = w33486 & ~w33489;
assign w45997 = ~w33486 & w33489;
assign w45998 = ~w33492 & w33493;
assign w45999 = w33492 & w33495;
assign w46000 = w33385 & w33501;
assign w46001 = ~w33385 & w33503;
assign w46002 = ~w31576 & ~w33512;
assign w46003 = w31576 & w33512;
assign w46004 = w33311 & w33525;
assign w46005 = ~w33313 & w33540;
assign w46006 = (~w33563 & w32698) | (~w33563 & w46970) | (w32698 & w46970);
assign w46007 = ~w32698 & w46971;
assign w46008 = (~w33569 & ~w33568) | (~w33569 & w46972) | (~w33568 & w46972);
assign w46009 = ~w3242 & w33571;
assign w46010 = w33574 & ~w32146;
assign w46011 = ~w32182 & ~w33570;
assign w46012 = ~w32182 & w33570;
assign w46013 = ~w33568 & w33601;
assign w46014 = (~w33603 & ~w33568) | (~w33603 & w46973) | (~w33568 & w46973);
assign w46015 = w33605 & ~w33606;
assign w46016 = ~w33605 & w33606;
assign w46017 = ~w33584 & w46974;
assign w46018 = ~w32921 & ~w32128;
assign w46019 = ~w32129 & ~w4430;
assign w46020 = w33605 & w33623;
assign w46021 = ~w33605 & w33625;
assign w46022 = ~w33479 & ~w33481;
assign w46023 = ~w33475 & ~w7924;
assign w46024 = w33492 & ~w33661;
assign w46025 = ~w33492 & w33661;
assign w46026 = ~w33414 & w46975;
assign w46027 = (w33672 & w33414) | (w33672 & w46976) | (w33414 & w46976);
assign w46028 = w33693 & w33631;
assign w46029 = ~w33556 & w33696;
assign w46030 = ~w33616 & ~w33618;
assign w46031 = w33574 & w33712;
assign w46032 = ~w33574 & w33714;
assign w46033 = ~w2285 & ~w33724;
assign w46034 = (w32995 & ~w32994) | (w32995 & w46977) | (~w32994 & w46977);
assign w46035 = w32977 & w32830;
assign w46036 = ~w42686 & w33798;
assign w46037 = w42687 & w33808;
assign w46038 = ~w33730 & w49354;
assign w46039 = (w33730 & w49355) | (w33730 & w49356) | (w49355 & w49356);
assign w46040 = (w33730 & w49357) | (w33730 & w49358) | (w49357 & w49358);
assign w46041 = ~w33730 & w49359;
assign w46042 = ~w32994 & w49360;
assign w46043 = w33900 & ~w33697;
assign w46044 = w32996 & ~w33927;
assign w46045 = w32996 & w33945;
assign w46046 = w32996 & w20906;
assign w46047 = w32996 & ~w20906;
assign w46048 = ~w33978 & w25851;
assign w46049 = w32974 & w50239;
assign w46050 = ~w34750 & w34752;
assign w46051 = ~w33718 & ~w34762;
assign w46052 = ~w34750 & w33723;
assign w46053 = w34750 & ~w34811;
assign w46054 = w34812 & ~w2006;
assign w46055 = w34132 & ~w33992;
assign w46056 = ~w33963 & w46982;
assign w46057 = ~w35428 & w46983;
assign w46058 = ~w35442 & ~w35436;
assign w46059 = ~w35442 & w34899;
assign w46060 = w7924 & ~w35441;
assign w46061 = (w7924 & w34899) | (w7924 & w46984) | (w34899 & w46984);
assign w46062 = w35527 & w35452;
assign w46063 = w35568 & ~w35629;
assign w46064 = ~w35568 & w35649;
assign w46065 = ~w35652 & ~w35661;
assign w46066 = ~w35662 & ~w35664;
assign w46067 = w35634 & ~w35670;
assign w46068 = ~w35680 & w35683;
assign w46069 = w34780 & ~w35693;
assign w46070 = w34780 & w42935;
assign w46071 = ~w35696 & w42937;
assign w46072 = ~w35705 & ~w35693;
assign w46073 = ~w35705 & w42935;
assign w46074 = ~w33855 & ~w35710;
assign w46075 = w35711 & ~w2006;
assign w46076 = ~w34740 & w34850;
assign w46077 = ~w35731 & ~w35732;
assign w46078 = w34715 & ~w2558;
assign w46079 = ~w35701 & w1738;
assign w46080 = w35747 & w35704;
assign w46081 = (~w35311 & ~w48036) | (~w35311 & w49941) | (~w48036 & w49941);
assign w46082 = w35605 & w35754;
assign w46083 = w33855 & ~w34834;
assign w46084 = ~w33855 & w1120;
assign w46085 = ~w34899 & w49362;
assign w46086 = (~w35776 & w34899) | (~w35776 & w49363) | (w34899 & w49363);
assign w46087 = ~w35784 & ~w35786;
assign w46088 = ~w42944 & w35786;
assign w46089 = ~w35788 & ~w35787;
assign w46090 = ~w35805 & ~w35804;
assign w46091 = w35671 & w35797;
assign w46092 = w35671 & w35775;
assign w46093 = ~w42945 & w33820;
assign w46094 = ~w42946 & w35842;
assign w46095 = w42946 & ~w35842;
assign w46096 = w35849 & ~w35848;
assign w46097 = ~w33855 & ~w34598;
assign w46098 = (w351 & w34899) | (w351 & w49364) | (w34899 & w49364);
assign w46099 = (w34881 & w49365) | (w34881 & w49366) | (w49365 & w49366);
assign w46100 = ~w34899 & w49367;
assign w46101 = (w34881 & w49942) | (w34881 & w49943) | (w49942 & w49943);
assign w46102 = ~w35966 & w35971;
assign w46103 = w35605 & w35984;
assign w46104 = w35099 & w36087;
assign w46105 = w35980 & ~w36093;
assign w46106 = w36092 & ~w28077;
assign w46107 = w36156 & w24874;
assign w46108 = ~w36173 & ~w36150;
assign w46109 = ~w35980 & w36404;
assign w46110 = ~w36397 & w35451;
assign w46111 = w36408 & w6769;
assign w46112 = ~w35980 & w7924;
assign w46113 = w36417 & ~w36411;
assign w46114 = ~w35980 & w35474;
assign w46115 = ~w35980 & ~w35462;
assign w46116 = w43022 & ~w35519;
assign w46117 = ~w36435 & w7924;
assign w46118 = ~w36408 & ~w6769;
assign w46119 = ~w35980 & ~w6769;
assign w46120 = w36441 & w36444;
assign w46121 = ~w36441 & w36446;
assign w46122 = ~w36461 & ~w36460;
assign w46123 = ~w35980 & ~w35515;
assign w46124 = w36491 & ~w9781;
assign w46125 = w36496 & ~w36549;
assign w46126 = w43045 & ~w36464;
assign w46127 = (~w36464 & w43045) | (~w36464 & w36547) | (w43045 & w36547);
assign w46128 = w35671 & w36617;
assign w46129 = w36027 & w36668;
assign w46130 = ~w36672 & w2006;
assign w46131 = ~w35980 & ~w2006;
assign w46132 = w36683 & w36686;
assign w46133 = ~w36683 & w36688;
assign w46134 = w36672 & ~w2006;
assign w46135 = w35671 & w43069;
assign w46136 = w43070 & w36741;
assign w46137 = (w36741 & w43070) | (w36741 & ~w35671) | (w43070 & ~w35671);
assign w46138 = w43071 & ~w35932;
assign w46139 = (~w35932 & w43071) | (~w35932 & ~w35671) | (w43071 & ~w35671);
assign w46140 = w43075 & ~w36764;
assign w46141 = (~w36764 & w43075) | (~w36764 & ~w35671) | (w43075 & ~w35671);
assign w46142 = w35980 & ~w36767;
assign w46143 = w35980 & w36767;
assign w46144 = w36786 & w36791;
assign w46145 = ~w36786 & w36793;
assign w46146 = w36786 & w36808;
assign w46147 = ~w36786 & w36810;
assign w46148 = ~w35802 & w36822;
assign w46149 = ~w36823 & w3646;
assign w46150 = w43079 & w35392;
assign w46151 = (w35392 & w43079) | (w35392 & ~w36823) | (w43079 & ~w36823);
assign w46152 = ~w36825 & ~w36828;
assign w46153 = w36827 & w35392;
assign w46154 = ~w36827 & ~w35392;
assign w46155 = w36857 & ~w36858;
assign w46156 = w36441 & w36443;
assign w46157 = w36861 & ~w6264;
assign w46158 = ~w35980 & ~w35537;
assign w46159 = ~w35980 & ~w35591;
assign w46160 = w36888 & w4838;
assign w46161 = w35671 & w36975;
assign w46162 = w43103 & ~w35859;
assign w46163 = (~w35859 & w43103) | (~w35859 & ~w35671) | (w43103 & ~w35671);
assign w46164 = w36976 & ~w80;
assign w46165 = ~w35858 & ~w80;
assign w46166 = ~w35980 & ~w80;
assign w46167 = ~w36976 & w80;
assign w46168 = w35671 & w37000;
assign w46169 = w35671 & w43108;
assign w46170 = ~w35980 & ~w35840;
assign w46171 = w35980 & w37023;
assign w46172 = ~w35980 & w35840;
assign w46173 = ~w36872 & ~w5745;
assign w46174 = ~w36888 & ~w4838;
assign w46175 = w36571 & w37110;
assign w46176 = w37114 & w37109;
assign w46177 = w37114 & ~w43114;
assign w46178 = ~w37106 & w37116;
assign w46179 = w36968 & w37140;
assign w46180 = ~w37142 & ~w37141;
assign w46181 = ~w37142 & ~w43115;
assign w46182 = ~w37106 & w37155;
assign w46183 = w36968 & w37167;
assign w46184 = w37106 & ~w37180;
assign w46185 = ~w37106 & ~w37183;
assign w46186 = ~w37170 & ~w37168;
assign w46187 = ~w37170 & ~w43117;
assign w46188 = w37106 & ~w37202;
assign w46189 = w37106 & ~w37212;
assign w46190 = w37173 & w1120;
assign w46191 = w37218 & ~w1120;
assign w46192 = w36968 & ~w36697;
assign w46193 = w37226 & ~w36682;
assign w46194 = w37106 & ~w1738;
assign w46195 = w37226 & w37235;
assign w46196 = w37106 & w1541;
assign w46197 = w37240 & w37242;
assign w46198 = ~w37240 & w37244;
assign w46199 = w37106 & w36681;
assign w46200 = w37250 & ~w37225;
assign w46201 = w37250 & ~w43121;
assign w46202 = w36968 & w37255;
assign w46203 = w37106 & ~w36126;
assign w46204 = ~w37106 & w37351;
assign w46205 = w37106 & w37373;
assign w46206 = ~w37106 & w37375;
assign w46207 = w37106 & w37391;
assign w46208 = ~w37106 & w37390;
assign w46209 = w37106 & w37397;
assign w46210 = ~w37106 & w37400;
assign w46211 = ~w37106 & w37409;
assign w46212 = w37106 & w37424;
assign w46213 = ~w37106 & w37426;
assign w46214 = w37106 & w37456;
assign w46215 = ~w37106 & w37458;
assign w46216 = w36118 & w36221;
assign w46217 = w37106 & w24874;
assign w46218 = ~w37106 & w37526;
assign w46219 = w37540 & w36203;
assign w46220 = w37106 & w37550;
assign w46221 = ~w37106 & w37552;
assign w46222 = w37106 & w37561;
assign w46223 = w37106 & w37567;
assign w46224 = ~w37106 & w37569;
assign w46225 = ~w37540 & ~w36202;
assign w46226 = ~w37554 & w37571;
assign w46227 = w37106 & w36384;
assign w46228 = ~w37106 & ~w37644;
assign w46229 = w37106 & w36237;
assign w46230 = w37656 & w19040;
assign w46231 = w37106 & w36148;
assign w46232 = ~w37106 & ~w37670;
assign w46233 = ~w37674 & ~w37675;
assign w46234 = w36564 & ~w36385;
assign w46235 = w36386 & w37698;
assign w46236 = w37106 & ~w36524;
assign w46237 = w37706 & w11138;
assign w46238 = ~w37715 & ~w37714;
assign w46239 = w37106 & ~w36532;
assign w46240 = w37106 & w37731;
assign w46241 = ~w37741 & ~w37742;
assign w46242 = ~w36375 & ~w12666;
assign w46243 = w37106 & ~w36379;
assign w46244 = ~w37751 & w13384;
assign w46245 = w36564 & w37757;
assign w46246 = ~w37106 & w37763;
assign w46247 = w37106 & w36352;
assign w46248 = ~w37724 & w11870;
assign w46249 = ~w37706 & ~w11138;
assign w46250 = w37106 & w15681;
assign w46251 = w37791 & w37796;
assign w46252 = ~w37791 & w37798;
assign w46253 = w37791 & w37811;
assign w46254 = ~w37791 & w37813;
assign w46255 = ~w37781 & w37818;
assign w46256 = ~w37842 & w37844;
assign w46257 = w37106 & w37875;
assign w46258 = w36863 & w37882;
assign w46259 = w37106 & w36436;
assign w46260 = w37896 & w7315;
assign w46261 = ~w37917 & w37919;
assign w46262 = ~w37921 & ~w37922;
assign w46263 = ~w37915 & w36496;
assign w46264 = w37697 & ~w37946;
assign w46265 = ~w37697 & ~w37949;
assign w46266 = ~w37945 & w9781;
assign w46267 = ~w37915 & w37968;
assign w46268 = ~w37967 & ~w37970;
assign w46269 = w37106 & ~w36494;
assign w46270 = w37973 & w9195;
assign w46271 = ~w37106 & w37959;
assign w46272 = ~w10419 & ~w37955;
assign w46273 = w37935 & w8666;
assign w46274 = ~w38001 & ~w37099;
assign w46275 = ~w38020 & w38022;
assign w46276 = w37994 & ~w38000;
assign w46277 = ~w38037 & w3242;
assign w46278 = w38060 & w38022;
assign w46279 = w43139 & w38094;
assign w46280 = (w38094 & w43139) | (w38094 & ~w36571) | (w43139 & ~w36571);
assign w46281 = w37106 & ~w36891;
assign w46282 = w43140 & w38100;
assign w46283 = (w38100 & w43140) | (w38100 & ~w36571) | (w43140 & ~w36571);
assign w46284 = ~w38103 & w4430;
assign w46285 = ~w38105 & ~w4056;
assign w46286 = ~w37883 & ~w36876;
assign w46287 = w38124 & w38174;
assign w46288 = w38338 & ~w38424;
assign w46289 = w37446 & ~w38433;
assign w46290 = w37446 & w43167;
assign w46291 = ~w38454 & w38452;
assign w46292 = ~w38454 & w43168;
assign w46293 = ~w38463 & ~w38461;
assign w46294 = ~w38472 & w38469;
assign w46295 = ~w38472 & w43171;
assign w46296 = w38338 & ~w28077;
assign w46297 = w37377 & w43172;
assign w46298 = w25851 & ~w38501;
assign w46299 = w25851 & ~w43175;
assign w46300 = w38511 & ~w38509;
assign w46301 = w38511 & ~w43176;
assign w46302 = w38513 & w38509;
assign w46303 = w38513 & w43176;
assign w46304 = w37492 & w38452;
assign w46305 = w37492 & w43168;
assign w46306 = ~w37824 & ~w38525;
assign w46307 = ~w37824 & w43178;
assign w46308 = ~w38541 & ~w37829;
assign w46309 = ~w38541 & w43182;
assign w46310 = w38548 & w38526;
assign w46311 = w38548 & w43181;
assign w46312 = w38551 & w38526;
assign w46313 = w38551 & w43181;
assign w46314 = ~w38338 & w38566;
assign w46315 = ~w37695 & w38572;
assign w46316 = w43188 | ~w37823;
assign w46317 = (~w37823 & w43188) | (~w37823 & w38573) | (w43188 & w38573);
assign w46318 = w43190 | w38585;
assign w46319 = (w38585 & w43190) | (w38585 & w38573) | (w43190 & w38573);
assign w46320 = ~w38338 & w38588;
assign w46321 = ~w38338 & w38591;
assign w46322 = w38589 & ~w12666;
assign w46323 = w38338 & w37822;
assign w46324 = ~w38609 & w13384;
assign w46325 = ~w43195 & ~w37621;
assign w46326 = ~w37659 & ~w37639;
assign w46327 = ~w37659 & w43199;
assign w46328 = w38700 & ~w38701;
assign w46329 = w22767 & w38723;
assign w46330 = ~w38338 & w38764;
assign w46331 = w38338 & w38767;
assign w46332 = w38773 & ~w38775;
assign w46333 = w37789 & w38555;
assign w46334 = w37789 & ~w43185;
assign w46335 = w38829 & ~w37639;
assign w46336 = w38829 & w43199;
assign w46337 = w38838 & ~w38824;
assign w46338 = w38338 & ~w38856;
assign w46339 = ~w38338 & ~w38868;
assign w46340 = ~w37835 & w10419;
assign w46341 = ~w38874 & ~w38875;
assign w46342 = ~w38874 & w43201;
assign w46343 = ~w38589 & w12666;
assign w46344 = w38338 & ~w11870;
assign w46345 = w38895 & w38900;
assign w46346 = ~w38895 & w38902;
assign w46347 = ~w38895 & ~w38899;
assign w46348 = w43204 | w38162;
assign w46349 = (w38162 & w43204) | (w38162 & w37835) | (w43204 & w37835);
assign w46350 = w38338 & ~w38944;
assign w46351 = w43206 | ~w38159;
assign w46352 = (~w38159 & w43206) | (~w38159 & w37835) | (w43206 & w37835);
assign w46353 = ~w37928 & w43207;
assign w46354 = w37835 & w38959;
assign w46355 = ~w37899 & w38962;
assign w46356 = ~w37899 & w43208;
assign w46357 = w37835 & w39028;
assign w46358 = ~w37835 & w37993;
assign w46359 = ~w38338 & ~w3242;
assign w46360 = ~w38338 & ~w38115;
assign w46361 = w38338 & w38116;
assign w46362 = ~w38338 & w39109;
assign w46363 = ~w43219 & w2006;
assign w46364 = ~w39170 & ~w39176;
assign w46365 = w1738 & ~w43220;
assign w46366 = ~w38338 & ~w2558;
assign w46367 = ~w38338 & w2558;
assign w46368 = ~w38338 & w39302;
assign w46369 = ~w37316 & ~w38254;
assign w46370 = w38195 & ~w37300;
assign w46371 = ~w37247 & ~w37205;
assign w46372 = ~w37288 & w39424;
assign w46373 = ~w38338 & ~w39426;
assign w46374 = ~w38190 & ~w37192;
assign w46375 = ~w38338 & w754;
assign w46376 = ~w39450 & w945;
assign w46377 = ~w39167 & w43216;
assign w46378 = ~w39167 & ~w2285;
assign w46379 = ~w39167 & w43214;
assign w46380 = w39167 & w2285;
assign w46381 = w39167 & ~w43214;
assign w46382 = w38338 & ~w1320;
assign w46383 = w39515 & w39514;
assign w46384 = ~w39515 & ~w39514;
assign w46385 = ~w39525 & w400;
assign w46386 = ~w39523 & w39527;
assign w46387 = ~w39523 & w39546;
assign w46388 = ~w43218 & ~w39558;
assign w46389 = w43218 & ~w39560;
assign w46390 = ~w43239 & ~w39560;
assign w46391 = w43218 & ~w39176;
assign w46392 = w39567 & ~w1738;
assign w46393 = ~w39450 & ~w39587;
assign w46394 = w492 & w419;
assign w46395 = ~w492 & ~w419;
assign w46396 = w1134 & w252;
assign w46397 = w1160 & w1162;
assign w46398 = ~w1160 & w1164;
assign w46399 = ~w1160 & ~w1161;
assign w46400 = w1160 & w1161;
assign w46401 = ~w1224 & ~w1202;
assign w46402 = w1224 & ~w3;
assign w46403 = w1499 & ~w3;
assign w46404 = w1499 & w39824;
assign w46405 = ~w1120 & w1554;
assign w46406 = ~w1120 & w39831;
assign w46407 = w1559 & w1555;
assign w46408 = w1559 & ~w39832;
assign w46409 = ~w1370 & ~w1590;
assign w46410 = ~w1370 & ~w39840;
assign w46411 = w1603 & ~w1602;
assign w46412 = w1603 & ~w39844;
assign w46413 = w1605 & w1602;
assign w46414 = w1605 & w39844;
assign w46415 = w1608 & ~w1590;
assign w46416 = w1608 & ~w39840;
assign w46417 = w1610 & w1590;
assign w46418 = w1610 & w39840;
assign w46419 = w1641 & ~w1602;
assign w46420 = w1641 & ~w39844;
assign w46421 = w1643 & w1602;
assign w46422 = w1643 & w39844;
assign w46423 = ~w1493 & w42;
assign w46424 = (~w3 & ~w1699) | (~w3 & w51402) | (~w1699 & w51402);
assign w46425 = (w3 & ~w1699) | (w3 & w51403) | (~w1699 & w51403);
assign w46426 = w1699 & w51404;
assign w46427 = (w1764 & ~w1699) | (w1764 & w51405) | (~w1699 & w51405);
assign w46428 = w1699 & w51406;
assign w46429 = (w1778 & ~w1699) | (w1778 & w51407) | (~w1699 & w51407);
assign w46430 = w1699 & w51408;
assign w46431 = (w1784 & ~w1699) | (w1784 & w51409) | (~w1699 & w51409);
assign w46432 = w1699 & w51410;
assign w46433 = w1699 & w51411;
assign w46434 = (w1775 & ~w1699) | (w1775 & w51412) | (~w1699 & w51412);
assign w46435 = w1725 & ~w1806;
assign w46436 = w1699 & w51413;
assign w46437 = (w1814 & ~w1699) | (w1814 & w51414) | (~w1699 & w51414);
assign w46438 = ~w1691 & w43288;
assign w46439 = w1699 & w51415;
assign w46440 = (w1934 & ~w1699) | (w1934 & w51416) | (~w1699 & w51416);
assign w46441 = w1699 & w51417;
assign w46442 = (w1943 & ~w1699) | (w1943 & w51418) | (~w1699 & w51418);
assign w46443 = ~w2897 & ~w400;
assign w46444 = ~w2680 & w3226;
assign w46445 = w2922 & w3248;
assign w46446 = w2922 & w3269;
assign w46447 = w2922 & ~w3328;
assign w46448 = w3388 & w3385;
assign w46449 = ~w3388 & ~w3385;
assign w46450 = w2922 & ~w3424;
assign w46451 = w3425 & ~w493;
assign w46452 = w2922 & w3206;
assign w46453 = w2922 & w2981;
assign w46454 = w40076 & ~w754;
assign w46455 = w3443 & w612;
assign w46456 = ~w40076 & w754;
assign w46457 = w2922 & w400;
assign w46458 = ~w3508 & ~w3513;
assign w46459 = w2954 & w3554;
assign w46460 = ~w2954 & w3560;
assign w46461 = w3606 & w48473;
assign w46462 = w3607 & w3765;
assign w46463 = w3606 & w48474;
assign w46464 = w3606 & w48475;
assign w46465 = w3606 & w48476;
assign w46466 = w3606 & w48477;
assign w46467 = w3607 & w3579;
assign w46468 = w3607 & w3519;
assign w46469 = w4054 & ~w57;
assign w46470 = ~w4051 & w48478;
assign w46471 = (~w4080 & w50418) | (~w4080 & w50419) | (w50418 & w50419);
assign w46472 = ~w4051 & w48479;
assign w46473 = ~w4187 & ~w4186;
assign w46474 = w4054 & w4215;
assign w46475 = w4054 & w4233;
assign w46476 = ~w4054 & w4232;
assign w46477 = ~w4054 & ~w4243;
assign w46478 = w4054 & ~w4246;
assign w46479 = (w4269 & w4051) | (w4269 & w51419) | (w4051 & w51419);
assign w46480 = ~w4051 & w51420;
assign w46481 = (w4279 & w4051) | (w4279 & w51421) | (w4051 & w51421);
assign w46482 = (w4287 & w4051) | (w4287 & w51422) | (w4051 & w51422);
assign w46483 = ~w3878 & ~w1541;
assign w46484 = ~w4051 & w48480;
assign w46485 = w3878 & w1541;
assign w46486 = ~w4051 & w51423;
assign w46487 = ~w4051 & w51424;
assign w46488 = ~w4138 & ~w4407;
assign w46489 = w43361 | ~w4204;
assign w46490 = (~w4204 & w43361) | (~w4204 & ~w4401) | (w43361 & ~w4401);
assign w46491 = w4409 & ~w4715;
assign w46492 = ~w40251 & w5134;
assign w46493 = w5625 & ~w5640;
assign w46494 = ~w5763 & ~w351;
assign w46495 = ~w351 & ~w5640;
assign w46496 = ~w351 & w40294;
assign w46497 = ~w40299 & w5798;
assign w46498 = ~w40301 & w5802;
assign w46499 = w5763 & w351;
assign w46500 = ~w40301 & w5814;
assign w46501 = ~w5771 & ~w5791;
assign w46502 = w5743 & w5861;
assign w46503 = w5743 & w5869;
assign w46504 = w5743 & w5920;
assign w46505 = ~w40328 & ~w1738;
assign w46506 = w5743 & w5956;
assign w46507 = w5385 & w5875;
assign w46508 = w5385 & w40316;
assign w46509 = w5743 & w6080;
assign w46510 = ~w5743 & w6079;
assign w46511 = w5743 & w6096;
assign w46512 = w40328 & w1738;
assign w46513 = ~w5703 & w6125;
assign w46514 = w5743 & ~w5563;
assign w46515 = ~w5546 & ~w5502;
assign w46516 = w5546 & ~w5502;
assign w46517 = w5743 & w6214;
assign w46518 = w5743 & w6222;
assign w46519 = w40355 & w1120;
assign w46520 = ~w40378 & w945;
assign w46521 = w6113 & w5855;
assign w46522 = ~w6092 & w6269;
assign w46523 = ~w6092 & w6503;
assign w46524 = ~w6254 & ~w80;
assign w46525 = (w6735 & ~w6642) | (w6735 & w48481) | (~w6642 & w48481);
assign w46526 = ~w252 & w7835;
assign w46527 = w252 & w7837;
assign w46528 = w7935 & w8586;
assign w46529 = ~w7935 & w8588;
assign w46530 = ~w8189 & ~w7945;
assign w46531 = w8539 & w8682;
assign w46532 = ~w8687 & ~w8458;
assign w46533 = w8189 & w8977;
assign w46534 = ~w8189 & w8979;
assign w46535 = w8157 & ~w9102;
assign w46536 = ~w9064 & w8158;
assign w46537 = w9064 & ~w8158;
assign w46538 = w12255 & w12252;
assign w46539 = (w12255 & w12251) | (w12255 & w46538) | (w12251 & w46538);
assign w46540 = w12257 & ~w12252;
assign w46541 = ~w12251 & w46540;
assign w46542 = w12269 & w12266;
assign w46543 = (w12269 & w12265) | (w12269 & w46542) | (w12265 & w46542);
assign w46544 = w12271 & ~w12266;
assign w46545 = ~w12265 & w46544;
assign w46546 = ~w12179 & ~w12176;
assign w46547 = ~w12179 & w41030;
assign w46548 = w12560 & ~w12491;
assign w46549 = w12560 & w41083;
assign w46550 = ~w12254 & ~w12252;
assign w46551 = ~w12254 & w41044;
assign w46552 = w12254 & w12252;
assign w46553 = w12254 & ~w41044;
assign w46554 = w12043 & ~w12835;
assign w46555 = ~w12936 & ~w4430;
assign w46556 = ~w14652 & w351;
assign w46557 = w14652 & ~w351;
assign w46558 = ~w14069 & w14074;
assign w46559 = w14707 & ~w14767;
assign w46560 = ~w14707 & w14767;
assign w46561 = w15091 & ~w14297;
assign w46562 = w15091 & w41287;
assign w46563 = w4056 & ~w14297;
assign w46564 = ~w14213 & w46563;
assign w46565 = ~w4056 & w14297;
assign w46566 = (~w4056 & w14213) | (~w4056 & w46565) | (w14213 & w46565);
assign w46567 = w14761 & w48482;
assign w46568 = (w15268 & ~w14761) | (w15268 & w48483) | (~w14761 & w48483);
assign w46569 = w14761 & w48484;
assign w46570 = (w15358 & ~w14761) | (w15358 & w48485) | (~w14761 & w48485);
assign w46571 = w43502 | w16085;
assign w46572 = (w16085 & w43502) | (w16085 & w15551) | (w43502 & w15551);
assign w46573 = ~w15551 & w43503;
assign w46574 = w15679 & w14806;
assign w46575 = ~w16245 & w16538;
assign w46576 = ~w9195 & ~w20639;
assign w46577 = ~w20120 & ~w20226;
assign w46578 = ~w21241 & w22007;
assign w46579 = ~w21241 & w22050;
assign w46580 = w21241 & ~w21214;
assign w46581 = ~w41927 & ~w7315;
assign w46582 = w21241 & ~w21298;
assign w46583 = ~w41930 & ~w5745;
assign w46584 = w22558 & ~w6769;
assign w46585 = w21241 & ~w5330;
assign w46586 = ~w21241 & w22630;
assign w46587 = ~w21241 & w21772;
assign w46588 = w21241 & ~w4838;
assign w46589 = w41961 & w22734;
assign w46590 = ~w41961 & ~w22734;
assign w46591 = w23216 & ~w23219;
assign w46592 = ~w23216 & w23219;
assign w46593 = ~w12666 & ~w23265;
assign w46594 = ~w12666 & w42006;
assign w46595 = w23301 & w23304;
assign w46596 = ~w23301 & ~w23304;
assign w46597 = ~w23301 & w23316;
assign w46598 = w23301 & w23318;
assign w46599 = w22763 & w22137;
assign w46600 = ~w24913 & ~w24859;
assign w46601 = ~w24913 & w42085;
assign w46602 = w24912 & w10419;
assign w46603 = (~w12666 & w24865) | (~w12666 & w49368) | (w24865 & w49368);
assign w46604 = w24864 & w7315;
assign w46605 = w24864 & w24556;
assign w46606 = w25098 & w24158;
assign w46607 = ~w25098 & ~w24158;
assign w46608 = w20906 & ~w25204;
assign w46609 = ~w24870 & w25110;
assign w46610 = w24870 & ~w20000;
assign w46611 = ~w24232 & ~w25299;
assign w46612 = ~w42131 & w43586;
assign w46613 = ~w25394 & w48486;
assign w46614 = ~w5745 & w24561;
assign w46615 = ~w42166 & ~w25502;
assign w46616 = w6264 & ~w24859;
assign w46617 = w6264 & w42085;
assign w46618 = ~w5745 & w25516;
assign w46619 = w25529 & ~w2558;
assign w46620 = w3646 & w25559;
assign w46621 = w3646 & w24417;
assign w46622 = w3646 & w42188;
assign w46623 = ~w25357 & ~w2285;
assign w46624 = w42212 & w25727;
assign w46625 = w26950 & ~w26177;
assign w46626 = w26959 & ~w754;
assign w46627 = w754 & ~w26959;
assign w46628 = ~w26073 & w4430;
assign w46629 = w26076 & ~w27265;
assign w46630 = w26876 & ~w27265;
assign w46631 = ~w26073 & ~w27263;
assign w46632 = w27273 & ~w27276;
assign w46633 = ~w26073 & w27309;
assign w46634 = w26076 & w27314;
assign w46635 = w26076 & w27322;
assign w46636 = w26876 & w27374;
assign w46637 = w26076 & w27374;
assign w46638 = ~w27446 & ~w27447;
assign w46639 = w26078 & w26127;
assign w46640 = ~w26078 & ~w26127;
assign w46641 = ~w27339 & w27258;
assign w46642 = (w28412 & w28037) | (w28412 & w49944) | (w28037 & w49944);
assign w46643 = ~w28453 & ~w28456;
assign w46644 = ~w27253 & w28702;
assign w46645 = ~w28813 & w26973;
assign w46646 = w42420 & ~w2558;
assign w46647 = ~w27177 & w2896;
assign w46648 = ~w28929 & ~w30044;
assign w46649 = w28882 & w3;
assign w46650 = ~w28882 & w30058;
assign w46651 = ~w30034 & w43690;
assign w46652 = ~w30145 & ~w29977;
assign w46653 = w30287 & w30289;
assign w46654 = ~w30287 & w30291;
assign w46655 = w400 & w30294;
assign w46656 = ~w30145 & ~w29926;
assign w46657 = w30287 & w30317;
assign w46658 = ~w30287 & w30319;
assign w46659 = ~w30145 & ~w30525;
assign w46660 = w30531 & w28077;
assign w46661 = ~w30572 & w30576;
assign w46662 = w30560 & w30578;
assign w46663 = w30606 & w29484;
assign w46664 = ~w30606 & ~w29484;
assign w46665 = w30807 & ~w11870;
assign w46666 = ~w30807 & w11870;
assign w46667 = ~w30836 & ~w14766;
assign w46668 = ~w30836 & ~w42513;
assign w46669 = w30897 & ~w30836;
assign w46670 = ~w30897 & w30836;
assign w46671 = ~w30884 & w15681;
assign w46672 = ~w30182 & ~w4056;
assign w46673 = w29674 & w5745;
assign w46674 = w29736 & ~w5330;
assign w46675 = ~w29674 & ~w5745;
assign w46676 = w30182 & w4056;
assign w46677 = w2006 & ~w29823;
assign w46678 = ~w30145 & ~w31250;
assign w46679 = w2558 & w31271;
assign w46680 = ~w2558 & w31274;
assign w46681 = ~w2558 & w31280;
assign w46682 = w2558 & w31285;
assign w46683 = w30216 & w31298;
assign w46684 = ~w2896 & w31298;
assign w46685 = w2896 & w31304;
assign w46686 = w2896 & w31310;
assign w46687 = ~w2896 & w31313;
assign w46688 = w29821 & w29794;
assign w46689 = ~w31662 & w30877;
assign w46690 = ~w31772 & ~w31773;
assign w46691 = ~w31793 & ~w31794;
assign w46692 = ~w31811 & w50246;
assign w46693 = ~w31876 & ~w31877;
assign w46694 = ~w32392 & w57;
assign w46695 = w400 & w32444;
assign w46696 = w33001 & w31971;
assign w46697 = w33342 & ~w31668;
assign w46698 = ~w33435 & ~w6264;
assign w46699 = ~w32790 & ~w33734;
assign w46700 = ~w32790 & w33874;
assign w46701 = w32710 & ~w33937;
assign w46702 = ~w32710 & ~w33927;
assign w46703 = ~w32710 & w33945;
assign w46704 = w32710 & ~w33080;
assign w46705 = w32710 & w33098;
assign w46706 = ~w32790 & w33985;
assign w46707 = w32790 & w33987;
assign w46708 = w32710 & w34000;
assign w46709 = ~w32710 & w20906;
assign w46710 = ~w32710 & ~w20906;
assign w46711 = ~w32790 & w34126;
assign w46712 = w32790 & w34128;
assign w46713 = ~w32790 & w34140;
assign w46714 = ~w32790 & ~w33289;
assign w46715 = w33361 & ~w34209;
assign w46716 = w34313 & w34584;
assign w46717 = ~w33668 & ~w33450;
assign w46718 = ~w34320 & ~w33450;
assign w46719 = ~w34320 & w42764;
assign w46720 = ~w32790 & w34326;
assign w46721 = w34332 & w34331;
assign w46722 = ~w34332 & ~w34331;
assign w46723 = ~w33485 & ~w33659;
assign w46724 = ~w32790 & w34361;
assign w46725 = ~w33438 & w42764;
assign w46726 = ~w32790 & ~w33437;
assign w46727 = ~w32790 & w7315;
assign w46728 = ~w32790 & w4838;
assign w46729 = ~w33622 & ~w34423;
assign w46730 = ~w32790 & w33609;
assign w46731 = w33699 & w33702;
assign w46732 = w32710 & w34444;
assign w46733 = ~w33552 & ~w34469;
assign w46734 = w33552 & w34466;
assign w46735 = ~w32790 & w34533;
assign w46736 = ~w33634 & w9781;
assign w46737 = w33634 & ~w9781;
assign w46738 = ~w32790 & ~w34550;
assign w46739 = ~w32790 & w34560;
assign w46740 = ~w42686 & w34593;
assign w46741 = w32790 & w32807;
assign w46742 = w32790 & ~w34610;
assign w46743 = w32790 & w34610;
assign w46744 = w32710 & w2896;
assign w46745 = ~w42825 & w34671;
assign w46746 = ~w32790 & ~w2558;
assign w46747 = ~w32790 & w34711;
assign w46748 = ~w42824 & w34717;
assign w46749 = w42824 & w34720;
assign w46750 = ~w3646 & ~w34729;
assign w46751 = ~w3646 & ~w42844;
assign w46752 = ~w32790 & w34798;
assign w46753 = ~w32790 & w32962;
assign w46754 = ~w34812 & w2006;
assign w46755 = w8666 & w35423;
assign w46756 = ~w34168 & w49369;
assign w46757 = ~w8666 & ~w35423;
assign w46758 = (~w8666 & w34168) | (~w8666 & w49370) | (w34168 & w49370);
assign w46759 = w35639 & ~w35641;
assign w46760 = ~w35986 & ~w36020;
assign w46761 = ~w36838 & ~w37099;
assign w46762 = w36968 & ~w2285;
assign w46763 = w36968 & w36697;
assign w46764 = w36968 & ~w37327;
assign w46765 = w36968 & ~w37498;
assign w46766 = w36968 & ~w37507;
assign w46767 = w36968 & ~w37584;
assign w46768 = w36968 & w37600;
assign w46769 = w36968 & w37912;
assign w46770 = w36968 & w36935;
assign w46771 = w36968 & ~w36855;
assign w46772 = w36968 & ~w36958;
assign w46773 = ~w38140 & w39363;
assign w46774 = (w1877 & ~w1699) | (w1877 & w51425) | (~w1699 & w51425);
assign w46775 = w1699 & w51426;
assign w46776 = (w1892 & ~w1699) | (w1892 & w51427) | (~w1699 & w51427);
assign w46777 = w1699 & w51428;
assign w46778 = w4378 & ~w1120;
assign w46779 = ~w14882 & ~w14966;
assign w46780 = ~w26316 & w26720;
assign w46781 = ~w26316 & w26718;
assign w46782 = ~w28143 & w27270;
assign w46783 = ~w28166 & ~w28193;
assign w46784 = ~w28313 & w48487;
assign w46785 = w43637 & w28528;
assign w46786 = ~w43637 & w28530;
assign w46787 = ~w43637 & ~w28527;
assign w46788 = w43637 & w28527;
assign w46789 = ~w43650 & w8666;
assign w46790 = w43653 & ~w28696;
assign w46791 = w43668 & w2006;
assign w46792 = w43676 & w29123;
assign w46793 = ~w43676 & w29125;
assign w46794 = ~w43676 & ~w29122;
assign w46795 = w43676 & w29122;
assign w46796 = ~w30230 & ~w2006;
assign w46797 = w30516 & ~w31966;
assign w46798 = ~w4838 & ~w30517;
assign w46799 = w5745 & ~w32236;
assign w46800 = ~w32710 & ~w32717;
assign w46801 = ~w32710 & w32842;
assign w46802 = w32710 & w34745;
assign w46803 = w32710 & ~w1541;
assign w46804 = w43774 & w34793;
assign w46805 = ~w43788 & w8666;
assign w46806 = w1138 & ~w57;
assign w46807 = w1323 & w80;
assign w46808 = ~w1138 & w57;
assign w46809 = ~w1224 & w1486;
assign w46810 = ~w1224 & ~w80;
assign w46811 = w1636 & ~w1671;
assign w46812 = ~w2134 & ~w2344;
assign w46813 = ~w2134 & ~w2185;
assign w46814 = w2134 & w1120;
assign w46815 = w2284 & w2420;
assign w46816 = ~w2284 & w2422;
assign w46817 = w2134 & w612;
assign w46818 = ~w2284 & w2439;
assign w46819 = w2284 & w2441;
assign w46820 = ~w2284 & w2452;
assign w46821 = w2284 & w2454;
assign w46822 = w2284 & ~w2451;
assign w46823 = ~w2284 & w2451;
assign w46824 = ~w2134 & w2099;
assign w46825 = ~w2134 & ~w2519;
assign w46826 = ~w2134 & w2519;
assign w46827 = w2134 & w80;
assign w46828 = w2792 & w43309;
assign w46829 = ~w2805 & ~w43312;
assign w46830 = ~a[95] & ~w44019;
assign w46831 = ~a[95] & ~w44020;
assign w46832 = ~w2611 & w2589;
assign w46833 = w2986 & ~w945;
assign w46834 = ~w3029 & w3032;
assign w46835 = w3029 & w3034;
assign w46836 = ~w3057 & ~w3058;
assign w46837 = ~w2986 & w945;
assign w46838 = w3099 & ~w3100;
assign w46839 = ~w3132 & ~w2589;
assign w46840 = ~w3132 & ~w44031;
assign w46841 = w3766 & w2896;
assign w46842 = ~w3765 & ~w2896;
assign w46843 = ~w44088 & ~w2558;
assign w46844 = w44088 & w2558;
assign w46845 = ~w400 & w3907;
assign w46846 = w400 & w3910;
assign w46847 = w42 & ~w3952;
assign w46848 = w42 & w40135;
assign w46849 = ~w80 & w3983;
assign w46850 = w80 & w3986;
assign w46851 = ~w3597 & w57;
assign w46852 = ~w80 & w4030;
assign w46853 = w80 & w4033;
assign w46854 = (w3646 & w4418) | (w3646 & w48488) | (w4418 & w48488);
assign w46855 = w4418 & w48489;
assign w46856 = (~w1738 & ~w4418) | (~w1738 & w48490) | (~w4418 & w48490);
assign w46857 = ~w4660 & ~w754;
assign w46858 = w4660 & w754;
assign w46859 = w40210 & ~w4387;
assign w46860 = ~w4387 & w1120;
assign w46861 = (w4372 & w46860) | (w4372 & w48491) | (w46860 & w48491);
assign w46862 = w4418 & w48492;
assign w46863 = (w4810 & ~w4418) | (w4810 & w48493) | (~w4418 & w48493);
assign w46864 = (w4824 & ~w4418) | (w4824 & w48494) | (~w4418 & w48494);
assign w46865 = w4418 & w48495;
assign w46866 = a[79] & w5346;
assign w46867 = ~a[79] & w5351;
assign w46868 = a[79] & w5362;
assign w46869 = ~a[79] & a[78];
assign w46870 = ~w1120 & ~w5161;
assign w46871 = ~w1120 & w44187;
assign w46872 = ~w1320 & w5150;
assign w46873 = ~w1320 & w44194;
assign w46874 = w5559 & ~w754;
assign w46875 = ~w5854 & ~w6256;
assign w46876 = ~w5854 & w6297;
assign w46877 = ~w6536 & w6562;
assign w46878 = ~w6536 & w6556;
assign w46879 = w7425 & w612;
assign w46880 = ~w7425 & ~w612;
assign w46881 = w7923 & w252;
assign w46882 = ~w7909 & w8296;
assign w46883 = w8568 & w8612;
assign w46884 = w8568 & ~w8612;
assign w46885 = ~w8568 & w8612;
assign w46886 = w44409 & w8982;
assign w46887 = ~w44409 & ~w8982;
assign w46888 = ~w44416 & w9033;
assign w46889 = w9077 & w8983;
assign w46890 = ~w44416 & w9081;
assign w46891 = w44498 & ~w1541;
assign w46892 = w44502 & ~w1320;
assign w46893 = ~w44498 & w1541;
assign w46894 = w80 & w13896;
assign w46895 = ~w80 & ~w13896;
assign w46896 = w80 & ~w14792;
assign w46897 = ~w14500 & w493;
assign w46898 = w14500 & ~w493;
assign w46899 = ~w80 & w14600;
assign w46900 = ~w14203 & ~w4430;
assign w46901 = ~w14203 & w15184;
assign w46902 = w5745 & w15224;
assign w46903 = ~w5745 & w15227;
assign w46904 = ~w14125 & ~w14126;
assign w46905 = w15361 & w5745;
assign w46906 = w14203 & w4430;
assign w46907 = w14777 & ~w15718;
assign w46908 = w14777 & w15719;
assign w46909 = w14777 & w15707;
assign w46910 = w14777 & w15744;
assign w46911 = w14777 & ~w15514;
assign w46912 = ~w15271 & w15233;
assign w46913 = w14777 & ~w15195;
assign w46914 = w14777 & ~w3646;
assign w46915 = w14777 & w16016;
assign w46916 = ~w15618 & w16310;
assign w46917 = ~w15537 & w16310;
assign w46918 = w14777 & w400;
assign w46919 = w16948 & w17367;
assign w46920 = w17042 & ~w17357;
assign w46921 = (w17042 & w17365) | (w17042 & w49371) | (w17365 & w49371);
assign w46922 = w21241 & ~w21283;
assign w46923 = w45244 & w5330;
assign w46924 = w41942 & w22603;
assign w46925 = ~w41942 & ~w22603;
assign w46926 = w13384 & ~w23294;
assign w46927 = ~w24237 & ~w24161;
assign w46928 = w24568 & ~w24540;
assign w46929 = ~w45412 & ~w7924;
assign w46930 = ~w45414 & ~w9195;
assign w46931 = w45414 & w9195;
assign w46932 = w45412 & w7924;
assign w46933 = w25113 & w24142;
assign w46934 = w24556 & w4056;
assign w46935 = ~w26052 & ~w26053;
assign w46936 = ~w26729 & w1738;
assign w46937 = ~w26729 & ~w45586;
assign w46938 = w26729 & ~w1738;
assign w46939 = w26729 & w45586;
assign w46940 = ~w26377 & w3646;
assign w46941 = ~w27109 & ~w4056;
assign w46942 = w27109 & w4056;
assign w46943 = ~w27116 & w4056;
assign w46944 = ~w27298 & ~w25945;
assign w46945 = ~w27298 & w45513;
assign w46946 = w28107 & w24874;
assign w46947 = w28133 & w24874;
assign w46948 = ~w28133 & ~w24874;
assign w46949 = w27484 & ~w27636;
assign w46950 = ~w27250 & w28002;
assign w46951 = ~w28498 & w28677;
assign w46952 = w29657 & w29363;
assign w46953 = ~w351 & w30263;
assign w46954 = w351 & w30265;
assign w46955 = w351 & ~w30262;
assign w46956 = ~w351 & w30262;
assign w46957 = w31174 & w31179;
assign w46958 = ~w1738 & w31234;
assign w46959 = w1738 & w31236;
assign w46960 = ~w1738 & w31368;
assign w46961 = w1738 & w31370;
assign w46962 = w1738 & ~w31233;
assign w46963 = ~w1738 & w31233;
assign w46964 = w2285 & w31391;
assign w46965 = ~w32392 & ~w32614;
assign w46966 = ~w32392 & w32622;
assign w46967 = w80 & w32621;
assign w46968 = ~w80 & ~w32621;
assign w46969 = w32415 & w32323;
assign w46970 = ~w2896 & ~w33563;
assign w46971 = w2896 & w33563;
assign w46972 = ~w32097 & ~w33569;
assign w46973 = ~w4430 & ~w33603;
assign w46974 = ~w32096 & ~w3646;
assign w46975 = w32416 & w5745;
assign w46976 = w32415 & w33672;
assign w46977 = ~w32786 & w32995;
assign w46978 = ~w252 & w33816;
assign w46979 = w252 & w33818;
assign w46980 = w252 & ~w33815;
assign w46981 = ~w252 & w33815;
assign w46982 = ~w34121 & w49372;
assign w46983 = w35434 & ~w35441;
assign w46984 = w33855 & w7924;
assign w46985 = ~w53 & ~w55;
assign w46986 = ~w56 & w219;
assign w46987 = w56 & ~w219;
assign w46988 = ~w263 & ~w264;
assign w46989 = w251 & w271;
assign w46990 = w309 & w269;
assign w46991 = w751 & ~w796;
assign w46992 = w1335 & ~w80;
assign w46993 = ~w43939 & ~w1202;
assign w46994 = ~w43940 & ~w1485;
assign w46995 = ~w43941 & w1203;
assign w46996 = w1498 & w1493;
assign w46997 = w1492 & w3;
assign w46998 = ~w1492 & ~w3;
assign w46999 = w1474 & w80;
assign w47000 = ~w1474 & ~w80;
assign w47001 = ~w1479 & ~w57;
assign w47002 = w1479 & w57;
assign w47003 = ~w754 & w1370;
assign w47004 = (w1477 & w51429) | (w1477 & w51430) | (w51429 & w51430);
assign w47005 = (w1549 & w1698) | (w1549 & w51479) | (w1698 & w51479);
assign w47006 = w1705 & w1549;
assign w47007 = ~w1699 & ~w1748;
assign w47008 = ~w1647 & w1845;
assign w47009 = w1647 & ~w1845;
assign w47010 = w1594 & w1612;
assign w47011 = w43959 | w1645;
assign w47012 = (w1645 & w43959) | (w1645 & ~w1854) | (w43959 & ~w1854);
assign w47013 = w1612 & w52333;
assign w47014 = ~w1648 & w1902;
assign w47015 = ~w1906 & w39890;
assign w47016 = ~w1921 & w252;
assign w47017 = w1921 & ~w252;
assign w47018 = ~w1964 & ~w1757;
assign w47019 = ~w1862 & ~w1917;
assign w47020 = ~w2028 & w2022;
assign w47021 = w2028 & ~w2022;
assign w47022 = ~w2000 & ~w2093;
assign w47023 = ~w2241 & w1826;
assign w47024 = w2113 & a[97];
assign w47025 = ~w2113 & ~a[97];
assign w47026 = w2245 & ~w945;
assign w47027 = ~w2245 & w945;
assign w47028 = w39956 & w2389;
assign w47029 = ~w39956 & ~w2389;
assign w47030 = ~w2232 & w2278;
assign w47031 = ~w2399 & w2198;
assign w47032 = ~w2126 & ~w351;
assign w47033 = ~w2429 & w2259;
assign w47034 = ~w2457 & ~w2458;
assign w47035 = ~w2462 & ~w493;
assign w47036 = w2478 & w2130;
assign w47037 = ~w2298 & w57;
assign w47038 = ~w2680 & w80;
assign w47039 = w2571 & w52334;
assign w47040 = (w2864 & w48496) | (w2864 & w48497) | (w48496 & w48497);
assign w47041 = ~w2648 & ~w2643;
assign w47042 = w2785 & w351;
assign w47043 = ~w2785 & ~w351;
assign w47044 = w2680 & ~w2670;
assign w47045 = w2949 & w2670;
assign w47046 = w2958 & w52334;
assign w47047 = (w2864 & w51432) | (w2864 & w51433) | (w51432 & w51433);
assign w47048 = ~w2971 & w2771;
assign w47049 = ~w2977 & ~w2978;
assign w47050 = ~w2680 & ~w754;
assign w47051 = w2680 & w3006;
assign w47052 = w2971 & ~w1320;
assign w47053 = ~w3087 & w3086;
assign w47054 = w2680 & w3117;
assign w47055 = ~w3214 & ~w351;
assign w47056 = ~w3235 & w3234;
assign w47057 = w40046 | ~w1541;
assign w47058 = (~w1541 & w40046) | (~w1541 & w3115) | (w40046 & w3115);
assign w47059 = ~w3015 & w3234;
assign w47060 = w3163 & ~w3209;
assign w47061 = w2962 & w40091;
assign w47062 = ~w2944 & ~w2962;
assign w47063 = w3083 & w40102;
assign w47064 = w40103 & w3560;
assign w47065 = (w3560 & w40103) | (w3560 & ~w3083) | (w40103 & ~w3083);
assign w47066 = w3083 & ~w3573;
assign w47067 = ~w2876 & w51434;
assign w47068 = ~w40111 & w3491;
assign w47069 = ~w40110 & w3491;
assign w47070 = w40112 & w252;
assign w47071 = w40113 & w252;
assign w47072 = ~w40110 & w3490;
assign w47073 = ~w3631 & ~w3624;
assign w47074 = w3635 & ~w252;
assign w47075 = (~w3658 & w3645) | (~w3658 & w51435) | (w3645 & w51435);
assign w47076 = ~w3645 & w51436;
assign w47077 = w3846 & w3620;
assign w47078 = w3846 & ~w3464;
assign w47079 = w3857 & w3861;
assign w47080 = ~w3857 & w3863;
assign w47081 = w3884 & ~w3383;
assign w47082 = ~w3884 & w3383;
assign w47083 = ~w3857 & ~w3860;
assign w47084 = w3857 & w3860;
assign w47085 = w3910 & w3654;
assign w47086 = w3910 & w40115;
assign w47087 = w3519 & ~w3952;
assign w47088 = w3519 & w40135;
assign w47089 = w3409 & ~w3616;
assign w47090 = w4001 & w80;
assign w47091 = ~w3645 & w51437;
assign w47092 = w4140 & w4184;
assign w47093 = w4055 & w4327;
assign w47094 = w4185 & w40199;
assign w47095 = w4185 & ~w44129;
assign w47096 = (~w4436 & w4418) | (~w4436 & w48498) | (w4418 & w48498);
assign w47097 = ~w40202 & w4141;
assign w47098 = w4424 & ~w2285;
assign w47099 = w4531 & w2006;
assign w47100 = ~w4305 & w51438;
assign w47101 = ~w4372 & w4541;
assign w47102 = ~w4531 & ~w2006;
assign w47103 = w4558 & w4617;
assign w47104 = ~w4558 & w4619;
assign w47105 = ~w4390 & w4638;
assign w47106 = (w945 & w4681) | (w945 & w49373) | (w4681 & w49373);
assign w47107 = (w351 & w4689) | (w351 & w48499) | (w4689 & w48499);
assign w47108 = ~w4689 & w48500;
assign w47109 = ~w4430 & w48501;
assign w47110 = ~w4387 & ~w945;
assign w47111 = w4649 & w4739;
assign w47112 = ~w4114 & ~w42;
assign w47113 = w4114 & w42;
assign w47114 = w4754 & w48502;
assign w47115 = w4752 & w4111;
assign w47116 = (w4752 & w4443) | (w4752 & w48503) | (w4443 & w48503);
assign w47117 = w4794 & ~w4168;
assign w47118 = w4794 & ~w40217;
assign w47119 = ~w4794 & w4168;
assign w47120 = (w4693 & w47119) | (w4693 & w48504) | (w47119 & w48504);
assign w47121 = (~w252 & w4430) | (~w252 & w48505) | (w4430 & w48505);
assign w47122 = ~w44163 & ~w5350;
assign w47123 = ~w44167 & w5365;
assign w47124 = ~w5366 & w4056;
assign w47125 = ~w44168 & w5354;
assign w47126 = w44169 & ~w5372;
assign w47127 = ~w5329 & w5378;
assign w47128 = w5329 & w5354;
assign w47129 = w5366 & ~w4056;
assign w47130 = ~w5164 & ~w5503;
assign w47131 = w5931 & ~w2006;
assign w47132 = (w5705 & w6116) | (w5705 & w5719) | (w6116 & w5719);
assign w47133 = w6155 & ~w5691;
assign w47134 = (w6155 & w6116) | (w6155 & w47133) | (w6116 & w47133);
assign w47135 = ~w6123 & ~w44232;
assign w47136 = ~w6165 & ~w6297;
assign w47137 = ~w6165 & ~w44233;
assign w47138 = w6243 & w6056;
assign w47139 = ~w6243 & ~w6056;
assign w47140 = ~w6265 & w5960;
assign w47141 = ~w1120 & ~w6594;
assign w47142 = (w6254 & ~w6287) | (w6254 & w49374) | (~w6287 & w49374);
assign w47143 = ~w6673 & ~w6674;
assign w47144 = w6736 & ~w6538;
assign w47145 = (~w1320 & w6804) | (~w1320 & w49375) | (w6804 & w49375);
assign w47146 = ~w6834 & ~w6832;
assign w47147 = (~w6834 & ~w47144) | (~w6834 & w49376) | (~w47144 & w49376);
assign w47148 = w6829 & w6835;
assign w47149 = w6854 & ~w6853;
assign w47150 = (w6854 & ~w47144) | (w6854 & w49377) | (~w47144 & w49377);
assign w47151 = w47144 & w49378;
assign w47152 = w6880 & w6878;
assign w47153 = (w6880 & ~w47144) | (w6880 & w49379) | (~w47144 & w49379);
assign w47154 = a[75] & ~w6853;
assign w47155 = (a[75] & ~w47144) | (a[75] & w49380) | (~w47144 & w49380);
assign w47156 = w47144 & w49381;
assign w47157 = ~w5330 & ~w6883;
assign w47158 = (~w5330 & ~w47144) | (~w5330 & w49382) | (~w47144 & w49382);
assign w47159 = w6390 & w6878;
assign w47160 = (w6390 & ~w47144) | (w6390 & w49383) | (~w47144 & w49383);
assign w47161 = w47144 & w49384;
assign w47162 = w6441 & w6426;
assign w47163 = w6441 & ~w40449;
assign w47164 = ~w6432 & w6969;
assign w47165 = w47144 & w49385;
assign w47166 = w7016 & w2558;
assign w47167 = w7063 & w50165;
assign w47168 = ~w6985 & w7067;
assign w47169 = w7075 & w7081;
assign w47170 = ~w6457 & w50420;
assign w47171 = (w7093 & w6457) | (w7093 & w50421) | (w6457 & w50421);
assign w47172 = (w6737 & w49386) | (w6737 & w49387) | (w49386 & w49387);
assign w47173 = ~w6754 & ~w6769;
assign w47174 = ~w7145 & ~w6538;
assign w47175 = ~w7151 & w7150;
assign w47176 = w6538 & w47175;
assign w47177 = w7151 & ~w7150;
assign w47178 = (w7151 & ~w6538) | (w7151 & w47177) | (~w6538 & w47177);
assign w47179 = w7231 & ~w7229;
assign w47180 = (w7231 & ~w47144) | (w7231 & w49388) | (~w47144 & w49388);
assign w47181 = ~w7316 & ~w7314;
assign w47182 = ~w7316 & w7139;
assign w47183 = w7075 & w7331;
assign w47184 = w7333 & ~w7340;
assign w47185 = ~w7333 & w7340;
assign w47186 = ~w7343 & w7344;
assign w47187 = ~w7346 & w7314;
assign w47188 = ~w7346 & ~w7139;
assign w47189 = w7343 & ~w7009;
assign w47190 = w7343 & w7363;
assign w47191 = (w1320 & ~w7313) | (w1320 & w49389) | (~w7313 & w49389);
assign w47192 = ~w7068 & w48506;
assign w47193 = ~w7376 & ~w7378;
assign w47194 = (w7082 & w48507) | (w7082 & w48508) | (w48507 & w48508);
assign w47195 = (w7278 & w40479) | (w7278 & w7396) | (w40479 & w7396);
assign w47196 = ~w7396 & w40480;
assign w47197 = w7313 & w49390;
assign w47198 = (~w7276 & w7068) | (~w7276 & w48509) | (w7068 & w48509);
assign w47199 = w7418 & ~w7314;
assign w47200 = w7418 & w7139;
assign w47201 = w7343 & w7533;
assign w47202 = w6862 & ~w4056;
assign w47203 = ~w7139 & w48510;
assign w47204 = (w7747 & w7139) | (w7747 & w48511) | (w7139 & w48511);
assign w47205 = ~w7138 & w48512;
assign w47206 = ~w7784 & ~w400;
assign w47207 = w7784 & w400;
assign w47208 = (~w7846 & ~w7313) | (~w7846 & w49391) | (~w7313 & w49391);
assign w47209 = ~w7068 & w48513;
assign w47210 = w7241 & ~w44341;
assign w47211 = w7241 & ~w44342;
assign w47212 = w40540 & w7888;
assign w47213 = (w7138 & w48514) | (w7138 & w48515) | (w48514 & w48515);
assign w47214 = w7819 & ~w7900;
assign w47215 = ~w7923 & ~w7903;
assign w47216 = ~w7923 & ~w7543;
assign w47217 = ~w7374 & w7450;
assign w47218 = ~w7954 & ~w7955;
assign w47219 = w252 & ~w7439;
assign w47220 = (w252 & w7928) | (w252 & w48516) | (w7928 & w48516);
assign w47221 = (~w47216 & w48517) | (~w47216 & w48518) | (w48517 & w48518);
assign w47222 = w8148 & ~w7903;
assign w47223 = w8148 & ~w7543;
assign w47224 = w5745 & ~w44363;
assign w47225 = ~w7543 & w48519;
assign w47226 = w8597 & ~w8618;
assign w47227 = w8627 & ~w8631;
assign w47228 = ~w8621 & ~w8584;
assign w47229 = ~w8621 & w48520;
assign w47230 = (w8448 & w8621) | (w8448 & w48521) | (w8621 & w48521);
assign w47231 = w8694 & w8721;
assign w47232 = ~w8621 & w48522;
assign w47233 = (w8743 & w8621) | (w8743 & w48523) | (w8621 & w48523);
assign w47234 = w8188 & ~w8777;
assign w47235 = (w5745 & w8187) | (w5745 & w48524) | (w8187 & w48524);
assign w47236 = ~w8275 & w48525;
assign w47237 = ~w8793 & w44405;
assign w47238 = (w8793 & w8275) | (w8793 & w48526) | (w8275 & w48526);
assign w47239 = w8793 & ~w44405;
assign w47240 = ~w8621 & w48527;
assign w47241 = (~w8379 & w8621) | (~w8379 & w48528) | (w8621 & w48528);
assign w47242 = w8385 & w8276;
assign w47243 = w8385 & w44405;
assign w47244 = (w4056 & w8187) | (w4056 & w48529) | (w8187 & w48529);
assign w47245 = ~w8820 & w48530;
assign w47246 = (w8826 & w8820) | (w8826 & w48531) | (w8820 & w48531);
assign w47247 = ~w8621 & w48532;
assign w47248 = (w8848 & w8820) | (w8848 & w48533) | (w8820 & w48533);
assign w47249 = ~w8820 & w48534;
assign w47250 = ~w8621 & w49392;
assign w47251 = (w8858 & w8621) | (w8858 & w48535) | (w8621 & w48535);
assign w47252 = w8831 & w8880;
assign w47253 = ~w8187 & w48536;
assign w47254 = (~w8891 & w8187) | (~w8891 & w49945) | (w8187 & w49945);
assign w47255 = ~w8970 & ~w8735;
assign w47256 = ~w8882 & w8974;
assign w47257 = ~w8155 & ~w351;
assign w47258 = w9042 & w9105;
assign w47259 = w47258 & w49946;
assign w47260 = w9126 & ~w9028;
assign w47261 = ~w9175 & w9192;
assign w47262 = ~w8882 & w9210;
assign w47263 = ~w8882 & w9227;
assign w47264 = w8831 & ~w8867;
assign w47265 = ~w8855 & w48537;
assign w47266 = (~w9496 & w8855) | (~w9496 & w48538) | (w8855 & w48538);
assign w47267 = w8680 & ~w9178;
assign w47268 = ~w10467 & ~w10510;
assign w47269 = w10673 & ~w400;
assign w47270 = w11163 & ~w11166;
assign w47271 = w11163 & w11184;
assign w47272 = ~w11163 & w11186;
assign w47273 = ~w11204 & ~w493;
assign w47274 = ~w10673 & w10530;
assign w47275 = ~w11930 & w12039;
assign w47276 = ~w12336 & w12304;
assign w47277 = ~w12421 & w12413;
assign w47278 = w12421 & w12609;
assign w47279 = (~w10419 & ~w50187) | (~w10419 & w50592) | (~w50187 & w50592);
assign w47280 = w50187 & w50593;
assign w47281 = w12662 & w12675;
assign w47282 = w12065 & ~w12797;
assign w47283 = w12065 & ~w12583;
assign w47284 = ~w12065 & w12797;
assign w47285 = ~w12065 & w12583;
assign w47286 = ~w12030 & ~w12736;
assign w47287 = ~w12868 & w3646;
assign w47288 = w12839 & w3242;
assign w47289 = ~w12802 & w12827;
assign w47290 = ~w12112 & ~w12421;
assign w47291 = ~w12112 & ~w12613;
assign w47292 = ~w12862 & w12112;
assign w47293 = (w12960 & w50594) | (w12960 & w50595) | (w50594 & w50595);
assign w47294 = w12868 & ~w3646;
assign w47295 = ~w12985 & ~w12995;
assign w47296 = ~w12770 & ~w13102;
assign w47297 = ~w12583 & w50596;
assign w47298 = w400 & w13108;
assign w47299 = w12583 & w13240;
assign w47300 = w12583 & ~w13240;
assign w47301 = w13292 & w2006;
assign w47302 = ~w13292 & ~w2006;
assign w47303 = w12616 & w13362;
assign w47304 = ~w13363 & ~w400;
assign w47305 = (~w6769 & ~w12996) | (~w6769 & w50422) | (~w12996 & w50422);
assign w47306 = w12996 & w50423;
assign w47307 = (w13454 & ~w12996) | (w13454 & w50424) | (~w12996 & w50424);
assign w47308 = w12996 & w50425;
assign w47309 = (w12953 & ~w12996) | (w12953 & w50597) | (~w12996 & w50597);
assign w47310 = w47309 & w49393;
assign w47311 = (~w12824 & ~w12996) | (~w12824 & w50598) | (~w12996 & w50598);
assign w47312 = w47311 & w49394;
assign w47313 = (~w2558 & ~w12996) | (~w2558 & w50599) | (~w12996 & w50599);
assign w47314 = w13383 & w13539;
assign w47315 = (w13548 & ~w12996) | (w13548 & w50600) | (~w12996 & w50600);
assign w47316 = (w13555 & ~w12996) | (w13555 & w50601) | (~w12996 & w50601);
assign w47317 = (~w12855 & ~w12996) | (~w12855 & w50602) | (~w12996 & w50602);
assign w47318 = ~w13565 & ~w2558;
assign w47319 = (w13577 & ~w12996) | (w13577 & w50603) | (~w12996 & w50603);
assign w47320 = w13578 & ~w2896;
assign w47321 = w13565 & w2558;
assign w47322 = (w4838 & ~w47311) | (w4838 & w49395) | (~w47311 & w49395);
assign w47323 = (~w12980 & ~w12996) | (~w12980 & w50604) | (~w12996 & w50604);
assign w47324 = (~w4056 & ~w47323) | (~w4056 & w49396) | (~w47323 & w49396);
assign w47325 = (~w12871 & ~w12996) | (~w12871 & w50605) | (~w12996 & w50605);
assign w47326 = (w3242 & ~w47325) | (w3242 & w49397) | (~w47325 & w49397);
assign w47327 = (~w4430 & ~w47309) | (~w4430 & w49398) | (~w47309 & w49398);
assign w47328 = (w13649 & ~w12996) | (w13649 & w50426) | (~w12996 & w50426);
assign w47329 = w12996 & w50427;
assign w47330 = (w13664 & ~w12996) | (w13664 & w50428) | (~w12996 & w50428);
assign w47331 = w12996 & w50429;
assign w47332 = w47323 & w49399;
assign w47333 = (~w754 & ~w12996) | (~w754 & w50606) | (~w12996 & w50606);
assign w47334 = w47333 & w49400;
assign w47335 = (w13762 & ~w47333) | (w13762 & w49401) | (~w47333 & w49401);
assign w47336 = (~w13759 & ~w47333) | (~w13759 & w49402) | (~w47333 & w49402);
assign w47337 = w47333 & w49403;
assign w47338 = (~w493 & ~w12996) | (~w493 & w50607) | (~w12996 & w50607);
assign w47339 = w47338 & w49404;
assign w47340 = (w13796 & ~w47338) | (w13796 & w49405) | (~w47338 & w49405);
assign w47341 = w47338 & w49406;
assign w47342 = (w13802 & ~w47338) | (w13802 & w49407) | (~w47338 & w49407);
assign w47343 = (~w612 & ~w12996) | (~w612 & w50608) | (~w12996 & w50608);
assign w47344 = w47343 & w49408;
assign w47345 = (w13813 & ~w47343) | (w13813 & w49409) | (~w47343 & w49409);
assign w47346 = w12996 & w50609;
assign w47347 = (w13376 & ~w12996) | (w13376 & w50610) | (~w12996 & w50610);
assign w47348 = (~w351 & ~w12996) | (~w351 & w50611) | (~w12996 & w50611);
assign w47349 = w47348 & w49410;
assign w47350 = (w13891 & ~w47348) | (w13891 & w49411) | (~w47348 & w49411);
assign w47351 = w12996 & w50430;
assign w47352 = (w13198 & w48539) | (w13198 & w13471) | (w48539 & w13471);
assign w47353 = (~w3 & ~w12996) | (~w3 & w50431) | (~w12996 & w50431);
assign w47354 = (~w13267 & ~w12996) | (~w13267 & w50432) | (~w12996 & w50432);
assign w47355 = w47354 & w49412;
assign w47356 = (~w13302 & ~w12996) | (~w13302 & w50433) | (~w12996 & w50433);
assign w47357 = w47356 & w49413;
assign w47358 = (w13974 & ~w12996) | (w13974 & w50434) | (~w12996 & w50434);
assign w47359 = (~w1541 & ~w47354) | (~w1541 & w49414) | (~w47354 & w49414);
assign w47360 = (~w1738 & ~w47356) | (~w1738 & w49415) | (~w47356 & w49415);
assign w47361 = w47358 & w49416;
assign w47362 = (~w13888 & ~w47348) | (~w13888 & w50435) | (~w47348 & w50435);
assign w47363 = w47348 & w50436;
assign w47364 = ~w13932 & ~w14034;
assign w47365 = w13818 & ~w14031;
assign w47366 = ~w14075 & w13458;
assign w47367 = ~w14110 & ~w6264;
assign w47368 = w14116 & w14114;
assign w47369 = w14116 & w41193;
assign w47370 = ~w14119 & ~w14114;
assign w47371 = ~w14119 & ~w41193;
assign w47372 = w41194 & w6769;
assign w47373 = (w44745 & w49417) | (w44745 & w49418) | (w49417 & w49418);
assign w47374 = w14038 & w14132;
assign w47375 = w14139 & w5330;
assign w47376 = ~w14139 & ~w5330;
assign w47377 = w13417 & ~w5745;
assign w47378 = ~w13417 & w5745;
assign w47379 = w14038 & w14175;
assign w47380 = ~w14177 & ~w14135;
assign w47381 = w14197 & ~w4430;
assign w47382 = ~w14038 & w41209;
assign w47383 = ~w14533 & ~w14536;
assign w47384 = w14564 & ~w14550;
assign w47385 = w14519 & w14566;
assign w47386 = ~w13857 & w14037;
assign w47387 = w41261 & w14074;
assign w47388 = (w14074 & w41261) | (w14074 & ~w14568) | (w41261 & ~w14568);
assign w47389 = (w14033 & w13856) | (w14033 & w50612) | (w13856 & w50612);
assign w47390 = w41262 | ~w13932;
assign w47391 = (~w13932 & w41262) | (~w13932 & w14709) | (w41262 & w14709);
assign w47392 = ~w14728 & ~w44840;
assign w47393 = ~w14728 & ~w44841;
assign w47394 = w14038 & ~w13921;
assign w47395 = w14038 & w13921;
assign w47396 = w14766 & ~w14775;
assign w47397 = ~w14582 & w14778;
assign w47398 = ~w14796 & ~w14795;
assign w47399 = w14788 & w14798;
assign w47400 = ~w14783 & w48540;
assign w47401 = (w14804 & w14783) | (w14804 & w48541) | (w14783 & w48541);
assign w47402 = ~w14582 & w14686;
assign w47403 = w41270 & ~w14656;
assign w47404 = (~w252 & ~w47403) | (~w252 & w48542) | (~w47403 & w48542);
assign w47405 = ~w14823 & w14826;
assign w47406 = w14823 & w14828;
assign w47407 = w14580 & w14565;
assign w47408 = ~w14865 & w14879;
assign w47409 = ~w612 & ~w14885;
assign w47410 = ~w612 & ~w41275;
assign w47411 = ~w14872 & w41276;
assign w47412 = ~w14917 & ~w1120;
assign w47413 = w14832 & w14900;
assign w47414 = w14832 & ~w14966;
assign w47415 = w14819 & w252;
assign w47416 = ~w14783 & w48543;
assign w47417 = w14788 & ~w80;
assign w47418 = w14823 & w14989;
assign w47419 = ~w14823 & w14991;
assign w47420 = ~w15000 & w14737;
assign w47421 = w14974 & ~w14777;
assign w47422 = ~w14549 & w14763;
assign w47423 = w15028 & ~w1320;
assign w47424 = ~w41283 & w15034;
assign w47425 = ~w14545 & w14763;
assign w47426 = w15036 & w1541;
assign w47427 = ~w15035 & ~w1541;
assign w47428 = ~w14136 & ~w14184;
assign w47429 = ~w15181 & w4056;
assign w47430 = ~w15188 & w15187;
assign w47431 = w15188 & ~w15187;
assign w47432 = ~w15214 & w4838;
assign w47433 = w14170 & w15227;
assign w47434 = ~w14177 & ~w14103;
assign w47435 = ~w14177 & w44911;
assign w47436 = ~w15245 & ~w15246;
assign w47437 = w14097 & w15275;
assign w47438 = w14097 & ~w14418;
assign w47439 = ~w9781 & w14395;
assign w47440 = ~w9781 & w41299;
assign w47441 = ~w15331 & w8666;
assign w47442 = w15331 & ~w8666;
assign w47443 = w14759 & w15403;
assign w47444 = ~w15397 & ~w11870;
assign w47445 = ~w14582 & ~w15453;
assign w47446 = w15465 & ~w15460;
assign w47447 = ~w15450 & w15518;
assign w47448 = ~w15193 & w4056;
assign w47449 = w15624 & ~w14832;
assign w47450 = w15624 & ~w15621;
assign w47451 = ~w15058 & w15623;
assign w47452 = ~w15624 & ~w14777;
assign w47453 = (w15682 & w15677) | (w15682 & w48544) | (w15677 & w48544);
assign w47454 = (w15687 & w15677) | (w15687 & w48545) | (w15677 & w48545);
assign w47455 = ~w15677 & w48546;
assign w47456 = (w15694 & w15677) | (w15694 & w48547) | (w15677 & w48547);
assign w47457 = ~w15722 & w15721;
assign w47458 = ~w15724 & ~w11870;
assign w47459 = ~w15730 & w15729;
assign w47460 = w15680 & w15732;
assign w47461 = w15680 & w15719;
assign w47462 = ~w15680 & w15742;
assign w47463 = ~w15746 & ~w15745;
assign w47464 = w15680 & w15750;
assign w47465 = ~w15680 & w15752;
assign w47466 = ~w15761 & w15764;
assign w47467 = ~w15766 & ~w11138;
assign w47468 = w15680 & w15770;
assign w47469 = ~w15680 & w15772;
assign w47470 = w15766 & w11138;
assign w47471 = ~w15761 & w15779;
assign w47472 = ~w15788 & ~w15787;
assign w47473 = ~w14832 & ~w14995;
assign w47474 = ~w15680 & w15740;
assign w47475 = ~w15680 & ~w15820;
assign w47476 = ~w15680 & w15828;
assign w47477 = ~w15677 & w48548;
assign w47478 = ~w15832 & ~w15539;
assign w47479 = ~w15677 & w48549;
assign w47480 = ~w15672 & w48550;
assign w47481 = ~w15874 & w15876;
assign w47482 = w15874 & w15878;
assign w47483 = (~w7924 & w15672) | (~w7924 & w48551) | (w15672 & w48551);
assign w47484 = ~w15874 & w15908;
assign w47485 = w15874 & w15910;
assign w47486 = w15832 & w15183;
assign w47487 = w15832 & ~w15186;
assign w47488 = w15832 & w15196;
assign w47489 = w15943 & ~w3646;
assign w47490 = ~w15983 & ~w15985;
assign w47491 = w15680 & w4430;
assign w47492 = ~w15680 & w15980;
assign w47493 = ~w15271 & w15373;
assign w47494 = ~w16025 & ~w4838;
assign w47495 = w15680 & ~w15371;
assign w47496 = ~w16022 & w4838;
assign w47497 = w16114 & ~w15939;
assign w47498 = w15680 & ~w14881;
assign w47499 = w15058 & w16318;
assign w47500 = w15058 & w16317;
assign w47501 = ~w15680 & w16338;
assign w47502 = w15680 & w16341;
assign w47503 = ~w15680 & w16348;
assign w47504 = w15680 & w16351;
assign w47505 = ~w16359 & ~w16360;
assign w47506 = w15680 & w16363;
assign w47507 = ~w16305 & w16312;
assign w47508 = ~w16373 & ~w16374;
assign w47509 = w16390 & ~w16389;
assign w47510 = w16390 & ~w15575;
assign w47511 = w16397 & ~w16394;
assign w47512 = w16397 & ~w15575;
assign w47513 = ~w16391 & ~w16398;
assign w47514 = w15680 & w252;
assign w47515 = ~w16411 & w16413;
assign w47516 = w16411 & w16415;
assign w47517 = w16420 & w16428;
assign w47518 = ~w16420 & w16430;
assign w47519 = ~w16419 & ~w16435;
assign w47520 = w16419 & ~w16437;
assign w47521 = ~w16437 & ~w16423;
assign w47522 = ~w16437 & w15575;
assign w47523 = ~w16411 & w16446;
assign w47524 = w16556 & w400;
assign w47525 = ~w16556 & w57;
assign w47526 = w16727 & w16731;
assign w47527 = ~w16727 & w16733;
assign w47528 = ~w16751 & w3;
assign w47529 = ~w16772 & w57;
assign w47530 = w16727 & w16776;
assign w47531 = ~w16727 & w16778;
assign w47532 = ~w16750 & w48552;
assign w47533 = (w16788 & w16791) | (w16788 & w48553) | (w16791 & w48553);
assign w47534 = ~w16791 & w48554;
assign w47535 = ~w16757 & w49419;
assign w47536 = ~w16821 & ~w16823;
assign w47537 = w16556 & ~w16869;
assign w47538 = ~w16875 & w4430;
assign w47539 = w16556 & w41394;
assign w47540 = ~w16556 & w4430;
assign w47541 = ~w16978 & w16900;
assign w47542 = w16556 & ~w17001;
assign w47543 = w16556 & w17011;
assign w47544 = w16556 & w17035;
assign w47545 = w17048 & ~w17060;
assign w47546 = w16541 & w41413;
assign w47547 = w16541 & w41414;
assign w47548 = w17069 & ~w15824;
assign w47549 = ~w17075 & w6769;
assign w47550 = ~w17085 & ~w7315;
assign w47551 = ~w16556 & ~w15853;
assign w47552 = w17099 & w6264;
assign w47553 = ~w17118 & ~w17112;
assign w47554 = w41417 & w17112;
assign w47555 = w16556 & ~w17127;
assign w47556 = ~w17138 & w9781;
assign w47557 = ~w17118 & w17180;
assign w47558 = ~w17223 & w14039;
assign w47559 = ~w16799 & w16813;
assign w47560 = ~w16766 & w48555;
assign w47561 = w17354 & ~w17379;
assign w47562 = w17341 & w48556;
assign w47563 = w17345 & w17560;
assign w47564 = w17341 & w48557;
assign w47565 = w17580 & w17582;
assign w47566 = (w15681 & w17379) | (w15681 & w48558) | (w17379 & w48558);
assign w47567 = (w17598 & ~w17346) | (w17598 & w48559) | (~w17346 & w48559);
assign w47568 = (~w17607 & w17379) | (~w17607 & w48560) | (w17379 & w48560);
assign w47569 = ~w17644 & w16830;
assign w47570 = (w17651 & w17379) | (w17651 & w48561) | (w17379 & w48561);
assign w47571 = (w17659 & w17379) | (w17659 & w48562) | (w17379 & w48562);
assign w47572 = ~w17379 & w48563;
assign w47573 = (w17667 & w17379) | (w17667 & w48564) | (w17379 & w48564);
assign w47574 = ~w17379 & w48565;
assign w47575 = (w17672 & w17379) | (w17672 & w48566) | (w17379 & w48566);
assign w47576 = ~w17379 & w48567;
assign w47577 = (w17321 & w17379) | (w17321 & w48568) | (w17379 & w48568);
assign w47578 = ~w17666 & w17264;
assign w47579 = ~w17379 & w48569;
assign w47580 = w16891 & w17041;
assign w47581 = ~w17741 & ~w16968;
assign w47582 = ~w17354 & w16948;
assign w47583 = ~w17760 & ~w17044;
assign w47584 = ~w17776 & ~w17029;
assign w47585 = w17345 & w17779;
assign w47586 = w17769 & w2285;
assign w47587 = ~w17753 & w17810;
assign w47588 = ~w17740 & w48570;
assign w47589 = ~w17752 & w48571;
assign w47590 = ~w17849 & w17819;
assign w47591 = w17346 & w48572;
assign w47592 = w17849 & ~w17819;
assign w47593 = (w17849 & ~w17346) | (w17849 & w48573) | (~w17346 & w48573);
assign w47594 = (w17846 & w17752) | (w17846 & w48574) | (w17752 & w48574);
assign w47595 = w17753 & w17865;
assign w47596 = w17878 & w18155;
assign w47597 = ~w18172 & ~w18164;
assign w47598 = ~w18453 & w17887;
assign w47599 = ~w18453 & ~w17880;
assign w47600 = ~w18052 & ~w17861;
assign w47601 = w17878 & w18125;
assign w47602 = w17878 & w41578;
assign w47603 = w41579 & ~w18174;
assign w47604 = (~w18174 & w41579) | (~w18174 & ~w17878) | (w41579 & ~w17878);
assign w47605 = w17878 & w41580;
assign w47606 = w41581 & ~w18121;
assign w47607 = (~w18121 & w41581) | (~w18121 & ~w17878) | (w41581 & ~w17878);
assign w47608 = w18906 & w57;
assign w47609 = ~w18906 & ~w57;
assign w47610 = w19229 & w19237;
assign w47611 = w19229 & w18812;
assign w47612 = ~w20911 & ~w21542;
assign w47613 = ~w21777 & ~w2006;
assign w47614 = w21241 & w1320;
assign w47615 = w22011 & w22018;
assign w47616 = w22002 & w22005;
assign w47617 = ~w22002 & w22027;
assign w47618 = w22022 & w22007;
assign w47619 = w22022 & w41847;
assign w47620 = ~w22030 & ~w22038;
assign w47621 = w21709 & w22542;
assign w47622 = ~w21343 & w48575;
assign w47623 = w22629 & w21771;
assign w47624 = ~w21709 & ~w2558;
assign w47625 = w21709 & ~w22662;
assign w47626 = w22531 & w7315;
assign w47627 = w22744 & w22764;
assign w47628 = ~w22001 & ~w22066;
assign w47629 = ~w22203 & w48576;
assign w47630 = ~w252 & ~w22765;
assign w47631 = ~w22774 & w21821;
assign w47632 = w22774 & ~w21821;
assign w47633 = (~w22880 & w22835) | (~w22880 & w49420) | (w22835 & w49420);
assign w47634 = ~w22835 & w49421;
assign w47635 = w22879 & w22899;
assign w47636 = ~w22879 & w22901;
assign w47637 = w22906 & ~w22908;
assign w47638 = w23051 & w23057;
assign w47639 = ~w23246 & ~w23223;
assign w47640 = w23293 & ~w13384;
assign w47641 = ~w23293 & w13384;
assign w47642 = w22910 & ~w22815;
assign w47643 = w23416 & w23410;
assign w47644 = ~w23416 & ~w23410;
assign w47645 = ~w23425 & w2285;
assign w47646 = w23491 & w23496;
assign w47647 = ~w23503 & w23502;
assign w47648 = ~w23580 & ~w23631;
assign w47649 = ~w23641 & ~w21820;
assign w47650 = (~w23646 & w22203) | (~w23646 & w48577) | (w22203 & w48577);
assign w47651 = ~w23646 & w22765;
assign w47652 = (~w23689 & w22203) | (~w23689 & w48578) | (w22203 & w48578);
assign w47653 = ~w23689 & w22765;
assign w47654 = (w23689 & w22203) | (w23689 & w48579) | (w22203 & w48579);
assign w47655 = w23689 & w22765;
assign w47656 = ~w22203 & w48580;
assign w47657 = w493 & ~w22765;
assign w47658 = w23701 & w23700;
assign w47659 = ~w23701 & ~w23700;
assign w47660 = w23514 & ~w23748;
assign w47661 = ~w23767 & w23825;
assign w47662 = w23802 & w23741;
assign w47663 = ~w23320 & w23310;
assign w47664 = w23803 & ~w23912;
assign w47665 = w23842 & w23992;
assign w47666 = w23993 & ~w14039;
assign w47667 = w24001 & w23294;
assign w47668 = w24009 & w12666;
assign w47669 = ~w24009 & ~w12666;
assign w47670 = w24190 & w24185;
assign w47671 = w23842 & w24202;
assign w47672 = ~w23842 & ~w24205;
assign w47673 = ~w23842 & w23189;
assign w47674 = w24231 & ~w17380;
assign w47675 = w18183 & ~w23153;
assign w47676 = w18183 & ~w45336;
assign w47677 = w23153 & ~w18183;
assign w47678 = ~w24231 & w17380;
assign w47679 = (~w23499 & w45343) | (~w23499 & w24264) | (w45343 & w24264);
assign w47680 = (~w23499 & w45343) | (~w23499 & w23330) | (w45343 & w23330);
assign w47681 = ~w23355 & ~w23485;
assign w47682 = (~w22871 & w45355) | (~w22871 & w23051) | (w45355 & w23051);
assign w47683 = (~w22871 & w45355) | (~w22871 & w23330) | (w45355 & w23330);
assign w47684 = ~w24039 & ~w24540;
assign w47685 = ~w24976 & ~w24545;
assign w47686 = w24998 & ~w9195;
assign w47687 = ~w24998 & w9195;
assign w47688 = ~w25008 & ~w42109;
assign w47689 = ~w25008 & w24865;
assign w47690 = ~w25072 & w6264;
assign w47691 = ~w24985 & ~w6769;
assign w47692 = w24870 & ~w24176;
assign w47693 = w24871 & ~w25122;
assign w47694 = ~w25114 & w25104;
assign w47695 = w24870 & ~w25148;
assign w47696 = ~w24250 & ~w24198;
assign w47697 = w24871 & w25272;
assign w47698 = ~w42131 & ~w25303;
assign w47699 = ~w25305 & w16559;
assign w47700 = w25317 & w25323;
assign w47701 = ~w25332 & w42164;
assign w47702 = ~w25497 & w5330;
assign w47703 = w24864 & ~w25594;
assign w47704 = w24864 & w25594;
assign w47705 = w4056 & w24423;
assign w47706 = w4056 & w42192;
assign w47707 = w25607 & ~w25589;
assign w47708 = ~w25630 & ~w25632;
assign w47709 = ~w25728 & w24632;
assign w47710 = ~w25734 & ~w493;
assign w47711 = w25734 & w493;
assign w47712 = w25788 & w25840;
assign w47713 = w7924 & ~w26231;
assign w47714 = w26167 & w25319;
assign w47715 = ~w26167 & ~w25319;
assign w47716 = (~w25789 & w25056) | (~w25789 & w49947) | (w25056 & w49947);
assign w47717 = ~w26338 & ~w25611;
assign w47718 = ~w26347 & w4056;
assign w47719 = w26347 & ~w4056;
assign w47720 = w26382 & w26389;
assign w47721 = ~w26382 & w26391;
assign w47722 = w26382 & w26416;
assign w47723 = ~w26382 & w26418;
assign w47724 = w26459 & w26487;
assign w47725 = ~w26459 & w26486;
assign w47726 = ~w26459 & w26497;
assign w47727 = ~w25264 & ~w16559;
assign w47728 = w25264 & w16559;
assign w47729 = w25842 & w25283;
assign w47730 = ~w25842 & ~w25283;
assign w47731 = ~w25842 & ~w26612;
assign w47732 = w25842 & w26612;
assign w47733 = (~w26662 & w49948) | (~w26662 & w49949) | (w49948 & w49949);
assign w47734 = w25842 & w26681;
assign w47735 = ~w25842 & w26683;
assign w47736 = w26651 & ~w26664;
assign w47737 = w26771 & w25540;
assign w47738 = ~w26771 & w26772;
assign w47739 = ~w26771 & ~w2558;
assign w47740 = w26771 & w2558;
assign w47741 = ~w26077 & w48581;
assign w47742 = w26878 & ~w26707;
assign w47743 = ~w26048 & ~w42247;
assign w47744 = (~w26048 & w26894) | (~w26048 & w48582) | (w26894 & w48582);
assign w47745 = w26707 & w42249;
assign w47746 = w26707 & w27033;
assign w47747 = w26707 & ~w27037;
assign w47748 = (w27072 & ~w27008) | (w27072 & w48583) | (~w27008 & w48583);
assign w47749 = ~w27088 & w27091;
assign w47750 = w27088 & w26423;
assign w47751 = ~w27088 & w27094;
assign w47752 = w27088 & w26378;
assign w47753 = w26415 & ~w27109;
assign w47754 = w27008 & w48584;
assign w47755 = (w3242 & w26879) | (w3242 & w48585) | (w26879 & w48585);
assign w47756 = ~w26077 & w49950;
assign w47757 = w27267 & ~w26707;
assign w47758 = ~w27281 & ~w27280;
assign w47759 = ~w27335 & ~w27334;
assign w47760 = w22767 & w27336;
assign w47761 = ~w27358 & ~w27357;
assign w47762 = ~w27370 & ~w27369;
assign w47763 = ~w26077 & w49951;
assign w47764 = w27375 & ~w26707;
assign w47765 = ~w27376 & w49952;
assign w47766 = ~w27406 & ~w27405;
assign w47767 = ~w27432 & ~w27431;
assign w47768 = ~w27440 & w27439;
assign w47769 = ~w27493 & ~w27492;
assign w47770 = ~w27503 & ~w27502;
assign w47771 = ~w27609 & ~w27608;
assign w47772 = ~w27787 & ~w27786;
assign w47773 = ~w26077 & w48586;
assign w47774 = w27809 & ~w26707;
assign w47775 = w27105 & ~w27202;
assign w47776 = ~w27875 & w27905;
assign w47777 = ~w27954 & ~w27953;
assign w47778 = ~w26077 & w48587;
assign w47779 = w27957 & ~w26707;
assign w47780 = ~w26077 & w48588;
assign w47781 = w27971 & ~w26707;
assign w47782 = w27345 & ~w27385;
assign w47783 = w28297 & w28336;
assign w47784 = w28297 & w28341;
assign w47785 = ~w27746 & w49953;
assign w47786 = w28509 & ~w45703;
assign w47787 = ~w27746 & w49422;
assign w47788 = w27785 & ~w45703;
assign w47789 = ~w27746 & w49954;
assign w47790 = w27779 & ~w45705;
assign w47791 = ~w28564 & ~w27689;
assign w47792 = w28644 & ~w8666;
assign w47793 = ~w28607 & ~w28669;
assign w47794 = ~w28050 & w28964;
assign w47795 = ~w28973 & w28970;
assign w47796 = w28973 & ~w28970;
assign w47797 = ~w27823 & w49955;
assign w47798 = w29009 & w29011;
assign w47799 = w29023 & w2006;
assign w47800 = w28050 & w27190;
assign w47801 = ~w29017 & w27139;
assign w47802 = w29009 & w29050;
assign w47803 = ~w29051 & w29055;
assign w47804 = w29009 & w27893;
assign w47805 = w29010 & w27177;
assign w47806 = w29064 & w29068;
assign w47807 = w29044 & w2285;
assign w47808 = w29047 & w29035;
assign w47809 = ~w29010 & w29118;
assign w47810 = ~w29099 & ~w4056;
assign w47811 = ~w29354 & ~w28472;
assign w47812 = ~w29371 & ~w29370;
assign w47813 = ~w28311 & ~w11138;
assign w47814 = w28311 & w11138;
assign w47815 = ~w28328 & ~w28361;
assign w47816 = ~w29157 & ~w28372;
assign w47817 = w29624 & ~w9781;
assign w47818 = ~w29624 & w9781;
assign w47819 = w29586 & ~w9195;
assign w47820 = ~w29157 & w6769;
assign w47821 = ~w29669 & ~w29671;
assign w47822 = w29669 & w29671;
assign w47823 = w45798 & w29765;
assign w47824 = ~w29775 & ~w2558;
assign w47825 = w45807 & w29139;
assign w47826 = ~w29854 & w1541;
assign w47827 = w45820 & w29137;
assign w47828 = ~w30037 & w30038;
assign w47829 = ~w29159 & w30073;
assign w47830 = ~w30074 & w30072;
assign w47831 = ~w30074 & w30087;
assign w47832 = ~w29372 & w30095;
assign w47833 = w29372 & w30097;
assign w47834 = w29166 & ~w28738;
assign w47835 = ~w29157 & ~w28870;
assign w47836 = w29372 & ~w30094;
assign w47837 = ~w29372 & w30094;
assign w47838 = w30080 & w30132;
assign w47839 = ~w30080 & w30134;
assign w47840 = w30103 & w30138;
assign w47841 = ~w30103 & w30140;
assign w47842 = ~w42465 & w57;
assign w47843 = w29823 & w30339;
assign w47844 = ~w30303 & ~w29956;
assign w47845 = w30455 & ~w80;
assign w47846 = w30485 & w30487;
assign w47847 = ~w30485 & w30489;
assign w47848 = w30485 & w30493;
assign w47849 = ~w30485 & w30495;
assign w47850 = w30503 & w1120;
assign w47851 = w30351 & ~w612;
assign w47852 = ~w30145 & w30559;
assign w47853 = ~w30563 & w30560;
assign w47854 = ~w30145 & w30605;
assign w47855 = ~w30148 & ~w30621;
assign w47856 = w30629 & w30636;
assign w47857 = ~w30821 & w12666;
assign w47858 = ~w30841 & w30919;
assign w47859 = w30841 & w30921;
assign w47860 = w30947 & ~w29633;
assign w47861 = w30947 & ~w42522;
assign w47862 = w30958 & w45862;
assign w47863 = w30958 & w45863;
assign w47864 = ~w29664 & w30956;
assign w47865 = ~w29626 & w45870;
assign w47866 = ~w29626 & w45871;
assign w47867 = ~w29676 & w31076;
assign w47868 = ~w29676 & ~w31094;
assign w47869 = ~w29676 & ~w31112;
assign w47870 = ~w29676 & w31131;
assign w47871 = ~w29676 & ~w31133;
assign w47872 = w29823 & ~w2006;
assign w47873 = w29636 & w31248;
assign w47874 = ~w29793 & ~w31253;
assign w47875 = w29764 & ~w29808;
assign w47876 = w29636 & ~w31290;
assign w47877 = w29636 & w42568;
assign w47878 = w31355 & w31357;
assign w47879 = ~w31379 & ~w31380;
assign w47880 = w31379 & w31380;
assign w47881 = ~w31481 & ~w31406;
assign w47882 = w31364 & w31481;
assign w47883 = w31491 & w31493;
assign w47884 = ~w31491 & w30355;
assign w47885 = ~w31517 & ~w31520;
assign w47886 = ~w30353 & ~w31436;
assign w47887 = ~w30353 & w42591;
assign w47888 = ~w31536 & w31519;
assign w47889 = ~w31620 & w31622;
assign w47890 = w31620 & w31624;
assign w47891 = ~w31630 & w30811;
assign w47892 = w31630 & ~w30811;
assign w47893 = ~w31620 & w31647;
assign w47894 = w31620 & w31649;
assign w47895 = ~w31630 & w31652;
assign w47896 = w31630 & w31654;
assign w47897 = ~w31708 & w31709;
assign w47898 = w31708 & w31711;
assign w47899 = ~w31708 & w30892;
assign w47900 = w31708 & ~w30892;
assign w47901 = ~w31738 & w30932;
assign w47902 = w31738 & ~w30932;
assign w47903 = w30516 & w31436;
assign w47904 = w30516 & ~w31490;
assign w47905 = ~w31801 & w31814;
assign w47906 = ~w30457 & ~w30514;
assign w47907 = w31535 & w31845;
assign w47908 = ~w31842 & ~w31809;
assign w47909 = w31853 & ~w24874;
assign w47910 = w31825 & ~w23843;
assign w47911 = w31780 & w31863;
assign w47912 = ~w31780 & w31865;
assign w47913 = w31754 & w31884;
assign w47914 = ~w31754 & w31886;
assign w47915 = ~w30518 & w31900;
assign w47916 = w31475 & ~w31927;
assign w47917 = w31850 & w31920;
assign w47918 = ~w31849 & w31944;
assign w47919 = ~w31801 & w31949;
assign w47920 = ~w30518 & ~w31920;
assign w47921 = ~w31940 & w28077;
assign w47922 = ~w31491 & w31964;
assign w47923 = ~w30518 & a[15];
assign w47924 = ~w31491 & w31972;
assign w47925 = w31940 & ~w28077;
assign w47926 = ~w31853 & w24874;
assign w47927 = w31896 & ~w30750;
assign w47928 = ~w31896 & w30750;
assign w47929 = ~w31444 & w31404;
assign w47930 = w32078 & w32087;
assign w47931 = w32078 & w32098;
assign w47932 = ~w32151 & w32152;
assign w47933 = w32151 & w32154;
assign w47934 = ~w32151 & w32175;
assign w47935 = w32151 & w32177;
assign w47936 = ~w45927 & w32617;
assign w47937 = w45928 & ~w32627;
assign w47938 = ~w45928 & w32627;
assign w47939 = ~w32996 & ~w32790;
assign w47940 = w33088 & ~w33091;
assign w47941 = ~w33088 & w33091;
assign w47942 = ~w33149 & w33168;
assign w47943 = w33226 & ~w18183;
assign w47944 = ~w33239 & ~w33240;
assign w47945 = ~w33275 & ~w33247;
assign w47946 = ~w33226 & w18183;
assign w47947 = ~w31733 & ~w31576;
assign w47948 = w33510 & w33512;
assign w47949 = ~w32200 & w33572;
assign w47950 = ~w2896 & w32146;
assign w47951 = ~w2896 & ~w33573;
assign w47952 = w33718 & w33726;
assign w47953 = ~w33738 & ~w33737;
assign w47954 = w32998 & ~w3;
assign w47955 = ~w33754 & ~w33755;
assign w47956 = w33754 & w33755;
assign w47957 = w32719 & ~w32995;
assign w47958 = (w32994 & w47957) | (w32994 & w49423) | (w47957 & w49423);
assign w47959 = w33731 & w49424;
assign w47960 = (~w33766 & ~w33731) | (~w33766 & w49425) | (~w33731 & w49425);
assign w47961 = ~w33738 & w42686;
assign w47962 = ~w33738 & w42687;
assign w47963 = ~w32998 & ~w32750;
assign w47964 = ~w32998 & w351;
assign w47965 = ~w33993 & w33144;
assign w47966 = ~w33993 & ~w42713;
assign w47967 = w24874 & w33144;
assign w47968 = w24874 & ~w42713;
assign w47969 = w32996 & ~w34016;
assign w47970 = w32996 & w34019;
assign w47971 = w32996 & w34031;
assign w47972 = w33299 & w34141;
assign w47973 = ~w33299 & ~w34141;
assign w47974 = w33731 & ~w34195;
assign w47975 = ~w42744 & ~w33351;
assign w47976 = w34344 & ~w33659;
assign w47977 = w34344 & w42773;
assign w47978 = ~w42776 & ~w33670;
assign w47979 = ~w34426 & ~w34423;
assign w47980 = ~w34426 & w42789;
assign w47981 = w34434 & ~w33622;
assign w47982 = w34353 & w7924;
assign w47983 = ~w34353 & ~w7924;
assign w47984 = w32998 & ~w754;
assign w47985 = w32998 & ~w34640;
assign w47986 = w34622 & w34651;
assign w47987 = ~w34622 & w34653;
assign w47988 = ~w34637 & w34608;
assign w47989 = w32996 & w34687;
assign w47990 = w33453 & w34729;
assign w47991 = w33723 & w34769;
assign w47992 = ~w33718 & ~w34781;
assign w47993 = w34750 & w34808;
assign w47994 = ~w34870 & w34896;
assign w47995 = ~w34897 & ~w33855;
assign w47996 = ~w34897 & w34930;
assign w47997 = ~w34897 & w42876;
assign w47998 = ~w34931 & w49426;
assign w47999 = w42878 & w34949;
assign w48000 = (w34949 & w42878) | (w34949 & w34897) | (w42878 & w34897);
assign w48001 = ~w34897 & w42879;
assign w48002 = ~w34983 & w42881;
assign w48003 = ~w34983 & ~w34965;
assign w48004 = w34998 & ~w34892;
assign w48005 = w34998 & ~w42882;
assign w48006 = ~w35005 & ~w35003;
assign w48007 = ~w34871 & w35007;
assign w48008 = w35003 & ~w35014;
assign w48009 = w42884 & ~a[9];
assign w48010 = (~a[9] & w42884) | (~a[9] & w34897) | (w42884 & w34897);
assign w48011 = (w35029 & w34871) | (w35029 & w49427) | (w34871 & w49427);
assign w48012 = ~w35044 & w32698;
assign w48013 = w35044 & ~w32698;
assign w48014 = (w35060 & w35056) | (w35060 & w49428) | (w35056 & w49428);
assign w48015 = ~w35056 & w35067;
assign w48016 = ~w34897 & w42887;
assign w48017 = w33915 & w35079;
assign w48018 = ~w42888 & ~w33909;
assign w48019 = ~w42888 & w33909;
assign w48020 = (w29158 & w35056) | (w29158 & w49429) | (w35056 & w49429);
assign w48021 = w34988 & ~w35103;
assign w48022 = ~w34974 & ~w34959;
assign w48023 = ~w35092 & w35111;
assign w48024 = ~w35091 & w35135;
assign w48025 = w35057 & w35182;
assign w48026 = w42892 | ~w19040;
assign w48027 = (~w19040 & w42892) | (~w19040 & ~w35057) | (w42892 & ~w35057);
assign w48028 = ~w35192 & ~w35191;
assign w48029 = ~w34897 & w35198;
assign w48030 = ~w34897 & w42895;
assign w48031 = (w48030 & w49956) | (w48030 & w49957) | (w49956 & w49957);
assign w48032 = ~w34897 & w42900;
assign w48033 = (~w48030 & w49958) | (~w48030 & w49959) | (w49958 & w49959);
assign w48034 = ~w35266 & w35272;
assign w48035 = (~w35296 & w35282) | (~w35296 & w49430) | (w35282 & w49430);
assign w48036 = (w35311 & w35266) | (w35311 & w50166) | (w35266 & w50166);
assign w48037 = ~w34279 & w35314;
assign w48038 = w34878 & w34588;
assign w48039 = (~w34316 & w48038) | (~w34316 & w49431) | (w48038 & w49431);
assign w48040 = ~w34897 & w42905;
assign w48041 = (w48040 & w49960) | (w48040 & w49961) | (w49960 & w49961);
assign w48042 = (~w48040 & w49962) | (~w48040 & w49963) | (w49962 & w49963);
assign w48043 = w34900 & w49432;
assign w48044 = (w35449 & ~w34900) | (w35449 & w49433) | (~w34900 & w49433);
assign w48045 = ~w9781 & ~w34588;
assign w48046 = ~w9781 & w42903;
assign w48047 = w35496 & w35494;
assign w48048 = w35496 & ~w42920;
assign w48049 = w35498 & ~w35494;
assign w48050 = w35498 & w42920;
assign w48051 = w35520 & w35494;
assign w48052 = w35520 & ~w42920;
assign w48053 = w35522 & ~w35494;
assign w48054 = w35522 & w42920;
assign w48055 = w35540 & ~w35452;
assign w48056 = w35540 & w35481;
assign w48057 = ~w34216 & w35550;
assign w48058 = (~w34216 & w35550) | (~w34216 & w49435) | (w35550 & w49435);
assign w48059 = w34216 & ~w35550;
assign w48060 = ~w35550 & w49436;
assign w48061 = w35325 & w35611;
assign w48062 = ~w35136 & ~w35312;
assign w48063 = ~w35751 & ~w35750;
assign w48064 = w42954 & w35882;
assign w48065 = (w35882 & w42954) | (w35882 & w34897) | (w42954 & w34897);
assign w48066 = ~w34897 & w42955;
assign w48067 = w42959 & ~w34650;
assign w48068 = (~w34650 & w42959) | (~w34650 & w34897) | (w42959 & w34897);
assign w48069 = ~w34897 & w42960;
assign w48070 = w42961 & w35925;
assign w48071 = (w35925 & w42961) | (w35925 & w34897) | (w42961 & w34897);
assign w48072 = ~w35883 & w35938;
assign w48073 = ~w35982 & w35755;
assign w48074 = w35612 & w49437;
assign w48075 = w43023 | w36411;
assign w48076 = (w36411 & w43023) | (w36411 & w35980) | (w43023 & w35980);
assign w48077 = ~w36419 & ~w7315;
assign w48078 = w38338 & ~w38391;
assign w48079 = w38338 & w38495;
assign w48080 = w38609 & ~w13384;
assign w48081 = ~w39536 & w39542;
assign w48082 = ~w1302 & w400;
assign w48083 = ~w1867 & w612;
assign w48084 = w1867 & ~w612;
assign w48085 = w2034 & w80;
assign w48086 = ~w2034 & ~w80;
assign w48087 = w3730 & w3888;
assign w48088 = ~w4284 & w1738;
assign w48089 = w4431 & ~w4413;
assign w48090 = ~w40299 & w5811;
assign w48091 = w5743 & w6104;
assign w48092 = ~w40437 & ~w6822;
assign w48093 = ~w6767 & w6840;
assign w48094 = ~w6767 & w6969;
assign w48095 = ~w40451 & ~w7013;
assign w48096 = ~w6767 & w7140;
assign w48097 = w7333 & w49438;
assign w48098 = w8043 & ~w400;
assign w48099 = ~w8043 & w400;
assign w48100 = ~w8043 & w7439;
assign w48101 = ~w7775 & w7482;
assign w48102 = w8189 & w7945;
assign w48103 = ~w10868 & w11140;
assign w48104 = ~w12120 & w12123;
assign w48105 = w12182 & ~w12176;
assign w48106 = w12182 & w41030;
assign w48107 = ~w12318 & ~w12324;
assign w48108 = ~w12318 & w41060;
assign w48109 = (~w12624 & ~w12621) | (~w12624 & w50613) | (~w12621 & w50613);
assign w48110 = w12611 & w50437;
assign w48111 = ~w12614 & w12705;
assign w48112 = ~w12719 & ~w12720;
assign w48113 = (~w12736 & ~w12611) | (~w12736 & w50438) | (~w12611 & w50438);
assign w48114 = w12614 & w12915;
assign w48115 = w12614 & ~w12401;
assign w48116 = ~w12614 & w400;
assign w48117 = (w13171 & ~w12611) | (w13171 & w50439) | (~w12611 & w50439);
assign w48118 = ~w12614 & w12542;
assign w48119 = (w12527 & ~w12611) | (w12527 & w50440) | (~w12611 & w50440);
assign w48120 = w12614 & w13238;
assign w48121 = w12611 & w50441;
assign w48122 = w12611 & w50442;
assign w48123 = ~w12892 & w13333;
assign w48124 = ~w13981 & w14441;
assign w48125 = w46558 & w14074;
assign w48126 = (w14074 & w46558) | (w14074 & ~w14707) | (w46558 & ~w14707);
assign w48127 = w14616 & ~w14615;
assign w48128 = (~w14615 & w14616) | (~w14615 & ~w14779) | (w14616 & ~w14779);
assign w48129 = ~w14845 & w351;
assign w48130 = w12666 & w15640;
assign w48131 = ~w16643 & ~w945;
assign w48132 = w16643 & w945;
assign w48133 = w16082 & ~w16916;
assign w48134 = ~w17183 & ~w17123;
assign w48135 = ~w17413 & ~w9195;
assign w48136 = w17192 & w17351;
assign w48137 = w17192 & ~w17350;
assign w48138 = w17192 & ~w17531;
assign w48139 = ~w17192 & w17531;
assign w48140 = w17535 & ~w4838;
assign w48141 = w17192 & w17570;
assign w48142 = w17062 & w17819;
assign w48143 = w17062 & w17365;
assign w48144 = w17062 & ~w17361;
assign w48145 = w18451 & w18942;
assign w48146 = ~w18451 & w18023;
assign w48147 = w18451 & w18945;
assign w48148 = ~w18451 & w18165;
assign w48149 = w19870 & ~w19818;
assign w48150 = w19870 & w41728;
assign w48151 = ~w19764 & w19949;
assign w48152 = w19764 & w19951;
assign w48153 = ~w21241 & ~w21802;
assign w48154 = w21241 & w493;
assign w48155 = ~w21241 & ~w21858;
assign w48156 = ~w21241 & w21858;
assign w48157 = ~w21241 & w21419;
assign w48158 = w21587 & ~w21756;
assign w48159 = ~w21452 & ~w21792;
assign w48160 = w21877 & w21380;
assign w48161 = ~w21241 & w21824;
assign w48162 = w21241 & w57;
assign w48163 = w41831 & w21904;
assign w48164 = ~w41831 & ~w21904;
assign w48165 = w21241 & w22216;
assign w48166 = ~w21241 & w22218;
assign w48167 = w21241 & w22225;
assign w48168 = ~w21241 & w22224;
assign w48169 = ~w21241 & w22229;
assign w48170 = w21241 & w22221;
assign w48171 = ~w21241 & ~w22239;
assign w48172 = ~w21241 & ~w22255;
assign w48173 = w21241 & w21120;
assign w48174 = ~w21241 & w22280;
assign w48175 = ~w21241 & ~w22294;
assign w48176 = ~w21241 & ~w22457;
assign w48177 = ~w21241 & w22464;
assign w48178 = w21241 & ~w22659;
assign w48179 = w21584 & w22661;
assign w48180 = ~w21709 & w22681;
assign w48181 = w21709 & w22683;
assign w48182 = ~w21709 & w22691;
assign w48183 = w21709 & w22693;
assign w48184 = w21241 & ~w21350;
assign w48185 = w41958 & w3646;
assign w48186 = ~w22783 & w22791;
assign w48187 = ~w6264 & w5745;
assign w48188 = w22497 & ~w22479;
assign w48189 = w22852 & ~w6769;
assign w48190 = w23066 & w23071;
assign w48191 = ~w23066 & w22291;
assign w48192 = ~w21969 & ~w23108;
assign w48193 = ~w23150 & w22228;
assign w48194 = w23150 & ~w22228;
assign w48195 = w23160 & w23169;
assign w48196 = ~w23347 & w23051;
assign w48197 = ~w21970 & w43573;
assign w48198 = ~w21970 & w43574;
assign w48199 = ~w21970 & w43577;
assign w48200 = ~w21970 & w43578;
assign w48201 = ~w24684 & ~w24678;
assign w48202 = w24313 & w25387;
assign w48203 = ~w24864 & w1120;
assign w48204 = ~w24864 & w1541;
assign w48205 = w25504 & w25512;
assign w48206 = ~w24870 & ~w80;
assign w48207 = w24864 & w80;
assign w48208 = ~w26316 & w27143;
assign w48209 = w26316 & ~w27161;
assign w48210 = ~w42268 & w27163;
assign w48211 = w26067 & w26066;
assign w48212 = w26067 & w26826;
assign w48213 = w26938 & ~w26975;
assign w48214 = w43671 | w29054;
assign w48215 = (w29054 & w43671) | (w29054 & w29051) | (w43671 & w29051);
assign w48216 = ~w30145 & w30547;
assign w48217 = w30873 & w16559;
assign w48218 = ~w23843 & ~w34019;
assign w48219 = ~w23843 & ~w42718;
assign w48220 = w34034 & w34031;
assign w48221 = w34034 & w42721;
assign w48222 = w34036 & ~w34031;
assign w48223 = w34036 & ~w42721;
assign w48224 = w33129 & w34031;
assign w48225 = w33129 & w42721;
assign w48226 = ~w33129 & ~w34031;
assign w48227 = ~w33129 & ~w42721;
assign w48228 = w23843 & w34019;
assign w48229 = w23843 & w42718;
assign w48230 = w33855 & ~w34895;
assign w48231 = w33855 & ~w35002;
assign w48232 = w35022 & w35978;
assign w48233 = (w35022 & ~w35612) | (w35022 & w49439) | (~w35612 & w49439);
assign w48234 = w35612 & w49440;
assign w48235 = w35612 & w49441;
assign w48236 = w35612 & w49442;
assign w48237 = w36065 & w35978;
assign w48238 = (w36065 & ~w35612) | (w36065 & w49443) | (~w35612 & w49443);
assign w48239 = w35612 & w49444;
assign w48240 = w35612 & w49445;
assign w48241 = w35612 & w49446;
assign w48242 = w28077 & w35978;
assign w48243 = (w28077 & ~w35612) | (w28077 & w49447) | (~w35612 & w49447);
assign w48244 = w35612 & w49448;
assign w48245 = w35612 & w49449;
assign w48246 = w25851 & w35978;
assign w48247 = (w25851 & ~w35612) | (w25851 & w49450) | (~w35612 & w49450);
assign w48248 = w35612 & w49451;
assign w48249 = w35257 & w35978;
assign w48250 = (w35257 & ~w35612) | (w35257 & w49452) | (~w35612 & w49452);
assign w48251 = ~w35120 & w35978;
assign w48252 = (~w35120 & ~w35612) | (~w35120 & w49453) | (~w35612 & w49453);
assign w48253 = ~w36180 & ~w35978;
assign w48254 = ~w36180 & w35613;
assign w48255 = w35612 & w49454;
assign w48256 = w35612 & w49455;
assign w48257 = ~w2558 & w35978;
assign w48258 = (~w2558 & ~w35612) | (~w2558 & w49456) | (~w35612 & w49456);
assign w48259 = w43063 & w36692;
assign w48260 = ~w43063 & ~w36692;
assign w48261 = w35612 & w49457;
assign w48262 = ~w36754 & w35978;
assign w48263 = (~w36754 & ~w35612) | (~w36754 & w49458) | (~w35612 & w49458);
assign w48264 = w36754 & w35978;
assign w48265 = (w36754 & ~w35612) | (w36754 & w49459) | (~w35612 & w49459);
assign w48266 = w35612 & w49460;
assign w48267 = w4408 & ~w4111;
assign w48268 = w4670 & ~w4663;
assign w48269 = ~w43379 & w1320;
assign w48270 = w43378 & w6250;
assign w48271 = ~w43378 & w6252;
assign w48272 = w43389 & ~w754;
assign w48273 = (w7278 & ~w7100) | (w7278 & w49964) | (~w7100 & w49964);
assign w48274 = w7100 & w52104;
assign w48275 = w12896 & w4838;
assign w48276 = ~w16245 & w16565;
assign w48277 = w25352 & w2285;
assign w48278 = ~w26928 & w26065;
assign w48279 = ~w28036 & w49965;
assign w48280 = (~w27616 & w28036) | (~w27616 & w49966) | (w28036 & w49966);
assign w48281 = w28036 & ~w29092;
assign w48282 = w1507 & ~w1476;
assign w48283 = w1674 & w1687;
assign w48284 = ~w1674 & w1689;
assign w48285 = ~w2288 & ~w57;
assign w48286 = ~w43313 & w2808;
assign w48287 = a[95] & ~w2808;
assign w48288 = a[95] & ~w44021;
assign w48289 = ~w2845 & w2878;
assign w48290 = ~w2974 & w3060;
assign w48291 = ~w3507 & ~w2962;
assign w48292 = w3400 & ~w3663;
assign w48293 = w3400 & w3666;
assign w48294 = w3400 & ~w3675;
assign w48295 = w754 & w3704;
assign w48296 = w3813 & w3818;
assign w48297 = ~w3813 & ~w3818;
assign w48298 = w3871 & w3304;
assign w48299 = w3 & ~w3944;
assign w48300 = ~w3 & w3944;
assign w48301 = ~w4050 & w4083;
assign w48302 = ~w4050 & w3638;
assign w48303 = w3929 & w57;
assign w48304 = ~w4049 & w51332;
assign w48305 = w4319 & w4373;
assign w48306 = ~w4319 & w4375;
assign w48307 = ~w3929 & ~w57;
assign w48308 = ~w4445 & ~w42;
assign w48309 = w46875 | ~w6256;
assign w48310 = (~w6256 & w46875) | (~w6256 & w5833) | (w46875 & w5833);
assign w48311 = w6077 & ~w6228;
assign w48312 = ~w6243 & w4056;
assign w48313 = ~w7001 & w1541;
assign w48314 = w6767 & ~w7154;
assign w48315 = w7163 & w7197;
assign w48316 = ~w7163 & w7199;
assign w48317 = w7163 & w7212;
assign w48318 = ~w7163 & w7214;
assign w48319 = ~w6764 & ~w7246;
assign w48320 = ~w7247 & ~w42;
assign w48321 = w6318 & w49967;
assign w48322 = w7247 & w42;
assign w48323 = (w6796 & w40471) | (w6796 & ~w7086) | (w40471 & ~w7086);
assign w48324 = w7217 & w49461;
assign w48325 = ~w612 & ~w7267;
assign w48326 = (~w612 & ~w7217) | (~w612 & w49462) | (~w7217 & w49462);
assign w48327 = w7114 & ~w7267;
assign w48328 = (w7114 & ~w7217) | (w7114 & w49463) | (~w7217 & w49463);
assign w48329 = ~w7416 & ~w43405;
assign w48330 = ~w2558 & ~w7267;
assign w48331 = (~w2558 & ~w7217) | (~w2558 & w49464) | (~w7217 & w49464);
assign w48332 = w2285 & ~w7267;
assign w48333 = (w2285 & ~w7217) | (w2285 & w49465) | (~w7217 & w49465);
assign w48334 = w7555 & ~w7267;
assign w48335 = (w7555 & ~w7217) | (w7555 & w49466) | (~w7217 & w49466);
assign w48336 = ~w7584 & ~w7267;
assign w48337 = ~w7584 & ~w7218;
assign w48338 = w7595 & ~w7267;
assign w48339 = w7595 & ~w7218;
assign w48340 = w7606 & ~w7267;
assign w48341 = (w7606 & ~w7217) | (w7606 & w49467) | (~w7217 & w49467);
assign w48342 = w7617 & ~w7267;
assign w48343 = (w7617 & ~w7217) | (w7617 & w49468) | (~w7217 & w49468);
assign w48344 = w7630 & ~w7267;
assign w48345 = (w7630 & ~w7217) | (w7630 & w49469) | (~w7217 & w49469);
assign w48346 = w7652 & ~w7267;
assign w48347 = (w7652 & ~w7217) | (w7652 & w49470) | (~w7217 & w49470);
assign w48348 = ~w7660 & ~w7267;
assign w48349 = (~w7660 & ~w7217) | (~w7660 & w49471) | (~w7217 & w49471);
assign w48350 = ~w7718 & ~w7267;
assign w48351 = (~w7718 & ~w7217) | (~w7718 & w49472) | (~w7217 & w49472);
assign w48352 = w7728 & ~w7267;
assign w48353 = (w7728 & ~w7217) | (w7728 & w49473) | (~w7217 & w49473);
assign w48354 = w7797 & w7267;
assign w48355 = w7797 & w7218;
assign w48356 = (w7194 & w40526) | (w7194 & ~w7267) | (w40526 & ~w7267);
assign w48357 = (w7194 & w40526) | (w7194 & ~w7218) | (w40526 & ~w7218);
assign w48358 = w7290 & ~w7267;
assign w48359 = (w7290 & ~w7217) | (w7290 & w49474) | (~w7217 & w49474);
assign w48360 = ~w7444 & ~w7783;
assign w48361 = ~w7909 & ~w7820;
assign w48362 = w7904 & ~w2896;
assign w48363 = w44471 & w10464;
assign w48364 = ~w44471 & ~w10464;
assign w48365 = w11381 & w1738;
assign w48366 = w12227 & ~w945;
assign w48367 = ~w11489 & w754;
assign w48368 = w12614 & w13118;
assign w48369 = ~w13348 & w13256;
assign w48370 = w13491 & w13593;
assign w48371 = ~w13637 & ~w11870;
assign w48372 = w13637 & w11870;
assign w48373 = w13339 & w13088;
assign w48374 = w13876 & ~w13879;
assign w48375 = ~w13471 & w50443;
assign w48376 = (~w13917 & w13471) | (~w13917 & w50444) | (w13471 & w50444);
assign w48377 = w13849 & ~w14031;
assign w48378 = w41269 | ~w14615;
assign w48379 = (~w14615 & w41269) | (~w14615 & ~w14567) | (w41269 & ~w14567);
assign w48380 = w14567 & w14705;
assign w48381 = w41271 | w14670;
assign w48382 = (w14670 & w41271) | (w14670 & ~w14567) | (w41271 & ~w14567);
assign w48383 = ~w14567 & w14704;
assign w48384 = ~w1120 & w14905;
assign w48385 = w1120 & w14908;
assign w48386 = ~w1120 & w14927;
assign w48387 = w1120 & w14930;
assign w48388 = w945 & w14947;
assign w48389 = ~w945 & w14950;
assign w48390 = w14562 & w1738;
assign w48391 = w14223 & w2285;
assign w48392 = ~w14282 & w3242;
assign w48393 = w14282 & ~w3242;
assign w48394 = ~w15158 & w15173;
assign w48395 = w15158 & w15204;
assign w48396 = ~w15158 & w15206;
assign w48397 = ~w15158 & ~w14113;
assign w48398 = ~w14096 & ~w15305;
assign w48399 = w12666 & w15441;
assign w48400 = ~w14112 & ~w5745;
assign w48401 = ~w5745 & w15557;
assign w48402 = (w15608 & w41321) | (w15608 & w15602) | (w41321 & w15602);
assign w48403 = (w15605 & w41322) | (w15605 & w15602) | (w41322 & w15602);
assign w48404 = w15334 & ~w15374;
assign w48405 = ~w16510 & w3;
assign w48406 = w16510 & ~w3;
assign w48407 = ~w16530 & ~w16234;
assign w48408 = ~w17354 & w2285;
assign w48409 = ~w17062 & ~w17819;
assign w48410 = ~w18348 & ~w5330;
assign w48411 = ~w17879 & ~w1541;
assign w48412 = w20287 & w5330;
assign w48413 = ~w23527 & ~w23514;
assign w48414 = w23539 & w945;
assign w48415 = ~w612 & w23712;
assign w48416 = w612 & w23714;
assign w48417 = ~w21983 & w612;
assign w48418 = w612 & w23732;
assign w48419 = ~w612 & w23734;
assign w48420 = ~w23913 & ~w17380;
assign w48421 = w24271 & w43582;
assign w48422 = w23487 & ~w23488;
assign w48423 = (~w23996 & w42097) | (~w23996 & ~w24254) | (w42097 & ~w24254);
assign w48424 = ~w45434 & w14039;
assign w48425 = ~w25669 & w80;
assign w48426 = w25914 & ~w57;
assign w48427 = ~w25784 & w25429;
assign w48428 = ~w25970 & w400;
assign w48429 = ~w25990 & w25994;
assign w48430 = w25776 & w25748;
assign w48431 = ~w400 & ~w26006;
assign w48432 = ~w25435 & ~w26056;
assign w48433 = ~w22767 & ~w26495;
assign w48434 = ~w22767 & w45558;
assign w48435 = w26569 & w25306;
assign w48436 = ~w26569 & ~w25306;
assign w48437 = w25844 & w25093;
assign w48438 = ~w16559 & w25093;
assign w48439 = ~w16559 & w45577;
assign w48440 = ~w26707 & w26002;
assign w48441 = ~w26914 & w493;
assign w48442 = ~w26750 & ~w26078;
assign w48443 = ~w26750 & w45600;
assign w48444 = ~w945 & ~w26750;
assign w48445 = (w48443 & w49968) | (w48443 & w49969) | (w49968 & w49969);
assign w48446 = w27044 & w26078;
assign w48447 = w27044 & ~w45600;
assign w48448 = w1320 & ~w27062;
assign w48449 = w1320 & w45613;
assign w48450 = ~w26668 & w50167;
assign w48451 = ~w26668 & w50168;
assign w48452 = w27225 & w26078;
assign w48453 = w27225 & ~w45600;
assign w48454 = w26890 & w11870;
assign w48455 = w9781 & w27686;
assign w48456 = ~w26965 & w49970;
assign w48457 = w26876 & ~w26264;
assign w48458 = w26700 & w49971;
assign w48459 = w26700 & w49972;
assign w48460 = w26876 & ~w26038;
assign w48461 = w26876 & w27969;
assign w48462 = ~w25925 & w27929;
assign w48463 = ~w25925 & ~w45676;
assign w48464 = ~w80 & w28022;
assign w48465 = ~w27723 & w28508;
assign w48466 = (w28508 & w27605) | (w28508 & w49973) | (w27605 & w49973);
assign w48467 = ~w27723 & ~w27880;
assign w48468 = (~w27880 & w27605) | (~w27880 & w49974) | (w27605 & w49974);
assign w48469 = w26994 & w26939;
assign w48470 = ~w29016 & ~w27191;
assign w48471 = w29023 & ~w2285;
assign w48472 = ~w30145 & w28077;
assign w48473 = ~w3598 & w3759;
assign w48474 = ~w3598 & ~a[89];
assign w48475 = ~w3598 & w3786;
assign w48476 = ~w3598 & w3792;
assign w48477 = ~w3598 & w2558;
assign w48478 = ~w4049 & w51439;
assign w48479 = ~w4049 & w51440;
assign w48480 = ~w4049 & w51441;
assign w48481 = w6623 & w6735;
assign w48482 = w6769 & w15266;
assign w48483 = ~w6769 & w15268;
assign w48484 = w6769 & w15356;
assign w48485 = ~w6769 & w15358;
assign w48486 = ~w25393 & w1120;
assign w48487 = w28319 & w11138;
assign w48488 = ~w4463 & w3646;
assign w48489 = ~w4583 & w1738;
assign w48490 = w4583 & ~w1738;
assign w48491 = ~w4387 & w43360;
assign w48492 = ~w57 & w4808;
assign w48493 = w57 & w4810;
assign w48494 = w57 & w4824;
assign w48495 = ~w57 & w4826;
assign w48496 = ~w2571 & w80;
assign w48497 = ~w2571 & w47038;
assign w48498 = a[83] & ~w4436;
assign w48499 = ~w4405 & w351;
assign w48500 = w4405 & ~w351;
assign w48501 = w4714 & w252;
assign w48502 = w4114 & w4769;
assign w48503 = ~w43363 & w4752;
assign w48504 = ~w4794 & w43364;
assign w48505 = ~w4714 & ~w252;
assign w48506 = w7138 & w1320;
assign w48507 = w7394 & w49975;
assign w48508 = w7278 & w43401;
assign w48509 = ~w7138 & ~w7276;
assign w48510 = w7303 & w49475;
assign w48511 = (w7747 & ~w7303) | (w7747 & w49476) | (~w7303 & w49476);
assign w48512 = ~w7285 & w49477;
assign w48513 = w7138 & ~w7846;
assign w48514 = w40540 | w7888;
assign w48515 = (w7888 & w40540) | (w7888 & ~w7286) | (w40540 & ~w7286);
assign w48516 = ~w8038 & w252;
assign w48517 = ~w7438 & w44344;
assign w48518 = ~w7438 & ~w47215;
assign w48519 = ~w7781 & w5745;
assign w48520 = w8596 & w8428;
assign w48521 = ~w8596 & w8448;
assign w48522 = w8596 & w8741;
assign w48523 = ~w8596 & w8743;
assign w48524 = ~w8185 & w5745;
assign w48525 = ~w8274 & ~w8793;
assign w48526 = w8274 & w8793;
assign w48527 = w8596 & w8379;
assign w48528 = ~w8596 & ~w8379;
assign w48529 = ~w8185 & w4056;
assign w48530 = ~w8818 & w8824;
assign w48531 = w8818 & w8826;
assign w48532 = w8596 & ~w8316;
assign w48533 = w8818 & w8848;
assign w48534 = ~w8818 & w8850;
assign w48535 = ~w8596 & w8858;
assign w48536 = w8185 & w8886;
assign w48537 = w9500 & w9496;
assign w48538 = ~w9500 & ~w9496;
assign w48539 = w13353 & w13198;
assign w48540 = w14786 & w14802;
assign w48541 = ~w14786 & w14804;
assign w48542 = w14810 & ~w252;
assign w48543 = w14786 & w14985;
assign w48544 = w15679 & w15682;
assign w48545 = w15679 & w15687;
assign w48546 = ~w15679 & ~w15691;
assign w48547 = w15679 & w15694;
assign w48548 = ~w15679 & ~w15291;
assign w48549 = ~w15679 & w15333;
assign w48550 = w47479 & w7924;
assign w48551 = ~w47479 & ~w7924;
assign w48552 = w16751 & ~w3;
assign w48553 = ~w16792 & w16788;
assign w48554 = w16792 & ~w16788;
assign w48555 = ~w16758 & ~w57;
assign w48556 = w17344 & w16863;
assign w48557 = w17344 & ~w17569;
assign w48558 = ~w17590 & w15681;
assign w48559 = ~w17353 & w17598;
assign w48560 = w17610 & ~w17607;
assign w48561 = w17641 & w17651;
assign w48562 = w17656 & w17659;
assign w48563 = ~w17656 & w17661;
assign w48564 = ~w17665 & w17667;
assign w48565 = w17665 & w17669;
assign w48566 = w17656 & w17672;
assign w48567 = ~w17656 & w17674;
assign w48568 = w17641 & w17321;
assign w48569 = w17665 & ~w17264;
assign w48570 = w17046 & w16931;
assign w48571 = w17376 & ~w1738;
assign w48572 = w17353 & ~w17849;
assign w48573 = ~w17353 & w17849;
assign w48574 = ~w17376 & w17846;
assign w48575 = w21357 & w21584;
assign w48576 = w21970 & ~w252;
assign w48577 = ~w21970 & ~w23646;
assign w48578 = ~w21970 & ~w23689;
assign w48579 = ~w21970 & w23689;
assign w48580 = w21970 & w493;
assign w48581 = w26877 & ~w26826;
assign w48582 = ~w26002 & ~w26048;
assign w48583 = (w27072 & w26668) | (w27072 & w50169) | (w26668 & w50169);
assign w48584 = ~w26668 & w50170;
assign w48585 = (w3242 & w26078) | (w3242 & w49976) | (w26078 & w49976);
assign w48586 = w45648 & ~w26826;
assign w48587 = w45669 & ~w26826;
assign w48588 = w45670 & ~w26826;
assign w48589 = w1336 & ~w43942;
assign w48590 = w1336 & ~w1508;
assign w48591 = ~w44030 & w2880;
assign w48592 = w2882 & w2886;
assign w48593 = ~w2882 & w2888;
assign w48594 = ~w3668 & w3669;
assign w48595 = w3668 & w3671;
assign w48596 = w3546 & w3465;
assign w48597 = ~w3645 & w51442;
assign w48598 = (w3696 & w3645) | (w3696 & w51443) | (w3645 & w51443);
assign w48599 = w3689 & w3702;
assign w48600 = ~w3735 & w945;
assign w48601 = w3741 & ~w754;
assign w48602 = w3546 & w3755;
assign w48603 = ~w3921 & ~w945;
assign w48604 = ~w3546 & w3579;
assign w48605 = ~w4055 & w3685;
assign w48606 = w400 & ~w4179;
assign w48607 = ~w4055 & ~w612;
assign w48608 = w4055 & w40168;
assign w48609 = ~w4055 & w3743;
assign w48610 = w4201 & w612;
assign w48611 = ~w4319 & w4322;
assign w48612 = w4319 & w4325;
assign w48613 = w40187 | w3887;
assign w48614 = (w3887 & w40187) | (w3887 & ~w4055) | (w40187 & ~w4055);
assign w48615 = ~w945 & ~w4349;
assign w48616 = (w48614 & w51444) | (w48614 & w51445) | (w51444 & w51445);
assign w48617 = ~w612 & ~w4201;
assign w48618 = w3685 & w52335;
assign w48619 = ~w4092 & ~w4413;
assign w48620 = ~w4275 & ~w4268;
assign w48621 = ~w4448 & ~w4442;
assign w48622 = w4465 & ~w3646;
assign w48623 = ~w4418 & w4479;
assign w48624 = w4418 & w4481;
assign w48625 = ~w4418 & w4475;
assign w48626 = w4418 & ~w4478;
assign w48627 = w4275 & ~w4519;
assign w48628 = ~w4275 & w4519;
assign w48629 = ~w4497 & w4535;
assign w48630 = ~w4342 & w47101;
assign w48631 = w4418 & ~w4548;
assign w48632 = w4558 & w4560;
assign w48633 = ~w4558 & w4562;
assign w48634 = w4306 & w4292;
assign w48635 = ~w4299 & ~w4575;
assign w48636 = ~w4339 & ~w1541;
assign w48637 = w4418 & w4633;
assign w48638 = ~w4635 & w612;
assign w48639 = ~w4342 & w40210;
assign w48640 = w4418 & ~w4198;
assign w48641 = ~w4709 & w400;
assign w48642 = ~w4694 & w4718;
assign w48643 = w4549 & w1120;
assign w48644 = w4709 & ~w400;
assign w48645 = ~w40202 & w4755;
assign w48646 = ~w4765 & w4127;
assign w48647 = w4772 & ~w42;
assign w48648 = w4418 & w4150;
assign w48649 = ~w5330 & w49478;
assign w48650 = ~w5626 & ~w5629;
assign w48651 = w5329 & w754;
assign w48652 = w5642 & w5610;
assign w48653 = ~w5642 & ~w5610;
assign w48654 = ~w5527 & w5819;
assign w48655 = w5745 & w49479;
assign w48656 = w6065 & ~w6201;
assign w48657 = ~w6204 & ~w6203;
assign w48658 = ~w5843 & ~w6123;
assign w48659 = (~w6248 & w6255) | (~w6248 & w52105) | (w6255 & w52105);
assign w48660 = ~w6244 & w47136;
assign w48661 = ~w6244 & ~w6285;
assign w48662 = w6281 & w42;
assign w48663 = ~w6301 & w6308;
assign w48664 = ~w6262 & ~a[75];
assign w48665 = ~w6262 & ~w6368;
assign w48666 = w6243 & w6374;
assign w48667 = ~w6262 & w6378;
assign w48668 = ~w6262 & w6400;
assign w48669 = ~w6262 & w6419;
assign w48670 = ~w6262 & w6422;
assign w48671 = w6262 & w2285;
assign w48672 = ~w6262 & ~w6467;
assign w48673 = ~w6262 & ~w6481;
assign w48674 = w6262 & w2558;
assign w48675 = w6262 & ~w1738;
assign w48676 = ~w6509 & w6514;
assign w48677 = w6509 & w6516;
assign w48678 = w6262 & ~w2896;
assign w48679 = w6528 & ~w6531;
assign w48680 = ~w6528 & w6531;
assign w48681 = ~w6509 & w6545;
assign w48682 = w6509 & w6547;
assign w48683 = ~w6528 & w6552;
assign w48684 = w6528 & w6554;
assign w48685 = w6262 & w6073;
assign w48686 = w6262 & ~w1320;
assign w48687 = w6262 & ~w351;
assign w48688 = ~w6635 & w6638;
assign w48689 = w6635 & w6640;
assign w48690 = ~w6262 & ~w6648;
assign w48691 = ~w6635 & w6660;
assign w48692 = w6635 & w6662;
assign w48693 = ~w6575 & w754;
assign w48694 = ~w6599 & w6740;
assign w48695 = w6599 & w6742;
assign w48696 = ~w6774 & w6778;
assign w48697 = w6774 & w6780;
assign w48698 = w6784 & w6318;
assign w48699 = w6784 & w40434;
assign w48700 = ~w6774 & w6787;
assign w48701 = w6774 & w6789;
assign w48702 = w6793 & w6318;
assign w48703 = w6793 & w40434;
assign w48704 = w6817 & w6318;
assign w48705 = w6817 & w40434;
assign w48706 = ~w6425 & w6318;
assign w48707 = ~w6425 & w40434;
assign w48708 = ~w44258 & w6494;
assign w48709 = ~w6989 & w6318;
assign w48710 = (~w6762 & w48709) | (~w6762 & w52121) | (w48709 & w52121);
assign w48711 = (~w6737 & w52122) | (~w6737 & w52123) | (w52122 & w52123);
assign w48712 = ~w44258 & w7003;
assign w48713 = ~w7005 & ~w7006;
assign w48714 = w6521 & w7022;
assign w48715 = ~w6521 & ~w7022;
assign w48716 = w7035 & w6318;
assign w48717 = w7035 & w40434;
assign w48718 = w44261 & ~w7040;
assign w48719 = ~w44261 & w7040;
assign w48720 = w6995 & w1738;
assign w48721 = ~w7080 & ~w7081;
assign w48722 = ~w7080 & ~w7077;
assign w48723 = w7138 & ~w7067;
assign w48724 = w7138 & ~w6943;
assign w48725 = w6307 & w6622;
assign w48726 = ~w6717 & w6680;
assign w48727 = (w44307 & w44308) | (w44307 & ~w7067) | (w44308 & ~w7067);
assign w48728 = (w44307 & w44308) | (w44307 & ~w6943) | (w44308 & ~w6943);
assign w48729 = ~w7337 & ~w7331;
assign w48730 = ~w7337 & ~w7077;
assign w48731 = (w44316 & w44317) | (w44316 & ~w7067) | (w44317 & ~w7067);
assign w48732 = (w44316 & w44317) | (w44316 & ~w6943) | (w44317 & ~w6943);
assign w48733 = ~w40941 & ~w11142;
assign w48734 = w10673 & ~w351;
assign w48735 = w11154 & w11150;
assign w48736 = ~w11154 & ~w11150;
assign w48737 = w11333 & ~w3242;
assign w48738 = ~w40941 & w11791;
assign w48739 = ~w11794 & ~w11796;
assign w48740 = w11143 & w10464;
assign w48741 = ~w12076 & w12096;
assign w48742 = w41034 & ~w12204;
assign w48743 = (~w12204 & w41034) | (~w12204 & w11813) | (w41034 & w11813);
assign w48744 = ~w11424 & w11414;
assign w48745 = w11738 & w2006;
assign w48746 = ~w12721 & w7924;
assign w48747 = w12709 & ~w12809;
assign w48748 = w12203 & w12897;
assign w48749 = w12203 & w12901;
assign w48750 = w12203 & w12407;
assign w48751 = w12919 & w4430;
assign w48752 = (w12543 & w13161) | (w12543 & w50614) | (w13161 & w50614);
assign w48753 = w13175 & ~w13159;
assign w48754 = ~w13348 & w13257;
assign w48755 = ~w12693 & w44676;
assign w48756 = ~w12744 & w13407;
assign w48757 = ~w13471 & w13476;
assign w48758 = ~w13504 & ~w13507;
assign w48759 = w44700 & ~w13596;
assign w48760 = ~w44700 & w13596;
assign w48761 = ~w13655 & w11138;
assign w48762 = ~w13670 & w13678;
assign w48763 = (w13384 & w50445) | (w13384 & w50446) | (w50445 & w50446);
assign w48764 = ~w13471 & ~w13688;
assign w48765 = w754 & w13384;
assign w48766 = (w13779 & w13371) | (w13779 & w50447) | (w13371 & w50447);
assign w48767 = (w13781 & w13371) | (w13781 & w50448) | (w13371 & w50448);
assign w48768 = w13787 & w13780;
assign w48769 = w13787 & ~w44726;
assign w48770 = (w13820 & ~w13819) | (w13820 & w50449) | (~w13819 & w50449);
assign w48771 = w13913 & w13198;
assign w48772 = w13913 & w47352;
assign w48773 = (w41184 & ~w13819) | (w41184 & w50450) | (~w13819 & w50450);
assign w48774 = (~w252 & ~w13880) | (~w252 & w376) | (~w13880 & w376);
assign w48775 = w13679 & w14128;
assign w48776 = w14038 & w14180;
assign w48777 = ~w14456 & ~w14441;
assign w48778 = ~w14456 & ~w41223;
assign w48779 = ~w14038 & ~w14010;
assign w48780 = ~w14038 & w13969;
assign w48781 = w14532 & ~w14529;
assign w48782 = (w14532 & ~w13738) | (w14532 & w48781) | (~w13738 & w48781);
assign w48783 = w14038 & ~w14533;
assign w48784 = ~w41226 & w14535;
assign w48785 = ~w14528 & w1541;
assign w48786 = ~w14019 & w50621;
assign w48787 = ~w14650 & w14633;
assign w48788 = ~w14657 & ~w14691;
assign w48789 = ~w14766 & ~w14788;
assign w48790 = ~w400 & w14840;
assign w48791 = ~w400 & ~w44859;
assign w48792 = ~w14877 & w1120;
assign w48793 = w41279 | w14517;
assign w48794 = (w14517 & w41279) | (w14517 & w14872) | (w41279 & w14872);
assign w48795 = w400 & ~w14840;
assign w48796 = w400 & w44859;
assign w48797 = ~w15105 & ~w2558;
assign w48798 = ~w14263 & w44896;
assign w48799 = ~w14263 & ~w41288;
assign w48800 = ~w15088 & w15117;
assign w48801 = ~w6769 & w14765;
assign w48802 = ~w15245 & w15256;
assign w48803 = ~w15306 & ~w7924;
assign w48804 = w15160 & ~w15363;
assign w48805 = ~w15160 & w15363;
assign w48806 = w15306 & w7924;
assign w48807 = w15599 & ~w1738;
assign w48808 = w15015 & w15634;
assign w48809 = ~w15015 & w15636;
assign w48810 = ~w15643 & ~w15013;
assign w48811 = ~w15644 & w15647;
assign w48812 = ~w15684 & w14039;
assign w48813 = w14039 & w15687;
assign w48814 = w14039 & w47454;
assign w48815 = w15680 & w15707;
assign w48816 = ~w15817 & w7924;
assign w48817 = w15817 & ~w7924;
assign w48818 = w15533 & ~w15565;
assign w48819 = w15533 & w15566;
assign w48820 = ~w15833 & w15836;
assign w48821 = ~w15852 & ~w6769;
assign w48822 = w15856 & w15353;
assign w48823 = ~w15680 & ~w15867;
assign w48824 = w15902 & w15816;
assign w48825 = ~w15727 & w15777;
assign w48826 = ~w15854 & ~w15871;
assign w48827 = ~w15671 & w15539;
assign w48828 = ~w15671 & ~w5330;
assign w48829 = w15680 & w15578;
assign w48830 = w16061 & w2285;
assign w48831 = w16067 & ~w2558;
assign w48832 = w15680 & w16092;
assign w48833 = ~w16066 & w2558;
assign w48834 = ~w15680 & w15965;
assign w48835 = w15680 & ~w15152;
assign w48836 = ~w15680 & w16105;
assign w48837 = w15660 & w16118;
assign w48838 = w15680 & w15043;
assign w48839 = ~w16147 & w1320;
assign w48840 = ~w15680 & ~w16152;
assign w48841 = ~w16176 & ~w1541;
assign w48842 = ~w15680 & ~w16142;
assign w48843 = ~w15680 & w14968;
assign w48844 = ~w16196 & w945;
assign w48845 = w15680 & w16215;
assign w48846 = w16209 & w16214;
assign w48847 = ~w16209 & w16220;
assign w48848 = w15680 & w16223;
assign w48849 = w16176 & w1541;
assign w48850 = w15680 & ~w1320;
assign w48851 = w16235 & w16238;
assign w48852 = ~w16235 & w16240;
assign w48853 = ~w16032 & ~w16034;
assign w48854 = w15680 & ~w16259;
assign w48855 = ~w16266 & ~w16267;
assign w48856 = w15680 & w15576;
assign w48857 = w15680 & w16284;
assign w48858 = w15680 & w16289;
assign w48859 = ~w16083 & ~w16110;
assign w48860 = ~w16277 & ~w2006;
assign w48861 = ~w16359 & w16533;
assign w48862 = w16417 & ~w16526;
assign w48863 = ~w16366 & w16560;
assign w48864 = w16556 & w16571;
assign w48865 = ~w16556 & ~w16370;
assign w48866 = ~w16542 & w16433;
assign w48867 = ~w16585 & w351;
assign w48868 = w16556 & ~w16560;
assign w48869 = w16556 & ~w16566;
assign w48870 = w16114 & w41359;
assign w48871 = ~w16629 & w16623;
assign w48872 = w16556 & w16622;
assign w48873 = ~w16556 & w16673;
assign w48874 = ~w16669 & w16678;
assign w48875 = ~w16556 & w16685;
assign w48876 = ~w16669 & w16690;
assign w48877 = ~w41373 & w16697;
assign w48878 = w41373 & w16699;
assign w48879 = ~w16556 & w16269;
assign w48880 = ~w41373 & w16713;
assign w48881 = w41373 & w16715;
assign w48882 = ~w16667 & w16609;
assign w48883 = w16585 & ~w351;
assign w48884 = ~w41396 & w16896;
assign w48885 = w41396 & w16898;
assign w48886 = w16541 & ~w2285;
assign w48887 = w16523 & ~w16063;
assign w48888 = ~w16906 & ~w2006;
assign w48889 = w16556 & w16991;
assign w48890 = ~w17026 & w2896;
assign w48891 = w16964 & w2558;
assign w48892 = w16556 & w17168;
assign w48893 = w16541 & ~w17234;
assign w48894 = ~w17237 & ~w17236;
assign w48895 = w16541 & ~w17244;
assign w48896 = w16523 & ~w15681;
assign w48897 = w16523 & a[47];
assign w48898 = ~w16554 & ~w11138;
assign w48899 = w11138 & w15736;
assign w48900 = w11138 & w41353;
assign w48901 = w41352 & w11138;
assign w48902 = w16523 & w11870;
assign w48903 = w15714 & w11870;
assign w48904 = ~w16556 & ~w16269;
assign w48905 = w17275 & w17381;
assign w48906 = ~w17402 & w17159;
assign w48907 = w17402 & ~w17159;
assign w48908 = ~w17402 & w17417;
assign w48909 = w17402 & w17419;
assign w48910 = ~w17396 & w17426;
assign w48911 = ~w17442 & ~w17190;
assign w48912 = ~w17191 & ~w17089;
assign w48913 = w17491 & w17493;
assign w48914 = ~w17491 & w17495;
assign w48915 = w17491 & w17500;
assign w48916 = ~w17491 & w17502;
assign w48917 = w17559 & ~w17560;
assign w48918 = w17559 & w41450;
assign w48919 = ~w17559 & w17560;
assign w48920 = ~w17559 & ~w41450;
assign w48921 = ~w17504 & w17497;
assign w48922 = w17594 & w14766;
assign w48923 = ~w17643 & w16592;
assign w48924 = w17378 & w17665;
assign w48925 = ~w17679 & ~w11870;
assign w48926 = ~w17693 & w17217;
assign w48927 = w17693 & ~w17217;
assign w48928 = w16891 & ~w16998;
assign w48929 = ~w17778 & ~w17779;
assign w48930 = ~w17778 & w41450;
assign w48931 = w17354 & ~w17753;
assign w48932 = w45004 & ~w17779;
assign w48933 = w45004 & w41450;
assign w48934 = ~w47587 & ~w17809;
assign w48935 = ~w17811 & ~w2896;
assign w48936 = ~w17852 & w1120;
assign w48937 = ~w17859 & w17876;
assign w48938 = w17998 & w18000;
assign w48939 = ~w17998 & w18002;
assign w48940 = w17998 & w18007;
assign w48941 = ~w17998 & w18009;
assign w48942 = w17842 & w18053;
assign w48943 = ~w17380 & w16655;
assign w48944 = ~w18094 & w612;
assign w48945 = ~w18102 & w16692;
assign w48946 = w19039 & ~w18788;
assign w48947 = ~w19052 & w19054;
assign w48948 = w18840 & ~w18844;
assign w48949 = w19039 & w18845;
assign w48950 = ~w19858 & w19860;
assign w48951 = w19858 & w19862;
assign w48952 = ~w41730 & w19866;
assign w48953 = w41730 & w19869;
assign w48954 = ~w19894 & ~w252;
assign w48955 = ~w19285 & w1320;
assign w48956 = w19061 & w612;
assign w48957 = ~w19799 & ~w19977;
assign w48958 = w19799 & w19977;
assign w48959 = ~w19998 & w20455;
assign w48960 = ~w20561 & w20618;
assign w48961 = ~w20913 & w20967;
assign w48962 = ~w20913 & w20978;
assign w48963 = ~w20979 & w12666;
assign w48964 = ~w20913 & w20995;
assign w48965 = ~w20996 & w14039;
assign w48966 = w20979 & ~w12666;
assign w48967 = ~w20913 & ~w21090;
assign w48968 = ~w20913 & w21096;
assign w48969 = ~w21105 & w20525;
assign w48970 = w21105 & ~w20525;
assign w48971 = w21100 & w15681;
assign w48972 = w20996 & ~w14039;
assign w48973 = w21217 & ~w21238;
assign w48974 = ~w21709 & w20923;
assign w48975 = ~w21803 & ~w21815;
assign w48976 = w21822 & ~w21747;
assign w48977 = ~w21850 & ~w21852;
assign w48978 = w21850 & w21852;
assign w48979 = w21859 & w351;
assign w48980 = w21241 & ~w612;
assign w48981 = w21358 & w21874;
assign w48982 = ~w21822 & w21703;
assign w48983 = ~w21893 & w21899;
assign w48984 = w21893 & w21901;
assign w48985 = ~w21906 & w21909;
assign w48986 = ~w21859 & ~w351;
assign w48987 = w21709 & w21973;
assign w48988 = w21709 & w21980;
assign w48989 = ~w21038 & ~w22255;
assign w48990 = ~w21038 & w41890;
assign w48991 = w22297 & ~w22294;
assign w48992 = w22297 & w41893;
assign w48993 = ~w21709 & w20960;
assign w48994 = ~w41909 & w22434;
assign w48995 = w21709 & w22440;
assign w48996 = ~w22443 & ~w22444;
assign w48997 = w22461 & ~w22457;
assign w48998 = w22461 & w41913;
assign w48999 = w22468 & w22464;
assign w49000 = w22468 & w41914;
assign w49001 = w22394 & w11138;
assign w49002 = ~w22479 & ~w22433;
assign w49003 = w41949 & ~w2896;
assign w49004 = ~w21251 & w21749;
assign w49005 = ~w21709 & ~w21352;
assign w49006 = ~w22701 & ~w3646;
assign w49007 = w22783 & ~w22304;
assign w49008 = ~w22796 & ~w22797;
assign w49009 = w22818 & w22820;
assign w49010 = w22823 & w6264;
assign w49011 = w22070 & ~w22546;
assign w49012 = w21970 & ~w5330;
assign w49013 = w22897 & w6027;
assign w49014 = ~w22897 & ~w4838;
assign w49015 = w21970 & ~w22924;
assign w49016 = ~w10419 & w22479;
assign w49017 = ~w10419 & ~w41976;
assign w49018 = ~w21969 & w22939;
assign w49019 = ~w22497 & w22387;
assign w49020 = ~w22955 & ~w22954;
assign w49021 = w21970 & ~w22964;
assign w49022 = ~w21969 & w22971;
assign w49023 = ~w23007 & ~w23006;
assign w49024 = w6027 | w4838;
assign w49025 = (w4838 & w6027) | (w4838 & w22897) | (w6027 & w22897);
assign w49026 = w21970 & w23095;
assign w49027 = w21931 & w21952;
assign w49028 = ~w23098 & w21968;
assign w49029 = w23099 & ~w23102;
assign w49030 = ~w41995 & ~w23109;
assign w49031 = ~w21970 & w23122;
assign w49032 = w21970 & w23118;
assign w49033 = ~w21970 & ~w23160;
assign w49034 = w22070 & ~w23208;
assign w49035 = w42020 & w23412;
assign w49036 = (w23412 & w42020) | (w23412 & ~w22477) | (w42020 & ~w22477);
assign w49037 = w21970 & w3242;
assign w49038 = ~w22740 & ~w23478;
assign w49039 = w22740 & w23478;
assign w49040 = w23482 & w3646;
assign w49041 = w23466 & ~w23469;
assign w49042 = ~w22897 & w42024;
assign w49043 = w23509 & w23506;
assign w49044 = ~w23509 & ~w23506;
assign w49045 = ~w23520 & ~w22135;
assign w49046 = ~w23540 & w1009;
assign w49047 = ~w23540 & ~w945;
assign w49048 = ~w23641 & w21931;
assign w49049 = w23665 & w3;
assign w49050 = w22064 & w21891;
assign w49051 = ~w23743 & ~w23684;
assign w49052 = w400 & ~w45296;
assign w49053 = w45282 & ~w23750;
assign w49054 = w23449 & ~w24263;
assign w49055 = ~w24275 & ~w24276;
assign w49056 = w24284 & w23420;
assign w49057 = ~w24284 & ~w23420;
assign w49058 = ~w23842 & w1541;
assign w49059 = w23842 & w24292;
assign w49060 = ~w24301 & ~w24302;
assign w49061 = ~w23842 & w24308;
assign w49062 = w24306 & w1541;
assign w49063 = ~w24320 & w24318;
assign w49064 = w24320 & ~w24318;
assign w49065 = ~w23842 & w23393;
assign w49066 = w23487 & ~w24267;
assign w49067 = w23487 & w42050;
assign w49068 = ~w3242 & ~w23485;
assign w49069 = ~w3242 & ~w45344;
assign w49070 = ~w23914 & w24334;
assign w49071 = w24335 & ~w23487;
assign w49072 = ~w23348 & w23052;
assign w49073 = ~w24399 & ~w24402;
assign w49074 = ~w23842 & w22799;
assign w49075 = ~w24415 & ~w4056;
assign w49076 = ~w24324 & ~w1738;
assign w49077 = ~w24305 & ~w1541;
assign w49078 = w24594 & ~w24596;
assign w49079 = ~w23808 & w23696;
assign w49080 = w24870 & w23986;
assign w49081 = w25173 & ~w25226;
assign w49082 = w24871 & w25229;
assign w49083 = ~w24357 & ~w24343;
assign w49084 = ~w24489 & ~w24424;
assign w49085 = ~w25352 & ~w25350;
assign w49086 = ~w25352 & ~w42136;
assign w49087 = w25364 & ~w24288;
assign w49088 = w25364 & w42139;
assign w49089 = ~w24871 & w24279;
assign w49090 = ~w25370 & w1738;
assign w49091 = ~w25377 & w1541;
assign w49092 = w24864 & ~w24299;
assign w49093 = w42146 & w1120;
assign w49094 = (w1120 & w42146) | (w1120 & ~w24557) | (w42146 & ~w24557);
assign w49095 = w25370 & ~w1738;
assign w49096 = w25399 & ~w25401;
assign w49097 = w25641 & w3;
assign w49098 = ~w24783 & ~w3;
assign w49099 = w24783 & ~w3;
assign w49100 = ~w25710 & w25709;
assign w49101 = w25785 & ~w25720;
assign w49102 = w24831 & w23863;
assign w49103 = w24831 & ~w42072;
assign w49104 = ~w25860 & w25699;
assign w49105 = ~w24885 & ~w25833;
assign w49106 = ~w25901 & w25904;
assign w49107 = w25900 & ~w25765;
assign w49108 = ~w25900 & w25765;
assign w49109 = ~w25967 & ~w25766;
assign w49110 = ~w25844 & w25776;
assign w49111 = w25850 & ~w351;
assign w49112 = w26023 & w26026;
assign w49113 = ~w26023 & w26028;
assign w49114 = w26023 & w26039;
assign w49115 = ~w26023 & w26041;
assign w49116 = w25842 & w24956;
assign w49117 = ~w25842 & ~w24956;
assign w49118 = ~w25325 & ~w24966;
assign w49119 = w25788 & w26162;
assign w49120 = w25788 & w26212;
assign w49121 = w25788 & w26220;
assign w49122 = w25788 & w26383;
assign w49123 = ~w26395 & w25514;
assign w49124 = ~w26395 & w26410;
assign w49125 = w26411 & ~w4838;
assign w49126 = w25802 & w25849;
assign w49127 = ~w25844 & w25212;
assign w49128 = w45555 | w26447;
assign w49129 = (w26447 & w45555) | (w26447 & w26459) | (w45555 & w26459);
assign w49130 = w25788 & w45556;
assign w49131 = ~w26574 & w25312;
assign w49132 = ~w26574 & ~w42229;
assign w49133 = ~w26587 & ~w26586;
assign w49134 = w25259 & w25128;
assign w49135 = w25788 & w26630;
assign w49136 = w25788 & w26633;
assign w49137 = ~w26643 & w17380;
assign w49138 = ~w26804 & ~w26805;
assign w49139 = w26838 & w26802;
assign w49140 = ~w26907 & w26994;
assign w49141 = w42256 & w27027;
assign w49142 = (w27027 & w42256) | (w27027 & ~w26722) | (w42256 & ~w26722);
assign w49143 = w26722 & w42257;
assign w49144 = w26877 & ~w26306;
assign w49145 = ~w26295 & ~w27789;
assign w49146 = ~w27790 & w49145;
assign w49147 = ~w27794 & w27786;
assign w49148 = ~w27794 & ~w26827;
assign w49149 = ~w27796 & w27799;
assign w49150 = w27796 & w27802;
assign w49151 = ~w27812 & w27814;
assign w49152 = w27808 & w27818;
assign w49153 = w27812 & w27817;
assign w49154 = w27822 & ~w27831;
assign w49155 = w27808 & w27842;
assign w49156 = w27823 & w49977;
assign w49157 = w27784 & w49978;
assign w49158 = w26877 & ~w26021;
assign w49159 = w27906 & ~w28050;
assign w49160 = w28085 & w52336;
assign w49161 = w28067 & w28039;
assign w49162 = w28067 & w27258;
assign w49163 = ~w28102 & ~w28091;
assign w49164 = w25851 & w24874;
assign w49165 = w27339 & w28039;
assign w49166 = w27339 & w27258;
assign w49167 = w27949 & ~w27339;
assign w49168 = (~w28049 & w50171) | (~w28049 & w50172) | (w50171 & w50172);
assign w49169 = w27311 & w28039;
assign w49170 = w27311 & w27258;
assign w49171 = ~w22767 & w28193;
assign w49172 = (~w22767 & w28192) | (~w22767 & w49979) | (w28192 & w49979);
assign w49173 = w22767 & ~w28193;
assign w49174 = ~w28192 & w49980;
assign w49175 = w15681 & w27646;
assign w49176 = ~w15681 & w27585;
assign w49177 = ~w42351 & ~w28351;
assign w49178 = ~w12666 & w28352;
assign w49179 = w27585 & w28039;
assign w49180 = w26978 & w50248;
assign w49181 = w27401 & w28039;
assign w49182 = w26978 & w50249;
assign w49183 = w28467 & ~w16559;
assign w49184 = w27822 & w47786;
assign w49185 = w27822 & ~w45704;
assign w49186 = w42367 & ~w28511;
assign w49187 = w28516 & ~w4838;
assign w49188 = (w28516 & w28049) | (w28516 & w49983) | (w28049 & w49983);
assign w49189 = w28519 & w4838;
assign w49190 = ~w28049 & w49984;
assign w49191 = w28534 & ~w4838;
assign w49192 = (w28534 & w28049) | (w28534 & w49985) | (w28049 & w49985);
assign w49193 = w28537 & w4838;
assign w49194 = ~w28049 & w49986;
assign w49195 = ~w42376 & w27722;
assign w49196 = w28582 & w47790;
assign w49197 = w28582 & ~w45706;
assign w49198 = w28588 & ~w28598;
assign w49199 = w28562 & ~w28612;
assign w49200 = w28683 & ~w28066;
assign w49201 = w28695 & w28697;
assign w49202 = ~w28695 & w28699;
assign w49203 = w27906 & ~w28745;
assign w49204 = ~w28714 & ~w252;
assign w49205 = w28010 & w52337;
assign w49206 = ~w28946 & ~w28947;
assign w49207 = w28946 & w28947;
assign w49208 = ~w42415 & w28994;
assign w49209 = ~w28990 & ~w1320;
assign w49210 = ~w29005 & ~w28951;
assign w49211 = ~w28998 & ~w28951;
assign w49212 = ~w29026 & ~w29022;
assign w49213 = w29136 & ~w29138;
assign w49214 = (w28884 & ~w28855) | (w28884 & w49987) | (~w28855 & w49987);
assign w49215 = ~w28920 & w49988;
assign w49216 = (~w29208 & w28920) | (~w29208 & w42435) | (w28920 & w42435);
assign w49217 = w29157 & w29245;
assign w49218 = ~w28920 & w49989;
assign w49219 = ~w29559 & w29561;
assign w49220 = w29559 & w29564;
assign w49221 = ~w29559 & w29571;
assign w49222 = w29559 & w29574;
assign w49223 = ~w28920 & w49990;
assign w49224 = ~w28920 & w49991;
assign w49225 = ~w29781 & w2285;
assign w49226 = ~w28920 & w49992;
assign w49227 = ~w29864 & ~w1738;
assign w49228 = ~w29895 & w2006;
assign w49229 = ~w28920 & w49993;
assign w49230 = ~w29986 & w29988;
assign w49231 = w29986 & w29991;
assign w49232 = ~w29986 & w30015;
assign w49233 = w29986 & w30018;
assign w49234 = (~w30044 & w28920) | (~w30044 & w49994) | (w28920 & w49994);
assign w49235 = (w3 & ~w28855) | (w3 & w49995) | (~w28855 & w49995);
assign w49236 = ~w28920 & w49996;
assign w49237 = ~w30079 & w30082;
assign w49238 = w30079 & w30085;
assign w49239 = ~w28920 & w49997;
assign w49240 = ~w30158 & w5330;
assign w49241 = w30158 & ~w5330;
assign w49242 = ~w30160 & w4838;
assign w49243 = ~w29678 & w30184;
assign w49244 = w29678 & w30187;
assign w49245 = ~w29962 & w30236;
assign w49246 = w29963 & w30034;
assign w49247 = w29963 & ~w30032;
assign w49248 = w30972 & w7924;
assign w49249 = ~w31484 & w31486;
assign w49250 = w31540 & ~w31849;
assign w49251 = ~w31986 & w31988;
assign w49252 = ~a[8] & ~w34895;
assign w49253 = ~a[8] & w42874;
assign w49254 = w34617 & w35002;
assign w49255 = w34617 & ~w42883;
assign w49256 = ~w35872 & w400;
assign w49257 = w35872 & w400;
assign w49258 = ~w34897 & w42956;
assign w49259 = w33765 & w612;
assign w49260 = w34912 & ~w754;
assign w49261 = ~w35760 & ~w35745;
assign w49262 = w35994 & ~w36737;
assign w49263 = ~w36778 & w252;
assign w49264 = ~w36978 & ~w36985;
assign w49265 = w37004 & ~w37008;
assign w49266 = ~w37143 & ~w36572;
assign w49267 = ~w37143 & w46180;
assign w49268 = w36732 & ~w36572;
assign w49269 = w36732 & w46180;
assign w49270 = ~w37166 & ~w36572;
assign w49271 = ~w37166 & w46186;
assign w49272 = w37058 & ~w37614;
assign w49273 = w37058 & ~w37628;
assign w49274 = w4164 & w400;
assign w49275 = w4164 & w40160;
assign w49276 = w4170 & w400;
assign w49277 = w4170 & w40160;
assign w49278 = w4377 & ~w4351;
assign w49279 = w5743 & ~w5339;
assign w49280 = ~w7401 & w612;
assign w49281 = ~w7430 & ~w400;
assign w49282 = w6997 & ~w1541;
assign w49283 = ~w7640 & w7642;
assign w49284 = w7640 & w7644;
assign w49285 = w7675 & w7678;
assign w49286 = ~w7675 & w7680;
assign w49287 = w3646 & w3242;
assign w49288 = (w7814 & w43409) | (w7814 & ~w7314) | (w43409 & ~w7314);
assign w49289 = (w7814 & w43409) | (w7814 & w7139) | (w43409 & w7139);
assign w49290 = (w7837 & w46527) | (w7837 & ~w7314) | (w46527 & ~w7314);
assign w49291 = (w7837 & w46527) | (w7837 & w7139) | (w46527 & w7139);
assign w49292 = ~w7220 & ~w7843;
assign w49293 = w1320 & ~w7933;
assign w49294 = ~w11861 & w12147;
assign w49295 = ~w11861 & w12185;
assign w49296 = w11435 & ~w40955;
assign w49297 = w12354 & ~w11865;
assign w49298 = (w12626 & ~w12611) | (w12626 & w50451) | (~w12611 & w50451);
assign w49299 = (w1120 & w14458) | (w1120 & w50452) | (w14458 & w50452);
assign w49300 = ~w14458 & w50453;
assign w49301 = w15736 & w16515;
assign w49302 = w15736 & w16521;
assign w49303 = w22932 & w22939;
assign w49304 = w22932 & w22971;
assign w49305 = ~w23413 & ~w22705;
assign w49306 = ~w26076 & ~w252;
assign w49307 = w27949 & w27216;
assign w49308 = w30248 & ~w29963;
assign w49309 = w43779 & w34892;
assign w49310 = (w34892 & w43779) | (w34892 & ~w34996) | (w43779 & ~w34996);
assign w49311 = ~w35025 & ~a[9];
assign w49312 = ~w33855 & w35039;
assign w49313 = w33855 & w43780;
assign w49314 = w35193 & ~w20906;
assign w49315 = ~w35193 & w20906;
assign w49316 = ~w34897 & w43783;
assign w49317 = ~w34897 & w43797;
assign w49318 = ~w35640 & w43798;
assign w49319 = ~w34664 & w33850;
assign w49320 = ~w34664 & ~w33845;
assign w49321 = ~w34897 & w43804;
assign w49322 = ~w34897 & w43806;
assign w49323 = w4838 & ~w43381;
assign w49324 = w4430 & ~w43382;
assign w49325 = w4430 & ~w43383;
assign w49326 = ~w7277 & w7278;
assign w49327 = w7277 & w7399;
assign w49328 = ~w32966 & w32872;
assign w49329 = ~w34830 & ~w34821;
assign w49330 = ~w4342 & w4211;
assign w49331 = ~w5064 & ~w5133;
assign w49332 = w5597 & w493;
assign w49333 = w5622 & ~w493;
assign w49334 = w5622 & w44213;
assign w49335 = w5632 & w400;
assign w49336 = w5632 & w44216;
assign w49337 = w6262 & ~w6361;
assign w49338 = w6262 & w6413;
assign w49339 = ~w6262 & w6415;
assign w49340 = w6262 & w6436;
assign w49341 = ~w6262 & w6438;
assign w49342 = w6262 & ~w6694;
assign w49343 = w6262 & w6726;
assign w49344 = w6698 & ~w351;
assign w49345 = w7151 & w6642;
assign w49346 = w7151 & w44283;
assign w49347 = ~w7325 & w945;
assign w49348 = w2285 & ~w43475;
assign w49349 = w2285 & ~w43474;
assign w49350 = w15671 & w16482;
assign w49351 = ~w25454 & ~w25783;
assign w49352 = w25971 & ~w351;
assign w49353 = w945 & w32849;
assign w49354 = w32998 & w46978;
assign w49355 = w46979 | w33818;
assign w49356 = (w33818 & w46979) | (w33818 & ~w32998) | (w46979 & ~w32998);
assign w49357 = w46980 | ~w33815;
assign w49358 = (~w33815 & w46980) | (~w33815 & ~w32998) | (w46980 & ~w32998);
assign w49359 = w32998 & w46981;
assign w49360 = w32996 & w33900;
assign w49361 = ~w35652 & ~w35649;
assign w49362 = w46084 & w35776;
assign w49363 = ~w46084 & ~w35776;
assign w49364 = ~w46097 & w351;
assign w49365 = w35887 & ~w43777;
assign w49366 = w35887 & ~w34906;
assign w49367 = w46097 & ~w351;
assign w49368 = ~w24951 & ~w12666;
assign w49369 = ~w34282 & w8666;
assign w49370 = w34282 & ~w8666;
assign w49371 = ~w17366 & w17042;
assign w49372 = w34131 & ~w33935;
assign w49373 = w4682 & w51447;
assign w49374 = ~w5853 & w6254;
assign w49375 = ~w6814 & ~w1320;
assign w49376 = ~w6609 & ~w6834;
assign w49377 = ~w6609 & w6854;
assign w49378 = w6609 & w6857;
assign w49379 = ~w6609 & w6880;
assign w49380 = ~w6609 & a[75];
assign w49381 = w6609 & ~a[75];
assign w49382 = ~w6609 & ~w5330;
assign w49383 = ~w6609 & w6390;
assign w49384 = w6609 & ~w6390;
assign w49385 = w6609 & ~w6432;
assign w49386 = w6754 & w6318;
assign w49387 = w6754 & w40434;
assign w49388 = ~w6609 & w7231;
assign w49389 = w7268 & w1320;
assign w49390 = ~w7268 & ~w7276;
assign w49391 = w7268 & ~w7846;
assign w49392 = w8596 & w8856;
assign w49393 = ~w13350 & w50454;
assign w49394 = ~w13350 & w50455;
assign w49395 = (w4838 & w13350) | (w4838 & w50456) | (w13350 & w50456);
assign w49396 = (~w4056 & w13350) | (~w4056 & w50457) | (w13350 & w50457);
assign w49397 = (w3242 & w13350) | (w3242 & w50458) | (w13350 & w50458);
assign w49398 = (~w4430 & w13350) | (~w4430 & w50459) | (w13350 & w50459);
assign w49399 = w13382 & w4056;
assign w49400 = ~w13350 & w50460;
assign w49401 = (w13762 & w13350) | (w13762 & w50461) | (w13350 & w50461);
assign w49402 = (~w13759 & w13350) | (~w13759 & w50462) | (w13350 & w50462);
assign w49403 = ~w13350 & w50463;
assign w49404 = ~w13350 & w50464;
assign w49405 = (w13796 & w13350) | (w13796 & w50465) | (w13350 & w50465);
assign w49406 = ~w13350 & w50466;
assign w49407 = (w13802 & w13350) | (w13802 & w50467) | (w13350 & w50467);
assign w49408 = ~w13350 & w50468;
assign w49409 = (w13813 & w13350) | (w13813 & w50469) | (w13350 & w50469);
assign w49410 = ~w13350 & w50470;
assign w49411 = (w13891 & w13350) | (w13891 & w50471) | (w13350 & w50471);
assign w49412 = ~w13350 & w50472;
assign w49413 = ~w13350 & w50473;
assign w49414 = (~w1541 & w13350) | (~w1541 & w50474) | (w13350 & w50474);
assign w49415 = (~w1738 & w13350) | (~w1738 & w50475) | (w13350 & w50475);
assign w49416 = ~w13350 & w50476;
assign w49417 = (w6769 & w41194) | (w6769 & w14037) | (w41194 & w14037);
assign w49418 = (w6769 & w41194) | (w6769 & ~w13935) | (w41194 & ~w13935);
assign w49419 = w16756 & w16820;
assign w49420 = ~w22878 & ~w22880;
assign w49421 = w22878 & w22880;
assign w49422 = (w27785 & w27873) | (w27785 & w49998) | (w27873 & w49998);
assign w49423 = w32719 & ~w46977;
assign w49424 = ~w80 & w33766;
assign w49425 = w80 & ~w33766;
assign w49426 = w34929 & ~w26880;
assign w49427 = ~w33854 & w35029;
assign w49428 = w34895 & w35060;
assign w49429 = ~w35095 & w29158;
assign w49430 = ~w35158 & ~w35296;
assign w49431 = w34878 & ~w43784;
assign w49432 = ~w7924 & w35447;
assign w49433 = w7924 & w35449;
assign w49434 = w34279 & w34239;
assign w49435 = ~w33855 & ~w34216;
assign w49436 = w33855 & w34216;
assign w49437 = w35297 & w36014;
assign w49438 = w7010 & ~w1120;
assign w49439 = ~w35297 & w35022;
assign w49440 = w35297 & ~w36016;
assign w49441 = w35297 & w36038;
assign w49442 = w35297 & ~w36057;
assign w49443 = ~w35297 & w36065;
assign w49444 = w35297 & w36075;
assign w49445 = w35297 & w36103;
assign w49446 = w35297 & w36123;
assign w49447 = ~w35297 & w28077;
assign w49448 = w35297 & w36130;
assign w49449 = w35297 & w36145;
assign w49450 = ~w35297 & w25851;
assign w49451 = w35297 & w36152;
assign w49452 = ~w35297 & w35257;
assign w49453 = ~w35297 & ~w35120;
assign w49454 = w35297 & w36190;
assign w49455 = w35297 & ~w35463;
assign w49456 = ~w35297 & ~w2558;
assign w49457 = w35297 & w36750;
assign w49458 = ~w35297 & ~w36754;
assign w49459 = ~w35297 & w36754;
assign w49460 = w35297 & ~w35946;
assign w49461 = ~w7202 & ~w7115;
assign w49462 = w7202 & ~w612;
assign w49463 = w7202 & w7114;
assign w49464 = w7202 & ~w2558;
assign w49465 = w7202 & w2285;
assign w49466 = w7202 & w7555;
assign w49467 = w7202 & w7606;
assign w49468 = w7202 & w7617;
assign w49469 = w7202 & w7630;
assign w49470 = w7202 & w7652;
assign w49471 = w7202 & ~w7660;
assign w49472 = w7202 & ~w7718;
assign w49473 = w7202 & w7728;
assign w49474 = w7202 & w7290;
assign w49475 = ~w7268 & w7745;
assign w49476 = w7268 & w7747;
assign w49477 = w7284 & ~w7301;
assign w49478 = ~w5559 & w754;
assign w49479 = w5839 & w57;
assign w49480 = ~w4627 & ~w4625;
assign w49481 = ~w4626 & w49480;
assign w49482 = w4627 & w4625;
assign w49483 = (w4627 & w4626) | (w4627 & w49482) | (w4626 & w49482);
assign w49484 = w4688 & w40245;
assign w49485 = w5170 & ~w4703;
assign w49486 = w5180 & w252;
assign w49487 = ~w5180 & ~w252;
assign w49488 = w40257 & w5202;
assign w49489 = (w5202 & w40257) | (w5202 & w5168) | (w40257 & w5168);
assign w49490 = ~w5168 & w40258;
assign w49491 = w40259 & w5208;
assign w49492 = (w5208 & w40259) | (w5208 & w5168) | (w40259 & w5168);
assign w49493 = ~w5168 & w40260;
assign w49494 = w5217 & ~w5168;
assign w49495 = ~w5692 & w5267;
assign w49496 = w5757 & ~w1541;
assign w49497 = w5718 & ~w5986;
assign w49498 = w5718 & ~w4838;
assign w49499 = w6152 & ~w6157;
assign w49500 = ~w5934 & ~w5963;
assign w49501 = ~w40390 & ~w6268;
assign w49502 = ~w6265 & w5962;
assign w49503 = ~w5917 & w6086;
assign w49504 = w5854 & w2285;
assign w49505 = w5854 & w2558;
assign w49506 = w5854 & ~w1738;
assign w49507 = w5854 & ~w2896;
assign w49508 = w5854 & ~w351;
assign w49509 = ~w6262 & w6648;
assign w49510 = ~w6262 & ~w351;
assign w49511 = w6695 & ~w400;
assign w49512 = w6752 & w612;
assign w49513 = ~w6309 & ~w6764;
assign w49514 = ~w6307 & w6319;
assign w49515 = w6307 & w6264;
assign w49516 = w6307 & w6863;
assign w49517 = w6307 & w2896;
assign w49518 = ~w6543 & w7002;
assign w49519 = w6543 & ~w7002;
assign w49520 = w7026 & w6318;
assign w49521 = w7026 & w40434;
assign w49522 = w6799 & w6318;
assign w49523 = w6799 & w40434;
assign w49524 = ~w7083 & w1320;
assign w49525 = ~w6698 & w6318;
assign w49526 = ~w6698 & w40434;
assign w49527 = ~w6710 & w6318;
assign w49528 = ~w6710 & w40434;
assign w49529 = ~w6796 & w6821;
assign w49530 = ~w6796 & w44273;
assign w49531 = (~w945 & w44309) | (~w945 & ~w7314) | (w44309 & ~w7314);
assign w49532 = (~w945 & w44309) | (~w945 & w7139) | (w44309 & w7139);
assign w49533 = (~w1120 & w44310) | (~w1120 & ~w7314) | (w44310 & ~w7314);
assign w49534 = (~w1120 & w44310) | (~w1120 & w7139) | (w44310 & w7139);
assign w49535 = ~w7268 & ~w612;
assign w49536 = ~w7268 & w7114;
assign w49537 = w754 & ~w44318;
assign w49538 = w754 & ~w44319;
assign w49539 = ~w40489 & w7454;
assign w49540 = w40489 & ~w7454;
assign w49541 = ~w7268 & ~w6997;
assign w49542 = ~w6985 & w7063;
assign w49543 = ~w7268 & ~w2558;
assign w49544 = ~w7268 & w2285;
assign w49545 = ~w7030 & w7039;
assign w49546 = ~w7520 & w1738;
assign w49547 = ~w7466 & w1541;
assign w49548 = ~w7268 & w7555;
assign w49549 = w7268 & ~w7552;
assign w49550 = a[71] & w6318;
assign w49551 = a[71] & w40434;
assign w49552 = w7268 & ~w7575;
assign w49553 = ~w7568 & w6318;
assign w49554 = ~w7568 & w40434;
assign w49555 = ~w7268 & ~w7584;
assign w49556 = w7268 & w7592;
assign w49557 = ~w7268 & w7595;
assign w49558 = w7268 & w40495;
assign w49559 = w40496 & w7606;
assign w49560 = (w7606 & w40496) | (w7606 & ~w7268) | (w40496 & ~w7268);
assign w49561 = w7268 & w40497;
assign w49562 = w40498 & w7617;
assign w49563 = (w7617 & w40498) | (w7617 & ~w7268) | (w40498 & ~w7268);
assign w49564 = ~w4838 & ~w7637;
assign w49565 = ~w4838 & w40501;
assign w49566 = w4838 & w7637;
assign w49567 = w4838 & ~w40501;
assign w49568 = w6895 & ~w6903;
assign w49569 = w6837 & w7685;
assign w49570 = ~w7268 & ~w7718;
assign w49571 = ~w7305 & ~w7744;
assign w49572 = w7305 & w7744;
assign w49573 = w7268 & ~w351;
assign w49574 = w40525 | ~w7194;
assign w49575 = (~w7194 & w40525) | (~w7194 & w7784) | (w40525 & w7784);
assign w49576 = w7268 & ~w7195;
assign w49577 = w7178 & w50250;
assign w49578 = (w7784 & w44337) | (w7784 & w44338) | (w44337 & w44338);
assign w49579 = ~w7268 & w7290;
assign w49580 = w7268 & ~w7863;
assign w49581 = w7268 & w7863;
assign w49582 = ~w7879 & w47211;
assign w49583 = ~w7879 & w47210;
assign w49584 = w7893 & ~w7898;
assign w49585 = w7848 & ~w3;
assign w49586 = ~w7949 & w7959;
assign w49587 = ~w7451 & w8040;
assign w49588 = w7783 & w8057;
assign w49589 = w252 & ~w44344;
assign w49590 = w252 & w47215;
assign w49591 = ~w8044 & w400;
assign w49592 = w8070 & w8071;
assign w49593 = w8072 & ~w7831;
assign w49594 = w8117 & w3;
assign w49595 = w8123 & ~w8120;
assign w49596 = w8123 & ~w44359;
assign w49597 = w8130 & ~w8127;
assign w49598 = w8130 & ~w44360;
assign w49599 = ~w8133 & ~w8134;
assign w49600 = ~w8133 & ~w44361;
assign w49601 = ~w7854 & ~w8127;
assign w49602 = ~w7854 & ~w44360;
assign w49603 = w8177 & ~w42;
assign w49604 = ~w8118 & ~w3;
assign w49605 = w8291 & w8287;
assign w49606 = w8291 & w40604;
assign w49607 = w6264 & ~w8294;
assign w49608 = w7759 & w8527;
assign w49609 = ~w8555 & w8557;
assign w49610 = ~w40649 & w8018;
assign w49611 = w8157 & ~w8585;
assign w49612 = ~w8189 & w8511;
assign w49613 = w8672 & ~w1541;
assign w49614 = ~w8189 & w8719;
assign w49615 = w8728 & w2285;
assign w49616 = ~w8720 & ~w2006;
assign w49617 = ~w8672 & w1541;
assign w49618 = ~w8189 & ~w8331;
assign w49619 = w8189 & ~w8771;
assign w49620 = ~w8101 & w5745;
assign w49621 = w8776 & ~w8775;
assign w49622 = ~w8189 & w8315;
assign w49623 = ~w8403 & ~w8316;
assign w49624 = ~w8101 & w8889;
assign w49625 = ~w8189 & w8901;
assign w49626 = w8189 & w8903;
assign w49627 = ~w8189 & w8900;
assign w49628 = w8189 & ~w8914;
assign w49629 = w8189 & ~w8219;
assign w49630 = w8189 & w8927;
assign w49631 = w8189 & w8941;
assign w49632 = ~w9016 & w8099;
assign w49633 = ~w9016 & w44414;
assign w49634 = ~w44418 & w8033;
assign w49635 = ~w8189 & w80;
assign w49636 = w9119 & w9121;
assign w49637 = ~w9119 & w9123;
assign w49638 = w13894 & ~w13875;
assign w49639 = w14043 & w14056;
assign w49640 = ~w14310 & ~w14311;
assign w49641 = (w14328 & w14027) | (w14328 & w50477) | (w14027 & w50477);
assign w49642 = ~w14333 & ~w14331;
assign w49643 = (w13681 & w14027) | (w13681 & w50478) | (w14027 & w50478);
assign w49644 = ~w14027 & w50479;
assign w49645 = w14334 & w50480;
assign w49646 = w14375 & ~w14389;
assign w49647 = (w14402 & w14027) | (w14402 & w50481) | (w14027 & w50481);
assign w49648 = ~w14027 & w50482;
assign w49649 = w41221 & w14416;
assign w49650 = (w14416 & w41221) | (w14416 & ~w14375) | (w41221 & ~w14375);
assign w49651 = (~w13709 & w14027) | (~w13709 & w50483) | (w14027 & w50483);
assign w49652 = ~w14027 & w50484;
assign w49653 = ~w14444 & ~w13954;
assign w49654 = (~w13982 & w14027) | (~w13982 & w50485) | (w14027 & w50485);
assign w49655 = ~w14484 & w14488;
assign w49656 = (~w14491 & w14486) | (~w14491 & w50486) | (w14486 & w50486);
assign w49657 = (~w14491 & w41231) | (~w14491 & w14484) | (w41231 & w14484);
assign w49658 = (~w13880 & w14027) | (~w13880 & w50487) | (w14027 & w50487);
assign w49659 = ~w13584 & w14620;
assign w49660 = ~w14630 & w50488;
assign w49661 = ~w14634 & w252;
assign w49662 = w14043 & ~w14709;
assign w49663 = ~w15174 & w15172;
assign w49664 = ~w15174 & w41320;
assign w49665 = w41354 & w11138;
assign w49666 = w26044 & ~w25947;
assign w49667 = (~w28076 & w50173) | (~w28076 & w50174) | (w50173 & w50174);
assign w49668 = (w28076 & w50175) | (w28076 & w50176) | (w50175 & w50176);
assign w49669 = ~w28589 & w28599;
assign w49670 = w28589 & w28593;
assign w49671 = ~w27861 & ~w28608;
assign w49672 = w28562 & w28624;
assign w49673 = w28562 & ~w28635;
assign w49674 = ~w28562 & ~w27859;
assign w49675 = w28619 & ~w7315;
assign w49676 = ~w28491 & w28671;
assign w49677 = w28491 & w28673;
assign w49678 = ~w27949 & w27999;
assign w49679 = ~w28695 & w28696;
assign w49680 = ~w28077 & ~w28771;
assign w49681 = ~w28800 & ~w26992;
assign w49682 = ~w27949 & ~w754;
assign w49683 = w28820 & ~w493;
assign w49684 = ~w28755 & w28848;
assign w49685 = w28755 & w28850;
assign w49686 = w28865 & ~w3;
assign w49687 = ~w28019 & ~w28075;
assign w49688 = ~w28894 & ~w28893;
assign w49689 = w28888 & w28904;
assign w49690 = w28788 & ~w28793;
assign w49691 = ~w28967 & w1541;
assign w49692 = w28967 & ~w1541;
assign w49693 = w27847 & w27900;
assign w49694 = ~w27949 & ~w29023;
assign w49695 = ~w29008 & ~w29006;
assign w49696 = ~w29230 & ~w29225;
assign w49697 = ~w29234 & ~w28176;
assign w49698 = w28273 & w28504;
assign w49699 = w28273 & ~w16559;
assign w49700 = ~w28273 & w16559;
assign w49701 = ~w32704 & ~w47957;
assign w49702 = ~w32704 & ~w47958;
assign w49703 = ~w42 & w33783;
assign w49704 = w32988 & ~w32983;
assign w49705 = w33803 & ~w33787;
assign w49706 = ~w32998 & w33837;
assign w49707 = ~w33792 & w32808;
assign w49708 = ~w33840 & w252;
assign w49709 = w33773 & w33786;
assign w49710 = w33978 & ~w25851;
assign w49711 = w32998 & w493;
assign w49712 = w34594 & w34592;
assign w49713 = ~w34594 & ~w34592;
assign w49714 = w32998 & w400;
assign w49715 = ~w34600 & ~w34603;
assign w49716 = w34600 & w34603;
assign w49717 = ~w34611 & ~w493;
assign w49718 = w34622 & w34624;
assign w49719 = ~w34622 & w34626;
assign w49720 = w34611 & w493;
assign w49721 = w34594 & w34630;
assign w49722 = ~w34594 & w34632;
assign w49723 = w34655 & ~w34618;
assign w49724 = ~w34869 & w34664;
assign w49725 = ~w34885 & w34887;
assign w49726 = w33765 & w33784;
assign w49727 = w34590 & ~w34871;
assign w49728 = ~w34916 & w34918;
assign w49729 = w42874 & ~w34895;
assign w49730 = (~w34895 & w42874) | (~w34895 & w34916) | (w42874 & w34916);
assign w49731 = ~w33962 & ~w33954;
assign w49732 = ~w33979 & w34898;
assign w49733 = ~w33979 & ~w47999;
assign w49734 = w33979 & ~w34898;
assign w49735 = w33979 & w47999;
assign w49736 = ~w34916 & ~w34871;
assign w49737 = w42883 & ~w35002;
assign w49738 = (~w35002 & w42883) | (~w35002 & w34916) | (w42883 & w34916);
assign w49739 = ~w34916 & w48007;
assign w49740 = ~w34916 & w42886;
assign w49741 = w48012 | w32698;
assign w49742 = (w32698 & w48012) | (w32698 & w35040) | (w48012 & w35040);
assign w49743 = ~w35040 & w48013;
assign w49744 = ~w28077 & ~w42887;
assign w49745 = ~w28077 & ~w34898;
assign w49746 = ~w35103 & w35110;
assign w49747 = ~w23843 & ~w33855;
assign w49748 = ~w23843 & w34898;
assign w49749 = w35122 & w26445;
assign w49750 = w34220 & ~w35145;
assign w49751 = ~w35153 & ~w33855;
assign w49752 = ~w35153 & w34898;
assign w49753 = ~w34040 & w34102;
assign w49754 = ~w34162 & w34898;
assign w49755 = w35211 & ~w18183;
assign w49756 = ~w35155 & ~w14766;
assign w49757 = w34574 & ~w48038;
assign w49758 = w34574 & ~w48039;
assign w49759 = ~w3646 & w33855;
assign w49760 = ~w3646 & ~w34898;
assign w49761 = w34224 & ~w33855;
assign w49762 = w34224 & w34898;
assign w49763 = w35562 & w11870;
assign w49764 = ~w35596 & ~w35599;
assign w49765 = ~w35609 & ~w35408;
assign w49766 = ~w35633 & ~w35409;
assign w49767 = ~w35642 & w4838;
assign w49768 = ~w34836 & ~w35683;
assign w49769 = ~w34836 & ~w46068;
assign w49770 = w35730 & w34850;
assign w49771 = w35730 & w46076;
assign w49772 = w34838 & ~w35683;
assign w49773 = w34838 & ~w46068;
assign w49774 = ~w80 & w33820;
assign w49775 = ~w80 & w46093;
assign w49776 = ~w35845 & w80;
assign w49777 = w35845 & ~w80;
assign w49778 = w35851 & w35853;
assign w49779 = ~w34885 & w35869;
assign w49780 = w34900 & w46098;
assign w49781 = w46100 & ~w351;
assign w49782 = (~w351 & w46100) | (~w351 & ~w34900) | (w46100 & ~w34900);
assign w49783 = (~w400 & w42962) | (~w400 & w35887) | (w42962 & w35887);
assign w49784 = (~w400 & w42962) | (~w400 & w46099) | (w42962 & w46099);
assign w49785 = w42967 & w35936;
assign w49786 = (w35936 & w42967) | (w35936 & w35633) | (w42967 & w35633);
assign w49787 = w36041 & w36038;
assign w49788 = w36041 & w42980;
assign w49789 = w36072 & w36038;
assign w49790 = w36072 & w42980;
assign w49791 = w36078 & w36075;
assign w49792 = w36078 & w42983;
assign w49793 = ~w35070 & w36103;
assign w49794 = ~w35070 & w42985;
assign w49795 = ~w35021 & w36075;
assign w49796 = ~w35021 & w42983;
assign w49797 = ~w34934 & w36123;
assign w49798 = ~w34934 & w42986;
assign w49799 = w36138 & w36123;
assign w49800 = w36138 & w42986;
assign w49801 = ~w36141 & ~w36127;
assign w49802 = ~w34952 & w36145;
assign w49803 = ~w34952 & w42989;
assign w49804 = w36150 & ~w36149;
assign w49805 = w36194 & w36190;
assign w49806 = w36194 & w42996;
assign w49807 = w36199 & w36190;
assign w49808 = w36199 & w42996;
assign w49809 = w36202 & ~w36173;
assign w49810 = w36990 & ~w35946;
assign w49811 = w36990 & w43104;
assign w49812 = w5894 & w5875;
assign w49813 = w5894 & w40316;
assign w49814 = ~w4838 & ~w5981;
assign w49815 = ~w4838 & w40335;
assign w49816 = w6043 & w6039;
assign w49817 = w6043 & w40345;
assign w49818 = ~w6120 & ~w80;
assign w49819 = ~w6619 & ~w57;
assign w49820 = w6619 & w57;
assign w49821 = ~w6727 & ~w6212;
assign w49822 = ~w6727 & w40428;
assign w49823 = w6727 & w6212;
assign w49824 = w6727 & ~w40428;
assign w49825 = w7401 & ~w612;
assign w49826 = ~w41234 & ~w612;
assign w49827 = w14634 & ~w252;
assign w49828 = w26073 & ~w1120;
assign w49829 = ~w26073 & w27288;
assign w49830 = w27776 & ~w27752;
assign w49831 = w28077 & w252;
assign w49832 = w33855 & ~w8666;
assign w49833 = w33855 & ~w42910;
assign w49834 = ~w27949 & w28080;
assign w49835 = w46782 & w27270;
assign w49836 = (w27270 & w46782) | (w27270 & w27949) | (w46782 & w27949);
assign w49837 = w27949 & w14039;
assign w49838 = w28444 & ~w27482;
assign w49839 = ~w27949 & ~w28512;
assign w49840 = w27949 & w4838;
assign w49841 = w27949 & ~w5330;
assign w49842 = ~w27949 & w7315;
assign w49843 = w27949 & ~w6769;
assign w49844 = w27949 & w252;
assign w49845 = ~w27949 & ~w80;
assign w49846 = ~w27949 & w28001;
assign w49847 = w27949 & w27196;
assign w49848 = w27949 & w3646;
assign w49849 = w5974 & w6237;
assign w49850 = ~w8179 & ~w8890;
assign w49851 = w13713 & ~w14037;
assign w49852 = w13857 & w50489;
assign w49853 = w13391 & ~w14037;
assign w49854 = w13857 & w50490;
assign w49855 = w13469 & ~w14037;
assign w49856 = w13857 & w50491;
assign w49857 = ~w14167 & ~w14037;
assign w49858 = w13857 & w50492;
assign w49859 = w6264 & w13391;
assign w49860 = w6264 & w44756;
assign w49861 = w14173 & ~w14037;
assign w49862 = w13857 & w50493;
assign w49863 = w13516 & ~w14037;
assign w49864 = w13857 & w50494;
assign w49865 = w5745 & ~w14167;
assign w49866 = w5745 & w44759;
assign w49867 = ~w13579 & ~w14037;
assign w49868 = w13857 & w50495;
assign w49869 = w14237 & ~w14037;
assign w49870 = w13857 & w50496;
assign w49871 = ~w14259 & ~w14037;
assign w49872 = w13857 & w50497;
assign w49873 = ~w3242 & ~w14259;
assign w49874 = ~w3242 & w44774;
assign w49875 = w13612 & ~w14037;
assign w49876 = w13857 & w50498;
assign w49877 = w3646 & w13612;
assign w49878 = w3646 & w44782;
assign w49879 = ~w13500 & ~w14037;
assign w49880 = w13857 & w50499;
assign w49881 = w4056 & ~w13500;
assign w49882 = w4056 & w44784;
assign w49883 = w13979 & ~w14037;
assign w49884 = w13857 & w50500;
assign w49885 = w1738 & w13979;
assign w49886 = w1738 & w44813;
assign w49887 = ~w13544 & ~w14037;
assign w49888 = w13857 & w50501;
assign w49889 = w493 & ~w14037;
assign w49890 = w13857 & w50502;
assign w49891 = w14668 & w493;
assign w49892 = w14668 & w44827;
assign w49893 = w14674 & w493;
assign w49894 = w14674 & w44827;
assign w49895 = ~w612 & ~w14037;
assign w49896 = w13857 & w50503;
assign w49897 = w14682 & ~w612;
assign w49898 = w14682 & w44832;
assign w49899 = w14700 & ~w612;
assign w49900 = w14700 & w44832;
assign w49901 = ~w3 & ~w14037;
assign w49902 = w13857 & w50504;
assign w49903 = ~w14738 & ~w3;
assign w49904 = ~w14738 & w44837;
assign w49905 = w9781 & ~w26089;
assign w49906 = w25844 & w24929;
assign w49907 = w26181 & ~w25326;
assign w49908 = w25844 & w25020;
assign w49909 = ~w25837 & ~w26206;
assign w49910 = ~w25837 & w26217;
assign w49911 = ~w7315 & w25020;
assign w49912 = ~w7315 & w45528;
assign w49913 = w25844 & w6264;
assign w49914 = ~w25837 & w26362;
assign w49915 = ~w26524 & w26527;
assign w49916 = w26524 & w26529;
assign w49917 = ~w26536 & w26542;
assign w49918 = w26536 & w26544;
assign w49919 = w25844 & w25292;
assign w49920 = ~w26536 & ~w26541;
assign w49921 = w25844 & ~w1738;
assign w49922 = ~w25844 & ~w25426;
assign w49923 = ~w25844 & ~w25434;
assign w49924 = w25844 & w2896;
assign w49925 = ~w25837 & ~w25621;
assign w49926 = ~w26760 & ~w26958;
assign w49927 = ~w26706 & w27180;
assign w49928 = w26706 & ~w27180;
assign w49929 = w26557 & w25945;
assign w49930 = w26557 & ~w45513;
assign w49931 = w27659 & w8666;
assign w49932 = ~w26154 & ~w9195;
assign w49933 = w26229 & ~w7315;
assign w49934 = ~w27909 & w25899;
assign w49935 = ~w27909 & w25898;
assign w49936 = ~w26021 & ~w25945;
assign w49937 = ~w26021 & w45513;
assign w49938 = w80 & w28020;
assign w49939 = w28113 & w27256;
assign w49940 = w28769 & w28701;
assign w49941 = ~w35262 & ~w35311;
assign w49942 = ~w34866 & ~w43777;
assign w49943 = ~w34866 & ~w34906;
assign w49944 = ~w14766 & w28412;
assign w49945 = ~w44408 & ~w8891;
assign w49946 = w9075 & ~w9028;
assign w49947 = ~w25079 & ~w25789;
assign w49948 = ~w17380 & w16559;
assign w49949 = ~w17380 & ~w45578;
assign w49950 = w42275 & ~w26826;
assign w49951 = w42284 & ~w26826;
assign w49952 = w27380 & ~w21801;
assign w49953 = ~w27874 & w28509;
assign w49954 = ~w27874 & w27779;
assign w49955 = ~w27880 & w27900;
assign w49956 = w15681 & w42895;
assign w49957 = w15681 & w34898;
assign w49958 = ~w15681 & ~w42895;
assign w49959 = ~w15681 & ~w34898;
assign w49960 = w35410 & w42905;
assign w49961 = w35410 & w34898;
assign w49962 = ~w35410 & ~w42905;
assign w49963 = ~w35410 & ~w34898;
assign w49964 = w7086 & w7278;
assign w49965 = w27949 & w27616;
assign w49966 = ~w27949 & ~w27616;
assign w49967 = ~w6767 & ~w6605;
assign w49968 = ~w945 & w26827;
assign w49969 = ~w945 & w48442;
assign w49970 = w27685 & w9781;
assign w49971 = w26706 & w25899;
assign w49972 = w26706 & w25898;
assign w49973 = ~w27638 & w28508;
assign w49974 = ~w27638 & ~w27880;
assign w49975 = w48273 & w7278;
assign w49976 = ~w27167 & w3242;
assign w49977 = ~w27847 & w27880;
assign w49978 = ~w27780 & w27880;
assign w49979 = ~w43624 & ~w22767;
assign w49980 = w43624 & w22767;
assign w49981 = w27585 & w27256;
assign w49982 = w27401 & w27256;
assign w49983 = ~w43636 & w28516;
assign w49984 = w43636 & w28519;
assign w49985 = ~w43636 & w28534;
assign w49986 = w43636 & w28537;
assign w49987 = ~w28854 & w28884;
assign w49988 = ~w28930 & w28232;
assign w49989 = ~w28930 & ~w9195;
assign w49990 = ~w28930 & w4430;
assign w49991 = ~w28930 & w29061;
assign w49992 = ~w28930 & ~w29037;
assign w49993 = ~w28930 & ~w493;
assign w49994 = w28930 & ~w30044;
assign w49995 = ~w28854 & w3;
assign w49996 = ~w28930 & w57;
assign w49997 = ~w28930 & w30157;
assign w49998 = w27723 & w27785;
assign w49999 = w7001 & w6318;
assign w50000 = w7001 & w40434;
assign w50001 = w7007 & ~w1541;
assign w50002 = ~w8189 & w400;
assign w50003 = w9035 & w9038;
assign w50004 = ~w9035 & w9040;
assign w50005 = w9035 & w9146;
assign w50006 = ~w9035 & w9148;
assign w50007 = w24857 & ~w49102;
assign w50008 = w24857 & ~w49103;
assign w50009 = w24879 & ~w42;
assign w50010 = ~w25826 & ~w23863;
assign w50011 = ~w25826 & w42072;
assign w50012 = ~w25831 & w50251;
assign w50013 = ~w25771 & ~w25816;
assign w50014 = ~w25846 & ~w25845;
assign w50015 = w26054 & w26053;
assign w50016 = w26054 & ~w45508;
assign w50017 = ~w26091 & w26095;
assign w50018 = ~w26091 & ~w26094;
assign w50019 = ~w11870 & ~w24966;
assign w50020 = ~w11870 & w49118;
assign w50021 = w25837 & ~w13384;
assign w50022 = w25844 & ~w13384;
assign w50023 = ~w26196 & ~w25062;
assign w50024 = ~w26198 & ~w26199;
assign w50025 = w25837 & ~w26211;
assign w50026 = w25844 & ~w26211;
assign w50027 = w25837 & w25024;
assign w50028 = w25844 & w25024;
assign w50029 = ~w26256 & ~w26255;
assign w50030 = ~w26204 & w26265;
assign w50031 = ~w47716 & w26307;
assign w50032 = w47716 & ~w26307;
assign w50033 = w25850 & w25793;
assign w50034 = ~w26311 & w5330;
assign w50035 = ~w26322 & w26321;
assign w50036 = ~w26324 & w26329;
assign w50037 = w25850 & w25588;
assign w50038 = ~w26593 & ~w26688;
assign w50039 = ~w25844 & ~w25363;
assign w50040 = w25850 & w1541;
assign w50041 = ~w26738 & w26740;
assign w50042 = w26738 & w26742;
assign w50043 = ~w26054 & ~w26053;
assign w50044 = ~w26054 & w45508;
assign w50045 = w25850 & w1120;
assign w50046 = w26752 & w26756;
assign w50047 = ~w26752 & w26758;
assign w50048 = w25966 & w25987;
assign w50049 = w26888 & ~w400;
assign w50050 = w26920 & ~w26907;
assign w50051 = w26745 & ~w42251;
assign w50052 = w26745 & ~w26951;
assign w50053 = ~w26953 & w26956;
assign w50054 = w26877 & ~w26980;
assign w50055 = ~w26953 & w26955;
assign w50056 = w26952 & ~w26860;
assign w50057 = ~w27018 & w27022;
assign w50058 = w27018 & w27024;
assign w50059 = w26783 & ~w26855;
assign w50060 = w26880 & w27080;
assign w50061 = ~w26880 & w27082;
assign w50062 = ~w26719 & w26394;
assign w50063 = w26423 & ~w3646;
assign w50064 = ~w27160 & ~w26356;
assign w50065 = w26880 & w26782;
assign w50066 = ~w26880 & ~w26782;
assign w50067 = ~w26851 & ~w27021;
assign w50068 = w26880 & ~w1320;
assign w50069 = ~w26979 & w945;
assign w50070 = w26877 & w27279;
assign w50071 = w42275 & ~w24874;
assign w50072 = ~w26074 & w27301;
assign w50073 = w26877 & ~w27315;
assign w50074 = w26877 & w27322;
assign w50075 = w26521 & ~w27364;
assign w50076 = ~w18183 & w27389;
assign w50077 = ~w18183 & w42286;
assign w50078 = w26877 & ~w27392;
assign w50079 = ~w26073 & ~w26615;
assign w50080 = w26073 & w26615;
assign w50081 = w42284 & w27421;
assign w50082 = w26877 & ~w27403;
assign w50083 = ~w26073 & ~w27475;
assign w50084 = ~w27469 & w16559;
assign w50085 = w26877 & ~w27672;
assign w50086 = ~w27702 & w26114;
assign w50087 = ~w27702 & w45643;
assign w50088 = w27716 & ~w26292;
assign w50089 = w27716 & ~w45646;
assign w50090 = ~w27749 & ~w27748;
assign w50091 = ~w27749 & ~w42319;
assign w50092 = ~w27753 & ~w27754;
assign w50093 = ~w27753 & ~w42320;
assign w50094 = w27793 & ~w49145;
assign w50095 = w27793 & ~w49146;
assign w50096 = w25936 & ~w45663;
assign w50097 = w25936 & ~w45662;
assign w50098 = w27933 & ~w27935;
assign w50099 = ~w27945 & w42;
assign w50100 = ~w27963 & ~w27964;
assign w50101 = w27963 & w27964;
assign w50102 = w27963 & w28012;
assign w50103 = ~w27963 & w28014;
assign w50104 = w27968 & w28017;
assign w50105 = ~w27253 & w28046;
assign w50106 = ~w28050 & w28090;
assign w50107 = w28050 & w28160;
assign w50108 = w27291 & w23843;
assign w50109 = ~w27291 & ~w23843;
assign w50110 = w28050 & w28195;
assign w50111 = ~w27458 & ~w27461;
assign w50112 = ~w28242 & w17380;
assign w50113 = w28242 & ~w17380;
assign w50114 = ~w28302 & w28301;
assign w50115 = w28307 & ~w28075;
assign w50116 = w28325 & ~w11138;
assign w50117 = ~w11138 & w28370;
assign w50118 = ~w28371 & w10419;
assign w50119 = ~w28352 & w12666;
assign w50120 = w28394 & w28401;
assign w50121 = ~w28402 & ~w13384;
assign w50122 = w28402 & w13384;
assign w50123 = ~w27485 & w28427;
assign w50124 = w28407 & w28498;
assign w50125 = ~w28441 & w28426;
assign w50126 = ~w28067 & ~w27260;
assign w50127 = w28562 & w27862;
assign w50128 = w28576 & ~w6769;
assign w50129 = w28585 & ~w5745;
assign w50130 = ~w28585 & w5745;
assign w50131 = ~w28576 & w6769;
assign w50132 = w28677 & w28658;
assign w50133 = ~w27255 & ~w28717;
assign w50134 = w28825 & w28820;
assign w50135 = ~w29025 & ~w29024;
assign w50136 = ~w30259 & w30260;
assign w50137 = w35269 & ~w35237;
assign w50138 = w35545 & w35568;
assign w50139 = w35570 & w35609;
assign w50140 = w7279 & w7011;
assign w50141 = ~w42270 & ~w27184;
assign w50142 = ~w28144 & w43622;
assign w50143 = ~w28419 & w14039;
assign w50144 = w43635 & ~w28512;
assign w50145 = (~w28512 & w43635) | (~w28512 & w28038) | (w43635 & w28038);
assign w50146 = ~w28038 & w43648;
assign w50147 = w43662 & w28001;
assign w50148 = (w28001 & w43662) | (w28001 & w28038) | (w43662 & w28038);
assign w50149 = w42407 & w28877;
assign w50150 = ~w28037 & ~w27874;
assign w50151 = ~w28037 & w27640;
assign w50152 = w945 & ~w44301;
assign w50153 = w945 & ~w44302;
assign w50154 = ~w7277 & w7011;
assign w50155 = w26962 & ~w25945;
assign w50156 = w26962 & w45513;
assign w50157 = w23843 & w27270;
assign w50158 = w23843 & w42339;
assign w50159 = w21801 & ~w28170;
assign w50160 = w21801 & ~w45694;
assign w50161 = ~w23843 & ~w27270;
assign w50162 = ~w23843 & ~w42339;
assign w50163 = ~w21801 & w28170;
assign w50164 = ~w21801 & w45694;
assign w50165 = w7052 & w7011;
assign w50166 = ~w35299 & w35311;
assign w50167 = w26699 & w27151;
assign w50168 = w26699 & ~w27153;
assign w50169 = ~w26699 & w27072;
assign w50170 = w26699 & ~w27072;
assign w50171 = w28186 & ~w28183;
assign w50172 = w28186 & ~w43623;
assign w50173 = ~w28594 & w6769;
assign w50174 = ~w28594 & ~w42378;
assign w50175 = w28594 & ~w6769;
assign w50176 = w28594 & w42378;
assign w50177 = ~w7085 & ~w7082;
assign w50178 = ~w7085 & w44311;
assign w50179 = w26877 & w27474;
assign w50180 = w28440 & ~w28424;
assign w50181 = (w2729 & ~w2381) | (w2729 & ~w39990) | (~w2381 & ~w39990);
assign w50182 = (~w4154 & ~w40165) | (~w4154 & ~w3890) | (~w40165 & ~w3890);
assign w50183 = (w4724 & ~w4623) | (w4724 & ~w40245) | (~w4623 & ~w40245);
assign w50184 = (~w8682 & ~w8390) | (~w8682 & ~w40653) | (~w8390 & ~w40653);
assign w50185 = (w9609 & w43428) | (w9609 & ~w9349) | (w43428 & ~w9349);
assign w50186 = (~w11152 & ~w44474) | (~w11152 & ~w11136) | (~w44474 & ~w11136);
assign w50187 = (w11888 & ~w12583) | (w11888 & ~w41103) | (~w12583 & ~w41103);
assign w50188 = (w12753 & ~w12583) | (w12753 & ~w41117) | (~w12583 & ~w41117);
assign w50189 = (~w12785 & ~w12583) | (~w12785 & ~w41119) | (~w12583 & ~w41119);
assign w50190 = (w945 & ~w12583) | (w945 & ~w41139) | (~w12583 & ~w41139);
assign w50191 = (~w945 & ~w12583) | (~w945 & ~w41143) | (~w12583 & ~w41143);
assign w50192 = (w13868 & ~w13372) | (w13868 & w50505) | (~w13372 & w50505);
assign w50193 = (w14607 & ~w13895) | (w14607 & w50506) | (~w13895 & w50506);
assign w50194 = (~w14764 & ~w14549) | (~w14764 & w47422) | (~w14549 & w47422);
assign w50195 = (~w14764 & ~w14545) | (~w14764 & w47425) | (~w14545 & w47425);
assign w50196 = (~w15240 & ~w6769) | (~w15240 & w48801) | (~w6769 & w48801);
assign w50197 = (~w14395 & ~w41299) | (~w14395 & ~w14383) | (~w41299 & ~w14383);
assign w50198 = (~w15574 & w15625) | (~w15574 & w44931) | (w15625 & w44931);
assign w50199 = (w14974 & ~w15643) | (w14974 & w48810) | (~w15643 & w48810);
assign w50200 = (~w15687 & ~w47454) | (~w15687 & ~w15672) | (~w47454 & ~w15672);
assign w50201 = (~w15537 & w16056) | (~w15537 & w44956) | (w16056 & w44956);
assign w50202 = (w16226 & ~w16531) | (w16226 & ~w41368) | (~w16531 & ~w41368);
assign w50203 = (~w17541 & w17341) | (~w17541 & ~w41458) | (w17341 & ~w41458);
assign w50204 = (~w18470 & ~w41526) | (~w18470 & ~w18158) | (~w41526 & ~w18158);
assign w50205 = (~w18866 & ~w18450) | (~w18866 & ~w41591) | (~w18450 & ~w41591);
assign w50206 = (w41531 & ~w45042) | (w41531 & ~w45043) | (~w45042 & ~w45043);
assign w50207 = (~w22229 & ~w41887) | (~w22229 & ~w21800) | (~w41887 & ~w21800);
assign w50208 = (w22255 & ~w41890) | (w22255 & ~w21800) | (~w41890 & ~w21800);
assign w50209 = (~w22137 & ~w42026) | (~w22137 & ~w22745) | (~w42026 & ~w22745);
assign w50210 = (~w23998 & ~w45319) | (~w23998 & ~w23640) | (~w45319 & ~w23640);
assign w50211 = (~w24264 & ~w23330) | (~w24264 & ~w42049) | (~w23330 & ~w42049);
assign w50212 = (w24288 & ~w42139) | (w24288 & ~w25340) | (~w42139 & ~w25340);
assign w50213 = (w24966 & ~w49118) | (w24966 & ~w25316) | (~w49118 & ~w25316);
assign w50214 = (~w14039 & ~w42352) | (~w14039 & ~w28076) | (~w42352 & ~w28076);
assign w50215 = (~w47790 & w45706) | (~w47790 & ~w47789) | (w45706 & ~w47789);
assign w50216 = (w27906 & ~w28019) | (w27906 & w49687) | (~w28019 & w49687);
assign w50217 = (w28473 & ~w28286) | (w28473 & ~w45748) | (~w28286 & ~w45748);
assign w50218 = (~w28677 & ~w45767) | (~w28677 & ~w29527) | (~w45767 & ~w29527);
assign w50219 = (~w30303 & ~w42473) | (~w30303 & ~w30308) | (~w42473 & ~w30308);
assign w50220 = (~w30246 & ~w30308) | (~w30246 & ~w29677) | (~w30308 & ~w29677);
assign w50221 = (~w45862 & ~w45863) | (~w45862 & ~w30946) | (~w45863 & ~w30946);
assign w50222 = (~w32849 & ~w45960) | (~w32849 & ~w32846) | (~w45960 & ~w32846);
assign w50223 = (w35180 & ~w42891) | (w35180 & ~w34899) | (~w42891 & ~w34899);
assign w50224 = (~w34897 & ~w34162) | (~w34897 & w49754) | (~w34162 & w49754);
assign w50225 = (w35693 & ~w42935) | (w35693 & ~w34591) | (~w42935 & ~w34591);
assign w50226 = (~w43108 & w36972) | (~w43108 & ~w46169) | (w36972 & ~w46169);
assign w50227 = (~w37168 & ~w43117) | (~w37168 & ~w36572) | (~w43117 & ~w36572);
assign w50228 = (w3525 & ~w40094) | (w3525 & ~w3241) | (~w40094 & ~w3241);
assign w50229 = w9862 & ~w10431;
assign w50230 = (w12176 & ~w41030) | (w12176 & ~w11814) | (~w41030 & ~w11814);
assign w50231 = (~w19016 & ~w41719) | (~w19016 & ~w18860) | (~w41719 & ~w18860);
assign w50232 = ~w33704 & ~w33628;
assign w50233 = (~w34830 & w49329) | (~w34830 & ~w34881) | (w49329 & ~w34881);
assign w50234 = w35640 & ~w35582;
assign w50235 = (~w35979 & ~w35463) | (~w35979 & w48256) | (~w35463 & w48256);
assign w50236 = ~w16517 & ~w16282;
assign w50237 = ~w23411 & ~w22723;
assign w50238 = (w33869 & ~w43752) | (w33869 & ~w32789) | (~w43752 & ~w32789);
assign w50239 = (~w32870 & ~w43769) | (~w32870 & ~w33736) | (~w43769 & ~w33736);
assign w50240 = (~w2789 & ~w43309) | (~w2789 & ~w2554) | (~w43309 & ~w2554);
assign w50241 = (w7519 & ~w43414) | (w7519 & ~w43415) | (~w43414 & ~w43415);
assign w50242 = (w14763 & w12666) | (w14763 & w48399) | (w12666 & w48399);
assign w50243 = (~w17374 & w16948) | (~w17374 & w46919) | (w16948 & w46919);
assign w50244 = (w25315 & w26181) | (w25315 & w49907) | (w26181 & w49907);
assign w50245 = (~w26995 & w28113) | (~w26995 & w49939) | (w28113 & w49939);
assign w50246 = ~w31823 & w30654;
assign w50247 = ~w24394 & ~w24577;
assign w50248 = (~w26995 & w27585) | (~w26995 & w49981) | (w27585 & w49981);
assign w50249 = (~w26995 & w27401) | (~w26995 & w49982) | (w27401 & w49982);
assign w50250 = ~w40537 | ~w7844;
assign w50251 = w42 & ~w25809;
assign w50252 = ~w957 & ~w1114;
assign w50253 = w957 & ~w1114;
assign w50254 = w1317 & ~w1323;
assign w50255 = ~w351 & w1314;
assign w50256 = ~w351 & ~w39799;
assign w50257 = ~w43938 & ~w1202;
assign w50258 = w1453 & ~w1445;
assign w50259 = w1453 & ~w1449;
assign w50260 = w3246 & w2967;
assign w50261 = ~w3239 & w51448;
assign w50262 = w40087 & ~w2946;
assign w50263 = (~w2946 & w40087) | (~w2946 & ~w3083) | (w40087 & ~w3083);
assign w50264 = w3833 & w3620;
assign w50265 = w3833 & ~w3464;
assign w50266 = w3845 & w3620;
assign w50267 = w3845 & ~w3464;
assign w50268 = w3965 & w3952;
assign w50269 = (w3937 & w51449) | (w3937 & w50268) | (w51449 & w50268);
assign w50270 = w4038 & ~w4115;
assign w50271 = w4038 & ~w40154;
assign w50272 = w5745 & w5827;
assign w50273 = ~w5745 & w5829;
assign w50274 = w5745 & w6167;
assign w50275 = ~w5745 & w6169;
assign w50276 = w40416 | ~w6074;
assign w50277 = (~w6074 & w40416) | (~w6074 & w6262) | (w40416 & w6262);
assign w50278 = ~w6586 & w40418;
assign w50279 = w5854 & ~w1320;
assign w50280 = ~w6262 & w6270;
assign w50281 = w6853 & w6857;
assign w50282 = w6853 & ~a[75];
assign w50283 = ~w6878 & ~w6390;
assign w50284 = ~w7132 & w493;
assign w50285 = ~w6720 & w48314;
assign w50286 = ~w7819 & w7839;
assign w50287 = (w7927 & w40545) | (w7927 & w7903) | (w40545 & w7903);
assign w50288 = (w7927 & w40545) | (w7927 & w7543) | (w40545 & w7543);
assign w50289 = w7954 & w7955;
assign w50290 = (w7807 & w40579) | (w7807 & w7903) | (w40579 & w7903);
assign w50291 = (w7807 & w40579) | (w7807 & w7543) | (w40579 & w7543);
assign w50292 = (~w7831 & w40590) | (~w7831 & w7903) | (w40590 & w7903);
assign w50293 = (~w7831 & w40590) | (~w7831 & w7543) | (w40590 & w7543);
assign w50294 = (w8246 & w40599) | (w8246 & w7903) | (w40599 & w7903);
assign w50295 = (w8246 & w40599) | (w8246 & w7543) | (w40599 & w7543);
assign w50296 = (w3646 & w40609) | (w3646 & w7903) | (w40609 & w7903);
assign w50297 = (w3646 & w40609) | (w3646 & w7543) | (w40609 & w7543);
assign w50298 = w8125 & ~w8183;
assign w50299 = w8125 & ~w44415;
assign w50300 = w11293 & w11298;
assign w50301 = w11296 & w4838;
assign w50302 = ~w10673 & ~w11310;
assign w50303 = ~w11303 & w11316;
assign w50304 = w40955 & ~w11343;
assign w50305 = (~w11343 & w40955) | (~w11343 & ~w11331) | (w40955 & ~w11331);
assign w50306 = ~w11303 & ~w11577;
assign w50307 = w11506 & w5745;
assign w50308 = ~w11151 & w10570;
assign w50309 = w11706 & w11781;
assign w50310 = ~w12121 & ~w12123;
assign w50311 = ~w12329 & w2285;
assign w50312 = w12399 & w5330;
assign w50313 = ~w12228 & w945;
assign w50314 = ~w7924 & w12034;
assign w50315 = ~w7924 & ~w12049;
assign w50316 = ~w11922 & ~w12747;
assign w50317 = ~w11922 & ~w12049;
assign w50318 = w12637 & ~w6769;
assign w50319 = w12637 & ~w11902;
assign w50320 = ~w12637 & w6769;
assign w50321 = ~w12581 & w12787;
assign w50322 = ~w12854 & w2896;
assign w50323 = ~w12288 & w12259;
assign w50324 = ~w12352 & w12335;
assign w50325 = w12999 & w12998;
assign w50326 = (w13010 & w12580) | (w13010 & w50507) | (w12580 & w50507);
assign w50327 = (w12602 & w12580) | (w12602 & w50508) | (w12580 & w50508);
assign w50328 = ~w13112 & ~w12465;
assign w50329 = ~w13112 & w44645;
assign w50330 = ~w13112 & w12471;
assign w50331 = (~w12573 & w12580) | (~w12573 & w50509) | (w12580 & w50509);
assign w50332 = w13220 & w12412;
assign w50333 = w13220 & w12724;
assign w50334 = ~w13244 & w13246;
assign w50335 = ~w13260 & w13262;
assign w50336 = ~w13305 & w13306;
assign w50337 = w13229 & w252;
assign w50338 = w12666 & ~w493;
assign w50339 = ~w13754 & w754;
assign w50340 = ~w13379 & w13779;
assign w50341 = ~w13379 & w13781;
assign w50342 = ~w14590 & ~w14583;
assign w50343 = w15906 & w41393;
assign w50344 = w17188 & w17191;
assign w50345 = w17357 & ~w17752;
assign w50346 = w22477 & w22802;
assign w50347 = ~w25690 & ~w57;
assign w50348 = w25690 & w57;
assign w50349 = (~w25062 & w50023) | (~w25062 & w25059) | (w50023 & w25059);
assign w50350 = (~w25062 & w50023) | (~w25062 & w25818) | (w50023 & w25818);
assign w50351 = (~w26255 & w50029) | (~w26255 & w25059) | (w50029 & w25059);
assign w50352 = (~w26255 & w50029) | (~w26255 & w25818) | (w50029 & w25818);
assign w50353 = w25850 & ~w25359;
assign w50354 = w26832 & w26838;
assign w50355 = w27164 & w27167;
assign w50356 = ~w27146 & ~w3646;
assign w50357 = ~w27509 & w11870;
assign w50358 = ~w27521 & ~w15681;
assign w50359 = w27521 & w15681;
assign w50360 = w27577 & w27642;
assign w50361 = ~w27577 & w27644;
assign w50362 = ~w27537 & w27646;
assign w50363 = ~w25851 & w42336;
assign w50364 = ~w25851 & ~w45688;
assign w50365 = (w24874 & w49164) | (w24874 & ~w42336) | (w49164 & ~w42336);
assign w50366 = (w24874 & w49164) | (w24874 & w45688) | (w49164 & w45688);
assign w50367 = w25851 & ~w42336;
assign w50368 = w25851 & w45688;
assign w50369 = w49164 & ~w42336;
assign w50370 = w49164 & w45688;
assign w50371 = ~w22767 & ~w42336;
assign w50372 = ~w22767 & w49169;
assign w50373 = ~w21801 & ~w42336;
assign w50374 = ~w21801 & w49165;
assign w50375 = ~w28050 & w28307;
assign w50376 = ~w27742 & w27487;
assign w50377 = w28418 & w42336;
assign w50378 = w28418 & ~w49179;
assign w50379 = ~w28691 & ~w28690;
assign w50380 = w29188 & w28250;
assign w50381 = ~w29188 & ~w28250;
assign w50382 = ~w29157 & ~w28207;
assign w50383 = w29157 & w29242;
assign w50384 = w29265 & w29202;
assign w50385 = ~w30803 & ~w29276;
assign w50386 = w32192 & ~w33569;
assign w50387 = w32192 & w46008;
assign w50388 = ~w35130 & w24874;
assign w50389 = w35130 & ~w24874;
assign w50390 = w35325 & w35567;
assign w50391 = w35980 & w43022;
assign w50392 = w36420 & w7315;
assign w50393 = ~w38060 & ~w38063;
assign w50394 = w43354 & w252;
assign w50395 = (w252 & w43354) | (w252 & w4055) | (w43354 & w4055);
assign w50396 = w4166 & ~w400;
assign w50397 = w4166 & ~w40160;
assign w50398 = w4172 & ~w400;
assign w50399 = w4172 & ~w40160;
assign w50400 = w29093 & ~w28038;
assign w50401 = ~w35978 & ~w36016;
assign w50402 = ~w35978 & w36038;
assign w50403 = ~w35978 & ~w36057;
assign w50404 = ~w35978 & w36075;
assign w50405 = ~w35978 & w36103;
assign w50406 = ~w35978 & w36123;
assign w50407 = ~w35978 & w36130;
assign w50408 = ~w35978 & w36145;
assign w50409 = ~w35978 & w36152;
assign w50410 = ~w35978 & w36190;
assign w50411 = ~w35978 & w36750;
assign w50412 = ~w35978 & ~w35946;
assign w50413 = w6262 & w6178;
assign w50414 = w6178 & ~w6263;
assign w50415 = w7267 & ~w7115;
assign w50416 = w8380 & ~w8391;
assign w50417 = w8303 & ~w8391;
assign w50418 = w3 & w4003;
assign w50419 = w3 & ~w40149;
assign w50420 = w6537 & w7091;
assign w50421 = ~w6537 & w7093;
assign w50422 = ~w13337 & ~w6769;
assign w50423 = w13337 & w13409;
assign w50424 = ~w13337 & w13454;
assign w50425 = w13337 & w13456;
assign w50426 = ~w13337 & w13649;
assign w50427 = w13337 & w13648;
assign w50428 = ~w13337 & w13664;
assign w50429 = w13337 & w13663;
assign w50430 = w13337 & ~w13377;
assign w50431 = ~w13337 & ~w3;
assign w50432 = ~w13337 & ~w13267;
assign w50433 = ~w13337 & ~w13302;
assign w50434 = ~w13337 & w13974;
assign w50435 = ~w13382 & ~w13888;
assign w50436 = w13382 & w13888;
assign w50437 = w12613 & w12027;
assign w50438 = ~w12613 & ~w12736;
assign w50439 = ~w12613 & w13171;
assign w50440 = ~w12613 & w12527;
assign w50441 = w12613 & ~w2006;
assign w50442 = w12613 & w2558;
assign w50443 = ~w13355 & w13917;
assign w50444 = w13355 & ~w13917;
assign w50445 = ~w11138 & w13654;
assign w50446 = ~w11138 & w44709;
assign w50447 = w13369 & w13779;
assign w50448 = w13369 & w13781;
assign w50449 = ~w13280 & w13820;
assign w50450 = ~w13985 & w41184;
assign w50451 = ~w12613 & w12626;
assign w50452 = w14457 & w1120;
assign w50453 = ~w14457 & ~w1120;
assign w50454 = ~w13381 & w4430;
assign w50455 = ~w13381 & ~w4838;
assign w50456 = w13381 & w4838;
assign w50457 = w13381 & ~w4056;
assign w50458 = w13381 & w3242;
assign w50459 = w13381 & ~w4430;
assign w50460 = ~w13381 & w13760;
assign w50461 = w13381 & w13762;
assign w50462 = w13381 & ~w13759;
assign w50463 = ~w13381 & w13759;
assign w50464 = ~w13381 & w13794;
assign w50465 = w13381 & w13796;
assign w50466 = ~w13381 & w13800;
assign w50467 = w13381 & w13802;
assign w50468 = ~w13381 & w13811;
assign w50469 = w13381 & w13813;
assign w50470 = ~w13381 & w13889;
assign w50471 = w13381 & w13891;
assign w50472 = ~w13381 & w1541;
assign w50473 = ~w13381 & w1738;
assign w50474 = w13381 & ~w1541;
assign w50475 = w13381 & ~w1738;
assign w50476 = ~w13381 & ~w2006;
assign w50477 = ~w14327 & w14328;
assign w50478 = ~w14360 & w13681;
assign w50479 = w14360 & w14364;
assign w50480 = ~w14329 & w11870;
assign w50481 = ~w14401 & w14402;
assign w50482 = w14401 & w14404;
assign w50483 = ~w14401 & ~w13709;
assign w50484 = w14401 & w13709;
assign w50485 = ~w14448 & ~w13982;
assign w50486 = w43487 & ~w14491;
assign w50487 = ~w14058 & ~w13880;
assign w50488 = ~w14628 & w13804;
assign w50489 = ~w13934 & w13713;
assign w50490 = ~w13934 & w13391;
assign w50491 = ~w13934 & w13469;
assign w50492 = ~w13934 & ~w14167;
assign w50493 = ~w13934 & w14173;
assign w50494 = ~w13934 & w13516;
assign w50495 = ~w13934 & ~w13579;
assign w50496 = ~w13934 & w14237;
assign w50497 = ~w13934 & ~w14259;
assign w50498 = ~w13934 & w13612;
assign w50499 = ~w13934 & ~w13500;
assign w50500 = ~w13934 & w13979;
assign w50501 = ~w13934 & ~w13544;
assign w50502 = ~w13934 & w493;
assign w50503 = ~w13934 & ~w612;
assign w50504 = ~w13934 & ~w3;
assign w50505 = w13868 & ~w13380;
assign w50506 = w14607 & ~w13930;
assign w50507 = ~w12421 & w13010;
assign w50508 = ~w12421 & w12602;
assign w50509 = ~w12421 & ~w12573;
assign w50510 = ~w11064 & w11304;
assign w50511 = ~w10673 & w11312;
assign w50512 = w11748 & w11781;
assign w50513 = (~w11874 & w40985) | (~w11874 & ~w11148) | (w40985 & ~w11148);
assign w50514 = (~w11874 & w40985) | (~w11874 & w11787) | (w40985 & w11787);
assign w50515 = ~w11813 & w11880;
assign w50516 = w11705 & w11344;
assign w50517 = ~w12463 & w612;
assign w50518 = w41094 & w12544;
assign w50519 = (w12544 & w41094) | (w12544 & w11813) | (w41094 & w11813);
assign w50520 = ~w11770 & w12548;
assign w50521 = ~w12050 & ~w12028;
assign w50522 = ~w12710 & w8666;
assign w50523 = w12710 & ~w8666;
assign w50524 = ~w12743 & ~w12700;
assign w50525 = ~w12032 & w12042;
assign w50526 = w41114 & w47286;
assign w50527 = (w47286 & w41114) | (w47286 & ~w12030) | (w41114 & ~w12030);
assign w50528 = w12822 & w5330;
assign w50529 = ~w5745 & w12184;
assign w50530 = ~w3646 & w12159;
assign w50531 = ~w3646 & w41121;
assign w50532 = ~w12640 & w12392;
assign w50533 = ~w12822 & ~w5330;
assign w50534 = ~w12090 & w12192;
assign w50535 = ~w12666 & w493;
assign w50536 = w12772 & w12612;
assign w50537 = ~w12533 & w12565;
assign w50538 = ~w13166 & ~w12534;
assign w50539 = w13202 & w126;
assign w50540 = w13202 & w161;
assign w50541 = w13211 & ~w57;
assign w50542 = ~w13211 & w57;
assign w50543 = ~w13232 & ~w252;
assign w50544 = w12695 & w13396;
assign w50545 = w12665 & ~w13450;
assign w50546 = ~w12665 & w13450;
assign w50547 = w13432 & w13459;
assign w50548 = ~w13823 & w13837;
assign w50549 = ~w13756 & ~w754;
assign w50550 = ~w13783 & w13129;
assign w50551 = w13783 & ~w13129;
assign w50552 = ~w13799 & ~w13849;
assign w50553 = w13367 & ~w13146;
assign w50554 = ~w13832 & ~w13838;
assign w50555 = ~w13082 & ~w1120;
assign w50556 = ~w13823 & ~w13939;
assign w50557 = ~w13447 & w13438;
assign w50558 = w13447 & ~w13438;
assign w50559 = w14453 & ~w1320;
assign w50560 = ~w14453 & w1320;
assign w50561 = w11277 & w4430;
assign w50562 = ~w11861 & w12085;
assign w50563 = ~w11861 & w12107;
assign w50564 = ~w11861 & w12138;
assign w50565 = ~w11861 & w1541;
assign w50566 = w46541 & w46540;
assign w50567 = (w46540 & w46541) | (w46540 & w11813) | (w46541 & w11813);
assign w50568 = ~w12434 & ~w493;
assign w50569 = w12434 & ~w493;
assign w50570 = w12434 & w493;
assign w50571 = ~w12434 & w493;
assign w50572 = w12497 & ~w12491;
assign w50573 = w12497 & w41083;
assign w50574 = ~w12268 & ~w12266;
assign w50575 = ~w12268 & w41049;
assign w50576 = w12635 & ~w7924;
assign w50577 = ~w12052 & ~w12034;
assign w50578 = ~w12052 & w12747;
assign w50579 = w41160 & w13258;
assign w50580 = ~w41160 & ~w13258;
assign w50581 = w41166 & w13312;
assign w50582 = ~w41166 & w13314;
assign w50583 = w41160 & w13319;
assign w50584 = ~w41160 & w13321;
assign w50585 = ~w41166 & w13329;
assign w50586 = (~w14491 & w43487) | (~w14491 & ~w14021) | (w43487 & ~w14021);
assign w50587 = (~w14491 & w43487) | (~w14491 & w41230) | (w43487 & w41230);
assign w50588 = w12584 & ~w12393;
assign w50589 = w12887 & w2558;
assign w50590 = ~w12595 & w12331;
assign w50591 = ~w12887 & ~w2558;
assign w50592 = w12648 & ~w10419;
assign w50593 = ~w12648 & w10419;
assign w50594 = ~w4056 & ~w12961;
assign w50595 = ~w4056 & w41135;
assign w50596 = ~w12615 & ~w12464;
assign w50597 = ~w13337 & w12953;
assign w50598 = ~w13337 & ~w12824;
assign w50599 = ~w13337 & ~w2558;
assign w50600 = ~w13337 & w13548;
assign w50601 = ~w13337 & w13555;
assign w50602 = ~w13337 & ~w12855;
assign w50603 = ~w13337 & w13577;
assign w50604 = ~w13337 & ~w12980;
assign w50605 = ~w13337 & ~w12871;
assign w50606 = ~w13337 & ~w754;
assign w50607 = ~w13337 & ~w493;
assign w50608 = ~w13337 & ~w612;
assign w50609 = w13337 & w13863;
assign w50610 = ~w13337 & w13376;
assign w50611 = ~w13337 & ~w351;
assign w50612 = ~w13855 & w14033;
assign w50613 = ~w12623 & ~w12624;
assign w50614 = ~w13165 & w12543;
assign w50615 = w13540 & w13532;
assign w50616 = ~w13540 & ~w13532;
assign w50617 = w44729 | ~w493;
assign w50618 = (~w493 & w44729) | (~w493 & w13808) | (w44729 & w13808);
assign w50619 = w13808 & w13810;
assign w50620 = w41166 & w13327;
assign w50621 = ~w13738 & w14619;
assign w50622 = ~a[120] & a[121];
assign w50623 = w106 & ~w18;
assign w50624 = a[122] & ~w3;
assign w50625 = ~w39648 & w111;
assign w50626 = ~w39648 & w109;
assign w50627 = ~w155 & w3;
assign w50628 = ~w113 & ~w157;
assign w50629 = ~w211 & ~w42;
assign w50630 = ~w410 & ~w409;
assign w50631 = (~w410 & ~w398) | (~w410 & w50687) | (~w398 & w50687);
assign w50632 = (~w50631 & w50781) | (~w50631 & w50782) | (w50781 & w50782);
assign w50633 = w420 & ~w409;
assign w50634 = (w420 & ~w398) | (w420 & w50749) | (~w398 & w50749);
assign w50635 = w431 & ~w427;
assign w50636 = (w431 & ~w398) | (w431 & w50688) | (~w398 & w50688);
assign w50637 = w433 & w427;
assign w50638 = w398 & w50689;
assign w50639 = w460 & w427;
assign w50640 = w398 & w50750;
assign w50641 = w462 & ~w427;
assign w50642 = (w462 & ~w398) | (w462 & w50751) | (~w398 & w50751);
assign w50643 = ~w443 & w479;
assign w50644 = (~w50643 & w50690) | (~w50643 & w50691) | (w50690 & w50691);
assign w50645 = (~w50643 & w50692) | (~w50643 & w50693) | (w50692 & w50693);
assign w50646 = (~w50643 & w50694) | (~w50643 & w50695) | (w50694 & w50695);
assign w50647 = ~w492 & w50752;
assign w50648 = ~w492 & w50783;
assign w50649 = (w408 & w50739) | (w408 & w50784) | (w50739 & w50784);
assign w50650 = (~w408 & w50740) | (~w408 & w50785) | (w50740 & w50785);
assign w50651 = w39703 & w524;
assign w50652 = (w524 & w39703) | (w524 & w480) | (w39703 & w480);
assign w50653 = (w419 & w46394) | (w419 & w50697) | (w46394 & w50697);
assign w50654 = (w419 & w39707) | (w419 & w480) | (w39707 & w480);
assign w50655 = ~w480 & w39708;
assign w50656 = w39712 & w572;
assign w50657 = (w572 & w39712) | (w572 & w480) | (w39712 & w480);
assign w50658 = w39713 & ~w577;
assign w50659 = (~w577 & w39713) | (~w577 & w480) | (w39713 & w480);
assign w50660 = ~w480 & w39714;
assign w50661 = w39716 & w586;
assign w50662 = (w586 & w39716) | (w586 & w480) | (w39716 & w480);
assign w50663 = ~w480 & w39719;
assign w50664 = w39720 & w596;
assign w50665 = (w596 & w39720) | (w596 & w480) | (w39720 & w480);
assign w50666 = ~w609 & ~w552;
assign w50667 = ~w609 & w558;
assign w50668 = (~w3 & ~w612) | (~w3 & w50753) | (~w612 & w50753);
assign w50669 = w612 & w50754;
assign w50670 = ~a[125] & ~a[122];
assign w50671 = w103 & ~w3;
assign w50672 = ~w375 & w43247;
assign w50673 = w404 & w330;
assign w50674 = (w404 & w370) | (w404 & w50755) | (w370 & w50755);
assign w50675 = ~w370 & w50756;
assign w50676 = ~w370 & w50757;
assign w50677 = w427 & w371;
assign w50678 = w449 & ~w330;
assign w50679 = w449 & w371;
assign w50680 = ~w452 & w330;
assign w50681 = (~w452 & w370) | (~w452 & w50842) | (w370 & w50842);
assign w50682 = ~w369 & w273;
assign w50683 = ~w155 & w42;
assign w50684 = w231 & w346;
assign w50685 = w231 & a[118];
assign w50686 = a[115] & w371;
assign w50687 = w388 & ~w410;
assign w50688 = w388 & w431;
assign w50689 = ~w388 & w433;
assign w50690 = ~w492 & ~w479;
assign w50691 = ~w492 & ~w465;
assign w50692 = (w3 & ~w478) | (w3 & w50758) | (~w478 & w50758);
assign w50693 = (w3 & w459) | (w3 & w50759) | (w459 & w50759);
assign w50694 = (~w3 & ~w478) | (~w3 & w50760) | (~w478 & w50760);
assign w50695 = (~w3 & w459) | (~w3 & w50761) | (w459 & w50761);
assign w50696 = w3 & w464;
assign w50697 = ~w548 & w419;
assign w50698 = ~w56 & ~a[120];
assign w50699 = ~w43866 & ~w3;
assign w50700 = w56 & w39663;
assign w50701 = ~w242 & ~w245;
assign w50702 = w56 & a[120];
assign w50703 = ~w199 & w285;
assign w50704 = w199 & w286;
assign w50705 = w274 & w329;
assign w50706 = w199 & w335;
assign w50707 = w199 & a[118];
assign w50708 = ~w199 & ~a[118];
assign w50709 = w199 & ~w57;
assign w50710 = ~w199 & w57;
assign w50711 = ~w39694 & w42;
assign w50712 = ~w475 & ~w42;
assign w50713 = ~w441 & ~w3;
assign w50714 = w545 & w512;
assign w50715 = ~w528 & w3;
assign w50716 = ~w547 & w639;
assign w50717 = w547 & w606;
assign w50718 = w39729 & ~w661;
assign w50719 = (~w661 & w39729) | (~w661 & ~w547) | (w39729 & ~w547);
assign w50720 = ~w547 & w657;
assign w50721 = w547 & w668;
assign w50722 = ~w547 & w667;
assign w50723 = w547 & w673;
assign w50724 = ~w547 & w675;
assign w50725 = ~w512 & ~w80;
assign w50726 = w721 & ~w558;
assign w50727 = w721 & ~w603;
assign w50728 = w724 & w725;
assign w50729 = w724 & ~w535;
assign w50730 = w734 & w839;
assign w50731 = ~w734 & ~w839;
assign w50732 = ~w752 & w849;
assign w50733 = w734 & w857;
assign w50734 = ~w734 & w859;
assign w50735 = w752 & w870;
assign w50736 = ~w752 & w882;
assign w50737 = w752 & w917;
assign w50738 = ~w752 & ~w909;
assign w50739 = w252 & ~w57;
assign w50740 = ~w252 & w57;
assign w50741 = ~w80 & w551;
assign w50742 = w557 & w3;
assign w50743 = w163 & w714;
assign w50744 = w747 & ~w750;
assign w50745 = w43251 & w80;
assign w50746 = (w80 & w43251) | (w80 & ~w752) | (w43251 & ~w752);
assign w50747 = w747 & w895;
assign w50748 = w752 & w936;
assign w50749 = w388 & w420;
assign w50750 = ~w388 & w460;
assign w50751 = w388 & w462;
assign w50752 = ~w441 & w50696;
assign w50753 = ~w39746 & ~w3;
assign w50754 = w39746 & w3;
assign w50755 = ~w369 & w404;
assign w50756 = w369 & w406;
assign w50757 = w369 & w409;
assign w50758 = w472 & w3;
assign w50759 = ~w464 & w3;
assign w50760 = w472 & ~w3;
assign w50761 = ~w464 & ~w3;
assign w50762 = ~w234 & a[117];
assign w50763 = ~w443 & ~w473;
assign w50764 = w43884 | ~w42;
assign w50765 = (~w42 & w43884) | (~w42 & ~w507) | (w43884 & ~w507);
assign w50766 = ~w507 & w490;
assign w50767 = w397 & w562;
assign w50768 = w39723 | w630;
assign w50769 = (w630 & w39723) | (w630 & w547) | (w39723 & w547);
assign w50770 = ~w547 & w39724;
assign w50771 = w39727 | w644;
assign w50772 = (w644 & w39727) | (w644 & w547) | (w39727 & w547);
assign w50773 = ~w547 & w39728;
assign w50774 = w39730 | w678;
assign w50775 = (w678 & w39730) | (w678 & w547) | (w39730 & w547);
assign w50776 = w547 & w39731;
assign w50777 = ~w80 & w547;
assign w50778 = w709 & w3;
assign w50779 = w752 & w642;
assign w50780 = w521 & w700;
assign w50781 = ~w252 & ~w50630;
assign w50782 = ~w252 & w39688;
assign w50783 = w50713 & ~w464;
assign w50784 = ~w57 & ~w50632;
assign w50785 = w57 & w50632;
assign w50786 = ~w155 & ~w161;
assign w50787 = ~w113 & ~w162;
assign w50788 = w6 & w171;
assign w50789 = ~a[123] & w19;
assign w50790 = w182 & ~w188;
assign w50791 = w90 & w163;
assign w50792 = ~w87 & w163;
assign w50793 = w56 & ~w236;
assign w50794 = ~w56 & w236;
assign w50795 = w199 & w254;
assign w50796 = ~w199 & w256;
assign w50797 = w216 & w3;
assign w50798 = ~w254 & w3;
assign w50799 = w189 & w279;
assign w50800 = w199 & w287;
assign w50801 = w189 & w278;
assign w50802 = w254 & ~w3;
assign w50803 = w199 & w299;
assign w50804 = ~w199 & w301;
assign w50805 = ~w199 & ~w335;
assign w50806 = w56 & ~w353;
assign w50807 = ~w56 & w353;
assign w50808 = ~w196 & ~w57;
assign w50809 = ~w234 & ~w402;
assign w50810 = w234 & w402;
assign w50811 = w234 & ~a[116];
assign w50812 = ~w234 & a[116];
assign w50813 = ~w349 & ~w57;
assign w50814 = w349 & w57;
assign w50815 = w234 & w353;
assign w50816 = ~w467 & w329;
assign w50817 = ~w305 & w228;
assign w50818 = ~a[113] & ~w401;
assign w50819 = w563 & w351;
assign w50820 = w397 & a[114];
assign w50821 = ~w397 & ~a[114];
assign w50822 = ~w563 & ~w351;
assign w50823 = a[114] & ~w409;
assign w50824 = w252 & ~w409;
assign w50825 = w252 & w50823;
assign w50826 = a[112] & a[113];
assign w50827 = w547 & ~w624;
assign w50828 = ~w547 & w628;
assign w50829 = w654 & a[111];
assign w50830 = ~w652 & ~a[111];
assign w50831 = ~w652 & ~w50829;
assign w50832 = ~w400 & ~w50830;
assign w50833 = ~w400 & ~w50831;
assign w50834 = ~a[111] & ~w400;
assign w50835 = w654 & ~w400;
assign w50836 = ~w654 & w400;
assign w50837 = w528 & w42;
assign w50838 = ~w528 & w42;
assign w50839 = w738 & w42;
assign w50840 = ~w3 & w714;
assign w50841 = ~w738 & ~w42;
assign w50842 = ~w369 & ~w452;
assign w50843 = w654 & ~a[111];
assign w50844 = w654 & w50834;
assign w50845 = w776 & ~w720;
assign w50846 = w776 & ~w39750;
assign w50847 = w743 & w714;
assign w50848 = w738 & ~w42;
assign w50849 = w547 & a[111];
assign w50850 = ~w547 & ~a[111];
assign w50851 = a[110] & ~w652;
assign w50852 = w547 & ~w880;
assign w50853 = ~a[109] & ~w653;
assign w50854 = ~w547 & w880;
assign w50855 = ~w650 & ~w886;
assign w50856 = w752 & w885;
assign w50857 = w863 & ~w400;
assign w50858 = ~w547 & ~w903;
assign w50859 = w493 & ~w905;
assign w50860 = ~w547 & ~a[110];
assign w50861 = ~a[109] & a[110];
assign w50862 = ~w911 & ~w916;
assign w50863 = ~w771 & w963;
assign w50864 = w771 & ~w806;
assign w50865 = ~w986 & a[107];
assign w50866 = ~w50865 & ~w879;
assign w50867 = w986 & ~a[107];
assign w50868 = w547 & ~w1001;
assign w50869 = a[108] & a[109];
assign w50870 = ~w547 & w1001;
assign w50871 = ~w884 & ~w493;
assign w50872 = ~w876 & w351;
assign w50873 = w876 & ~w351;
assign w50874 = w57 & ~w792;
assign w50875 = ~w1079 & w1106;
assign w50876 = ~w966 & w956;
assign w50877 = w984 & w1208;
assign w50878 = w1216 & ~w1114;
assign w50879 = w1216 & w50253;
assign w50880 = a[104] & a[105];
assign w50881 = w1228 & ~w1229;
assign w50882 = w1227 & ~w1231;
assign w50883 = ~w983 & ~w1241;
assign w50884 = w984 & w1250;
assign w50885 = ~w984 & w1252;
assign w50886 = ~w983 & ~w1257;
assign w50887 = ~w983 & w1271;
assign w50888 = w984 & ~w1149;
assign w50889 = ~w1322 & ~w57;
assign w50890 = ~w1166 & w1332;
assign w50891 = ~w1331 & ~w1333;
assign w50892 = ~w984 & ~a[104];
assign w50893 = w984 & ~w945;
assign w50894 = ~w984 & w945;
assign w50895 = a[102] & a[103];
assign w50896 = ~w984 & ~w1354;
assign w50897 = w984 & ~w1356;
assign w50898 = w1358 & w945;
assign w50899 = ~w1352 & w945;
assign w50900 = w984 & a[104];
assign w50901 = w1352 & ~w945;
assign w50902 = ~w1358 & ~w945;
assign w50903 = w984 & ~w1240;
assign w50904 = ~w984 & w1244;
assign w50905 = w1276 & ~w493;
assign w50906 = w1254 & ~w612;
assign w50907 = ~w1254 & w612;
assign w50908 = w1292 & ~w1428;
assign w50909 = w1308 & ~w1314;
assign w50910 = w1317 & w1305;
assign w50911 = w1429 & ~w1431;
assign w50912 = w1437 & w1432;
assign w50913 = w1317 & w1138;
assign w50914 = w1200 & w80;
assign w50915 = w1178 & ~w1187;
assign w50916 = ~w1178 & ~w1220;
assign w50917 = ~w1497 & ~w42;
assign w50918 = (w1504 & w51450) | (w1504 & w51451) | (w51450 & w51451);
assign w50919 = w42 & w1516;
assign w50920 = ~w1525 & ~w1524;
assign w50921 = w1467 & w80;
assign w50922 = ~w1467 & w80;
assign w50923 = w1317 & ~w1551;
assign w50924 = ~a[101] & ~w1351;
assign w50925 = ~w1317 & w1551;
assign w50926 = ~w1552 & ~w1120;
assign w50927 = ~w1317 & ~a[102];
assign w50928 = w1317 & a[102];
assign w50929 = ~w984 & w1577;
assign w50930 = w984 & ~w1577;
assign w50931 = ~w1317 & ~w1580;
assign w50932 = w1317 & w1580;
assign w50933 = ~w1376 & w754;
assign w50934 = ~w1393 & ~w1613;
assign w50935 = w1393 & w1613;
assign w50936 = ~w1418 & ~w1626;
assign w50937 = w1418 & w1626;
assign w50938 = (w1465 & w51452) | (w1465 & w51453) | (w51452 & w51453);
assign w50939 = w1629 & ~w1526;
assign w50940 = ~w1632 & w1509;
assign w50941 = ~w1632 & w1526;
assign w50942 = w400 & ~w50258;
assign w50943 = w400 & ~w50259;
assign w50944 = ~w1674 & ~w43942;
assign w50945 = ~w1674 & ~w1508;
assign w50946 = ~w1671 & w1680;
assign w50947 = w1683 & w57;
assign w50948 = ~w1467 & ~w80;
assign w50949 = w1467 & ~w80;
assign w50950 = ~w1686 & w1704;
assign w50951 = w1510 & ~w1483;
assign w50952 = w1510 & ~w39863;
assign w50953 = w1513 & ~w1483;
assign w50954 = w1513 & ~w39863;
assign w50955 = ~w1512 & w1514;
assign w50956 = w1506 & w1514;
assign w50957 = w1506 & w50955;
assign w50958 = ~w1504 & ~w42;
assign w50959 = w1721 & ~w42;
assign w50960 = w1721 & ~w39864;
assign w50961 = w1704 & w1722;
assign w50962 = w1724 & ~w1681;
assign w50963 = ~w1497 & w1514;
assign w50964 = ~w1497 & w50955;
assign w50965 = w1724 & w1648;
assign w50966 = w1735 & w1706;
assign w50967 = w1735 & ~w1706;
assign w50968 = ~w1544 & w1473;
assign w50969 = w1544 & ~w1473;
assign w50970 = ~a[100] & ~w1526;
assign w50971 = w1771 & ~w1553;
assign w50972 = ~w1774 & w1120;
assign w50973 = w1805 & ~w1526;
assign w50974 = ~w1320 & ~w1806;
assign w50975 = ~w1320 & ~w1809;
assign w50976 = w1841 & w80;
assign w50977 = ~w1853 & w47011;
assign w50978 = ~w1853 & w1595;
assign w50979 = w1570 & ~w1599;
assign w50980 = ~w1722 & ~w1868;
assign w50981 = ~w1612 & w612;
assign w50982 = w1612 & w612;
assign w50983 = (~w80 & w1738) | (~w80 & w51454) | (w1738 & w51454);
assign w50984 = w1675 & w1435;
assign w50985 = ~w1675 & ~w1435;
assign w50986 = ~w493 & ~w612;
assign w50987 = ~w1612 & ~w612;
assign w50988 = w1612 & ~w612;
assign w50989 = ~w1844 & ~w1955;
assign w50990 = w1968 & ~w1757;
assign w50991 = w1968 & w47018;
assign w50992 = w1723 & ~w1727;
assign w50993 = ~w1716 & ~w1970;
assign w50994 = ~w1975 & ~w1974;
assign w50995 = w1716 & ~w42;
assign w50996 = w1995 & ~w1757;
assign w50997 = ~w1844 & w3;
assign w50998 = w1844 & ~w3;
assign w50999 = w2005 & w1926;
assign w51000 = w2033 & w57;
assign w51001 = w1921 & ~w57;
assign w51002 = w1927 & ~w1956;
assign w51003 = w57 & w1915;
assign w51004 = w2089 & ~w80;
assign w51005 = ~w2000 & w2097;
assign w51006 = ~w2157 & ~w1541;
assign w51007 = ~w1875 & ~w1876;
assign w51008 = w1875 & w1876;
assign w51009 = ~w1803 & w2222;
assign w51010 = w2005 & w1851;
assign w51011 = ~w2005 & ~a[96];
assign w51012 = w2005 & a[96];
assign w51013 = ~w2005 & w2313;
assign w51014 = w2005 & ~w2313;
assign w51015 = ~a[95] & ~w2156;
assign w51016 = ~w1981 & w2302;
assign w51017 = w2100 & w2337;
assign w51018 = ~w2005 & w1738;
assign w51019 = w2340 & w2157;
assign w51020 = ~w2340 & ~w2157;
assign w51021 = ~w2035 & ~a[97];
assign w51022 = w2005 & w1801;
assign w51023 = ~w2005 & w2234;
assign w51024 = ~w2232 & w2277;
assign w51025 = ~w1981 & ~w493;
assign w51026 = ~w2239 & w2264;
assign w51027 = ~w1981 & ~w754;
assign w51028 = w2433 & w2259;
assign w51029 = w2433 & w47033;
assign w51030 = w2005 & w1866;
assign w51031 = ~w2005 & w2226;
assign w51032 = w2482 & ~w2484;
assign w51033 = w2111 & w2100;
assign w51034 = ~w2103 & ~w2100;
assign w51035 = ~w2103 & ~w51033;
assign w51036 = w2512 & ~w51034;
assign w51037 = w2512 & ~w51035;
assign w51038 = ~w2517 & ~w2499;
assign w51039 = ~w2301 & ~w57;
assign w51040 = ~w2301 & ~w44002;
assign w51041 = w2550 & ~w2564;
assign w51042 = ~w2566 & ~w80;
assign w51043 = ~w2573 & ~w2572;
assign w51044 = ~w2491 & w2576;
assign w51045 = w2528 & ~w2530;
assign w51046 = ~w2528 & w2530;
assign w51047 = w2516 & ~w2585;
assign w51048 = w2106 & ~w51034;
assign w51049 = w2106 & ~w51035;
assign w51050 = w2600 & ~w42;
assign w51051 = w1965 & w51048;
assign w51052 = w1965 & w51049;
assign w51053 = ~w2604 & ~w2605;
assign w51054 = w2517 & w2493;
assign w51055 = ~w39975 & ~w2658;
assign w51056 = ~w2654 & ~w2659;
assign w51057 = ~w2407 & ~w252;
assign w51058 = w2407 & ~w252;
assign w51059 = w2516 & ~w2392;
assign w51060 = w2359 & ~w2379;
assign w51061 = ~w2456 & ~w2474;
assign w51062 = w2456 & w2474;
assign w51063 = w2717 & w493;
assign w51064 = w2431 & ~w2433;
assign w51065 = ~w2431 & w2433;
assign w51066 = w2555 & ~w2726;
assign w51067 = w2732 & ~w400;
assign w51068 = w1320 & w2765;
assign w51069 = w1320 & w39996;
assign w51070 = w2357 & w52338;
assign w51071 = w2769 & ~w39997;
assign w51072 = w2776 & w2771;
assign w51073 = ~w2732 & w400;
assign w51074 = w351 & ~w2785;
assign w51075 = w2006 & w2313;
assign w51076 = ~w2006 & w2313;
assign w51077 = w2516 & w2813;
assign w51078 = ~w2005 & w2818;
assign w51079 = ~w2825 & a[93];
assign w51080 = ~w51079 & ~w2312;
assign w51081 = w2825 & ~a[93];
assign w51082 = w2850 & w2786;
assign w51083 = w2849 & w2763;
assign w51084 = w2736 & w2860;
assign w51085 = w2854 & ~w2862;
assign w51086 = ~w2643 & w3;
assign w51087 = ~w44030 & w2883;
assign w51088 = ~w2631 & w2901;
assign w51089 = ~w2648 & w2902;
assign w51090 = ~w2619 & w2589;
assign w51091 = ~w2619 & w44031;
assign w51092 = (w2643 & w2909) | (w2643 & w51455) | (w2909 & w51455);
assign w51093 = (~w47041 & w2909) | (~w47041 & w51456) | (w2909 & w51456);
assign w51094 = ~w2680 & ~w2630;
assign w51095 = w2910 & ~w2912;
assign w51096 = ~w2900 & w2914;
assign w51097 = w2591 & ~w2601;
assign w51098 = ~w2918 & ~w2914;
assign w51099 = ~w2918 & ~w51096;
assign w51100 = w2589 & w2914;
assign w51101 = w2589 & w51096;
assign w51102 = w2627 & w2924;
assign w51103 = w2858 & ~w2665;
assign w51104 = w2680 & w2928;
assign w51105 = ~w2626 & w51457;
assign w51106 = (w2671 & w2930) | (w2671 & w51458) | (w2930 & w51458);
assign w51107 = ~w2931 & ~w44032;
assign w51108 = (~w80 & w2935) | (~w80 & w51459) | (w2935 & w51459);
assign w51109 = ~w2951 & w252;
assign w51110 = ~w2890 & w2922;
assign w51111 = w2962 & w2922;
assign w51112 = w2555 & w2378;
assign w51113 = ~w2555 & w2742;
assign w51114 = w47048 & w2776;
assign w51115 = ~w2757 & w2976;
assign w51116 = w2757 & ~w2976;
assign w51117 = w2680 & w47049;
assign w51118 = ~w2980 & w754;
assign w51119 = w2555 & w2333;
assign w51120 = ~w2555 & w2752;
assign w51121 = ~w47048 & ~w2776;
assign w51122 = ~w2985 & ~w2986;
assign w51123 = ~w47048 & ~w2757;
assign w51124 = ~w2995 & w2988;
assign w51125 = ~w2982 & w945;
assign w51126 = ~w2982 & ~w44034;
assign w51127 = w2980 & ~w754;
assign w51128 = ~w2849 & w2796;
assign w51129 = w2839 & ~w3003;
assign w51130 = w2897 & w3029;
assign w51131 = ~w2895 & w3030;
assign w51132 = w2841 & w1541;
assign w51133 = ~w2841 & ~w1541;
assign w51134 = w2866 & w2795;
assign w51135 = w2897 & w3044;
assign w51136 = ~w3053 & ~w3051;
assign w51137 = ~w2796 & ~w2771;
assign w51138 = ~w2796 & w2848;
assign w51139 = ~w2895 & w3045;
assign w51140 = ~w2555 & ~a[92];
assign w51141 = ~w2555 & w2828;
assign w51142 = w2648 & w3084;
assign w51143 = ~w2824 & a[93];
assign w51144 = w2676 & w3090;
assign w51145 = ~w2555 & w2285;
assign w51146 = w40003 & w2825;
assign w51147 = w2825 & ~w3098;
assign w51148 = ~w2858 & w3102;
assign w51149 = ~w2558 & w2677;
assign w51150 = ~w2824 & ~w3109;
assign w51151 = ~w2312 & w2677;
assign w51152 = w2858 & w2312;
assign w51153 = ~w2555 & w3119;
assign w51154 = w2555 & w3124;
assign w51155 = w2866 & ~w3125;
assign w51156 = a[90] & a[91];
assign w51157 = w2555 & ~w2824;
assign w51158 = w2866 & ~w3132;
assign w51159 = w2866 & w2558;
assign w51160 = w2866 & w44057;
assign w51161 = w3116 & ~w2006;
assign w51162 = w2708 & ~w3003;
assign w51163 = ~w2723 & ~w3175;
assign w51164 = ~w2723 & w3174;
assign w51165 = w2680 & w3177;
assign w51166 = w2720 & ~w3174;
assign w51167 = w2723 & ~w3174;
assign w51168 = w2866 & ~w2719;
assign w51169 = w3178 & ~w400;
assign w51170 = ~w3178 & w400;
assign w51171 = w2778 & ~w2707;
assign w51172 = w2897 & w3202;
assign w51173 = (~w2720 & w40021) | (~w2720 & w3175) | (w40021 & w3175);
assign w51174 = (~w2720 & w40021) | (~w2720 & ~w3174) | (w40021 & ~w3174);
assign w51175 = ~w3211 & w51173;
assign w51176 = ~w3211 & w51174;
assign w51177 = ~w2680 & ~w3244;
assign w51178 = ~a[89] & ~w3119;
assign w51179 = w2680 & ~a[90];
assign w51180 = ~w2680 & a[90];
assign w51181 = w2555 & ~w3257;
assign w51182 = w2680 & ~w2558;
assign w51183 = ~w2680 & w2558;
assign w51184 = ~w2555 & w3257;
assign w51185 = ~w2558 & w2285;
assign w51186 = w2558 & ~w2285;
assign w51187 = ~w3155 & w3265;
assign w51188 = ~w3155 & w40042;
assign w51189 = w3310 & w3028;
assign w51190 = ~w3162 & ~w3315;
assign w51191 = ~w3317 & ~w3319;
assign w51192 = w1738 & w1541;
assign w51193 = w3027 & ~w3116;
assign w51194 = w3027 & ~w47057;
assign w51195 = ~w3329 & ~w1738;
assign w51196 = w3330 & ~w3326;
assign w51197 = ~w3168 & ~w3028;
assign w51198 = w1541 & ~w3028;
assign w51199 = w1541 & w51197;
assign w51200 = ~w1541 & w3028;
assign w51201 = ~w1541 & ~w51197;
assign w51202 = w40049 & w2967;
assign w51203 = w40049 & w3240;
assign w51204 = (w3350 & w40050) | (w3350 & ~w2967) | (w40050 & ~w2967);
assign w51205 = (w3350 & w40050) | (w3350 & ~w3240) | (w40050 & ~w3240);
assign w51206 = ~w3339 & w3352;
assign w51207 = w3073 & ~w1120;
assign w51208 = w3359 & w3361;
assign w51209 = ~w3073 & ~w1120;
assign w51210 = ~w3359 & w3363;
assign w51211 = w3162 & w1738;
assign w51212 = ~w3162 & ~w1738;
assign w51213 = w3375 & ~w3372;
assign w51214 = w3375 & w40057;
assign w51215 = w2680 & w3044;
assign w51216 = w3168 & w3036;
assign w51217 = ~w3073 & w1120;
assign w51218 = w3073 & w1120;
assign w51219 = ~w3164 & ~w3054;
assign w51220 = w3455 & w3453;
assign w51221 = ~w3455 & ~w3453;
assign w51222 = w3500 & w3502;
assign w51223 = ~w3500 & w3504;
assign w51224 = w3190 & ~w2954;
assign w51225 = w80 & ~w2946;
assign w51226 = w2882 & ~w2630;
assign w51227 = ~w2882 & w2630;
assign w51228 = ~w3524 & w42;
assign w51229 = ~w2962 & ~w2876;
assign w51230 = ~w3536 & ~w3535;
assign w51231 = ~w3536 & w40096;
assign w51232 = ~w2921 & ~w42;
assign w51233 = w3533 & ~w3528;
assign w51234 = ~w3506 & ~w3545;
assign w51235 = w80 & w57;
assign w51236 = ~w2954 & ~w3221;
assign w51237 = w3219 & ~w3240;
assign w51238 = ~w3595 & ~w252;
assign w51239 = ~w3605 & ~w3598;
assign w51240 = w3589 & ~w3607;
assign w51241 = w3595 & w252;
assign w51242 = w351 & ~w3615;
assign w51243 = w3618 & ~w3546;
assign w51244 = w3445 & ~w493;
assign w51245 = ~w3445 & w493;
assign w51246 = ~w3446 & ~w3428;
assign w51247 = w3446 & ~w493;
assign w51248 = w3426 & w400;
assign w51249 = ~w3426 & w400;
assign w51250 = w3680 & ~w3647;
assign w51251 = w3399 & w51460;
assign w51252 = ~w3682 & ~w3681;
assign w51253 = w3683 & w493;
assign w51254 = ~w3683 & ~w493;
assign w51255 = w3359 & w3355;
assign w51256 = ~w3359 & ~w3355;
assign w51257 = w754 & ~w945;
assign w51258 = ~w3710 & ~w3711;
assign w51259 = ~w3713 & w3716;
assign w51260 = w3713 & ~w3716;
assign w51261 = w3733 & w3620;
assign w51262 = w3733 & ~w3464;
assign w51263 = ~w3701 & ~w3687;
assign w51264 = ~w3750 & ~w3240;
assign w51265 = a[87] & ~w3751;
assign w51266 = a[88] & ~w3240;
assign w51267 = w3774 & w3464;
assign w51268 = ~w3783 & ~w3240;
assign w51269 = ~w44090 & w2285;
assign w51270 = w3255 & ~w3240;
assign w51271 = ~w3027 & ~w3372;
assign w51272 = ~w3027 & w40057;
assign w51273 = w3264 & w2006;
assign w51274 = ~w3264 & ~w2006;
assign w51275 = ~w3872 & ~w3875;
assign w51276 = ~w3379 & w3340;
assign w51277 = ~w1320 & w3340;
assign w51278 = ~w1320 & w51276;
assign w51279 = w3866 & ~w3888;
assign w51280 = w3810 & w3889;
assign w51281 = ~w3668 & ~w3427;
assign w51282 = w3668 & w3427;
assign w51283 = w3687 & ~w3888;
assign w51284 = (~w3888 & w51283) | (~w3888 & w3701) | (w51283 & w3701);
assign w51285 = w3953 & ~w3519;
assign w51286 = ~w3617 & w3996;
assign w51287 = w3995 & w3464;
assign w51288 = w3993 & w3933;
assign w51289 = w3969 & w3630;
assign w51290 = w4062 & ~w57;
assign w51291 = w4062 & w4029;
assign w51292 = (~w3888 & w4024) | (~w3888 & w51543) | (w4024 & w51543);
assign w51293 = ~w4074 & ~w4075;
assign w51294 = ~w4074 & ~w3747;
assign w51295 = w4097 & ~w57;
assign w51296 = w4097 & w4029;
assign w51297 = ~w4103 & ~w4104;
assign w51298 = ~w4115 & w3925;
assign w51299 = w3981 & w3982;
assign w51300 = ~w3981 & ~w3982;
assign w51301 = w4134 & w50270;
assign w51302 = w4134 & ~w4116;
assign w51303 = w3745 & w3698;
assign w51304 = w3969 & ~w3686;
assign w51305 = ~w3673 & ~w351;
assign w51306 = w3673 & ~w351;
assign w51307 = w3673 & w351;
assign w51308 = ~w3673 & w351;
assign w51309 = ~w3741 & w754;
assign w51310 = ~w4213 & w3464;
assign w51311 = ~a[85] & ~w3749;
assign w51312 = a[86] & w3464;
assign w51313 = ~w4240 & w3464;
assign w51314 = w3969 & w4251;
assign w51315 = w2285 & ~w2807;
assign w51316 = w4029 & w4280;
assign w51317 = ~w4029 & w4282;
assign w51318 = ~w3805 & ~w2558;
assign w51319 = w3805 & w2558;
assign w51320 = w4029 & w4288;
assign w51321 = ~w4029 & w4290;
assign w51322 = w4029 & w3829;
assign w51323 = ~w4029 & w4296;
assign w51324 = w4029 & w4300;
assign w51325 = ~w4029 & w4302;
assign w51326 = w40180 & w1738;
assign w51327 = (w1738 & w40180) | (w1738 & ~w3810) | (w40180 & ~w3810);
assign w51328 = w3810 & w40181;
assign w51329 = w40183 | ~w1541;
assign w51330 = (~w1541 & w40183) | (~w1541 & ~w4055) | (w40183 & ~w4055);
assign w51331 = w4029 & ~w3878;
assign w51332 = ~w3969 & w1541;
assign w51333 = w4316 & w3933;
assign w51334 = w3895 & w4325;
assign w51335 = w4277 & w3821;
assign w51336 = ~w4344 & ~w4345;
assign w51337 = w4352 & w4356;
assign w51338 = ~w4352 & w4358;
assign w51339 = w4055 & w40190;
assign w51340 = w4029 & w4363;
assign w51341 = w40194 & w3896;
assign w51342 = (w3896 & w40194) | (w3896 & ~w3810) | (w40194 & ~w3810);
assign w51343 = w3852 & ~w4378;
assign w51344 = ~w3852 & w4378;
assign w51345 = ~w4342 & w4390;
assign w51346 = w4352 & w4397;
assign w51347 = ~w4352 & w4399;
assign w51348 = w4147 & ~w252;
assign w51349 = ~w4262 & w4273;
assign w51350 = w4250 & w4419;
assign w51351 = ~w4136 & w4447;
assign w51352 = w4055 & ~a[85];
assign w51353 = a[84] & a[85];
assign w51354 = w4225 & w2896;
assign w51355 = ~w4225 & ~w2896;
assign w51356 = w4055 & ~w4243;
assign w51357 = ~w4055 & ~w4246;
assign w51358 = w4029 & w3801;
assign w51359 = ~w4029 & ~w3801;
assign w51360 = w47100 & ~w1738;
assign w51361 = (~w1738 & w47100) | (~w1738 & w4294) | (w47100 & w4294);
assign w51362 = ~w4294 & w40204;
assign w51363 = ~w40204 & ~w4339;
assign w51364 = (~w4339 & w51363) | (~w4339 & w4294) | (w51363 & w4294);
assign w51365 = ~w4320 & w4321;
assign w51366 = w4320 & ~w4321;
assign w51367 = ~w4549 & ~w1120;
assign w51368 = w4029 & w3821;
assign w51369 = ~w4029 & ~w3821;
assign w51370 = ~w4352 & ~w4355;
assign w51371 = w4352 & w4355;
assign w51372 = w612 & w4638;
assign w51373 = w612 & w47105;
assign w51374 = w4640 & ~w4638;
assign w51375 = w4640 & ~w47105;
assign w51376 = ~w4351 & ~w4625;
assign w51377 = ~w4351 & w40207;
assign w51378 = ~w3320 & w2967;
assign w51379 = ~w3320 & w3240;
assign w51380 = w3161 & w1541;
assign w51381 = w3969 & w4217;
assign w51382 = w4222 & w4226;
assign w51383 = w4182 & w4717;
assign w51384 = ~w4649 & w4729;
assign w51385 = ~w1507 & w1554;
assign w51386 = ~w1507 & ~w1555;
assign w51387 = ~w1507 & w1590;
assign w51388 = ~w1507 & w1602;
assign w51389 = w2517 & w2772;
assign w51390 = ~w3 & w4073;
assign w51391 = w4344 & w3888;
assign w51392 = ~w1155 & ~w1212;
assign w51393 = w2099 & ~w2035;
assign w51394 = ~w42 & w2578;
assign w51395 = ~w42 & ~w44005;
assign w51396 = w3162 & w3234;
assign w51397 = w3305 & ~w3369;
assign w51398 = w44094 & w1738;
assign w51399 = ~w3662 & ~w3920;
assign w51400 = ~w3737 & w43355;
assign w51401 = ~w3737 & w43356;
assign w51402 = ~w1724 & ~w3;
assign w51403 = ~w1724 & w3;
assign w51404 = w1724 & w1762;
assign w51405 = ~w1724 & w1764;
assign w51406 = w1724 & w1776;
assign w51407 = ~w1724 & w1778;
assign w51408 = w1724 & w1782;
assign w51409 = ~w1724 & w1784;
assign w51410 = w1724 & w1792;
assign w51411 = w1724 & ~w1770;
assign w51412 = ~w1724 & w1775;
assign w51413 = w1724 & w1812;
assign w51414 = ~w1724 & w1814;
assign w51415 = w1724 & w1931;
assign w51416 = ~w1724 & w1934;
assign w51417 = w1724 & w1940;
assign w51418 = ~w1724 & w1943;
assign w51419 = ~w4050 & w4269;
assign w51420 = w4050 & w4271;
assign w51421 = ~w4050 & w4279;
assign w51422 = ~w4050 & w4287;
assign w51423 = w4050 & w3901;
assign w51424 = w4050 & ~w3901;
assign w51425 = ~w1724 & w1877;
assign w51426 = w1724 & w1879;
assign w51427 = ~w1724 & w1892;
assign w51428 = w1724 & w1894;
assign w51429 = ~w754 & ~w46409;
assign w51430 = ~w754 & ~w46410;
assign w51431 = w1621 & ~w1599;
assign w51432 = w2960 & w80;
assign w51433 = w2960 & w47038;
assign w51434 = w2890 & w2954;
assign w51435 = ~w3657 & ~w3658;
assign w51436 = w3657 & w3658;
assign w51437 = w4014 & ~w57;
assign w51438 = w4284 & ~w1738;
assign w51439 = ~w3969 & ~w4003;
assign w51440 = ~w3969 & w400;
assign w51441 = ~w3969 & w945;
assign w51442 = w3688 & w3694;
assign w51443 = ~w3688 & w3696;
assign w51444 = w945 & w4029;
assign w51445 = w945 & w48613;
assign w51446 = ~w400 & w4029;
assign w51447 = w4387 & w945;
assign w51448 = w3237 & w3246;
assign w51449 = w3965 & w3506;
assign w51450 = w1516 & ~w50917;
assign w51451 = w1516 & w1498;
assign w51452 = w1629 & ~w43942;
assign w51453 = w1629 & ~w1508;
assign w51454 = ~w1685 & ~w80;
assign w51455 = w2907 & w2643;
assign w51456 = w2907 & ~w47041;
assign w51457 = ~w2611 & w252;
assign w51458 = ~w2665 & w2671;
assign w51459 = w57 & ~w80;
assign w51460 = w3400 & w3680;
assign w51461 = w39840 & w1590;
assign w51462 = (w1590 & w39840) | (w1590 & w1476) | (w39840 & w1476);
assign w51463 = ~w2005 & w2229;
assign w51464 = ~w2005 & w2275;
assign w51465 = w42 & ~w51093;
assign w51466 = w42 & ~w51092;
assign w51467 = w3418 & w3014;
assign w51468 = ~w3418 & w3429;
assign w51469 = w3418 & ~w3429;
assign w51470 = w3287 & ~w50265;
assign w51471 = w3287 & ~w50264;
assign w51472 = ~w3287 & w50265;
assign w51473 = ~w3287 & w50264;
assign w51474 = ~w3830 & ~w3837;
assign w51475 = ~w3888 & ~w3662;
assign w51476 = ~w3969 & w3881;
assign w51477 = (w1120 & w43358) | (w1120 & w3901) | (w43358 & w3901);
assign w51478 = (w1120 & w43358) | (w1120 & w40193) | (w43358 & w40193);
assign w51479 = ~w50950 & w1549;
assign w51480 = w547 & a[110];
assign w51481 = ~w983 & ~w1232;
assign w51482 = (~w1187 & w50915) | (~w1187 & w1203) | (w50915 & w1203);
assign w51483 = (~w1187 & w50915) | (~w1187 & w46995) | (w50915 & w46995);
assign w51484 = ~w1492 & ~w1707;
assign w51485 = ~w1772 & ~w1526;
assign w51486 = ~w1594 & w754;
assign w51487 = w1972 & w1973;
assign w51488 = w1993 & w52339;
assign w51489 = w1993 & w52340;
assign w51490 = w2005 & ~w1738;
assign w51491 = ~w2591 & w2594;
assign w51492 = ~w42 & ~w51100;
assign w51493 = ~w42 & ~w51101;
assign w51494 = ~w2680 & ~w2970;
assign w51495 = w2897 & w2991;
assign w51496 = ~w2895 & w2992;
assign w51497 = ~w44006 & w3089;
assign w51498 = w2680 & w3215;
assign w51499 = w2680 & w3244;
assign w51500 = w3162 & w3168;
assign w51501 = w40082 | ~w3235;
assign w51502 = (~w3235 & w40082) | (~w3235 & w3418) | (w40082 & w3418);
assign w51503 = (~w3383 & w47081) | (~w3383 & ~w3620) | (w47081 & ~w3620);
assign w51504 = (~w3383 & w47081) | (~w3383 & w3464) | (w47081 & w3464);
assign w51505 = w47082 & w3620;
assign w51506 = w47082 & ~w3464;
assign w51507 = ~w3662 & ~w4022;
assign w51508 = ~w3698 & ~w493;
assign w51509 = w3698 & ~w493;
assign w51510 = w4222 & ~w4223;
assign w51511 = w4393 & ~w4351;
assign w51512 = w4418 & w4666;
assign w51513 = ~w4409 & ~w4182;
assign w51514 = w4692 & ~w4701;
assign w51515 = w4413 & w4102;
assign w51516 = ~w4114 & w4414;
assign w51517 = ~w42 & w4136;
assign w51518 = w4418 & ~w4091;
assign w51519 = ~w4772 & ~w4773;
assign w51520 = ~w40216 & w4780;
assign w51521 = w4418 & ~w4785;
assign w51522 = w4418 & w40220;
assign w51523 = ~w4822 & ~w4821;
assign w51524 = w4603 & w4839;
assign w51525 = ~w4603 & ~w4839;
assign w51526 = ~w1320 & w1541;
assign w51527 = ~w4610 & w4869;
assign w51528 = w4793 & ~w2558;
assign w51529 = ~w4497 & w4503;
assign w51530 = ~w4484 & ~w4496;
assign w51531 = w4466 & ~w4468;
assign w51532 = w4450 & ~w3646;
assign w51533 = ~w4450 & w3646;
assign w51534 = ~w4793 & ~w4934;
assign w51535 = w4465 & w3242;
assign w51536 = ~w4465 & w3242;
assign w51537 = ~w4418 & ~a[82];
assign w51538 = w3477 & w2967;
assign w51539 = w3477 & w3240;
assign w51540 = ~w3489 & ~w351;
assign w51541 = w3489 & w351;
assign w51542 = w3409 & ~w3934;
assign w51543 = w4022 & ~w3888;
assign w51544 = w1971 & w52339;
assign w51545 = w1971 & w52340;
assign w51546 = ~w3489 & w252;
assign w51547 = w3489 & ~w351;
assign w51548 = w4793 & w4956;
assign w51549 = ~w4418 & ~w4972;
assign w51550 = w4418 & w4972;
assign w51551 = w4793 & w40234;
assign w51552 = ~w4793 & w4979;
assign w51553 = ~w4418 & w4989;
assign w51554 = w4793 & ~w4990;
assign w51555 = w4418 & ~w4989;
assign w51556 = w4793 & w4993;
assign w51557 = w4793 & w4430;
assign w51558 = ~w4833 & w5012;
assign w51559 = a[82] & w4434;
assign w51560 = ~w4833 & w5025;
assign w51561 = ~w4465 & ~w3242;
assign w51562 = w4465 & ~w3242;
assign w51563 = w4793 & ~w4662;
assign w51564 = w4793 & ~w4685;
assign w51565 = w4549 & ~w945;
assign w51566 = ~w4549 & ~w945;
assign w51567 = w4793 & w5097;
assign w51568 = ~w4549 & w945;
assign w51569 = w4549 & w945;
assign w51570 = w4793 & w5107;
assign w51571 = ~w4558 & ~w4559;
assign w51572 = w4558 & w4559;
assign w51573 = w4882 & w4518;
assign w51574 = w4882 & ~w4605;
assign w51575 = w4669 & ~w4724;
assign w51576 = ~w4709 & ~w351;
assign w51577 = w4709 & w351;
assign w51578 = w400 & ~w5194;
assign w51579 = ~w4669 & ~w4637;
assign w51580 = ~w5193 & ~w5198;
assign w51581 = ~w4823 & ~w42;
assign w51582 = w4823 & ~w42;
assign w51583 = w4418 & w252;
assign w51584 = ~w5253 & w4794;
assign w51585 = w5253 & ~w4794;
assign w51586 = ~w5193 & ~w5194;
assign w51587 = ~w5214 & ~w5168;
assign w51588 = ~w5273 & ~w5274;
assign w51589 = w5344 & w4430;
assign w51590 = ~w4418 & a[78];
assign w51591 = ~w5344 & ~w4430;
assign w51592 = w4430 & ~w4988;
assign w51593 = ~w47127 & ~w5001;
assign w51594 = w44169 & ~w5380;
assign w51595 = ~w4987 & ~w5404;
assign w51596 = w4987 & w5404;
assign w51597 = w4913 & w4931;
assign w51598 = ~w44176 & ~w5424;
assign w51599 = ~w5432 & ~w5433;
assign w51600 = ~w5434 & ~w2285;
assign w51601 = ~w4892 & ~w4898;
assign w51602 = w4892 & w4898;
assign w51603 = ~w5442 & w5441;
assign w51604 = w5442 & ~w5441;
assign w51605 = ~w5329 & w5448;
assign w51606 = ~w5329 & w5459;
assign w51607 = ~w40270 & w5466;
assign w51608 = w5157 & w4868;
assign w51609 = ~w4987 & w5045;
assign w51610 = w4920 & w4495;
assign w51611 = ~w4920 & ~w4495;
assign w51612 = ~w44189 & w5289;
assign w51613 = ~w5128 & w5290;
assign w51614 = w4876 & w5290;
assign w51615 = ~w5048 & w5553;
assign w51616 = w5329 & ~w5559;
assign w51617 = ~w5329 & ~w5555;
assign w51618 = w4913 & w2285;
assign w51619 = ~w4913 & w2285;
assign w51620 = w5082 & w5078;
assign w51621 = ~w5062 & ~w493;
assign w51622 = ~w5608 & ~w5598;
assign w51623 = ~w5612 & ~w5613;
assign w51624 = ~w5329 & ~w5611;
assign w51625 = w5329 & w351;
assign w51626 = ~w5271 & ~w252;
assign w51627 = w5653 & w5655;
assign w51628 = w5271 & ~w252;
assign w51629 = ~w5653 & w5657;
assign w51630 = ~w5676 & w5659;
assign w51631 = ~w5692 & w5266;
assign w51632 = w5329 & w5260;
assign w51633 = ~w5693 & ~w5694;
assign w51634 = w5693 & w5694;
assign w51635 = w57 & ~w5181;
assign w51636 = w57 & w40280;
assign w51637 = ~w5702 & ~w5701;
assign w51638 = w5676 & ~w5700;
assign w51639 = w5294 & w5707;
assign w51640 = ~w5294 & ~w5707;
assign w51641 = w5329 & ~w5713;
assign w51642 = w5710 & w5715;
assign w51643 = w5695 & ~w3;
assign w51644 = w5271 & w252;
assign w51645 = ~w5271 & w252;
assign w51646 = ~w5300 & w5246;
assign w51647 = w5738 & w5246;
assign w51648 = w5738 & w51646;
assign w51649 = w5710 & ~w5714;
assign w51650 = ~w42 & ~w5740;
assign w51651 = w5718 & ~w5640;
assign w51652 = ~w5771 & w5646;
assign w51653 = w5609 & ~w400;
assign w51654 = ~w5609 & ~w400;
assign w51655 = ~w5609 & w400;
assign w51656 = w5609 & w400;
assign w51657 = ~w5835 & w5834;
assign w51658 = w5744 & w5839;
assign w51659 = ~w5836 & ~w5837;
assign w51660 = w5844 & ~w5843;
assign w51661 = w5857 & ~w3242;
assign w51662 = ~w5401 & ~w5865;
assign w51663 = w5401 & w5865;
assign w51664 = ~w5744 & w5871;
assign w51665 = w5718 & w5875;
assign w51666 = w5384 & w3646;
assign w51667 = ~w5876 & w5892;
assign w51668 = ~w5895 & ~w5893;
assign w51669 = w3646 & ~w5420;
assign w51670 = ~w5744 & w5912;
assign w51671 = w5898 & ~w5419;
assign w51672 = w5437 & w5586;
assign w51673 = ~w5422 & w5928;
assign w51674 = w5329 & w5440;
assign w51675 = ~w5329 & ~w5445;
assign w51676 = w5451 & ~w5464;
assign w51677 = ~w5329 & w5978;
assign w51678 = ~w51677 & ~w5980;
assign w51679 = w5718 & ~w5981;
assign w51680 = w5329 & ~w5978;
assign w51681 = ~w5329 & ~a[78];
assign w51682 = w5329 & a[78];
assign w51683 = w5718 & w6006;
assign w51684 = ~w51681 & a[79];
assign w51685 = w51681 & ~a[79];
assign w51686 = w5329 & w4838;
assign w51687 = w6024 & w51686;
assign w51688 = w5744 & ~w6021;
assign w51689 = ~w5744 & w6030;
assign w51690 = w5718 & w6039;
assign w51691 = w5874 & ~w6053;
assign w51692 = w6078 & ~w5529;
assign w51693 = w6078 & w40320;
assign w51694 = w2896 & ~w2558;
assign w51695 = ~w5744 & w5955;
assign w51696 = w5744 & w6089;
assign w51697 = w6083 & ~w6091;
assign w51698 = w5929 & w2006;
assign w51699 = ~w5744 & w6094;
assign w51700 = w6115 & ~w5659;
assign w51701 = w6115 & ~w40363;
assign w51702 = w5744 & w6120;
assign w51703 = ~w6119 & ~w6117;
assign w51704 = ~w5703 & ~w5689;
assign w51705 = w5744 & ~w80;
assign w51706 = w6127 & w6129;
assign w51707 = ~w6127 & w6131;
assign w51708 = ~w5717 & ~w5719;
assign w51709 = ~w5717 & ~w47132;
assign w51710 = ~w5321 & w5246;
assign w51711 = ~w5321 & w51646;
assign w51712 = w5321 & w5318;
assign w51713 = ~w6138 & ~w5742;
assign w51714 = w5676 & ~w6149;
assign w51715 = w6150 & ~w5691;
assign w51716 = w6150 & ~w40367;
assign w51717 = w5744 & ~w3;
assign w51718 = w5676 & ~w3;
assign w51719 = ~w5743 & ~w47133;
assign w51720 = ~w5743 & ~w47134;
assign w51721 = w5699 & w42;
assign w51722 = w6152 & w6158;
assign w51723 = w6127 & w6124;
assign w51724 = ~w6127 & ~w6124;
assign w51725 = w5513 & ~w754;
assign w51726 = w5544 & w5546;
assign w51727 = ~w5513 & ~w754;
assign w51728 = ~w5513 & w754;
assign w51729 = w5513 & w754;
assign w51730 = w6121 & w80;
assign w51731 = w6092 & w5897;
assign w51732 = w6099 & ~w5963;
assign w51733 = w6108 & w6268;
assign w51734 = w6108 & ~w6267;
assign w51735 = ~w6248 & ~w42;
assign w51736 = ~w6163 & ~w42;
assign w51737 = w5744 & ~w6320;
assign w51738 = w5854 & w6324;
assign w51739 = ~w5744 & w6320;
assign w51740 = ~w6343 & w6347;
assign w51741 = ~w5744 & ~a[76];
assign w51742 = w5744 & a[76];
assign w51743 = w5744 & ~w6362;
assign w51744 = ~w5744 & w6362;
assign w51745 = ~a[77] & ~w4838;
assign w51746 = ~w6385 & ~w6386;
assign w51747 = ~w6387 & w4838;
assign w51748 = ~w6059 & w6480;
assign w51749 = ~w6262 & w6505;
assign w51750 = ~w5947 & w1541;
assign w51751 = w5947 & w1541;
assign w51752 = w5947 & ~w1541;
assign w51753 = ~w5947 & ~w1541;
assign w51754 = ~w6569 & w945;
assign w51755 = ~w6571 & ~w6573;
assign w51756 = ~w6586 & ~w6584;
assign w51757 = w6593 & ~w6605;
assign w51758 = ~w5833 & w6610;
assign w51759 = w5833 & ~w6610;
assign w51760 = ~w6114 & ~w6614;
assign w51761 = ~w5845 & ~w5848;
assign w51762 = w5845 & w5848;
assign w51763 = ~w5817 & w6625;
assign w51764 = w6061 & ~w6627;
assign w51765 = ~w5833 & w5853;
assign w51766 = ~w5817 & ~w351;
assign w51767 = w6200 & w6683;
assign w51768 = ~w6200 & ~w6683;
assign w51769 = w6061 & w6690;
assign w51770 = w5744 & w945;
assign w51771 = ~w5744 & w6185;
assign w51772 = w6656 & w80;
assign w51773 = w6805 & w6807;
assign w51774 = ~w44258 & w6814;
assign w51775 = w6307 & a[73];
assign w51776 = w6307 & w6831;
assign w51777 = ~w5329 & ~a[75];
assign w51778 = ~w5329 & a[75];
assign w51779 = ~w6346 & ~w4838;
assign w51780 = w6346 & w4838;
assign w51781 = ~w6307 & ~w6877;
assign w51782 = ~w6387 & w4430;
assign w51783 = w6387 & w4430;
assign w51784 = w6425 & w3646;
assign w51785 = w6421 & w3646;
assign w51786 = w6392 & ~w6916;
assign w51787 = w6359 & ~w6391;
assign w51788 = ~w6421 & ~w3646;
assign w51789 = w6425 & ~w3646;
assign w51790 = w6946 & w6382;
assign w51791 = ~w6425 & ~w3646;
assign w51792 = w6951 & ~w6952;
assign w51793 = ~w6953 & w4056;
assign w51794 = w6435 & w6973;
assign w51795 = ~w6435 & ~w6973;
assign w51796 = ~w6979 & w6318;
assign w51797 = ~w6979 & w40434;
assign w51798 = w6461 & w5933;
assign w51799 = ~w6461 & ~w5933;
assign w51800 = w6744 & ~w945;
assign w51801 = ~w6744 & ~w945;
assign w51802 = ~w7119 & ~w7117;
assign w51803 = ~w6644 & w6735;
assign w51804 = w6307 & ~w6622;
assign w51805 = w7155 & ~w50285;
assign w51806 = w7155 & ~w7153;
assign w51807 = w7159 & ~w80;
assign w51808 = ~w6713 & ~w351;
assign w51809 = ~w51808 & ~w6715;
assign w51810 = w6735 & ~w6715;
assign w51811 = w6713 & w351;
assign w51812 = w7162 & w7174;
assign w51813 = ~w7162 & w7176;
assign w51814 = ~w44289 & w7187;
assign w51815 = w7191 & ~w7188;
assign w51816 = w7170 & w7208;
assign w51817 = ~w6309 & w80;
assign w51818 = ~w6656 & ~w3;
assign w51819 = ~w6307 & w7224;
assign w51820 = ~w6307 & w80;
assign w51821 = w6656 & ~w3;
assign w51822 = ~w7243 & w6735;
assign w51823 = w6305 & ~w3;
assign w51824 = ~w6281 & ~w42;
assign w51825 = (~w7260 & w40464) | (~w7260 & ~w6316) | (w40464 & ~w6316);
assign w51826 = (~w7260 & w40464) | (~w7260 & w40462) | (w40464 & w40462);
assign w51827 = w7132 & ~w493;
assign w51828 = w6735 & ~w7296;
assign w51829 = ~w7297 & ~w7298;
assign w51830 = w7299 & w400;
assign w51831 = w6774 & ~w6777;
assign w51832 = ~w6774 & w6777;
assign w51833 = w6280 & w6318;
assign w51834 = w6280 & w40434;
assign w51835 = ~w7007 & w1120;
assign w51836 = ~w7007 & ~w1120;
assign w51837 = w7111 & w754;
assign w51838 = ~w7111 & ~w754;
assign w51839 = ~w40486 & ~w7282;
assign w51840 = w7268 & w7430;
assign w51841 = w7429 & ~w7430;
assign w51842 = ~w754 & ~w47198;
assign w51843 = ~w754 & ~w47197;
assign w51844 = w7046 & w6318;
assign w51845 = w7046 & w40434;
assign w51846 = ~w7007 & w1320;
assign w51847 = ~w6264 & w6318;
assign w51848 = ~w6264 & w40434;
assign w51849 = a[70] & a[73];
assign w51850 = ~a[70] & ~a[73];
assign w51851 = ~w7565 & w7569;
assign w51852 = ~a[72] & ~w6828;
assign w51853 = w7563 & w7573;
assign w51854 = w7574 & ~w5745;
assign w51855 = a[70] & a[71];
assign w51856 = ~w6264 & w7577;
assign w51857 = w7563 & ~w7578;
assign w51858 = ~w7574 & w5745;
assign w51859 = w7268 & w7601;
assign w51860 = w6837 & w5330;
assign w51861 = ~w6837 & ~w5330;
assign w51862 = w7268 & ~w7625;
assign w51863 = w7268 & w40499;
assign w51864 = w40500 & w7630;
assign w51865 = (w7630 & w40500) | (w7630 & ~w7268) | (w40500 & ~w7268);
assign w51866 = w7268 & w7640;
assign w51867 = w7268 & w40504;
assign w51868 = w40505 & w7652;
assign w51869 = (w7652 & w40505) | (w7652 & ~w7268) | (w40505 & ~w7268);
assign w51870 = w2896 & w7063;
assign w51871 = w2896 & w49542;
assign w51872 = w2896 & ~w7701;
assign w51873 = w6972 & w7063;
assign w51874 = w6972 & w49542;
assign w51875 = ~w7469 & ~w7704;
assign w51876 = w7705 & ~w2558;
assign w51877 = ~w7703 & w7055;
assign w51878 = w7743 & ~w3242;
assign w51879 = ~w7743 & ~w3242;
assign w51880 = ~w7703 & w7766;
assign w51881 = ~w7437 & w400;
assign w51882 = w7268 & ~w7789;
assign w51883 = ~w7192 & w351;
assign w51884 = w493 & w6318;
assign w51885 = w493 & w40434;
assign w51886 = ~w7824 & w7296;
assign w51887 = w7824 & ~w7296;
assign w51888 = ~w7195 & ~w7301;
assign w51889 = w7217 & ~w7220;
assign w51890 = ~w6281 & w6301;
assign w51891 = ~w7878 & ~w42;
assign w51892 = ~w7881 & w47210;
assign w51893 = ~w7881 & w47211;
assign w51894 = w7308 & w7216;
assign w51895 = ~w7162 & ~w7173;
assign w51896 = w7162 & w7173;
assign w51897 = w7343 & w7009;
assign w51898 = ~w7343 & ~w7009;
assign w51899 = w7467 & ~w1320;
assign w51900 = ~w7427 & ~w7413;
assign w51901 = ~w7326 & w754;
assign w51902 = w7326 & w754;
assign w51903 = w7326 & ~w754;
assign w51904 = ~w7326 & ~w754;
assign w51905 = ~w234 & w252;
assign w51906 = ~w7437 & ~w351;
assign w51907 = w7450 & ~w7783;
assign w51908 = w7909 & ~w7915;
assign w51909 = w7839 & ~w8115;
assign w51910 = ~w7916 & w3;
assign w51911 = ~w7916 & ~w7920;
assign w51912 = ~w8128 & ~w7854;
assign w51913 = ~w8128 & w7854;
assign w51914 = w7872 & w49601;
assign w51915 = w7872 & w49602;
assign w51916 = ~w42 & w7908;
assign w51917 = w8121 & ~w8120;
assign w51918 = w8121 & ~w44359;
assign w51919 = w8198 & w7139;
assign w51920 = a[71] & ~w8196;
assign w51921 = w8195 & w6264;
assign w51922 = ~w44345 & w8199;
assign w51923 = w8207 & w7564;
assign w51924 = ~w7887 & w8209;
assign w51925 = ~w8212 & ~w8211;
assign w51926 = w8218 & w7139;
assign w51927 = w8220 & w7139;
assign w51928 = ~w6769 & w7139;
assign w51929 = a[68] & w6318;
assign w51930 = a[68] & w40434;
assign w51931 = w8266 & w8267;
assign w51932 = ~w8271 & ~w8272;
assign w51933 = w8195 & ~w8197;
assign w51934 = w8288 & a[72];
assign w51935 = ~w8288 & ~a[72];
assign w51936 = ~w7668 & w7694;
assign w51937 = ~w7636 & w7657;
assign w51938 = ~w7641 & w6873;
assign w51939 = w7641 & ~w6873;
assign w51940 = w8348 & ~w8344;
assign w51941 = w8348 & ~w40611;
assign w51942 = w8350 & w8344;
assign w51943 = w8350 & w40611;
assign w51944 = w7622 & ~w4838;
assign w51945 = ~w7622 & w4838;
assign w51946 = ~w7626 & w6895;
assign w51947 = w7626 & ~w6895;
assign w51948 = ~w7602 & w6845;
assign w51949 = w7602 & ~w6845;
assign w51950 = ~w2896 & w7713;
assign w51951 = ~w8413 & ~w8414;
assign w51952 = ~w7899 & ~w2558;
assign w51953 = w7909 & w8417;
assign w51954 = w7841 & w8418;
assign w51955 = w7708 & ~w2285;
assign w51956 = ~w7708 & ~w2285;
assign w51957 = w7708 & w2285;
assign w51958 = ~w7708 & w2285;
assign w51959 = ~w8406 & ~w3242;
assign w51960 = w8406 & w3242;
assign w51961 = w8452 & w7762;
assign w51962 = ~w8452 & ~w7762;
assign w51963 = ~w2896 & ~w7713;
assign w51964 = w3278 & ~w3277;
assign w51965 = ~w7502 & ~w8522;
assign w51966 = ~w7900 & w7522;
assign w51967 = w7522 & ~w7922;
assign w51968 = ~w8529 & w8531;
assign w51969 = w8322 & w3242;
assign w51970 = w51966 & w1541;
assign w51971 = w7841 & w8563;
assign w51972 = w7781 & w8564;
assign w51973 = ~w8576 & ~w8580;
assign w51974 = ~w8541 & w8581;
assign w51975 = ~w8576 & w8580;
assign w51976 = w8590 & w945;
assign w51977 = w8540 & ~w8602;
assign w51978 = w1120 & w8554;
assign w51979 = ~w44387 & ~w8619;
assign w51980 = w8390 & ~w8646;
assign w51981 = ~w8469 & w8479;
assign w51982 = w8459 & ~w44344;
assign w51983 = w8459 & w47215;
assign w51984 = w8455 & w2558;
assign w51985 = ~w8455 & w2558;
assign w51986 = ~w8189 & w8706;
assign w51987 = w8748 & ~w1738;
assign w51988 = ~w8680 & ~w8633;
assign w51989 = w8275 & w8337;
assign w51990 = ~w8359 & w8356;
assign w51991 = ~w8359 & w40612;
assign w51992 = w8275 & w8339;
assign w51993 = ~w8101 & w4056;
assign w51994 = w8365 & ~w8302;
assign w51995 = ~w8365 & ~w8401;
assign w51996 = ~w8841 & ~w8842;
assign w51997 = ~w3242 & w8842;
assign w51998 = ~w3242 & ~w51996;
assign w51999 = ~a[67] & ~w8218;
assign w52000 = w8884 & ~w44344;
assign w52001 = w8884 & w47215;
assign w52002 = ~a[68] & ~w44344;
assign w52003 = ~a[68] & w47215;
assign w52004 = ~w8911 & ~w44344;
assign w52005 = ~w8911 & w47215;
assign w52006 = w6769 & ~w6264;
assign w52007 = ~w8278 & ~w8940;
assign w52008 = ~w8765 & ~w8611;
assign w52009 = ~w7943 & ~w754;
assign w52010 = ~w7983 & w7445;
assign w52011 = w7983 & ~w7445;
assign w52012 = w8075 & w8153;
assign w52013 = ~w8189 & w8181;
assign w52014 = ~w8666 & ~w9020;
assign w52015 = w8113 & ~w8177;
assign w52016 = w9024 & ~w50298;
assign w52017 = w9024 & ~w50299;
assign w52018 = ~w8027 & ~w7971;
assign w52019 = ~w57 & ~w9046;
assign w52020 = ~w9077 & w8027;
assign w52021 = ~w8013 & w8027;
assign w52022 = ~w8074 & w8087;
assign w52023 = ~w40678 & w9116;
assign w52024 = w57 & ~w9046;
assign w52025 = w44427 & ~w80;
assign w52026 = (~w80 & w44427) | (~w80 & w40678) | (w44427 & w40678);
assign w52027 = ~w9119 & w9120;
assign w52028 = w9182 & w49601;
assign w52029 = w9182 & w49602;
assign w52030 = (w42 & w40688) | (w42 & ~w50298) | (w40688 & ~w50298);
assign w52031 = (w42 & w40688) | (w42 & ~w50299) | (w40688 & ~w50299);
assign w52032 = ~w8762 & w8981;
assign w52033 = w8762 & ~w9198;
assign w52034 = ~w9200 & ~w9199;
assign w52035 = ~w9197 & ~w8976;
assign w52036 = w9207 & w612;
assign w52037 = w8756 & ~w8675;
assign w52038 = ~w9226 & w8665;
assign w52039 = w40691 | w9252;
assign w52040 = (w9252 & w40691) | (w9252 & w8882) | (w40691 & w8882);
assign w52041 = ~w9255 & ~w9254;
assign w52042 = w9255 & ~w9252;
assign w52043 = ~w9175 & w9262;
assign w52044 = w9256 & w1541;
assign w52045 = ~w8882 & w8973;
assign w52046 = w40693 | w9229;
assign w52047 = (w9229 & w40693) | (w9229 & w8882) | (w40693 & w8882);
assign w52048 = ~w9225 & ~w9271;
assign w52049 = ~w9175 & w9278;
assign w52050 = w8756 & ~w9286;
assign w52051 = ~w8756 & w9286;
assign w52052 = w9272 & ~w1120;
assign w52053 = w40699 | ~w8747;
assign w52054 = (~w8747 & w40699) | (~w8747 & w8882) | (w40699 & w8882);
assign w52055 = w40700 | w8745;
assign w52056 = (w8745 & w40700) | (w8745 & w8882) | (w40700 & w8882);
assign w52057 = w40701 | w9339;
assign w52058 = (w9339 & w40701) | (w9339 & w8882) | (w40701 & w8882);
assign w52059 = ~w9340 & ~w9338;
assign w52060 = w8189 & w9351;
assign w52061 = ~w8189 & ~w9351;
assign w52062 = ~w9175 & w9357;
assign w52063 = ~w8189 & a[66];
assign w52064 = w8189 & ~a[66];
assign w52065 = ~w8189 & w7924;
assign w52066 = w8189 & ~w7924;
assign w52067 = w8935 & w9398;
assign w52068 = ~w8935 & ~w9398;
assign w52069 = ~w9028 & w9421;
assign w52070 = ~w8948 & ~w8957;
assign w52071 = ~w9443 & ~w8957;
assign w52072 = ~w9443 & w52070;
assign w52073 = w8947 & w9463;
assign w52074 = ~w8947 & ~w9463;
assign w52075 = w8957 & w9485;
assign w52076 = ~w9486 & w9480;
assign w52077 = w9486 & ~w9480;
assign w52078 = ~w8957 & ~w8867;
assign w52079 = ~w8828 & w8852;
assign w52080 = w8814 & w8860;
assign w52081 = ~w9526 & w40723;
assign w52082 = ~w9175 & w9532;
assign w52083 = ~w7705 & w2558;
assign w52084 = ~w8453 & ~w8456;
assign w52085 = ~w9175 & w9546;
assign w52086 = ~w9175 & w9627;
assign w52087 = ~w9207 & ~w612;
assign w52088 = ~w6767 & w6824;
assign w52089 = ~w7853 & w7886;
assign w52090 = ~w8077 & ~w7911;
assign w52091 = w8424 & ~w8420;
assign w52092 = w8424 & w40618;
assign w52093 = w8426 & w8420;
assign w52094 = w8426 & ~w40618;
assign w52095 = w8444 & w8420;
assign w52096 = w8444 & ~w40618;
assign w52097 = w8446 & ~w8420;
assign w52098 = w8446 & w40618;
assign w52099 = w5898 & w5907;
assign w52100 = ~w5898 & w5909;
assign w52101 = ~w6003 & ~w4430;
assign w52102 = w9079 & ~w44421;
assign w52103 = w9079 & w9078;
assign w52104 = ~w7086 & w7399;
assign w52105 = ~w48658 & ~w6248;
assign w52106 = ~w5855 & ~w6262;
assign w52107 = ~w6263 & w5759;
assign w52108 = w6263 & w6277;
assign w52109 = ~w6263 & w80;
assign w52110 = w6311 & w6310;
assign w52111 = ~w6311 & ~w6310;
assign w52112 = ~w6263 & w6451;
assign w52113 = ~w6453 & ~w2896;
assign w52114 = ~w6263 & w5842;
assign w52115 = ~w6263 & w6666;
assign w52116 = w6714 & w351;
assign w52117 = ~w6263 & w6731;
assign w52118 = ~w6609 & w40457;
assign w52119 = w40458 & w7224;
assign w52120 = (w7224 & w40458) | (w7224 & w6609) | (w40458 & w6609);
assign w52121 = ~w6989 & w43393;
assign w52122 = ~w1738 & ~w48709;
assign w52123 = ~w1738 & ~w48710;
assign w52124 = w7152 & ~w7156;
assign w52125 = ~w7158 & w80;
assign w52126 = ~w48711 & w1541;
assign w52127 = w48711 & ~w1541;
assign w52128 = (~a[123] & ~w39652) | (~a[123] & ~w75) | (~w39652 & ~w75);
assign w52129 = (w456 & ~w39701) | (w456 & ~w424) | (~w39701 & ~w424);
assign w52130 = (w693 & ~w80) | (w693 & w50777) | (~w80 & w50777);
assign w52131 = (w552 & ~w603) | (w552 & ~w50666) | (~w603 & ~w50666);
assign w52132 = (w716 & ~w3) | (w716 & w50840) | (~w3 & w50840);
assign w52133 = (w720 & w39750) | (w720 & ~w758) | (w39750 & ~w758);
assign w52134 = (w716 & w743) | (w716 & w50847) | (w743 & w50847);
assign w52135 = (w905 & ~w50859) | (w905 & ~w904) | (~w50859 & ~w904);
assign w52136 = (~w942 & w57) | (~w942 & w50874) | (w57 & w50874);
assign w52137 = (w1114 & ~w50253) | (w1114 & ~w1179) | (~w50253 & ~w1179);
assign w52138 = (~w1203 & ~w46995) | (~w1203 & ~w1328) | (~w46995 & ~w1328);
assign w52139 = (w50258 & w50259) | (w50258 & ~w1395) | (w50259 & ~w1395);
assign w52140 = (w1483 & w39863) | (w1483 & ~w1465) | (w39863 & ~w1465);
assign w52141 = (~w1514 & ~w50955) | (~w1514 & ~w1465) | (~w50955 & ~w1465);
assign w52142 = (w1528 & ~a[100]) | (w1528 & w50970) | (~a[100] & w50970);
assign w52143 = (w1528 & ~w1772) | (w1528 & w51485) | (~w1772 & w51485);
assign w52144 = (w1528 & w1805) | (w1528 & w50973) | (w1805 & w50973);
assign w52145 = (~w47011 & ~w1595) | (~w47011 & ~w47012) | (~w1595 & ~w47012);
assign w52146 = (w1757 & ~w47018) | (w1757 & ~w1954) | (~w47018 & ~w1954);
assign w52147 = ~w2103 & w52341;
assign w52148 = (~w2535 & ~w44004) | (~w2535 & ~w2517) | (~w44004 & ~w2517);
assign w52149 = (w2548 & ~w2517) | (w2548 & ~w2537) | (~w2517 & ~w2537);
assign w52150 = (w3002 & w2720) | (w3002 & w51166) | (w2720 & w51166);
assign w52151 = (w3002 & w2723) | (w3002 & w51167) | (w2723 & w51167);
assign w52152 = (~w3265 & ~w40042) | (~w3265 & ~w3241) | (~w40042 & ~w3241);
assign w52153 = (~w1541 & ~w51192) | (~w1541 & ~w3161) | (~w51192 & ~w3161);
assign w52154 = (w3372 & ~w40057) | (w3372 & ~w3241) | (~w40057 & ~w3241);
assign w52155 = (~w3049 & w3168) | (~w3049 & w51216) | (w3168 & w51216);
assign w52156 = (w3055 & ~w3164) | (w3055 & w51219) | (~w3164 & w51219);
assign w52157 = w3536 & ~w3494;
assign w52158 = (w3236 & ~w2954) | (w3236 & w51236) | (~w2954 & w51236);
assign w52159 = (w3224 & w3221) | (w3224 & ~w40106) | (w3221 & ~w40106);
assign w52160 = (w3223 & w3219) | (w3223 & w51237) | (w3219 & w51237);
assign w52161 = (~w3647 & w3401) | (~w3647 & ~w40118) | (w3401 & ~w40118);
assign w52162 = (w3223 & ~w3750) | (w3223 & w51264) | (~w3750 & w51264);
assign w52163 = (~w3754 & ~w40120) | (~w3754 & ~w3619) | (~w40120 & ~w3619);
assign w52164 = (w3223 & a[88]) | (w3223 & w51266) | (a[88] & w51266);
assign w52165 = (~w3644 & w3774) | (~w3644 & w51267) | (w3774 & w51267);
assign w52166 = (~w3771 & ~w40123) | (~w3771 & ~w3619) | (~w40123 & ~w3619);
assign w52167 = (w3223 & ~w3783) | (w3223 & w51268) | (~w3783 & w51268);
assign w52168 = (w3247 & ~w40125) | (w3247 & ~w3619) | (~w40125 & ~w3619);
assign w52169 = (w3223 & w3255) | (w3223 & w51270) | (w3255 & w51270);
assign w52170 = (~w3340 & ~w51276) | (~w3340 & ~w3309) | (~w51276 & ~w3309);
assign w52171 = (~w3644 & w3995) | (~w3644 & w51287) | (w3995 & w51287);
assign w52172 = (w3597 & ~w40144) | (w3597 & ~w3608) | (~w40144 & ~w3608);
assign w52173 = (~w4019 & ~w4115) | (~w4019 & w51298) | (~w4115 & w51298);
assign w52174 = (~w50270 & w4116) | (~w50270 & ~w50271) | (w4116 & ~w50271);
assign w52175 = (~w3644 & ~w4213) | (~w3644 & w51310) | (~w4213 & w51310);
assign w52176 = (~w3644 & a[86]) | (~w3644 & w51312) | (a[86] & w51312);
assign w52177 = (~w3644 & ~w4240) | (~w3644 & w51313) | (~w4240 & w51313);
assign w52178 = (~w3901 & ~w40193) | (~w3901 & ~w4080) | (~w40193 & ~w4080);
assign w52179 = (w4407 & ~w4432) | (w4407 & ~w44132) | (~w4432 & ~w44132);
assign w52180 = (~w47101 & ~w4295) | (~w47101 & ~w48630) | (~w4295 & ~w48630);
assign w52181 = w40205 & ~w4264;
assign w52182 = w4390 & ~w4343;
assign w52183 = (~w4112 & ~w40214) | (~w4112 & ~w4446) | (~w40214 & ~w4446);
assign w52184 = w40216 & ~w4446;
assign w52185 = (~w40222 & w4850) | (~w40222 & ~w4843) | (w4850 & ~w4843);
assign w52186 = (~w4746 & w5168) | (~w4746 & ~w40255) | (w5168 & ~w40255);
assign w52187 = (~w5175 & w5168) | (~w5175 & ~w40256) | (w5168 & ~w40256);
assign w52188 = (~w5213 & w5168) | (~w5213 & ~w40261) | (w5168 & ~w40261);
assign w52189 = (w4962 & w5217) | (w4962 & w49494) | (w5217 & w49494);
assign w52190 = (w4962 & ~w5214) | (w4962 & w51587) | (~w5214 & w51587);
assign w52191 = (~w4835 & ~w40267) | (~w4835 & ~w5225) | (~w40267 & ~w5225);
assign w52192 = (~w5354 & ~w47128) | (~w5354 & ~w5328) | (~w47128 & ~w5328);
assign w52193 = (~w5509 & ~w44190) | (~w5509 & ~w5328) | (~w44190 & ~w5328);
assign w52194 = (~w5615 & ~w44212) | (~w5615 & ~w5328) | (~w44212 & ~w5328);
assign w52195 = (~w5224 & ~w40274) | (~w5224 & ~w5293) | (~w40274 & ~w5293);
assign w52196 = (~w5967 & ~w5400) | (~w5967 & ~w40332) | (~w5400 & ~w40332);
assign w52197 = (~w47136 & w6285) | (~w47136 & ~w47137) | (w6285 & ~w47137);
assign w52198 = (~w1120 & w6593) | (~w1120 & w51757) | (w6593 & w51757);
assign w52199 = (w6674 & ~w6061) | (w6674 & ~w47143) | (~w6061 & ~w47143);
assign w52200 = (~w6197 & ~w6701) | (~w6197 & ~w40427) | (~w6701 & ~w40427);
assign w52201 = (~w47162 & w6910) | (~w47162 & ~w47163) | (w6910 & ~w47163);
assign w52202 = (w6592 & ~w44279) | (w6592 & ~w7107) | (~w44279 & ~w7107);
assign w52203 = (~w7252 & ~w40463) | (~w7252 & ~w6737) | (~w40463 & ~w6737);
assign w52204 = (~w7269 & ~w40484) | (~w7269 & ~w7068) | (~w40484 & ~w7068);
assign w52205 = (w47198 & w47197) | (w47198 & ~w40470) | (w47197 & ~w40470);
assign w52206 = (~w47210 & ~w47211) | (~w47210 & ~w7787) | (~w47211 & ~w7787);
assign w52207 = (w7955 & ~w7951) | (w7955 & ~w47218) | (~w7951 & ~w47218);
assign w52208 = (w7832 & ~w8079) | (w7832 & ~w40577) | (~w8079 & ~w40577);
assign w52209 = (~w49601 & ~w49602) | (~w49601 & ~w8103) | (~w49602 & ~w8103);
assign w52210 = (~w7304 & w8198) | (~w7304 & w51919) | (w8198 & w51919);
assign w52211 = (~w8209 & ~w51924) | (~w8209 & ~w8127) | (~w51924 & ~w8127);
assign w52212 = (~w7304 & w8218) | (~w7304 & w51926) | (w8218 & w51926);
assign w52213 = (~w7304 & w8220) | (~w7304 & w51927) | (w8220 & w51927);
assign w52214 = (~w8250 & ~w40600) | (~w8250 & ~w7782) | (~w40600 & ~w7782);
assign w52215 = (~w7304 & ~w6769) | (~w7304 & w51928) | (~w6769 & w51928);
assign w52216 = (~w8260 & ~w40602) | (~w8260 & ~w7782) | (~w40602 & ~w7782);
assign w52217 = (~w8270 & ~w40603) | (~w8270 & ~w7782) | (~w40603 & ~w7782);
assign w52218 = (~w8297 & ~w40605) | (~w8297 & ~w7782) | (~w40605 & ~w7782);
assign w52219 = (~w8344 & ~w40611) | (~w8344 & ~w7782) | (~w40611 & ~w7782);
assign w52220 = (w7914 & w7522) | (w7914 & w51967) | (w7522 & w51967);
assign w52221 = (w8512 & ~w40648) | (w8512 & ~w8615) | (~w40648 & ~w8615);
assign w52222 = (~w8583 & w1120) | (~w8583 & w51978) | (w1120 & w51978);
assign w52223 = (~w8356 & ~w40612) | (~w8356 & ~w7782) | (~w40612 & ~w7782);
assign w52224 = (~w8099 & ~w44414) | (~w8099 & ~w9013) | (~w44414 & ~w9013);
assign w52225 = (w50298 & w50299) | (w50298 & ~w9013) | (w50299 & ~w9013);
assign w52226 = ~w9119 & ~w9112;
assign w52227 = (~w8183 & ~w44415) | (~w8183 & ~w9013) | (~w44415 & ~w9013);
assign w52228 = (w8957 & ~w52070) | (w8957 & ~w8937) | (~w52070 & ~w8937);
assign w52229 = (~w9452 & ~w40716) | (~w9452 & ~w8937) | (~w40716 & ~w8937);
assign w52230 = (w9862 & w50229) | (w9862 & ~w10421) | (w50229 & ~w10421);
assign w52231 = (w10389 & ~w40892) | (w10389 & ~w10074) | (~w40892 & ~w10074);
assign w52232 = (w9850 & ~w40893) | (w9850 & ~w10396) | (~w40893 & ~w10396);
assign w52233 = (w11310 & ~w50302) | (w11310 & ~w11137) | (~w50302 & ~w11137);
assign w52234 = (w11346 & w40956) | (w11346 & ~w11221) | (w40956 & ~w11221);
assign w52235 = (w11148 & ~w11787) | (w11148 & ~w44540) | (~w11787 & ~w44540);
assign w52236 = (~w12249 & ~w41042) | (~w12249 & ~w12246) | (~w41042 & ~w12246);
assign w52237 = (~w12263 & ~w41047) | (~w12263 & ~w12246) | (~w41047 & ~w12246);
assign w52238 = (~w11358 & ~w41063) | (~w11358 & ~w12246) | (~w41063 & ~w12246);
assign w52239 = (~w12385 & w12076) | (~w12385 & ~w41068) | (w12076 & ~w41068);
assign w52240 = (~w12159 & ~w41121) | (~w12159 & ~w12833) | (~w41121 & ~w12833);
assign w52241 = (~w12598 & ~w12637) | (~w12598 & ~w44637) | (~w12637 & ~w44637);
assign w52242 = w13166 & ~w13160;
assign w52243 = (~w12527 & ~w41158) | (~w12527 & ~w12583) | (~w41158 & ~w12583);
assign w52244 = (~w13407 & w12696) | (~w13407 & ~w48756) | (w12696 & ~w48756);
assign w52245 = (~w13722 & ~w44808) | (~w13722 & ~w44809) | (~w44808 & ~w44809);
assign w52246 = (~w44896 & w41288) | (~w44896 & ~w44897) | (w41288 & ~w44897);
assign w52247 = (~w16704 & ~w15938) | (~w16704 & ~w41395) | (~w15938 & ~w41395);
assign w52248 = (~w21497 & ~w21256) | (~w21497 & ~w41807) | (~w21256 & ~w41807);
assign w52249 = (w21491 & ~w21256) | (w21491 & ~w41808) | (~w21256 & ~w41808);
assign w52250 = (w22294 & ~w41893) | (w22294 & ~w21800) | (~w41893 & ~w21800);
assign w52251 = (~w21237 & ~w41921) | (~w21237 & ~w21140) | (~w41921 & ~w21140);
assign w52252 = (~w22479 & w41976) | (~w22479 & ~w22416) | (w41976 & ~w22416);
assign w52253 = (w22118 & ~w42027) | (w22118 & ~w22745) | (~w42027 & ~w22745);
assign w52254 = (~w45403 & ~w45404) | (~w45403 & ~w24258) | (~w45404 & ~w24258);
assign w52255 = (w24557 & w25439) | (w24557 & w42154) | (w25439 & w42154);
assign w52256 = (w80 & ~w42200) | (w80 & ~w24901) | (~w42200 & ~w24901);
assign w52257 = (~w25312 & w42229) | (~w25312 & ~w25237) | (w42229 & ~w25237);
assign w52258 = (w25821 & w26051) | (w25821 & w45585) | (w26051 & w45585);
assign w52259 = (w26950 & w46625) | (w26950 & ~w26949) | (w46625 & ~w26949);
assign w52260 = (~w26750 & w26073) | (~w26750 & ~w42253) | (w26073 & ~w42253);
assign w52261 = (w42235 & ~w47756) | (w42235 & ~w47757) | (~w47756 & ~w47757);
assign w52262 = (~w27389 & ~w42286) | (~w27389 & ~w26517) | (~w42286 & ~w26517);
assign w52263 = (~w26622 & ~w42291) | (~w26622 & ~w26517) | (~w42291 & ~w26517);
assign w52264 = (~w26114 & ~w45643) | (~w26114 & ~w27654) | (~w45643 & ~w27654);
assign w52265 = (w26292 & w45646) | (w26292 & ~w26949) | (w45646 & ~w26949);
assign w52266 = (w27786 & ~w26827) | (w27786 & ~w47772) | (~w26827 & ~w47772);
assign w52267 = (~w27951 & ~w42333) | (~w27951 & ~w26885) | (~w42333 & ~w26885);
assign w52268 = (~w27639 & ~w27742) | (~w27639 & w50376) | (~w27742 & w50376);
assign w52269 = (w28696 & ~w42394) | (w28696 & ~w28694) | (~w42394 & ~w28694);
assign w52270 = (~w28783 & ~w42398) | (~w28783 & ~w27876) | (~w42398 & ~w27876);
assign w52271 = (~w28472 & ~w42436) | (~w28472 & ~w29353) | (~w42436 & ~w29353);
assign w52272 = (~w33798 & ~w46036) | (~w33798 & ~w33739) | (~w46036 & ~w33739);
assign w52273 = (~w33144 & w42713) | (~w33144 & ~w33084) | (w42713 & ~w33084);
assign w52274 = (~w34671 & ~w42826) | (~w34671 & ~w33557) | (~w42826 & ~w33557);
assign w52275 = ~w34750 & ~w34749;
assign w52276 = (w32964 & ~w42862) | (w32964 & ~w34787) | (~w42862 & ~w34787);
assign w52277 = (~w35029 & ~w48011) | (~w35029 & ~w34917) | (~w48011 & ~w34917);
assign w52278 = w49434 & ~w34168;
assign w52279 = (~w35652 & w49361) | (~w35652 & ~w35631) | (w49361 & ~w35631);
assign w52280 = (~w34850 & ~w46076) | (~w34850 & ~w35371) | (~w46076 & ~w35371);
assign w52281 = (~w35754 & ~w46082) | (~w35754 & ~w35631) | (~w46082 & ~w35631);
assign w52282 = (~w33820 & ~w46093) | (~w33820 & ~w34917) | (~w46093 & ~w34917);
assign w52283 = (~w36038 & ~w42980) | (~w36038 & ~w35993) | (~w42980 & ~w35993);
assign w52284 = (~w36075 & ~w42983) | (~w36075 & ~w35993) | (~w42983 & ~w35993);
assign w52285 = (~w36103 & ~w42985) | (~w36103 & ~w35993) | (~w42985 & ~w35993);
assign w52286 = (~w36123 & ~w42986) | (~w36123 & ~w35993) | (~w42986 & ~w35993);
assign w52287 = (~w36145 & ~w42989) | (~w36145 & ~w35993) | (~w42989 & ~w35993);
assign w52288 = (w36572 & ~w46180) | (w36572 & ~w46181) | (~w46180 & ~w46181);
assign w52289 = (w36572 & ~w46200) | (w36572 & ~w46201) | (~w46200 & ~w46201);
assign w52290 = (~w38328 & ~w43162) | (~w38328 & ~w38197) | (~w43162 & ~w38197);
assign w52291 = (w38403 & ~w43166) | (w38403 & ~w38336) | (~w43166 & ~w38336);
assign w52292 = (w38433 & ~w43167) | (w38433 & ~w38336) | (~w43167 & ~w38336);
assign w52293 = (~w38469 & ~w43171) | (~w38469 & ~w38336) | (~w43171 & ~w38336);
assign w52294 = (w37829 & ~w43182) | (w37829 & ~w37663) | (~w43182 & ~w37663);
assign w52295 = (~w38526 & ~w43181) | (~w38526 & ~w38336) | (~w43181 & ~w38336);
assign w52296 = (~w38962 & ~w43208) | (~w38962 & ~w37836) | (~w43208 & ~w37836);
assign w52297 = (~w38271 & ~w43226) | (~w38271 & ~w38197) | (~w43226 & ~w38197);
assign w52298 = (~w38291 & ~w43228) | (~w38291 & ~w38197) | (~w43228 & ~w38197);
assign w52299 = (~w39431 & ~w43232) | (~w39431 & ~w38142) | (~w43232 & ~w38142);
assign w52300 = w375 & ~w374;
assign w52301 = (~w332 & w406) | (~w332 & w50675) | (w406 & w50675);
assign w52302 = (~w332 & w409) | (~w332 & w50676) | (w409 & w50676);
assign w52303 = (~w332 & w427) | (~w332 & w50677) | (w427 & w50677);
assign w52304 = (w716 & w163) | (w716 & w50743) | (w163 & w50743);
assign w52305 = (w3 & ~w39824) | (w3 & ~w1319) | (~w39824 & ~w1319);
assign w52306 = (~w1554 & ~w39831) | (~w1554 & ~w1477) | (~w39831 & ~w1477);
assign w52307 = (w5628 & ~w40288) | (w5628 & ~w5590) | (~w40288 & ~w5590);
assign w52308 = (w5981 & ~w40335) | (w5981 & ~w5732) | (~w40335 & ~w5732);
assign w52309 = (w9090 & ~w40668) | (w9090 & ~w8985) | (~w40668 & ~w8985);
assign w52310 = (~w9094 & ~w40670) | (~w9094 & ~w8985) | (~w40670 & ~w8985);
assign w52311 = (~w1120 & ~w40881) | (~w1120 & ~w10396) | (~w40881 & ~w10396);
assign w52312 = (w12266 & ~w41049) | (w12266 & ~w11814) | (~w41049 & ~w11814);
assign w52313 = (~w19819 & ~w41720) | (~w19819 & ~w18827) | (~w41720 & ~w18827);
assign w52314 = (~w23411 & w50237) | (~w23411 & ~w22762) | (w50237 & ~w22762);
assign w52315 = (~w24394 & w50247) | (~w24394 & ~w24573) | (w50247 & ~w24573);
assign w52316 = (~w3242 & ~w42196) | (~w3242 & ~w24873) | (~w42196 & ~w24873);
assign w52317 = (w252 & ~w42207) | (w252 & ~w24873) | (~w42207 & ~w24873);
assign w52318 = (w27260 & w29093) | (w27260 & w50400) | (w29093 & w50400);
assign w52319 = w30034 & ~w30250;
assign w52320 = (w34016 & ~w42717) | (w34016 & ~w32997) | (~w42717 & ~w32997);
assign w52321 = (w33450 & ~w42764) | (w33450 & ~w33555) | (~w42764 & ~w33555);
assign w52322 = (w34729 & w42844) | (w34729 & ~w33695) | (w42844 & ~w33695);
assign w52323 = (~w332 & a[115]) | (~w332 & w50686) | (a[115] & w50686);
assign w52324 = (w1555 & ~w39832) | (w1555 & ~w1477) | (~w39832 & ~w1477);
assign w52325 = (w493 & ~w44213) | (w493 & ~w5328) | (~w44213 & ~w5328);
assign w52326 = (~w400 & ~w44216) | (~w400 & ~w5328) | (~w44216 & ~w5328);
assign w52327 = (w6243 & w6178) | (w6243 & w50414) | (w6178 & w50414);
assign w52328 = (w44337 & w44338) | (w44337 & ~w7787) | (w44338 & ~w7787);
assign w52329 = (~w11864 & w11815) | (~w11864 & ~w11869) | (w11815 & ~w11869);
assign w52330 = (w43475 & w43474) | (w43475 & ~w11332) | (w43474 & ~w11332);
assign w52331 = (w12334 & ~w12595) | (w12334 & w50590) | (~w12595 & w50590);
assign w52332 = (w14167 & ~w44759) | (w14167 & ~w14025) | (~w44759 & ~w14025);
assign w52333 = (w1594 & w1621) | (w1594 & w51431) | (w1621 & w51431);
assign w52334 = (~w80 & ~w47038) | (~w80 & ~w2864) | (~w47038 & ~w2864);
assign w52335 = (~w4055 & ~w400) | (~w4055 & w51446) | (~w400 & w51446);
assign w52336 = (~w28080 & ~w43620) | (~w28080 & ~w28049) | (~w43620 & ~w28049);
assign w52337 = (w80 & ~w43659) | (w80 & ~w28049) | (~w43659 & ~w28049);
assign w52338 = ~w2764 & w1320;
assign w52339 = (~w1727 & w50992) | (~w1727 & w1549) | (w50992 & w1549);
assign w52340 = (~w1727 & w50992) | (~w1727 & w47005) | (w50992 & w47005);
assign w52341 = (~w2100 & ~w51033) | (~w2100 & ~w2336) | (~w51033 & ~w2336);
assign w52342 = (w1727 & ~w50992) | (w1727 & ~w1706) | (~w50992 & ~w1706);
assign w52343 = (~w24394 & w52315) | (~w24394 & ~w24706) | (w52315 & ~w24706);
assign one = 1;
assign asqrt[0] = w39640;// level 690
assign asqrt[1] = ~w38339;// level 677
assign asqrt[2] = w37107;// level 663
assign asqrt[3] = ~w35994;// level 649
assign asqrt[4] = ~w34900;// level 632
assign asqrt[5] = ~w33731;// level 618
assign asqrt[6] = w32698;// level 605
assign asqrt[7] = ~w31477;// level 591
assign asqrt[8] = ~w30239;// level 576
assign asqrt[9] = ~w29158;// level 563
assign asqrt[10] = w28077;// level 549
assign asqrt[11] = ~w26880;// level 536
assign asqrt[12] = w25851;// level 523
assign asqrt[13] = w24874;// level 510
assign asqrt[14] = w23843;// level 497
assign asqrt[15] = w22767;// level 480
assign asqrt[16] = ~w21801;// level 467
assign asqrt[17] = w20906;// level 453
assign asqrt[18] = ~w20000;// level 440
assign asqrt[19] = ~w19040;// level 427
assign asqrt[20] = ~w18183;// level 414
assign asqrt[21] = w17380;// level 401
assign asqrt[22] = ~w16559;// level 389
assign asqrt[23] = ~w15681;// level 376
assign asqrt[24] = ~w14766;// level 363
assign asqrt[25] = w14039;// level 352
assign asqrt[26] = ~w13384;// level 340
assign asqrt[27] = w12666;// level 328
assign asqrt[28] = w11870;// level 315
assign asqrt[29] = ~w11138;// level 304
assign asqrt[30] = w10419;// level 292
assign asqrt[31] = w9781;// level 280
assign asqrt[32] = ~w9195;// level 268
assign asqrt[33] = w8666;// level 257
assign asqrt[34] = w7924;// level 246
assign asqrt[35] = w7315;// level 235
assign asqrt[36] = ~w6769;// level 224
assign asqrt[37] = w6264;// level 213
assign asqrt[38] = ~w5745;// level 202
assign asqrt[39] = w5330;// level 191
assign asqrt[40] = ~w4838;// level 180
assign asqrt[41] = w4430;// level 170
assign asqrt[42] = w4056;// level 160
assign asqrt[43] = ~w3646;// level 150
assign asqrt[44] = ~w3242;// level 140
assign asqrt[45] = w2896;// level 129
assign asqrt[46] = ~w2558;// level 119
assign asqrt[47] = w2285;// level 109
assign asqrt[48] = w2006;// level 100
assign asqrt[49] = w1738;// level 90
assign asqrt[50] = w1541;// level 82
assign asqrt[51] = w1320;// level 71
assign asqrt[52] = ~w1120;// level 62
assign asqrt[53] = ~w945;// level 54
assign asqrt[54] = w754;// level 46
assign asqrt[55] = w612;// level 39
assign asqrt[56] = w493;// level 31
assign asqrt[57] = ~w400;// level 25
assign asqrt[58] = w351;// level 18
assign asqrt[59] = ~w252;// level 13
assign asqrt[60] = ~w57;// level 8
assign asqrt[61] = w80;// level 4
assign asqrt[62] = ~w3;// level 3
assign asqrt[63] = ~w42;// level 1
endmodule

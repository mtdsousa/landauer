// Benchmark "t481" written by ABC on Sun Apr 22 21:43:14 2018

module t481 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15,
    po0  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15;
  output po0;
  wire n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
    n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
    n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890;
  assign n18 = ~pi01 & ~pi08;
  assign n19 = ~pi02 & n18;
  assign n20 = ~pi10 & n19;
  assign n21 = pi09 & n20;
  assign n22 = ~pi01 & ~pi09;
  assign n23 = ~pi02 & n22;
  assign n24 = ~pi11 & n23;
  assign n25 = pi10 & n24;
  assign n26 = ~pi01 & ~pi02;
  assign n27 = ~pi13 & ~pi14;
  assign n28 = n26 & n27;
  assign n29 = ~pi13 & pi15;
  assign n30 = n26 & n29;
  assign n31 = ~n21 & ~n25;
  assign n32 = ~n28 & ~n30;
  assign n33 = n31 & n32;
  assign n34 = pi08 & n26;
  assign n35 = pi10 & ~pi11;
  assign n36 = n34 & n35;
  assign n37 = pi09 & n19;
  assign n38 = pi11 & n37;
  assign n39 = pi12 & pi15;
  assign n40 = n26 & n39;
  assign n41 = ~pi01 & ~pi12;
  assign n42 = ~pi02 & n41;
  assign n43 = ~pi15 & n42;
  assign n44 = pi13 & pi14;
  assign n45 = n43 & n44;
  assign n46 = ~n36 & ~n38;
  assign n47 = ~n40 & ~n45;
  assign n48 = n46 & n47;
  assign n49 = pi12 & ~pi14;
  assign n50 = n26 & n49;
  assign n51 = ~pi02 & ~pi08;
  assign n52 = pi00 & n51;
  assign n53 = ~pi10 & n52;
  assign n54 = pi09 & n53;
  assign n55 = ~pi02 & ~pi09;
  assign n56 = pi00 & n55;
  assign n57 = ~pi11 & n56;
  assign n58 = pi10 & n57;
  assign n59 = pi00 & ~pi02;
  assign n60 = n27 & n59;
  assign n61 = ~n50 & ~n54;
  assign n62 = ~n58 & ~n60;
  assign n63 = n61 & n62;
  assign n64 = n29 & n59;
  assign n65 = pi08 & n35;
  assign n66 = n59 & n65;
  assign n67 = pi09 & n52;
  assign n68 = pi11 & n67;
  assign n69 = n39 & n59;
  assign n70 = ~n64 & ~n66;
  assign n71 = ~n68 & ~n69;
  assign n72 = n70 & n71;
  assign n73 = n33 & n48;
  assign n74 = n63 & n73;
  assign n75 = n72 & n74;
  assign n76 = pi04 & ~pi07;
  assign n77 = pi06 & n76;
  assign n78 = pi15 & n77;
  assign n79 = pi12 & n78;
  assign n80 = pi04 & pi06;
  assign n81 = ~pi07 & n80;
  assign n82 = ~pi12 & n81;
  assign n83 = ~pi15 & n82;
  assign n84 = n44 & n83;
  assign n85 = ~pi07 & n49;
  assign n86 = n80 & n85;
  assign n87 = pi03 & n18;
  assign n88 = ~pi10 & n87;
  assign n89 = pi09 & n88;
  assign n90 = ~n79 & ~n84;
  assign n91 = ~n86 & ~n89;
  assign n92 = n90 & n91;
  assign n93 = ~pi01 & pi03;
  assign n94 = ~pi13 & n93;
  assign n95 = pi15 & n94;
  assign n96 = ~pi09 & n35;
  assign n97 = ~pi01 & n96;
  assign n98 = pi03 & n97;
  assign n99 = ~pi14 & n94;
  assign n100 = n92 & ~n95;
  assign n101 = ~n98 & n100;
  assign n102 = ~n99 & n101;
  assign n103 = pi13 & ~pi15;
  assign n104 = pi14 & n103;
  assign n105 = ~pi12 & n104;
  assign n106 = ~pi02 & n105;
  assign n107 = pi00 & n106;
  assign n108 = ~pi14 & n59;
  assign n109 = pi12 & n108;
  assign n110 = ~pi10 & n77;
  assign n111 = ~pi08 & n110;
  assign n112 = pi09 & n111;
  assign n113 = ~pi11 & n77;
  assign n114 = ~pi09 & n113;
  assign n115 = pi10 & n114;
  assign n116 = ~n107 & ~n109;
  assign n117 = ~n112 & n116;
  assign n118 = ~n115 & n117;
  assign n119 = ~pi13 & n81;
  assign n120 = ~pi14 & n119;
  assign n121 = pi15 & n119;
  assign n122 = pi08 & n113;
  assign n123 = pi10 & n122;
  assign n124 = pi11 & n77;
  assign n125 = ~pi08 & n124;
  assign n126 = pi09 & n125;
  assign n127 = ~n120 & ~n121;
  assign n128 = ~n123 & n127;
  assign n129 = ~n126 & n128;
  assign n130 = n75 & n102;
  assign n131 = n118 & n129;
  assign n132 = n130 & n131;
  assign n133 = ~pi04 & ~pi06;
  assign n134 = pi05 & n133;
  assign n135 = ~pi10 & n134;
  assign n136 = ~pi08 & n135;
  assign n137 = pi09 & n136;
  assign n138 = ~pi11 & n134;
  assign n139 = ~pi09 & n138;
  assign n140 = pi10 & n139;
  assign n141 = ~pi04 & pi05;
  assign n142 = ~pi06 & n141;
  assign n143 = ~pi13 & n142;
  assign n144 = ~pi14 & n143;
  assign n145 = pi15 & n143;
  assign n146 = ~n137 & ~n140;
  assign n147 = ~n144 & n146;
  assign n148 = ~n145 & n147;
  assign n149 = pi15 & n134;
  assign n150 = pi12 & n149;
  assign n151 = pi08 & pi10;
  assign n152 = n138 & n151;
  assign n153 = pi11 & n134;
  assign n154 = ~pi08 & pi09;
  assign n155 = n153 & n154;
  assign n156 = n148 & ~n150;
  assign n157 = ~n152 & ~n155;
  assign n158 = n156 & n157;
  assign n159 = ~pi05 & ~pi07;
  assign n160 = pi06 & n159;
  assign n161 = ~pi11 & n160;
  assign n162 = ~pi09 & pi10;
  assign n163 = n161 & n162;
  assign n164 = ~pi07 & n27;
  assign n165 = ~pi05 & pi06;
  assign n166 = n164 & n165;
  assign n167 = ~pi13 & n160;
  assign n168 = pi15 & n167;
  assign n169 = n151 & n161;
  assign n170 = ~n163 & ~n166;
  assign n171 = ~n168 & ~n169;
  assign n172 = n170 & n171;
  assign n173 = pi11 & n160;
  assign n174 = n154 & n173;
  assign n175 = pi15 & n160;
  assign n176 = pi12 & n175;
  assign n177 = ~pi07 & n165;
  assign n178 = ~pi12 & n177;
  assign n179 = ~pi15 & n178;
  assign n180 = n44 & n179;
  assign n181 = ~pi14 & n160;
  assign n182 = pi12 & n181;
  assign n183 = ~n174 & ~n176;
  assign n184 = ~n180 & ~n182;
  assign n185 = n183 & n184;
  assign n186 = n158 & n172;
  assign n187 = n185 & n186;
  assign n188 = pi00 & pi03;
  assign n189 = n29 & n188;
  assign n190 = n65 & n188;
  assign n191 = pi00 & ~pi08;
  assign n192 = pi03 & n191;
  assign n193 = pi09 & n192;
  assign n194 = pi11 & n193;
  assign n195 = n39 & n188;
  assign n196 = ~n189 & ~n190;
  assign n197 = ~n194 & ~n195;
  assign n198 = n196 & n197;
  assign n199 = ~pi10 & n160;
  assign n200 = ~pi08 & n199;
  assign n201 = pi09 & n200;
  assign n202 = pi00 & ~pi12;
  assign n203 = pi03 & n202;
  assign n204 = ~pi15 & n203;
  assign n205 = pi13 & n204;
  assign n206 = pi14 & n205;
  assign n207 = ~pi14 & n188;
  assign n208 = pi12 & n207;
  assign n209 = n198 & ~n201;
  assign n210 = ~n206 & n209;
  assign n211 = ~n208 & n210;
  assign n212 = ~pi01 & pi08;
  assign n213 = pi03 & n212;
  assign n214 = ~pi11 & n213;
  assign n215 = pi10 & n214;
  assign n216 = pi09 & pi11;
  assign n217 = ~pi08 & n216;
  assign n218 = ~pi01 & n217;
  assign n219 = pi03 & n218;
  assign n220 = pi15 & n93;
  assign n221 = pi12 & n220;
  assign n222 = ~pi01 & n105;
  assign n223 = pi03 & n222;
  assign n224 = ~n215 & ~n219;
  assign n225 = ~n221 & n224;
  assign n226 = ~n223 & n225;
  assign n227 = ~pi14 & n93;
  assign n228 = pi12 & n227;
  assign n229 = ~pi08 & n188;
  assign n230 = ~pi10 & n229;
  assign n231 = pi09 & n230;
  assign n232 = ~pi09 & n188;
  assign n233 = ~pi11 & n232;
  assign n234 = pi10 & n233;
  assign n235 = ~pi13 & n188;
  assign n236 = ~pi14 & n235;
  assign n237 = ~n228 & ~n231;
  assign n238 = ~n234 & n237;
  assign n239 = ~n236 & n238;
  assign n240 = n187 & n211;
  assign n241 = n226 & n239;
  assign n242 = n240 & n241;
  assign n243 = ~pi00 & pi03;
  assign n244 = pi01 & n243;
  assign n245 = ~pi04 & pi06;
  assign n246 = pi05 & n245;
  assign n247 = ~pi07 & pi11;
  assign n248 = pi08 & n247;
  assign n249 = pi14 & ~pi15;
  assign n250 = pi12 & n249;
  assign n251 = n244 & n246;
  assign n252 = n248 & n251;
  assign n253 = n250 & n252;
  assign n254 = ~pi05 & ~pi06;
  assign n255 = ~pi02 & n254;
  assign n256 = ~pi00 & pi01;
  assign n257 = n255 & n256;
  assign n258 = pi08 & pi12;
  assign n259 = pi11 & n258;
  assign n260 = n257 & n259;
  assign n261 = ~pi15 & n260;
  assign n262 = pi14 & n261;
  assign n263 = pi03 & n254;
  assign n264 = n256 & n263;
  assign n265 = n259 & n264;
  assign n266 = ~pi15 & n265;
  assign n267 = pi14 & n266;
  assign n268 = ~pi00 & ~pi02;
  assign n269 = pi01 & n268;
  assign n270 = ~pi06 & n269;
  assign n271 = pi04 & n270;
  assign n272 = n259 & n271;
  assign n273 = ~pi15 & n272;
  assign n274 = pi14 & n273;
  assign n275 = ~n253 & ~n262;
  assign n276 = ~n267 & n275;
  assign n277 = ~n274 & n276;
  assign n278 = ~pi15 & n259;
  assign n279 = pi14 & n278;
  assign n280 = n244 & n279;
  assign n281 = ~pi05 & pi07;
  assign n282 = n280 & n281;
  assign n283 = pi04 & ~pi06;
  assign n284 = n280 & n283;
  assign n285 = n269 & n279;
  assign n286 = n281 & n285;
  assign n287 = n277 & ~n282;
  assign n288 = ~n284 & ~n286;
  assign n289 = n287 & n288;
  assign n290 = ~pi03 & n256;
  assign n291 = pi02 & n290;
  assign n292 = ~pi11 & n291;
  assign n293 = n151 & n292;
  assign n294 = pi11 & n291;
  assign n295 = n154 & n294;
  assign n296 = ~pi00 & pi02;
  assign n297 = pi01 & n296;
  assign n298 = pi15 & n297;
  assign n299 = ~pi03 & pi12;
  assign n300 = n298 & n299;
  assign n301 = ~pi12 & pi13;
  assign n302 = ~pi15 & n301;
  assign n303 = pi14 & n302;
  assign n304 = n291 & n303;
  assign n305 = ~n293 & ~n295;
  assign n306 = ~n300 & ~n304;
  assign n307 = n305 & n306;
  assign n308 = ~pi03 & ~pi14;
  assign n309 = pi12 & n308;
  assign n310 = pi02 & n309;
  assign n311 = n256 & n310;
  assign n312 = pi04 & pi07;
  assign n313 = n285 & n312;
  assign n314 = n280 & n312;
  assign n315 = ~pi02 & n246;
  assign n316 = ~pi00 & n315;
  assign n317 = pi01 & n316;
  assign n318 = ~pi15 & n248;
  assign n319 = pi14 & n318;
  assign n320 = pi12 & n319;
  assign n321 = n317 & n320;
  assign n322 = ~n311 & ~n313;
  assign n323 = ~n314 & ~n321;
  assign n324 = n322 & n323;
  assign n325 = n289 & n307;
  assign n326 = n324 & n325;
  assign n327 = pi07 & n141;
  assign n328 = n39 & n327;
  assign n329 = ~pi12 & n141;
  assign n330 = pi07 & n329;
  assign n331 = ~pi15 & n330;
  assign n332 = n44 & n331;
  assign n333 = n49 & n327;
  assign n334 = ~pi10 & n291;
  assign n335 = n154 & n334;
  assign n336 = ~n328 & ~n332;
  assign n337 = ~n333 & ~n335;
  assign n338 = n336 & n337;
  assign n339 = ~pi03 & n298;
  assign n340 = ~pi13 & n339;
  assign n341 = pi02 & ~pi03;
  assign n342 = n256 & n341;
  assign n343 = ~pi11 & n342;
  assign n344 = ~pi09 & n343;
  assign n345 = pi10 & n344;
  assign n346 = ~pi14 & n297;
  assign n347 = ~pi03 & n346;
  assign n348 = ~pi13 & n347;
  assign n349 = n338 & ~n340;
  assign n350 = ~n345 & n349;
  assign n351 = ~n348 & n350;
  assign n352 = ~pi06 & ~pi12;
  assign n353 = n141 & n352;
  assign n354 = ~pi15 & n353;
  assign n355 = pi13 & n354;
  assign n356 = pi14 & n355;
  assign n357 = ~pi14 & n142;
  assign n358 = pi12 & n357;
  assign n359 = ~pi04 & pi07;
  assign n360 = pi05 & n359;
  assign n361 = ~pi10 & n360;
  assign n362 = ~pi08 & n361;
  assign n363 = pi09 & n362;
  assign n364 = ~pi11 & n360;
  assign n365 = ~pi09 & n364;
  assign n366 = pi10 & n365;
  assign n367 = ~n356 & ~n358;
  assign n368 = ~n363 & n367;
  assign n369 = ~n366 & n368;
  assign n370 = ~pi13 & n360;
  assign n371 = ~pi14 & n370;
  assign n372 = pi15 & n370;
  assign n373 = pi08 & n364;
  assign n374 = pi10 & n373;
  assign n375 = pi11 & n360;
  assign n376 = ~pi08 & n375;
  assign n377 = pi09 & n376;
  assign n378 = ~n371 & ~n372;
  assign n379 = ~n374 & n378;
  assign n380 = ~n377 & n379;
  assign n381 = n326 & n351;
  assign n382 = n369 & n380;
  assign n383 = n381 & n382;
  assign n384 = ~pi03 & n283;
  assign n385 = pi00 & pi02;
  assign n386 = n384 & n385;
  assign n387 = ~pi10 & pi12;
  assign n388 = pi08 & n387;
  assign n389 = n386 & n388;
  assign n390 = ~pi15 & n389;
  assign n391 = pi14 & n390;
  assign n392 = ~pi07 & ~pi10;
  assign n393 = pi08 & n392;
  assign n394 = ~pi15 & n393;
  assign n395 = pi12 & pi14;
  assign n396 = n394 & n395;
  assign n397 = ~pi01 & pi02;
  assign n398 = n246 & n396;
  assign n399 = ~pi03 & n398;
  assign n400 = n397 & n399;
  assign n401 = n385 & n399;
  assign n402 = ~pi01 & ~pi03;
  assign n403 = pi02 & n402;
  assign n404 = ~pi05 & n403;
  assign n405 = pi07 & n404;
  assign n406 = n388 & n405;
  assign n407 = ~pi15 & n406;
  assign n408 = pi14 & n407;
  assign n409 = ~n391 & ~n400;
  assign n410 = ~n401 & n409;
  assign n411 = ~n408 & n410;
  assign n412 = ~pi15 & n388;
  assign n413 = pi14 & n412;
  assign n414 = n403 & n413;
  assign n415 = n312 & n414;
  assign n416 = ~pi03 & n385;
  assign n417 = ~pi05 & n416;
  assign n418 = pi07 & n417;
  assign n419 = n388 & n418;
  assign n420 = n249 & n419;
  assign n421 = ~pi02 & n312;
  assign n422 = ~pi00 & n421;
  assign n423 = pi01 & n422;
  assign n424 = ~pi09 & pi12;
  assign n425 = ~pi10 & n424;
  assign n426 = n423 & n425;
  assign n427 = n249 & n426;
  assign n428 = n411 & ~n415;
  assign n429 = ~n420 & ~n427;
  assign n430 = n428 & n429;
  assign n431 = ~pi05 & n244;
  assign n432 = ~pi06 & n431;
  assign n433 = n388 & n432;
  assign n434 = n249 & n433;
  assign n435 = n269 & n413;
  assign n436 = n283 & n435;
  assign n437 = n244 & n413;
  assign n438 = n283 & n437;
  assign n439 = n281 & n435;
  assign n440 = ~n434 & ~n436;
  assign n441 = ~n438 & ~n439;
  assign n442 = n440 & n441;
  assign n443 = n281 & n437;
  assign n444 = ~pi03 & n397;
  assign n445 = ~pi05 & n444;
  assign n446 = ~pi06 & n445;
  assign n447 = n388 & n446;
  assign n448 = n249 & n447;
  assign n449 = ~pi06 & n417;
  assign n450 = n388 & n449;
  assign n451 = n249 & n450;
  assign n452 = n283 & n414;
  assign n453 = ~n443 & ~n448;
  assign n454 = ~n451 & ~n452;
  assign n455 = n453 & n454;
  assign n456 = n430 & n442;
  assign n457 = n455 & n456;
  assign n458 = n312 & n435;
  assign n459 = n279 & n403;
  assign n460 = n312 & n459;
  assign n461 = pi00 & n341;
  assign n462 = n279 & n461;
  assign n463 = n312 & n462;
  assign n464 = n312 & n437;
  assign n465 = ~n458 & ~n460;
  assign n466 = ~n463 & ~n464;
  assign n467 = n465 & n466;
  assign n468 = n257 & n388;
  assign n469 = ~pi15 & n468;
  assign n470 = pi14 & n469;
  assign n471 = ~pi02 & n398;
  assign n472 = n256 & n471;
  assign n473 = n244 & n396;
  assign n474 = n246 & n473;
  assign n475 = n467 & ~n470;
  assign n476 = ~n472 & n475;
  assign n477 = ~n474 & n476;
  assign n478 = ~pi03 & n254;
  assign n479 = n397 & n478;
  assign n480 = n259 & n479;
  assign n481 = ~pi15 & n480;
  assign n482 = pi14 & n481;
  assign n483 = n385 & n478;
  assign n484 = n259 & n483;
  assign n485 = ~pi15 & n484;
  assign n486 = pi14 & n485;
  assign n487 = ~pi06 & n403;
  assign n488 = pi04 & n487;
  assign n489 = n259 & n488;
  assign n490 = ~pi15 & n489;
  assign n491 = pi14 & n490;
  assign n492 = n259 & n386;
  assign n493 = ~pi15 & n492;
  assign n494 = pi14 & n493;
  assign n495 = ~n482 & ~n486;
  assign n496 = ~n491 & n495;
  assign n497 = ~n494 & n496;
  assign n498 = pi06 & n403;
  assign n499 = n141 & n498;
  assign n500 = n248 & n499;
  assign n501 = ~pi15 & n500;
  assign n502 = n395 & n501;
  assign n503 = n246 & n461;
  assign n504 = n248 & n503;
  assign n505 = n250 & n504;
  assign n506 = n259 & n405;
  assign n507 = ~pi15 & n506;
  assign n508 = pi14 & n507;
  assign n509 = ~pi03 & n281;
  assign n510 = n385 & n509;
  assign n511 = n259 & n510;
  assign n512 = ~pi15 & n511;
  assign n513 = pi14 & n512;
  assign n514 = ~n502 & ~n505;
  assign n515 = ~n508 & n514;
  assign n516 = ~n513 & n515;
  assign n517 = n457 & n477;
  assign n518 = n497 & n516;
  assign n519 = n517 & n518;
  assign n520 = n132 & n242;
  assign n521 = n383 & n520;
  assign n522 = n519 & n521;
  assign n523 = ~pi10 & n250;
  assign n524 = ~pi07 & n523;
  assign n525 = ~pi09 & n524;
  assign n526 = n461 & n525;
  assign n527 = pi06 & n141;
  assign n528 = n526 & n527;
  assign n529 = ~pi01 & n509;
  assign n530 = pi02 & n529;
  assign n531 = n425 & n530;
  assign n532 = n249 & n531;
  assign n533 = n418 & n425;
  assign n534 = n249 & n533;
  assign n535 = ~pi09 & ~pi13;
  assign n536 = ~pi10 & n535;
  assign n537 = n423 & n536;
  assign n538 = n249 & n537;
  assign n539 = ~n528 & ~n532;
  assign n540 = ~n534 & ~n538;
  assign n541 = n539 & n540;
  assign n542 = ~pi03 & n312;
  assign n543 = ~pi01 & n542;
  assign n544 = pi02 & n543;
  assign n545 = n425 & n544;
  assign n546 = n249 & n545;
  assign n547 = pi02 & n542;
  assign n548 = pi00 & n547;
  assign n549 = n425 & n548;
  assign n550 = n249 & n549;
  assign n551 = pi03 & n312;
  assign n552 = ~pi00 & n551;
  assign n553 = pi01 & n552;
  assign n554 = n536 & n553;
  assign n555 = n249 & n554;
  assign n556 = ~pi09 & n392;
  assign n557 = ~pi13 & ~pi15;
  assign n558 = pi14 & n557;
  assign n559 = n317 & n556;
  assign n560 = n558 & n559;
  assign n561 = ~n546 & ~n550;
  assign n562 = ~n555 & ~n560;
  assign n563 = n561 & n562;
  assign n564 = pi03 & n246;
  assign n565 = ~pi00 & n564;
  assign n566 = pi01 & n565;
  assign n567 = n556 & n566;
  assign n568 = n558 & n567;
  assign n569 = ~pi02 & n256;
  assign n570 = ~pi05 & n569;
  assign n571 = ~pi06 & n570;
  assign n572 = n536 & n571;
  assign n573 = n249 & n572;
  assign n574 = n432 & n536;
  assign n575 = n249 & n574;
  assign n576 = ~pi02 & n283;
  assign n577 = ~pi00 & n576;
  assign n578 = pi01 & n577;
  assign n579 = n536 & n578;
  assign n580 = n249 & n579;
  assign n581 = ~n568 & ~n573;
  assign n582 = ~n575 & ~n580;
  assign n583 = n581 & n582;
  assign n584 = pi07 & n431;
  assign n585 = n536 & n584;
  assign n586 = n249 & n585;
  assign n587 = ~pi06 & n244;
  assign n588 = pi04 & n587;
  assign n589 = n536 & n588;
  assign n590 = n249 & n589;
  assign n591 = ~pi02 & n281;
  assign n592 = ~pi00 & n591;
  assign n593 = pi01 & n592;
  assign n594 = n536 & n593;
  assign n595 = n249 & n594;
  assign n596 = ~n586 & ~n590;
  assign n597 = ~n595 & n596;
  assign n598 = n541 & n563;
  assign n599 = n583 & n598;
  assign n600 = n597 & n599;
  assign n601 = n425 & n593;
  assign n602 = n249 & n601;
  assign n603 = n425 & n584;
  assign n604 = n249 & n603;
  assign n605 = n425 & n446;
  assign n606 = n249 & n605;
  assign n607 = n425 & n449;
  assign n608 = n249 & n607;
  assign n609 = ~n602 & ~n604;
  assign n610 = ~n606 & ~n608;
  assign n611 = n609 & n610;
  assign n612 = ~pi15 & n556;
  assign n613 = n395 & n612;
  assign n614 = n246 & n613;
  assign n615 = ~pi03 & n614;
  assign n616 = n397 & n615;
  assign n617 = ~pi09 & ~pi10;
  assign n618 = pi12 & n617;
  assign n619 = n249 & n618;
  assign n620 = n403 & n619;
  assign n621 = ~pi06 & n620;
  assign n622 = pi04 & n621;
  assign n623 = n461 & n619;
  assign n624 = ~pi06 & n623;
  assign n625 = pi04 & n624;
  assign n626 = n611 & ~n616;
  assign n627 = ~n622 & n626;
  assign n628 = ~n625 & n627;
  assign n629 = pi07 & n461;
  assign n630 = pi04 & n629;
  assign n631 = n388 & n630;
  assign n632 = ~pi15 & n631;
  assign n633 = pi14 & n632;
  assign n634 = n244 & n619;
  assign n635 = pi07 & n634;
  assign n636 = pi04 & n635;
  assign n637 = ~pi02 & n614;
  assign n638 = n256 & n637;
  assign n639 = n244 & n613;
  assign n640 = n246 & n639;
  assign n641 = ~n633 & ~n636;
  assign n642 = ~n638 & n641;
  assign n643 = ~n640 & n642;
  assign n644 = n269 & n619;
  assign n645 = ~pi05 & n644;
  assign n646 = ~pi06 & n645;
  assign n647 = ~pi05 & n634;
  assign n648 = ~pi06 & n647;
  assign n649 = ~pi06 & n644;
  assign n650 = pi04 & n649;
  assign n651 = ~pi06 & n634;
  assign n652 = pi04 & n651;
  assign n653 = ~n646 & ~n648;
  assign n654 = ~n650 & n653;
  assign n655 = ~n652 & n654;
  assign n656 = n600 & n628;
  assign n657 = n643 & n655;
  assign n658 = n656 & n657;
  assign n659 = ~pi09 & ~pi12;
  assign n660 = ~pi10 & n659;
  assign n661 = n432 & n660;
  assign n662 = pi13 & ~pi14;
  assign n663 = n661 & n662;
  assign n664 = n578 & n660;
  assign n665 = n662 & n664;
  assign n666 = n588 & n660;
  assign n667 = n662 & n666;
  assign n668 = n593 & n660;
  assign n669 = n662 & n668;
  assign n670 = ~n663 & ~n665;
  assign n671 = ~n667 & ~n669;
  assign n672 = n670 & n671;
  assign n673 = n584 & n660;
  assign n674 = n662 & n673;
  assign n675 = n446 & n660;
  assign n676 = n662 & n675;
  assign n677 = n449 & n660;
  assign n678 = n662 & n677;
  assign n679 = ~pi01 & n384;
  assign n680 = pi02 & n679;
  assign n681 = n660 & n680;
  assign n682 = n662 & n681;
  assign n683 = ~n674 & ~n676;
  assign n684 = ~n678 & ~n682;
  assign n685 = n683 & n684;
  assign n686 = ~pi06 & n416;
  assign n687 = pi04 & n686;
  assign n688 = n660 & n687;
  assign n689 = n662 & n688;
  assign n690 = ~pi03 & n246;
  assign n691 = ~pi01 & n690;
  assign n692 = pi02 & n691;
  assign n693 = ~pi12 & ~pi14;
  assign n694 = pi13 & n693;
  assign n695 = n556 & n692;
  assign n696 = n694 & n695;
  assign n697 = pi02 & n690;
  assign n698 = pi00 & n697;
  assign n699 = n556 & n698;
  assign n700 = n694 & n699;
  assign n701 = n530 & n660;
  assign n702 = n662 & n701;
  assign n703 = ~n689 & ~n696;
  assign n704 = ~n700 & ~n702;
  assign n705 = n703 & n704;
  assign n706 = n548 & n660;
  assign n707 = n662 & n706;
  assign n708 = n418 & n660;
  assign n709 = n662 & n708;
  assign n710 = n544 & n660;
  assign n711 = n662 & n710;
  assign n712 = ~n707 & ~n709;
  assign n713 = ~n711 & n712;
  assign n714 = n672 & n685;
  assign n715 = n705 & n714;
  assign n716 = n713 & n715;
  assign n717 = n423 & n660;
  assign n718 = n662 & n717;
  assign n719 = n536 & n544;
  assign n720 = n249 & n719;
  assign n721 = n536 & n548;
  assign n722 = n249 & n721;
  assign n723 = n553 & n660;
  assign n724 = n662 & n723;
  assign n725 = ~n718 & ~n720;
  assign n726 = ~n722 & ~n724;
  assign n727 = n725 & n726;
  assign n728 = ~pi14 & n660;
  assign n729 = pi13 & n728;
  assign n730 = n269 & n729;
  assign n731 = ~pi05 & n730;
  assign n732 = ~pi06 & n731;
  assign n733 = ~pi14 & n556;
  assign n734 = n301 & n733;
  assign n735 = n246 & n734;
  assign n736 = ~pi02 & n735;
  assign n737 = n256 & n736;
  assign n738 = n244 & n734;
  assign n739 = n246 & n738;
  assign n740 = n727 & ~n732;
  assign n741 = ~n737 & n740;
  assign n742 = ~n739 & n741;
  assign n743 = ~pi15 & n536;
  assign n744 = pi14 & n743;
  assign n745 = n403 & n744;
  assign n746 = ~pi05 & n745;
  assign n747 = ~pi06 & n746;
  assign n748 = n461 & n744;
  assign n749 = ~pi05 & n748;
  assign n750 = ~pi06 & n749;
  assign n751 = ~pi06 & n745;
  assign n752 = pi04 & n751;
  assign n753 = ~pi06 & n748;
  assign n754 = pi04 & n753;
  assign n755 = ~n747 & ~n750;
  assign n756 = ~n752 & n755;
  assign n757 = ~n754 & n756;
  assign n758 = ~pi13 & pi14;
  assign n759 = n612 & n758;
  assign n760 = n246 & n759;
  assign n761 = ~pi03 & n760;
  assign n762 = n397 & n761;
  assign n763 = n385 & n761;
  assign n764 = pi07 & n746;
  assign n765 = pi07 & n749;
  assign n766 = ~n762 & ~n763;
  assign n767 = ~n764 & n766;
  assign n768 = ~n765 & n767;
  assign n769 = n716 & n742;
  assign n770 = n757 & n768;
  assign n771 = n769 & n770;
  assign n772 = pi11 & n558;
  assign n773 = ~pi07 & pi08;
  assign n774 = n772 & n773;
  assign n775 = n244 & n774;
  assign n776 = n246 & n775;
  assign n777 = pi08 & ~pi13;
  assign n778 = pi11 & n777;
  assign n779 = n257 & n778;
  assign n780 = ~pi15 & n779;
  assign n781 = pi14 & n780;
  assign n782 = n264 & n778;
  assign n783 = ~pi15 & n782;
  assign n784 = pi14 & n783;
  assign n785 = n271 & n778;
  assign n786 = ~pi15 & n785;
  assign n787 = pi14 & n786;
  assign n788 = ~n776 & ~n781;
  assign n789 = ~n784 & n788;
  assign n790 = ~n787 & n789;
  assign n791 = pi08 & pi11;
  assign n792 = ~pi13 & n791;
  assign n793 = ~pi15 & n792;
  assign n794 = pi14 & n793;
  assign n795 = n244 & n794;
  assign n796 = n281 & n795;
  assign n797 = n283 & n795;
  assign n798 = n269 & n794;
  assign n799 = n281 & n798;
  assign n800 = n790 & ~n796;
  assign n801 = ~n797 & ~n799;
  assign n802 = n800 & n801;
  assign n803 = ~pi07 & ~pi09;
  assign n804 = n250 & n698;
  assign n805 = pi11 & n803;
  assign n806 = n804 & n805;
  assign n807 = pi11 & n424;
  assign n808 = ~pi15 & n807;
  assign n809 = pi14 & n808;
  assign n810 = n403 & n809;
  assign n811 = n281 & n810;
  assign n812 = n418 & n807;
  assign n813 = n249 & n812;
  assign n814 = n312 & n810;
  assign n815 = ~n806 & ~n811;
  assign n816 = ~n813 & ~n814;
  assign n817 = n815 & n816;
  assign n818 = n461 & n809;
  assign n819 = n312 & n818;
  assign n820 = n312 & n798;
  assign n821 = n312 & n795;
  assign n822 = ~pi13 & n318;
  assign n823 = pi14 & n822;
  assign n824 = n317 & n823;
  assign n825 = ~n819 & ~n820;
  assign n826 = ~n821 & ~n824;
  assign n827 = n825 & n826;
  assign n828 = n802 & n817;
  assign n829 = n827 & n828;
  assign n830 = n269 & n809;
  assign n831 = n281 & n830;
  assign n832 = n244 & n809;
  assign n833 = n281 & n832;
  assign n834 = n446 & n807;
  assign n835 = n249 & n834;
  assign n836 = n449 & n807;
  assign n837 = n249 & n836;
  assign n838 = ~n831 & ~n833;
  assign n839 = ~n835 & ~n837;
  assign n840 = n838 & n839;
  assign n841 = ~pi09 & n247;
  assign n842 = ~pi15 & n841;
  assign n843 = n395 & n842;
  assign n844 = n246 & n843;
  assign n845 = ~pi03 & n844;
  assign n846 = n397 & n845;
  assign n847 = n488 & n807;
  assign n848 = ~pi15 & n847;
  assign n849 = pi14 & n848;
  assign n850 = n386 & n807;
  assign n851 = ~pi15 & n850;
  assign n852 = pi14 & n851;
  assign n853 = n840 & ~n846;
  assign n854 = ~n849 & n853;
  assign n855 = ~n852 & n854;
  assign n856 = pi07 & n269;
  assign n857 = pi04 & n856;
  assign n858 = n807 & n857;
  assign n859 = ~pi15 & n858;
  assign n860 = pi14 & n859;
  assign n861 = pi03 & n256;
  assign n862 = n312 & n861;
  assign n863 = n807 & n862;
  assign n864 = ~pi15 & n863;
  assign n865 = pi14 & n864;
  assign n866 = ~pi02 & n844;
  assign n867 = n256 & n866;
  assign n868 = n244 & n843;
  assign n869 = n246 & n868;
  assign n870 = ~n860 & ~n865;
  assign n871 = ~n867 & n870;
  assign n872 = ~n869 & n871;
  assign n873 = n257 & n807;
  assign n874 = ~pi15 & n873;
  assign n875 = pi14 & n874;
  assign n876 = n264 & n807;
  assign n877 = ~pi15 & n876;
  assign n878 = pi14 & n877;
  assign n879 = n271 & n807;
  assign n880 = ~pi15 & n879;
  assign n881 = pi14 & n880;
  assign n882 = pi03 & n283;
  assign n883 = n256 & n882;
  assign n884 = n807 & n883;
  assign n885 = ~pi15 & n884;
  assign n886 = pi14 & n885;
  assign n887 = ~n875 & ~n878;
  assign n888 = ~n881 & n887;
  assign n889 = ~n886 & n888;
  assign n890 = n829 & n855;
  assign n891 = n872 & n889;
  assign n892 = n890 & n891;
  assign n893 = ~pi10 & ~pi13;
  assign n894 = pi08 & n893;
  assign n895 = n432 & n894;
  assign n896 = n249 & n895;
  assign n897 = n578 & n894;
  assign n898 = n249 & n897;
  assign n899 = n588 & n894;
  assign n900 = n249 & n899;
  assign n901 = n593 & n894;
  assign n902 = n249 & n901;
  assign n903 = ~n896 & ~n898;
  assign n904 = ~n900 & ~n902;
  assign n905 = n903 & n904;
  assign n906 = n584 & n894;
  assign n907 = n249 & n906;
  assign n908 = n446 & n894;
  assign n909 = n249 & n908;
  assign n910 = n449 & n894;
  assign n911 = n249 & n910;
  assign n912 = n680 & n894;
  assign n913 = n249 & n912;
  assign n914 = ~n907 & ~n909;
  assign n915 = ~n911 & ~n913;
  assign n916 = n914 & n915;
  assign n917 = n687 & n894;
  assign n918 = n249 & n917;
  assign n919 = n393 & n692;
  assign n920 = n558 & n919;
  assign n921 = n393 & n698;
  assign n922 = n558 & n921;
  assign n923 = n530 & n894;
  assign n924 = n249 & n923;
  assign n925 = ~n918 & ~n920;
  assign n926 = ~n922 & ~n924;
  assign n927 = n925 & n926;
  assign n928 = n548 & n894;
  assign n929 = n249 & n928;
  assign n930 = n418 & n894;
  assign n931 = n249 & n930;
  assign n932 = n544 & n894;
  assign n933 = n249 & n932;
  assign n934 = ~n929 & ~n931;
  assign n935 = ~n933 & n934;
  assign n936 = n905 & n916;
  assign n937 = n927 & n936;
  assign n938 = n935 & n937;
  assign n939 = n423 & n894;
  assign n940 = n249 & n939;
  assign n941 = n403 & n794;
  assign n942 = n312 & n941;
  assign n943 = n461 & n794;
  assign n944 = n312 & n943;
  assign n945 = n553 & n894;
  assign n946 = n249 & n945;
  assign n947 = ~n940 & ~n942;
  assign n948 = ~n944 & ~n946;
  assign n949 = n947 & n948;
  assign n950 = ~pi15 & n894;
  assign n951 = pi14 & n950;
  assign n952 = n269 & n951;
  assign n953 = ~pi05 & n952;
  assign n954 = ~pi06 & n953;
  assign n955 = n394 & n758;
  assign n956 = n246 & n955;
  assign n957 = ~pi02 & n956;
  assign n958 = n256 & n957;
  assign n959 = n244 & n955;
  assign n960 = n246 & n959;
  assign n961 = n949 & ~n954;
  assign n962 = ~n958 & n961;
  assign n963 = ~n960 & n962;
  assign n964 = n479 & n778;
  assign n965 = ~pi15 & n964;
  assign n966 = pi14 & n965;
  assign n967 = n483 & n778;
  assign n968 = ~pi15 & n967;
  assign n969 = pi14 & n968;
  assign n970 = n488 & n778;
  assign n971 = ~pi15 & n970;
  assign n972 = pi14 & n971;
  assign n973 = n386 & n778;
  assign n974 = ~pi15 & n973;
  assign n975 = pi14 & n974;
  assign n976 = ~n966 & ~n969;
  assign n977 = ~n972 & n976;
  assign n978 = ~n975 & n977;
  assign n979 = n499 & n774;
  assign n980 = n246 & n774;
  assign n981 = ~pi03 & n980;
  assign n982 = n385 & n981;
  assign n983 = n405 & n778;
  assign n984 = ~pi15 & n983;
  assign n985 = pi14 & n984;
  assign n986 = n510 & n778;
  assign n987 = ~pi15 & n986;
  assign n988 = pi14 & n987;
  assign n989 = ~n979 & ~n982;
  assign n990 = ~n985 & n989;
  assign n991 = ~n988 & n990;
  assign n992 = n938 & n963;
  assign n993 = n978 & n991;
  assign n994 = n992 & n993;
  assign n995 = n658 & n771;
  assign n996 = n892 & n995;
  assign n997 = n994 & n996;
  assign n998 = pi11 & n535;
  assign n999 = n423 & n998;
  assign n1000 = n249 & n999;
  assign n1001 = n553 & n998;
  assign n1002 = n249 & n1001;
  assign n1003 = n317 & n558;
  assign n1004 = n805 & n1003;
  assign n1005 = n558 & n566;
  assign n1006 = n805 & n1005;
  assign n1007 = ~n1000 & ~n1002;
  assign n1008 = ~n1004 & ~n1006;
  assign n1009 = n1007 & n1008;
  assign n1010 = n571 & n998;
  assign n1011 = n249 & n1010;
  assign n1012 = n432 & n998;
  assign n1013 = n249 & n1012;
  assign n1014 = n578 & n998;
  assign n1015 = n249 & n1014;
  assign n1016 = n588 & n998;
  assign n1017 = n249 & n1016;
  assign n1018 = ~n1011 & ~n1013;
  assign n1019 = ~n1015 & ~n1017;
  assign n1020 = n1018 & n1019;
  assign n1021 = n593 & n998;
  assign n1022 = n249 & n1021;
  assign n1023 = n584 & n998;
  assign n1024 = n249 & n1023;
  assign n1025 = n446 & n998;
  assign n1026 = n249 & n1025;
  assign n1027 = n449 & n998;
  assign n1028 = n249 & n1027;
  assign n1029 = ~n1022 & ~n1024;
  assign n1030 = ~n1026 & ~n1028;
  assign n1031 = n1029 & n1030;
  assign n1032 = n558 & n692;
  assign n1033 = n805 & n1032;
  assign n1034 = n680 & n998;
  assign n1035 = n249 & n1034;
  assign n1036 = n687 & n998;
  assign n1037 = n249 & n1036;
  assign n1038 = ~n1033 & ~n1035;
  assign n1039 = ~n1037 & n1038;
  assign n1040 = n1009 & n1020;
  assign n1041 = n1031 & n1040;
  assign n1042 = n1039 & n1041;
  assign n1043 = n566 & n694;
  assign n1044 = n805 & n1043;
  assign n1045 = pi11 & n659;
  assign n1046 = n571 & n1045;
  assign n1047 = n662 & n1046;
  assign n1048 = n432 & n1045;
  assign n1049 = n662 & n1048;
  assign n1050 = n578 & n1045;
  assign n1051 = n662 & n1050;
  assign n1052 = ~n1044 & ~n1047;
  assign n1053 = ~n1049 & ~n1051;
  assign n1054 = n1052 & n1053;
  assign n1055 = ~pi14 & n1045;
  assign n1056 = pi13 & n1055;
  assign n1057 = n244 & n1056;
  assign n1058 = ~pi05 & n1057;
  assign n1059 = pi07 & n1058;
  assign n1060 = ~pi06 & n1057;
  assign n1061 = pi04 & n1060;
  assign n1062 = n269 & n1056;
  assign n1063 = ~pi05 & n1062;
  assign n1064 = pi07 & n1063;
  assign n1065 = n1054 & ~n1059;
  assign n1066 = ~n1061 & n1065;
  assign n1067 = ~n1064 & n1066;
  assign n1068 = n758 & n842;
  assign n1069 = n246 & n1068;
  assign n1070 = ~pi03 & n1069;
  assign n1071 = n385 & n1070;
  assign n1072 = ~pi15 & n998;
  assign n1073 = pi14 & n1072;
  assign n1074 = n403 & n1073;
  assign n1075 = ~pi05 & n1074;
  assign n1076 = pi07 & n1075;
  assign n1077 = n461 & n1073;
  assign n1078 = ~pi05 & n1077;
  assign n1079 = pi07 & n1078;
  assign n1080 = n857 & n1045;
  assign n1081 = ~pi14 & n1080;
  assign n1082 = pi13 & n1081;
  assign n1083 = ~n1071 & ~n1076;
  assign n1084 = ~n1079 & n1083;
  assign n1085 = ~n1082 & n1084;
  assign n1086 = pi07 & n403;
  assign n1087 = pi04 & n1086;
  assign n1088 = n998 & n1087;
  assign n1089 = ~pi15 & n1088;
  assign n1090 = pi14 & n1089;
  assign n1091 = n630 & n998;
  assign n1092 = ~pi15 & n1091;
  assign n1093 = pi14 & n1092;
  assign n1094 = n862 & n1045;
  assign n1095 = ~pi14 & n1094;
  assign n1096 = pi13 & n1095;
  assign n1097 = ~pi14 & n841;
  assign n1098 = n301 & n1097;
  assign n1099 = n246 & n1098;
  assign n1100 = ~pi02 & n1099;
  assign n1101 = n256 & n1100;
  assign n1102 = ~n1090 & ~n1093;
  assign n1103 = ~n1096 & n1102;
  assign n1104 = ~n1101 & n1103;
  assign n1105 = n1042 & n1067;
  assign n1106 = n1085 & n1104;
  assign n1107 = n1105 & n1106;
  assign n1108 = n1045 & n1087;
  assign n1109 = ~pi14 & n1108;
  assign n1110 = pi13 & n1109;
  assign n1111 = n630 & n1045;
  assign n1112 = ~pi14 & n1111;
  assign n1113 = pi13 & n1112;
  assign n1114 = ~pi08 & n269;
  assign n1115 = n312 & n1114;
  assign n1116 = pi09 & pi10;
  assign n1117 = n250 & n1115;
  assign n1118 = ~pi11 & n1117;
  assign n1119 = n1116 & n1118;
  assign n1120 = ~pi08 & n244;
  assign n1121 = n312 & n1120;
  assign n1122 = n250 & n1121;
  assign n1123 = ~pi11 & n1122;
  assign n1124 = n1116 & n1123;
  assign n1125 = ~n1110 & ~n1113;
  assign n1126 = ~n1119 & n1125;
  assign n1127 = ~n1124 & n1126;
  assign n1128 = pi09 & ~pi11;
  assign n1129 = pi10 & n1128;
  assign n1130 = ~pi15 & n1129;
  assign n1131 = pi14 & n1130;
  assign n1132 = pi12 & n1131;
  assign n1133 = ~pi05 & ~pi08;
  assign n1134 = ~pi06 & n1133;
  assign n1135 = n269 & n1132;
  assign n1136 = n1134 & n1135;
  assign n1137 = n35 & n154;
  assign n1138 = ~pi15 & n1137;
  assign n1139 = pi14 & n1138;
  assign n1140 = pi12 & n1139;
  assign n1141 = ~pi04 & n569;
  assign n1142 = pi06 & ~pi07;
  assign n1143 = pi05 & n1142;
  assign n1144 = n1140 & n1141;
  assign n1145 = n1143 & n1144;
  assign n1146 = ~pi04 & n256;
  assign n1147 = pi03 & n1146;
  assign n1148 = n1140 & n1147;
  assign n1149 = n1143 & n1148;
  assign n1150 = n1127 & ~n1136;
  assign n1151 = ~n1145 & ~n1149;
  assign n1152 = n1150 & n1151;
  assign n1153 = n446 & n1045;
  assign n1154 = n662 & n1153;
  assign n1155 = n449 & n1045;
  assign n1156 = n662 & n1155;
  assign n1157 = n680 & n1045;
  assign n1158 = n662 & n1157;
  assign n1159 = n687 & n1045;
  assign n1160 = n662 & n1159;
  assign n1161 = ~n1154 & ~n1156;
  assign n1162 = ~n1158 & ~n1160;
  assign n1163 = n1161 & n1162;
  assign n1164 = n692 & n694;
  assign n1165 = n805 & n1164;
  assign n1166 = n694 & n698;
  assign n1167 = n805 & n1166;
  assign n1168 = n530 & n1045;
  assign n1169 = n662 & n1168;
  assign n1170 = n418 & n1045;
  assign n1171 = n662 & n1170;
  assign n1172 = ~n1165 & ~n1167;
  assign n1173 = ~n1169 & ~n1171;
  assign n1174 = n1172 & n1173;
  assign n1175 = n1152 & n1163;
  assign n1176 = n1174 & n1175;
  assign n1177 = ~pi08 & n461;
  assign n1178 = ~pi06 & n1177;
  assign n1179 = pi04 & n1178;
  assign n1180 = n1132 & n1179;
  assign n1181 = ~pi04 & n444;
  assign n1182 = n1140 & n1181;
  assign n1183 = n1143 & n1182;
  assign n1184 = ~pi04 & n416;
  assign n1185 = n1140 & n1184;
  assign n1186 = n1143 & n1185;
  assign n1187 = pi07 & n1133;
  assign n1188 = n403 & n1132;
  assign n1189 = n1187 & n1188;
  assign n1190 = ~n1180 & ~n1183;
  assign n1191 = ~n1186 & ~n1189;
  assign n1192 = n1190 & n1191;
  assign n1193 = ~pi08 & n403;
  assign n1194 = n312 & n1193;
  assign n1195 = n250 & n1194;
  assign n1196 = ~pi11 & n1195;
  assign n1197 = n1116 & n1196;
  assign n1198 = ~pi03 & n1187;
  assign n1199 = n385 & n1198;
  assign n1200 = n250 & n1199;
  assign n1201 = ~pi11 & n1200;
  assign n1202 = n1116 & n1201;
  assign n1203 = n558 & n1115;
  assign n1204 = ~pi11 & n1203;
  assign n1205 = n1116 & n1204;
  assign n1206 = n1192 & ~n1197;
  assign n1207 = ~n1202 & n1206;
  assign n1208 = ~n1205 & n1207;
  assign n1209 = pi03 & n1134;
  assign n1210 = n256 & n1209;
  assign n1211 = n250 & n1210;
  assign n1212 = ~pi11 & n1211;
  assign n1213 = n1116 & n1212;
  assign n1214 = ~pi06 & ~pi08;
  assign n1215 = pi04 & n1214;
  assign n1216 = ~pi02 & n1215;
  assign n1217 = n256 & n1216;
  assign n1218 = n250 & n1217;
  assign n1219 = ~pi11 & n1218;
  assign n1220 = n1116 & n1219;
  assign n1221 = pi03 & n1215;
  assign n1222 = n256 & n1221;
  assign n1223 = n250 & n1222;
  assign n1224 = ~pi11 & n1223;
  assign n1225 = n1116 & n1224;
  assign n1226 = ~pi02 & n1187;
  assign n1227 = n256 & n1226;
  assign n1228 = n250 & n1227;
  assign n1229 = ~pi11 & n1228;
  assign n1230 = n1116 & n1229;
  assign n1231 = ~n1213 & ~n1220;
  assign n1232 = ~n1225 & n1231;
  assign n1233 = ~n1230 & n1232;
  assign n1234 = pi03 & n1187;
  assign n1235 = n256 & n1234;
  assign n1236 = n250 & n1235;
  assign n1237 = ~pi11 & n1236;
  assign n1238 = n1116 & n1237;
  assign n1239 = ~pi03 & n1134;
  assign n1240 = n397 & n1239;
  assign n1241 = n250 & n1240;
  assign n1242 = ~pi11 & n1241;
  assign n1243 = n1116 & n1242;
  assign n1244 = n385 & n1239;
  assign n1245 = n250 & n1244;
  assign n1246 = ~pi11 & n1245;
  assign n1247 = n1116 & n1246;
  assign n1248 = ~pi03 & n1215;
  assign n1249 = n397 & n1248;
  assign n1250 = n250 & n1249;
  assign n1251 = ~pi11 & n1250;
  assign n1252 = n1116 & n1251;
  assign n1253 = ~n1238 & ~n1243;
  assign n1254 = ~n1247 & n1253;
  assign n1255 = ~n1252 & n1254;
  assign n1256 = n1176 & n1208;
  assign n1257 = n1233 & n1255;
  assign n1258 = n1256 & n1257;
  assign n1259 = ~pi13 & n1138;
  assign n1260 = pi14 & n1259;
  assign n1261 = n1184 & n1260;
  assign n1262 = n1143 & n1261;
  assign n1263 = ~pi13 & n1130;
  assign n1264 = pi14 & n1263;
  assign n1265 = n403 & n1264;
  assign n1266 = n1187 & n1265;
  assign n1267 = ~pi05 & n1177;
  assign n1268 = pi07 & n1267;
  assign n1269 = n1264 & n1268;
  assign n1270 = pi07 & ~pi08;
  assign n1271 = pi04 & n1270;
  assign n1272 = ~pi03 & n1271;
  assign n1273 = ~pi01 & n1272;
  assign n1274 = pi02 & n1273;
  assign n1275 = n1264 & n1274;
  assign n1276 = ~n1262 & ~n1266;
  assign n1277 = ~n1269 & ~n1275;
  assign n1278 = n1276 & n1277;
  assign n1279 = pi02 & n1272;
  assign n1280 = pi00 & n1279;
  assign n1281 = n1264 & n1280;
  assign n1282 = ~pi12 & n791;
  assign n1283 = pi13 & n1282;
  assign n1284 = pi15 & n1283;
  assign n1285 = n269 & n1284;
  assign n1286 = n312 & n1285;
  assign n1287 = n244 & n1284;
  assign n1288 = n312 & n1287;
  assign n1289 = pi15 & n248;
  assign n1290 = ~pi12 & n1289;
  assign n1291 = pi13 & n1290;
  assign n1292 = n317 & n1291;
  assign n1293 = ~n1281 & ~n1286;
  assign n1294 = ~n1288 & ~n1292;
  assign n1295 = n1293 & n1294;
  assign n1296 = n566 & n1291;
  assign n1297 = pi08 & ~pi12;
  assign n1298 = pi11 & n1297;
  assign n1299 = n571 & n1298;
  assign n1300 = pi13 & pi15;
  assign n1301 = n1299 & n1300;
  assign n1302 = n432 & n1298;
  assign n1303 = n1300 & n1302;
  assign n1304 = n283 & n1285;
  assign n1305 = ~n1296 & ~n1301;
  assign n1306 = ~n1303 & ~n1304;
  assign n1307 = n1305 & n1306;
  assign n1308 = n584 & n1298;
  assign n1309 = n1300 & n1308;
  assign n1310 = n588 & n1298;
  assign n1311 = n1300 & n1310;
  assign n1312 = n281 & n1285;
  assign n1313 = ~n1309 & ~n1311;
  assign n1314 = ~n1312 & n1313;
  assign n1315 = n1278 & n1295;
  assign n1316 = n1307 & n1315;
  assign n1317 = n1314 & n1316;
  assign n1318 = n269 & n1264;
  assign n1319 = n1187 & n1318;
  assign n1320 = n1187 & n1264;
  assign n1321 = n861 & n1320;
  assign n1322 = n1134 & n1265;
  assign n1323 = ~pi06 & n1267;
  assign n1324 = n1264 & n1323;
  assign n1325 = ~n1319 & ~n1321;
  assign n1326 = ~n1322 & ~n1324;
  assign n1327 = n1325 & n1326;
  assign n1328 = ~pi07 & n1181;
  assign n1329 = pi05 & pi06;
  assign n1330 = n1328 & n1329;
  assign n1331 = n1137 & n1330;
  assign n1332 = ~pi15 & n1331;
  assign n1333 = n758 & n1332;
  assign n1334 = n558 & n1249;
  assign n1335 = ~pi11 & n1334;
  assign n1336 = n1116 & n1335;
  assign n1337 = n385 & n1248;
  assign n1338 = n558 & n1337;
  assign n1339 = ~pi11 & n1338;
  assign n1340 = n1116 & n1339;
  assign n1341 = n1327 & ~n1333;
  assign n1342 = ~n1336 & n1341;
  assign n1343 = ~n1340 & n1342;
  assign n1344 = n312 & n1177;
  assign n1345 = n250 & n1344;
  assign n1346 = ~pi11 & n1345;
  assign n1347 = n1116 & n1346;
  assign n1348 = ~pi11 & n558;
  assign n1349 = n1116 & n1348;
  assign n1350 = n244 & n1349;
  assign n1351 = ~pi08 & n1350;
  assign n1352 = n312 & n1351;
  assign n1353 = ~pi07 & n1141;
  assign n1354 = n1329 & n1353;
  assign n1355 = n1137 & n1354;
  assign n1356 = ~pi15 & n1355;
  assign n1357 = n758 & n1356;
  assign n1358 = ~pi11 & n154;
  assign n1359 = pi10 & n1358;
  assign n1360 = ~pi15 & n1359;
  assign n1361 = n758 & n1360;
  assign n1362 = pi03 & ~pi04;
  assign n1363 = n256 & n1362;
  assign n1364 = n1361 & n1363;
  assign n1365 = ~pi07 & n1364;
  assign n1366 = n1329 & n1365;
  assign n1367 = ~n1347 & ~n1352;
  assign n1368 = ~n1357 & n1367;
  assign n1369 = ~n1366 & n1368;
  assign n1370 = ~pi02 & n1134;
  assign n1371 = n256 & n1370;
  assign n1372 = n558 & n1371;
  assign n1373 = ~pi11 & n1372;
  assign n1374 = n1116 & n1373;
  assign n1375 = n558 & n1210;
  assign n1376 = ~pi11 & n1375;
  assign n1377 = n1116 & n1376;
  assign n1378 = n558 & n1217;
  assign n1379 = ~pi11 & n1378;
  assign n1380 = n1116 & n1379;
  assign n1381 = n558 & n1222;
  assign n1382 = ~pi11 & n1381;
  assign n1383 = n1116 & n1382;
  assign n1384 = ~n1374 & ~n1377;
  assign n1385 = ~n1380 & n1384;
  assign n1386 = ~n1383 & n1385;
  assign n1387 = n1317 & n1343;
  assign n1388 = n1369 & n1386;
  assign n1389 = n1387 & n1388;
  assign n1390 = ~pi10 & ~pi12;
  assign n1391 = pi08 & n1390;
  assign n1392 = n432 & n1391;
  assign n1393 = n1300 & n1392;
  assign n1394 = ~pi12 & n1300;
  assign n1395 = ~pi10 & n1394;
  assign n1396 = pi08 & n1395;
  assign n1397 = n269 & n1396;
  assign n1398 = n283 & n1397;
  assign n1399 = n588 & n1391;
  assign n1400 = n1300 & n1399;
  assign n1401 = n281 & n1397;
  assign n1402 = ~n1393 & ~n1398;
  assign n1403 = ~n1400 & ~n1401;
  assign n1404 = n1402 & n1403;
  assign n1405 = n584 & n1391;
  assign n1406 = n1300 & n1405;
  assign n1407 = n446 & n1391;
  assign n1408 = n1300 & n1407;
  assign n1409 = n449 & n1391;
  assign n1410 = n1300 & n1409;
  assign n1411 = n403 & n1396;
  assign n1412 = n283 & n1411;
  assign n1413 = ~n1406 & ~n1408;
  assign n1414 = ~n1410 & ~n1412;
  assign n1415 = n1413 & n1414;
  assign n1416 = n687 & n1391;
  assign n1417 = n1300 & n1416;
  assign n1418 = pi15 & n301;
  assign n1419 = n919 & n1418;
  assign n1420 = n921 & n1418;
  assign n1421 = n281 & n1411;
  assign n1422 = ~n1417 & ~n1419;
  assign n1423 = ~n1420 & ~n1421;
  assign n1424 = n1422 & n1423;
  assign n1425 = n312 & n1411;
  assign n1426 = n418 & n1391;
  assign n1427 = n1300 & n1426;
  assign n1428 = ~pi09 & n1394;
  assign n1429 = ~pi10 & n1428;
  assign n1430 = n269 & n1429;
  assign n1431 = n312 & n1430;
  assign n1432 = ~n1425 & ~n1427;
  assign n1433 = ~n1431 & n1432;
  assign n1434 = n1404 & n1415;
  assign n1435 = n1424 & n1434;
  assign n1436 = n1433 & n1435;
  assign n1437 = n312 & n1397;
  assign n1438 = n403 & n1284;
  assign n1439 = n312 & n1438;
  assign n1440 = n461 & n1284;
  assign n1441 = n312 & n1440;
  assign n1442 = n244 & n1396;
  assign n1443 = n312 & n1442;
  assign n1444 = ~n1437 & ~n1439;
  assign n1445 = ~n1441 & ~n1443;
  assign n1446 = n1444 & n1445;
  assign n1447 = pi13 & n1391;
  assign n1448 = pi15 & n1447;
  assign n1449 = n269 & n1448;
  assign n1450 = ~pi05 & n1449;
  assign n1451 = ~pi06 & n1450;
  assign n1452 = pi15 & n393;
  assign n1453 = n301 & n1452;
  assign n1454 = n246 & n1453;
  assign n1455 = ~pi02 & n1454;
  assign n1456 = n256 & n1455;
  assign n1457 = n244 & n1453;
  assign n1458 = n246 & n1457;
  assign n1459 = n1446 & ~n1451;
  assign n1460 = ~n1456 & n1459;
  assign n1461 = ~n1458 & n1460;
  assign n1462 = pi13 & n1298;
  assign n1463 = pi15 & n1462;
  assign n1464 = n403 & n1463;
  assign n1465 = ~pi05 & n1464;
  assign n1466 = ~pi06 & n1465;
  assign n1467 = n461 & n1463;
  assign n1468 = ~pi05 & n1467;
  assign n1469 = ~pi06 & n1468;
  assign n1470 = n488 & n1298;
  assign n1471 = pi13 & n1470;
  assign n1472 = pi15 & n1471;
  assign n1473 = ~pi06 & n1467;
  assign n1474 = pi04 & n1473;
  assign n1475 = ~n1466 & ~n1469;
  assign n1476 = ~n1472 & n1475;
  assign n1477 = ~n1474 & n1476;
  assign n1478 = ~pi12 & pi15;
  assign n1479 = pi13 & n1478;
  assign n1480 = n500 & n1479;
  assign n1481 = n504 & n1479;
  assign n1482 = n405 & n1298;
  assign n1483 = pi13 & n1482;
  assign n1484 = pi15 & n1483;
  assign n1485 = pi07 & n1468;
  assign n1486 = ~n1480 & ~n1481;
  assign n1487 = ~n1484 & n1486;
  assign n1488 = ~n1485 & n1487;
  assign n1489 = n1436 & n1461;
  assign n1490 = n1477 & n1488;
  assign n1491 = n1489 & n1490;
  assign n1492 = n1107 & n1258;
  assign n1493 = n1389 & n1492;
  assign n1494 = n1491 & n1493;
  assign n1495 = ~pi10 & n1479;
  assign n1496 = ~pi07 & n1495;
  assign n1497 = ~pi09 & n1496;
  assign n1498 = n461 & n1497;
  assign n1499 = n527 & n1498;
  assign n1500 = n403 & n1429;
  assign n1501 = n281 & n1500;
  assign n1502 = n708 & n1300;
  assign n1503 = n312 & n1500;
  assign n1504 = ~n1499 & ~n1501;
  assign n1505 = ~n1502 & ~n1503;
  assign n1506 = n1504 & n1505;
  assign n1507 = n461 & n1429;
  assign n1508 = n312 & n1507;
  assign n1509 = pi11 & n1428;
  assign n1510 = n269 & n1509;
  assign n1511 = n312 & n1510;
  assign n1512 = n244 & n1509;
  assign n1513 = n312 & n1512;
  assign n1514 = n317 & n1479;
  assign n1515 = n805 & n1514;
  assign n1516 = ~n1508 & ~n1511;
  assign n1517 = ~n1513 & ~n1515;
  assign n1518 = n1516 & n1517;
  assign n1519 = n566 & n1479;
  assign n1520 = n805 & n1519;
  assign n1521 = n1046 & n1300;
  assign n1522 = n1048 & n1300;
  assign n1523 = n283 & n1510;
  assign n1524 = ~n1520 & ~n1521;
  assign n1525 = ~n1522 & ~n1523;
  assign n1526 = n1524 & n1525;
  assign n1527 = n584 & n1045;
  assign n1528 = n1300 & n1527;
  assign n1529 = n588 & n1045;
  assign n1530 = n1300 & n1529;
  assign n1531 = n281 & n1510;
  assign n1532 = ~n1528 & ~n1530;
  assign n1533 = ~n1531 & n1532;
  assign n1534 = n1506 & n1518;
  assign n1535 = n1526 & n1534;
  assign n1536 = n1533 & n1535;
  assign n1537 = n281 & n1430;
  assign n1538 = n673 & n1300;
  assign n1539 = n675 & n1300;
  assign n1540 = n677 & n1300;
  assign n1541 = ~n1537 & ~n1538;
  assign n1542 = ~n1539 & ~n1540;
  assign n1543 = n1541 & n1542;
  assign n1544 = pi15 & n556;
  assign n1545 = n301 & n1544;
  assign n1546 = n246 & n1545;
  assign n1547 = ~pi03 & n1546;
  assign n1548 = n397 & n1547;
  assign n1549 = pi13 & n660;
  assign n1550 = pi15 & n1549;
  assign n1551 = n403 & n1550;
  assign n1552 = ~pi06 & n1551;
  assign n1553 = pi04 & n1552;
  assign n1554 = n461 & n1550;
  assign n1555 = ~pi06 & n1554;
  assign n1556 = pi04 & n1555;
  assign n1557 = n1543 & ~n1548;
  assign n1558 = ~n1553 & n1557;
  assign n1559 = ~n1556 & n1558;
  assign n1560 = n461 & n1448;
  assign n1561 = pi07 & n1560;
  assign n1562 = pi04 & n1561;
  assign n1563 = n244 & n1550;
  assign n1564 = pi07 & n1563;
  assign n1565 = pi04 & n1564;
  assign n1566 = ~pi02 & n1546;
  assign n1567 = n256 & n1566;
  assign n1568 = n244 & n1545;
  assign n1569 = n246 & n1568;
  assign n1570 = ~n1562 & ~n1565;
  assign n1571 = ~n1567 & n1570;
  assign n1572 = ~n1569 & n1571;
  assign n1573 = n269 & n1550;
  assign n1574 = ~pi05 & n1573;
  assign n1575 = ~pi06 & n1574;
  assign n1576 = ~pi05 & n1563;
  assign n1577 = ~pi06 & n1576;
  assign n1578 = ~pi06 & n1573;
  assign n1579 = pi04 & n1578;
  assign n1580 = ~pi06 & n1563;
  assign n1581 = pi04 & n1580;
  assign n1582 = ~n1575 & ~n1577;
  assign n1583 = ~n1579 & n1582;
  assign n1584 = ~n1581 & n1583;
  assign n1585 = n1536 & n1559;
  assign n1586 = n1572 & n1584;
  assign n1587 = n1585 & n1586;
  assign n1588 = n386 & n1298;
  assign n1589 = ~pi14 & n1588;
  assign n1590 = pi13 & n1589;
  assign n1591 = pi11 & n694;
  assign n1592 = n773 & n1591;
  assign n1593 = n499 & n1592;
  assign n1594 = n246 & n1592;
  assign n1595 = ~pi03 & n1594;
  assign n1596 = n385 & n1595;
  assign n1597 = ~pi14 & n1482;
  assign n1598 = pi13 & n1597;
  assign n1599 = ~n1590 & ~n1593;
  assign n1600 = ~n1596 & n1599;
  assign n1601 = ~n1598 & n1600;
  assign n1602 = ~pi14 & n1282;
  assign n1603 = pi13 & n1602;
  assign n1604 = n403 & n1603;
  assign n1605 = n312 & n1604;
  assign n1606 = n461 & n1603;
  assign n1607 = n281 & n1606;
  assign n1608 = n423 & n1391;
  assign n1609 = n662 & n1608;
  assign n1610 = n1601 & ~n1605;
  assign n1611 = ~n1607 & ~n1609;
  assign n1612 = n1610 & n1611;
  assign n1613 = n662 & n1302;
  assign n1614 = n269 & n1603;
  assign n1615 = n283 & n1614;
  assign n1616 = n244 & n1603;
  assign n1617 = n283 & n1616;
  assign n1618 = n281 & n1614;
  assign n1619 = ~n1613 & ~n1615;
  assign n1620 = ~n1617 & ~n1618;
  assign n1621 = n1619 & n1620;
  assign n1622 = n281 & n1616;
  assign n1623 = n254 & n1604;
  assign n1624 = n449 & n1298;
  assign n1625 = n662 & n1624;
  assign n1626 = n283 & n1604;
  assign n1627 = ~n1622 & ~n1623;
  assign n1628 = ~n1625 & ~n1626;
  assign n1629 = n1627 & n1628;
  assign n1630 = n1612 & n1621;
  assign n1631 = n1629 & n1630;
  assign n1632 = n403 & n1509;
  assign n1633 = n312 & n1632;
  assign n1634 = n461 & n1509;
  assign n1635 = n312 & n1634;
  assign n1636 = n312 & n1614;
  assign n1637 = n312 & n1616;
  assign n1638 = ~n1633 & ~n1635;
  assign n1639 = ~n1636 & ~n1637;
  assign n1640 = n1638 & n1639;
  assign n1641 = n257 & n1298;
  assign n1642 = ~pi14 & n1641;
  assign n1643 = pi13 & n1642;
  assign n1644 = pi06 & n269;
  assign n1645 = n141 & n1644;
  assign n1646 = n1592 & n1645;
  assign n1647 = n244 & n1592;
  assign n1648 = n246 & n1647;
  assign n1649 = n1640 & ~n1643;
  assign n1650 = ~n1646 & n1649;
  assign n1651 = ~n1648 & n1650;
  assign n1652 = pi13 & n1045;
  assign n1653 = pi15 & n1652;
  assign n1654 = n403 & n1653;
  assign n1655 = ~pi05 & n1654;
  assign n1656 = ~pi06 & n1655;
  assign n1657 = n461 & n1653;
  assign n1658 = ~pi05 & n1657;
  assign n1659 = ~pi06 & n1658;
  assign n1660 = ~pi06 & n1654;
  assign n1661 = pi04 & n1660;
  assign n1662 = ~pi06 & n1657;
  assign n1663 = pi04 & n1662;
  assign n1664 = ~n1656 & ~n1659;
  assign n1665 = ~n1661 & n1664;
  assign n1666 = ~n1663 & n1665;
  assign n1667 = pi15 & n841;
  assign n1668 = n301 & n1667;
  assign n1669 = n246 & n1668;
  assign n1670 = ~pi03 & n1669;
  assign n1671 = n397 & n1670;
  assign n1672 = n385 & n1670;
  assign n1673 = pi07 & n1655;
  assign n1674 = pi07 & n1658;
  assign n1675 = ~n1671 & ~n1672;
  assign n1676 = ~n1673 & n1675;
  assign n1677 = ~n1674 & n1676;
  assign n1678 = n1631 & n1651;
  assign n1679 = n1666 & n1677;
  assign n1680 = n1678 & n1679;
  assign n1681 = n312 & n1606;
  assign n1682 = n553 & n1391;
  assign n1683 = n662 & n1682;
  assign n1684 = n317 & n393;
  assign n1685 = n694 & n1684;
  assign n1686 = n393 & n566;
  assign n1687 = n694 & n1686;
  assign n1688 = ~n1681 & ~n1683;
  assign n1689 = ~n1685 & ~n1687;
  assign n1690 = n1688 & n1689;
  assign n1691 = n571 & n1391;
  assign n1692 = n662 & n1691;
  assign n1693 = n662 & n1392;
  assign n1694 = n578 & n1391;
  assign n1695 = n662 & n1694;
  assign n1696 = n662 & n1399;
  assign n1697 = ~n1692 & ~n1693;
  assign n1698 = ~n1695 & ~n1696;
  assign n1699 = n1697 & n1698;
  assign n1700 = n593 & n1391;
  assign n1701 = n662 & n1700;
  assign n1702 = n662 & n1405;
  assign n1703 = n662 & n1407;
  assign n1704 = n662 & n1409;
  assign n1705 = ~n1701 & ~n1702;
  assign n1706 = ~n1703 & ~n1704;
  assign n1707 = n1705 & n1706;
  assign n1708 = n694 & n919;
  assign n1709 = n680 & n1391;
  assign n1710 = n662 & n1709;
  assign n1711 = n662 & n1416;
  assign n1712 = ~n1708 & ~n1710;
  assign n1713 = ~n1711 & n1712;
  assign n1714 = n1690 & n1699;
  assign n1715 = n1707 & n1714;
  assign n1716 = n1713 & n1715;
  assign n1717 = ~pi07 & n1363;
  assign n1718 = pi06 & n1717;
  assign n1719 = pi05 & n1718;
  assign n1720 = n1359 & n1719;
  assign n1721 = n1418 & n1720;
  assign n1722 = pi15 & n1129;
  assign n1723 = ~pi12 & n1722;
  assign n1724 = pi13 & n1723;
  assign n1725 = n269 & n1724;
  assign n1726 = n1134 & n1725;
  assign n1727 = n1134 & n1724;
  assign n1728 = n861 & n1727;
  assign n1729 = n1215 & n1725;
  assign n1730 = ~n1721 & ~n1726;
  assign n1731 = ~n1728 & ~n1729;
  assign n1732 = n1730 & n1731;
  assign n1733 = n1235 & n1479;
  assign n1734 = ~pi11 & n1733;
  assign n1735 = n1116 & n1734;
  assign n1736 = n1222 & n1479;
  assign n1737 = ~pi11 & n1736;
  assign n1738 = n1116 & n1737;
  assign n1739 = n1227 & n1479;
  assign n1740 = ~pi11 & n1739;
  assign n1741 = n1116 & n1740;
  assign n1742 = n1732 & ~n1735;
  assign n1743 = ~n1738 & n1742;
  assign n1744 = ~n1741 & n1743;
  assign n1745 = ~pi14 & n393;
  assign n1746 = n301 & n1745;
  assign n1747 = n246 & n1746;
  assign n1748 = ~pi03 & n1747;
  assign n1749 = n385 & n1748;
  assign n1750 = ~pi14 & n1391;
  assign n1751 = pi13 & n1750;
  assign n1752 = n403 & n1751;
  assign n1753 = ~pi05 & n1752;
  assign n1754 = pi07 & n1753;
  assign n1755 = n461 & n1751;
  assign n1756 = ~pi05 & n1755;
  assign n1757 = pi07 & n1756;
  assign n1758 = n1087 & n1391;
  assign n1759 = ~pi14 & n1758;
  assign n1760 = pi13 & n1759;
  assign n1761 = ~n1749 & ~n1754;
  assign n1762 = ~n1757 & n1761;
  assign n1763 = ~n1760 & n1762;
  assign n1764 = n630 & n1391;
  assign n1765 = ~pi14 & n1764;
  assign n1766 = pi13 & n1765;
  assign n1767 = n1115 & n1479;
  assign n1768 = ~pi11 & n1767;
  assign n1769 = n1116 & n1768;
  assign n1770 = n1121 & n1479;
  assign n1771 = ~pi11 & n1770;
  assign n1772 = n1116 & n1771;
  assign n1773 = pi15 & n1359;
  assign n1774 = n301 & n1773;
  assign n1775 = n1354 & n1774;
  assign n1776 = ~n1766 & ~n1769;
  assign n1777 = ~n1772 & n1776;
  assign n1778 = ~n1775 & n1777;
  assign n1779 = n1716 & n1744;
  assign n1780 = n1763 & n1778;
  assign n1781 = n1779 & n1780;
  assign n1782 = n694 & n1337;
  assign n1783 = ~pi11 & n1782;
  assign n1784 = n1116 & n1783;
  assign n1785 = ~pi14 & n1331;
  assign n1786 = n301 & n1785;
  assign n1787 = ~pi14 & n1359;
  assign n1788 = n301 & n1787;
  assign n1789 = ~pi03 & ~pi04;
  assign n1790 = n385 & n1789;
  assign n1791 = n1788 & n1790;
  assign n1792 = ~pi07 & n1791;
  assign n1793 = n1329 & n1792;
  assign n1794 = n397 & n1198;
  assign n1795 = n694 & n1794;
  assign n1796 = ~pi11 & n1795;
  assign n1797 = n1116 & n1796;
  assign n1798 = ~n1784 & ~n1786;
  assign n1799 = ~n1793 & n1798;
  assign n1800 = ~n1797 & n1799;
  assign n1801 = ~pi14 & n1129;
  assign n1802 = ~pi12 & n1801;
  assign n1803 = pi13 & n1802;
  assign n1804 = n1280 & n1803;
  assign n1805 = n1268 & n1803;
  assign n1806 = n1274 & n1803;
  assign n1807 = n1800 & ~n1804;
  assign n1808 = ~n1805 & ~n1806;
  assign n1809 = n1807 & n1808;
  assign n1810 = n1134 & n1803;
  assign n1811 = n861 & n1810;
  assign n1812 = n269 & n1803;
  assign n1813 = n1215 & n1812;
  assign n1814 = n1215 & n1803;
  assign n1815 = n861 & n1814;
  assign n1816 = n1187 & n1812;
  assign n1817 = ~n1811 & ~n1813;
  assign n1818 = ~n1815 & ~n1816;
  assign n1819 = n1817 & n1818;
  assign n1820 = n1187 & n1803;
  assign n1821 = n861 & n1820;
  assign n1822 = n403 & n1803;
  assign n1823 = n1134 & n1822;
  assign n1824 = n1323 & n1803;
  assign n1825 = n1215 & n1822;
  assign n1826 = ~n1821 & ~n1823;
  assign n1827 = ~n1824 & ~n1825;
  assign n1828 = n1826 & n1827;
  assign n1829 = n1809 & n1819;
  assign n1830 = n1828 & n1829;
  assign n1831 = ~pi02 & n1271;
  assign n1832 = ~pi00 & n1831;
  assign n1833 = pi01 & n1832;
  assign n1834 = n1803 & n1833;
  assign n1835 = n1274 & n1724;
  assign n1836 = n1280 & n1724;
  assign n1837 = pi03 & n1271;
  assign n1838 = ~pi00 & n1837;
  assign n1839 = pi01 & n1838;
  assign n1840 = n1803 & n1839;
  assign n1841 = ~n1834 & ~n1835;
  assign n1842 = ~n1836 & ~n1840;
  assign n1843 = n1841 & n1842;
  assign n1844 = n694 & n1371;
  assign n1845 = ~pi11 & n1844;
  assign n1846 = n1116 & n1845;
  assign n1847 = ~pi14 & n1355;
  assign n1848 = n301 & n1847;
  assign n1849 = n1363 & n1788;
  assign n1850 = ~pi07 & n1849;
  assign n1851 = n1329 & n1850;
  assign n1852 = n1843 & ~n1846;
  assign n1853 = ~n1848 & n1852;
  assign n1854 = ~n1851 & n1853;
  assign n1855 = n1240 & n1479;
  assign n1856 = ~pi11 & n1855;
  assign n1857 = n1116 & n1856;
  assign n1858 = n1244 & n1479;
  assign n1859 = ~pi11 & n1858;
  assign n1860 = n1116 & n1859;
  assign n1861 = n1249 & n1479;
  assign n1862 = ~pi11 & n1861;
  assign n1863 = n1116 & n1862;
  assign n1864 = n1337 & n1479;
  assign n1865 = ~pi11 & n1864;
  assign n1866 = n1116 & n1865;
  assign n1867 = ~n1857 & ~n1860;
  assign n1868 = ~n1863 & n1867;
  assign n1869 = ~n1866 & n1868;
  assign n1870 = n1330 & n1774;
  assign n1871 = n1774 & n1790;
  assign n1872 = ~pi07 & n1871;
  assign n1873 = n1329 & n1872;
  assign n1874 = n1479 & n1794;
  assign n1875 = ~pi11 & n1874;
  assign n1876 = n1116 & n1875;
  assign n1877 = n1199 & n1479;
  assign n1878 = ~pi11 & n1877;
  assign n1879 = n1116 & n1878;
  assign n1880 = ~n1870 & ~n1873;
  assign n1881 = ~n1876 & n1880;
  assign n1882 = ~n1879 & n1881;
  assign n1883 = n1830 & n1854;
  assign n1884 = n1869 & n1882;
  assign n1885 = n1883 & n1884;
  assign n1886 = n1587 & n1680;
  assign n1887 = n1781 & n1886;
  assign n1888 = n1885 & n1887;
  assign n1889 = n522 & n997;
  assign n1890 = n1494 & n1888;
  assign po0 = ~n1889 | ~n1890;
endmodule



module top (
            a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, a_64, a_65, a_66, a_67, a_68, a_69, a_70, a_71, a_72, a_73, a_74, a_75, a_76, a_77, a_78, a_79, a_80, a_81, a_82, a_83, a_84, a_85, a_86, a_87, a_88, a_89, a_90, a_91, a_92, a_93, a_94, a_95, a_96, a_97, a_98, a_99, a_100, a_101, a_102, a_103, a_104, a_105, a_106, a_107, a_108, a_109, a_110, a_111, a_112, a_113, a_114, a_115, a_116, a_117, a_118, a_119, a_120, a_121, a_122, a_123, a_124, a_125, a_126, a_127, b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, b_8, b_9, b_10, b_11, b_12, b_13, b_14, b_15, b_16, b_17, b_18, b_19, b_20, b_21, b_22, b_23, b_24, b_25, b_26, b_27, b_28, b_29, b_30, b_31, b_32, b_33, b_34, b_35, b_36, b_37, b_38, b_39, b_40, b_41, b_42, b_43, b_44, b_45, b_46, b_47, b_48, b_49, b_50, b_51, b_52, b_53, b_54, b_55, b_56, b_57, b_58, b_59, b_60, b_61, b_62, b_63, b_64, b_65, b_66, b_67, b_68, b_69, b_70, b_71, b_72, b_73, b_74, b_75, b_76, b_77, b_78, b_79, b_80, b_81, b_82, b_83, b_84, b_85, b_86, b_87, b_88, b_89, b_90, b_91, b_92, b_93, b_94, b_95, b_96, b_97, b_98, b_99, b_100, b_101, b_102, b_103, b_104, b_105, b_106, b_107, b_108, b_109, b_110, b_111, b_112, b_113, b_114, b_115, b_116, b_117, b_118, b_119, b_120, b_121, b_122, b_123, b_124, b_125, b_126, b_127, 
            f_0, f_1, f_2, f_3, f_4, f_5, f_6, f_7, f_8, f_9, f_10, f_11, f_12, f_13, f_14, f_15, f_16, f_17, f_18, f_19, f_20, f_21, f_22, f_23, f_24, f_25, f_26, f_27, f_28, f_29, f_30, f_31, f_32, f_33, f_34, f_35, f_36, f_37, f_38, f_39, f_40, f_41, f_42, f_43, f_44, f_45, f_46, f_47, f_48, f_49, f_50, f_51, f_52, f_53, f_54, f_55, f_56, f_57, f_58, f_59, f_60, f_61, f_62, f_63, f_64, f_65, f_66, f_67, f_68, f_69, f_70, f_71, f_72, f_73, f_74, f_75, f_76, f_77, f_78, f_79, f_80, f_81, f_82, f_83, f_84, f_85, f_86, f_87, f_88, f_89, f_90, f_91, f_92, f_93, f_94, f_95, f_96, f_97, f_98, f_99, f_100, f_101, f_102, f_103, f_104, f_105, f_106, f_107, f_108, f_109, f_110, f_111, f_112, f_113, f_114, f_115, f_116, f_117, f_118, f_119, f_120, f_121, f_122, f_123, f_124, f_125, f_126, f_127, cOut);
input a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, a_64, a_65, a_66, a_67, a_68, a_69, a_70, a_71, a_72, a_73, a_74, a_75, a_76, a_77, a_78, a_79, a_80, a_81, a_82, a_83, a_84, a_85, a_86, a_87, a_88, a_89, a_90, a_91, a_92, a_93, a_94, a_95, a_96, a_97, a_98, a_99, a_100, a_101, a_102, a_103, a_104, a_105, a_106, a_107, a_108, a_109, a_110, a_111, a_112, a_113, a_114, a_115, a_116, a_117, a_118, a_119, a_120, a_121, a_122, a_123, a_124, a_125, a_126, a_127, b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, b_8, b_9, b_10, b_11, b_12, b_13, b_14, b_15, b_16, b_17, b_18, b_19, b_20, b_21, b_22, b_23, b_24, b_25, b_26, b_27, b_28, b_29, b_30, b_31, b_32, b_33, b_34, b_35, b_36, b_37, b_38, b_39, b_40, b_41, b_42, b_43, b_44, b_45, b_46, b_47, b_48, b_49, b_50, b_51, b_52, b_53, b_54, b_55, b_56, b_57, b_58, b_59, b_60, b_61, b_62, b_63, b_64, b_65, b_66, b_67, b_68, b_69, b_70, b_71, b_72, b_73, b_74, b_75, b_76, b_77, b_78, b_79, b_80, b_81, b_82, b_83, b_84, b_85, b_86, b_87, b_88, b_89, b_90, b_91, b_92, b_93, b_94, b_95, b_96, b_97, b_98, b_99, b_100, b_101, b_102, b_103, b_104, b_105, b_106, b_107, b_108, b_109, b_110, b_111, b_112, b_113, b_114, b_115, b_116, b_117, b_118, b_119, b_120, b_121, b_122, b_123, b_124, b_125, b_126, b_127;
output f_0, f_1, f_2, f_3, f_4, f_5, f_6, f_7, f_8, f_9, f_10, f_11, f_12, f_13, f_14, f_15, f_16, f_17, f_18, f_19, f_20, f_21, f_22, f_23, f_24, f_25, f_26, f_27, f_28, f_29, f_30, f_31, f_32, f_33, f_34, f_35, f_36, f_37, f_38, f_39, f_40, f_41, f_42, f_43, f_44, f_45, f_46, f_47, f_48, f_49, f_50, f_51, f_52, f_53, f_54, f_55, f_56, f_57, f_58, f_59, f_60, f_61, f_62, f_63, f_64, f_65, f_66, f_67, f_68, f_69, f_70, f_71, f_72, f_73, f_74, f_75, f_76, f_77, f_78, f_79, f_80, f_81, f_82, f_83, f_84, f_85, f_86, f_87, f_88, f_89, f_90, f_91, f_92, f_93, f_94, f_95, f_96, f_97, f_98, f_99, f_100, f_101, f_102, f_103, f_104, f_105, f_106, f_107, f_108, f_109, f_110, f_111, f_112, f_113, f_114, f_115, f_116, f_117, f_118, f_119, f_120, f_121, f_122, f_123, f_124, f_125, f_126, f_127, cOut;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981;
assign w0 = a_0 & ~b_0;
assign w1 = ~a_0 & b_0;
assign w2 = ~w0 & ~w1;
assign w3 = a_0 & b_0;
assign w4 = ~a_1 & ~b_1;
assign w5 = a_1 & b_1;
assign w6 = ~w4 & ~w5;
assign w7 = w3 & ~w6;
assign w8 = ~w3 & w6;
assign w9 = ~w7 & ~w8;
assign w10 = w3 & ~w4;
assign w11 = ~w5 & ~w10;
assign w12 = ~a_2 & ~b_2;
assign w13 = a_2 & b_2;
assign w14 = ~w12 & ~w13;
assign w15 = w11 & ~w14;
assign w16 = ~w11 & w14;
assign w17 = ~w15 & ~w16;
assign w18 = (~w12 & w10) | (~w12 & w815) | (w10 & w815);
assign w19 = ~a_3 & ~b_3;
assign w20 = a_3 & b_3;
assign w21 = ~w19 & ~w20;
assign w22 = ~w18 & w1261;
assign w23 = (w21 & w18) | (w21 & w1262) | (w18 & w1262);
assign w24 = ~w22 & ~w23;
assign w25 = (~w18 & w817) | (~w18 & w818) | (w817 & w818);
assign w26 = ~a_4 & ~b_4;
assign w27 = a_4 & b_4;
assign w28 = ~w26 & ~w27;
assign w29 = w25 & ~w28;
assign w30 = ~w25 & w28;
assign w31 = ~w29 & ~w30;
assign w32 = ~a_5 & ~b_5;
assign w33 = a_5 & b_5;
assign w34 = ~w32 & ~w33;
assign w35 = (w25 & w1263) | (w25 & w1264) | (w1263 & w1264);
assign w36 = w34 & w2786;
assign w37 = ~w35 & ~w36;
assign w38 = (w25 & w821) | (w25 & w822) | (w821 & w822);
assign w39 = ~a_6 & ~b_6;
assign w40 = a_6 & b_6;
assign w41 = ~w39 & ~w40;
assign w42 = (w25 & w1265) | (w25 & w1266) | (w1265 & w1266);
assign w43 = w41 & ~w38;
assign w44 = ~w42 & ~w43;
assign w45 = (w25 & w1267) | (w25 & w1268) | (w1267 & w1268);
assign w46 = ~a_7 & ~b_7;
assign w47 = a_7 & b_7;
assign w48 = ~w46 & ~w47;
assign w49 = w45 & ~w48;
assign w50 = ~w45 & w48;
assign w51 = ~w49 & ~w50;
assign w52 = (w25 & w1269) | (w25 & w1270) | (w1269 & w1270);
assign w53 = ~a_8 & ~b_8;
assign w54 = a_8 & b_8;
assign w55 = ~w53 & ~w54;
assign w56 = w52 & ~w55;
assign w57 = ~w52 & w55;
assign w58 = ~w56 & ~w57;
assign w59 = (~w38 & w827) | (~w38 & w828) | (w827 & w828);
assign w60 = ~a_9 & ~b_9;
assign w61 = a_9 & b_9;
assign w62 = ~w60 & ~w61;
assign w63 = (w38 & w1995) | (w38 & w1996) | (w1995 & w1996);
assign w64 = (~w38 & w1997) | (~w38 & w1998) | (w1997 & w1998);
assign w65 = ~w63 & ~w64;
assign w66 = (w38 & w1271) | (w38 & w1272) | (w1271 & w1272);
assign w67 = ~a_10 & ~b_10;
assign w68 = a_10 & b_10;
assign w69 = ~w67 & ~w68;
assign w70 = w66 & ~w69;
assign w71 = ~w66 & w69;
assign w72 = ~w70 & ~w71;
assign w73 = (w38 & w1273) | (w38 & w1274) | (w1273 & w1274);
assign w74 = ~a_11 & ~b_11;
assign w75 = a_11 & b_11;
assign w76 = ~w74 & ~w75;
assign w77 = w73 & ~w76;
assign w78 = ~w73 & w76;
assign w79 = ~w77 & ~w78;
assign w80 = (~w38 & w1887) | (~w38 & w1888) | (w1887 & w1888);
assign w81 = (w38 & w1999) | (w38 & w2000) | (w1999 & w2000);
assign w82 = ~a_12 & ~b_12;
assign w83 = a_12 & b_12;
assign w84 = ~w82 & ~w83;
assign w85 = w81 & ~w84;
assign w86 = ~w81 & w84;
assign w87 = ~w85 & ~w86;
assign w88 = ~a_13 & ~b_13;
assign w89 = a_13 & b_13;
assign w90 = ~w88 & ~w89;
assign w91 = ~w90 & w2937;
assign w92 = (w59 & w2001) | (w59 & w2002) | (w2001 & w2002);
assign w93 = ~w91 & ~w92;
assign w94 = ~a_14 & ~b_14;
assign w95 = a_14 & b_14;
assign w96 = ~w94 & ~w95;
assign w97 = ~w96 & w2788;
assign w98 = (w59 & w2003) | (w59 & w2004) | (w2003 & w2004);
assign w99 = ~w97 & ~w98;
assign w100 = (~w80 & w843) | (~w80 & w844) | (w843 & w844);
assign w101 = ~a_15 & ~b_15;
assign w102 = a_15 & b_15;
assign w103 = ~w101 & ~w102;
assign w104 = (~w80 & w1279) | (~w80 & w1280) | (w1279 & w1280);
assign w105 = (w80 & w1281) | (w80 & w1282) | (w1281 & w1282);
assign w106 = ~w104 & ~w105;
assign w107 = ~a_16 & ~b_16;
assign w108 = a_16 & b_16;
assign w109 = ~w107 & ~w108;
assign w110 = ~w109 & w2938;
assign w111 = (w80 & w2005) | (w80 & w2006) | (w2005 & w2006);
assign w112 = ~w110 & ~w111;
assign w113 = ~a_17 & ~b_17;
assign w114 = a_17 & b_17;
assign w115 = ~w113 & ~w114;
assign w116 = (~w80 & w2007) | (~w80 & w2008) | (w2007 & w2008);
assign w117 = (w80 & w2009) | (w80 & w2010) | (w2009 & w2010);
assign w118 = ~w116 & ~w117;
assign w119 = ~a_18 & ~b_18;
assign w120 = a_18 & b_18;
assign w121 = ~w119 & ~w120;
assign w122 = ~w121 & w2789;
assign w123 = (w80 & w2011) | (w80 & w2012) | (w2011 & w2012);
assign w124 = ~w122 & ~w123;
assign w125 = (~w80 & w1889) | (~w80 & w1890) | (w1889 & w1890);
assign w126 = ~a_19 & ~b_19;
assign w127 = a_19 & b_19;
assign w128 = ~w126 & ~w127;
assign w129 = (w1288 & w1287) | (w1288 & w100) | (w1287 & w100);
assign w130 = (w80 & w2013) | (w80 & w2014) | (w2013 & w2014);
assign w131 = ~w129 & ~w130;
assign w132 = (w1292 & w1291) | (w1292 & w100) | (w1291 & w100);
assign w133 = ~a_20 & ~b_20;
assign w134 = a_20 & b_20;
assign w135 = ~w133 & ~w134;
assign w136 = w132 & ~w135;
assign w137 = ~w132 & w135;
assign w138 = ~w136 & ~w137;
assign w139 = (w1294 & w1293) | (w1294 & w100) | (w1293 & w100);
assign w140 = ~a_21 & ~b_21;
assign w141 = a_21 & b_21;
assign w142 = ~w140 & ~w141;
assign w143 = w139 & ~w142;
assign w144 = ~w139 & w142;
assign w145 = ~w143 & ~w144;
assign w146 = ~a_22 & ~b_22;
assign w147 = a_22 & b_22;
assign w148 = ~w146 & ~w147;
assign w149 = (w100 & w2015) | (w100 & w2016) | (w2015 & w2016);
assign w150 = (~w100 & w2017) | (~w100 & w2018) | (w2017 & w2018);
assign w151 = ~w149 & ~w150;
assign w152 = ~a_23 & ~b_23;
assign w153 = a_23 & b_23;
assign w154 = ~w152 & ~w153;
assign w155 = (w100 & w2019) | (w100 & w2020) | (w2019 & w2020);
assign w156 = w154 & w2939;
assign w157 = ~w155 & ~w156;
assign w158 = ~a_24 & ~b_24;
assign w159 = a_24 & b_24;
assign w160 = ~w158 & ~w159;
assign w161 = (w125 & w2021) | (w125 & w2022) | (w2021 & w2022);
assign w162 = (~w125 & w2023) | (~w125 & w2024) | (w2023 & w2024);
assign w163 = ~w161 & ~w162;
assign w164 = ~a_25 & ~b_25;
assign w165 = a_25 & b_25;
assign w166 = ~w164 & ~w165;
assign w167 = (w125 & w2025) | (w125 & w2026) | (w2025 & w2026);
assign w168 = w166 & w2790;
assign w169 = ~w167 & ~w168;
assign w170 = ~a_26 & ~b_26;
assign w171 = a_26 & b_26;
assign w172 = ~w170 & ~w171;
assign w173 = (w125 & w2027) | (w125 & w2028) | (w2027 & w2028);
assign w174 = (w2445 & w2708) | (w2445 & w2792) | (w2708 & w2792);
assign w175 = ~w173 & ~w174;
assign w176 = ~a_27 & ~b_27;
assign w177 = a_27 & b_27;
assign w178 = ~w176 & ~w177;
assign w179 = (w125 & w2029) | (w125 & w2030) | (w2029 & w2030);
assign w180 = (~w125 & w2031) | (~w125 & w2032) | (w2031 & w2032);
assign w181 = ~w179 & ~w180;
assign w182 = ~a_28 & ~b_28;
assign w183 = a_28 & b_28;
assign w184 = ~w182 & ~w183;
assign w185 = (w125 & w2033) | (w125 & w2034) | (w2033 & w2034);
assign w186 = w184 & w2791;
assign w187 = ~w185 & ~w186;
assign w188 = ~a_29 & ~b_29;
assign w189 = a_29 & b_29;
assign w190 = ~w188 & ~w189;
assign w191 = (w125 & w2628) | (w125 & w2629) | (w2628 & w2629);
assign w192 = w190 & w2793;
assign w193 = ~w191 & ~w192;
assign w194 = (w125 & w2037) | (w125 & w2038) | (w2037 & w2038);
assign w195 = ~a_30 & ~b_30;
assign w196 = a_30 & b_30;
assign w197 = ~w195 & ~w196;
assign w198 = w194 & ~w197;
assign w199 = ~w194 & w197;
assign w200 = ~w198 & ~w199;
assign w201 = (w125 & w2039) | (w125 & w2040) | (w2039 & w2040);
assign w202 = ~a_31 & ~b_31;
assign w203 = a_31 & b_31;
assign w204 = ~w202 & ~w203;
assign w205 = w201 & ~w204;
assign w206 = ~w201 & w204;
assign w207 = ~w205 & ~w206;
assign w208 = (w125 & w2041) | (w125 & w2042) | (w2041 & w2042);
assign w209 = ~a_32 & ~b_32;
assign w210 = a_32 & b_32;
assign w211 = ~w209 & ~w210;
assign w212 = w208 & ~w211;
assign w213 = ~w208 & w211;
assign w214 = ~w212 & ~w213;
assign w215 = (w125 & w2043) | (w125 & w2044) | (w2043 & w2044);
assign w216 = ~a_33 & ~b_33;
assign w217 = a_33 & b_33;
assign w218 = ~w216 & ~w217;
assign w219 = w215 & ~w218;
assign w220 = ~w215 & w218;
assign w221 = ~w219 & ~w220;
assign w222 = (w125 & w2045) | (w125 & w2046) | (w2045 & w2046);
assign w223 = ~a_34 & ~b_34;
assign w224 = a_34 & b_34;
assign w225 = ~w223 & ~w224;
assign w226 = (w125 & w2047) | (w125 & w2048) | (w2047 & w2048);
assign w227 = (w1310 & w1309) | (w1310 & w2794) | (w1309 & w2794);
assign w228 = ~w226 & ~w227;
assign w229 = (w125 & w2049) | (w125 & w2050) | (w2049 & w2050);
assign w230 = ~a_35 & ~b_35;
assign w231 = a_35 & b_35;
assign w232 = ~w230 & ~w231;
assign w233 = w229 & ~w232;
assign w234 = ~w229 & w232;
assign w235 = ~w233 & ~w234;
assign w236 = (w125 & w2051) | (w125 & w2052) | (w2051 & w2052);
assign w237 = ~a_36 & ~b_36;
assign w238 = a_36 & b_36;
assign w239 = ~w237 & ~w238;
assign w240 = w236 & ~w239;
assign w241 = ~w236 & w239;
assign w242 = ~w240 & ~w241;
assign w243 = (w125 & w2053) | (w125 & w2054) | (w2053 & w2054);
assign w244 = ~a_37 & ~b_37;
assign w245 = a_37 & b_37;
assign w246 = ~w244 & ~w245;
assign w247 = w243 & ~w246;
assign w248 = ~w243 & w246;
assign w249 = ~w247 & ~w248;
assign w250 = ~a_38 & ~b_38;
assign w251 = a_38 & b_38;
assign w252 = ~w250 & ~w251;
assign w253 = ~w252 & w2795;
assign w254 = (w2794 & w2055) | (w2794 & w2056) | (w2055 & w2056);
assign w255 = ~w253 & ~w254;
assign w256 = ~a_39 & ~b_39;
assign w257 = a_39 & b_39;
assign w258 = ~w256 & ~w257;
assign w259 = ~w258 & w2796;
assign w260 = (w2794 & w2057) | (w2794 & w2058) | (w2057 & w2058);
assign w261 = ~w259 & ~w260;
assign w262 = (w125 & w2622) | (w125 & w2623) | (w2622 & w2623);
assign w263 = ~a_40 & ~b_40;
assign w264 = a_40 & b_40;
assign w265 = ~w263 & ~w264;
assign w266 = (w222 & w1319) | (w222 & w1320) | (w1319 & w1320);
assign w267 = (~w222 & w1321) | (~w222 & w1322) | (w1321 & w1322);
assign w268 = ~w266 & ~w267;
assign w269 = ~a_41 & ~b_41;
assign w270 = a_41 & b_41;
assign w271 = ~w269 & ~w270;
assign w272 = (w222 & w2059) | (w222 & w2060) | (w2059 & w2060);
assign w273 = w271 & w2797;
assign w274 = ~w272 & ~w273;
assign w275 = ~a_42 & ~b_42;
assign w276 = a_42 & b_42;
assign w277 = ~w275 & ~w276;
assign w278 = (w222 & w2061) | (w222 & w2062) | (w2061 & w2062);
assign w279 = (~w222 & w2063) | (~w222 & w2064) | (w2063 & w2064);
assign w280 = ~w278 & ~w279;
assign w281 = ~a_43 & ~b_43;
assign w282 = a_43 & b_43;
assign w283 = ~w281 & ~w282;
assign w284 = (w222 & w2065) | (w222 & w2066) | (w2065 & w2066);
assign w285 = w283 & w2798;
assign w286 = ~w284 & ~w285;
assign w287 = ~a_44 & ~b_44;
assign w288 = a_44 & b_44;
assign w289 = ~w287 & ~w288;
assign w290 = (w222 & w2067) | (w222 & w2068) | (w2067 & w2068);
assign w291 = w289 & w2799;
assign w292 = ~w290 & ~w291;
assign w293 = ~a_45 & ~b_45;
assign w294 = a_45 & b_45;
assign w295 = ~w293 & ~w294;
assign w296 = (w222 & w2069) | (w222 & w2070) | (w2069 & w2070);
assign w297 = w295 & w2800;
assign w298 = ~w296 & ~w297;
assign w299 = ~a_46 & ~b_46;
assign w300 = a_46 & b_46;
assign w301 = ~w299 & ~w300;
assign w302 = (w222 & w2071) | (w222 & w2072) | (w2071 & w2072);
assign w303 = w301 & w2801;
assign w304 = ~w302 & ~w303;
assign w305 = (w2794 & w2073) | (w2794 & w2074) | (w2073 & w2074);
assign w306 = ~a_47 & ~b_47;
assign w307 = a_47 & b_47;
assign w308 = ~w306 & ~w307;
assign w309 = (w2738 & w2739) | (w2738 & w2802) | (w2739 & w2802);
assign w310 = (w2794 & w2630) | (w2794 & w2631) | (w2630 & w2631);
assign w311 = ~w309 & ~w310;
assign w312 = ~a_48 & ~b_48;
assign w313 = a_48 & b_48;
assign w314 = ~w312 & ~w313;
assign w315 = ~w314 & w2803;
assign w316 = (w2794 & w2632) | (w2794 & w2633) | (w2632 & w2633);
assign w317 = ~w315 & ~w316;
assign w318 = ~a_49 & ~b_49;
assign w319 = a_49 & b_49;
assign w320 = ~w318 & ~w319;
assign w321 = ~w320 & w2804;
assign w322 = (w2794 & w2634) | (w2794 & w2635) | (w2634 & w2635);
assign w323 = ~w321 & ~w322;
assign w324 = ~a_50 & ~b_50;
assign w325 = a_50 & b_50;
assign w326 = ~w324 & ~w325;
assign w327 = ~w326 & w2805;
assign w328 = (w2794 & w2636) | (w2794 & w2637) | (w2636 & w2637);
assign w329 = ~w327 & ~w328;
assign w330 = (~w2794 & w2081) | (~w2794 & w2082) | (w2081 & w2082);
assign w331 = ~a_51 & ~b_51;
assign w332 = a_51 & b_51;
assign w333 = ~w331 & ~w332;
assign w334 = w330 & ~w333;
assign w335 = ~w330 & w333;
assign w336 = ~w334 & ~w335;
assign w337 = ~a_52 & ~b_52;
assign w338 = a_52 & b_52;
assign w339 = ~w337 & ~w338;
assign w340 = ~w339 & w2806;
assign w341 = (w2794 & w2638) | (w2794 & w2639) | (w2638 & w2639);
assign w342 = ~w340 & ~w341;
assign w343 = (~w2794 & w2085) | (~w2794 & w2086) | (w2085 & w2086);
assign w344 = ~a_53 & ~b_53;
assign w345 = a_53 & b_53;
assign w346 = ~w344 & ~w345;
assign w347 = w343 & ~w346;
assign w348 = ~w343 & w346;
assign w349 = ~w347 & ~w348;
assign w350 = (w2794 & w2087) | (w2794 & w2088) | (w2087 & w2088);
assign w351 = ~a_54 & ~b_54;
assign w352 = a_54 & b_54;
assign w353 = ~w351 & ~w352;
assign w354 = (w2089 & w2090) | (w2089 & ~w305) | (w2090 & ~w305);
assign w355 = (w2794 & w2640) | (w2794 & w2641) | (w2640 & w2641);
assign w356 = ~w354 & ~w355;
assign w357 = ~a_55 & ~b_55;
assign w358 = a_55 & b_55;
assign w359 = ~w357 & ~w358;
assign w360 = (w2093 & w2094) | (w2093 & ~w305) | (w2094 & ~w305);
assign w361 = (w2794 & w2642) | (w2794 & w2643) | (w2642 & w2643);
assign w362 = ~w360 & ~w361;
assign w363 = ~a_56 & ~b_56;
assign w364 = a_56 & b_56;
assign w365 = ~w363 & ~w364;
assign w366 = (w2098 & w2097) | (w2098 & ~w305) | (w2097 & ~w305);
assign w367 = (w2794 & w2644) | (w2794 & w2645) | (w2644 & w2645);
assign w368 = ~w366 & ~w367;
assign w369 = ~a_57 & ~b_57;
assign w370 = a_57 & b_57;
assign w371 = ~w369 & ~w370;
assign w372 = (w2100 & w2099) | (w2100 & ~w305) | (w2099 & ~w305);
assign w373 = (w2794 & w2646) | (w2794 & w2647) | (w2646 & w2647);
assign w374 = ~w372 & ~w373;
assign w375 = ~a_58 & ~b_58;
assign w376 = a_58 & b_58;
assign w377 = ~w375 & ~w376;
assign w378 = (~w305 & w2101) | (~w305 & w2102) | (w2101 & w2102);
assign w379 = (w305 & w2103) | (w305 & w2104) | (w2103 & w2104);
assign w380 = ~w378 & ~w379;
assign w381 = ~a_59 & ~b_59;
assign w382 = a_59 & b_59;
assign w383 = ~w381 & ~w382;
assign w384 = (w2106 & w2105) | (w2106 & ~w305) | (w2105 & ~w305);
assign w385 = (w2794 & w2751) | (w2794 & w2752) | (w2751 & w2752);
assign w386 = ~w384 & ~w385;
assign w387 = ~a_60 & ~b_60;
assign w388 = a_60 & b_60;
assign w389 = ~w387 & ~w388;
assign w390 = (~w305 & w2107) | (~w305 & w2108) | (w2107 & w2108);
assign w391 = (w305 & w2109) | (w305 & w2110) | (w2109 & w2110);
assign w392 = ~w390 & ~w391;
assign w393 = (w262 & w1897) | (w262 & w1898) | (w1897 & w1898);
assign w394 = ~a_61 & ~b_61;
assign w395 = a_61 & b_61;
assign w396 = ~w394 & ~w395;
assign w397 = (~w350 & w1351) | (~w350 & w1352) | (w1351 & w1352);
assign w398 = (w350 & w1353) | (w350 & w1354) | (w1353 & w1354);
assign w399 = ~w397 & ~w398;
assign w400 = ~a_62 & ~b_62;
assign w401 = a_62 & b_62;
assign w402 = ~w400 & ~w401;
assign w403 = (~w350 & w2111) | (~w350 & w2112) | (w2111 & w2112);
assign w404 = (w350 & w2113) | (w350 & w2114) | (w2113 & w2114);
assign w405 = ~w403 & ~w404;
assign w406 = ~a_63 & ~b_63;
assign w407 = a_63 & b_63;
assign w408 = ~w406 & ~w407;
assign w409 = (~w350 & w2115) | (~w350 & w2116) | (w2115 & w2116);
assign w410 = (w350 & w2117) | (w350 & w2118) | (w2117 & w2118);
assign w411 = ~w409 & ~w410;
assign w412 = ~a_64 & ~b_64;
assign w413 = a_64 & b_64;
assign w414 = ~w412 & ~w413;
assign w415 = (~w350 & w2119) | (~w350 & w2120) | (w2119 & w2120);
assign w416 = (w350 & w2121) | (w350 & w2122) | (w2121 & w2122);
assign w417 = ~w415 & ~w416;
assign w418 = ~a_65 & ~b_65;
assign w419 = a_65 & b_65;
assign w420 = ~w418 & ~w419;
assign w421 = (~w350 & w2123) | (~w350 & w2124) | (w2123 & w2124);
assign w422 = (w350 & w2125) | (w350 & w2126) | (w2125 & w2126);
assign w423 = ~w421 & ~w422;
assign w424 = ~a_66 & ~b_66;
assign w425 = a_66 & b_66;
assign w426 = ~w424 & ~w425;
assign w427 = (~w350 & w2127) | (~w350 & w2128) | (w2127 & w2128);
assign w428 = (w350 & w2129) | (w350 & w2130) | (w2129 & w2130);
assign w429 = ~w427 & ~w428;
assign w430 = ~a_67 & ~b_67;
assign w431 = a_67 & b_67;
assign w432 = ~w430 & ~w431;
assign w433 = (~w350 & w2131) | (~w350 & w2132) | (w2131 & w2132);
assign w434 = (w350 & w2133) | (w350 & w2134) | (w2133 & w2134);
assign w435 = ~w433 & ~w434;
assign w436 = ~a_68 & ~b_68;
assign w437 = a_68 & b_68;
assign w438 = ~w436 & ~w437;
assign w439 = (~w350 & w2135) | (~w350 & w2136) | (w2135 & w2136);
assign w440 = (w350 & w2137) | (w350 & w2138) | (w2137 & w2138);
assign w441 = ~w439 & ~w440;
assign w442 = (w262 & w1927) | (w262 & w1928) | (w1927 & w1928);
assign w443 = ~a_69 & ~b_69;
assign w444 = a_69 & b_69;
assign w445 = ~w443 & ~w444;
assign w446 = (w262 & w2139) | (w262 & w2140) | (w2139 & w2140);
assign w447 = (w2476 & w2477) | (w2476 & w2807) | (w2477 & w2807);
assign w448 = ~w446 & ~w447;
assign w449 = (w262 & w2141) | (w262 & w2142) | (w2141 & w2142);
assign w450 = ~a_70 & ~b_70;
assign w451 = a_70 & b_70;
assign w452 = ~w450 & ~w451;
assign w453 = w449 & ~w452;
assign w454 = ~w449 & w452;
assign w455 = ~w453 & ~w454;
assign w456 = (w262 & w2143) | (w262 & w2144) | (w2143 & w2144);
assign w457 = ~a_71 & ~b_71;
assign w458 = a_71 & b_71;
assign w459 = ~w457 & ~w458;
assign w460 = w456 & ~w459;
assign w461 = ~w456 & w459;
assign w462 = ~w460 & ~w461;
assign w463 = (w262 & w2145) | (w262 & w2146) | (w2145 & w2146);
assign w464 = ~a_72 & ~b_72;
assign w465 = a_72 & b_72;
assign w466 = ~w464 & ~w465;
assign w467 = w463 & ~w466;
assign w468 = ~w463 & w466;
assign w469 = ~w467 & ~w468;
assign w470 = (w262 & w2147) | (w262 & w2148) | (w2147 & w2148);
assign w471 = ~a_73 & ~b_73;
assign w472 = a_73 & b_73;
assign w473 = ~w471 & ~w472;
assign w474 = w470 & ~w473;
assign w475 = ~w470 & w473;
assign w476 = ~w474 & ~w475;
assign w477 = (w262 & w2149) | (w262 & w2150) | (w2149 & w2150);
assign w478 = ~a_74 & ~b_74;
assign w479 = a_74 & b_74;
assign w480 = ~w478 & ~w479;
assign w481 = w477 & ~w480;
assign w482 = ~w477 & w480;
assign w483 = ~w481 & ~w482;
assign w484 = (w262 & w2151) | (w262 & w2152) | (w2151 & w2152);
assign w485 = ~a_75 & ~b_75;
assign w486 = a_75 & b_75;
assign w487 = ~w485 & ~w486;
assign w488 = w484 & ~w487;
assign w489 = ~w484 & w487;
assign w490 = ~w488 & ~w489;
assign w491 = (w262 & w2153) | (w262 & w2154) | (w2153 & w2154);
assign w492 = ~a_76 & ~b_76;
assign w493 = a_76 & b_76;
assign w494 = ~w492 & ~w493;
assign w495 = w491 & ~w494;
assign w496 = ~w491 & w494;
assign w497 = ~w495 & ~w496;
assign w498 = (w262 & w2155) | (w262 & w2156) | (w2155 & w2156);
assign w499 = ~a_77 & ~b_77;
assign w500 = a_77 & b_77;
assign w501 = ~w499 & ~w500;
assign w502 = w498 & ~w501;
assign w503 = ~w498 & w501;
assign w504 = ~w502 & ~w503;
assign w505 = (~w262 & w1929) | (~w262 & w1930) | (w1929 & w1930);
assign w506 = ~a_78 & ~b_78;
assign w507 = a_78 & b_78;
assign w508 = ~w506 & ~w507;
assign w509 = (w442 & w2157) | (w442 & w2158) | (w2157 & w2158);
assign w510 = (~w442 & w2159) | (~w442 & w2160) | (w2159 & w2160);
assign w511 = ~w509 & ~w510;
assign w512 = ~a_79 & ~b_79;
assign w513 = a_79 & b_79;
assign w514 = ~w512 & ~w513;
assign w515 = (w442 & w2161) | (w442 & w2162) | (w2161 & w2162);
assign w516 = (~w442 & w2163) | (~w442 & w2164) | (w2163 & w2164);
assign w517 = ~w515 & ~w516;
assign w518 = ~a_80 & ~b_80;
assign w519 = a_80 & b_80;
assign w520 = ~w518 & ~w519;
assign w521 = (w442 & w2165) | (w442 & w2166) | (w2165 & w2166);
assign w522 = (~w442 & w2167) | (~w442 & w2168) | (w2167 & w2168);
assign w523 = ~w521 & ~w522;
assign w524 = ~a_81 & ~b_81;
assign w525 = a_81 & b_81;
assign w526 = ~w524 & ~w525;
assign w527 = (w442 & w2169) | (w442 & w2170) | (w2169 & w2170);
assign w528 = w526 & w2940;
assign w529 = ~w527 & ~w528;
assign w530 = ~a_82 & ~b_82;
assign w531 = a_82 & b_82;
assign w532 = ~w530 & ~w531;
assign w533 = (w442 & w2171) | (w442 & w2172) | (w2171 & w2172);
assign w534 = w532 & w2808;
assign w535 = ~w533 & ~w534;
assign w536 = ~a_83 & ~b_83;
assign w537 = a_83 & b_83;
assign w538 = ~w536 & ~w537;
assign w539 = (w442 & w2173) | (w442 & w2174) | (w2173 & w2174);
assign w540 = w538 & w2809;
assign w541 = ~w539 & ~w540;
assign w542 = ~a_84 & ~b_84;
assign w543 = a_84 & b_84;
assign w544 = ~w542 & ~w543;
assign w545 = (w442 & w2175) | (w442 & w2176) | (w2175 & w2176);
assign w546 = (~w442 & w2177) | (~w442 & w2178) | (w2177 & w2178);
assign w547 = ~w545 & ~w546;
assign w548 = ~a_85 & ~b_85;
assign w549 = a_85 & b_85;
assign w550 = ~w548 & ~w549;
assign w551 = (w442 & w2179) | (w442 & w2180) | (w2179 & w2180);
assign w552 = (~w442 & w2181) | (~w442 & w2182) | (w2181 & w2182);
assign w553 = ~w551 & ~w552;
assign w554 = ~a_86 & ~b_86;
assign w555 = a_86 & b_86;
assign w556 = ~w554 & ~w555;
assign w557 = (w442 & w2183) | (w442 & w2184) | (w2183 & w2184);
assign w558 = (~w442 & w2185) | (~w442 & w2186) | (w2185 & w2186);
assign w559 = ~w557 & ~w558;
assign w560 = (~w393 & w1901) | (~w393 & w1902) | (w1901 & w1902);
assign w561 = ~a_87 & ~b_87;
assign w562 = a_87 & b_87;
assign w563 = ~w561 & ~w562;
assign w564 = (~w505 & w2187) | (~w505 & w2188) | (w2187 & w2188);
assign w565 = (w505 & w2189) | (w505 & w2190) | (w2189 & w2190);
assign w566 = ~w564 & ~w565;
assign w567 = ~a_88 & ~b_88;
assign w568 = a_88 & b_88;
assign w569 = ~w567 & ~w568;
assign w570 = (~w505 & w2191) | (~w505 & w2192) | (w2191 & w2192);
assign w571 = (w505 & w2193) | (w505 & w2194) | (w2193 & w2194);
assign w572 = ~w570 & ~w571;
assign w573 = ~a_89 & ~b_89;
assign w574 = a_89 & b_89;
assign w575 = ~w573 & ~w574;
assign w576 = (~w505 & w2195) | (~w505 & w2196) | (w2195 & w2196);
assign w577 = (w505 & w2197) | (w505 & w2198) | (w2197 & w2198);
assign w578 = ~w576 & ~w577;
assign w579 = ~a_90 & ~b_90;
assign w580 = a_90 & b_90;
assign w581 = ~w579 & ~w580;
assign w582 = (~w505 & w2199) | (~w505 & w2200) | (w2199 & w2200);
assign w583 = (w505 & w2201) | (w505 & w2202) | (w2201 & w2202);
assign w584 = ~w582 & ~w583;
assign w585 = ~a_91 & ~b_91;
assign w586 = a_91 & b_91;
assign w587 = ~w585 & ~w586;
assign w588 = (~w505 & w2203) | (~w505 & w2204) | (w2203 & w2204);
assign w589 = (w505 & w2205) | (w505 & w2206) | (w2205 & w2206);
assign w590 = ~w588 & ~w589;
assign w591 = ~a_92 & ~b_92;
assign w592 = a_92 & b_92;
assign w593 = ~w591 & ~w592;
assign w594 = (~w505 & w2207) | (~w505 & w2208) | (w2207 & w2208);
assign w595 = (w505 & w2209) | (w505 & w2210) | (w2209 & w2210);
assign w596 = ~w594 & ~w595;
assign w597 = ~a_93 & ~b_93;
assign w598 = a_93 & b_93;
assign w599 = ~w597 & ~w598;
assign w600 = (~w505 & w2211) | (~w505 & w2212) | (w2211 & w2212);
assign w601 = (w505 & w2213) | (w505 & w2214) | (w2213 & w2214);
assign w602 = ~w600 & ~w601;
assign w603 = ~a_94 & ~b_94;
assign w604 = a_94 & b_94;
assign w605 = ~w603 & ~w604;
assign w606 = (~w505 & w2215) | (~w505 & w2216) | (w2215 & w2216);
assign w607 = (w505 & w2217) | (w505 & w2218) | (w2217 & w2218);
assign w608 = ~w606 & ~w607;
assign w609 = ~a_95 & ~b_95;
assign w610 = a_95 & b_95;
assign w611 = ~w609 & ~w610;
assign w612 = (~w505 & w2219) | (~w505 & w2220) | (w2219 & w2220);
assign w613 = (w505 & w2221) | (w505 & w2222) | (w2221 & w2222);
assign w614 = ~w612 & ~w613;
assign w615 = (w393 & w1931) | (w393 & w1932) | (w1931 & w1932);
assign w616 = ~a_96 & ~b_96;
assign w617 = a_96 & b_96;
assign w618 = ~w616 & ~w617;
assign w619 = (w393 & w2223) | (w393 & w2224) | (w2223 & w2224);
assign w620 = (w2526 & w2527) | (w2526 & w2810) | (w2527 & w2810);
assign w621 = ~w619 & ~w620;
assign w622 = ~a_97 & ~b_97;
assign w623 = a_97 & b_97;
assign w624 = ~w622 & ~w623;
assign w625 = (w393 & w2753) | (w393 & w2754) | (w2753 & w2754);
assign w626 = w624 & w2811;
assign w627 = ~w625 & ~w626;
assign w628 = ~a_98 & ~b_98;
assign w629 = a_98 & b_98;
assign w630 = ~w628 & ~w629;
assign w631 = (w393 & w2755) | (w393 & w2756) | (w2755 & w2756);
assign w632 = w630 & w2812;
assign w633 = ~w631 & ~w632;
assign w634 = (w393 & w1937) | (w393 & w1938) | (w1937 & w1938);
assign w635 = ~a_99 & ~b_99;
assign w636 = a_99 & b_99;
assign w637 = ~w635 & ~w636;
assign w638 = w634 & ~w637;
assign w639 = ~w634 & w637;
assign w640 = ~w638 & ~w639;
assign w641 = (w393 & w1939) | (w393 & w1940) | (w1939 & w1940);
assign w642 = ~a_100 & ~b_100;
assign w643 = a_100 & b_100;
assign w644 = ~w642 & ~w643;
assign w645 = w641 & ~w644;
assign w646 = ~w641 & w644;
assign w647 = ~w645 & ~w646;
assign w648 = (w393 & w1941) | (w393 & w1942) | (w1941 & w1942);
assign w649 = ~a_101 & ~b_101;
assign w650 = a_101 & b_101;
assign w651 = ~w649 & ~w650;
assign w652 = w648 & ~w651;
assign w653 = ~w648 & w651;
assign w654 = ~w652 & ~w653;
assign w655 = (w393 & w1943) | (w393 & w1944) | (w1943 & w1944);
assign w656 = ~a_102 & ~b_102;
assign w657 = a_102 & b_102;
assign w658 = ~w656 & ~w657;
assign w659 = w655 & ~w658;
assign w660 = ~w655 & w658;
assign w661 = ~w659 & ~w660;
assign w662 = ~a_103 & ~b_103;
assign w663 = a_103 & b_103;
assign w664 = ~w662 & ~w663;
assign w665 = (w393 & w2648) | (w393 & w2649) | (w2648 & w2649);
assign w666 = (w1948 & w1947) | (w1948 & w560) | (w1947 & w560);
assign w667 = ~w665 & ~w666;
assign w668 = ~a_104 & ~b_104;
assign w669 = a_104 & b_104;
assign w670 = ~w668 & ~w669;
assign w671 = (w393 & w2650) | (w393 & w2651) | (w2650 & w2651);
assign w672 = (w1952 & w1951) | (w1952 & w560) | (w1951 & w560);
assign w673 = ~w671 & ~w672;
assign w674 = ~a_105 & ~b_105;
assign w675 = a_105 & b_105;
assign w676 = ~w674 & ~w675;
assign w677 = (w393 & w2757) | (w393 & w2758) | (w2757 & w2758);
assign w678 = (w1956 & w1955) | (w1956 & w560) | (w1955 & w560);
assign w679 = ~w677 & ~w678;
assign w680 = (w393 & w2759) | (w393 & w2760) | (w2759 & w2760);
assign w681 = ~a_106 & ~b_106;
assign w682 = a_106 & b_106;
assign w683 = ~w681 & ~w682;
assign w684 = (~w560 & w1957) | (~w560 & w1958) | (w1957 & w1958);
assign w685 = (w560 & w1959) | (w560 & w1960) | (w1959 & w1960);
assign w686 = ~w684 & ~w685;
assign w687 = ~a_107 & ~b_107;
assign w688 = a_107 & b_107;
assign w689 = ~w687 & ~w688;
assign w690 = (w393 & w2761) | (w393 & w2762) | (w2761 & w2762);
assign w691 = (w1223 & w1224) | (w1223 & ~w615) | (w1224 & ~w615);
assign w692 = ~w690 & ~w691;
assign w693 = ~a_108 & ~b_108;
assign w694 = a_108 & b_108;
assign w695 = ~w693 & ~w694;
assign w696 = (w393 & w2763) | (w393 & w2764) | (w2763 & w2764);
assign w697 = (w1228 & w1227) | (w1228 & ~w615) | (w1227 & ~w615);
assign w698 = ~w696 & ~w697;
assign w699 = ~a_109 & ~b_109;
assign w700 = a_109 & b_109;
assign w701 = ~w699 & ~w700;
assign w702 = (w393 & w2765) | (w393 & w2766) | (w2765 & w2766);
assign w703 = (w1232 & w1231) | (w1232 & ~w615) | (w1231 & ~w615);
assign w704 = ~w702 & ~w703;
assign w705 = ~a_110 & ~b_110;
assign w706 = a_110 & b_110;
assign w707 = ~w705 & ~w706;
assign w708 = (w393 & w2767) | (w393 & w2768) | (w2767 & w2768);
assign w709 = (w1235 & w1236) | (w1235 & ~w615) | (w1236 & ~w615);
assign w710 = ~w708 & ~w709;
assign w711 = ~a_111 & ~b_111;
assign w712 = a_111 & b_111;
assign w713 = ~w711 & ~w712;
assign w714 = (w393 & w2769) | (w393 & w2770) | (w2769 & w2770);
assign w715 = (w1240 & w1239) | (w1240 & ~w615) | (w1239 & ~w615);
assign w716 = ~w714 & ~w715;
assign w717 = ~a_112 & ~b_112;
assign w718 = a_112 & b_112;
assign w719 = ~w717 & ~w718;
assign w720 = (w393 & w2771) | (w393 & w2772) | (w2771 & w2772);
assign w721 = (w1243 & w1244) | (w1243 & ~w615) | (w1244 & ~w615);
assign w722 = ~w720 & ~w721;
assign w723 = ~a_113 & ~b_113;
assign w724 = a_113 & b_113;
assign w725 = ~w723 & ~w724;
assign w726 = (w615 & w1245) | (w615 & w1246) | (w1245 & w1246);
assign w727 = (~w615 & w1247) | (~w615 & w1248) | (w1247 & w1248);
assign w728 = ~w726 & ~w727;
assign w729 = ~a_114 & ~b_114;
assign w730 = a_114 & b_114;
assign w731 = ~w729 & ~w730;
assign w732 = (w393 & w2773) | (w393 & w2774) | (w2773 & w2774);
assign w733 = (w1252 & w1251) | (w1252 & ~w615) | (w1251 & ~w615);
assign w734 = ~w732 & ~w733;
assign w735 = ~a_115 & ~b_115;
assign w736 = a_115 & b_115;
assign w737 = ~w735 & ~w736;
assign w738 = (w393 & w2775) | (w393 & w2776) | (w2775 & w2776);
assign w739 = (w1256 & w1255) | (w1256 & ~w615) | (w1255 & ~w615);
assign w740 = ~w738 & ~w739;
assign w741 = ~a_116 & ~b_116;
assign w742 = a_116 & b_116;
assign w743 = ~w741 & ~w742;
assign w744 = (w615 & w1257) | (w615 & w1258) | (w1257 & w1258);
assign w745 = (~w615 & w1259) | (~w615 & w1260) | (w1259 & w1260);
assign w746 = ~w744 & ~w745;
assign w747 = ~a_117 & ~b_117;
assign w748 = a_117 & b_117;
assign w749 = ~w747 & ~w748;
assign w750 = (~w560 & w1961) | (~w560 & w1962) | (w1961 & w1962);
assign w751 = (w560 & w1963) | (w560 & w1964) | (w1963 & w1964);
assign w752 = ~w750 & ~w751;
assign w753 = ~a_118 & ~b_118;
assign w754 = a_118 & b_118;
assign w755 = ~w753 & ~w754;
assign w756 = (~w560 & w1965) | (~w560 & w1966) | (w1965 & w1966);
assign w757 = (w560 & w1967) | (w560 & w1968) | (w1967 & w1968);
assign w758 = ~w756 & ~w757;
assign w759 = ~a_119 & ~b_119;
assign w760 = a_119 & b_119;
assign w761 = ~w759 & ~w760;
assign w762 = (~w560 & w1969) | (~w560 & w1970) | (w1969 & w1970);
assign w763 = (w560 & w1971) | (w560 & w1972) | (w1971 & w1972);
assign w764 = ~w762 & ~w763;
assign w765 = ~a_120 & ~b_120;
assign w766 = a_120 & b_120;
assign w767 = ~w765 & ~w766;
assign w768 = (~w560 & w1973) | (~w560 & w1974) | (w1973 & w1974);
assign w769 = (w560 & w1975) | (w560 & w1976) | (w1975 & w1976);
assign w770 = ~w768 & ~w769;
assign w771 = ~a_121 & ~b_121;
assign w772 = a_121 & b_121;
assign w773 = ~w771 & ~w772;
assign w774 = (~w560 & w1977) | (~w560 & w1978) | (w1977 & w1978);
assign w775 = (w560 & w1979) | (w560 & w1980) | (w1979 & w1980);
assign w776 = ~w774 & ~w775;
assign w777 = ~a_122 & ~b_122;
assign w778 = a_122 & b_122;
assign w779 = ~w777 & ~w778;
assign w780 = (~w560 & w1981) | (~w560 & w1982) | (w1981 & w1982);
assign w781 = (w560 & w1983) | (w560 & w1984) | (w1983 & w1984);
assign w782 = ~w780 & ~w781;
assign w783 = ~a_123 & ~b_123;
assign w784 = a_123 & b_123;
assign w785 = ~w783 & ~w784;
assign w786 = (~w560 & w1985) | (~w560 & w1986) | (w1985 & w1986);
assign w787 = (w560 & w1987) | (w560 & w1988) | (w1987 & w1988);
assign w788 = ~w786 & ~w787;
assign w789 = ~a_124 & ~b_124;
assign w790 = a_124 & b_124;
assign w791 = ~w789 & ~w790;
assign w792 = (~w560 & w1989) | (~w560 & w1990) | (w1989 & w1990);
assign w793 = (w560 & w1991) | (w560 & w1992) | (w1991 & w1992);
assign w794 = ~w792 & ~w793;
assign w795 = ~a_125 & ~b_125;
assign w796 = a_125 & b_125;
assign w797 = ~w795 & ~w796;
assign w798 = (w680 & w1191) | (w680 & w1192) | (w1191 & w1192);
assign w799 = (~w680 & w1193) | (~w680 & w1194) | (w1193 & w1194);
assign w800 = ~w798 & ~w799;
assign w801 = ~a_126 & ~b_126;
assign w802 = a_126 & b_126;
assign w803 = ~w801 & ~w802;
assign w804 = (~w560 & w1993) | (~w560 & w1994) | (w1993 & w1994);
assign w805 = (w560 & w2624) | (w560 & w2625) | (w2624 & w2625);
assign w806 = ~w804 & ~w805;
assign w807 = ~a_127 & ~b_127;
assign w808 = a_127 & b_127;
assign w809 = ~w807 & ~w808;
assign w810 = (w615 & w1903) | (w615 & w1904) | (w1903 & w1904);
assign w811 = (~w615 & w1905) | (~w615 & w1906) | (w1905 & w1906);
assign w812 = ~w810 & ~w811;
assign w813 = (~w615 & w1907) | (~w615 & w1908) | (w1907 & w1908);
assign w814 = ~w808 & ~w813;
assign w815 = w5 & ~w12;
assign w816 = w13 & ~w19;
assign w817 = ~w20 & w19;
assign w818 = ~w20 & ~w816;
assign w819 = w26 & ~w27;
assign w820 = ~w32 & w27;
assign w821 = ~w33 & ~w820;
assign w822 = (~w33 & w819) | (~w33 & w1122) | (w819 & w1122);
assign w823 = w39 & ~w40;
assign w824 = ~w46 & w40;
assign w825 = ~w47 & ~w824;
assign w826 = (~w47 & w823) | (~w47 & w1123) | (w823 & w1123);
assign w827 = (~w53 & w824) | (~w53 & w1405) | (w824 & w1405);
assign w828 = ~w53 & ~w826;
assign w829 = w54 & ~w60;
assign w830 = ~w61 & w60;
assign w831 = (~w67 & w829) | (~w67 & w1124) | (w829 & w1124);
assign w832 = (~w68 & w830) | (~w68 & w1406) | (w830 & w1406);
assign w833 = ~w68 & ~w831;
assign w834 = ~w74 & ~w832;
assign w835 = (~w74 & w831) | (~w74 & w1407) | (w831 & w1407);
assign w836 = w75 & ~w82;
assign w837 = ~w83 & w82;
assign w838 = ~w83 & ~w836;
assign w839 = (~w88 & w836) | (~w88 & w1125) | (w836 & w1125);
assign w840 = (~w89 & w837) | (~w89 & w1408) | (w837 & w1408);
assign w841 = ~w89 & ~w839;
assign w842 = (~w94 & w839) | (~w94 & w1409) | (w839 & w1409);
assign w843 = (~w95 & w840) | (~w95 & w1410) | (w840 & w1410);
assign w844 = ~w95 & ~w842;
assign w845 = w101 & ~w102;
assign w846 = ~w107 & w102;
assign w847 = ~w108 & ~w846;
assign w848 = (~w108 & w845) | (~w108 & w1126) | (w845 & w1126);
assign w849 = (~w113 & w846) | (~w113 & w1411) | (w846 & w1411);
assign w850 = ~w114 & ~w849;
assign w851 = (~w114 & w848) | (~w114 & w1412) | (w848 & w1412);
assign w852 = (~w848 & w1413) | (~w848 & w1414) | (w1413 & w1414);
assign w853 = (~w120 & w1415) | (~w120 & w850) | (w1415 & w850);
assign w854 = ~w120 & ~w852;
assign w855 = w126 & ~w127;
assign w856 = ~w133 & w127;
assign w857 = ~w134 & ~w856;
assign w858 = (~w134 & w855) | (~w134 & w1127) | (w855 & w1127);
assign w859 = (~w140 & w856) | (~w140 & w1416) | (w856 & w1416);
assign w860 = ~w141 & ~w859;
assign w861 = (~w141 & w858) | (~w141 & w1417) | (w858 & w1417);
assign w862 = (~w858 & w1418) | (~w858 & w1419) | (w1418 & w1419);
assign w863 = (~w147 & w1420) | (~w147 & w860) | (w1420 & w860);
assign w864 = ~w147 & ~w862;
assign w865 = (~w860 & w1421) | (~w860 & w1422) | (w1421 & w1422);
assign w866 = (~w152 & w862) | (~w152 & w1421) | (w862 & w1421);
assign w867 = w153 & ~w158;
assign w868 = ~w159 & w158;
assign w869 = (~w164 & w867) | (~w164 & w1128) | (w867 & w1128);
assign w870 = (~w165 & w868) | (~w165 & w1423) | (w868 & w1423);
assign w871 = (~w170 & w869) | (~w170 & w1424) | (w869 & w1424);
assign w872 = ~w171 & ~w871;
assign w873 = (~w870 & w1426) | (~w870 & w1427) | (w1426 & w1427);
assign w874 = ~w177 & ~w873;
assign w875 = (~w182 & w873) | (~w182 & w1837) | (w873 & w1837);
assign w876 = (w871 & w1429) | (w871 & w1430) | (w1429 & w1430);
assign w877 = w183 & ~w188;
assign w878 = ~w189 & w188;
assign w879 = (~w195 & w877) | (~w195 & w1129) | (w877 & w1129);
assign w880 = (~w196 & w878) | (~w196 & w1431) | (w878 & w1431);
assign w881 = ~w196 & ~w879;
assign w882 = (~w202 & w879) | (~w202 & w1432) | (w879 & w1432);
assign w883 = (~w203 & w880) | (~w203 & w1433) | (w880 & w1433);
assign w884 = ~w203 & ~w882;
assign w885 = (~w880 & w1434) | (~w880 & w1435) | (w1434 & w1435);
assign w886 = ~w210 & ~w885;
assign w887 = (w882 & w1437) | (w882 & w1438) | (w1437 & w1438);
assign w888 = (~w885 & w2225) | (~w885 & w2226) | (w2225 & w2226);
assign w889 = (~w882 & w2227) | (~w882 & w2228) | (w2227 & w2228);
assign w890 = w223 & ~w224;
assign w891 = ~w230 & w224;
assign w892 = ~w231 & ~w891;
assign w893 = (~w231 & w890) | (~w231 & w1130) | (w890 & w1130);
assign w894 = (~w237 & w891) | (~w237 & w1440) | (w891 & w1440);
assign w895 = ~w238 & ~w894;
assign w896 = (~w238 & w893) | (~w238 & w1441) | (w893 & w1441);
assign w897 = (~w893 & w1442) | (~w893 & w1443) | (w1442 & w1443);
assign w898 = (~w245 & w1444) | (~w245 & w895) | (w1444 & w895);
assign w899 = ~w245 & ~w897;
assign w900 = (w895 & w1446) | (w895 & w1447) | (w1446 & w1447);
assign w901 = ~w251 & w2815;
assign w902 = (w897 & w1909) | (w897 & w1910) | (w1909 & w1910);
assign w903 = (w895 & w2229) | (w895 & w2230) | (w2229 & w2230);
assign w904 = (~w897 & w2231) | (~w897 & w2232) | (w2231 & w2232);
assign w905 = w263 & ~w264;
assign w906 = ~w269 & w264;
assign w907 = ~w270 & ~w906;
assign w908 = (~w270 & w905) | (~w270 & w1131) | (w905 & w1131);
assign w909 = (~w275 & w906) | (~w275 & w1450) | (w906 & w1450);
assign w910 = ~w276 & ~w909;
assign w911 = (~w276 & w908) | (~w276 & w1451) | (w908 & w1451);
assign w912 = ~w281 & ~w911;
assign w913 = (~w282 & w1452) | (~w282 & w910) | (w1452 & w910);
assign w914 = ~w282 & ~w912;
assign w915 = (w910 & w1454) | (w910 & w1455) | (w1454 & w1455);
assign w916 = ~w288 & w2816;
assign w917 = (w912 & w1911) | (w912 & w1912) | (w1911 & w1912);
assign w918 = (w910 & w2233) | (w910 & w2234) | (w2233 & w2234);
assign w919 = ~w294 & ~w917;
assign w920 = (w1458 & w1459) | (w1458 & ~w915) | (w1459 & ~w915);
assign w921 = (w912 & w2235) | (w912 & w2236) | (w2235 & w2236);
assign w922 = w300 & ~w306;
assign w923 = ~w307 & w306;
assign w924 = ~w307 & ~w922;
assign w925 = (~w312 & w922) | (~w312 & w1132) | (w922 & w1132);
assign w926 = (~w313 & w923) | (~w313 & w1460) | (w923 & w1460);
assign w927 = ~w313 & ~w925;
assign w928 = (~w318 & w925) | (~w318 & w1461) | (w925 & w1461);
assign w929 = (~w319 & w926) | (~w319 & w1462) | (w926 & w1462);
assign w930 = ~w319 & ~w928;
assign w931 = (~w926 & w1463) | (~w926 & w1464) | (w1463 & w1464);
assign w932 = ~w325 & ~w931;
assign w933 = ~w325 & w2817;
assign w934 = (~w332 & w1468) | (~w332 & w932) | (w1468 & w932);
assign w935 = (~w928 & w2237) | (~w928 & w2238) | (w2237 & w2238);
assign w936 = (w928 & w1913) | (w928 & w1914) | (w1913 & w1914);
assign w937 = (w1471 & w1470) | (w1471 & w932) | (w1470 & w932);
assign w938 = ~w338 & ~w936;
assign w939 = (~w932 & w1472) | (~w932 & w1473) | (w1472 & w1473);
assign w940 = (~w344 & w936) | (~w344 & w1474) | (w936 & w1474);
assign w941 = w345 & ~w351;
assign w942 = ~w352 & w351;
assign w943 = ~w352 & ~w941;
assign w944 = (~w357 & w941) | (~w357 & w1133) | (w941 & w1133);
assign w945 = (~w358 & w942) | (~w358 & w1475) | (w942 & w1475);
assign w946 = ~w358 & ~w944;
assign w947 = (~w363 & w944) | (~w363 & w1476) | (w944 & w1476);
assign w948 = (~w364 & w945) | (~w364 & w1477) | (w945 & w1477);
assign w949 = ~w364 & ~w947;
assign w950 = (~w945 & w1478) | (~w945 & w1479) | (w1478 & w1479);
assign w951 = ~w370 & ~w950;
assign w952 = (~w947 & w2241) | (~w947 & w2242) | (w2241 & w2242);
assign w953 = (w947 & w2243) | (w947 & w2244) | (w2243 & w2244);
assign w954 = (w1487 & w1486) | (w1487 & w951) | (w1486 & w951);
assign w955 = ~w382 & ~w953;
assign w956 = (~w951 & w1488) | (~w951 & w1489) | (w1488 & w1489);
assign w957 = (w951 & w2245) | (w951 & w2246) | (w2245 & w2246);
assign w958 = (~w953 & w1491) | (~w953 & w1492) | (w1491 & w1492);
assign w959 = w394 & ~w395;
assign w960 = ~w400 & w395;
assign w961 = ~w401 & ~w960;
assign w962 = (~w401 & w959) | (~w401 & w1134) | (w959 & w1134);
assign w963 = (~w406 & w960) | (~w406 & w1493) | (w960 & w1493);
assign w964 = ~w407 & ~w963;
assign w965 = (~w407 & w962) | (~w407 & w1494) | (w962 & w1494);
assign w966 = (~w962 & w1495) | (~w962 & w1496) | (w1495 & w1496);
assign w967 = (~w413 & w1497) | (~w413 & w964) | (w1497 & w964);
assign w968 = ~w413 & ~w966;
assign w969 = (w964 & w1499) | (w964 & w1500) | (w1499 & w1500);
assign w970 = (w964 & w2247) | (w964 & w2248) | (w2247 & w2248);
assign w971 = ~w425 & w2941;
assign w972 = (w966 & w2249) | (w966 & w2250) | (w2249 & w2250);
assign w973 = (w964 & w2652) | (w964 & w2653) | (w2652 & w2653);
assign w974 = ~w431 & ~w972;
assign w975 = (~w969 & w1506) | (~w969 & w1507) | (w1506 & w1507);
assign w976 = (w969 & w2251) | (w969 & w2252) | (w2251 & w2252);
assign w977 = (~w972 & w1509) | (~w972 & w1510) | (w1509 & w1510);
assign w978 = w443 & ~w444;
assign w979 = ~w450 & w444;
assign w980 = ~w451 & ~w979;
assign w981 = (~w451 & w978) | (~w451 & w1135) | (w978 & w1135);
assign w982 = (~w457 & w979) | (~w457 & w1511) | (w979 & w1511);
assign w983 = ~w458 & ~w982;
assign w984 = (~w458 & w981) | (~w458 & w1512) | (w981 & w1512);
assign w985 = (~w981 & w1513) | (~w981 & w1514) | (w1513 & w1514);
assign w986 = (~w465 & w1515) | (~w465 & w983) | (w1515 & w983);
assign w987 = ~w465 & ~w985;
assign w988 = (w983 & w1517) | (w983 & w1518) | (w1517 & w1518);
assign w989 = ~w472 & w2819;
assign w990 = (w983 & w2253) | (w983 & w2254) | (w2253 & w2254);
assign w991 = ~w479 & w2942;
assign w992 = (w985 & w2255) | (w985 & w2256) | (w2255 & w2256);
assign w993 = (w983 & w2654) | (w983 & w2655) | (w2654 & w2655);
assign w994 = ~w486 & ~w992;
assign w995 = (w988 & w1919) | (w988 & w1920) | (w1919 & w1920);
assign w996 = ~w493 & w2820;
assign w997 = (~w988 & w2626) | (~w988 & w2627) | (w2626 & w2627);
assign w998 = (w992 & w1527) | (w992 & w1528) | (w1527 & w1528);
assign w999 = w500 & ~w506;
assign w1000 = ~w507 & w506;
assign w1001 = ~w507 & ~w999;
assign w1002 = (~w512 & w999) | (~w512 & w1136) | (w999 & w1136);
assign w1003 = (~w513 & w1000) | (~w513 & w1529) | (w1000 & w1529);
assign w1004 = ~w513 & ~w1002;
assign w1005 = (~w518 & w1002) | (~w518 & w1530) | (w1002 & w1530);
assign w1006 = (~w519 & w1003) | (~w519 & w1531) | (w1003 & w1531);
assign w1007 = ~w519 & ~w1005;
assign w1008 = ~w524 & ~w1006;
assign w1009 = ~w525 & ~w1008;
assign w1010 = (~w531 & w1536) | (~w531 & w1009) | (w1536 & w1009);
assign w1011 = (~w1005 & w2257) | (~w1005 & w2258) | (w2257 & w2258);
assign w1012 = (w1005 & w2259) | (w1005 & w2260) | (w2259 & w2260);
assign w1013 = (w1539 & w1538) | (w1539 & w1009) | (w1538 & w1009);
assign w1014 = ~w537 & ~w1012;
assign w1015 = (w1009 & w2261) | (w1009 & w2262) | (w2261 & w2262);
assign w1016 = (w1012 & w1544) | (w1012 & w1545) | (w1544 & w1545);
assign w1017 = (w1009 & w2656) | (w1009 & w2657) | (w2656 & w2657);
assign w1018 = (~w1012 & w2263) | (~w1012 & w2264) | (w2263 & w2264);
assign w1019 = (~w1009 & w2658) | (~w1009 & w2659) | (w2658 & w2659);
assign w1020 = (w1012 & w2265) | (w1012 & w2266) | (w2265 & w2266);
assign w1021 = w555 & ~w561;
assign w1022 = ~w562 & w561;
assign w1023 = ~w562 & ~w1021;
assign w1024 = (~w567 & w1021) | (~w567 & w1137) | (w1021 & w1137);
assign w1025 = (~w568 & w1022) | (~w568 & w1549) | (w1022 & w1549);
assign w1026 = ~w568 & ~w1024;
assign w1027 = (~w573 & w1024) | (~w573 & w1550) | (w1024 & w1550);
assign w1028 = (~w574 & w1025) | (~w574 & w1551) | (w1025 & w1551);
assign w1029 = ~w574 & ~w1027;
assign w1030 = (~w1025 & w1552) | (~w1025 & w1553) | (w1552 & w1553);
assign w1031 = ~w580 & ~w1030;
assign w1032 = (~w586 & w1557) | (~w586 & w1031) | (w1557 & w1031);
assign w1033 = (~w1027 & w2267) | (~w1027 & w2268) | (w2267 & w2268);
assign w1034 = (w1027 & w2269) | (w1027 & w2270) | (w2269 & w2270);
assign w1035 = (w1560 & w1559) | (w1560 & w1031) | (w1559 & w1031);
assign w1036 = ~w592 & ~w1034;
assign w1037 = (w1031 & w2271) | (w1031 & w2272) | (w2271 & w2272);
assign w1038 = (w1031 & w2660) | (w1031 & w2661) | (w2660 & w2661);
assign w1039 = (~w1034 & w2273) | (~w1034 & w2274) | (w2273 & w2274);
assign w1040 = (w1034 & w2275) | (w1034 & w2276) | (w2275 & w2276);
assign w1041 = (w1031 & w2662) | (w1031 & w2663) | (w2662 & w2663);
assign w1042 = (w1856 & w1569) | (w1856 & w2825) | (w1569 & w2825);
assign w1043 = w616 & ~w617;
assign w1044 = ~w622 & w617;
assign w1045 = ~w623 & ~w1044;
assign w1046 = (~w623 & w1043) | (~w623 & w1138) | (w1043 & w1138);
assign w1047 = (~w628 & w1044) | (~w628 & w1199) | (w1044 & w1199);
assign w1048 = ~w629 & ~w1047;
assign w1049 = (~w629 & w1046) | (~w629 & w1200) | (w1046 & w1200);
assign w1050 = (~w1046 & w1571) | (~w1046 & w1572) | (w1571 & w1572);
assign w1051 = (~w1047 & w1573) | (~w1047 & w1574) | (w1573 & w1574);
assign w1052 = ~w636 & ~w1050;
assign w1053 = (~w643 & w1051) | (~w643 & w1576) | (w1051 & w1576);
assign w1054 = (~w1050 & w1576) | (~w1050 & w2279) | (w1576 & w2279);
assign w1055 = (w1051 & w1578) | (w1051 & w1579) | (w1578 & w1579);
assign w1056 = (~w1050 & w2280) | (~w1050 & w2281) | (w2280 & w2281);
assign w1057 = (w1050 & w2282) | (w1050 & w2283) | (w2282 & w2283);
assign w1058 = (w1051 & w2664) | (w1051 & w2665) | (w2664 & w2665);
assign w1059 = ~w657 & ~w1057;
assign w1060 = (w1051 & w2284) | (w1051 & w2285) | (w2284 & w2285);
assign w1061 = ~w663 & w2826;
assign w1062 = (w1055 & w2286) | (w1055 & w2287) | (w2286 & w2287);
assign w1063 = (w1587 & w1588) | (w1587 & w2826) | (w1588 & w2826);
assign w1064 = (w1057 & w2288) | (w1057 & w2289) | (w2288 & w2289);
assign w1065 = (w1055 & w2666) | (w1055 & w2667) | (w2666 & w2667);
assign w1066 = ~w675 & ~w1064;
assign w1067 = w681 & ~w682;
assign w1068 = ~w687 & w682;
assign w1069 = ~w688 & ~w1068;
assign w1070 = (~w688 & w1067) | (~w688 & w1139) | (w1067 & w1139);
assign w1071 = (~w693 & w1068) | (~w693 & w1146) | (w1068 & w1146);
assign w1072 = ~w694 & ~w1071;
assign w1073 = (~w694 & w1070) | (~w694 & w1147) | (w1070 & w1147);
assign w1074 = ~w699 & ~w1073;
assign w1075 = ~w700 & w2827;
assign w1076 = ~w700 & ~w1074;
assign w1077 = (~w706 & w1075) | (~w706 & w1593) | (w1075 & w1593);
assign w1078 = (~w1074 & w1593) | (~w1074 & w2290) | (w1593 & w2290);
assign w1079 = (w1074 & w1923) | (w1074 & w1924) | (w1923 & w1924);
assign w1080 = (w1075 & w2390) | (w1075 & w1595) | (w2390 & w1595);
assign w1081 = (~w1074 & w2291) | (~w1074 & w2292) | (w2291 & w2292);
assign w1082 = (w1074 & w2293) | (w1074 & w2294) | (w2293 & w2294);
assign w1083 = (w1075 & w2295) | (w1075 & w2296) | (w2295 & w2296);
assign w1084 = (w1075 & w2297) | (w1075 & w2298) | (w2297 & w2298);
assign w1085 = (~w1082 & w1861) | (~w1082 & w1599) | (w1861 & w1599);
assign w1086 = (w1080 & w2299) | (w1080 & w2300) | (w2299 & w2300);
assign w1087 = (w1603 & w1604) | (w1603 & w2828) | (w1604 & w2828);
assign w1088 = (w1082 & w2301) | (w1082 & w2302) | (w2301 & w2302);
assign w1089 = (w1080 & w2668) | (w1080 & w2669) | (w2668 & w2669);
assign w1090 = ~w736 & ~w1088;
assign w1091 = (~w1080 & w2670) | (~w1080 & w2671) | (w2670 & w2671);
assign w1092 = (w1082 & w2303) | (w1082 & w2304) | (w2303 & w2304);
assign w1093 = w742 & ~w747;
assign w1094 = ~w748 & w747;
assign w1095 = ~w748 & ~w1093;
assign w1096 = (~w753 & w1093) | (~w753 & w1148) | (w1093 & w1148);
assign w1097 = (~w754 & w1094) | (~w754 & w1202) | (w1094 & w1202);
assign w1098 = ~w754 & ~w1096;
assign w1099 = (~w759 & w1096) | (~w759 & w1203) | (w1096 & w1203);
assign w1100 = (~w760 & w1097) | (~w760 & w1610) | (w1097 & w1610);
assign w1101 = ~w760 & ~w1099;
assign w1102 = (~w1097 & w1611) | (~w1097 & w1612) | (w1611 & w1612);
assign w1103 = ~w766 & ~w1102;
assign w1104 = ~w766 & w2829;
assign w1105 = (~w772 & w1616) | (~w772 & w1103) | (w1616 & w1103);
assign w1106 = (~w1099 & w2305) | (~w1099 & w2306) | (w2305 & w2306);
assign w1107 = (w1099 & w1925) | (w1099 & w1926) | (w1925 & w1926);
assign w1108 = (w1619 & w1618) | (w1619 & w1103) | (w1618 & w1103);
assign w1109 = ~w778 & ~w1107;
assign w1110 = (w1103 & w2307) | (w1103 & w2308) | (w2307 & w2308);
assign w1111 = (~w1107 & w1622) | (~w1107 & w1623) | (w1622 & w1623);
assign w1112 = (w1103 & w2672) | (w1103 & w2673) | (w2672 & w2673);
assign w1113 = (~w1107 & w2309) | (~w1107 & w2310) | (w2309 & w2310);
assign w1114 = (w1103 & w2674) | (w1103 & w2675) | (w2674 & w2675);
assign w1115 = ~w796 & w2943;
assign w1116 = (w1110 & w1632) | (w1110 & w1633) | (w1632 & w1633);
assign w1117 = w1634 & w2831;
assign w1118 = (~w1110 & w1635) | (~w1110 & w1636) | (w1635 & w1636);
assign w1119 = (w1107 & w2777) | (w1107 & w2778) | (w2777 & w2778);
assign w1120 = ~w807 & w2944;
assign w1121 = (w1107 & w2779) | (w1107 & w2780) | (w2779 & w2780);
assign w1122 = w32 & ~w33;
assign w1123 = w46 & ~w47;
assign w1124 = w61 & ~w67;
assign w1125 = w83 & ~w88;
assign w1126 = w107 & ~w108;
assign w1127 = w133 & ~w134;
assign w1128 = w159 & ~w164;
assign w1129 = w189 & ~w195;
assign w1130 = w230 & ~w231;
assign w1131 = w269 & ~w270;
assign w1132 = w307 & ~w312;
assign w1133 = w352 & ~w357;
assign w1134 = w400 & ~w401;
assign w1135 = w450 & ~w451;
assign w1136 = w507 & ~w512;
assign w1137 = w562 & ~w567;
assign w1138 = w622 & ~w623;
assign w1139 = w687 & ~w688;
assign w1140 = (w1638 & w1639) | (w1638 & ~w1088) | (w1639 & ~w1088);
assign w1141 = (w1642 & w1641) | (w1642 & ~w1088) | (w1641 & ~w1088);
assign w1142 = (~w1088 & w1647) | (~w1088 & w1648) | (w1647 & w1648);
assign w1143 = (w1086 & w1651) | (w1086 & w1652) | (w1651 & w1652);
assign w1144 = (w1112 & w1113) | (w1112 & w2832) | (w1113 & w2832);
assign w1145 = (w1112 & w1113) | (w1112 & ~w1091) | (w1113 & ~w1091);
assign w1146 = w688 & ~w693;
assign w1147 = w693 & ~w694;
assign w1148 = w748 & ~w753;
assign w1149 = (~w682 & w1067) | (~w682 & w1066) | (w1067 & w1066);
assign w1150 = (w1070 & w1069) | (w1070 & w1066) | (w1069 & w1066);
assign w1151 = ~w700 & w2945;
assign w1152 = (w1062 & w1663) | (w1062 & w1664) | (w1663 & w1664);
assign w1153 = (w1062 & w2315) | (w1062 & w2316) | (w2315 & w2316);
assign w1154 = (~w1064 & w1666) | (~w1064 & w1667) | (w1666 & w1667);
assign w1155 = (w1085 & w1084) | (w1085 & w1066) | (w1084 & w1066);
assign w1156 = (~w1088 & w1668) | (~w1088 & w1669) | (w1668 & w1669);
assign w1157 = (w1092 & w1091) | (w1092 & ~w1066) | (w1091 & ~w1066);
assign w1158 = (w1088 & w1670) | (w1088 & w1671) | (w1670 & w1671);
assign w1159 = (w1080 & w2676) | (w1080 & w2677) | (w2676 & w2677);
assign w1160 = ~w749 & w1140;
assign w1161 = w749 & w2946;
assign w1162 = w749 & ~w1140;
assign w1163 = (w1086 & w1672) | (w1086 & w1673) | (w1672 & w1673);
assign w1164 = (w1095 & w1877) | (w1095 & w2947) | (w1877 & w2947);
assign w1165 = w755 & w2948;
assign w1166 = w755 & ~w1141;
assign w1167 = (w1086 & w1674) | (w1086 & w1675) | (w1674 & w1675);
assign w1168 = (w1098 & w1880) | (w1098 & w2833) | (w1880 & w2833);
assign w1169 = (~w1098 & w1884) | (~w1098 & w2834) | (w1884 & w2834);
assign w1170 = (w1088 & w1676) | (w1088 & w2317) | (w1676 & w2317);
assign w1171 = (w1086 & w1677) | (w1086 & w1678) | (w1677 & w1678);
assign w1172 = ~w767 & w2835;
assign w1173 = w767 & w2836;
assign w1174 = (w1088 & w1679) | (w1088 & w2318) | (w1679 & w2318);
assign w1175 = (w1086 & w1680) | (w1086 & w1681) | (w1680 & w1681);
assign w1176 = (~w1088 & w1681) | (~w1088 & w1682) | (w1681 & w1682);
assign w1177 = (~w1086 & w1683) | (~w1086 & w1684) | (w1683 & w1684);
assign w1178 = w773 & ~w1142;
assign w1179 = ~w779 & w1143;
assign w1180 = (~w1088 & w1685) | (~w1088 & w1686) | (w1685 & w1686);
assign w1181 = w779 & ~w1143;
assign w1182 = (w1088 & w1687) | (w1088 & w1688) | (w1687 & w1688);
assign w1183 = (~w1091 & w2319) | (~w1091 & w2320) | (w2319 & w2320);
assign w1184 = (~w1088 & w1689) | (~w1088 & w1690) | (w1689 & w1690);
assign w1185 = (w1091 & w1691) | (w1091 & w1692) | (w1691 & w1692);
assign w1186 = (w1088 & w1693) | (w1088 & w1694) | (w1693 & w1694);
assign w1187 = (~w1091 & w2321) | (~w1091 & w2322) | (w2321 & w2322);
assign w1188 = (~w1088 & w1695) | (~w1088 & w1696) | (w1695 & w1696);
assign w1189 = (w1091 & w1697) | (w1091 & w1698) | (w1697 & w1698);
assign w1190 = (w1088 & w1699) | (w1088 & w1700) | (w1699 & w1700);
assign w1191 = ~w797 & w1145;
assign w1192 = ~w797 & w1144;
assign w1193 = w797 & ~w1145;
assign w1194 = w797 & ~w1144;
assign w1195 = (w1115 & w1701) | (w1115 & w1702) | (w1701 & w1702);
assign w1196 = (~w1092 & w1702) | (~w1092 & w1703) | (w1702 & w1703);
assign w1197 = (~w1115 & w1704) | (~w1115 & w1705) | (w1704 & w1705);
assign w1198 = (~w1114 & w2323) | (~w1114 & w2324) | (w2323 & w2324);
assign w1199 = w623 & ~w628;
assign w1200 = w628 & ~w629;
assign w1201 = w694 & ~w699;
assign w1202 = w753 & ~w754;
assign w1203 = w754 & ~w759;
assign w1204 = (w1707 & w1706) | (w1707 & ~w1040) | (w1706 & ~w1040);
assign w1205 = (w1031 & w2678) | (w1031 & w2679) | (w2678 & w2679);
assign w1206 = (w1709 & w1708) | (w1709 & ~w1040) | (w1708 & ~w1040);
assign w1207 = (w1031 & w2680) | (w1031 & w2681) | (w2680 & w2681);
assign w1208 = (~w1040 & w1710) | (~w1040 & w1711) | (w1710 & w1711);
assign w1209 = (w1037 & w1712) | (w1037 & w1713) | (w1712 & w1713);
assign w1210 = (~w1040 & w1714) | (~w1040 & w1715) | (w1714 & w1715);
assign w1211 = (w1037 & w1716) | (w1037 & w1717) | (w1716 & w1717);
assign w1212 = (~w1040 & w1718) | (~w1040 & w1719) | (w1718 & w1719);
assign w1213 = (w1037 & w1720) | (w1037 & w1721) | (w1720 & w1721);
assign w1214 = (~w1040 & w1722) | (~w1040 & w1723) | (w1722 & w1723);
assign w1215 = (w1037 & w2325) | (w1037 & w2326) | (w2325 & w2326);
assign w1216 = (w1059 & w1058) | (w1059 & w1042) | (w1058 & w1042);
assign w1217 = (w1061 & w1060) | (w1061 & w1042) | (w1060 & w1042);
assign w1218 = (w1063 & w1062) | (w1063 & w1041) | (w1062 & w1041);
assign w1219 = (w1066 & w1065) | (w1066 & w1042) | (w1065 & w1042);
assign w1220 = (~w1064 & w1724) | (~w1064 & w1725) | (w1724 & w1725);
assign w1221 = (w1055 & w2682) | (w1055 & w2683) | (w2682 & w2683);
assign w1222 = ~w689 & w2949;
assign w1223 = w689 & w2950;
assign w1224 = w689 & ~w1149;
assign w1225 = (w1062 & w1726) | (w1062 & w1727) | (w1726 & w1727);
assign w1226 = ~w695 & w1150;
assign w1227 = w695 & w2837;
assign w1228 = w695 & ~w1150;
assign w1229 = (w1062 & w1728) | (w1062 & w1729) | (w1728 & w1729);
assign w1230 = ~w701 & w2838;
assign w1231 = w701 & w2839;
assign w1232 = (w1064 & w1730) | (w1064 & w2327) | (w1730 & w2327);
assign w1233 = (w1062 & w1731) | (w1062 & w1732) | (w1731 & w1732);
assign w1234 = (w2383 & w1076) | (w2383 & w2840) | (w1076 & w2840);
assign w1235 = w707 & w2951;
assign w1236 = w707 & ~w1151;
assign w1237 = ~w713 & w1152;
assign w1238 = (~w1064 & w1733) | (~w1064 & w1734) | (w1733 & w1734);
assign w1239 = w713 & ~w1152;
assign w1240 = (w1064 & w1735) | (w1064 & w1736) | (w1735 & w1736);
assign w1241 = ~w719 & w1153;
assign w1242 = (~w1064 & w1737) | (~w1064 & w1738) | (w1737 & w1738);
assign w1243 = w719 & w2952;
assign w1244 = (w1064 & w1739) | (w1064 & w1740) | (w1739 & w1740);
assign w1245 = (w1065 & w2328) | (w1065 & w2329) | (w2328 & w2329);
assign w1246 = ~w725 & w1154;
assign w1247 = (~w1065 & w2330) | (~w1065 & w2331) | (w2330 & w2331);
assign w1248 = w725 & ~w1154;
assign w1249 = (w1065 & w2332) | (w1065 & w2333) | (w2332 & w2333);
assign w1250 = (w1066 & w1741) | (w1066 & w1742) | (w1741 & w1742);
assign w1251 = w731 & w2953;
assign w1252 = w731 & ~w1155;
assign w1253 = (w1087 & w1743) | (w1087 & w1744) | (w1743 & w1744);
assign w1254 = (w1066 & w1743) | (w1066 & w1745) | (w1743 & w1745);
assign w1255 = (~w1087 & w1746) | (~w1087 & w1747) | (w1746 & w1747);
assign w1256 = (~w1087 & w2334) | (~w1087 & w1746) | (w2334 & w1746);
assign w1257 = ~w743 & w1156;
assign w1258 = (w1089 & w2335) | (w1089 & w2336) | (w2335 & w2336);
assign w1259 = w743 & ~w1156;
assign w1260 = (~w1089 & w2337) | (~w1089 & w2338) | (w2337 & w2338);
assign w1261 = ~w13 & ~w21;
assign w1262 = w13 & w21;
assign w1263 = ~w34 & ~w27;
assign w1264 = ~w34 & w819;
assign w1265 = ~w41 & w822;
assign w1266 = ~w41 & w821;
assign w1267 = (~w40 & w823) | (~w40 & w822) | (w823 & w822);
assign w1268 = (~w40 & w823) | (~w40 & w821) | (w823 & w821);
assign w1269 = (w826 & w825) | (w826 & w822) | (w825 & w822);
assign w1270 = (w826 & w825) | (w826 & w821) | (w825 & w821);
assign w1271 = ~w61 & w2841;
assign w1272 = ~w61 & w2842;
assign w1273 = (w833 & w832) | (w833 & ~w828) | (w832 & ~w828);
assign w1274 = (w833 & w832) | (w833 & ~w827) | (w832 & ~w827);
assign w1275 = ~w75 & ~w835;
assign w1276 = (~w75 & w832) | (~w75 & w1749) | (w832 & w1749);
assign w1277 = (w841 & w840) | (w841 & ~w835) | (w840 & ~w835);
assign w1278 = (w841 & w840) | (w841 & ~w834) | (w840 & ~w834);
assign w1279 = ~w842 & w1750;
assign w1280 = (w840 & w1750) | (w840 & w1751) | (w1750 & w1751);
assign w1281 = (w103 & w842) | (w103 & w1752) | (w842 & w1752);
assign w1282 = w103 & ~w843;
assign w1283 = (w840 & w1754) | (w840 & w1755) | (w1754 & w1755);
assign w1284 = (w848 & w847) | (w848 & w844) | (w847 & w844);
assign w1285 = (w851 & w850) | (w851 & w844) | (w850 & w844);
assign w1286 = (w851 & w850) | (w851 & w843) | (w850 & w843);
assign w1287 = ~w852 & w1756;
assign w1288 = (w850 & w1756) | (w850 & w1757) | (w1756 & w1757);
assign w1289 = (w128 & w852) | (w128 & w1758) | (w852 & w1758);
assign w1290 = w128 & ~w853;
assign w1291 = (~w127 & w855) | (~w127 & w854) | (w855 & w854);
assign w1292 = (w850 & w1759) | (w850 & w1760) | (w1759 & w1760);
assign w1293 = (w858 & w857) | (w858 & w854) | (w857 & w854);
assign w1294 = (w850 & w1761) | (w850 & w1762) | (w1761 & w1762);
assign w1295 = (w861 & w860) | (w861 & w853) | (w860 & w853);
assign w1296 = (w864 & w863) | (w864 & w854) | (w863 & w854);
assign w1297 = ~w159 & w2954;
assign w1298 = (w860 & w1766) | (w860 & w1767) | (w1766 & w1767);
assign w1299 = ~w177 & w2843;
assign w1300 = ~w177 & w2844;
assign w1301 = (~w871 & w2339) | (~w871 & w2340) | (w2339 & w2340);
assign w1302 = (~w183 & w1768) | (~w183 & w874) | (w1768 & w874);
assign w1303 = ~w189 & w2955;
assign w1304 = (w874 & w1769) | (w874 & w1770) | (w1769 & w1770);
assign w1305 = (w881 & w880) | (w881 & ~w876) | (w880 & ~w876);
assign w1306 = (w874 & w1771) | (w874 & w1772) | (w1771 & w1772);
assign w1307 = w1773 & ~w887;
assign w1308 = ~w225 & w2956;
assign w1309 = (w882 & w2341) | (w882 & w2342) | (w2341 & w2342);
assign w1310 = (w885 & w2343) | (w885 & w2344) | (w2343 & w2344);
assign w1311 = (w893 & w892) | (w893 & w2845) | (w892 & w2845);
assign w1312 = (w886 & w1775) | (w886 & w1776) | (w1775 & w1776);
assign w1313 = (w896 & w895) | (w896 & w2845) | (w895 & w2845);
assign w1314 = (w886 & w1777) | (w886 & w1778) | (w1777 & w1778);
assign w1315 = (w899 & w898) | (w899 & w889) | (w898 & w889);
assign w1316 = (w899 & w898) | (w899 & w888) | (w898 & w888);
assign w1317 = (w901 & w900) | (w901 & w889) | (w900 & w889);
assign w1318 = (w901 & w900) | (w901 & w888) | (w900 & w888);
assign w1319 = w1779 & ~w902;
assign w1320 = (w895 & w2345) | (w895 & w2346) | (w2345 & w2346);
assign w1321 = (w897 & w2347) | (w897 & w2348) | (w2347 & w2348);
assign w1322 = w265 & w2957;
assign w1323 = (~w264 & w905) | (~w264 & w2846) | (w905 & w2846);
assign w1324 = (w895 & w2349) | (w895 & w2350) | (w2349 & w2350);
assign w1325 = (w911 & w910) | (w911 & w2846) | (w910 & w2846);
assign w1326 = (w900 & w1784) | (w900 & w1785) | (w1784 & w1785);
assign w1327 = (w914 & w913) | (w914 & w2846) | (w913 & w2846);
assign w1328 = (w914 & w913) | (w914 & w903) | (w913 & w903);
assign w1329 = (w916 & w915) | (w916 & w904) | (w915 & w904);
assign w1330 = (w916 & w915) | (w916 & w903) | (w915 & w903);
assign w1331 = (w919 & w918) | (w919 & w904) | (w918 & w904);
assign w1332 = (w919 & w918) | (w919 & w903) | (w918 & w903);
assign w1333 = ~w300 & w2847;
assign w1334 = (w910 & w2684) | (w910 & w2685) | (w2684 & w2685);
assign w1335 = (w923 & w924) | (w923 & w2847) | (w924 & w2847);
assign w1336 = (w915 & w1789) | (w915 & w1790) | (w1789 & w1790);
assign w1337 = (w926 & w927) | (w926 & w2847) | (w927 & w2847);
assign w1338 = (w915 & w1791) | (w915 & w1792) | (w1791 & w1792);
assign w1339 = (w929 & w930) | (w929 & w2847) | (w930 & w2847);
assign w1340 = (w930 & w929) | (w930 & ~w920) | (w929 & ~w920);
assign w1341 = (~w917 & w1793) | (~w917 & w1794) | (w1793 & w1794);
assign w1342 = ~w325 & w2848;
assign w1343 = (w932 & w2351) | (w932 & w2352) | (w2351 & w2352);
assign w1344 = (w945 & w946) | (w945 & ~w940) | (w946 & ~w940);
assign w1345 = (w932 & w2353) | (w932 & w2354) | (w2353 & w2354);
assign w1346 = (w948 & w949) | (w948 & ~w940) | (w949 & ~w940);
assign w1347 = (w932 & w2355) | (w932 & w2356) | (w2355 & w2356);
assign w1348 = ~w370 & w2958;
assign w1349 = (w955 & w954) | (w955 & ~w940) | (w954 & ~w940);
assign w1350 = (w955 & w954) | (w955 & ~w939) | (w954 & ~w939);
assign w1351 = ~w396 & w958;
assign w1352 = (w951 & w2357) | (w951 & w2358) | (w2357 & w2358);
assign w1353 = (w953 & w1798) | (w953 & w1799) | (w1798 & w1799);
assign w1354 = (w396 & w1800) | (w396 & w956) | (w1800 & w956);
assign w1355 = (w951 & w2359) | (w951 & w2360) | (w2359 & w2360);
assign w1356 = (w951 & w2361) | (w951 & w2362) | (w2361 & w2362);
assign w1357 = (w965 & w964) | (w965 & w958) | (w964 & w958);
assign w1358 = (w968 & w967) | (w968 & w958) | (w967 & w958);
assign w1359 = (w968 & w967) | (w968 & w2849) | (w967 & w2849);
assign w1360 = (w974 & w973) | (w974 & w958) | (w973 & w958);
assign w1361 = (w974 & w973) | (w974 & w957) | (w973 & w957);
assign w1362 = ~w445 & w977;
assign w1363 = (w969 & w2363) | (w969 & w2364) | (w2363 & w2364);
assign w1364 = (w972 & w1807) | (w972 & w1808) | (w1807 & w1808);
assign w1365 = (w445 & w1809) | (w445 & w975) | (w1809 & w975);
assign w1366 = (~w444 & w978) | (~w444 & w977) | (w978 & w977);
assign w1367 = (w969 & w2365) | (w969 & w2366) | (w2365 & w2366);
assign w1368 = (w981 & w980) | (w981 & w977) | (w980 & w977);
assign w1369 = (w969 & w2367) | (w969 & w2368) | (w2367 & w2368);
assign w1370 = (w984 & w983) | (w984 & w977) | (w983 & w977);
assign w1371 = (w984 & w983) | (w984 & w2850) | (w983 & w2850);
assign w1372 = (w987 & w986) | (w987 & w977) | (w986 & w977);
assign w1373 = (w987 & w986) | (w987 & w2850) | (w986 & w2850);
assign w1374 = (~w972 & w1810) | (~w972 & w1811) | (w1810 & w1811);
assign w1375 = (w989 & w988) | (w989 & w976) | (w988 & w976);
assign w1376 = (w991 & w990) | (w991 & w977) | (w990 & w977);
assign w1377 = (w991 & w990) | (w991 & w976) | (w990 & w976);
assign w1378 = (w994 & w993) | (w994 & w977) | (w993 & w977);
assign w1379 = (w994 & w993) | (w994 & w976) | (w993 & w976);
assign w1380 = (w996 & w995) | (w996 & w977) | (w995 & w977);
assign w1381 = (w996 & w995) | (w996 & w976) | (w995 & w976);
assign w1382 = (w1003 & w1004) | (w1003 & ~w998) | (w1004 & ~w998);
assign w1383 = (w1006 & w1007) | (w1006 & ~w998) | (w1007 & ~w998);
assign w1384 = ~w525 & w2959;
assign w1385 = (w995 & w1818) | (w995 & w1819) | (w1818 & w1819);
assign w1386 = (~w992 & w1820) | (~w992 & w1821) | (w1820 & w1821);
assign w1387 = (w995 & w1822) | (w995 & w1823) | (w1822 & w1823);
assign w1388 = (w1014 & w1013) | (w1014 & ~w998) | (w1013 & ~w998);
assign w1389 = (w2910 & w1015) | (w2910 & ~w998) | (w1015 & ~w998);
assign w1390 = (w1018 & w1017) | (w1018 & ~w997) | (w1017 & ~w997);
assign w1391 = (w1009 & w2686) | (w1009 & w2687) | (w2686 & w2687);
assign w1392 = ~w562 & w2960;
assign w1393 = (w1009 & w2688) | (w1009 & w2689) | (w2688 & w2689);
assign w1394 = ~w580 & w2961;
assign w1395 = (w1015 & w1831) | (w1015 & w1832) | (w1831 & w1832);
assign w1396 = (w1033 & w1032) | (w1033 & w2851) | (w1032 & w2851);
assign w1397 = (w1015 & w1833) | (w1015 & w1834) | (w1833 & w1834);
assign w1398 = (w1036 & w1035) | (w1036 & ~w1020) | (w1035 & ~w1020);
assign w1399 = (w2913 & w1037) | (w2913 & ~w1020) | (w1037 & ~w1020);
assign w1400 = (w1039 & w1038) | (w1039 & ~w1019) | (w1038 & ~w1019);
assign w1401 = w1835 & ~w1040;
assign w1402 = (w1031 & w2690) | (w1031 & w2691) | (w2690 & w2691);
assign w1403 = (w1034 & w2371) | (w1034 & w2372) | (w2371 & w2372);
assign w1404 = w618 & w2962;
assign w1405 = w47 & ~w53;
assign w1406 = w67 & ~w68;
assign w1407 = w68 & ~w74;
assign w1408 = w88 & ~w89;
assign w1409 = w89 & ~w94;
assign w1410 = w94 & ~w95;
assign w1411 = w108 & ~w113;
assign w1412 = w113 & ~w114;
assign w1413 = ~w119 & w114;
assign w1414 = ~w119 & ~w1412;
assign w1415 = w119 & ~w120;
assign w1416 = w134 & ~w140;
assign w1417 = w140 & ~w141;
assign w1418 = ~w146 & w141;
assign w1419 = ~w146 & ~w1417;
assign w1420 = w146 & ~w147;
assign w1421 = ~w152 & w147;
assign w1422 = ~w152 & ~w1420;
assign w1423 = w164 & ~w165;
assign w1424 = w165 & ~w170;
assign w1425 = w170 & ~w171;
assign w1426 = ~w176 & w171;
assign w1427 = ~w176 & ~w1425;
assign w1428 = ~w177 & w176;
assign w1429 = ~w182 & ~w1428;
assign w1430 = (~w182 & w1426) | (~w182 & w1837) | (w1426 & w1837);
assign w1431 = w195 & ~w196;
assign w1432 = w196 & ~w202;
assign w1433 = w202 & ~w203;
assign w1434 = ~w209 & w203;
assign w1435 = ~w209 & ~w1433;
assign w1436 = ~w210 & w209;
assign w1437 = ~w216 & ~w1436;
assign w1438 = (~w216 & w1434) | (~w216 & w1838) | (w1434 & w1838);
assign w1439 = w216 & ~w217;
assign w1440 = w231 & ~w237;
assign w1441 = w237 & ~w238;
assign w1442 = ~w244 & w238;
assign w1443 = ~w244 & ~w1441;
assign w1444 = w244 & ~w245;
assign w1445 = ~w250 & w245;
assign w1446 = ~w251 & ~w1445;
assign w1447 = (~w251 & w1444) | (~w251 & w1839) | (w1444 & w1839);
assign w1448 = w251 & ~w256;
assign w1449 = w256 & ~w257;
assign w1450 = w270 & ~w275;
assign w1451 = w275 & ~w276;
assign w1452 = w281 & ~w282;
assign w1453 = ~w287 & w282;
assign w1454 = ~w288 & ~w1453;
assign w1455 = (~w288 & w1452) | (~w288 & w1840) | (w1452 & w1840);
assign w1456 = w288 & ~w293;
assign w1457 = w293 & ~w294;
assign w1458 = ~w299 & w294;
assign w1459 = ~w299 & ~w1457;
assign w1460 = w312 & ~w313;
assign w1461 = w313 & ~w318;
assign w1462 = w318 & ~w319;
assign w1463 = ~w324 & w319;
assign w1464 = ~w324 & ~w1462;
assign w1465 = ~w325 & w324;
assign w1466 = ~w331 & ~w1465;
assign w1467 = (~w331 & w1463) | (~w331 & w1841) | (w1463 & w1841);
assign w1468 = w331 & ~w332;
assign w1469 = ~w337 & w332;
assign w1470 = ~w338 & ~w1469;
assign w1471 = (~w338 & w1468) | (~w338 & w1842) | (w1468 & w1842);
assign w1472 = (~w344 & w1469) | (~w344 & w1474) | (w1469 & w1474);
assign w1473 = ~w344 & ~w1471;
assign w1474 = w338 & ~w344;
assign w1475 = w357 & ~w358;
assign w1476 = w358 & ~w363;
assign w1477 = w363 & ~w364;
assign w1478 = ~w369 & w364;
assign w1479 = ~w369 & ~w1477;
assign w1480 = ~w370 & w369;
assign w1481 = ~w370 & ~w1478;
assign w1482 = ~w375 & ~w1480;
assign w1483 = (~w375 & w1478) | (~w375 & w1843) | (w1478 & w1843);
assign w1484 = w375 & ~w376;
assign w1485 = ~w381 & w376;
assign w1486 = ~w382 & ~w1485;
assign w1487 = (~w382 & w1484) | (~w382 & w1844) | (w1484 & w1844);
assign w1488 = (~w387 & w1485) | (~w387 & w1490) | (w1485 & w1490);
assign w1489 = ~w387 & ~w1487;
assign w1490 = w382 & ~w387;
assign w1491 = ~w388 & w387;
assign w1492 = ~w388 & ~w1490;
assign w1493 = w401 & ~w406;
assign w1494 = w406 & ~w407;
assign w1495 = ~w412 & w407;
assign w1496 = ~w412 & ~w1494;
assign w1497 = w412 & ~w413;
assign w1498 = ~w418 & w413;
assign w1499 = ~w419 & ~w1498;
assign w1500 = (~w419 & w1497) | (~w419 & w1845) | (w1497 & w1845);
assign w1501 = w419 & ~w424;
assign w1502 = w424 & ~w425;
assign w1503 = ~w430 & w425;
assign w1504 = ~w431 & ~w1503;
assign w1505 = (~w431 & w1502) | (~w431 & w1846) | (w1502 & w1846);
assign w1506 = (~w436 & w1503) | (~w436 & w1508) | (w1503 & w1508);
assign w1507 = ~w436 & ~w1505;
assign w1508 = w431 & ~w436;
assign w1509 = ~w437 & w436;
assign w1510 = ~w437 & ~w1508;
assign w1511 = w451 & ~w457;
assign w1512 = w457 & ~w458;
assign w1513 = ~w464 & w458;
assign w1514 = ~w464 & ~w1512;
assign w1515 = w464 & ~w465;
assign w1516 = ~w471 & w465;
assign w1517 = ~w472 & ~w1516;
assign w1518 = (~w472 & w1515) | (~w472 & w1847) | (w1515 & w1847);
assign w1519 = w472 & ~w478;
assign w1520 = w478 & ~w479;
assign w1521 = ~w485 & w479;
assign w1522 = ~w486 & ~w1521;
assign w1523 = (~w486 & w1520) | (~w486 & w1848) | (w1520 & w1848);
assign w1524 = (~w492 & w1521) | (~w492 & w1525) | (w1521 & w1525);
assign w1525 = w486 & ~w492;
assign w1526 = ~w493 & w492;
assign w1527 = ~w499 & ~w1526;
assign w1528 = (~w499 & w1525) | (~w499 & w1849) | (w1525 & w1849);
assign w1529 = w512 & ~w513;
assign w1530 = w513 & ~w518;
assign w1531 = w518 & ~w519;
assign w1532 = ~w524 & w519;
assign w1533 = ~w525 & w524;
assign w1534 = ~w530 & ~w1533;
assign w1535 = (~w530 & w1532) | (~w530 & w1850) | (w1532 & w1850);
assign w1536 = w530 & ~w531;
assign w1537 = ~w536 & w531;
assign w1538 = ~w537 & ~w1537;
assign w1539 = (~w537 & w1536) | (~w537 & w1851) | (w1536 & w1851);
assign w1540 = (~w542 & w1537) | (~w542 & w1541) | (w1537 & w1541);
assign w1541 = w537 & ~w542;
assign w1542 = ~w543 & w542;
assign w1543 = ~w543 & ~w1541;
assign w1544 = ~w548 & ~w1542;
assign w1545 = (~w548 & w1541) | (~w548 & w1852) | (w1541 & w1852);
assign w1546 = w548 & ~w549;
assign w1547 = ~w554 & w549;
assign w1548 = ~w554 & ~w1546;
assign w1549 = w567 & ~w568;
assign w1550 = w568 & ~w573;
assign w1551 = w573 & ~w574;
assign w1552 = ~w579 & w574;
assign w1553 = ~w579 & ~w1551;
assign w1554 = ~w580 & w579;
assign w1555 = ~w585 & ~w1554;
assign w1556 = (~w585 & w1552) | (~w585 & w1853) | (w1552 & w1853);
assign w1557 = w585 & ~w586;
assign w1558 = ~w591 & w586;
assign w1559 = ~w592 & ~w1558;
assign w1560 = (~w592 & w1557) | (~w592 & w1854) | (w1557 & w1854);
assign w1561 = (~w597 & w1558) | (~w597 & w1562) | (w1558 & w1562);
assign w1562 = w592 & ~w597;
assign w1563 = ~w598 & w597;
assign w1564 = ~w598 & ~w1562;
assign w1565 = ~w603 & ~w1563;
assign w1566 = (~w603 & w1562) | (~w603 & w1855) | (w1562 & w1855);
assign w1567 = w603 & ~w604;
assign w1568 = ~w609 & w604;
assign w1569 = ~w610 & ~w1568;
assign w1570 = (~w610 & w1567) | (~w610 & w1856) | (w1567 & w1856);
assign w1571 = w629 & ~w635;
assign w1572 = ~w635 & ~w1200;
assign w1573 = ~w636 & w635;
assign w1574 = ~w636 & ~w1571;
assign w1575 = w636 & ~w642;
assign w1576 = w642 & ~w643;
assign w1577 = ~w649 & w643;
assign w1578 = ~w650 & ~w1577;
assign w1579 = (~w650 & w1576) | (~w650 & w1857) | (w1576 & w1857);
assign w1580 = w650 & ~w656;
assign w1581 = w656 & ~w657;
assign w1582 = ~w662 & w657;
assign w1583 = ~w663 & ~w1582;
assign w1584 = (~w663 & w1581) | (~w663 & w1858) | (w1581 & w1858);
assign w1585 = (~w668 & w1582) | (~w668 & w1586) | (w1582 & w1586);
assign w1586 = w663 & ~w668;
assign w1587 = ~w669 & w668;
assign w1588 = ~w669 & ~w1586;
assign w1589 = ~w674 & ~w1587;
assign w1590 = (~w674 & w1586) | (~w674 & w1859) | (w1586 & w1859);
assign w1591 = w674 & ~w675;
assign w1592 = w700 & ~w705;
assign w1593 = w705 & ~w706;
assign w1594 = ~w711 & w706;
assign w1595 = (~w712 & w1593) | (~w712 & w1860) | (w1593 & w1860);
assign w1596 = w712 & ~w717;
assign w1597 = w717 & ~w718;
assign w1598 = ~w723 & w718;
assign w1599 = ~w724 & ~w1598;
assign w1600 = (~w724 & w1597) | (~w724 & w1861) | (w1597 & w1861);
assign w1601 = (~w729 & w1598) | (~w729 & w1602) | (w1598 & w1602);
assign w1602 = w724 & ~w729;
assign w1603 = ~w730 & w729;
assign w1604 = ~w730 & ~w1602;
assign w1605 = ~w735 & ~w1603;
assign w1606 = (~w735 & w1602) | (~w735 & w1862) | (w1602 & w1862);
assign w1607 = w735 & ~w736;
assign w1608 = ~w741 & w736;
assign w1609 = ~w741 & ~w1607;
assign w1610 = w759 & ~w760;
assign w1611 = ~w765 & w760;
assign w1612 = ~w765 & ~w1610;
assign w1613 = ~w766 & w765;
assign w1614 = ~w771 & ~w1613;
assign w1615 = (~w771 & w1611) | (~w771 & w1863) | (w1611 & w1863);
assign w1616 = w771 & ~w772;
assign w1617 = ~w777 & w772;
assign w1618 = ~w778 & ~w1617;
assign w1619 = (~w778 & w1616) | (~w778 & w1864) | (w1616 & w1864);
assign w1620 = (~w783 & w1617) | (~w783 & w1621) | (w1617 & w1621);
assign w1621 = w778 & ~w783;
assign w1622 = ~w784 & w783;
assign w1623 = ~w784 & ~w1621;
assign w1624 = ~w789 & ~w1622;
assign w1625 = (~w789 & w1621) | (~w789 & w1865) | (w1621 & w1865);
assign w1626 = w789 & ~w790;
assign w1627 = ~w795 & w790;
assign w1628 = ~w796 & ~w1627;
assign w1629 = (~w796 & w1626) | (~w796 & w1866) | (w1626 & w1866);
assign w1630 = ~w801 & ~w1629;
assign w1631 = w796 & ~w801;
assign w1632 = (w1628 & w1634) | (w1628 & w1868) | (w1634 & w1868);
assign w1633 = ~w1630 & w1634;
assign w1634 = ~w802 & ~w809;
assign w1635 = w809 & w2852;
assign w1636 = (w809 & w1630) | (w809 & w1637) | (w1630 & w1637);
assign w1637 = w802 & w809;
assign w1638 = ~w742 & w741;
assign w1639 = ~w742 & ~w1608;
assign w1640 = (~w742 & w1607) | (~w742 & w1638) | (w1607 & w1638);
assign w1641 = ~w748 & w2853;
assign w1642 = ~w748 & w2854;
assign w1643 = ~w748 & w2855;
assign w1644 = (w1100 & w1101) | (w1100 & w741) | (w1101 & w741);
assign w1645 = (w1100 & w1101) | (w1100 & ~w1608) | (w1101 & ~w1608);
assign w1646 = (w1100 & w1101) | (w1100 & ~w1609) | (w1101 & ~w1609);
assign w1647 = (w1103 & w1104) | (w1103 & w741) | (w1104 & w741);
assign w1648 = (w1103 & w1104) | (w1103 & ~w1608) | (w1104 & ~w1608);
assign w1649 = (w1103 & w1104) | (w1103 & ~w1609) | (w1104 & ~w1609);
assign w1650 = (w1105 & w1106) | (w1105 & w741) | (w1106 & w741);
assign w1651 = (w1105 & w1106) | (w1105 & ~w1608) | (w1106 & ~w1608);
assign w1652 = (w1105 & w1106) | (w1105 & ~w1609) | (w1106 & ~w1609);
assign w1653 = (w1110 & w1111) | (w1110 & w741) | (w1111 & w741);
assign w1654 = (w1110 & w1111) | (w1110 & ~w1608) | (w1111 & ~w1608);
assign w1655 = (~w682 & w1067) | (~w682 & ~w675) | (w1067 & ~w675);
assign w1656 = (~w682 & w1067) | (~w682 & w1591) | (w1067 & w1591);
assign w1657 = (w1070 & w1069) | (w1070 & ~w675) | (w1069 & ~w675);
assign w1658 = (w1070 & w1069) | (w1070 & w1591) | (w1069 & w1591);
assign w1659 = w1072 & w1073;
assign w1660 = (w1073 & w1072) | (w1073 & ~w675) | (w1072 & ~w675);
assign w1661 = (w1073 & w1072) | (w1073 & w1591) | (w1072 & w1591);
assign w1662 = w1078 & w1077;
assign w1663 = (w1077 & w1078) | (w1077 & ~w675) | (w1078 & ~w675);
assign w1664 = (w1077 & w1078) | (w1077 & w1591) | (w1078 & w1591);
assign w1665 = (~w1079 & w1871) | (~w1079 & w1872) | (w1871 & w1872);
assign w1666 = ~w1082 & w1873;
assign w1667 = (~w1082 & w1874) | (~w1082 & w1875) | (w1874 & w1875);
assign w1668 = w1089 & w1065;
assign w1669 = (w1065 & w1089) | (w1065 & ~w736) | (w1089 & ~w736);
assign w1670 = (~w1065 & w1091) | (~w1065 & ~w741) | (w1091 & ~w741);
assign w1671 = (~w1065 & w1091) | (~w1065 & w1608) | (w1091 & w1608);
assign w1672 = ~w755 & w1643;
assign w1673 = (w1095 & w1876) | (w1095 & w1877) | (w1876 & w1877);
assign w1674 = (w1098 & w1879) | (w1098 & w1880) | (w1879 & w1880);
assign w1675 = (w1098 & w1881) | (w1098 & w1880) | (w1881 & w1880);
assign w1676 = w761 & w2857;
assign w1677 = (w1101 & w1885) | (w1101 & w1886) | (w1885 & w1886);
assign w1678 = ~w767 & w1645;
assign w1679 = w767 & ~w1645;
assign w1680 = ~w773 & w1649;
assign w1681 = ~w773 & w1648;
assign w1682 = ~w773 & w1647;
assign w1683 = w773 & ~w1649;
assign w1684 = w773 & ~w1648;
assign w1685 = ~w779 & w1651;
assign w1686 = ~w779 & w1650;
assign w1687 = w779 & ~w1651;
assign w1688 = w779 & ~w1650;
assign w1689 = (w1109 & w2374) | (w1109 & w2319) | (w2374 & w2319);
assign w1690 = (w1109 & w2375) | (w1109 & w2319) | (w2375 & w2319);
assign w1691 = w785 & ~w1108;
assign w1692 = (w785 & w1107) | (w785 & w2376) | (w1107 & w2376);
assign w1693 = (~w1109 & w2377) | (~w1109 & w1691) | (w2377 & w1691);
assign w1694 = (~w1109 & w2692) | (~w1109 & w1691) | (w2692 & w1691);
assign w1695 = ~w791 & w1654;
assign w1696 = ~w791 & w1653;
assign w1697 = (~w1103 & w2693) | (~w1103 & w2694) | (w2693 & w2694);
assign w1698 = (w1107 & w2378) | (w1107 & w2379) | (w2378 & w2379);
assign w1699 = w791 & ~w1654;
assign w1700 = w791 & ~w1653;
assign w1701 = (w1080 & w2695) | (w1080 & w2696) | (w2695 & w2696);
assign w1702 = (w1103 & w2697) | (w1103 & w2698) | (w2697 & w2698);
assign w1703 = ~w803 & w2858;
assign w1704 = (w2380 & w2381) | (w2380 & ~w1086) | (w2381 & ~w1086);
assign w1705 = w803 & w2963;
assign w1706 = w1043 & ~w617;
assign w1707 = (~w617 & w1043) | (~w617 & ~w610) | (w1043 & ~w610);
assign w1708 = w1045 & w1046;
assign w1709 = (w1046 & w1045) | (w1046 & ~w610) | (w1045 & ~w610);
assign w1710 = w1048 & w1049;
assign w1711 = (w1049 & w1048) | (w1049 & ~w610) | (w1048 & ~w610);
assign w1712 = (w1049 & w1048) | (w1049 & w1569) | (w1048 & w1569);
assign w1713 = (w1049 & w1048) | (w1049 & w1570) | (w1048 & w1570);
assign w1714 = w1052 & w1051;
assign w1715 = (w1051 & w1052) | (w1051 & ~w610) | (w1052 & ~w610);
assign w1716 = (w1051 & w1052) | (w1051 & w1569) | (w1052 & w1569);
assign w1717 = (w1051 & w1052) | (w1051 & w1570) | (w1052 & w1570);
assign w1718 = w1054 & w1053;
assign w1719 = (w1053 & w1054) | (w1053 & ~w610) | (w1054 & ~w610);
assign w1720 = (w1053 & w1054) | (w1053 & w1569) | (w1054 & w1569);
assign w1721 = (w1053 & w1054) | (w1053 & w1570) | (w1054 & w1570);
assign w1722 = w1056 & w1055;
assign w1723 = (w1055 & w1056) | (w1055 & ~w610) | (w1056 & ~w610);
assign w1724 = w1065 & w1041;
assign w1725 = (w1041 & w1065) | (w1041 & ~w675) | (w1065 & ~w675);
assign w1726 = ~w695 & w1658;
assign w1727 = ~w695 & w1657;
assign w1728 = ~w701 & w1661;
assign w1729 = ~w701 & w1660;
assign w1730 = w701 & ~w1660;
assign w1731 = (w1076 & w2382) | (w1076 & w2383) | (w2382 & w2383);
assign w1732 = (w1076 & w2384) | (w1076 & w2383) | (w2384 & w2383);
assign w1733 = ~w713 & w1663;
assign w1734 = ~w713 & w1662;
assign w1735 = w713 & ~w1663;
assign w1736 = w713 & ~w1662;
assign w1737 = ~w719 & w1665;
assign w1738 = w1870 & w2385;
assign w1739 = w719 & ~w1665;
assign w1740 = (w719 & ~w1870) | (w719 & w2386) | (~w1870 & w2386);
assign w1741 = ~w731 & w1084;
assign w1742 = ~w731 & w1085;
assign w1743 = (w1080 & w2699) | (w1080 & w2700) | (w2699 & w2700);
assign w1744 = (w1055 & w2701) | (w1055 & w2702) | (w2701 & w2702);
assign w1745 = (w2387 & w2388) | (w2387 & w2828) | (w2388 & w2828);
assign w1746 = (~w1080 & w2781) | (~w1080 & w2782) | (w2781 & w2782);
assign w1747 = w737 & w2931;
assign w1748 = w53 & ~w54;
assign w1749 = ~w75 & w74;
assign w1750 = ~w95 & ~w103;
assign w1751 = ~w103 & w1410;
assign w1752 = w95 & w103;
assign w1753 = w845 & ~w102;
assign w1754 = (~w102 & w845) | (~w102 & ~w95) | (w845 & ~w95);
assign w1755 = (~w102 & w845) | (~w102 & w1410) | (w845 & w1410);
assign w1756 = ~w120 & ~w128;
assign w1757 = ~w128 & w1415;
assign w1758 = w120 & w128;
assign w1759 = (~w127 & w855) | (~w127 & ~w120) | (w855 & ~w120);
assign w1760 = (~w127 & w855) | (~w127 & w1415) | (w855 & w1415);
assign w1761 = (w858 & w857) | (w858 & ~w120) | (w857 & ~w120);
assign w1762 = (w858 & w857) | (w858 & w1415) | (w857 & w1415);
assign w1763 = ~w153 & w152;
assign w1764 = ~w153 & ~w1421;
assign w1765 = (~w153 & w1420) | (~w153 & w1763) | (w1420 & w1763);
assign w1766 = ~w159 & w2859;
assign w1767 = ~w159 & w2860;
assign w1768 = w182 & ~w183;
assign w1769 = ~w189 & w2861;
assign w1770 = ~w189 & w2862;
assign w1771 = w881 | w880;
assign w1772 = (w880 & w881) | (w880 & w182) | (w881 & w182);
assign w1773 = ~w217 & ~w225;
assign w1774 = w217 & w225;
assign w1775 = (w893 & w892) | (w893 & ~w217) | (w892 & ~w217);
assign w1776 = (w893 & w892) | (w893 & w1439) | (w892 & w1439);
assign w1777 = (w896 & w895) | (w896 & ~w217) | (w895 & ~w217);
assign w1778 = (w896 & w895) | (w896 & w1439) | (w895 & w1439);
assign w1779 = ~w257 & ~w265;
assign w1780 = w257 & w265;
assign w1781 = w907 & w908;
assign w1782 = (w908 & w907) | (w908 & ~w257) | (w907 & ~w257);
assign w1783 = (w908 & w907) | (w908 & w1449) | (w907 & w1449);
assign w1784 = (w911 & w910) | (w911 & ~w257) | (w910 & ~w257);
assign w1785 = (w911 & w910) | (w911 & w1449) | (w910 & w1449);
assign w1786 = ~w300 & w299;
assign w1787 = ~w300 & ~w1458;
assign w1788 = (~w300 & w1457) | (~w300 & w1786) | (w1457 & w1786);
assign w1789 = ~w307 & w2863;
assign w1790 = ~w307 & w2864;
assign w1791 = (w926 & w927) | (w926 & ~w1458) | (w927 & ~w1458);
assign w1792 = (w926 & w927) | (w926 & ~w1459) | (w927 & ~w1459);
assign w1793 = (w933 & w932) | (w933 & w299) | (w932 & w299);
assign w1794 = (w933 & w932) | (w933 & ~w1458) | (w932 & ~w1458);
assign w1795 = ~w345 & w344;
assign w1796 = ~w345 & ~w1474;
assign w1797 = ~w388 & ~w396;
assign w1798 = w396 & ~w1491;
assign w1799 = w396 & ~w1492;
assign w1800 = w388 & w396;
assign w1801 = (~w395 & w959) | (~w395 & w1491) | (w959 & w1491);
assign w1802 = (w962 & w961) | (w962 & w1491) | (w961 & w1491);
assign w1803 = (w962 & w961) | (w962 & w1492) | (w961 & w1492);
assign w1804 = w964 & w965;
assign w1805 = (w965 & w964) | (w965 & ~w388) | (w964 & ~w388);
assign w1806 = ~w437 & ~w445;
assign w1807 = w445 & ~w1509;
assign w1808 = w445 & ~w1510;
assign w1809 = w437 & w445;
assign w1810 = (w988 & w989) | (w988 & w1509) | (w989 & w1509);
assign w1811 = (w988 & w989) | (w988 & w1510) | (w989 & w1510);
assign w1812 = (~w500 & w1526) | (~w500 & w1813) | (w1526 & w1813);
assign w1813 = w499 & ~w500;
assign w1814 = ~w507 & w2865;
assign w1815 = ~w507 & w2866;
assign w1816 = w1007 | w1006;
assign w1817 = (w1006 & w1007) | (w1006 & w499) | (w1007 & w499);
assign w1818 = ~w525 & w2867;
assign w1819 = ~w525 & w2868;
assign w1820 = (w1011 & w1010) | (w1011 & ~w1527) | (w1010 & ~w1527);
assign w1821 = (w1011 & w1010) | (w1011 & ~w1528) | (w1010 & ~w1528);
assign w1822 = w1010 | w1011;
assign w1823 = (w1011 & w1010) | (w1011 & w499) | (w1010 & w499);
assign w1824 = ~w555 & w554;
assign w1825 = ~w555 & ~w1547;
assign w1826 = (~w555 & w1546) | (~w555 & w1824) | (w1546 & w1824);
assign w1827 = ~w562 & w2869;
assign w1828 = (w1028 & w1029) | (w1028 & w554) | (w1029 & w554);
assign w1829 = (w1028 & w1029) | (w1028 & ~w1547) | (w1029 & ~w1547);
assign w1830 = (w1028 & w1029) | (w1028 & ~w1548) | (w1029 & ~w1548);
assign w1831 = ~w580 & w2870;
assign w1832 = ~w580 & w2871;
assign w1833 = (w1033 & w1032) | (w1033 & ~w1547) | (w1032 & ~w1547);
assign w1834 = (w1033 & w1032) | (w1033 & ~w1548) | (w1032 & ~w1548);
assign w1835 = ~w610 & ~w618;
assign w1836 = w610 & w618;
assign w1837 = w177 & ~w182;
assign w1838 = w210 & ~w216;
assign w1839 = w250 & ~w251;
assign w1840 = w287 & ~w288;
assign w1841 = w325 & ~w331;
assign w1842 = w337 & ~w338;
assign w1843 = w370 & ~w375;
assign w1844 = w381 & ~w382;
assign w1845 = w418 & ~w419;
assign w1846 = w430 & ~w431;
assign w1847 = w471 & ~w472;
assign w1848 = w485 & ~w486;
assign w1849 = w493 & ~w499;
assign w1850 = w525 & ~w530;
assign w1851 = w536 & ~w537;
assign w1852 = w543 & ~w548;
assign w1853 = w580 & ~w585;
assign w1854 = w591 & ~w592;
assign w1855 = w598 & ~w603;
assign w1856 = w609 & ~w610;
assign w1857 = w649 & ~w650;
assign w1858 = w662 & ~w663;
assign w1859 = w669 & ~w674;
assign w1860 = w711 & ~w712;
assign w1861 = w723 & ~w724;
assign w1862 = w730 & ~w735;
assign w1863 = w766 & ~w771;
assign w1864 = w777 & ~w778;
assign w1865 = w784 & ~w789;
assign w1866 = w795 & ~w796;
assign w1867 = w801 & ~w802;
assign w1868 = ~w809 & w1867;
assign w1869 = ~w807 & w802;
assign w1870 = (w1075 & w2389) | (w1075 & w2390) | (w2389 & w2390);
assign w1871 = (w1075 & w2391) | (w1075 & w2392) | (w2391 & w2392);
assign w1872 = (w1075 & w2393) | (w1075 & w2394) | (w2393 & w2394);
assign w1873 = ~w718 & w1083;
assign w1874 = w1083 & ~w675;
assign w1875 = (~w675 & w1083) | (~w675 & ~w718) | (w1083 & ~w718);
assign w1876 = ~w755 & ~w1608;
assign w1877 = ~w755 & w1094;
assign w1878 = ~w755 & w741;
assign w1879 = ~w761 & ~w1609;
assign w1880 = ~w761 & w1097;
assign w1881 = ~w761 & ~w1608;
assign w1882 = ~w761 & w741;
assign w1883 = w761 & w1609;
assign w1884 = w761 & ~w1097;
assign w1885 = ~w767 & ~w1609;
assign w1886 = (w1097 & w2395) | (w1097 & w2396) | (w2395 & w2396);
assign w1887 = (w835 & w834) | (w835 & w827) | (w834 & w827);
assign w1888 = (w835 & w834) | (w835 & w828) | (w834 & w828);
assign w1889 = (w854 & w853) | (w854 & w843) | (w853 & w843);
assign w1890 = (w854 & w853) | (w854 & w844) | (w853 & w844);
assign w1891 = (w876 & w875) | (w876 & w866) | (w875 & w866);
assign w1892 = (w876 & w875) | (w876 & w865) | (w875 & w865);
assign w1893 = (w903 & w904) | (w903 & w889) | (w904 & w889);
assign w1894 = (w903 & w904) | (w903 & w888) | (w904 & w888);
assign w1895 = (w939 & w940) | (w939 & w920) | (w940 & w920);
assign w1896 = (w939 & w940) | (w939 & w921) | (w940 & w921);
assign w1897 = (w958 & w957) | (w958 & ~w1896) | (w957 & ~w1896);
assign w1898 = (w958 & w957) | (w958 & ~w1895) | (w957 & ~w1895);
assign w1899 = (w998 & w997) | (w998 & ~w976) | (w997 & ~w976);
assign w1900 = (w998 & w997) | (w998 & ~w977) | (w997 & ~w977);
assign w1901 = (w1020 & w1019) | (w1020 & w1900) | (w1019 & w1900);
assign w1902 = (w1020 & w1019) | (w1020 & w1899) | (w1019 & w1899);
assign w1903 = (w1116 & w1117) | (w1116 & ~w1158) | (w1117 & ~w1158);
assign w1904 = (w1116 & w1117) | (w1116 & ~w1157) | (w1117 & ~w1157);
assign w1905 = (w1118 & w1119) | (w1118 & w1158) | (w1119 & w1158);
assign w1906 = (w1118 & w1119) | (w1118 & w1157) | (w1119 & w1157);
assign w1907 = (w1120 & w1121) | (w1120 & w1158) | (w1121 & w1158);
assign w1908 = (w1120 & w1121) | (w1120 & w1157) | (w1121 & w1157);
assign w1909 = (~w256 & w1448) | (~w256 & ~w250) | (w1448 & ~w250);
assign w1910 = (~w256 & w1448) | (~w256 & w1445) | (w1448 & w1445);
assign w1911 = (~w293 & w1456) | (~w293 & ~w287) | (w1456 & ~w287);
assign w1912 = (~w293 & w1456) | (~w293 & w1453) | (w1456 & w1453);
assign w1913 = (~w337 & w1469) | (~w337 & w1467) | (w1469 & w1467);
assign w1914 = (~w337 & w1469) | (~w337 & w1466) | (w1469 & w1466);
assign w1915 = (~w424 & w1501) | (~w424 & ~w418) | (w1501 & ~w418);
assign w1916 = (~w424 & w1501) | (~w424 & w1498) | (w1501 & w1498);
assign w1917 = (~w478 & w1519) | (~w478 & ~w471) | (w1519 & ~w471);
assign w1918 = (~w478 & w1519) | (~w478 & w1516) | (w1519 & w1516);
assign w1919 = (~w493 & w1523) | (~w493 & w1526) | (w1523 & w1526);
assign w1920 = ~w493 & ~w1524;
assign w1921 = (~w649 & w1577) | (~w649 & ~w642) | (w1577 & ~w642);
assign w1922 = (~w649 & w1577) | (~w649 & w1575) | (w1577 & w1575);
assign w1923 = (~w711 & w1594) | (~w711 & ~w705) | (w1594 & ~w705);
assign w1924 = (~w711 & w1594) | (~w711 & w1592) | (w1594 & w1592);
assign w1925 = (~w777 & w1617) | (~w777 & w1615) | (w1617 & w1615);
assign w1926 = (~w777 & w1617) | (~w777 & w1614) | (w1617 & w1614);
assign w1927 = (~w1895 & w2397) | (~w1895 & w2398) | (w2397 & w2398);
assign w1928 = (~w1896 & w2397) | (~w1896 & w2398) | (w2397 & w2398);
assign w1929 = (w1900 & w1899) | (w1900 & ~w1898) | (w1899 & ~w1898);
assign w1930 = (w1900 & w1899) | (w1900 & ~w1897) | (w1899 & ~w1897);
assign w1931 = (~w1899 & w2399) | (~w1899 & w2400) | (w2399 & w2400);
assign w1932 = (~w1900 & w2399) | (~w1900 & w2400) | (w2399 & w2400);
assign w1933 = (~w1899 & w2401) | (~w1899 & w2402) | (w2401 & w2402);
assign w1934 = (~w1900 & w2401) | (~w1900 & w2402) | (w2401 & w2402);
assign w1935 = (~w1899 & w2403) | (~w1899 & w2404) | (w2403 & w2404);
assign w1936 = (~w1900 & w2403) | (~w1900 & w2404) | (w2403 & w2404);
assign w1937 = (~w1899 & w2405) | (~w1899 & w2406) | (w2405 & w2406);
assign w1938 = (~w1900 & w2405) | (~w1900 & w2406) | (w2405 & w2406);
assign w1939 = (~w1899 & w2407) | (~w1899 & w2408) | (w2407 & w2408);
assign w1940 = (~w1900 & w2407) | (~w1900 & w2408) | (w2407 & w2408);
assign w1941 = (~w1899 & w2409) | (~w1899 & w2410) | (w2409 & w2410);
assign w1942 = (~w1900 & w2409) | (~w1900 & w2410) | (w2409 & w2410);
assign w1943 = (~w1899 & w2411) | (~w1899 & w2412) | (w2411 & w2412);
assign w1944 = (~w1900 & w2411) | (~w1900 & w2412) | (w2411 & w2412);
assign w1945 = (w1041 & w2413) | (w1041 & w2414) | (w2413 & w2414);
assign w1946 = ~w664 & w1216;
assign w1947 = (~w1041 & w2415) | (~w1041 & w2416) | (w2415 & w2416);
assign w1948 = w664 & ~w1216;
assign w1949 = (w1041 & w2417) | (w1041 & w2418) | (w2417 & w2418);
assign w1950 = ~w670 & w1217;
assign w1951 = (~w1041 & w2419) | (~w1041 & w2420) | (w2419 & w2420);
assign w1952 = w670 & ~w1217;
assign w1953 = ~w676 & w1218;
assign w1954 = (w1063 & w2421) | (w1063 & w2422) | (w2421 & w2422);
assign w1955 = w676 & ~w1218;
assign w1956 = (~w1063 & w2423) | (~w1063 & w2424) | (w2423 & w2424);
assign w1957 = ~w683 & w1220;
assign w1958 = (w1065 & w2425) | (w1065 & w2426) | (w2425 & w2426);
assign w1959 = w683 & ~w1220;
assign w1960 = (~w1065 & w2427) | (~w1065 & w2428) | (w2427 & w2428);
assign w1961 = (w1159 & w1160) | (w1159 & w1220) | (w1160 & w1220);
assign w1962 = (w1159 & w1160) | (w1159 & w1219) | (w1160 & w1219);
assign w1963 = (w1161 & w1162) | (w1161 & ~w1220) | (w1162 & ~w1220);
assign w1964 = (w1161 & w1162) | (w1161 & ~w1219) | (w1162 & ~w1219);
assign w1965 = (w1163 & w1164) | (w1163 & w1220) | (w1164 & w1220);
assign w1966 = (w1163 & w1164) | (w1163 & w1219) | (w1164 & w1219);
assign w1967 = (w1165 & w1166) | (w1165 & ~w1220) | (w1166 & ~w1220);
assign w1968 = (w1165 & w1166) | (w1165 & ~w1219) | (w1166 & ~w1219);
assign w1969 = (w1167 & w1168) | (w1167 & w1220) | (w1168 & w1220);
assign w1970 = (w1167 & w1168) | (w1167 & w1219) | (w1168 & w1219);
assign w1971 = (w1169 & w1170) | (w1169 & ~w1220) | (w1170 & ~w1220);
assign w1972 = (w1169 & w1170) | (w1169 & ~w1219) | (w1170 & ~w1219);
assign w1973 = (w1171 & w1172) | (w1171 & w1220) | (w1172 & w1220);
assign w1974 = (w1171 & w1172) | (w1171 & w1219) | (w1172 & w1219);
assign w1975 = (w1173 & w1174) | (w1173 & ~w1220) | (w1174 & ~w1220);
assign w1976 = (w1173 & w1174) | (w1173 & ~w1219) | (w1174 & ~w1219);
assign w1977 = (w1175 & w1176) | (w1175 & w1220) | (w1176 & w1220);
assign w1978 = (w1175 & w1176) | (w1175 & w1219) | (w1176 & w1219);
assign w1979 = (w1177 & w1178) | (w1177 & ~w1220) | (w1178 & ~w1220);
assign w1980 = (w1177 & w1178) | (w1177 & ~w1219) | (w1178 & ~w1219);
assign w1981 = (w1180 & w1179) | (w1180 & w1220) | (w1179 & w1220);
assign w1982 = (w1180 & w1179) | (w1180 & w1219) | (w1179 & w1219);
assign w1983 = (w1182 & w1181) | (w1182 & ~w1220) | (w1181 & ~w1220);
assign w1984 = (w1182 & w1181) | (w1182 & ~w1219) | (w1181 & ~w1219);
assign w1985 = (w1184 & w1183) | (w1184 & w1220) | (w1183 & w1220);
assign w1986 = (w1184 & w1183) | (w1184 & w1219) | (w1183 & w1219);
assign w1987 = (w1186 & w1185) | (w1186 & ~w1220) | (w1185 & ~w1220);
assign w1988 = (w1186 & w1185) | (w1186 & ~w1219) | (w1185 & ~w1219);
assign w1989 = (w1188 & w1187) | (w1188 & w1220) | (w1187 & w1220);
assign w1990 = (w1188 & w1187) | (w1188 & w1219) | (w1187 & w1219);
assign w1991 = (w1189 & w1190) | (w1189 & ~w1220) | (w1190 & ~w1220);
assign w1992 = (w1189 & w1190) | (w1189 & ~w1219) | (w1190 & ~w1219);
assign w1993 = (w1196 & w1195) | (w1196 & w1220) | (w1195 & w1220);
assign w1994 = (w1196 & w1195) | (w1196 & w1219) | (w1195 & w1219);
assign w1995 = ~w827 & w2429;
assign w1996 = (w826 & w2429) | (w826 & w2430) | (w2429 & w2430);
assign w1997 = (w62 & w827) | (w62 & w2431) | (w827 & w2431);
assign w1998 = w62 & w2872;
assign w1999 = (w1276 & w1275) | (w1276 & ~w827) | (w1275 & ~w827);
assign w2000 = (w1276 & w1275) | (w1276 & ~w828) | (w1275 & ~w828);
assign w2001 = (w834 & w2432) | (w834 & w2433) | (w2432 & w2433);
assign w2002 = (w835 & w2432) | (w835 & w2433) | (w2432 & w2433);
assign w2003 = w96 & ~w1278;
assign w2004 = w96 & ~w1277;
assign w2005 = w109 & ~w1283;
assign w2006 = (w842 & w2434) | (w842 & w2435) | (w2434 & w2435);
assign w2007 = (w843 & w2703) | (w843 & w2704) | (w2703 & w2704);
assign w2008 = ~w115 & w1284;
assign w2009 = w115 & w2874;
assign w2010 = w115 & ~w1284;
assign w2011 = w121 & ~w1286;
assign w2012 = w121 & ~w1285;
assign w2013 = (w1290 & w1289) | (w1290 & ~w844) | (w1289 & ~w844);
assign w2014 = (w1290 & w1289) | (w1290 & ~w843) | (w1289 & ~w843);
assign w2015 = ~w148 & w1295;
assign w2016 = (w854 & w2436) | (w854 & w2437) | (w2436 & w2437);
assign w2017 = w148 & ~w1295;
assign w2018 = (~w854 & w2438) | (~w854 & w2439) | (w2438 & w2439);
assign w2019 = (w864 & w2705) | (w864 & w2706) | (w2705 & w2706);
assign w2020 = ~w154 & w1296;
assign w2021 = (w860 & w2440) | (w860 & w2441) | (w2440 & w2441);
assign w2022 = ~w160 & w2876;
assign w2023 = w160 & w2877;
assign w2024 = (w862 & w2707) | (w862 & w2442) | (w2707 & w2442);
assign w2025 = ~w166 & w1298;
assign w2026 = ~w166 & w1297;
assign w2027 = (~w865 & w2443) | (~w865 & w2444) | (w2443 & w2444);
assign w2028 = (~w866 & w2443) | (~w866 & w2444) | (w2443 & w2444);
assign w2029 = (~w865 & w2446) | (~w865 & w2447) | (w2446 & w2447);
assign w2030 = (~w866 & w2446) | (~w866 & w2447) | (w2446 & w2447);
assign w2031 = (w865 & w2448) | (w865 & w2449) | (w2448 & w2449);
assign w2032 = (w866 & w2448) | (w866 & w2709) | (w2448 & w2709);
assign w2033 = ~w184 & w1300;
assign w2034 = ~w184 & w1299;
assign w2035 = (w1302 & w1301) | (w1302 & ~w866) | (w1301 & ~w866);
assign w2036 = (w1302 & w1301) | (w1302 & ~w865) | (w1301 & ~w865);
assign w2037 = (w1304 & w1303) | (w1304 & ~w866) | (w1303 & ~w866);
assign w2038 = (w1304 & w1303) | (w1304 & ~w865) | (w1303 & ~w865);
assign w2039 = (w1306 & w1305) | (w1306 & ~w866) | (w1305 & ~w866);
assign w2040 = (w1306 & w1305) | (w1306 & ~w865) | (w1305 & ~w865);
assign w2041 = (w884 & w883) | (w884 & ~w1891) | (w883 & ~w1891);
assign w2042 = (w884 & w883) | (w884 & ~w1892) | (w883 & ~w1892);
assign w2043 = ~w210 & w2964;
assign w2044 = ~w210 & w2965;
assign w2045 = (w889 & w888) | (w889 & ~w1892) | (w888 & ~w1892);
assign w2046 = (w889 & w888) | (w889 & ~w1891) | (w888 & ~w1891);
assign w2047 = (w1308 & w1307) | (w1308 & ~w1892) | (w1307 & ~w1892);
assign w2048 = (w1308 & w1307) | (w1308 & ~w1891) | (w1307 & ~w1891);
assign w2049 = (~w224 & w890) | (~w224 & w2966) | (w890 & w2966);
assign w2050 = (~w224 & w890) | (~w224 & w2967) | (w890 & w2967);
assign w2051 = (w1312 & w1311) | (w1312 & ~w1892) | (w1311 & ~w1892);
assign w2052 = (w1312 & w1311) | (w1312 & ~w1891) | (w1311 & ~w1891);
assign w2053 = (w1314 & w1313) | (w1314 & ~w1892) | (w1313 & ~w1892);
assign w2054 = (w1314 & w1313) | (w1314 & ~w1891) | (w1313 & ~w1891);
assign w2055 = w252 & ~w1316;
assign w2056 = w252 & ~w1315;
assign w2057 = w258 & ~w1318;
assign w2058 = w258 & ~w1317;
assign w2059 = ~w271 & w1324;
assign w2060 = ~w271 & w1323;
assign w2061 = (w900 & w2450) | (w900 & w2451) | (w2450 & w2451);
assign w2062 = ~w277 & w2878;
assign w2063 = w277 & w2879;
assign w2064 = (w902 & w2452) | (w902 & w2710) | (w2452 & w2710);
assign w2065 = ~w283 & w1326;
assign w2066 = ~w283 & w1325;
assign w2067 = ~w289 & w1328;
assign w2068 = ~w289 & w1327;
assign w2069 = ~w295 & w1330;
assign w2070 = ~w295 & w1329;
assign w2071 = ~w301 & w1332;
assign w2072 = ~w301 & w1331;
assign w2073 = (w921 & w920) | (w921 & ~w1894) | (w920 & ~w1894);
assign w2074 = (w921 & w920) | (w921 & ~w1893) | (w920 & ~w1893);
assign w2075 = (w1336 & w1335) | (w1336 & w1894) | (w1335 & w1894);
assign w2076 = (w1336 & w1335) | (w1336 & w1893) | (w1335 & w1893);
assign w2077 = (w1338 & w1337) | (w1338 & w1894) | (w1337 & w1894);
assign w2078 = (w1338 & w1337) | (w1338 & w1893) | (w1337 & w1893);
assign w2079 = (w1340 & w1339) | (w1340 & w1894) | (w1339 & w1894);
assign w2080 = (w1340 & w1339) | (w1340 & w1893) | (w1339 & w1893);
assign w2081 = (w1342 & w1341) | (w1342 & w1894) | (w1341 & w1894);
assign w2082 = (w1342 & w1341) | (w1342 & w1893) | (w1341 & w1893);
assign w2083 = (w935 & w934) | (w935 & ~w2073) | (w934 & ~w2073);
assign w2084 = (w935 & w934) | (w935 & ~w2074) | (w934 & ~w2074);
assign w2085 = (w938 & w937) | (w938 & ~w2073) | (w937 & ~w2073);
assign w2086 = (w938 & w937) | (w938 & ~w2074) | (w937 & ~w2074);
assign w2087 = (w939 & w940) | (w939 & w2073) | (w940 & w2073);
assign w2088 = (w939 & w940) | (w939 & w2074) | (w940 & w2074);
assign w2089 = ~w353 & w2880;
assign w2090 = (w932 & w2711) | (w932 & w2712) | (w2711 & w2712);
assign w2091 = (w936 & w2454) | (w936 & w2455) | (w2454 & w2455);
assign w2092 = (~w932 & w2713) | (~w932 & w2714) | (w2713 & w2714);
assign w2093 = (w943 & w2560) | (w943 & w2881) | (w2560 & w2881);
assign w2094 = ~w359 & w1343;
assign w2095 = (w936 & w2456) | (w936 & w2457) | (w2456 & w2457);
assign w2096 = w359 & ~w1343;
assign w2097 = ~w365 & w1344;
assign w2098 = ~w365 & w1345;
assign w2099 = ~w371 & w1347;
assign w2100 = ~w371 & w1346;
assign w2101 = (~w939 & w2458) | (~w939 & w2459) | (w2458 & w2459);
assign w2102 = ~w377 & w1348;
assign w2103 = (w939 & w2460) | (w939 & w2461) | (w2460 & w2461);
assign w2104 = w377 & ~w1348;
assign w2105 = ~w383 & w2968;
assign w2106 = ~w383 & w2969;
assign w2107 = ~w389 & w1350;
assign w2108 = ~w389 & w1349;
assign w2109 = w389 & ~w1350;
assign w2110 = w389 & ~w1349;
assign w2111 = ~w402 & w1355;
assign w2112 = (~w953 & w2463) | (~w953 & w2464) | (w2463 & w2464);
assign w2113 = w402 & ~w1355;
assign w2114 = (w953 & w2465) | (w953 & w2466) | (w2465 & w2466);
assign w2115 = ~w408 & w1356;
assign w2116 = ~w408 & w2882;
assign w2117 = w408 & ~w1356;
assign w2118 = (w953 & w2467) | (w953 & w2468) | (w2467 & w2468);
assign w2119 = ~w414 & w2883;
assign w2120 = ~w414 & w1357;
assign w2121 = (w956 & w2469) | (w956 & w2470) | (w2469 & w2470);
assign w2122 = w414 & ~w1357;
assign w2123 = ~w420 & w1359;
assign w2124 = ~w420 & w1358;
assign w2125 = w420 & ~w1359;
assign w2126 = w420 & ~w1358;
assign w2127 = (w957 & w2471) | (w957 & w2472) | (w2471 & w2472);
assign w2128 = (w958 & w2471) | (w958 & w2472) | (w2471 & w2472);
assign w2129 = (~w957 & w2716) | (~w957 & w2473) | (w2716 & w2473);
assign w2130 = (~w958 & w2716) | (~w958 & w2717) | (w2716 & w2717);
assign w2131 = (w957 & w2474) | (w957 & w2475) | (w2474 & w2475);
assign w2132 = (w958 & w2474) | (w958 & w2475) | (w2474 & w2475);
assign w2133 = w432 & w2884;
assign w2134 = w432 & w2885;
assign w2135 = ~w438 & w1361;
assign w2136 = ~w438 & w1360;
assign w2137 = w438 & ~w1361;
assign w2138 = w438 & ~w1360;
assign w2139 = (w1363 & w1362) | (w1363 & w1898) | (w1362 & w1898);
assign w2140 = (w1363 & w1362) | (w1363 & w1897) | (w1362 & w1897);
assign w2141 = (~w1895 & w2478) | (~w1895 & w2479) | (w2478 & w2479);
assign w2142 = (~w1896 & w2478) | (~w1896 & w2479) | (w2478 & w2479);
assign w2143 = (~w1895 & w2480) | (~w1895 & w2481) | (w2480 & w2481);
assign w2144 = (~w1896 & w2480) | (~w1896 & w2481) | (w2480 & w2481);
assign w2145 = (w1371 & w1370) | (w1371 & w1898) | (w1370 & w1898);
assign w2146 = (w1371 & w1370) | (w1371 & w1897) | (w1370 & w1897);
assign w2147 = (w1373 & w1372) | (w1373 & w1898) | (w1372 & w1898);
assign w2148 = (w1373 & w1372) | (w1373 & w1897) | (w1372 & w1897);
assign w2149 = (w1375 & w1374) | (w1375 & w1898) | (w1374 & w1898);
assign w2150 = (w1375 & w1374) | (w1375 & w1897) | (w1374 & w1897);
assign w2151 = (w1377 & w1376) | (w1377 & w1898) | (w1376 & w1898);
assign w2152 = (w1377 & w1376) | (w1377 & w1897) | (w1376 & w1897);
assign w2153 = (w1379 & w1378) | (w1379 & w1898) | (w1378 & w1898);
assign w2154 = (w1379 & w1378) | (w1379 & w1897) | (w1378 & w1897);
assign w2155 = (w1381 & w1380) | (w1381 & w1898) | (w1380 & w1898);
assign w2156 = (w1381 & w1380) | (w1381 & w1897) | (w1380 & w1897);
assign w2157 = (w988 & w2718) | (w988 & w2719) | (w2718 & w2719);
assign w2158 = (~w992 & w2483) | (~w992 & w2484) | (w2483 & w2484);
assign w2159 = w508 & w2970;
assign w2160 = (w992 & w2720) | (w992 & w2721) | (w2720 & w2721);
assign w2161 = (w988 & w2783) | (w988 & w2784) | (w2783 & w2784);
assign w2162 = ~w514 & w2886;
assign w2163 = (w2489 & w2488) | (w2489 & ~w995) | (w2488 & ~w995);
assign w2164 = (w992 & w2722) | (w992 & w2723) | (w2722 & w2723);
assign w2165 = (w995 & w2490) | (w995 & w2491) | (w2490 & w2491);
assign w2166 = ~w520 & w1382;
assign w2167 = (w2579 & ~w1004) | (w2579 & w2887) | (~w1004 & w2887);
assign w2168 = w520 & ~w1382;
assign w2169 = (w995 & w2492) | (w995 & w2493) | (w2492 & w2493);
assign w2170 = ~w526 & w1383;
assign w2171 = ~w532 & w1385;
assign w2172 = ~w532 & w1384;
assign w2173 = ~w538 & w1387;
assign w2174 = ~w538 & w1386;
assign w2175 = (~w997 & w2494) | (~w997 & w2495) | (w2494 & w2495);
assign w2176 = ~w544 & w1388;
assign w2177 = (w997 & w2496) | (w997 & w2497) | (w2496 & w2497);
assign w2178 = w544 & ~w1388;
assign w2179 = (~w997 & w2498) | (~w997 & w2499) | (w2498 & w2499);
assign w2180 = ~w550 & w1389;
assign w2181 = (w997 & w2500) | (w997 & w2501) | (w2500 & w2501);
assign w2182 = w550 & ~w1389;
assign w2183 = ~w556 & w1390;
assign w2184 = (w1017 & w2502) | (w1017 & w2503) | (w2502 & w2503);
assign w2185 = w556 & ~w1390;
assign w2186 = (~w1017 & w2504) | (~w1017 & w2505) | (w2504 & w2505);
assign w2187 = ~w563 & w1391;
assign w2188 = ~w563 & w2889;
assign w2189 = w563 & w2971;
assign w2190 = (w1012 & w2506) | (w1012 & w2507) | (w2506 & w2507);
assign w2191 = ~w569 & w1393;
assign w2192 = ~w569 & w1392;
assign w2193 = w569 & w2972;
assign w2194 = w569 & ~w1392;
assign w2195 = (w1015 & w2508) | (w1015 & w2509) | (w2508 & w2509);
assign w2196 = (w1026 & w2598) | (w1026 & w2890) | (w2598 & w2890);
assign w2197 = (~w1026 & w2600) | (~w1026 & w2891) | (w2600 & w2891);
assign w2198 = (w1016 & w2510) | (w1016 & w2724) | (w2510 & w2724);
assign w2199 = (w1015 & w2511) | (w1015 & w2512) | (w2511 & w2512);
assign w2200 = ~w581 & w2892;
assign w2201 = w581 & w2893;
assign w2202 = (w1016 & w2513) | (w1016 & w2725) | (w2513 & w2725);
assign w2203 = ~w587 & w1395;
assign w2204 = ~w587 & w1394;
assign w2205 = w587 & ~w1395;
assign w2206 = w587 & ~w1394;
assign w2207 = ~w593 & w1397;
assign w2208 = ~w593 & w1396;
assign w2209 = w593 & ~w1397;
assign w2210 = w593 & ~w1396;
assign w2211 = (~w1019 & w2514) | (~w1019 & w2515) | (w2514 & w2515);
assign w2212 = ~w599 & w1398;
assign w2213 = (w1019 & w2516) | (w1019 & w2517) | (w2516 & w2517);
assign w2214 = w599 & ~w1398;
assign w2215 = (~w1019 & w2518) | (~w1019 & w2519) | (w2518 & w2519);
assign w2216 = ~w605 & w1399;
assign w2217 = (w1019 & w2520) | (w1019 & w2521) | (w2520 & w2521);
assign w2218 = w605 & ~w1399;
assign w2219 = ~w611 & w1400;
assign w2220 = (w1038 & w2522) | (w1038 & w2523) | (w2522 & w2523);
assign w2221 = w611 & ~w1400;
assign w2222 = (~w1038 & w2524) | (~w1038 & w2525) | (w2524 & w2525);
assign w2223 = (w1401 & w1402) | (w1401 & ~w1902) | (w1402 & ~w1902);
assign w2224 = (w1401 & w1402) | (w1401 & ~w1901) | (w1402 & ~w1901);
assign w2225 = w1439 & ~w217;
assign w2226 = (~w217 & w1439) | (~w217 & ~w210) | (w1439 & ~w210);
assign w2227 = ~w217 & ~w1438;
assign w2228 = (~w217 & w1436) | (~w217 & w1439) | (w1436 & w1439);
assign w2229 = (~w257 & w1449) | (~w257 & w1447) | (w1449 & w1447);
assign w2230 = (~w257 & w1449) | (~w257 & w1446) | (w1449 & w1446);
assign w2231 = ~w257 & ~w1910;
assign w2232 = ~w257 & ~w1909;
assign w2233 = (~w294 & w1457) | (~w294 & w1455) | (w1457 & w1455);
assign w2234 = (~w294 & w1457) | (~w294 & w1454) | (w1457 & w1454);
assign w2235 = (~w299 & w1458) | (~w299 & w1912) | (w1458 & w1912);
assign w2236 = (~w299 & w1458) | (~w299 & w1911) | (w1458 & w1911);
assign w2237 = ~w332 & ~w1467;
assign w2238 = (~w332 & w1465) | (~w332 & w1468) | (w1465 & w1468);
assign w2239 = w1484 & ~w376;
assign w2240 = (~w376 & w1484) | (~w376 & ~w370) | (w1484 & ~w370);
assign w2241 = ~w376 & ~w1483;
assign w2242 = (~w376 & w1480) | (~w376 & w1484) | (w1480 & w1484);
assign w2243 = (~w381 & w1485) | (~w381 & w1483) | (w1485 & w1483);
assign w2244 = (~w381 & w1485) | (~w381 & w1482) | (w1485 & w1482);
assign w2245 = (~w388 & w1487) | (~w388 & w1491) | (w1487 & w1491);
assign w2246 = ~w388 & ~w1488;
assign w2247 = (~w425 & w1502) | (~w425 & w1500) | (w1502 & w1500);
assign w2248 = (~w425 & w1502) | (~w425 & w1499) | (w1502 & w1499);
assign w2249 = (~w430 & w1503) | (~w430 & w1916) | (w1503 & w1916);
assign w2250 = (~w430 & w1503) | (~w430 & w1915) | (w1503 & w1915);
assign w2251 = (~w437 & w1505) | (~w437 & w1509) | (w1505 & w1509);
assign w2252 = ~w437 & ~w1506;
assign w2253 = (~w479 & w1520) | (~w479 & w1518) | (w1520 & w1518);
assign w2254 = (~w479 & w1520) | (~w479 & w1517) | (w1520 & w1517);
assign w2255 = (~w485 & w1521) | (~w485 & w1918) | (w1521 & w1918);
assign w2256 = (~w485 & w1521) | (~w485 & w1917) | (w1521 & w1917);
assign w2257 = ~w531 & ~w1535;
assign w2258 = (~w531 & w1533) | (~w531 & w1536) | (w1533 & w1536);
assign w2259 = (~w536 & w1537) | (~w536 & w1535) | (w1537 & w1535);
assign w2260 = (~w536 & w1537) | (~w536 & w1534) | (w1537 & w1534);
assign w2261 = (~w543 & w1539) | (~w543 & w1542) | (w1539 & w1542);
assign w2262 = ~w543 & ~w1540;
assign w2263 = ~w549 & ~w1545;
assign w2264 = (~w549 & w1542) | (~w549 & w1546) | (w1542 & w1546);
assign w2265 = (~w554 & w1547) | (~w554 & w1545) | (w1547 & w1545);
assign w2266 = (~w554 & w1547) | (~w554 & w1544) | (w1547 & w1544);
assign w2267 = ~w586 & ~w1556;
assign w2268 = (~w586 & w1554) | (~w586 & w1557) | (w1554 & w1557);
assign w2269 = (~w591 & w1558) | (~w591 & w1556) | (w1558 & w1556);
assign w2270 = (~w591 & w1558) | (~w591 & w1555) | (w1558 & w1555);
assign w2271 = (~w598 & w1560) | (~w598 & w1563) | (w1560 & w1563);
assign w2272 = ~w598 & ~w1561;
assign w2273 = ~w604 & ~w1566;
assign w2274 = (~w604 & w1563) | (~w604 & w1567) | (w1563 & w1567);
assign w2275 = (~w609 & w1568) | (~w609 & w1566) | (w1568 & w1566);
assign w2276 = (~w609 & w1568) | (~w609 & w1565) | (w1568 & w1565);
assign w2277 = ~w610 & ~w2276;
assign w2278 = ~w610 & ~w2275;
assign w2279 = ~w643 & ~w1575;
assign w2280 = ~w650 & ~w1922;
assign w2281 = ~w650 & ~w1921;
assign w2282 = (~w656 & w1580) | (~w656 & w1922) | (w1580 & w1922);
assign w2283 = (~w656 & w1580) | (~w656 & w1921) | (w1580 & w1921);
assign w2284 = (w1584 & w1583) | (w1584 & w1579) | (w1583 & w1579);
assign w2285 = (w1584 & w1583) | (w1584 & w1578) | (w1583 & w1578);
assign w2286 = (~w669 & w1584) | (~w669 & w1587) | (w1584 & w1587);
assign w2287 = ~w669 & ~w1585;
assign w2288 = (w1590 & w1589) | (w1590 & ~w662) | (w1589 & ~w662);
assign w2289 = (w1590 & w1589) | (w1590 & w1582) | (w1589 & w1582);
assign w2290 = ~w706 & ~w1592;
assign w2291 = ~w712 & ~w1924;
assign w2292 = ~w712 & ~w1923;
assign w2293 = (~w717 & w1596) | (~w717 & w1924) | (w1596 & w1924);
assign w2294 = (~w717 & w1596) | (~w717 & w1923) | (w1596 & w1923);
assign w2295 = (~w718 & w1597) | (~w718 & w1595) | (w1597 & w1595);
assign w2296 = (~w718 & w1597) | (~w718 & w2390) | (w1597 & w2390);
assign w2297 = (w1600 & w1599) | (w1600 & w1595) | (w1599 & w1595);
assign w2298 = (w1600 & w1599) | (w1600 & w2390) | (w1599 & w2390);
assign w2299 = (~w730 & w1600) | (~w730 & w1603) | (w1600 & w1603);
assign w2300 = ~w730 & ~w1601;
assign w2301 = (w1606 & w1605) | (w1606 & ~w723) | (w1605 & ~w723);
assign w2302 = (w1606 & w1605) | (w1606 & w1598) | (w1605 & w1598);
assign w2303 = (~w741 & w1608) | (~w741 & w2302) | (w1608 & w2302);
assign w2304 = (~w741 & w1608) | (~w741 & w2301) | (w1608 & w2301);
assign w2305 = ~w772 & ~w1615;
assign w2306 = (~w772 & w1613) | (~w772 & w1616) | (w1613 & w1616);
assign w2307 = (~w784 & w1619) | (~w784 & w1622) | (w1619 & w1622);
assign w2308 = ~w784 & ~w1620;
assign w2309 = ~w790 & ~w1625;
assign w2310 = (~w790 & w1622) | (~w790 & w1626) | (w1622 & w1626);
assign w2311 = ~w796 & w2894;
assign w2312 = ~w796 & w2895;
assign w2313 = (w1624 & w2528) | (w1624 & w2529) | (w2528 & w2529);
assign w2314 = (w1625 & w2528) | (w1625 & w2529) | (w2528 & w2529);
assign w2315 = (w1081 & w1080) | (w1081 & ~w675) | (w1080 & ~w675);
assign w2316 = (w1081 & w1080) | (w1081 & w1591) | (w1080 & w1591);
assign w2317 = w761 & w2896;
assign w2318 = w767 & ~w1644;
assign w2319 = ~w785 & w1108;
assign w2320 = ~w1107 & w2530;
assign w2321 = (w1103 & w2531) | (w1103 & w2532) | (w2531 & w2532);
assign w2322 = ~w791 & w1111;
assign w2323 = w803 & w1092;
assign w2324 = (w1107 & w2534) | (w1107 & w2535) | (w2534 & w2535);
assign w2325 = (w1056 & w1055) | (w1056 & w1570) | (w1055 & w1570);
assign w2326 = (w1056 & w1055) | (w1056 & w1569) | (w1055 & w1569);
assign w2327 = w701 & ~w1659;
assign w2328 = ~w725 & w1083;
assign w2329 = ~w1082 & w2536;
assign w2330 = w725 & ~w1083;
assign w2331 = (w725 & w1082) | (w725 & w2537) | (w1082 & w2537);
assign w2332 = w1741 & w1085;
assign w2333 = (w1085 & w1741) | (w1085 & ~w731) | (w1741 & ~w731);
assign w2334 = w737 & ~w1066;
assign w2335 = ~w743 & w1066;
assign w2336 = ~w743 & w1090;
assign w2337 = w743 & ~w1066;
assign w2338 = w743 & ~w1090;
assign w2339 = ~w183 & ~w1430;
assign w2340 = (~w183 & w1428) | (~w183 & w1768) | (w1428 & w1768);
assign w2341 = (w225 & w1774) | (w225 & w1438) | (w1774 & w1438);
assign w2342 = (w225 & w1774) | (w225 & w1437) | (w1774 & w1437);
assign w2343 = w225 & ~w2225;
assign w2344 = w225 & ~w2226;
assign w2345 = ~w265 & w2229;
assign w2346 = ~w265 & w2230;
assign w2347 = (w265 & w1780) | (w265 & w1910) | (w1780 & w1910);
assign w2348 = (w265 & w1780) | (w265 & w1909) | (w1780 & w1909);
assign w2349 = (~w264 & w905) | (~w264 & w2229) | (w905 & w2229);
assign w2350 = (~w264 & w905) | (~w264 & w2230) | (w905 & w2230);
assign w2351 = ~w352 & w2973;
assign w2352 = ~w352 & w2897;
assign w2353 = (w945 & w946) | (w945 & ~w1473) | (w946 & ~w1473);
assign w2354 = (w945 & w946) | (w945 & ~w1472) | (w946 & ~w1472);
assign w2355 = (w949 & w948) | (w949 & ~w1473) | (w948 & ~w1473);
assign w2356 = (w949 & w948) | (w949 & ~w1472) | (w948 & ~w1472);
assign w2357 = w1797 & ~w1489;
assign w2358 = w1797 & ~w1488;
assign w2359 = (~w395 & w959) | (~w395 & w2898) | (w959 & w2898);
assign w2360 = (~w395 & w959) | (~w395 & w2246) | (w959 & w2246);
assign w2361 = (w962 & w961) | (w962 & w2898) | (w961 & w2898);
assign w2362 = (w962 & w961) | (w962 & w2246) | (w961 & w2246);
assign w2363 = w1806 & ~w1507;
assign w2364 = w1806 & ~w1506;
assign w2365 = (~w444 & w978) | (~w444 & w2899) | (w978 & w2899);
assign w2366 = (~w444 & w978) | (~w444 & w2252) | (w978 & w2252);
assign w2367 = (w981 & w980) | (w981 & w2899) | (w980 & w2899);
assign w2368 = (w981 & w980) | (w981 & w2252) | (w980 & w2252);
assign w2369 = ~w555 & ~w2265;
assign w2370 = ~w555 & ~w2266;
assign w2371 = (w618 & w1836) | (w618 & w2276) | (w1836 & w2276);
assign w2372 = (w618 & w1836) | (w618 & w2275) | (w1836 & w2275);
assign w2373 = w761 & w1608;
assign w2374 = ~w785 & ~w1608;
assign w2375 = ~w785 & w741;
assign w2376 = w778 & w785;
assign w2377 = w785 & w1608;
assign w2378 = w791 & ~w1622;
assign w2379 = w791 & ~w1623;
assign w2380 = w803 & w1608;
assign w2381 = w803 & w1609;
assign w2382 = ~w707 & w1591;
assign w2383 = ~w707 & w1075;
assign w2384 = ~w707 & ~w675;
assign w2385 = ~w719 & ~w1079;
assign w2386 = (w1074 & w2538) | (w1074 & w2539) | (w2538 & w2539);
assign w2387 = ~w737 & w1603;
assign w2388 = ~w737 & w1604;
assign w2389 = ~w712 & w1595;
assign w2390 = ~w1594 & ~w712;
assign w2391 = ~w675 & w1595;
assign w2392 = ~w1594 & w2540;
assign w2393 = (~w712 & ~w675) | (~w712 & w1595) | (~w675 & w1595);
assign w2394 = (~w712 & ~w1594) | (~w712 & w2540) | (~w1594 & w2540);
assign w2395 = ~w767 & ~w760;
assign w2396 = ~w767 & w1610;
assign w2397 = (w977 & w976) | (w977 & w958) | (w976 & w958);
assign w2398 = (w977 & w976) | (w977 & w957) | (w976 & w957);
assign w2399 = (w1042 & w1041) | (w1042 & ~w1020) | (w1041 & ~w1020);
assign w2400 = (w1042 & w1041) | (w1042 & ~w1019) | (w1041 & ~w1019);
assign w2401 = (w1204 & w1205) | (w1204 & ~w1020) | (w1205 & ~w1020);
assign w2402 = (w1204 & w1205) | (w1204 & ~w1019) | (w1205 & ~w1019);
assign w2403 = (w1206 & w1207) | (w1206 & ~w1020) | (w1207 & ~w1020);
assign w2404 = (w1206 & w1207) | (w1206 & ~w1019) | (w1207 & ~w1019);
assign w2405 = (w1209 & w1208) | (w1209 & ~w1020) | (w1208 & ~w1020);
assign w2406 = (w1209 & w1208) | (w1209 & ~w1019) | (w1208 & ~w1019);
assign w2407 = (w1211 & w1210) | (w1211 & ~w1020) | (w1210 & ~w1020);
assign w2408 = (w1211 & w1210) | (w1211 & ~w1019) | (w1210 & ~w1019);
assign w2409 = (w1213 & w1212) | (w1213 & ~w1020) | (w1212 & ~w1020);
assign w2410 = (w1213 & w1212) | (w1213 & ~w1019) | (w1212 & ~w1019);
assign w2411 = (w1215 & w1214) | (w1215 & ~w1020) | (w1214 & ~w1020);
assign w2412 = (w1215 & w1214) | (w1215 & ~w1019) | (w1214 & ~w1019);
assign w2413 = ~w1057 & w2541;
assign w2414 = (w1051 & w2726) | (w1051 & w2727) | (w2726 & w2727);
assign w2415 = (w664 & w1057) | (w664 & w2542) | (w1057 & w2542);
assign w2416 = w664 & w2974;
assign w2417 = ~w670 & w1060;
assign w2418 = ~w670 & w2900;
assign w2419 = w670 & ~w1060;
assign w2420 = (w1057 & w2543) | (w1057 & w2544) | (w2543 & w2544);
assign w2421 = ~w676 & w2901;
assign w2422 = (w1055 & w2545) | (w1055 & w2546) | (w2545 & w2546);
assign w2423 = (w1034 & w2547) | (w1034 & w2548) | (w2547 & w2548);
assign w2424 = (~w1055 & w2549) | (~w1055 & w2550) | (w2549 & w2550);
assign w2425 = ~w683 & w2901;
assign w2426 = ~w683 & w1066;
assign w2427 = (w1034 & w2551) | (w1034 & w2552) | (w2551 & w2552);
assign w2428 = w683 & ~w1066;
assign w2429 = ~w54 & ~w62;
assign w2430 = ~w62 & w1748;
assign w2431 = w54 & w62;
assign w2432 = w90 & ~w837;
assign w2433 = w90 & ~w838;
assign w2434 = w109 & ~w1754;
assign w2435 = w109 & ~w1753;
assign w2436 = (w858 & w2553) | (w858 & w2554) | (w2553 & w2554);
assign w2437 = ~w859 & w2553;
assign w2438 = w148 & ~w861;
assign w2439 = (w148 & w859) | (w148 & w2555) | (w859 & w2555);
assign w2440 = ~w160 & w1765;
assign w2441 = ~w160 & w1764;
assign w2442 = w160 & ~w1764;
assign w2443 = ~w172 & w870;
assign w2444 = ~w869 & w2556;
assign w2445 = w172 & ~w870;
assign w2446 = ~w178 & w872;
assign w2447 = (w870 & w2558) | (w870 & w2559) | (w2558 & w2559);
assign w2448 = w178 & ~w872;
assign w2449 = w178 & w2902;
assign w2450 = ~w277 & w1783;
assign w2451 = ~w277 & w1782;
assign w2452 = w277 & ~w1782;
assign w2453 = ~w353 & w1795;
assign w2454 = w353 & ~w1795;
assign w2455 = w353 & ~w1796;
assign w2456 = w359 & w2903;
assign w2457 = w359 & w2904;
assign w2458 = ~w377 & w2905;
assign w2459 = ~w950 & w2561;
assign w2460 = (w947 & w2562) | (w947 & w2563) | (w2562 & w2563);
assign w2461 = (w377 & w950) | (w377 & w2564) | (w950 & w2564);
assign w2462 = w383 & ~w952;
assign w2463 = ~w402 & w1801;
assign w2464 = (w1492 & w2567) | (w1492 & w2568) | (w2567 & w2568);
assign w2465 = w402 & ~w1801;
assign w2466 = w402 & w2907;
assign w2467 = w408 & ~w1803;
assign w2468 = w408 & ~w1802;
assign w2469 = w414 & ~w1805;
assign w2470 = w414 & ~w1804;
assign w2471 = ~w426 & w2908;
assign w2472 = (w964 & w2570) | (w964 & w2569) | (w2570 & w2569);
assign w2473 = w426 & ~w969;
assign w2474 = ~w432 & w971;
assign w2475 = ~w432 & w970;
assign w2476 = (w1365 & w1364) | (w1365 & ~w958) | (w1364 & ~w958);
assign w2477 = (w1365 & w1364) | (w1365 & ~w957) | (w1364 & ~w957);
assign w2478 = (w1367 & w1366) | (w1367 & w958) | (w1366 & w958);
assign w2479 = (w1367 & w1366) | (w1367 & w957) | (w1366 & w957);
assign w2480 = (w1369 & w1368) | (w1369 & w958) | (w1368 & w958);
assign w2481 = (w1369 & w1368) | (w1369 & w957) | (w1368 & w957);
assign w2482 = ~w508 & ~w500;
assign w2483 = ~w508 & w1812;
assign w2484 = ~w1528 & w2482;
assign w2485 = w508 & w500;
assign w2486 = (w1001 & w2573) | (w1001 & w2574) | (w2573 & w2574);
assign w2487 = (~w514 & w1001) | (~w514 & w2574) | (w1001 & w2574);
assign w2488 = w514 & w2909;
assign w2489 = ~w1001 & w2575;
assign w2490 = (w1004 & w2576) | (w1004 & w2577) | (w2576 & w2577);
assign w2491 = (~w520 & w1004) | (~w520 & w2577) | (w1004 & w2577);
assign w2492 = ~w526 & w1817;
assign w2493 = ~w526 & w1816;
assign w2494 = ~w1012 & w2580;
assign w2495 = (w1009 & w2581) | (w1009 & w2582) | (w2581 & w2582);
assign w2496 = (w544 & w1012) | (w544 & w2583) | (w1012 & w2583);
assign w2497 = w544 & ~w1013;
assign w2498 = ~w550 & w2910;
assign w2499 = (w1009 & w2585) | (w1009 & w2586) | (w2585 & w2586);
assign w2500 = (w1012 & w2587) | (w1012 & w2588) | (w2587 & w2588);
assign w2501 = (~w1009 & w2589) | (~w1009 & w2590) | (w2589 & w2590);
assign w2502 = ~w556 & ~w998;
assign w2503 = (~w1012 & w2591) | (~w1012 & w2592) | (w2591 & w2592);
assign w2504 = (w992 & w2593) | (w992 & w2594) | (w2593 & w2594);
assign w2505 = (w1012 & w2595) | (w1012 & w2596) | (w2595 & w2596);
assign w2506 = w563 & ~w2370;
assign w2507 = w563 & ~w2369;
assign w2508 = (w1026 & w2597) | (w1026 & w2598) | (w2597 & w2598);
assign w2509 = (w1026 & w2599) | (w1026 & w2598) | (w2599 & w2598);
assign w2510 = w575 & w2912;
assign w2511 = ~w581 & w1830;
assign w2512 = ~w581 & w1829;
assign w2513 = w581 & ~w1829;
assign w2514 = ~w1034 & w2601;
assign w2515 = (w1031 & w2602) | (w1031 & w2603) | (w2602 & w2603);
assign w2516 = (w599 & w1034) | (w599 & w2604) | (w1034 & w2604);
assign w2517 = w599 & ~w1035;
assign w2518 = ~w605 & w2913;
assign w2519 = (w1031 & w2606) | (w1031 & w2607) | (w2606 & w2607);
assign w2520 = (w1034 & w2608) | (w1034 & w2609) | (w2608 & w2609);
assign w2521 = (~w1031 & w2610) | (~w1031 & w2611) | (w2610 & w2611);
assign w2522 = ~w611 & w2851;
assign w2523 = (~w1034 & w2612) | (~w1034 & w2613) | (w2612 & w2613);
assign w2524 = (w1012 & w2614) | (w1012 & w2615) | (w2614 & w2615);
assign w2525 = (w1034 & w2616) | (w1034 & w2617) | (w2616 & w2617);
assign w2526 = (w1403 & w1404) | (w1403 & w1020) | (w1404 & w1020);
assign w2527 = (w1403 & w1404) | (w1403 & w1019) | (w1404 & w1019);
assign w2528 = (~w801 & w1631) | (~w801 & ~w795) | (w1631 & ~w795);
assign w2529 = (~w801 & w1631) | (~w801 & w1627) | (w1631 & w1627);
assign w2530 = ~w778 & ~w785;
assign w2531 = ~w1620 & w2618;
assign w2532 = (w1619 & w2618) | (w1619 & w2533) | (w2618 & w2533);
assign w2533 = ~w791 & w1622;
assign w2534 = w803 & ~w2312;
assign w2535 = w803 & ~w2311;
assign w2536 = ~w718 & ~w725;
assign w2537 = w718 & w725;
assign w2538 = w719 & w1924;
assign w2539 = w719 & w1923;
assign w2540 = ~w712 & ~w675;
assign w2541 = ~w657 & ~w664;
assign w2542 = w657 & w664;
assign w2543 = w670 & ~w1858;
assign w2544 = w670 & ~w1583;
assign w2545 = ~w1585 & w2619;
assign w2546 = (w1584 & w2619) | (w1584 & w2620) | (w2619 & w2620);
assign w2547 = w676 & ~w2278;
assign w2548 = w676 & ~w2277;
assign w2549 = (w676 & w1585) | (w676 & w2621) | (w1585 & w2621);
assign w2550 = w676 & ~w2286;
assign w2551 = w683 & ~w2278;
assign w2552 = w683 & ~w2277;
assign w2553 = ~w148 & ~w141;
assign w2554 = ~w148 & w1417;
assign w2555 = w148 & w141;
assign w2556 = ~w165 & ~w172;
assign w2557 = w165 & w172;
assign w2558 = ~w178 & ~w171;
assign w2559 = ~w178 & w1425;
assign w2560 = ~w359 & w942;
assign w2561 = ~w370 & ~w377;
assign w2562 = w377 & ~w1480;
assign w2563 = w377 & ~w1481;
assign w2564 = w370 & w377;
assign w2565 = w383 & ~w2240;
assign w2566 = w383 & ~w2239;
assign w2567 = ~w402 & ~w395;
assign w2568 = ~w402 & w959;
assign w2569 = ~w426 & w1499;
assign w2570 = ~w426 & w1500;
assign w2571 = w426 & ~w1845;
assign w2572 = w426 & ~w1499;
assign w2573 = ~w514 & w499;
assign w2574 = ~w514 & w1000;
assign w2575 = w514 & ~w1000;
assign w2576 = ~w520 & w499;
assign w2577 = ~w520 & w1003;
assign w2578 = w520 & ~w499;
assign w2579 = w520 & ~w1003;
assign w2580 = ~w537 & ~w544;
assign w2581 = ~w544 & w1539;
assign w2582 = ~w544 & w1538;
assign w2583 = w537 & w544;
assign w2584 = ~w550 & w1542;
assign w2585 = ~w1540 & w2728;
assign w2586 = (w1539 & w2728) | (w1539 & w2584) | (w2728 & w2584);
assign w2587 = w550 & ~w1542;
assign w2588 = w550 & ~w1543;
assign w2589 = (w550 & w1540) | (w550 & w2729) | (w1540 & w2729);
assign w2590 = w550 & ~w2261;
assign w2591 = ~w556 & w2264;
assign w2592 = ~w1545 & w2730;
assign w2593 = w556 & w1528;
assign w2594 = w556 & w1527;
assign w2595 = w556 & ~w2264;
assign w2596 = (w556 & w1545) | (w556 & w2731) | (w1545 & w2731);
assign w2597 = ~w575 & ~w1548;
assign w2598 = ~w575 & w1025;
assign w2599 = ~w575 & ~w1547;
assign w2600 = w575 & ~w1025;
assign w2601 = ~w592 & ~w599;
assign w2602 = ~w599 & w1560;
assign w2603 = ~w599 & w1559;
assign w2604 = w592 & w599;
assign w2605 = ~w605 & w1563;
assign w2606 = ~w1561 & w2732;
assign w2607 = (w1560 & w2732) | (w1560 & w2605) | (w2732 & w2605);
assign w2608 = w605 & ~w1563;
assign w2609 = w605 & ~w1564;
assign w2610 = (w605 & w1561) | (w605 & w2733) | (w1561 & w2733);
assign w2611 = w605 & ~w2271;
assign w2612 = ~w611 & w2274;
assign w2613 = ~w1566 & w2734;
assign w2614 = (w1544 & w2735) | (w1544 & w2736) | (w2735 & w2736);
assign w2615 = (w1545 & w2735) | (w1545 & w2736) | (w2735 & w2736);
assign w2616 = w611 & ~w2274;
assign w2617 = (w611 & w1566) | (w611 & w2737) | (w1566 & w2737);
assign w2618 = ~w784 & ~w791;
assign w2619 = ~w669 & ~w676;
assign w2620 = ~w676 & w1587;
assign w2621 = w669 & w676;
assign w2622 = (w1894 & w1893) | (w1894 & ~w1892) | (w1893 & ~w1892);
assign w2623 = (w1894 & w1893) | (w1894 & ~w1891) | (w1893 & ~w1891);
assign w2624 = (w1198 & w1197) | (w1198 & ~w1219) | (w1197 & ~w1219);
assign w2625 = (w1198 & w1197) | (w1198 & ~w1220) | (w1197 & ~w1220);
assign w2626 = (~w499 & w1524) | (~w499 & w1849) | (w1524 & w1849);
assign w2627 = ~w499 & ~w1919;
assign w2628 = ~w190 & w2036;
assign w2629 = ~w190 & w2035;
assign w2630 = w308 & w2914;
assign w2631 = w308 & w2915;
assign w2632 = w314 & ~w2076;
assign w2633 = w314 & ~w2075;
assign w2634 = w320 & ~w2078;
assign w2635 = w320 & ~w2077;
assign w2636 = w326 & ~w2080;
assign w2637 = w326 & ~w2079;
assign w2638 = w339 & ~w2084;
assign w2639 = w339 & ~w2083;
assign w2640 = (w2091 & w2092) | (w2091 & w2074) | (w2092 & w2074);
assign w2641 = (w2091 & w2092) | (w2091 & w2073) | (w2092 & w2073);
assign w2642 = (w2095 & w2096) | (w2095 & w2074) | (w2096 & w2074);
assign w2643 = (w2095 & w2096) | (w2095 & w2073) | (w2096 & w2073);
assign w2644 = w365 & w2916;
assign w2645 = w365 & w2917;
assign w2646 = w371 & w2975;
assign w2647 = w371 & w2976;
assign w2648 = (w1946 & w1945) | (w1946 & ~w1902) | (w1945 & ~w1902);
assign w2649 = (w1946 & w1945) | (w1946 & ~w1901) | (w1945 & ~w1901);
assign w2650 = (w1950 & w1949) | (w1950 & ~w1902) | (w1949 & ~w1902);
assign w2651 = (w1950 & w1949) | (w1950 & ~w1901) | (w1949 & ~w1901);
assign w2652 = (w1505 & w1504) | (w1505 & w1500) | (w1504 & w1500);
assign w2653 = (w1505 & w1504) | (w1505 & w1499) | (w1504 & w1499);
assign w2654 = (w1523 & w1522) | (w1523 & w1518) | (w1522 & w1518);
assign w2655 = (w1523 & w1522) | (w1523 & w1517) | (w1522 & w1517);
assign w2656 = (~w549 & w1546) | (~w549 & w2262) | (w1546 & w2262);
assign w2657 = (w1539 & w2740) | (w1539 & w2264) | (w2740 & w2264);
assign w2658 = ~w554 & ~w2656;
assign w2659 = ~w554 & w2918;
assign w2660 = (~w604 & w1567) | (~w604 & w2272) | (w1567 & w2272);
assign w2661 = (w1560 & w2741) | (w1560 & w2274) | (w2741 & w2274);
assign w2662 = (w1570 & w1569) | (w1570 & w2272) | (w1569 & w2272);
assign w2663 = (w1570 & w1569) | (w1570 & w2271) | (w1569 & w2271);
assign w2664 = (~w657 & w1581) | (~w657 & w1579) | (w1581 & w1579);
assign w2665 = (~w657 & w1581) | (~w657 & w1578) | (w1581 & w1578);
assign w2666 = (~w675 & w1591) | (~w675 & w2287) | (w1591 & w2287);
assign w2667 = (w1584 & w2742) | (w1584 & w2743) | (w2742 & w2743);
assign w2668 = (~w736 & w1607) | (~w736 & w2300) | (w1607 & w2300);
assign w2669 = (w1600 & w2744) | (w1600 & w2745) | (w2744 & w2745);
assign w2670 = ~w741 & ~w2668;
assign w2671 = ~w741 & w2919;
assign w2672 = (~w790 & w1626) | (~w790 & w2308) | (w1626 & w2308);
assign w2673 = (w1619 & w2746) | (w1619 & w2310) | (w2746 & w2310);
assign w2674 = (w1629 & w1628) | (w1629 & w2308) | (w1628 & w2308);
assign w2675 = (w1629 & w1628) | (w1629 & w2307) | (w1628 & w2307);
assign w2676 = ~w749 & w2920;
assign w2677 = ~w749 & w2921;
assign w2678 = (~w617 & w1043) | (~w617 & w2662) | (w1043 & w2662);
assign w2679 = (~w617 & w1043) | (~w617 & w2663) | (w1043 & w2663);
assign w2680 = (w1046 & w1045) | (w1046 & w2662) | (w1045 & w2662);
assign w2681 = (w1046 & w1045) | (w1046 & w2663) | (w1045 & w2663);
assign w2682 = ~w689 & w2977;
assign w2683 = ~w689 & w2978;
assign w2684 = (w1788 & w1787) | (w1788 & w1455) | (w1787 & w1455);
assign w2685 = (w1788 & w1787) | (w1788 & w1454) | (w1787 & w1454);
assign w2686 = (w1826 & w1825) | (w1826 & w2262) | (w1825 & w2262);
assign w2687 = (w1826 & w1825) | (w1826 & w2261) | (w1825 & w2261);
assign w2688 = ~w562 & w2922;
assign w2689 = ~w562 & w2923;
assign w2690 = ~w618 & w2662;
assign w2691 = ~w618 & w2663;
assign w2692 = w785 & ~w741;
assign w2693 = (w791 & w1620) | (w791 & w2747) | (w1620 & w2747);
assign w2694 = w791 & ~w2307;
assign w2695 = ~w803 & w2924;
assign w2696 = ~w803 & w2925;
assign w2697 = ~w803 & w2674;
assign w2698 = ~w803 & w2675;
assign w2699 = ~w1601 & w2748;
assign w2700 = (w1600 & w2748) | (w1600 & w2387) | (w2748 & w2387);
assign w2701 = ~w737 & w2666;
assign w2702 = ~w737 & w2926;
assign w2703 = ~w115 & w848;
assign w2704 = ~w115 & w847;
assign w2705 = ~w154 & w853;
assign w2706 = ~w154 & w863;
assign w2707 = w160 & ~w1763;
assign w2708 = (w172 & w869) | (w172 & w2557) | (w869 & w2557);
assign w2709 = w178 & w2902;
assign w2710 = w277 & ~w1781;
assign w2711 = ~w1472 & w2749;
assign w2712 = (w1471 & w2749) | (w1471 & w2453) | (w2749 & w2453);
assign w2713 = (w353 & w1472) | (w353 & w2750) | (w1472 & w2750);
assign w2714 = w353 & w2927;
assign w2715 = (w950 & w2565) | (w950 & w2566) | (w2565 & w2566);
assign w2716 = (w966 & w2571) | (w966 & w2572) | (w2571 & w2572);
assign w2717 = w426 & ~w969;
assign w2718 = ~w508 & w2979;
assign w2719 = ~w508 & w2928;
assign w2720 = w508 & ~w1812;
assign w2721 = (w508 & w1528) | (w508 & w2485) | (w1528 & w2485);
assign w2722 = w514 & ~w1815;
assign w2723 = w514 & ~w1814;
assign w2724 = w575 & w2929;
assign w2725 = w581 & ~w1828;
assign w2726 = ~w664 & w2664;
assign w2727 = ~w664 & w2665;
assign w2728 = ~w543 & ~w550;
assign w2729 = w543 & w550;
assign w2730 = ~w549 & ~w556;
assign w2731 = w549 & w556;
assign w2732 = ~w598 & ~w605;
assign w2733 = w598 & w605;
assign w2734 = ~w604 & ~w611;
assign w2735 = w611 & ~w554;
assign w2736 = w611 & w1547;
assign w2737 = w604 & w611;
assign w2738 = ~w308 & w1334;
assign w2739 = ~w308 & w1333;
assign w2740 = (~w549 & w1546) | (~w549 & ~w543) | (w1546 & ~w543);
assign w2741 = (~w604 & w1567) | (~w604 & ~w598) | (w1567 & ~w598);
assign w2742 = (~w675 & w1591) | (~w675 & ~w669) | (w1591 & ~w669);
assign w2743 = (~w675 & w1591) | (~w675 & w1587) | (w1591 & w1587);
assign w2744 = (~w736 & w1607) | (~w736 & ~w730) | (w1607 & ~w730);
assign w2745 = (~w736 & w1607) | (~w736 & w1603) | (w1607 & w1603);
assign w2746 = (~w790 & w1626) | (~w790 & ~w784) | (w1626 & ~w784);
assign w2747 = w784 & w791;
assign w2748 = ~w730 & ~w737;
assign w2749 = ~w345 & ~w353;
assign w2750 = w345 & w353;
assign w2751 = (w2462 & w2715) | (w2462 & w2088) | (w2715 & w2088);
assign w2752 = (w2462 & w2715) | (w2462 & w2087) | (w2715 & w2087);
assign w2753 = ~w624 & w1934;
assign w2754 = ~w624 & w1933;
assign w2755 = ~w630 & w1936;
assign w2756 = ~w630 & w1935;
assign w2757 = (w1954 & w1953) | (w1954 & ~w1902) | (w1953 & ~w1902);
assign w2758 = (w1954 & w1953) | (w1954 & ~w1901) | (w1953 & ~w1901);
assign w2759 = (w1219 & w1220) | (w1219 & ~w1902) | (w1220 & ~w1902);
assign w2760 = (w1219 & w1220) | (w1219 & ~w1901) | (w1220 & ~w1901);
assign w2761 = (w1222 & w1221) | (w1222 & w1932) | (w1221 & w1932);
assign w2762 = (w1222 & w1221) | (w1222 & w1931) | (w1221 & w1931);
assign w2763 = (w1226 & w1225) | (w1226 & w1932) | (w1225 & w1932);
assign w2764 = (w1226 & w1225) | (w1226 & w1931) | (w1225 & w1931);
assign w2765 = (w1230 & w1229) | (w1230 & w1932) | (w1229 & w1932);
assign w2766 = (w1230 & w1229) | (w1230 & w1931) | (w1229 & w1931);
assign w2767 = (w1234 & w1233) | (w1234 & w1932) | (w1233 & w1932);
assign w2768 = (w1234 & w1233) | (w1234 & w1931) | (w1233 & w1931);
assign w2769 = (w1238 & w1237) | (w1238 & w1932) | (w1237 & w1932);
assign w2770 = (w1238 & w1237) | (w1238 & w1931) | (w1237 & w1931);
assign w2771 = (w1242 & w1241) | (w1242 & w1932) | (w1241 & w1932);
assign w2772 = (w1242 & w1241) | (w1242 & w1931) | (w1241 & w1931);
assign w2773 = (w1250 & w1249) | (w1250 & w1932) | (w1249 & w1932);
assign w2774 = (w1250 & w1249) | (w1250 & w1931) | (w1249 & w1931);
assign w2775 = (w1254 & w1253) | (w1254 & w1932) | (w1253 & w1932);
assign w2776 = (w1254 & w1253) | (w1254 & w1931) | (w1253 & w1931);
assign w2777 = (w809 & w1637) | (w809 & w2314) | (w1637 & w2314);
assign w2778 = (w809 & w1637) | (w809 & w2313) | (w1637 & w2313);
assign w2779 = (~w807 & w1869) | (~w807 & w2314) | (w1869 & w2314);
assign w2780 = (~w807 & w1869) | (~w807 & w2313) | (w1869 & w2313);
assign w2781 = (w737 & w1601) | (w737 & w2785) | (w1601 & w2785);
assign w2782 = w737 & ~w2299;
assign w2783 = (w2487 & w2486) | (w2487 & w1920) | (w2486 & w1920);
assign w2784 = (w2487 & w2486) | (w2487 & w1919) | (w2486 & w1919);
assign w2785 = w730 & w737;
assign w2786 = (w27 & ~w819) | (w27 & ~w25) | (~w819 & ~w25);
assign w2787 = (~w834 & ~w835) | (~w834 & ~w59) | (~w835 & ~w59);
assign w2788 = (w841 & w840) | (w841 & w2787) | (w840 & w2787);
assign w2789 = (w851 & w850) | (w851 & w100) | (w850 & w100);
assign w2790 = (~w1298 & ~w1297) | (~w1298 & ~w125) | (~w1297 & ~w125);
assign w2791 = (~w1300 & ~w1299) | (~w1300 & ~w125) | (~w1299 & ~w125);
assign w2792 = (w866 & w865) | (w866 & ~w125) | (w865 & ~w125);
assign w2793 = (~w2036 & ~w2035) | (~w2036 & ~w125) | (~w2035 & ~w125);
assign w2794 = (w876 & w875) | (w876 & w2792) | (w875 & w2792);
assign w2795 = (w1316 & w1315) | (w1316 & ~w2794) | (w1315 & ~w2794);
assign w2796 = (w1318 & w1317) | (w1318 & ~w2794) | (w1317 & ~w2794);
assign w2797 = (~w1324 & ~w1323) | (~w1324 & ~w222) | (~w1323 & ~w222);
assign w2798 = (~w1326 & ~w1325) | (~w1326 & ~w222) | (~w1325 & ~w222);
assign w2799 = (~w1328 & ~w1327) | (~w1328 & ~w222) | (~w1327 & ~w222);
assign w2800 = (~w1330 & ~w1329) | (~w1330 & ~w222) | (~w1329 & ~w222);
assign w2801 = (~w1332 & ~w1331) | (~w1332 & ~w222) | (~w1331 & ~w222);
assign w2802 = (w1893 & w1894) | (w1893 & ~w2794) | (w1894 & ~w2794);
assign w2803 = (w2076 & w2075) | (w2076 & ~w2794) | (w2075 & ~w2794);
assign w2804 = (w2078 & w2077) | (w2078 & ~w2794) | (w2077 & ~w2794);
assign w2805 = (w2080 & w2079) | (w2080 & ~w2794) | (w2079 & ~w2794);
assign w2806 = (w2084 & w2083) | (w2084 & ~w2794) | (w2083 & ~w2794);
assign w2807 = (w939 & w940) | (w939 & w2930) | (w940 & w2930);
assign w2808 = (~w1385 & ~w1384) | (~w1385 & ~w442) | (~w1384 & ~w442);
assign w2809 = (~w1387 & ~w1386) | (~w1387 & ~w442) | (~w1386 & ~w442);
assign w2810 = (w1899 & w1900) | (w1899 & ~w393) | (w1900 & ~w393);
assign w2811 = (~w1934 & ~w1933) | (~w1934 & ~w393) | (~w1933 & ~w393);
assign w2812 = (~w1936 & ~w1935) | (~w1936 & ~w393) | (~w1935 & ~w393);
assign w2813 = (w176 & ~w1426) | (w176 & ~w871) | (~w1426 & ~w871);
assign w2814 = (w209 & ~w1434) | (w209 & ~w882) | (~w1434 & ~w882);
assign w2815 = (w250 & ~w1445) | (w250 & ~w897) | (~w1445 & ~w897);
assign w2816 = (w287 & ~w1453) | (w287 & ~w912) | (~w1453 & ~w912);
assign w2817 = (w324 & ~w1463) | (w324 & ~w928) | (~w1463 & ~w928);
assign w2818 = (w369 & ~w1478) | (w369 & ~w947) | (~w1478 & ~w947);
assign w2819 = (w471 & ~w1516) | (w471 & ~w985) | (~w1516 & ~w985);
assign w2820 = (w492 & ~w1525) | (w492 & ~w992) | (~w1525 & ~w992);
assign w2821 = (w524 & ~w1532) | (w524 & ~w1005) | (~w1532 & ~w1005);
assign w2822 = (w542 & ~w1541) | (w542 & ~w1012) | (~w1541 & ~w1012);
assign w2823 = (w579 & ~w1552) | (w579 & ~w1027) | (~w1552 & ~w1027);
assign w2824 = (w597 & ~w1562) | (w597 & ~w1034) | (~w1562 & ~w1034);
assign w2825 = (~w1565 & ~w1566) | (~w1565 & ~w1034) | (~w1566 & ~w1034);
assign w2826 = (w662 & ~w1582) | (w662 & ~w1057) | (~w1582 & ~w1057);
assign w2827 = (w699 & ~w1201) | (w699 & ~w1071) | (~w1201 & ~w1071);
assign w2828 = (w723 & ~w1598) | (w723 & ~w1082) | (~w1598 & ~w1082);
assign w2829 = (w765 & ~w1611) | (w765 & ~w1099) | (~w1611 & ~w1099);
assign w2830 = (~w1624 & ~w1625) | (~w1624 & ~w1107) | (~w1625 & ~w1107);
assign w2831 = (~w2314 & ~w2313) | (~w2314 & ~w1107) | (~w2313 & ~w1107);
assign w2832 = (w741 & ~w1608) | (w741 & ~w1088) | (~w1608 & ~w1088);
assign w2833 = (w1881 & w1882) | (w1881 & ~w1088) | (w1882 & ~w1088);
assign w2834 = (w1883 & w2373) | (w1883 & ~w1086) | (w2373 & ~w1086);
assign w2835 = (w1645 & w1644) | (w1645 & ~w1088) | (w1644 & ~w1088);
assign w2836 = (~w1646 & ~w1645) | (~w1646 & ~w1086) | (~w1645 & ~w1086);
assign w2837 = (~w1658 & ~w1657) | (~w1658 & ~w1062) | (~w1657 & ~w1062);
assign w2838 = (w1073 & w1072) | (w1073 & w1066) | (w1072 & w1066);
assign w2839 = (~w1661 & ~w1660) | (~w1661 & ~w1062) | (~w1660 & ~w1062);
assign w2840 = w2384 & ~w1064;
assign w2841 = (w60 & ~w829) | (w60 & ~w828) | (~w829 & ~w828);
assign w2842 = (w60 & ~w829) | (w60 & ~w827) | (~w829 & ~w827);
assign w2843 = (w2813 & ~w873) | (w2813 & ~w866) | (~w873 & ~w866);
assign w2844 = (w2813 & ~w873) | (w2813 & ~w865) | (~w873 & ~w865);
assign w2845 = ~w217 & ~w887;
assign w2846 = ~w257 & ~w902;
assign w2847 = (w299 & ~w1458) | (w299 & ~w917) | (~w1458 & ~w917);
assign w2848 = (w2817 & ~w931) | (w2817 & ~w920) | (~w931 & ~w920);
assign w2849 = ~w388 & ~w956;
assign w2850 = ~w437 & ~w975;
assign w2851 = (w554 & ~w1547) | (w554 & ~w1016) | (~w1547 & ~w1016);
assign w2852 = (w802 & ~w1867) | (w802 & ~w1628) | (~w1867 & ~w1628);
assign w2853 = (w747 & ~w1093) | (w747 & w741) | (~w1093 & w741);
assign w2854 = (w747 & ~w1093) | (w747 & ~w1608) | (~w1093 & ~w1608);
assign w2855 = (w747 & ~w1093) | (w747 & ~w1609) | (~w1093 & ~w1609);
assign w2856 = (w1608 & ~w1094) | (w1608 & ~w1095) | (~w1094 & ~w1095);
assign w2857 = (w1608 & ~w1097) | (w1608 & ~w1098) | (~w1097 & ~w1098);
assign w2858 = ~w796 & w2932;
assign w2859 = (w158 & ~w867) | (w158 & ~w1421) | (~w867 & ~w1421);
assign w2860 = (w158 & ~w867) | (w158 & ~w1422) | (~w867 & ~w1422);
assign w2861 = ~w877 | w188;
assign w2862 = (w188 & ~w877) | (w188 & w182) | (~w877 & w182);
assign w2863 = (w306 & ~w922) | (w306 & ~w1458) | (~w922 & ~w1458);
assign w2864 = (w306 & ~w922) | (w306 & ~w1459) | (~w922 & ~w1459);
assign w2865 = (w506 & ~w999) | (w506 & ~w1527) | (~w999 & ~w1527);
assign w2866 = (w506 & ~w999) | (w506 & ~w1528) | (~w999 & ~w1528);
assign w2867 = ~w1008 | w2821;
assign w2868 = (w2821 & ~w1008) | (w2821 & w499) | (~w1008 & w499);
assign w2869 = (w561 & ~w1021) | (w561 & ~w1548) | (~w1021 & ~w1548);
assign w2870 = (w2823 & ~w1030) | (w2823 & ~w1547) | (~w1030 & ~w1547);
assign w2871 = (w2823 & ~w1030) | (w2823 & ~w1548) | (~w1030 & ~w1548);
assign w2872 = (w54 & ~w1748) | (w54 & ~w826) | (~w1748 & ~w826);
assign w2873 = (~w102 & w845) | (~w102 & w844) | (w845 & w844);
assign w2874 = (~w848 & ~w847) | (~w848 & ~w843) | (~w847 & ~w843);
assign w2875 = (~w853 & ~w863) | (~w853 & ~w864) | (~w863 & ~w864);
assign w2876 = ~w153 & ~w866;
assign w2877 = (~w1765 & ~w1764) | (~w1765 & ~w860) | (~w1764 & ~w860);
assign w2878 = (w908 & w907) | (w908 & w2846) | (w907 & w2846);
assign w2879 = (~w1783 & ~w1782) | (~w1783 & ~w900) | (~w1782 & ~w900);
assign w2880 = ~w345 & ~w940;
assign w2881 = ~w359 & ~w940;
assign w2882 = (w962 & w961) | (w962 & w958) | (w961 & w958);
assign w2883 = (w965 & w964) | (w965 & w2849) | (w964 & w2849);
assign w2884 = (~w971 & ~w970) | (~w971 & ~w957) | (~w970 & ~w957);
assign w2885 = (~w971 & ~w970) | (~w971 & ~w958) | (~w970 & ~w958);
assign w2886 = ~w507 & w2933;
assign w2887 = w2578 & ~w995;
assign w2888 = (~w1817 & ~w1816) | (~w1817 & ~w995) | (~w1816 & ~w995);
assign w2889 = ~w555 & ~w1020;
assign w2890 = ~w575 & w2851;
assign w2891 = w575 & w2980;
assign w2892 = (w1028 & w1029) | (w1028 & w2851) | (w1029 & w2851);
assign w2893 = (~w1830 & ~w1829) | (~w1830 & ~w1015) | (~w1829 & ~w1015);
assign w2894 = (w795 & ~w1627) | (w795 & ~w1624) | (~w1627 & ~w1624);
assign w2895 = (w795 & ~w1627) | (w795 & ~w1625) | (~w1627 & ~w1625);
assign w2896 = (~w741 & ~w1097) | (~w741 & ~w1098) | (~w1097 & ~w1098);
assign w2897 = (w351 & ~w941) | (w351 & ~w1472) | (~w941 & ~w1472);
assign w2898 = ~w388 & ~w1489;
assign w2899 = ~w437 & ~w1507;
assign w2900 = ~w663 & w2826;
assign w2901 = ~w610 & ~w1040;
assign w2902 = (w171 & ~w1425) | (w171 & ~w870) | (~w1425 & ~w870);
assign w2903 = (w1474 & ~w942) | (w1474 & ~w943) | (~w942 & ~w943);
assign w2904 = (~w344 & ~w942) | (~w344 & ~w943) | (~w942 & ~w943);
assign w2905 = ~w370 & w2818;
assign w2906 = (~w376 & w1484) | (~w376 & w951) | (w1484 & w951);
assign w2907 = (w395 & ~w959) | (w395 & ~w1492) | (~w959 & ~w1492);
assign w2908 = ~w419 & w2934;
assign w2909 = (~w499 & ~w1000) | (~w499 & ~w1001) | (~w1000 & ~w1001);
assign w2910 = ~w543 & w2822;
assign w2911 = (w1547 & ~w1022) | (w1547 & ~w1023) | (~w1022 & ~w1023);
assign w2912 = (w1547 & ~w1025) | (w1547 & ~w1026) | (~w1025 & ~w1026);
assign w2913 = ~w598 & w2824;
assign w2914 = (~w1334 & ~w1333) | (~w1334 & ~w1893) | (~w1333 & ~w1893);
assign w2915 = (~w1334 & ~w1333) | (~w1334 & ~w1894) | (~w1333 & ~w1894);
assign w2916 = (~w1345 & ~w1344) | (~w1345 & w2074) | (~w1344 & w2074);
assign w2917 = (~w1345 & ~w1344) | (~w1345 & w2073) | (~w1344 & w2073);
assign w2918 = (w549 & ~w1546) | (w549 & ~w2261) | (~w1546 & ~w2261);
assign w2919 = (w736 & ~w1607) | (w736 & ~w2299) | (~w1607 & ~w2299);
assign w2920 = (w1640 & w1639) | (w1640 & w2300) | (w1639 & w2300);
assign w2921 = (w1640 & w1639) | (w1640 & w2299) | (w1639 & w2299);
assign w2922 = (w561 & ~w1021) | (w561 & w2935) | (~w1021 & w2935);
assign w2923 = (w561 & ~w1021) | (w561 & w2936) | (~w1021 & w2936);
assign w2924 = (~w1608 & ~w1609) | (~w1608 & w2300) | (~w1609 & w2300);
assign w2925 = (~w1608 & ~w1609) | (~w1608 & w2299) | (~w1609 & w2299);
assign w2926 = (w1591 & ~w675) | (w1591 & w2286) | (~w675 & w2286);
assign w2927 = (w345 & ~w1795) | (w345 & ~w1471) | (~w1795 & ~w1471);
assign w2928 = (w1813 & ~w500) | (w1813 & w1919) | (~w500 & w1919);
assign w2929 = (~w554 & ~w1025) | (~w554 & ~w1026) | (~w1025 & ~w1026);
assign w2930 = (w920 & w921) | (w920 & ~w262) | (w921 & ~w262);
assign w2931 = (~w1591 & w675) | (~w1591 & ~w1062) | (w675 & ~w1062);
assign w2932 = (w2895 & w2894) | (w2895 & ~w1107) | (w2894 & ~w1107);
assign w2933 = (w506 & ~w999) | (w506 & ~w998) | (~w999 & ~w998);
assign w2934 = (w418 & ~w1498) | (w418 & ~w966) | (~w1498 & ~w966);
assign w2935 = (~w1548 & ~w1547) | (~w1548 & w2262) | (~w1547 & w2262);
assign w2936 = (~w1548 & ~w1547) | (~w1548 & w2261) | (~w1547 & w2261);
assign w2937 = ~w83 & w2981;
assign w2938 = (w1283 & w2873) | (w1283 & ~w80) | (w2873 & ~w80);
assign w2939 = (w2875 & ~w1296) | (w2875 & ~w100) | (~w1296 & ~w100);
assign w2940 = (w2888 & ~w1383) | (w2888 & ~w442) | (~w1383 & ~w442);
assign w2941 = (~w1916 & ~w1915) | (~w1916 & ~w966) | (~w1915 & ~w966);
assign w2942 = (~w1918 & ~w1917) | (~w1918 & ~w985) | (~w1917 & ~w985);
assign w2943 = (w795 & ~w1627) | (w795 & w2830) | (~w1627 & w2830);
assign w2944 = (w802 & ~w1867) | (w802 & w2963) | (~w1867 & w2963);
assign w2945 = (w2827 & ~w1074) | (w2827 & w1066) | (~w1074 & w1066);
assign w2946 = (~w1640 & ~w1639) | (~w1640 & ~w1086) | (~w1639 & ~w1086);
assign w2947 = (w1878 & w1876) | (w1878 & ~w1088) | (w1876 & ~w1088);
assign w2948 = (~w1643 & w2856) | (~w1643 & ~w1086) | (w2856 & ~w1086);
assign w2949 = (~w682 & w1067) | (~w682 & w1066) | (w1067 & w1066);
assign w2950 = (~w1655 & ~w1656) | (~w1655 & ~w1062) | (~w1656 & ~w1062);
assign w2951 = (~w1075 & w2931) | (~w1075 & ~w1076) | (w2931 & ~w1076);
assign w2952 = (~w1080 & ~w1081) | (~w1080 & ~w1065) | (~w1081 & ~w1065);
assign w2953 = (~w1084 & ~w1065) | (~w1084 & ~w1085) | (~w1065 & ~w1085);
assign w2954 = (w158 & ~w867) | (w158 & ~w866) | (~w867 & ~w866);
assign w2955 = (w188 & ~w877) | (w188 & ~w876) | (~w877 & ~w876);
assign w2956 = (w1439 & ~w217) | (w1439 & w886) | (~w217 & w886);
assign w2957 = (~w1449 & w257) | (~w1449 & ~w900) | (w257 & ~w900);
assign w2958 = (w2818 & ~w950) | (w2818 & ~w940) | (~w950 & ~w940);
assign w2959 = (w2821 & ~w1008) | (w2821 & ~w998) | (~w1008 & ~w998);
assign w2960 = (w561 & ~w1021) | (w561 & w2851) | (~w1021 & w2851);
assign w2961 = (w2823 & ~w1030) | (w2823 & w2851) | (~w1030 & w2851);
assign w2962 = (~w1570 & ~w1569) | (~w1570 & ~w1037) | (~w1569 & ~w1037);
assign w2963 = (~w1628 & ~w1629) | (~w1628 & ~w1110) | (~w1629 & ~w1110);
assign w2964 = (w2814 & ~w885) | (w2814 & ~w1891) | (~w885 & ~w1891);
assign w2965 = (w2814 & ~w885) | (w2814 & ~w1892) | (~w885 & ~w1892);
assign w2966 = (w2956 & w2845) | (w2956 & ~w1892) | (w2845 & ~w1892);
assign w2967 = (w2956 & w2845) | (w2956 & ~w1891) | (w2845 & ~w1891);
assign w2968 = (w952 & w2906) | (w952 & ~w939) | (w2906 & ~w939);
assign w2969 = (w952 & w2906) | (w952 & ~w940) | (w2906 & ~w940);
assign w2970 = (~w1813 & w500) | (~w1813 & ~w995) | (w500 & ~w995);
assign w2971 = (~w1825 & ~w1826) | (~w1825 & ~w1015) | (~w1826 & ~w1015);
assign w2972 = (~w1827 & w2911) | (~w1827 & ~w1015) | (w2911 & ~w1015);
assign w2973 = (w351 & ~w941) | (w351 & ~w1473) | (~w941 & ~w1473);
assign w2974 = (~w1581 & w657) | (~w1581 & ~w1055) | (w657 & ~w1055);
assign w2975 = (~w1346 & ~w1347) | (~w1346 & w2074) | (~w1347 & w2074);
assign w2976 = (~w1346 & ~w1347) | (~w1346 & w2073) | (~w1347 & w2073);
assign w2977 = (~w682 & w1067) | (~w682 & w2666) | (w1067 & w2666);
assign w2978 = (~w682 & w1067) | (~w682 & w2926) | (w1067 & w2926);
assign w2979 = (w1813 & ~w500) | (w1813 & w1920) | (~w500 & w1920);
assign w2980 = (w1548 & w1547) | (w1548 & ~w1015) | (w1547 & ~w1015);
assign w2981 = (w82 & ~w836) | (w82 & w2787) | (~w836 & w2787);
assign one = 1;
assign f_0 = ~w2;// level 2
assign f_1 = ~w9;// level 4
assign f_2 = w17;// level 5
assign f_3 = w24;// level 5
assign f_4 = w31;// level 6
assign f_5 = w37;// level 7
assign f_6 = w44;// level 7
assign f_7 = w51;// level 7
assign f_8 = w58;// level 7
assign f_9 = w65;// level 7
assign f_10 = w72;// level 9
assign f_11 = w79;// level 8
assign f_12 = w87;// level 9
assign f_13 = w93;// level 11
assign f_14 = w99;// level 10
assign f_15 = w106;// level 8
assign f_16 = w112;// level 9
assign f_17 = w118;// level 9
assign f_18 = w124;// level 10
assign f_19 = w131;// level 9
assign f_20 = w138;// level 10
assign f_21 = w145;// level 10
assign f_22 = w151;// level 9
assign f_23 = w157;// level 10
assign f_24 = w163;// level 9
assign f_25 = w169;// level 10
assign f_26 = w175;// level 10
assign f_27 = w181;// level 9
assign f_28 = w187;// level 10
assign f_29 = w193;// level 10
assign f_30 = w200;// level 11
assign f_31 = w207;// level 10
assign f_32 = w214;// level 10
assign f_33 = w221;// level 11
assign f_34 = w228;// level 11
assign f_35 = w235;// level 11
assign f_36 = w242;// level 11
assign f_37 = w249;// level 11
assign f_38 = w255;// level 12
assign f_39 = w261;// level 12
assign f_40 = w268;// level 10
assign f_41 = w274;// level 11
assign f_42 = w280;// level 10
assign f_43 = w286;// level 11
assign f_44 = w292;// level 11
assign f_45 = w298;// level 11
assign f_46 = w304;// level 11
assign f_47 = w311;// level 12
assign f_48 = w317;// level 12
assign f_49 = w323;// level 12
assign f_50 = w329;// level 12
assign f_51 = w336;// level 12
assign f_52 = w342;// level 12
assign f_53 = w349;// level 12
assign f_54 = w356;// level 12
assign f_55 = w362;// level 12
assign f_56 = w368;// level 12
assign f_57 = w374;// level 12
assign f_58 = w380;// level 12
assign f_59 = w386;// level 12
assign f_60 = w392;// level 12
assign f_61 = w399;// level 12
assign f_62 = w405;// level 12
assign f_63 = w411;// level 12
assign f_64 = w417;// level 12
assign f_65 = w423;// level 12
assign f_66 = w429;// level 12
assign f_67 = w435;// level 12
assign f_68 = w441;// level 12
assign f_69 = w448;// level 12
assign f_70 = w455;// level 12
assign f_71 = w462;// level 12
assign f_72 = w469;// level 12
assign f_73 = w476;// level 12
assign f_74 = w483;// level 12
assign f_75 = w490;// level 12
assign f_76 = w497;// level 12
assign f_77 = w504;// level 12
assign f_78 = w511;// level 11
assign f_79 = w517;// level 11
assign f_80 = w523;// level 11
assign f_81 = w529;// level 12
assign f_82 = w535;// level 12
assign f_83 = w541;// level 12
assign f_84 = w547;// level 11
assign f_85 = w553;// level 11
assign f_86 = w559;// level 11
assign f_87 = w566;// level 12
assign f_88 = w572;// level 12
assign f_89 = w578;// level 12
assign f_90 = w584;// level 12
assign f_91 = w590;// level 12
assign f_92 = w596;// level 12
assign f_93 = w602;// level 12
assign f_94 = w608;// level 12
assign f_95 = w614;// level 12
assign f_96 = w621;// level 12
assign f_97 = w627;// level 12
assign f_98 = w633;// level 12
assign f_99 = w640;// level 12
assign f_100 = w647;// level 12
assign f_101 = w654;// level 12
assign f_102 = w661;// level 12
assign f_103 = w667;// level 12
assign f_104 = w673;// level 12
assign f_105 = w679;// level 12
assign f_106 = w686;// level 12
assign f_107 = w692;// level 12
assign f_108 = w698;// level 12
assign f_109 = w704;// level 12
assign f_110 = w710;// level 12
assign f_111 = w716;// level 12
assign f_112 = w722;// level 12
assign f_113 = w728;// level 12
assign f_114 = w734;// level 12
assign f_115 = w740;// level 12
assign f_116 = w746;// level 12
assign f_117 = w752;// level 12
assign f_118 = w758;// level 12
assign f_119 = w764;// level 12
assign f_120 = w770;// level 12
assign f_121 = w776;// level 12
assign f_122 = w782;// level 12
assign f_123 = w788;// level 12
assign f_124 = w794;// level 12
assign f_125 = w800;// level 12
assign f_126 = w806;// level 12
assign f_127 = w812;// level 12
assign cOut = ~w814;// level 12
endmodule

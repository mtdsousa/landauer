module int2float_best_speed (
        pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, 
        po0, po1, po2, po3, po4, po5, po6);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10;
output po0, po1, po2, po3, po4, po5, po6;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245;
assign w0 = ~pi00 & pi01;
assign w1 = pi00 & ~pi01;
assign w2 = ~w0 & ~w1;
assign w3 = pi04 & ~w2;
assign w4 = pi00 & ~pi04;
assign w5 = ~pi08 & w4;
assign w6 = ~pi07 & w5;
assign w7 = (~pi07 & w3) | (~pi07 & w6) | (w3 & w6);
assign w8 = ~pi06 & w7;
assign w9 = pi04 & pi08;
assign w10 = ~pi04 & ~pi08;
assign w11 = pi03 & w10;
assign w12 = ~pi03 & pi04;
assign w13 = pi07 & w12;
assign w14 = (pi07 & w11) | (pi07 & w13) | (w11 & w13);
assign w15 = ~w9 & ~w14;
assign w16 = ~pi09 & ~w15;
assign w17 = (~pi09 & w8) | (~pi09 & w16) | (w8 & w16);
assign w18 = pi07 & pi10;
assign w19 = ~pi06 & ~w18;
assign w20 = pi02 & ~pi03;
assign w21 = ~pi02 & pi03;
assign w22 = ~w20 & ~w21;
assign w23 = ~pi07 & ~pi09;
assign w24 = ~pi08 & w23;
assign w25 = ~w22 & w24;
assign w26 = pi08 & pi09;
assign w27 = ~pi07 & pi10;
assign w28 = (pi10 & w26) | (pi10 & w27) | (w26 & w27);
assign w29 = pi06 & ~w28;
assign w30 = ~w25 & w29;
assign w31 = ~w19 & ~w30;
assign w32 = ~pi05 & ~pi10;
assign w33 = ~w31 & ~w32;
assign w34 = pi06 & pi09;
assign w35 = w32 & w34;
assign w36 = ~w31 & ~w35;
assign w37 = (~w17 & w33) | (~w17 & w36) | (w33 & w36);
assign w38 = ~pi04 & pi08;
assign w39 = pi04 & ~pi08;
assign w40 = ~pi03 & w39;
assign w41 = pi03 & ~pi04;
assign w42 = pi07 & w41;
assign w43 = (pi07 & w40) | (pi07 & w42) | (w40 & w42);
assign w44 = ~w38 & ~w43;
assign w45 = pi01 & ~pi02;
assign w46 = ~pi01 & pi02;
assign w47 = ~w45 & ~w46;
assign w48 = ~pi07 & ~pi08;
assign w49 = ~pi06 & w48;
assign w50 = ~w47 & w49;
assign w51 = ~pi09 & w50;
assign w52 = (~pi09 & ~w44) | (~pi09 & w51) | (~w44 & w51);
assign w53 = pi05 & ~pi10;
assign w54 = ~pi06 & pi09;
assign w55 = ~pi10 & w54;
assign w56 = pi05 & w55;
assign w57 = (w52 & w53) | (w52 & w56) | (w53 & w56);
assign w58 = w37 & ~w57;
assign w59 = pi02 & pi04;
assign w60 = pi03 & w59;
assign w61 = ~pi02 & ~pi04;
assign w62 = ~pi09 & w61;
assign w63 = (~pi09 & w60) | (~pi09 & w62) | (w60 & w62);
assign w64 = ~pi06 & ~pi10;
assign w65 = (~pi10 & ~w63) | (~pi10 & w64) | (~w63 & w64);
assign w66 = pi06 & ~pi09;
assign w67 = ~pi04 & w66;
assign w68 = pi01 & pi02;
assign w69 = pi05 & ~pi06;
assign w70 = ~w68 & w69;
assign w71 = ~w67 & ~w70;
assign w72 = ~pi03 & ~w71;
assign w73 = w65 & ~w72;
assign w74 = pi06 & pi07;
assign w75 = (pi07 & w64) | (pi07 & w74) | (w64 & w74);
assign w76 = ~pi08 & ~w75;
assign w77 = ~pi06 & pi10;
assign w78 = (~pi08 & w48) | (~pi08 & w77) | (w48 & w77);
assign w79 = (w63 & w76) | (w63 & w78) | (w76 & w78);
assign w80 = ~pi08 & w77;
assign w81 = ~pi06 & ~pi08;
assign w82 = ~w64 & w81;
assign w83 = (w63 & w80) | (w63 & w82) | (w80 & w82);
assign w84 = (~w73 & w79) | (~w73 & w83) | (w79 & w83);
assign w85 = ~pi06 & pi08;
assign w86 = pi07 & ~pi08;
assign w87 = ~pi03 & w86;
assign w88 = ~w85 & ~w87;
assign w89 = ~pi01 & ~pi06;
assign w90 = ~w86 & ~w89;
assign w91 = ~pi04 & ~w90;
assign w92 = w88 & ~w91;
assign w93 = ~pi09 & ~w92;
assign w94 = pi00 & ~pi02;
assign w95 = pi01 & ~pi04;
assign w96 = (pi01 & w94) | (pi01 & w95) | (w94 & w95);
assign w97 = pi00 & pi01;
assign w98 = pi02 & ~w97;
assign w99 = ~w96 & ~w98;
assign w100 = ~pi07 & pi09;
assign w101 = ~w66 & w100;
assign w102 = w32 & w101;
assign w103 = ~pi07 & ~w66;
assign w104 = w32 & w103;
assign w105 = (w99 & w102) | (w99 & w104) | (w102 & w104);
assign w106 = (w32 & w93) | (w32 & w105) | (w93 & w105);
assign w107 = pi06 & ~pi07;
assign w108 = pi09 & w107;
assign w109 = pi03 & pi07;
assign w110 = (pi03 & w68) | (pi03 & w109) | (w68 & w109);
assign w111 = ~pi08 & ~pi09;
assign w112 = ~w110 & w111;
assign w113 = ~w108 & ~w112;
assign w114 = pi04 & ~pi06;
assign w115 = pi08 & w114;
assign w116 = ~pi04 & pi06;
assign w117 = ~pi09 & w116;
assign w118 = (~pi09 & w115) | (~pi09 & w117) | (w115 & w117);
assign w119 = ~pi04 & ~pi09;
assign w120 = ~pi08 & w119;
assign w121 = pi07 & w54;
assign w122 = (pi07 & w120) | (pi07 & w121) | (w120 & w121);
assign w123 = ~w118 & ~w122;
assign w124 = w113 & w123;
assign w125 = w53 & w124;
assign w126 = ~w106 & ~w125;
assign w127 = ~w84 & w126;
assign w128 = pi08 & ~pi09;
assign w129 = w74 & w128;
assign w130 = pi10 & w129;
assign w131 = w127 & ~w130;
assign w132 = ~pi09 & ~pi10;
assign w133 = pi03 & pi04;
assign w134 = pi05 & pi06;
assign w135 = ~w133 & w134;
assign w136 = ~pi01 & w69;
assign w137 = ~pi05 & pi06;
assign w138 = pi02 & w137;
assign w139 = ~w136 & ~w138;
assign w140 = ~w133 & ~w135;
assign w141 = (~w135 & w139) | (~w135 & w140) | (w139 & w140);
assign w142 = ~pi08 & ~w141;
assign w143 = w69 & w133;
assign w144 = pi04 & pi05;
assign w145 = pi06 & ~w144;
assign w146 = ~w143 & ~w145;
assign w147 = pi07 & w132;
assign w148 = ~w146 & w147;
assign w149 = (w132 & w142) | (w132 & w148) | (w142 & w148);
assign w150 = pi01 & ~pi03;
assign w151 = ~pi00 & pi04;
assign w152 = (pi04 & ~w150) | (pi04 & w151) | (~w150 & w151);
assign w153 = pi02 & ~w152;
assign w154 = ~w97 & w133;
assign w155 = ~pi05 & w154;
assign w156 = (~pi05 & w153) | (~pi05 & w155) | (w153 & w155);
assign w157 = ~pi02 & ~pi06;
assign w158 = w133 & w157;
assign w159 = (~pi06 & w156) | (~pi06 & w158) | (w156 & w158);
assign w160 = pi02 & pi03;
assign w161 = w144 & ~w160;
assign w162 = pi04 & ~pi05;
assign w163 = ~pi01 & w162;
assign w164 = ~pi04 & pi05;
assign w165 = pi01 & w164;
assign w166 = ~w163 & ~w165;
assign w167 = ~w160 & ~w161;
assign w168 = (~w161 & w166) | (~w161 & w167) | (w166 & w167);
assign w169 = ~pi08 & ~w168;
assign w170 = (~pi08 & w159) | (~pi08 & w169) | (w159 & w169);
assign w171 = ~pi07 & w132;
assign w172 = w170 & w171;
assign w173 = ~w149 & ~w172;
assign w174 = pi07 & ~pi10;
assign w175 = ~pi06 & w174;
assign w176 = ~pi05 & pi09;
assign w177 = (pi09 & ~w174) | (pi09 & w176) | (~w174 & w176);
assign w178 = ~w175 & ~w177;
assign w179 = ~pi07 & ~pi10;
assign w180 = w144 & w179;
assign w181 = pi06 & w18;
assign w182 = (pi06 & w180) | (pi06 & w181) | (w180 & w181);
assign w183 = w178 & ~w182;
assign w184 = ~pi08 & pi09;
assign w185 = ~pi08 & pi10;
assign w186 = pi09 & w185;
assign w187 = (w183 & w184) | (w183 & w186) | (w184 & w186);
assign w188 = pi08 & ~w183;
assign w189 = ~w187 & ~w188;
assign w190 = w173 & w189;
assign w191 = pi07 & pi08;
assign w192 = pi06 & w191;
assign w193 = ~pi02 & w144;
assign w194 = w192 & w193;
assign w195 = ~pi04 & ~pi05;
assign w196 = w49 & w195;
assign w197 = ~w194 & ~w196;
assign w198 = w132 & ~w197;
assign w199 = ~pi03 & w198;
assign w200 = pi05 & w74;
assign w201 = ~pi06 & ~pi07;
assign w202 = w68 & w201;
assign w203 = ~w200 & ~w202;
assign w204 = ~pi05 & ~pi07;
assign w205 = pi04 & w204;
assign w206 = ~pi03 & ~w204;
assign w207 = pi04 & ~w206;
assign w208 = (~w203 & w205) | (~w203 & w207) | (w205 & w207);
assign w209 = ~pi04 & ~pi07;
assign w210 = (~pi07 & ~w160) | (~pi07 & w209) | (~w160 & w209);
assign w211 = (~pi08 & w81) | (~pi08 & ~w210) | (w81 & ~w210);
assign w212 = ~w208 & w211;
assign w213 = pi04 & w160;
assign w214 = ~pi05 & w97;
assign w215 = w213 & w214;
assign w216 = w81 & w215;
assign w217 = ~w212 & ~w216;
assign w218 = pi03 & pi08;
assign w219 = ~w20 & ~w218;
assign w220 = ~pi09 & ~w219;
assign w221 = pi07 & w134;
assign w222 = pi04 & w221;
assign w223 = w220 & w222;
assign w224 = w134 & w191;
assign w225 = pi09 & ~w224;
assign w226 = ~w223 & ~w225;
assign w227 = w217 & w226;
assign w228 = ~pi10 & ~w227;
assign w229 = ~pi02 & ~pi03;
assign w230 = w9 & ~w229;
assign w231 = w221 & w230;
assign w232 = ~pi05 & ~w97;
assign w233 = (~pi05 & ~w213) | (~pi05 & w232) | (~w213 & w232);
assign w234 = ~pi06 & ~w233;
assign w235 = w144 & w160;
assign w236 = pi06 & ~w235;
assign w237 = ~pi08 & w236;
assign w238 = (~pi08 & w234) | (~pi08 & w237) | (w234 & w237);
assign w239 = pi07 & ~w231;
assign w240 = (~w231 & ~w238) | (~w231 & w239) | (~w238 & w239);
assign w241 = w132 & w240;
assign w242 = pi06 & w235;
assign w243 = ~pi08 & ~w242;
assign w244 = ~pi07 & w243;
assign w245 = w132 & w244;
assign one = 1;
assign po0 = ~w58;
assign po1 = w131;
assign po2 = ~w190;
assign po3 = ~w199;
assign po4 = ~w228;
assign po5 = ~w241;
assign po6 = ~w245;
endmodule

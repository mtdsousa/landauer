module top (
            a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, 
            result_0, result_1, result_2, result_3, result_4, result_5, result_6, result_7, result_8, result_9, result_10, result_11, result_12, result_13, result_14, result_15, result_16, result_17, result_18, result_19, result_20, result_21, result_22, result_23, result_24, result_25, result_26, result_27, result_28, result_29, result_30, result_31);
input a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31;
output result_0, result_1, result_2, result_3, result_4, result_5, result_6, result_7, result_8, result_9, result_10, result_11, result_12, result_13, result_14, result_15, result_16, result_17, result_18, result_19, result_20, result_21, result_22, result_23, result_24, result_25, result_26, result_27, result_28, result_29, result_30, result_31;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583;
assign w0 = ~a_1 & ~a_2;
assign w1 = a_1 & a_2;
assign w2 = ~w0 & ~w1;
assign w3 = a_0 & ~w2;
assign w4 = a_24 & ~a_25;
assign w5 = ~a_23 & ~a_26;
assign w6 = w4 & w5;
assign w7 = ~a_27 & ~a_28;
assign w8 = a_29 & ~a_30;
assign w9 = w7 & w8;
assign w10 = w6 & w9;
assign w11 = ~a_29 & a_30;
assign w12 = a_27 & ~a_28;
assign w13 = w11 & w12;
assign w14 = ~a_24 & ~a_25;
assign w15 = w5 & w14;
assign w16 = w13 & w15;
assign w17 = ~w10 & ~w16;
assign w18 = w9 & w15;
assign w19 = w8 & w12;
assign w20 = a_23 & ~a_26;
assign w21 = ~a_24 & a_25;
assign w22 = w20 & w21;
assign w23 = w19 & w22;
assign w24 = ~w18 & ~w23;
assign w25 = ~a_23 & a_26;
assign w26 = w21 & w25;
assign w27 = ~a_27 & a_28;
assign w28 = a_29 & a_30;
assign w29 = w27 & w28;
assign w30 = w26 & w29;
assign w31 = a_27 & a_28;
assign w32 = w11 & w31;
assign w33 = w14 & w20;
assign w34 = w32 & w33;
assign w35 = ~a_29 & ~a_30;
assign w36 = w27 & w35;
assign w37 = a_24 & a_25;
assign w38 = w20 & w37;
assign w39 = w36 & w38;
assign w40 = w8 & w27;
assign w41 = w5 & w37;
assign w42 = w40 & w41;
assign w43 = ~w39 & ~w42;
assign w44 = w31 & w35;
assign w45 = w38 & w44;
assign w46 = w6 & w44;
assign w47 = w7 & w35;
assign w48 = a_23 & a_26;
assign w49 = w37 & w48;
assign w50 = w47 & w49;
assign w51 = ~w46 & ~w50;
assign w52 = ~w45 & w51;
assign w53 = w33 & w47;
assign w54 = w7 & w11;
assign w55 = w4 & w25;
assign w56 = w54 & w55;
assign w57 = ~w53 & ~w56;
assign w58 = w7 & w28;
assign w59 = w21 & w48;
assign w60 = w58 & w59;
assign w61 = w14 & w25;
assign w62 = w29 & w61;
assign w63 = ~w60 & ~w62;
assign w64 = w57 & w63;
assign w65 = w15 & w40;
assign w66 = w14 & w48;
assign w67 = w13 & w66;
assign w68 = w36 & w61;
assign w69 = ~w65 & ~w67;
assign w70 = ~w68 & w69;
assign w71 = w29 & w33;
assign w72 = w9 & w26;
assign w73 = ~w71 & ~w72;
assign w74 = w29 & w49;
assign w75 = w13 & w59;
assign w76 = w19 & w26;
assign w77 = ~w75 & ~w76;
assign w78 = ~w74 & w77;
assign w79 = w4 & w20;
assign w80 = w28 & w31;
assign w81 = w79 & w80;
assign w82 = w11 & w27;
assign w83 = w38 & w82;
assign w84 = ~w81 & ~w83;
assign w85 = w22 & w36;
assign w86 = w6 & w82;
assign w87 = w8 & w31;
assign w88 = w66 & w87;
assign w89 = w32 & w38;
assign w90 = ~w88 & ~w89;
assign w91 = ~w86 & w90;
assign w92 = w90 & w32636;
assign w93 = w25 & w37;
assign w94 = w9 & w93;
assign w95 = w32 & w41;
assign w96 = ~w94 & ~w95;
assign w97 = w58 & w61;
assign w98 = w26 & w80;
assign w99 = ~w97 & ~w98;
assign w100 = w84 & w96;
assign w101 = w99 & w100;
assign w102 = w101 & w32637;
assign w103 = ~w30 & ~w34;
assign w104 = w17 & w103;
assign w105 = w24 & w43;
assign w106 = w73 & w105;
assign w107 = w52 & w104;
assign w108 = w64 & w70;
assign w109 = w107 & w108;
assign w110 = w106 & w109;
assign w111 = w102 & w110;
assign w112 = w44 & w49;
assign w113 = w32 & w59;
assign w114 = ~w112 & ~w113;
assign w115 = w61 & w82;
assign w116 = w6 & w58;
assign w117 = w4 & w48;
assign w118 = w32 & w117;
assign w119 = ~w115 & ~w116;
assign w120 = ~w118 & w119;
assign w121 = w114 & w120;
assign w122 = w12 & w35;
assign w123 = w93 & w122;
assign w124 = w47 & w79;
assign w125 = w29 & w59;
assign w126 = w15 & w32;
assign w127 = w79 & w122;
assign w128 = w36 & w49;
assign w129 = ~w127 & ~w128;
assign w130 = w38 & w40;
assign w131 = w9 & w117;
assign w132 = ~w130 & ~w131;
assign w133 = w129 & w132;
assign w134 = w33 & w122;
assign w135 = w66 & w122;
assign w136 = w9 & w41;
assign w137 = ~w135 & ~w136;
assign w138 = w40 & w117;
assign w139 = w12 & w28;
assign w140 = w22 & w139;
assign w141 = ~w138 & ~w140;
assign w142 = w66 & w139;
assign w143 = w40 & w93;
assign w144 = w19 & w41;
assign w145 = ~w143 & ~w144;
assign w146 = w19 & w49;
assign w147 = w15 & w29;
assign w148 = ~w146 & ~w147;
assign w149 = w117 & w139;
assign w150 = w148 & ~w149;
assign w151 = w33 & w58;
assign w152 = w6 & w19;
assign w153 = w36 & w79;
assign w154 = ~w151 & ~w152;
assign w155 = ~w153 & w154;
assign w156 = w54 & w93;
assign w157 = w6 & w32;
assign w158 = ~w156 & ~w157;
assign w159 = w59 & w82;
assign w160 = w5 & w21;
assign w161 = w80 & w160;
assign w162 = ~w159 & ~w161;
assign w163 = w15 & w36;
assign w164 = w49 & w54;
assign w165 = ~w163 & ~w164;
assign w166 = w36 & w55;
assign w167 = w38 & w58;
assign w168 = ~w166 & ~w167;
assign w169 = w33 & w82;
assign w170 = w9 & w61;
assign w171 = ~w169 & ~w170;
assign w172 = w55 & w139;
assign w173 = w44 & w160;
assign w174 = ~w172 & ~w173;
assign w175 = w168 & w171;
assign w176 = w174 & w175;
assign w177 = w36 & w59;
assign w178 = w22 & w47;
assign w179 = ~w177 & ~w178;
assign w180 = w26 & w36;
assign w181 = w55 & w87;
assign w182 = ~w180 & ~w181;
assign w183 = w47 & w117;
assign w184 = ~a_24 & w25;
assign w185 = w13 & w184;
assign w186 = ~a_25 & w185;
assign w187 = ~w183 & ~w186;
assign w188 = w6 & w87;
assign w189 = ~w186 & w32638;
assign w190 = w9 & w22;
assign w191 = w22 & w87;
assign w192 = ~w190 & ~w191;
assign w193 = ~w6 & ~w38;
assign w194 = w54 & ~w193;
assign w195 = w13 & w160;
assign w196 = w59 & w87;
assign w197 = w54 & w117;
assign w198 = ~w196 & ~w197;
assign w199 = ~w194 & ~w195;
assign w200 = w198 & w199;
assign w201 = w179 & w182;
assign w202 = w192 & w201;
assign w203 = w189 & w202;
assign w204 = w200 & w203;
assign w205 = w44 & w55;
assign w206 = w13 & w79;
assign w207 = w22 & w80;
assign w208 = w87 & w93;
assign w209 = ~w207 & ~w208;
assign w210 = ~w206 & w209;
assign w211 = w209 & w32639;
assign w212 = w33 & w87;
assign w213 = w26 & w58;
assign w214 = w13 & w26;
assign w215 = ~w213 & ~w214;
assign w216 = w41 & w87;
assign w217 = w49 & w139;
assign w218 = w26 & w32;
assign w219 = ~w217 & ~w218;
assign w220 = w139 & w160;
assign w221 = w55 & w122;
assign w222 = ~w220 & ~w221;
assign w223 = ~w212 & ~w216;
assign w224 = w215 & w223;
assign w225 = w219 & w222;
assign w226 = w224 & w225;
assign w227 = w145 & w158;
assign w228 = w162 & w165;
assign w229 = w227 & w228;
assign w230 = w150 & w155;
assign w231 = w229 & w230;
assign w232 = w176 & w211;
assign w233 = w226 & w232;
assign w234 = w231 & w233;
assign w235 = w204 & w234;
assign w236 = w234 & w32640;
assign w237 = w47 & w59;
assign w238 = w82 & w117;
assign w239 = w13 & w93;
assign w240 = ~w238 & ~w239;
assign w241 = ~w237 & w240;
assign w242 = w19 & w61;
assign w243 = w9 & w66;
assign w244 = ~w242 & ~w243;
assign w245 = w80 & w117;
assign w246 = w38 & w122;
assign w247 = ~w245 & ~w246;
assign w248 = w41 & w82;
assign w249 = w9 & w79;
assign w250 = ~w248 & ~w249;
assign w251 = w19 & w66;
assign w252 = w38 & w47;
assign w253 = ~w251 & ~w252;
assign w254 = w26 & w82;
assign w255 = w33 & w54;
assign w256 = w41 & w54;
assign w257 = ~w255 & ~w256;
assign w258 = ~w254 & w257;
assign w259 = w253 & w258;
assign w260 = w58 & w93;
assign w261 = w29 & w38;
assign w262 = w26 & w122;
assign w263 = ~w261 & ~w262;
assign w264 = w41 & w80;
assign w265 = w44 & w59;
assign w266 = w47 & w66;
assign w267 = w9 & w49;
assign w268 = ~w266 & ~w267;
assign w269 = ~w260 & ~w264;
assign w270 = ~w265 & w269;
assign w271 = w263 & w268;
assign w272 = w270 & w271;
assign w273 = w244 & w247;
assign w274 = w250 & w273;
assign w275 = w241 & w274;
assign w276 = w259 & w272;
assign w277 = w275 & w276;
assign w278 = w29 & w41;
assign w279 = w58 & w79;
assign w280 = ~w278 & ~w279;
assign w281 = w29 & w93;
assign w282 = w22 & w44;
assign w283 = w79 & w139;
assign w284 = ~w282 & ~w283;
assign w285 = w280 & ~w281;
assign w286 = w284 & w285;
assign w287 = w40 & w55;
assign w288 = w40 & w79;
assign w289 = ~w287 & ~w288;
assign w290 = w22 & w122;
assign w291 = w59 & w80;
assign w292 = w79 & w82;
assign w293 = ~w291 & ~w292;
assign w294 = w289 & ~w290;
assign w295 = w293 & w294;
assign w296 = ~w123 & ~w124;
assign w297 = ~w125 & ~w126;
assign w298 = ~w134 & w297;
assign w299 = w137 & w296;
assign w300 = w141 & w299;
assign w301 = w133 & w298;
assign w302 = w300 & w301;
assign w303 = w121 & w286;
assign w304 = w295 & w303;
assign w305 = w302 & w304;
assign w306 = w277 & w305;
assign w307 = w111 & w306;
assign w308 = w236 & w307;
assign w309 = w54 & w59;
assign w310 = ~w94 & ~w309;
assign w311 = ~w34 & ~w177;
assign w312 = w36 & w93;
assign w313 = w32 & w79;
assign w314 = w38 & w139;
assign w315 = w117 & w122;
assign w316 = w6 & w122;
assign w317 = ~w10 & ~w316;
assign w318 = ~w123 & w317;
assign w319 = w6 & w80;
assign w320 = ~w125 & ~w319;
assign w321 = w40 & w59;
assign w322 = w15 & w82;
assign w323 = w44 & w93;
assign w324 = ~w322 & ~w323;
assign w325 = w6 & w47;
assign w326 = ~w144 & ~w321;
assign w327 = ~w325 & w326;
assign w328 = w324 & w327;
assign w329 = ~w312 & ~w313;
assign w330 = ~w314 & ~w315;
assign w331 = w329 & w330;
assign w332 = w310 & w311;
assign w333 = w320 & w332;
assign w334 = w318 & w331;
assign w335 = w333 & w334;
assign w336 = w328 & w335;
assign w337 = w9 & w55;
assign w338 = ~w98 & ~w248;
assign w339 = w19 & w38;
assign w340 = ~w23 & ~w339;
assign w341 = w36 & w66;
assign w342 = w55 & w82;
assign w343 = ~w188 & ~w342;
assign w344 = ~w341 & w343;
assign w345 = w41 & w139;
assign w346 = ~w138 & ~w170;
assign w347 = ~w56 & ~w345;
assign w348 = w346 & w347;
assign w349 = w29 & w160;
assign w350 = w19 & w93;
assign w351 = ~w349 & ~w350;
assign w352 = w87 & w160;
assign w353 = ~w288 & ~w352;
assign w354 = w351 & w353;
assign w355 = w49 & w122;
assign w356 = w44 & w66;
assign w357 = w32 & w160;
assign w358 = ~w356 & ~w357;
assign w359 = ~w76 & ~w167;
assign w360 = ~w113 & ~w245;
assign w361 = w359 & w360;
assign w362 = w13 & w22;
assign w363 = w13 & w41;
assign w364 = ~w362 & ~w363;
assign w365 = w19 & w59;
assign w366 = w29 & w79;
assign w367 = ~w365 & ~w366;
assign w368 = w44 & w79;
assign w369 = w40 & w160;
assign w370 = ~w368 & ~w369;
assign w371 = ~w71 & ~w355;
assign w372 = w358 & w371;
assign w373 = w364 & w367;
assign w374 = w370 & w373;
assign w375 = w354 & w372;
assign w376 = w361 & w375;
assign w377 = w374 & w376;
assign w378 = w13 & w49;
assign w379 = ~w115 & ~w378;
assign w380 = w66 & w82;
assign w381 = ~w287 & ~w380;
assign w382 = ~w134 & ~w218;
assign w383 = w379 & w382;
assign w384 = w381 & w383;
assign w385 = w15 & w19;
assign w386 = ~w265 & ~w385;
assign w387 = ~w46 & ~w153;
assign w388 = w19 & w33;
assign w389 = w58 & w66;
assign w390 = ~w249 & ~w389;
assign w391 = w61 & w139;
assign w392 = w15 & w58;
assign w393 = w41 & w47;
assign w394 = w22 & w40;
assign w395 = w58 & w117;
assign w396 = w80 & w93;
assign w397 = ~w30 & ~w396;
assign w398 = ~w118 & ~w237;
assign w399 = w54 & w79;
assign w400 = w47 & w93;
assign w401 = ~w53 & ~w399;
assign w402 = ~w400 & w401;
assign w403 = w26 & w54;
assign w404 = w49 & w80;
assign w405 = ~w403 & ~w404;
assign w406 = w26 & w40;
assign w407 = ~w97 & ~w406;
assign w408 = ~w135 & ~w391;
assign w409 = ~w392 & ~w393;
assign w410 = ~w394 & ~w395;
assign w411 = w409 & w410;
assign w412 = w397 & w408;
assign w413 = w398 & w405;
assign w414 = w407 & w413;
assign w415 = w411 & w412;
assign w416 = w402 & w415;
assign w417 = w414 & w416;
assign w418 = w54 & w160;
assign w419 = ~w157 & ~w418;
assign w420 = w36 & w160;
assign w421 = ~w180 & ~w420;
assign w422 = w6 & w29;
assign w423 = w22 & w54;
assign w424 = ~w422 & ~w423;
assign w425 = ~w255 & w419;
assign w426 = w421 & w424;
assign w427 = w425 & w426;
assign w428 = w15 & w80;
assign w429 = w32 & w49;
assign w430 = ~w428 & ~w429;
assign w431 = w9 & w160;
assign w432 = w13 & w38;
assign w433 = ~w431 & ~w432;
assign w434 = ~w197 & ~w217;
assign w435 = ~w281 & ~w388;
assign w436 = w434 & w435;
assign w437 = w386 & w387;
assign w438 = w390 & w430;
assign w439 = w433 & w438;
assign w440 = w436 & w437;
assign w441 = w439 & w440;
assign w442 = w384 & w427;
assign w443 = w441 & w442;
assign w444 = w417 & w443;
assign w445 = ~w126 & ~w283;
assign w446 = w26 & w87;
assign w447 = w22 & w29;
assign w448 = ~w446 & ~w447;
assign w449 = ~w220 & ~w243;
assign w450 = w55 & w58;
assign w451 = w32 & w93;
assign w452 = ~w291 & ~w451;
assign w453 = ~w75 & ~w195;
assign w454 = ~w206 & w453;
assign w455 = ~w266 & ~w450;
assign w456 = w452 & w455;
assign w457 = w454 & w456;
assign w458 = w41 & w122;
assign w459 = w47 & w55;
assign w460 = ~w290 & ~w459;
assign w461 = ~w68 & w460;
assign w462 = w460 & w31560;
assign w463 = w44 & w61;
assign w464 = ~w181 & ~w463;
assign w465 = ~w74 & ~w221;
assign w466 = ~w45 & ~w239;
assign w467 = ~w83 & ~w147;
assign w468 = w79 & w87;
assign w469 = ~w212 & ~w468;
assign w470 = w6 & w54;
assign w471 = ~w39 & ~w214;
assign w472 = ~w470 & w471;
assign w473 = w87 & w117;
assign w474 = ~w178 & ~w473;
assign w475 = w22 & w32;
assign w476 = w33 & w80;
assign w477 = ~w475 & ~w476;
assign w478 = ~w267 & w477;
assign w479 = w464 & w465;
assign w480 = w466 & w467;
assign w481 = w469 & w474;
assign w482 = w480 & w481;
assign w483 = w472 & w479;
assign w484 = w478 & w483;
assign w485 = w462 & w482;
assign w486 = w484 & w485;
assign w487 = ~w88 & ~w140;
assign w488 = ~w337 & w487;
assign w489 = w338 & w340;
assign w490 = w445 & w448;
assign w491 = w449 & w490;
assign w492 = w488 & w489;
assign w493 = w344 & w348;
assign w494 = w492 & w493;
assign w495 = w457 & w491;
assign w496 = w494 & w495;
assign w497 = w336 & w496;
assign w498 = w377 & w486;
assign w499 = w497 & w498;
assign w500 = w444 & w499;
assign w501 = ~w308 & ~w500;
assign w502 = ~a_20 & ~a_21;
assign w503 = a_20 & a_21;
assign w504 = ~w502 & ~w503;
assign w505 = ~a_21 & ~a_22;
assign w506 = a_21 & a_22;
assign w507 = ~w505 & ~w506;
assign w508 = ~w504 & ~w507;
assign w509 = a_23 & ~w508;
assign w510 = ~a_22 & w502;
assign w511 = (~w510 & w508) | (~w510 & w32641) | (w508 & w32641);
assign w512 = w308 & w500;
assign w513 = ~w501 & ~w512;
assign w514 = ~w511 & w513;
assign w515 = (~w501 & ~w513) | (~w501 & w32642) | (~w513 & w32642);
assign w516 = ~w188 & w469;
assign w517 = ~w39 & ~w264;
assign w518 = ~w38 & ~w61;
assign w519 = (w80 & ~w518) | (w80 & w81) | (~w518 & w81);
assign w520 = ~w161 & ~w476;
assign w521 = ~w519 & w520;
assign w522 = ~w74 & ~w428;
assign w523 = ~w207 & w320;
assign w524 = w522 & w523;
assign w525 = w521 & w524;
assign w526 = w516 & w517;
assign w527 = w525 & w526;
assign w528 = w525 & w32643;
assign w529 = ~w255 & ~w369;
assign w530 = w40 & w61;
assign w531 = w41 & w44;
assign w532 = ~w394 & ~w531;
assign w533 = ~w42 & ~w288;
assign w534 = w284 & ~w530;
assign w535 = w529 & w532;
assign w536 = w533 & w535;
assign w537 = w534 & w536;
assign w538 = w6 & w36;
assign w539 = ~w130 & ~w220;
assign w540 = w54 & w66;
assign w541 = w13 & w55;
assign w542 = ~w540 & ~w541;
assign w543 = w33 & w36;
assign w544 = w19 & w117;
assign w545 = ~w543 & ~w544;
assign w546 = w542 & w545;
assign w547 = w19 & w55;
assign w548 = ~w30 & ~w547;
assign w549 = ~w72 & ~w337;
assign w550 = ~w131 & ~w243;
assign w551 = ~w400 & ~w538;
assign w552 = w539 & w551;
assign w553 = w548 & w549;
assign w554 = w550 & w553;
assign w555 = w546 & w552;
assign w556 = w554 & w555;
assign w557 = ~w18 & ~w191;
assign w558 = w340 & w557;
assign w559 = w9 & w33;
assign w560 = ~w323 & ~w559;
assign w561 = ~w218 & ~w429;
assign w562 = w22 & w58;
assign w563 = w58 & w160;
assign w564 = ~w451 & ~w563;
assign w565 = w561 & ~w562;
assign w566 = w564 & w565;
assign w567 = ~w140 & ~w142;
assign w568 = w55 & w80;
assign w569 = ~w392 & ~w568;
assign w570 = ~w163 & ~w355;
assign w571 = ~w151 & ~w159;
assign w572 = w26 & w139;
assign w573 = ~w50 & ~w572;
assign w574 = ~w178 & ~w393;
assign w575 = ~w242 & w574;
assign w576 = ~w254 & w364;
assign w577 = w571 & w573;
assign w578 = w576 & w577;
assign w579 = w575 & w578;
assign w580 = w38 & w87;
assign w581 = ~w345 & ~w580;
assign w582 = w15 & w122;
assign w583 = w9 & w59;
assign w584 = ~w582 & ~w583;
assign w585 = w59 & w139;
assign w586 = ~w170 & ~w585;
assign w587 = ~w246 & ~w418;
assign w588 = ~w186 & w587;
assign w589 = w40 & w66;
assign w590 = w15 & w47;
assign w591 = ~w342 & ~w590;
assign w592 = ~w589 & w591;
assign w593 = w47 & w61;
assign w594 = ~w149 & ~w593;
assign w595 = ~w216 & w594;
assign w596 = ~w67 & ~w144;
assign w597 = w93 & w139;
assign w598 = ~w248 & ~w597;
assign w599 = ~w123 & w596;
assign w600 = w598 & w599;
assign w601 = w595 & w600;
assign w602 = ~w251 & ~w423;
assign w603 = ~w314 & ~w352;
assign w604 = ~w279 & ~w380;
assign w605 = ~w368 & ~w399;
assign w606 = ~w68 & w581;
assign w607 = w584 & w586;
assign w608 = w602 & w603;
assign w609 = w604 & w605;
assign w610 = w608 & w609;
assign w611 = w606 & w607;
assign w612 = w588 & w592;
assign w613 = w611 & w612;
assign w614 = w121 & w610;
assign w615 = w613 & w614;
assign w616 = w601 & w615;
assign w617 = ~w46 & ~w470;
assign w618 = ~w458 & w617;
assign w619 = w38 & w54;
assign w620 = ~w195 & ~w619;
assign w621 = ~w238 & w620;
assign w622 = w61 & w87;
assign w623 = w54 & w61;
assign w624 = ~w622 & ~w623;
assign w625 = ~w391 & w624;
assign w626 = w66 & w80;
assign w627 = ~w341 & ~w626;
assign w628 = ~w83 & ~w206;
assign w629 = w627 & w628;
assign w630 = ~w256 & ~w432;
assign w631 = w174 & w630;
assign w632 = w560 & w567;
assign w633 = w569 & w570;
assign w634 = w632 & w633;
assign w635 = w558 & w631;
assign w636 = w618 & w621;
assign w637 = w625 & w629;
assign w638 = w636 & w637;
assign w639 = w634 & w635;
assign w640 = w566 & w639;
assign w641 = w579 & w638;
assign w642 = w640 & w641;
assign w643 = w616 & w642;
assign w644 = w82 & w93;
assign w645 = w41 & w58;
assign w646 = ~w644 & ~w645;
assign w647 = w36 & w117;
assign w648 = ~w166 & ~w647;
assign w649 = w13 & w117;
assign w650 = ~w237 & ~w649;
assign w651 = ~w290 & w650;
assign w652 = w49 & w82;
assign w653 = w61 & w122;
assign w654 = ~w265 & ~w653;
assign w655 = ~w281 & ~w652;
assign w656 = w646 & w655;
assign w657 = w648 & w654;
assign w658 = w656 & w657;
assign w659 = w651 & w658;
assign w660 = w537 & w659;
assign w661 = w556 & w660;
assign w662 = w528 & w661;
assign w663 = w643 & w662;
assign w664 = ~w515 & w663;
assign w665 = w515 & ~w663;
assign w666 = ~w664 & ~w665;
assign w667 = ~a_31 & ~w35;
assign w668 = ~w28 & w667;
assign w669 = ~w45 & ~w190;
assign w670 = ~w342 & ~w652;
assign w671 = w15 & w54;
assign w672 = ~w65 & ~w671;
assign w673 = ~w134 & ~w207;
assign w674 = ~w319 & w673;
assign w675 = ~w136 & ~w400;
assign w676 = ~w81 & w675;
assign w677 = ~w151 & ~w180;
assign w678 = ~w356 & ~w541;
assign w679 = w677 & w678;
assign w680 = ~w125 & ~w246;
assign w681 = ~w220 & ~w589;
assign w682 = ~w178 & ~w218;
assign w683 = ~w403 & w682;
assign w684 = w340 & w669;
assign w685 = w670 & w672;
assign w686 = w680 & w681;
assign w687 = w685 & w686;
assign w688 = w683 & w684;
assign w689 = w674 & w676;
assign w690 = w679 & w689;
assign w691 = w687 & w688;
assign w692 = w690 & w691;
assign w693 = ~w161 & ~w355;
assign w694 = w13 & w33;
assign w695 = ~w590 & ~w694;
assign w696 = w6 & w40;
assign w697 = ~w170 & ~w216;
assign w698 = w33 & w139;
assign w699 = ~w647 & ~w698;
assign w700 = w697 & w699;
assign w701 = w33 & w40;
assign w702 = ~w53 & ~w701;
assign w703 = w693 & ~w696;
assign w704 = w695 & w702;
assign w705 = w703 & w704;
assign w706 = w700 & w705;
assign w707 = a_23 & w37;
assign w708 = w9 & w707;
assign w709 = ~w316 & ~w708;
assign w710 = w47 & w160;
assign w711 = ~w323 & ~w463;
assign w712 = ~w593 & w711;
assign w713 = ~w399 & ~w418;
assign w714 = w49 & w87;
assign w715 = ~w309 & ~w714;
assign w716 = w713 & w715;
assign w717 = ~w163 & ~w191;
assign w718 = ~w251 & w717;
assign w719 = w6 & w139;
assign w720 = w26 & w47;
assign w721 = ~w146 & ~w720;
assign w722 = ~w266 & ~w350;
assign w723 = ~w159 & ~w719;
assign w724 = w721 & w723;
assign w725 = w722 & w724;
assign w726 = ~w138 & ~w644;
assign w727 = ~w580 & w726;
assign w728 = ~w94 & ~w290;
assign w729 = ~w242 & w728;
assign w730 = w29 & w66;
assign w731 = ~w281 & ~w730;
assign w732 = w29 & w117;
assign w733 = ~w287 & ~w732;
assign w734 = w33 & w44;
assign w735 = ~w322 & ~w734;
assign w736 = ~w164 & ~w172;
assign w737 = w15 & w44;
assign w738 = ~w279 & ~w737;
assign w739 = ~w254 & ~w562;
assign w740 = w564 & w739;
assign w741 = w29 & w55;
assign w742 = ~w46 & ~w741;
assign w743 = ~w157 & ~w392;
assign w744 = ~w169 & ~w378;
assign w745 = ~w85 & w735;
assign w746 = w736 & w738;
assign w747 = w742 & w743;
assign w748 = w744 & w747;
assign w749 = w745 & w746;
assign w750 = w740 & w749;
assign w751 = w748 & w750;
assign w752 = ~w75 & ~w429;
assign w753 = ~w221 & ~w391;
assign w754 = ~w34 & ~w74;
assign w755 = ~w140 & ~w385;
assign w756 = ~w126 & ~w530;
assign w757 = ~w214 & ~w406;
assign w758 = ~w149 & ~w345;
assign w759 = ~w314 & w756;
assign w760 = w757 & w758;
assign w761 = w759 & w760;
assign w762 = w731 & w733;
assign w763 = w752 & w753;
assign w764 = w754 & w755;
assign w765 = w763 & w764;
assign w766 = w241 & w762;
assign w767 = w727 & w729;
assign w768 = w766 & w767;
assign w769 = w725 & w765;
assign w770 = w761 & w769;
assign w771 = w768 & w770;
assign w772 = w751 & w771;
assign w773 = ~w30 & ~w255;
assign w774 = ~w113 & ~w315;
assign w775 = ~w18 & ~w583;
assign w776 = w6 & w13;
assign w777 = ~w144 & ~w776;
assign w778 = ~w468 & ~w543;
assign w779 = ~w116 & ~w283;
assign w780 = ~w16 & ~w428;
assign w781 = ~w470 & w780;
assign w782 = w773 & w774;
assign w783 = w775 & w777;
assign w784 = w778 & w779;
assign w785 = w783 & w784;
assign w786 = w781 & w782;
assign w787 = w785 & w786;
assign w788 = ~w166 & ~w458;
assign w789 = w36 & w41;
assign w790 = ~w262 & ~w789;
assign w791 = ~w142 & ~w156;
assign w792 = ~w352 & ~w622;
assign w793 = ~w649 & w792;
assign w794 = ~w112 & ~w476;
assign w795 = ~w710 & w794;
assign w796 = w709 & w788;
assign w797 = w790 & w791;
assign w798 = w796 & w797;
assign w799 = w712 & w795;
assign w800 = w716 & w718;
assign w801 = w793 & w800;
assign w802 = w798 & w799;
assign w803 = w801 & w802;
assign w804 = w706 & w787;
assign w805 = w803 & w804;
assign w806 = w692 & w805;
assign w807 = w772 & w806;
assign w808 = ~w245 & ~w404;
assign w809 = ~w254 & ~w256;
assign w810 = ~w128 & ~w159;
assign w811 = ~w188 & w809;
assign w812 = w810 & w811;
assign w813 = ~w698 & ~w734;
assign w814 = ~w34 & ~w395;
assign w815 = w40 & w49;
assign w816 = ~w380 & ~w815;
assign w817 = ~w115 & ~w172;
assign w818 = w15 & w139;
assign w819 = ~w538 & ~w818;
assign w820 = ~w53 & ~w212;
assign w821 = ~w142 & ~w260;
assign w822 = ~w267 & ~w719;
assign w823 = ~w72 & ~w315;
assign w824 = ~w696 & w823;
assign w825 = w753 & w817;
assign w826 = w819 & w820;
assign w827 = w821 & w822;
assign w828 = w826 & w827;
assign w829 = w824 & w825;
assign w830 = w828 & w829;
assign w831 = a_27 & w35;
assign w832 = w26 & w831;
assign w833 = ~w85 & ~w146;
assign w834 = w15 & w87;
assign w835 = ~w94 & ~w834;
assign w836 = ~w191 & ~w580;
assign w837 = ~w216 & w836;
assign w838 = w49 & w58;
assign w839 = ~w131 & ~w838;
assign w840 = ~w694 & ~w776;
assign w841 = ~w140 & ~w197;
assign w842 = ~w291 & ~w423;
assign w843 = ~w450 & ~w653;
assign w844 = w842 & w843;
assign w845 = w833 & w841;
assign w846 = w835 & w839;
assign w847 = w840 & w846;
assign w848 = w844 & w845;
assign w849 = w837 & w848;
assign w850 = w847 & w849;
assign w851 = ~w337 & ~w832;
assign w852 = w849 & w32644;
assign w853 = ~w157 & ~w205;
assign w854 = ~w314 & w853;
assign w855 = ~w352 & ~w652;
assign w856 = w80 & w31561;
assign w857 = ~w16 & ~w164;
assign w858 = ~w18 & ~w396;
assign w859 = w449 & w591;
assign w860 = w855 & ~w856;
assign w861 = w857 & w858;
assign w862 = w860 & w861;
assign w863 = w854 & w859;
assign w864 = w862 & w863;
assign w865 = ~w60 & ~w238;
assign w866 = ~w167 & ~w389;
assign w867 = ~w248 & ~w737;
assign w868 = a_25 & w25;
assign w869 = w54 & w868;
assign w870 = w6 & w831;
assign w871 = ~w547 & ~w644;
assign w872 = ~w292 & w584;
assign w873 = w871 & w872;
assign w874 = ~w83 & ~w420;
assign w875 = ~w65 & ~w593;
assign w876 = ~w98 & ~w568;
assign w877 = ~w135 & ~w252;
assign w878 = w82 & w160;
assign w879 = ~w76 & ~w878;
assign w880 = w876 & w877;
assign w881 = w879 & w880;
assign w882 = ~w323 & ~w468;
assign w883 = ~w701 & ~w869;
assign w884 = ~w870 & w883;
assign w885 = w624 & w882;
assign w886 = w865 & w866;
assign w887 = w867 & w874;
assign w888 = w875 & w887;
assign w889 = w885 & w886;
assign w890 = w884 & w889;
assign w891 = w873 & w888;
assign w892 = w881 & w891;
assign w893 = w864 & w890;
assign w894 = w892 & w893;
assign w895 = w38 & w80;
assign w896 = w22 & w82;
assign w897 = ~w213 & ~w895;
assign w898 = ~w896 & w897;
assign w899 = ~w134 & ~w312;
assign w900 = ~w540 & w899;
assign w901 = w722 & w758;
assign w902 = w900 & w901;
assign w903 = w898 & w902;
assign w904 = w902 & w32645;
assign w905 = ~w365 & ~w544;
assign w906 = ~w645 & w905;
assign w907 = w44 & w117;
assign w908 = ~w50 & ~w177;
assign w909 = ~w619 & ~w907;
assign w910 = w908 & w909;
assign w911 = ~w112 & ~w143;
assign w912 = ~w309 & w911;
assign w913 = ~w153 & ~w393;
assign w914 = ~w264 & ~w789;
assign w915 = w913 & w914;
assign w916 = ~w56 & ~w86;
assign w917 = ~w321 & w916;
assign w918 = w386 & w445;
assign w919 = w808 & w813;
assign w920 = w814 & w816;
assign w921 = w919 & w920;
assign w922 = w917 & w918;
assign w923 = w906 & w910;
assign w924 = w912 & w915;
assign w925 = w923 & w924;
assign w926 = w921 & w922;
assign w927 = w812 & w926;
assign w928 = w830 & w925;
assign w929 = w927 & w928;
assign w930 = w904 & w929;
assign w931 = w852 & w894;
assign w932 = w930 & w931;
assign w933 = ~w807 & w932;
assign w934 = ~w714 & ~w838;
assign w935 = ~w216 & ~w896;
assign w936 = ~w127 & ~w708;
assign w937 = w935 & w936;
assign w938 = ~w393 & ~w450;
assign w939 = ~w152 & ~w696;
assign w940 = w938 & w939;
assign w941 = ~w256 & ~w391;
assign w942 = ~w188 & ~w404;
assign w943 = w941 & w942;
assign w944 = w87 & w868;
assign w945 = ~w341 & ~w349;
assign w946 = ~w246 & ~w815;
assign w947 = ~w143 & ~w582;
assign w948 = ~w76 & ~w169;
assign w949 = ~w97 & ~w345;
assign w950 = ~w126 & ~w249;
assign w951 = ~w547 & w950;
assign w952 = ~w149 & ~w281;
assign w953 = ~w262 & ~w420;
assign w954 = ~w136 & w952;
assign w955 = w953 & w954;
assign w956 = ~w72 & ~w245;
assign w957 = ~w357 & ~w622;
assign w958 = ~w265 & ~w626;
assign w959 = ~w42 & ~w50;
assign w960 = ~w68 & ~w647;
assign w961 = ~w157 & ~w243;
assign w962 = ~w447 & ~w593;
assign w963 = ~w473 & ~w597;
assign w964 = w956 & w963;
assign w965 = w957 & w958;
assign w966 = w959 & w960;
assign w967 = w961 & w962;
assign w968 = w966 & w967;
assign w969 = w964 & w965;
assign w970 = w968 & w969;
assign w971 = ~w65 & ~w944;
assign w972 = w934 & w971;
assign w973 = w945 & w946;
assign w974 = w947 & w948;
assign w975 = w949 & w974;
assign w976 = w972 & w973;
assign w977 = w937 & w940;
assign w978 = w943 & w951;
assign w979 = w977 & w978;
assign w980 = w975 & w976;
assign w981 = w955 & w980;
assign w982 = w970 & w979;
assign w983 = w981 & w982;
assign w984 = ~w197 & ~w312;
assign w985 = ~w544 & w984;
assign w986 = ~w403 & ~w540;
assign w987 = w628 & w986;
assign w988 = ~w170 & ~w431;
assign w989 = ~w583 & w988;
assign w990 = ~w283 & ~w362;
assign w991 = w520 & w990;
assign w992 = w122 & w160;
assign w993 = ~w818 & ~w992;
assign w994 = ~w71 & ~w135;
assign w995 = ~w458 & ~w701;
assign w996 = w61 & w80;
assign w997 = ~w907 & ~w996;
assign w998 = ~w45 & ~w62;
assign w999 = ~w116 & w998;
assign w1000 = ~w113 & ~w123;
assign w1001 = ~w531 & w1000;
assign w1002 = w993 & w994;
assign w1003 = w995 & w997;
assign w1004 = w1002 & w1003;
assign w1005 = w999 & w1001;
assign w1006 = w1004 & w1005;
assign w1007 = ~w75 & ~w776;
assign w1008 = ~w378 & w1007;
assign w1009 = ~w156 & ~w159;
assign w1010 = ~w238 & ~w319;
assign w1011 = ~w67 & ~w279;
assign w1012 = w1010 & w1011;
assign w1013 = w718 & w1012;
assign w1014 = ~w16 & ~w619;
assign w1015 = ~w732 & w1014;
assign w1016 = ~w131 & ~w221;
assign w1017 = ~w652 & w1016;
assign w1018 = ~w178 & ~w649;
assign w1019 = ~w60 & ~w207;
assign w1020 = ~w337 & w1019;
assign w1021 = w96 & w1018;
assign w1022 = w1020 & w1021;
assign w1023 = w1015 & w1017;
assign w1024 = w1022 & w1023;
assign w1025 = ~w392 & ~w789;
assign w1026 = ~w261 & ~w719;
assign w1027 = ~w380 & ~w418;
assign w1028 = ~w190 & ~w252;
assign w1029 = ~w46 & ~w138;
assign w1030 = ~w255 & w1029;
assign w1031 = w755 & w1009;
assign w1032 = w1025 & w1026;
assign w1033 = w1027 & w1028;
assign w1034 = w1032 & w1033;
assign w1035 = w1030 & w1031;
assign w1036 = w1008 & w1035;
assign w1037 = w1013 & w1034;
assign w1038 = w1036 & w1037;
assign w1039 = w1024 & w1038;
assign w1040 = w32 & w66;
assign w1041 = ~w128 & ~w1040;
assign w1042 = ~w388 & ~w538;
assign w1043 = w19 & w79;
assign w1044 = ~w292 & ~w432;
assign w1045 = ~w394 & ~w451;
assign w1046 = ~w167 & ~w180;
assign w1047 = ~w741 & ~w1043;
assign w1048 = w1046 & w1047;
assign w1049 = w1044 & w1045;
assign w1050 = w1048 & w1049;
assign w1051 = w26 & w44;
assign w1052 = ~w400 & ~w1051;
assign w1053 = ~w562 & w1052;
assign w1054 = ~w98 & ~w287;
assign w1055 = ~w88 & ~w118;
assign w1056 = ~w130 & w1055;
assign w1057 = w1041 & w1042;
assign w1058 = w1054 & w1057;
assign w1059 = w985 & w1056;
assign w1060 = w987 & w989;
assign w1061 = w991 & w1053;
assign w1062 = w1060 & w1061;
assign w1063 = w1058 & w1059;
assign w1064 = w1050 & w1063;
assign w1065 = w1006 & w1062;
assign w1066 = w1064 & w1065;
assign w1067 = w983 & w1066;
assign w1068 = w1039 & w1067;
assign w1069 = ~w149 & ~w470;
assign w1070 = ~w131 & w1069;
assign w1071 = ~w322 & ~w432;
assign w1072 = ~w239 & w1071;
assign w1073 = ~w315 & ~w644;
assign w1074 = ~w172 & ~w265;
assign w1075 = ~w81 & ~w406;
assign w1076 = ~w349 & ~w385;
assign w1077 = w9 & w38;
assign w1078 = ~w992 & ~w1077;
assign w1079 = ~w207 & ~w291;
assign w1080 = ~w563 & ~w701;
assign w1081 = ~w319 & ~w396;
assign w1082 = ~w153 & w948;
assign w1083 = ~w157 & w821;
assign w1084 = w1080 & w1081;
assign w1085 = w1083 & w1084;
assign w1086 = w1082 & w1085;
assign w1087 = w379 & ~w623;
assign w1088 = w1073 & w1074;
assign w1089 = w1075 & w1076;
assign w1090 = w1078 & w1079;
assign w1091 = w1089 & w1090;
assign w1092 = w1087 & w1088;
assign w1093 = w64 & w1070;
assign w1094 = w1072 & w1093;
assign w1095 = w1091 & w1092;
assign w1096 = w1094 & w1095;
assign w1097 = w1086 & w1096;
assign w1098 = ~w161 & ~w267;
assign w1099 = w874 & w1098;
assign w1100 = ~w128 & ~w543;
assign w1101 = ~w130 & ~w164;
assign w1102 = ~w118 & ~w213;
assign w1103 = ~w74 & ~w252;
assign w1104 = w32 & w55;
assign w1105 = ~w197 & ~w1104;
assign w1106 = w44 & w184;
assign w1107 = ~w89 & ~w696;
assign w1108 = ~w818 & w1107;
assign w1109 = ~w246 & ~w428;
assign w1110 = w790 & w1109;
assign w1111 = ~w261 & ~w622;
assign w1112 = ~w135 & ~w1043;
assign w1113 = ~w242 & ~w248;
assign w1114 = ~w237 & w1113;
assign w1115 = w1112 & w1114;
assign w1116 = ~w124 & ~w151;
assign w1117 = w19 & w160;
assign w1118 = ~w16 & ~w1117;
assign w1119 = ~w180 & ~w391;
assign w1120 = ~w562 & w1027;
assign w1121 = w1119 & w1120;
assign w1122 = ~w42 & ~w266;
assign w1123 = w32 & w61;
assign w1124 = ~w1040 & ~w1123;
assign w1125 = ~w67 & ~w404;
assign w1126 = ~w540 & ~w580;
assign w1127 = w1125 & w1126;
assign w1128 = ~w278 & ~w447;
assign w1129 = ~w399 & ~w476;
assign w1130 = ~w582 & ~w838;
assign w1131 = w1129 & w1130;
assign w1132 = w346 & w367;
assign w1133 = w840 & w1128;
assign w1134 = w1132 & w1133;
assign w1135 = w1127 & w1131;
assign w1136 = w1134 & w1135;
assign w1137 = ~w316 & ~w363;
assign w1138 = ~w531 & ~w834;
assign w1139 = w1137 & w1138;
assign w1140 = w814 & w1111;
assign w1141 = w1116 & w1118;
assign w1142 = w1122 & w1124;
assign w1143 = w1141 & w1142;
assign w1144 = w1139 & w1140;
assign w1145 = w1108 & w1110;
assign w1146 = w1144 & w1145;
assign w1147 = w1115 & w1143;
assign w1148 = w1121 & w1147;
assign w1149 = w1136 & w1146;
assign w1150 = w1148 & w1149;
assign w1151 = ~w112 & ~w196;
assign w1152 = ~w116 & ~w652;
assign w1153 = ~w123 & ~w356;
assign w1154 = ~w314 & ~w341;
assign w1155 = ~w400 & w1154;
assign w1156 = w1153 & w1155;
assign w1157 = ~w212 & ~w279;
assign w1158 = ~w178 & ~w282;
assign w1159 = w1157 & w1158;
assign w1160 = ~w46 & ~w422;
assign w1161 = ~w431 & w1160;
assign w1162 = w1151 & w1152;
assign w1163 = w1161 & w1162;
assign w1164 = w1159 & w1163;
assign w1165 = w1156 & w1164;
assign w1166 = ~w72 & ~w216;
assign w1167 = ~w339 & ~w944;
assign w1168 = w1166 & w1167;
assign w1169 = ~w18 & ~w251;
assign w1170 = ~w1106 & w1169;
assign w1171 = w950 & w1100;
assign w1172 = w1101 & w1102;
assign w1173 = w1103 & w1105;
assign w1174 = w1172 & w1173;
assign w1175 = w1170 & w1171;
assign w1176 = w1099 & w1168;
assign w1177 = w1175 & w1176;
assign w1178 = w189 & w1174;
assign w1179 = w1177 & w1178;
assign w1180 = w1165 & w1179;
assign w1181 = w1097 & w1180;
assign w1182 = w1150 & w1181;
assign w1183 = ~w1068 & ~w1182;
assign w1184 = w1068 & w1182;
assign w1185 = ~w1183 & ~w1184;
assign w1186 = ~a_26 & w1185;
assign w1187 = (~w1183 & ~w1185) | (~w1183 & w32646) | (~w1185 & w32646);
assign w1188 = w807 & ~w1187;
assign w1189 = ~w807 & w1187;
assign w1190 = ~w1188 & ~w1189;
assign w1191 = ~w153 & ~w420;
assign w1192 = w59 & w122;
assign w1193 = ~w10 & ~w1192;
assign w1194 = ~w315 & ~w337;
assign w1195 = w790 & w1194;
assign w1196 = ~w123 & ~w355;
assign w1197 = w1042 & ~w1117;
assign w1198 = ~w163 & ~w385;
assign w1199 = ~w94 & ~w1043;
assign w1200 = ~w152 & ~w543;
assign w1201 = w1196 & w1200;
assign w1202 = w1198 & w1199;
assign w1203 = w1201 & w1202;
assign w1204 = w1197 & w1203;
assign w1205 = ~w72 & ~w131;
assign w1206 = ~w190 & ~w249;
assign w1207 = ~w112 & ~w243;
assign w1208 = w1206 & w1207;
assign w1209 = ~w18 & ~w708;
assign w1210 = w560 & w1209;
assign w1211 = w1208 & w1210;
assign w1212 = ~w136 & w1205;
assign w1213 = w989 & w1212;
assign w1214 = w1211 & w1213;
assign w1215 = w1191 & w1193;
assign w1216 = w1195 & w1215;
assign w1217 = w1204 & w1216;
assign w1218 = w1214 & w1217;
assign w1219 = ~w39 & ~w339;
assign w1220 = a_23 & ~a_24;
assign w1221 = ~a_23 & a_24;
assign w1222 = ~w1220 & ~w1221;
assign w1223 = a_25 & ~a_26;
assign w1224 = ~a_25 & a_26;
assign w1225 = ~w1223 & ~w1224;
assign w1226 = ~w1222 & ~w1225;
assign w1227 = ~w20 & w1226;
assign w1228 = (w122 & w1227) | (w122 & w32647) | (w1227 & w32647);
assign w1229 = ~w115 & ~w159;
assign w1230 = ~w34 & ~w238;
assign w1231 = ~w248 & ~w644;
assign w1232 = ~w896 & w1231;
assign w1233 = w1229 & w1230;
assign w1234 = w1232 & w1233;
assign w1235 = ~w254 & w670;
assign w1236 = w1234 & w1235;
assign w1237 = ~w95 & w1124;
assign w1238 = ~w380 & ~w694;
assign w1239 = ~w126 & w1238;
assign w1240 = a_28 & w11;
assign w1241 = ~w193 & w1240;
assign w1242 = ~w67 & w364;
assign w1243 = ~w185 & ~w541;
assign w1244 = ~w649 & w1243;
assign w1245 = w744 & w1244;
assign w1246 = w454 & w1072;
assign w1247 = w1242 & w1246;
assign w1248 = w1245 & w1247;
assign w1249 = ~w313 & ~w357;
assign w1250 = ~w292 & ~w878;
assign w1251 = ~w776 & ~w1104;
assign w1252 = ~w1241 & w1249;
assign w1253 = w1250 & w1251;
assign w1254 = w1252 & w1253;
assign w1255 = w1237 & w1239;
assign w1256 = w1254 & w1255;
assign w1257 = w1236 & w1256;
assign w1258 = w1248 & w1257;
assign w1259 = w524 & w32648;
assign w1260 = ~w113 & ~w167;
assign w1261 = ~w392 & ~w645;
assign w1262 = ~w116 & ~w279;
assign w1263 = w1261 & w1262;
assign w1264 = w1260 & w1263;
assign w1265 = ~w71 & ~w572;
assign w1266 = ~w597 & ~w732;
assign w1267 = ~w585 & w1266;
assign w1268 = ~w349 & ~w730;
assign w1269 = ~w62 & ~w147;
assign w1270 = ~w217 & ~w366;
assign w1271 = w1269 & w1270;
assign w1272 = w1268 & w1271;
assign w1273 = ~w422 & ~w741;
assign w1274 = ~w261 & w1128;
assign w1275 = w1265 & w1273;
assign w1276 = w1274 & w1275;
assign w1277 = w1267 & w1276;
assign w1278 = w1272 & w1277;
assign w1279 = ~w389 & ~w698;
assign w1280 = ~w450 & ~w838;
assign w1281 = ~w260 & ~w719;
assign w1282 = ~w395 & w1281;
assign w1283 = ~w220 & w567;
assign w1284 = w758 & w1280;
assign w1285 = w1283 & w1284;
assign w1286 = w1282 & w1285;
assign w1287 = ~w124 & ~w325;
assign w1288 = ~a_26 & w14;
assign w1289 = w47 & w1288;
assign w1290 = w1287 & ~w1289;
assign w1291 = ~w283 & ~w818;
assign w1292 = ~w97 & ~w172;
assign w1293 = ~w60 & ~w314;
assign w1294 = w1292 & w1293;
assign w1295 = ~w213 & ~w391;
assign w1296 = w1291 & w1295;
assign w1297 = w1294 & w1296;
assign w1298 = w1279 & w1290;
assign w1299 = w1297 & w1298;
assign w1300 = w1286 & w1299;
assign w1301 = ~w118 & ~w151;
assign w1302 = ~w710 & w1301;
assign w1303 = w566 & w1302;
assign w1304 = w1264 & w1303;
assign w1305 = w1278 & w1304;
assign w1306 = w1300 & w1305;
assign w1307 = w1258 & w1259;
assign w1308 = w1306 & w1307;
assign w1309 = ~w144 & ~w544;
assign w1310 = ~w281 & ~w365;
assign w1311 = w1309 & w1310;
assign w1312 = ~w76 & ~w251;
assign w1313 = w548 & w1312;
assign w1314 = w575 & w1313;
assign w1315 = w1311 & w1314;
assign w1316 = ~w23 & ~w85;
assign w1317 = ~w252 & ~w475;
assign w1318 = w1316 & w1317;
assign w1319 = w1219 & w1318;
assign w1320 = ~w1228 & w1319;
assign w1321 = w1315 & w1320;
assign w1322 = w1218 & w1321;
assign w1323 = w1308 & w1322;
assign w1324 = (w668 & ~w1308) | (w668 & w32649) | (~w1308 & w32649);
assign w1325 = ~a_31 & ~w28;
assign w1326 = a_31 & ~w35;
assign w1327 = ~w1325 & ~w1326;
assign w1328 = w469 & w32650;
assign w1329 = ~w262 & ~w350;
assign w1330 = ~w400 & ~w696;
assign w1331 = ~w701 & ~w1192;
assign w1332 = ~w394 & ~w589;
assign w1333 = w627 & w1332;
assign w1334 = ~w10 & ~w177;
assign w1335 = w808 & w876;
assign w1336 = w36 & w184;
assign w1337 = ~w83 & ~w170;
assign w1338 = ~w246 & ~w1336;
assign w1339 = w1337 & w1338;
assign w1340 = ~w86 & ~w312;
assign w1341 = w132 & ~w321;
assign w1342 = w1340 & w1341;
assign w1343 = ~w653 & ~w878;
assign w1344 = ~w138 & ~w431;
assign w1345 = ~w737 & w756;
assign w1346 = ~w128 & ~w396;
assign w1347 = w533 & w1346;
assign w1348 = w549 & w788;
assign w1349 = w961 & w1343;
assign w1350 = w1344 & w1349;
assign w1351 = w1347 & w1348;
assign w1352 = w1345 & w1351;
assign w1353 = w1342 & w1350;
assign w1354 = w1352 & w1353;
assign w1355 = ~w190 & ~w1077;
assign w1356 = ~w292 & ~w734;
assign w1357 = ~w136 & ~w221;
assign w1358 = w1355 & w1357;
assign w1359 = w1356 & w1358;
assign w1360 = ~w143 & ~w369;
assign w1361 = ~w406 & ~w647;
assign w1362 = ~w249 & ~w291;
assign w1363 = ~w135 & w381;
assign w1364 = w1334 & w1360;
assign w1365 = w1361 & w1362;
assign w1366 = w1364 & w1365;
assign w1367 = w1333 & w1363;
assign w1368 = w1335 & w1339;
assign w1369 = w1367 & w1368;
assign w1370 = w1359 & w1366;
assign w1371 = w1369 & w1370;
assign w1372 = w1236 & w1371;
assign w1373 = w1354 & w1372;
assign w1374 = ~w459 & ~w815;
assign w1375 = ~w237 & ~w475;
assign w1376 = ~w18 & ~w834;
assign w1377 = ~w183 & ~w720;
assign w1378 = ~w112 & ~w266;
assign w1379 = w1374 & w1378;
assign w1380 = w1375 & w1376;
assign w1381 = w1377 & w1380;
assign w1382 = w1237 & w1379;
assign w1383 = w1381 & w1382;
assign w1384 = ~w146 & ~w315;
assign w1385 = ~w89 & w1384;
assign w1386 = ~w53 & w560;
assign w1387 = w840 & w875;
assign w1388 = w1249 & w1329;
assign w1389 = w1330 & w1331;
assign w1390 = w1388 & w1389;
assign w1391 = w1385 & w1387;
assign w1392 = w1386 & w1391;
assign w1393 = w1328 & w1390;
assign w1394 = w1392 & w1393;
assign w1395 = w1383 & w1394;
assign w1396 = w1248 & w1395;
assign w1397 = w1373 & w1396;
assign w1398 = w1327 & ~w1397;
assign w1399 = a_31 & w28;
assign w1400 = ~w134 & ~w710;
assign w1401 = ~w186 & ~w458;
assign w1402 = w114 & ~w696;
assign w1403 = w1279 & w1402;
assign w1404 = w1401 & w1403;
assign w1405 = ~w213 & ~w363;
assign w1406 = ~w65 & ~w396;
assign w1407 = w1405 & w1406;
assign w1408 = ~w216 & w1407;
assign w1409 = ~w10 & ~w459;
assign w1410 = ~w701 & w1409;
assign w1411 = w876 & w1410;
assign w1412 = ~w68 & ~w279;
assign w1413 = ~w446 & ~w562;
assign w1414 = ~w208 & ~w719;
assign w1415 = w1412 & w1414;
assign w1416 = w1413 & w1415;
assign w1417 = w793 & w1416;
assign w1418 = ~w362 & ~w818;
assign w1419 = ~w88 & ~w350;
assign w1420 = w560 & w627;
assign w1421 = ~w260 & ~w473;
assign w1422 = ~w541 & ~w714;
assign w1423 = ~w181 & ~w395;
assign w1424 = ~w116 & ~w249;
assign w1425 = ~w404 & ~w563;
assign w1426 = ~w653 & w1425;
assign w1427 = w1422 & w1423;
assign w1428 = w1424 & w1427;
assign w1429 = w1426 & w1428;
assign w1430 = ~w167 & ~w214;
assign w1431 = ~w86 & ~w196;
assign w1432 = w247 & w1430;
assign w1433 = w1431 & w1432;
assign w1434 = w1429 & w1433;
assign w1435 = ~w392 & ~w593;
assign w1436 = ~w322 & ~w838;
assign w1437 = ~w146 & ~w671;
assign w1438 = w561 & w1437;
assign w1439 = w1435 & w1436;
assign w1440 = w1438 & w1439;
assign w1441 = ~w67 & ~w135;
assign w1442 = ~w645 & w1441;
assign w1443 = w648 & w836;
assign w1444 = w1418 & w1419;
assign w1445 = w1421 & w1444;
assign w1446 = w1442 & w1443;
assign w1447 = w1420 & w1446;
assign w1448 = w457 & w1445;
assign w1449 = w1440 & w1448;
assign w1450 = w1447 & w1449;
assign w1451 = w1434 & w1450;
assign w1452 = ~w118 & ~w239;
assign w1453 = ~w151 & w1452;
assign w1454 = ~w18 & ~w97;
assign w1455 = ~w180 & w433;
assign w1456 = ~w60 & w744;
assign w1457 = w1454 & w1456;
assign w1458 = w1453 & w1455;
assign w1459 = w1457 & w1458;
assign w1460 = w1408 & w1411;
assign w1461 = w1459 & w1460;
assign w1462 = w1404 & w1417;
assign w1463 = w1461 & w1462;
assign w1464 = ~w173 & ~w368;
assign w1465 = ~w267 & w1464;
assign w1466 = w840 & ~w1104;
assign w1467 = w539 & w584;
assign w1468 = w1287 & w1400;
assign w1469 = w1467 & w1468;
assign w1470 = w52 & w1465;
assign w1471 = w1466 & w1470;
assign w1472 = w1469 & w1471;
assign w1473 = w537 & w1204;
assign w1474 = w1472 & w1473;
assign w1475 = w1451 & w32651;
assign w1476 = w1399 & ~w1475;
assign w1477 = ~w8 & ~w11;
assign w1478 = a_31 & ~w1477;
assign w1479 = ~w1397 & ~w1475;
assign w1480 = ~w321 & ~w356;
assign w1481 = ~w153 & ~w190;
assign w1482 = ~w138 & ~w708;
assign w1483 = ~w177 & ~w181;
assign w1484 = w1480 & w1483;
assign w1485 = w1481 & w1482;
assign w1486 = w1484 & w1485;
assign w1487 = ~w94 & ~w205;
assign w1488 = ~w127 & ~w147;
assign w1489 = ~w221 & ~w366;
assign w1490 = ~w65 & ~w291;
assign w1491 = ~w316 & ~w404;
assign w1492 = ~w136 & ~w245;
assign w1493 = ~w312 & ~w349;
assign w1494 = ~w71 & ~w124;
assign w1495 = ~w217 & w1494;
assign w1496 = ~w447 & ~w701;
assign w1497 = ~w896 & w1496;
assign w1498 = ~w266 & ~w463;
assign w1499 = w1054 & w1498;
assign w1500 = w1250 & w1493;
assign w1501 = w1499 & w1500;
assign w1502 = w1495 & w1497;
assign w1503 = w1501 & w1502;
assign w1504 = ~w385 & ~w696;
assign w1505 = ~w350 & ~w422;
assign w1506 = ~w88 & ~w325;
assign w1507 = ~w420 & w1506;
assign w1508 = w1505 & w1507;
assign w1509 = ~w396 & ~w406;
assign w1510 = w1377 & w1509;
assign w1511 = w1384 & w1487;
assign w1512 = w1488 & w1489;
assign w1513 = w1490 & w1491;
assign w1514 = w1492 & w1504;
assign w1515 = w1513 & w1514;
assign w1516 = w1511 & w1512;
assign w1517 = w1466 & w1510;
assign w1518 = w1516 & w1517;
assign w1519 = w1486 & w1515;
assign w1520 = w1508 & w1519;
assign w1521 = w1503 & w1518;
assign w1522 = w1520 & w1521;
assign w1523 = w643 & w1522;
assign w1524 = ~w126 & ~w196;
assign w1525 = ~w34 & w1524;
assign w1526 = w1208 & w1525;
assign w1527 = ~w115 & ~w221;
assign w1528 = ~w261 & ~w459;
assign w1529 = w1527 & w1528;
assign w1530 = w628 & w1491;
assign w1531 = w1529 & w1530;
assign w1532 = w1309 & w31562;
assign w1533 = ~w85 & ~w337;
assign w1534 = ~w282 & ~w568;
assign w1535 = w1533 & w1534;
assign w1536 = ~w50 & ~w992;
assign w1537 = ~w446 & w1536;
assign w1538 = ~w75 & ~w157;
assign w1539 = ~w292 & w1538;
assign w1540 = w1537 & w1539;
assign w1541 = ~w645 & ~w737;
assign w1542 = ~w125 & w1541;
assign w1543 = ~w166 & ~w694;
assign w1544 = ~w128 & ~w323;
assign w1545 = ~w649 & ~w832;
assign w1546 = w1544 & w1545;
assign w1547 = w1045 & w1543;
assign w1548 = w1546 & w1547;
assign w1549 = w1542 & w1548;
assign w1550 = ~w149 & ~w418;
assign w1551 = ~w183 & ~w776;
assign w1552 = ~w46 & ~w97;
assign w1553 = ~w118 & ~w463;
assign w1554 = w1552 & w1553;
assign w1555 = w215 & w1550;
assign w1556 = w1551 & w1555;
assign w1557 = w1535 & w1554;
assign w1558 = w1556 & w1557;
assign w1559 = w1532 & w1540;
assign w1560 = w1558 & w1559;
assign w1561 = w1549 & w1560;
assign w1562 = ~w56 & ~w287;
assign w1563 = ~w10 & ~w68;
assign w1564 = ~w237 & ~w470;
assign w1565 = ~w589 & w1564;
assign w1566 = w1563 & w1565;
assign w1567 = ~w325 & ~w458;
assign w1568 = ~w153 & ~w345;
assign w1569 = ~w429 & w1568;
assign w1570 = w1567 & w1569;
assign w1571 = ~w146 & ~w403;
assign w1572 = ~w278 & ~w583;
assign w1573 = ~w167 & ~w896;
assign w1574 = w63 & w1573;
assign w1575 = w141 & w360;
assign w1576 = w1343 & w1562;
assign w1577 = w1571 & w1572;
assign w1578 = w1576 & w1577;
assign w1579 = w1574 & w1575;
assign w1580 = w1578 & w1579;
assign w1581 = w1566 & w1570;
assign w1582 = w1580 & w1581;
assign w1583 = ~w177 & ~w593;
assign w1584 = ~w350 & ~w543;
assign w1585 = ~w388 & ~w815;
assign w1586 = ~w547 & w1360;
assign w1587 = w1585 & w1586;
assign w1588 = ~w291 & ~w626;
assign w1589 = ~w281 & w397;
assign w1590 = w1588 & w1589;
assign w1591 = w1587 & w1590;
assign w1592 = ~w123 & ~w178;
assign w1593 = ~w313 & ~w1104;
assign w1594 = w1592 & w1593;
assign w1595 = w353 & w1583;
assign w1596 = w1584 & w1595;
assign w1597 = w837 & w1594;
assign w1598 = w1596 & w1597;
assign w1599 = w1591 & w1598;
assign w1600 = ~w197 & ~w218;
assign w1601 = ~w239 & w1600;
assign w1602 = w1600 & w31563;
assign w1603 = ~w23 & w542;
assign w1604 = ~w391 & ~w741;
assign w1605 = ~w152 & ~w473;
assign w1606 = ~w907 & w1605;
assign w1607 = ~w172 & ~w572;
assign w1608 = ~w314 & ~w389;
assign w1609 = ~w395 & ~w652;
assign w1610 = w1608 & w1609;
assign w1611 = w338 & w1607;
assign w1612 = w1610 & w1611;
assign w1613 = w1606 & w1612;
assign w1614 = ~w136 & ~w644;
assign w1615 = ~w65 & ~w142;
assign w1616 = ~w195 & ~w730;
assign w1617 = w605 & w1616;
assign w1618 = w835 & w1604;
assign w1619 = w1614 & w1615;
assign w1620 = w1618 & w1619;
assign w1621 = w1603 & w1617;
assign w1622 = w1620 & w1621;
assign w1623 = w1526 & w1531;
assign w1624 = w1602 & w1623;
assign w1625 = w1613 & w1622;
assign w1626 = w1624 & w1625;
assign w1627 = w1582 & w1599;
assign w1628 = w1626 & w1627;
assign w1629 = w1561 & w1628;
assign w1630 = ~w1523 & ~w1629;
assign w1631 = ~w238 & ~w399;
assign w1632 = ~w153 & ~w543;
assign w1633 = ~w72 & ~w86;
assign w1634 = ~w131 & ~w392;
assign w1635 = w1631 & w1634;
assign w1636 = w1632 & w1633;
assign w1637 = w1635 & w1636;
assign w1638 = ~w365 & ~w559;
assign w1639 = ~w315 & ~w720;
assign w1640 = ~w205 & ~w260;
assign w1641 = ~w319 & ~w1123;
assign w1642 = ~w62 & w198;
assign w1643 = ~w95 & ~w531;
assign w1644 = ~w309 & ~w363;
assign w1645 = ~w156 & ~w212;
assign w1646 = ~w208 & ~w217;
assign w1647 = ~w838 & w1646;
assign w1648 = w755 & w871;
assign w1649 = w1638 & w1639;
assign w1650 = w1640 & w1641;
assign w1651 = w1643 & w1644;
assign w1652 = w1645 & w1651;
assign w1653 = w1649 & w1650;
assign w1654 = w1647 & w1648;
assign w1655 = w1642 & w1654;
assign w1656 = w1652 & w1653;
assign w1657 = w1655 & w1656;
assign w1658 = ~w151 & ~w393;
assign w1659 = ~w248 & w1658;
assign w1660 = ~w341 & w1615;
assign w1661 = ~w290 & ~w406;
assign w1662 = ~w279 & ~w388;
assign w1663 = ~w314 & ~w423;
assign w1664 = ~w267 & w620;
assign w1665 = ~w18 & ~w98;
assign w1666 = ~w88 & ~w169;
assign w1667 = ~w647 & w1666;
assign w1668 = w57 & w673;
assign w1669 = w813 & w1101;
assign w1670 = w1661 & w1662;
assign w1671 = w1663 & w1665;
assign w1672 = w1670 & w1671;
assign w1673 = w1668 & w1669;
assign w1674 = w1659 & w1667;
assign w1675 = w1660 & w1664;
assign w1676 = w1674 & w1675;
assign w1677 = w1672 & w1673;
assign w1678 = w1676 & w1677;
assign w1679 = ~w124 & ~w339;
assign w1680 = ~w428 & ~w622;
assign w1681 = ~w243 & ~w422;
assign w1682 = ~w626 & w1681;
assign w1683 = ~w256 & w986;
assign w1684 = w1682 & w1683;
assign w1685 = ~w94 & ~w283;
assign w1686 = ~w161 & ~w585;
assign w1687 = ~w68 & ~w895;
assign w1688 = ~w590 & w628;
assign w1689 = ~w562 & ~w583;
assign w1690 = ~w191 & ~w652;
assign w1691 = ~w278 & ~w362;
assign w1692 = ~w74 & ~w431;
assign w1693 = ~w355 & ~w589;
assign w1694 = ~w16 & ~w475;
assign w1695 = ~w404 & ~w623;
assign w1696 = w1691 & w1695;
assign w1697 = w1692 & w1693;
assign w1698 = w1694 & w1697;
assign w1699 = w354 & w1696;
assign w1700 = w1698 & w1699;
assign w1701 = ~w143 & w1028;
assign w1702 = w1679 & w1680;
assign w1703 = w1685 & w1686;
assign w1704 = w1687 & w1689;
assign w1705 = w1690 & w1704;
assign w1706 = w1702 & w1703;
assign w1707 = w1688 & w1701;
assign w1708 = w1706 & w1707;
assign w1709 = w1637 & w1705;
assign w1710 = w1684 & w1709;
assign w1711 = w1700 & w1708;
assign w1712 = w1710 & w1711;
assign w1713 = w1657 & w1678;
assign w1714 = w1712 & w1713;
assign w1715 = w1561 & w1714;
assign w1716 = w1266 & w1643;
assign w1717 = ~w538 & w1260;
assign w1718 = ~w169 & ~w540;
assign w1719 = ~w130 & ~w431;
assign w1720 = ~w245 & ~w1043;
assign w1721 = ~w153 & ~w339;
assign w1722 = ~w252 & ~w450;
assign w1723 = ~w316 & w1721;
assign w1724 = w1722 & w1723;
assign w1725 = ~w254 & ~w671;
assign w1726 = ~w468 & ~w568;
assign w1727 = ~w74 & ~w177;
assign w1728 = w1726 & w1727;
assign w1729 = ~w321 & ~w341;
assign w1730 = ~w352 & ~w563;
assign w1731 = ~w834 & w1730;
assign w1732 = w1725 & w1729;
assign w1733 = w1731 & w1732;
assign w1734 = w187 & w1728;
assign w1735 = w1733 & w1734;
assign w1736 = ~w541 & ~w734;
assign w1737 = ~w45 & ~w789;
assign w1738 = ~w476 & ~w585;
assign w1739 = ~w30 & ~w264;
assign w1740 = ~w292 & w1739;
assign w1741 = ~w205 & ~w248;
assign w1742 = ~w362 & ~w399;
assign w1743 = ~w907 & w1742;
assign w1744 = w1718 & w1741;
assign w1745 = w1719 & w1720;
assign w1746 = w1736 & w1737;
assign w1747 = w1738 & w1746;
assign w1748 = w1744 & w1745;
assign w1749 = w1740 & w1743;
assign w1750 = w1748 & w1749;
assign w1751 = w1724 & w1747;
assign w1752 = w1750 & w1751;
assign w1753 = w1735 & w1752;
assign w1754 = ~w404 & ~w626;
assign w1755 = ~w142 & ~w261;
assign w1756 = ~w140 & ~w357;
assign w1757 = ~w152 & ~w190;
assign w1758 = ~w400 & ~w710;
assign w1759 = ~w123 & w280;
assign w1760 = w1757 & w1758;
assign w1761 = w1759 & w1760;
assign w1762 = ~w206 & w1261;
assign w1763 = w1261 & w32652;
assign w1764 = ~w214 & ~w365;
assign w1765 = ~w173 & ~w473;
assign w1766 = ~w423 & ~w1117;
assign w1767 = w1764 & w1766;
assign w1768 = w1765 & w1767;
assign w1769 = ~w323 & ~w428;
assign w1770 = ~w164 & ~w197;
assign w1771 = ~w194 & w1770;
assign w1772 = ~w309 & ~w380;
assign w1773 = w673 & w1772;
assign w1774 = ~w112 & ~w644;
assign w1775 = ~w1077 & w1774;
assign w1776 = ~w172 & ~w378;
assign w1777 = ~w1104 & ~w1192;
assign w1778 = ~w366 & ~w878;
assign w1779 = w1122 & w1777;
assign w1780 = w1778 & w1779;
assign w1781 = ~w136 & ~w212;
assign w1782 = ~w23 & ~w76;
assign w1783 = ~w345 & w1782;
assign w1784 = w90 & w129;
assign w1785 = w289 & w1769;
assign w1786 = w1776 & w1781;
assign w1787 = w1785 & w1786;
assign w1788 = w1783 & w1784;
assign w1789 = w1282 & w1771;
assign w1790 = w1773 & w1775;
assign w1791 = w1789 & w1790;
assign w1792 = w1787 & w1788;
assign w1793 = w1780 & w1792;
assign w1794 = w1791 & w1793;
assign w1795 = ~w238 & ~w944;
assign w1796 = w145 & w1795;
assign w1797 = w1505 & w1754;
assign w1798 = w1755 & w1756;
assign w1799 = w1797 & w1798;
assign w1800 = w1716 & w1796;
assign w1801 = w1717 & w1800;
assign w1802 = w1761 & w1799;
assign w1803 = w1763 & w1768;
assign w1804 = w1802 & w1803;
assign w1805 = w706 & w1801;
assign w1806 = w1804 & w1805;
assign w1807 = w1753 & w1806;
assign w1808 = w1794 & w1807;
assign w1809 = w1715 & w1808;
assign w1810 = ~w149 & ~w459;
assign w1811 = ~w369 & ~w446;
assign w1812 = w1810 & w1811;
assign w1813 = ~w18 & ~w188;
assign w1814 = ~w177 & ~w896;
assign w1815 = ~w385 & ~w698;
assign w1816 = ~w400 & w602;
assign w1817 = w1400 & w1815;
assign w1818 = w1816 & w1817;
assign w1819 = ~w283 & ~w541;
assign w1820 = ~w181 & ~w292;
assign w1821 = ~w42 & ~w389;
assign w1822 = ~w195 & ~w342;
assign w1823 = ~w46 & ~w221;
assign w1824 = ~w216 & ~w544;
assign w1825 = w1823 & w1824;
assign w1826 = ~w135 & ~w173;
assign w1827 = w947 & w1826;
assign w1828 = w1819 & w1820;
assign w1829 = w1821 & w1822;
assign w1830 = w1828 & w1829;
assign w1831 = w1825 & w1827;
assign w1832 = w1830 & w1831;
assign w1833 = ~w53 & ~w345;
assign w1834 = ~w597 & ~w1104;
assign w1835 = w1833 & w1834;
assign w1836 = ~w363 & ~w996;
assign w1837 = w340 & w1836;
assign w1838 = w855 & w1260;
assign w1839 = w1533 & w1813;
assign w1840 = w1814 & w1839;
assign w1841 = w1837 & w1838;
assign w1842 = w999 & w1812;
assign w1843 = w1835 & w1842;
assign w1844 = w1840 & w1841;
assign w1845 = w1818 & w1844;
assign w1846 = w1832 & w1843;
assign w1847 = w1845 & w1846;
assign w1848 = ~w312 & ~w531;
assign w1849 = ~w147 & w317;
assign w1850 = ~w130 & ~w322;
assign w1851 = ~w140 & ~w671;
assign w1852 = w1850 & w1851;
assign w1853 = ~w75 & ~w458;
assign w1854 = ~w281 & ~w653;
assign w1855 = ~w196 & ~w314;
assign w1856 = ~w95 & w790;
assign w1857 = w1853 & w1854;
assign w1858 = w1855 & w1857;
assign w1859 = w1856 & w1858;
assign w1860 = ~w67 & ~w217;
assign w1861 = ~w278 & ~w719;
assign w1862 = ~w572 & ~w730;
assign w1863 = w1107 & w1862;
assign w1864 = w1333 & w1863;
assign w1865 = ~w593 & w1287;
assign w1866 = ~w243 & ~w393;
assign w1867 = w1865 & w1866;
assign w1868 = ~w350 & ~w1117;
assign w1869 = w289 & w1868;
assign w1870 = ~w112 & ~w734;
assign w1871 = ~w142 & ~w206;
assign w1872 = ~w97 & ~w720;
assign w1873 = ~w357 & ~w399;
assign w1874 = ~w451 & w839;
assign w1875 = w946 & w1111;
assign w1876 = w1662 & w1686;
assign w1877 = w1860 & w1861;
assign w1878 = w1870 & w1871;
assign w1879 = w1872 & w1873;
assign w1880 = w1878 & w1879;
assign w1881 = w1876 & w1877;
assign w1882 = w1874 & w1875;
assign w1883 = w1869 & w1882;
assign w1884 = w1880 & w1881;
assign w1885 = w1864 & w1867;
assign w1886 = w1884 & w1885;
assign w1887 = w1883 & w1886;
assign w1888 = ~w123 & ~w530;
assign w1889 = ~w714 & w1888;
assign w1890 = ~w266 & ~w418;
assign w1891 = w80 & w32653;
assign w1892 = ~w68 & ~w172;
assign w1893 = ~w220 & w1892;
assign w1894 = ~w391 & ~w645;
assign w1895 = ~w431 & ~w818;
assign w1896 = ~w267 & ~w362;
assign w1897 = w84 & w1896;
assign w1898 = w571 & w754;
assign w1899 = w1894 & w1895;
assign w1900 = w1898 & w1899;
assign w1901 = w1893 & w1897;
assign w1902 = w1900 & w1901;
assign w1903 = ~w180 & w1536;
assign w1904 = w1781 & w1848;
assign w1905 = w1890 & ~w1891;
assign w1906 = w1904 & w1905;
assign w1907 = w1849 & w1903;
assign w1908 = w1852 & w1889;
assign w1909 = w1907 & w1908;
assign w1910 = w1906 & w1909;
assign w1911 = w1859 & w1902;
assign w1912 = w1910 & w1911;
assign w1913 = w1847 & w1912;
assign w1914 = w1887 & w1913;
assign w1915 = ~w1715 & ~w1914;
assign w1916 = w1715 & w1914;
assign w1917 = ~w1915 & ~w1916;
assign w1918 = ~w458 & ~w815;
assign w1919 = ~w245 & ~w563;
assign w1920 = ~w34 & ~w694;
assign w1921 = ~w217 & ~w323;
assign w1922 = ~w94 & ~w146;
assign w1923 = ~w214 & ~w287;
assign w1924 = ~w362 & w1923;
assign w1925 = w713 & w1922;
assign w1926 = w1921 & w1925;
assign w1927 = w1924 & w1926;
assign w1928 = ~w186 & ~w380;
assign w1929 = ~w95 & ~w161;
assign w1930 = w1765 & w1929;
assign w1931 = ~w118 & ~w818;
assign w1932 = ~w147 & w680;
assign w1933 = w773 & w1280;
assign w1934 = w1918 & w1919;
assign w1935 = w1920 & w1931;
assign w1936 = w1934 & w1935;
assign w1937 = w1932 & w1933;
assign w1938 = w1928 & w1930;
assign w1939 = w1937 & w1938;
assign w1940 = w1936 & w1939;
assign w1941 = w1927 & w1940;
assign w1942 = ~w282 & ~w395;
assign w1943 = ~w76 & ~w583;
assign w1944 = ~w645 & w1943;
assign w1945 = w1010 & w1942;
assign w1946 = w1944 & w1945;
assign w1947 = ~w349 & ~w623;
assign w1948 = ~w113 & ~w730;
assign w1949 = ~w39 & ~w291;
assign w1950 = ~w288 & ~w292;
assign w1951 = ~w243 & ~w388;
assign w1952 = a_25 & w5;
assign w1953 = w36 & w1952;
assign w1954 = ~w23 & ~w585;
assign w1955 = ~w378 & ~w1953;
assign w1956 = w958 & w1955;
assign w1957 = w1848 & w1951;
assign w1958 = w1954 & w1957;
assign w1959 = w1956 & w1958;
assign w1960 = ~w696 & ~w1077;
assign w1961 = ~w221 & ~w429;
assign w1962 = ~w619 & w1961;
assign w1963 = w1960 & w1962;
assign w1964 = a_23 & w14;
assign w1965 = w47 & w1964;
assign w1966 = ~w188 & ~w475;
assign w1967 = ~w400 & ~w1043;
assign w1968 = ~w698 & w1967;
assign w1969 = ~w342 & ~w468;
assign w1970 = ~w256 & ~w447;
assign w1971 = ~w541 & w1970;
assign w1972 = w1969 & w1971;
assign w1973 = w1968 & w1972;
assign w1974 = ~w597 & ~w714;
assign w1975 = ~w18 & ~w459;
assign w1976 = ~w719 & ~w870;
assign w1977 = ~w1965 & w1976;
assign w1978 = w168 & w1975;
assign w1979 = w1480 & w1633;
assign w1980 = w1966 & w1974;
assign w1981 = w1979 & w1980;
assign w1982 = w1977 & w1978;
assign w1983 = w1981 & w1982;
assign w1984 = w1963 & w1983;
assign w1985 = w1973 & w1984;
assign w1986 = ~w1123 & w1687;
assign w1987 = ~w157 & ~w368;
assign w1988 = ~w363 & ~w463;
assign w1989 = ~w74 & ~w776;
assign w1990 = ~w404 & ~w944;
assign w1991 = w1989 & w1990;
assign w1992 = w677 & w1309;
assign w1993 = w1583 & w1693;
assign w1994 = w1947 & w1948;
assign w1995 = w1949 & w1950;
assign w1996 = w1987 & w1988;
assign w1997 = w1995 & w1996;
assign w1998 = w1993 & w1994;
assign w1999 = w1986 & w1992;
assign w2000 = w1991 & w1999;
assign w2001 = w1997 & w1998;
assign w2002 = w1946 & w2001;
assign w2003 = w1959 & w2000;
assign w2004 = w2002 & w2003;
assign w2005 = w1941 & w2004;
assign w2006 = w1985 & w2005;
assign w2007 = w1914 & w2006;
assign w2008 = ~w282 & ~w698;
assign w2009 = ~w530 & w2008;
assign w2010 = ~w261 & ~w671;
assign w2011 = ~w776 & w2010;
assign w2012 = ~w128 & ~w279;
assign w2013 = w1419 & w2012;
assign w2014 = ~w173 & ~w432;
assign w2015 = ~w563 & w935;
assign w2016 = ~w169 & ~w291;
assign w2017 = ~w392 & ~w1077;
assign w2018 = w2016 & w2017;
assign w2019 = ~w163 & ~w183;
assign w2020 = ~w42 & w1758;
assign w2021 = w1642 & w2019;
assign w2022 = w2020 & w2021;
assign w2023 = ~w283 & w346;
assign w2024 = w1633 & w2014;
assign w2025 = w2023 & w2024;
assign w2026 = w679 & w2009;
assign w2027 = w2011 & w2013;
assign w2028 = w2015 & w2018;
assign w2029 = w2027 & w2028;
assign w2030 = w2025 & w2026;
assign w2031 = w2029 & w2030;
assign w2032 = w2022 & w2031;
assign w2033 = ~w94 & ~w130;
assign w2034 = ~w23 & ~w429;
assign w2035 = ~w125 & ~w815;
assign w2036 = ~w394 & ~w720;
assign w2037 = ~w789 & w1607;
assign w2038 = ~w188 & w650;
assign w2039 = w1894 & w2033;
assign w2040 = w2034 & w2035;
assign w2041 = w2036 & w2040;
assign w2042 = w2038 & w2039;
assign w2043 = w2037 & w2042;
assign w2044 = w2041 & w2043;
assign w2045 = ~w208 & ~w447;
assign w2046 = ~w459 & w2045;
assign w2047 = ~w134 & ~w339;
assign w2048 = ~w732 & w2047;
assign w2049 = w122 & w868;
assign w2050 = ~w341 & ~w559;
assign w2051 = ~w2049 & w2050;
assign w2052 = ~w399 & ~w1043;
assign w2053 = ~w406 & w2052;
assign w2054 = ~w39 & ~w363;
assign w2055 = w693 & w2054;
assign w2056 = w1931 & w2055;
assign w2057 = ~w288 & ~w580;
assign w2058 = ~w719 & w2057;
assign w2059 = ~w319 & ~w538;
assign w2060 = w1193 & w2059;
assign w2061 = w1692 & w2060;
assign w2062 = w2058 & w2061;
assign w2063 = ~w265 & ~w895;
assign w2064 = ~w89 & ~w144;
assign w2065 = w587 & w2064;
assign w2066 = w2063 & w2065;
assign w2067 = w2046 & w2048;
assign w2068 = w2051 & w2053;
assign w2069 = w2067 & w2068;
assign w2070 = w2056 & w2066;
assign w2071 = w2069 & w2070;
assign w2072 = w2062 & w2071;
assign w2073 = w2044 & w2072;
assign w2074 = w894 & w2073;
assign w2075 = w2073 & w32654;
assign w2076 = ~w260 & ~w315;
assign w2077 = ~w647 & w2076;
assign w2078 = ~w127 & ~w544;
assign w2079 = ~w46 & w681;
assign w2080 = w2078 & w2079;
assign w2081 = w2077 & w2080;
assign w2082 = ~w252 & ~w267;
assign w2083 = ~w380 & ~w1965;
assign w2084 = w257 & w778;
assign w2085 = w853 & w2084;
assign w2086 = w317 & w1533;
assign w2087 = ~w645 & ~w996;
assign w2088 = ~w18 & ~w288;
assign w2089 = ~w71 & ~w143;
assign w2090 = ~w75 & ~w251;
assign w2091 = ~w325 & w2090;
assign w2092 = w460 & w2091;
assign w2093 = ~w734 & ~w1117;
assign w2094 = ~w580 & ~w818;
assign w2095 = ~w167 & ~w313;
assign w2096 = ~w352 & w2095;
assign w2097 = ~w34 & ~w262;
assign w2098 = w2094 & w2097;
assign w2099 = w2096 & w2098;
assign w2100 = ~w357 & ~w365;
assign w2101 = ~w547 & ~w1051;
assign w2102 = ~w213 & ~w254;
assign w2103 = ~w186 & ~w585;
assign w2104 = w867 & w2100;
assign w2105 = w2101 & w2102;
assign w2106 = w2104 & w2105;
assign w2107 = w2103 & w2106;
assign w2108 = ~w206 & w938;
assign w2109 = w1219 & w1644;
assign w2110 = w2087 & w2088;
assign w2111 = w2089 & w2093;
assign w2112 = w2110 & w2111;
assign w2113 = w2108 & w2109;
assign w2114 = w2086 & w2113;
assign w2115 = w2092 & w2112;
assign w2116 = w2099 & w2115;
assign w2117 = w2107 & w2114;
assign w2118 = w2116 & w2117;
assign w2119 = ~w218 & ~w694;
assign w2120 = ~w242 & w2119;
assign w2121 = ~w131 & ~w741;
assign w2122 = ~w159 & ~w389;
assign w2123 = ~w834 & w939;
assign w2124 = w939 & w32655;
assign w2125 = ~w45 & ~w81;
assign w2126 = ~w126 & ~w1104;
assign w2127 = w2125 & w2126;
assign w2128 = w240 & w2121;
assign w2129 = w2122 & w2128;
assign w2130 = w2120 & w2127;
assign w2131 = w2129 & w2130;
assign w2132 = w2124 & w2131;
assign w2133 = w137 & ~w345;
assign w2134 = w40 & w1288;
assign w2135 = w584 & ~w2134;
assign w2136 = ~w142 & ~w281;
assign w2137 = ~w714 & w2136;
assign w2138 = w857 & w2082;
assign w2139 = w2083 & w2138;
assign w2140 = w910 & w2137;
assign w2141 = w2133 & w2135;
assign w2142 = w2140 & w2141;
assign w2143 = w2085 & w2139;
assign w2144 = w2142 & w2143;
assign w2145 = w2081 & w2144;
assign w2146 = w2132 & w2145;
assign w2147 = w2032 & w2118;
assign w2148 = w2146 & w2147;
assign w2149 = ~w2075 & ~w2148;
assign w2150 = ~w72 & ~w323;
assign w2151 = ~w267 & ~w698;
assign w2152 = ~w256 & ~w547;
assign w2153 = ~w350 & ~w368;
assign w2154 = ~w562 & ~w626;
assign w2155 = ~w992 & ~w1192;
assign w2156 = w945 & w2155;
assign w2157 = w2154 & w2156;
assign w2158 = w2048 & w2157;
assign w2159 = ~w737 & ~w878;
assign w2160 = ~w42 & w2159;
assign w2161 = ~w264 & ~w380;
assign w2162 = ~w450 & w2161;
assign w2163 = w755 & w808;
assign w2164 = ~w255 & w646;
assign w2165 = ~w39 & w1152;
assign w2166 = w1737 & w1873;
assign w2167 = w2150 & w2151;
assign w2168 = w2152 & w2153;
assign w2169 = w2167 & w2168;
assign w2170 = w2165 & w2166;
assign w2171 = w2160 & w2162;
assign w2172 = w2163 & w2164;
assign w2173 = w2171 & w2172;
assign w2174 = w2169 & w2170;
assign w2175 = w2173 & w2174;
assign w2176 = w2158 & w2175;
assign w2177 = ~w126 & ~w316;
assign w2178 = ~w418 & w672;
assign w2179 = ~w10 & ~w694;
assign w2180 = w2177 & w2179;
assign w2181 = w2178 & w2180;
assign w2182 = ~w161 & ~w422;
assign w2183 = ~w159 & ~w178;
assign w2184 = ~w60 & ~w205;
assign w2185 = ~w83 & ~w363;
assign w2186 = w2182 & w2183;
assign w2187 = w2184 & w2185;
assign w2188 = w2186 & w2187;
assign w2189 = ~w118 & ~w647;
assign w2190 = ~w432 & w1823;
assign w2191 = ~w183 & ~w459;
assign w2192 = ~w313 & ~w530;
assign w2193 = ~w321 & ~w818;
assign w2194 = ~w146 & ~w163;
assign w2195 = ~w153 & ~w342;
assign w2196 = ~w389 & ~w701;
assign w2197 = w2195 & w2196;
assign w2198 = w2192 & w2193;
assign w2199 = w2194 & w2198;
assign w2200 = w2197 & w2199;
assign w2201 = ~w62 & ~w212;
assign w2202 = ~w291 & w2201;
assign w2203 = w158 & w2202;
assign w2204 = ~w86 & ~w541;
assign w2205 = ~w996 & w2204;
assign w2206 = w876 & w1643;
assign w2207 = w1764 & w2189;
assign w2208 = w2191 & w2207;
assign w2209 = w2205 & w2206;
assign w2210 = w1893 & w2190;
assign w2211 = w2209 & w2210;
assign w2212 = w2203 & w2208;
assign w2213 = w2211 & w2212;
assign w2214 = w2200 & w2213;
assign w2215 = w2213 & w32656;
assign w2216 = ~w262 & ~w315;
assign w2217 = ~w128 & w2216;
assign w2218 = w137 & w728;
assign w2219 = ~w151 & ~w1117;
assign w2220 = ~w237 & ~w572;
assign w2221 = ~w1051 & w2220;
assign w2222 = w171 & w792;
assign w2223 = w2219 & w2222;
assign w2224 = w2221 & w2223;
assign w2225 = ~w85 & ~w261;
assign w2226 = ~w378 & w2225;
assign w2227 = w182 & w2035;
assign w2228 = w2226 & w2227;
assign w2229 = w621 & w2217;
assign w2230 = w2218 & w2229;
assign w2231 = w2181 & w2228;
assign w2232 = w2188 & w2231;
assign w2233 = w2224 & w2230;
assign w2234 = w2232 & w2233;
assign w2235 = w2176 & w2234;
assign w2236 = w2215 & w2235;
assign w2237 = ~w2148 & ~w2236;
assign w2238 = ~w2149 & ~w2237;
assign w2239 = ~w60 & ~w355;
assign w2240 = ~w131 & ~w406;
assign w2241 = ~w166 & ~w313;
assign w2242 = ~w585 & w2241;
assign w2243 = ~w85 & ~w389;
assign w2244 = w2239 & w2243;
assign w2245 = w2240 & w2244;
assign w2246 = w2242 & w2245;
assign w2247 = ~w213 & ~w366;
assign w2248 = ~w10 & ~w278;
assign w2249 = ~w543 & ~w701;
assign w2250 = ~w369 & ~w623;
assign w2251 = ~w39 & ~w1123;
assign w2252 = ~w290 & ~w403;
assign w2253 = w2250 & w2251;
assign w2254 = w2252 & w2253;
assign w2255 = ~w337 & ~w476;
assign w2256 = ~w23 & ~w56;
assign w2257 = ~w180 & w2256;
assign w2258 = w1638 & w2249;
assign w2259 = w2255 & w2258;
assign w2260 = w2257 & w2259;
assign w2261 = w2254 & w2260;
assign w2262 = ~w88 & w1343;
assign w2263 = ~w218 & ~w572;
assign w2264 = ~w378 & ~w737;
assign w2265 = w469 & w1112;
assign w2266 = w2247 & w2248;
assign w2267 = w2263 & w2264;
assign w2268 = w2266 & w2267;
assign w2269 = ~w519 & w2265;
assign w2270 = w2262 & w2269;
assign w2271 = w2268 & w2270;
assign w2272 = w2246 & w2271;
assign w2273 = w2261 & w2272;
assign w2274 = ~w115 & ~w205;
assign w2275 = ~w282 & ~w325;
assign w2276 = ~w197 & ~w589;
assign w2277 = ~w181 & w673;
assign w2278 = ~w1104 & ~w1117;
assign w2279 = ~w173 & ~w652;
assign w2280 = ~w74 & ~w645;
assign w2281 = ~w130 & ~w1192;
assign w2282 = w620 & ~w710;
assign w2283 = w735 & w1309;
assign w2284 = w2281 & w2283;
assign w2285 = w2282 & w2284;
assign w2286 = ~w53 & ~w342;
assign w2287 = ~w316 & w2286;
assign w2288 = ~w86 & ~w264;
assign w2289 = ~w394 & ~w470;
assign w2290 = w2288 & w2289;
assign w2291 = w1376 & w1662;
assign w2292 = w1721 & w2185;
assign w2293 = w2274 & w2275;
assign w2294 = w2276 & w2278;
assign w2295 = w2279 & w2280;
assign w2296 = w2294 & w2295;
assign w2297 = w2292 & w2293;
assign w2298 = w2290 & w2291;
assign w2299 = w2277 & w2287;
assign w2300 = w2298 & w2299;
assign w2301 = w2296 & w2297;
assign w2302 = w2300 & w2301;
assign w2303 = w1927 & w2285;
assign w2304 = w2302 & w2303;
assign w2305 = w983 & w2304;
assign w2306 = w2273 & w2305;
assign w2307 = ~w172 & ~w239;
assign w2308 = ~w144 & w2307;
assign w2309 = ~w432 & ~w590;
assign w2310 = w1375 & w2309;
assign w2311 = w343 & w2052;
assign w2312 = ~w75 & w1633;
assign w2313 = w1689 & w2312;
assign w2314 = ~w255 & ~w696;
assign w2315 = w1266 & w2314;
assign w2316 = ~w355 & ~w838;
assign w2317 = ~w115 & ~w1117;
assign w2318 = w346 & w2317;
assign w2319 = w1105 & w1412;
assign w2320 = w2194 & w2316;
assign w2321 = w2319 & w2320;
assign w2322 = w2308 & w2310;
assign w2323 = w2311 & w2315;
assign w2324 = w2318 & w2323;
assign w2325 = w2321 & w2322;
assign w2326 = w2254 & w2313;
assign w2327 = w2325 & w2326;
assign w2328 = w2324 & w2327;
assign w2329 = ~w81 & ~w264;
assign w2330 = ~w147 & w2329;
assign w2331 = w40 & w184;
assign w2332 = ~w71 & ~w423;
assign w2333 = ~w126 & ~w378;
assign w2334 = ~w116 & ~w737;
assign w2335 = ~w368 & w948;
assign w2336 = ~w281 & ~w1051;
assign w2337 = ~w30 & ~w834;
assign w2338 = ~w161 & ~w181;
assign w2339 = ~w196 & ~w719;
assign w2340 = w2338 & w2339;
assign w2341 = w2087 & w2336;
assign w2342 = w2337 & w2341;
assign w2343 = w2051 & w2340;
assign w2344 = w2335 & w2343;
assign w2345 = w2342 & w2344;
assign w2346 = ~w185 & ~w190;
assign w2347 = ~w319 & ~w1953;
assign w2348 = ~w2331 & w2347;
assign w2349 = w137 & w2346;
assign w2350 = w1009 & w2008;
assign w2351 = w2332 & w2333;
assign w2352 = w2334 & w2351;
assign w2353 = w2349 & w2350;
assign w2354 = w2096 & w2348;
assign w2355 = w2330 & w2354;
assign w2356 = w2352 & w2353;
assign w2357 = w2355 & w2356;
assign w2358 = w2345 & w2357;
assign w2359 = ~w245 & w1758;
assign w2360 = w2358 & w2359;
assign w2361 = ~w50 & ~w422;
assign w2362 = ~w242 & ~w315;
assign w2363 = w1755 & w2362;
assign w2364 = ~w60 & ~w83;
assign w2365 = ~w388 & w2364;
assign w2366 = w99 & w648;
assign w2367 = w2361 & w2366;
assign w2368 = w2363 & w2365;
assign w2369 = w2367 & w2368;
assign w2370 = ~w164 & ~w463;
assign w2371 = ~w291 & ~w404;
assign w2372 = ~w252 & ~w321;
assign w2373 = w24 & w474;
assign w2374 = w561 & w1738;
assign w2375 = w2370 & w2371;
assign w2376 = w2372 & w2375;
assign w2377 = w2373 & w2374;
assign w2378 = w2376 & w2377;
assign w2379 = ~w322 & ~w450;
assign w2380 = ~w394 & w1890;
assign w2381 = ~w653 & w1685;
assign w2382 = ~w220 & ~w396;
assign w2383 = ~w543 & w2382;
assign w2384 = w358 & w386;
assign w2385 = w1769 & w2379;
assign w2386 = w2384 & w2385;
assign w2387 = w2380 & w2383;
assign w2388 = w2381 & w2387;
assign w2389 = w2386 & w2388;
assign w2390 = w2369 & w2378;
assign w2391 = w2389 & w2390;
assign w2392 = w2328 & w2391;
assign w2393 = w2360 & w2392;
assign w2394 = ~w2306 & ~w2393;
assign w2395 = ~w243 & ~w568;
assign w2396 = w906 & w2395;
assign w2397 = ~w221 & ~w262;
assign w2398 = ~w56 & ~w714;
assign w2399 = ~w140 & ~w741;
assign w2400 = ~w531 & ~w563;
assign w2401 = w2399 & w2400;
assign w2402 = ~w251 & ~w834;
assign w2403 = ~w400 & w2402;
assign w2404 = ~w42 & ~w163;
assign w2405 = ~w214 & ~w468;
assign w2406 = w162 & ~w547;
assign w2407 = w1340 & w2397;
assign w2408 = w2398 & w2404;
assign w2409 = w2405 & w2408;
assign w2410 = w2406 & w2407;
assign w2411 = w2401 & w2403;
assign w2412 = w2410 & w2411;
assign w2413 = w2396 & w2409;
assign w2414 = w2412 & w2413;
assign w2415 = w2378 & w2414;
assign w2416 = ~w115 & ~w173;
assign w2417 = ~w88 & ~w265;
assign w2418 = ~w128 & ~w313;
assign w2419 = ~w125 & ~w406;
assign w2420 = ~w281 & ~w562;
assign w2421 = ~w180 & ~w249;
assign w2422 = ~w396 & ~w1040;
assign w2423 = w2421 & w2422;
assign w2424 = w2094 & w2416;
assign w2425 = w2417 & w2418;
assign w2426 = w2419 & w2420;
assign w2427 = w2425 & w2426;
assign w2428 = w2423 & w2424;
assign w2429 = w2427 & w2428;
assign w2430 = w584 & w866;
assign w2431 = ~w341 & ~w710;
assign w2432 = w77 & w2431;
assign w2433 = ~w112 & ~w540;
assign w2434 = ~w65 & w2433;
assign w2435 = w2433 & w31564;
assign w2436 = ~w878 & w2276;
assign w2437 = w2011 & w2436;
assign w2438 = ~w345 & ~w644;
assign w2439 = ~w144 & ~w701;
assign w2440 = ~w30 & ~w459;
assign w2441 = ~w323 & ~w530;
assign w2442 = ~w170 & ~w451;
assign w2443 = ~w195 & ~w996;
assign w2444 = ~w266 & ~w694;
assign w2445 = ~w698 & ~w992;
assign w2446 = ~w279 & ~w403;
assign w2447 = w2443 & w2446;
assign w2448 = w2444 & w2445;
assign w2449 = w2447 & w2448;
assign w2450 = ~w420 & ~w538;
assign w2451 = ~w1117 & w2450;
assign w2452 = w1205 & w2451;
assign w2453 = w2077 & w2452;
assign w2454 = ~w146 & ~w357;
assign w2455 = w257 & w2454;
assign w2456 = ~w737 & w1265;
assign w2457 = w1757 & w2441;
assign w2458 = w2442 & w2457;
assign w2459 = w210 & w2456;
assign w2460 = w625 & w2310;
assign w2461 = w2455 & w2460;
assign w2462 = w2458 & w2459;
assign w2463 = w2449 & w2462;
assign w2464 = w2453 & w2461;
assign w2465 = w2463 & w2464;
assign w2466 = ~w123 & ~w212;
assign w2467 = ~w245 & ~w815;
assign w2468 = w2466 & w2467;
assign w2469 = w310 & w2438;
assign w2470 = w2439 & w2440;
assign w2471 = w2469 & w2470;
assign w2472 = w2430 & w2468;
assign w2473 = w2432 & w2472;
assign w2474 = w1272 & w2471;
assign w2475 = w2435 & w2437;
assign w2476 = w2474 & w2475;
assign w2477 = w2429 & w2473;
assign w2478 = w2476 & w2477;
assign w2479 = w2415 & w2478;
assign w2480 = w2465 & w2479;
assign w2481 = ~w30 & ~w1192;
assign w2482 = ~w163 & w1102;
assign w2483 = ~w85 & ~w95;
assign w2484 = ~w246 & w2483;
assign w2485 = ~w207 & ~w309;
assign w2486 = ~w312 & ~w341;
assign w2487 = ~w143 & ~w196;
assign w2488 = w814 & w2481;
assign w2489 = w2485 & w2486;
assign w2490 = w2487 & w2489;
assign w2491 = w2482 & w2488;
assign w2492 = w2484 & w2491;
assign w2493 = w2490 & w2492;
assign w2494 = ~w39 & ~w159;
assign w2495 = ~w218 & ~w563;
assign w2496 = ~w146 & ~w186;
assign w2497 = ~w714 & ~w1077;
assign w2498 = w2496 & w2497;
assign w2499 = ~w255 & ~w321;
assign w2500 = ~w451 & w2499;
assign w2501 = ~w116 & ~w450;
assign w2502 = ~w56 & ~w214;
assign w2503 = ~w319 & ~w339;
assign w2504 = ~w531 & w2503;
assign w2505 = w1489 & w2501;
assign w2506 = w2502 & w2505;
assign w2507 = w2500 & w2504;
assign w2508 = w2506 & w2507;
assign w2509 = w2498 & w2508;
assign w2510 = w13 & w1952;
assign w2511 = ~w432 & ~w671;
assign w2512 = ~w264 & ~w392;
assign w2513 = w774 & ~w2331;
assign w2514 = w2512 & w2513;
assign w2515 = ~w88 & ~w357;
assign w2516 = ~w89 & ~w287;
assign w2517 = ~w112 & ~w2510;
assign w2518 = w731 & w2517;
assign w2519 = w998 & w1125;
assign w2520 = w2511 & w2515;
assign w2521 = w2516 & w2520;
assign w2522 = w2518 & w2519;
assign w2523 = w2521 & w2522;
assign w2524 = w462 & w2514;
assign w2525 = w2523 & w2524;
assign w2526 = w2509 & w2525;
assign w2527 = ~w385 & ~w399;
assign w2528 = ~w217 & ~w647;
assign w2529 = w522 & w2528;
assign w2530 = ~w178 & ~w365;
assign w2531 = ~w418 & w2530;
assign w2532 = w1481 & w2527;
assign w2533 = w2531 & w2532;
assign w2534 = w2529 & w2533;
assign w2535 = ~w42 & w1421;
assign w2536 = w1052 & w1488;
assign w2537 = w2248 & w2317;
assign w2538 = w2494 & w2495;
assign w2539 = w2537 & w2538;
assign w2540 = w1267 & w2536;
assign w2541 = w2535 & w2540;
assign w2542 = w2539 & w2541;
assign w2543 = w2534 & w2542;
assign w2544 = w2493 & w2543;
assign w2545 = w894 & w2526;
assign w2546 = w2544 & w2545;
assign w2547 = ~w2480 & ~w2546;
assign w2548 = ~w355 & ~w388;
assign w2549 = ~w431 & ~w543;
assign w2550 = ~w130 & ~w323;
assign w2551 = w564 & w2550;
assign w2552 = ~w45 & ~w593;
assign w2553 = ~w56 & ~w249;
assign w2554 = w2552 & w2553;
assign w2555 = ~w267 & ~w590;
assign w2556 = w654 & w2555;
assign w2557 = ~w468 & ~w815;
assign w2558 = ~w97 & ~w357;
assign w2559 = ~w394 & ~w403;
assign w2560 = ~w86 & w2559;
assign w2561 = ~w254 & w1205;
assign w2562 = w2189 & w2557;
assign w2563 = w2558 & w2562;
assign w2564 = w1082 & w2561;
assign w2565 = w2560 & w2564;
assign w2566 = w2563 & w2565;
assign w2567 = w1355 & w1819;
assign w2568 = w1889 & w2567;
assign w2569 = ~w142 & ~w321;
assign w2570 = ~w313 & ~w878;
assign w2571 = ~w220 & ~w264;
assign w2572 = ~w143 & w2569;
assign w2573 = w2570 & w2571;
assign w2574 = w2572 & w2573;
assign w2575 = w1309 & w32657;
assign w2576 = ~w136 & ~w463;
assign w2577 = ~w458 & ~w720;
assign w2578 = w1152 & w2577;
assign w2579 = ~w98 & ~w239;
assign w2580 = w1009 & w2579;
assign w2581 = w997 & w2486;
assign w2582 = w2576 & w2581;
assign w2583 = w1930 & w2578;
assign w2584 = w2580 & w2583;
assign w2585 = w2568 & w2582;
assign w2586 = w2574 & w2575;
assign w2587 = w2585 & w2586;
assign w2588 = w2584 & w2587;
assign w2589 = w289 & w1356;
assign w2590 = w2034 & w2399;
assign w2591 = w2548 & w2549;
assign w2592 = w2590 & w2591;
assign w2593 = w150 & w2589;
assign w2594 = w1717 & w2551;
assign w2595 = w2554 & w2556;
assign w2596 = w2594 & w2595;
assign w2597 = w2592 & w2593;
assign w2598 = w2596 & w2597;
assign w2599 = w2566 & w2598;
assign w2600 = w1150 & w2599;
assign w2601 = w2588 & w2600;
assign w2602 = w2547 & ~w2601;
assign w2603 = ~w422 & ~w562;
assign w2604 = ~w112 & ~w597;
assign w2605 = ~w325 & ~w451;
assign w2606 = ~w815 & w2605;
assign w2607 = ~w30 & ~w582;
assign w2608 = ~w362 & w2607;
assign w2609 = ~w138 & ~w288;
assign w2610 = ~w125 & ~w838;
assign w2611 = w311 & w2610;
assign w2612 = w2177 & w2609;
assign w2613 = w2611 & w2612;
assign w2614 = w187 & w2613;
assign w2615 = ~w205 & ~w538;
assign w2616 = ~w720 & w2615;
assign w2617 = ~w190 & w617;
assign w2618 = w2052 & w2617;
assign w2619 = ~w39 & ~w1040;
assign w2620 = ~w287 & ~w622;
assign w2621 = ~w206 & ~w730;
assign w2622 = ~w385 & ~w389;
assign w2623 = w182 & w2622;
assign w2624 = w1435 & w2619;
assign w2625 = w2620 & w2621;
assign w2626 = w2624 & w2625;
assign w2627 = w2616 & w2623;
assign w2628 = w2626 & w2627;
assign w2629 = w2618 & w2628;
assign w2630 = ~w356 & ~w649;
assign w2631 = w836 & w2630;
assign w2632 = w1607 & w1942;
assign w2633 = w2279 & w2454;
assign w2634 = w2559 & w2603;
assign w2635 = w2604 & w2634;
assign w2636 = w2632 & w2633;
assign w2637 = w2606 & w2631;
assign w2638 = w2608 & w2637;
assign w2639 = w2635 & w2636;
assign w2640 = w2638 & w2639;
assign w2641 = w2614 & w2640;
assign w2642 = w2629 & w2641;
assign w2643 = ~w113 & ~w789;
assign w2644 = w2264 & w2643;
assign w2645 = ~w339 & ~w380;
assign w2646 = ~w363 & ~w432;
assign w2647 = ~w50 & ~w136;
assign w2648 = ~w319 & w2286;
assign w2649 = w2645 & w2646;
assign w2650 = w2647 & w2649;
assign w2651 = w2648 & w2650;
assign w2652 = ~w67 & ~w153;
assign w2653 = w1986 & w2652;
assign w2654 = ~w322 & ~w626;
assign w2655 = ~w95 & ~w292;
assign w2656 = ~w242 & ~w907;
assign w2657 = w17 & w2656;
assign w2658 = w2654 & w2655;
assign w2659 = w2657 & w2658;
assign w2660 = w2653 & w2659;
assign w2661 = w620 & ~w719;
assign w2662 = w1109 & w2661;
assign w2663 = ~w559 & ~w896;
assign w2664 = ~w89 & ~w446;
assign w2665 = w988 & w2664;
assign w2666 = w1533 & w2281;
assign w2667 = w2441 & w2487;
assign w2668 = w2663 & w2667;
assign w2669 = w2665 & w2666;
assign w2670 = w258 & w2644;
assign w2671 = w2669 & w2670;
assign w2672 = w2662 & w2668;
assign w2673 = w2671 & w2672;
assign w2674 = w2651 & w2660;
assign w2675 = w2673 & w2674;
assign w2676 = w2415 & w2675;
assign w2677 = w2642 & w2676;
assign w2678 = w2480 & w2546;
assign w2679 = ~w2677 & ~w2678;
assign w2680 = ~w2602 & ~w2679;
assign w2681 = ~w339 & ~w368;
assign w2682 = ~w127 & ~w1104;
assign w2683 = w1631 & w2682;
assign w2684 = ~w283 & ~w403;
assign w2685 = ~w312 & w2684;
assign w2686 = w2683 & w2685;
assign w2687 = w139 & ~w518;
assign w2688 = ~w53 & ~w337;
assign w2689 = ~w142 & ~w251;
assign w2690 = w179 & w1536;
assign w2691 = w1737 & w1772;
assign w2692 = w2557 & w2681;
assign w2693 = ~w2687 & w2688;
assign w2694 = w2689 & w2693;
assign w2695 = w2691 & w2692;
assign w2696 = w1311 & w2690;
assign w2697 = w2695 & w2696;
assign w2698 = w2686 & w2694;
assign w2699 = w2697 & w2698;
assign w2700 = ~w321 & ~w395;
assign w2701 = ~w345 & ~w568;
assign w2702 = ~w1043 & w2701;
assign w2703 = w532 & w2700;
assign w2704 = w2702 & w2703;
assign w2705 = ~w75 & ~w116;
assign w2706 = w93 & w831;
assign w2707 = ~w140 & ~w406;
assign w2708 = ~w260 & ~w559;
assign w2709 = ~w237 & ~w582;
assign w2710 = ~w23 & ~w239;
assign w2711 = ~w76 & ~w282;
assign w2712 = ~w538 & ~w563;
assign w2713 = w2711 & w2712;
assign w2714 = w2710 & w2713;
assign w2715 = ~w183 & ~w583;
assign w2716 = w58 & w707;
assign w2717 = ~w734 & ~w896;
assign w2718 = ~w56 & w2717;
assign w2719 = ~w95 & ~w153;
assign w2720 = ~w188 & ~w644;
assign w2721 = ~w2716 & w2720;
assign w2722 = w2715 & w2719;
assign w2723 = w2721 & w2722;
assign w2724 = w1495 & w2011;
assign w2725 = w2482 & w2718;
assign w2726 = w2724 & w2725;
assign w2727 = w2714 & w2723;
assign w2728 = w2726 & w2727;
assign w2729 = ~w89 & ~w316;
assign w2730 = ~w205 & ~w590;
assign w2731 = ~w245 & ~w463;
assign w2732 = w517 & w2731;
assign w2733 = w1454 & w2729;
assign w2734 = w2730 & w2733;
assign w2735 = w2732 & w2734;
assign w2736 = w2728 & w2735;
assign w2737 = w137 & w773;
assign w2738 = ~w83 & w1658;
assign w2739 = ~w291 & ~w420;
assign w2740 = ~w730 & ~w895;
assign w2741 = w2739 & w2740;
assign w2742 = ~w701 & ~w834;
assign w2743 = ~w156 & ~w1117;
assign w2744 = ~w254 & ~w366;
assign w2745 = ~w392 & w2744;
assign w2746 = w728 & w1193;
assign w2747 = w1690 & w2742;
assign w2748 = w2743 & w2747;
assign w2749 = w2745 & w2746;
assign w2750 = w2737 & w2738;
assign w2751 = w2741 & w2750;
assign w2752 = w2748 & w2749;
assign w2753 = w2751 & w2752;
assign w2754 = ~w267 & ~w2706;
assign w2755 = w1041 & w2754;
assign w2756 = w2397 & w2705;
assign w2757 = w2707 & w2708;
assign w2758 = w2709 & w2757;
assign w2759 = w2755 & w2756;
assign w2760 = w2758 & w2759;
assign w2761 = w200 & w2704;
assign w2762 = w2760 & w2761;
assign w2763 = w1404 & w1700;
assign w2764 = w2762 & w2763;
assign w2765 = w2699 & w2753;
assign w2766 = w2764 & w2765;
assign w2767 = w2736 & w2766;
assign w2768 = w2734 & w31565;
assign w2769 = w2728 & w2768;
assign w2770 = w293 & ~w593;
assign w2771 = ~w46 & ~w157;
assign w2772 = ~w366 & ~w447;
assign w2773 = ~w197 & ~w393;
assign w2774 = ~w418 & ~w653;
assign w2775 = ~w352 & ~w473;
assign w2776 = w2771 & w2775;
assign w2777 = w2772 & w2773;
assign w2778 = w2774 & w2777;
assign w2779 = w2770 & w2776;
assign w2780 = w2778 & w2779;
assign w2781 = ~w212 & ~w470;
assign w2782 = ~w597 & ~w1077;
assign w2783 = ~w138 & w2250;
assign w2784 = ~w388 & ~w396;
assign w2785 = ~w314 & ~w325;
assign w2786 = ~w86 & ~w530;
assign w2787 = w596 & w1464;
assign w2788 = w2119 & w2334;
assign w2789 = w2784 & w2785;
assign w2790 = w2786 & w2789;
assign w2791 = w2787 & w2788;
assign w2792 = w1053 & w2783;
assign w2793 = w2791 & w2792;
assign w2794 = w1684 & w2790;
assign w2795 = w2793 & w2794;
assign w2796 = ~w378 & ~w450;
assign w2797 = ~w568 & w2796;
assign w2798 = ~w190 & ~w878;
assign w2799 = w129 & w2798;
assign w2800 = ~w265 & ~w451;
assign w2801 = ~w75 & ~w81;
assign w2802 = ~w312 & w2800;
assign w2803 = w2801 & w2802;
assign w2804 = ~w428 & ~w1104;
assign w2805 = ~w719 & ~w992;
assign w2806 = w1871 & w2805;
assign w2807 = ~w459 & ~w652;
assign w2808 = ~w339 & w2807;
assign w2809 = ~w42 & ~w208;
assign w2810 = w950 & w1334;
assign w2811 = w1764 & w2607;
assign w2812 = w2804 & w2809;
assign w2813 = w2811 & w2812;
assign w2814 = w2797 & w2810;
assign w2815 = w2799 & w2806;
assign w2816 = w2808 & w2815;
assign w2817 = w2813 & w2814;
assign w2818 = w2803 & w2817;
assign w2819 = w2816 & w2818;
assign w2820 = ~w62 & ~w287;
assign w2821 = ~w1953 & ~w1965;
assign w2822 = w2820 & w2821;
assign w2823 = w253 & w754;
assign w2824 = w833 & w1584;
assign w2825 = w1607 & w2781;
assign w2826 = w2782 & w2825;
assign w2827 = w2823 & w2824;
assign w2828 = w700 & w2822;
assign w2829 = w2827 & w2828;
assign w2830 = w1115 & w2826;
assign w2831 = w2829 & w2830;
assign w2832 = w2780 & w2831;
assign w2833 = w2795 & w2832;
assign w2834 = w2769 & w2819;
assign w2835 = w2833 & w2834;
assign w2836 = ~w2767 & ~w2835;
assign w2837 = ~w2546 & ~w2767;
assign w2838 = ~w2836 & ~w2837;
assign w2839 = ~w42 & ~w248;
assign w2840 = ~w349 & ~w389;
assign w2841 = ~w626 & w2840;
assign w2842 = ~w446 & ~w1043;
assign w2843 = w2839 & w2842;
assign w2844 = w2841 & w2843;
assign w2845 = ~w213 & ~w323;
assign w2846 = ~w265 & ~w429;
assign w2847 = ~w352 & w2846;
assign w2848 = ~w262 & ~w355;
assign w2849 = ~w365 & w2848;
assign w2850 = ~w113 & w137;
assign w2851 = w726 & w1422;
assign w2852 = w1929 & w2152;
assign w2853 = w2845 & w2852;
assign w2854 = w2850 & w2851;
assign w2855 = w2847 & w2849;
assign w2856 = w2854 & w2855;
assign w2857 = w2449 & w2853;
assign w2858 = w2844 & w2857;
assign w2859 = w2856 & w2858;
assign w2860 = ~w125 & w1153;
assign w2861 = w179 & ~w395;
assign w2862 = ~w239 & ~w369;
assign w2863 = ~w538 & w2862;
assign w2864 = w465 & w586;
assign w2865 = w1640 & w2416;
assign w2866 = w2619 & w2865;
assign w2867 = w2863 & w2864;
assign w2868 = w2860 & w2861;
assign w2869 = w2867 & w2868;
assign w2870 = w2866 & w2869;
assign w2871 = ~w212 & ~w543;
assign w2872 = ~w196 & ~w431;
assign w2873 = ~w183 & ~w428;
assign w2874 = ~w237 & ~w243;
assign w2875 = ~w580 & ~w619;
assign w2876 = ~w789 & w2875;
assign w2877 = w99 & w2516;
assign w2878 = w2873 & w2874;
assign w2879 = w2877 & w2878;
assign w2880 = w2876 & w2879;
assign w2881 = ~w283 & ~w531;
assign w2882 = ~w23 & ~w319;
assign w2883 = ~w325 & w2882;
assign w2884 = w2881 & w2883;
assign w2885 = w80 & w31566;
assign w2886 = ~w191 & ~w322;
assign w2887 = ~w730 & w1918;
assign w2888 = ~w152 & ~w207;
assign w2889 = ~w282 & ~w420;
assign w2890 = ~w1123 & w2889;
assign w2891 = w1776 & w2888;
assign w2892 = w2189 & ~w2885;
assign w2893 = w2886 & w2892;
assign w2894 = w2890 & w2891;
assign w2895 = w937 & w2500;
assign w2896 = w2887 & w2895;
assign w2897 = w2893 & w2894;
assign w2898 = w761 & w2437;
assign w2899 = w2884 & w2898;
assign w2900 = w2896 & w2897;
assign w2901 = w2899 & w2900;
assign w2902 = ~w85 & ~w249;
assign w2903 = ~w476 & ~w1104;
assign w2904 = w2902 & w2903;
assign w2905 = w17 & w158;
assign w2906 = w584 & w911;
assign w2907 = w1435 & w2036;
assign w2908 = w2871 & w2872;
assign w2909 = w2907 & w2908;
assign w2910 = w2905 & w2906;
assign w2911 = w1660 & w2904;
assign w2912 = w2910 & w2911;
assign w2913 = w2909 & w2912;
assign w2914 = w2880 & w2913;
assign w2915 = w2870 & w2914;
assign w2916 = w2859 & w2901;
assign w2917 = w2915 & w2916;
assign w2918 = ~w2835 & ~w2917;
assign w2919 = w2838 & ~w2918;
assign w2920 = w2680 & w2919;
assign w2921 = w2767 & w2835;
assign w2922 = w2546 & w2767;
assign w2923 = ~w2921 & ~w2922;
assign w2924 = ~w2918 & ~w2923;
assign w2925 = ~w123 & ~w585;
assign w2926 = w1266 & w2925;
assign w2927 = ~w156 & ~w896;
assign w2928 = w1464 & w2927;
assign w2929 = ~w248 & ~w895;
assign w2930 = ~w60 & w2929;
assign w2931 = ~w180 & ~w710;
assign w2932 = ~w218 & w1632;
assign w2933 = w2438 & w2705;
assign w2934 = w2931 & w2933;
assign w2935 = w2930 & w2932;
assign w2936 = w2934 & w2935;
assign w2937 = ~w113 & ~w128;
assign w2938 = ~w246 & ~w422;
assign w2939 = w2937 & w2938;
assign w2940 = ~w98 & ~w470;
assign w2941 = ~w134 & ~w720;
assign w2942 = ~w252 & ~w838;
assign w2943 = ~w261 & ~w647;
assign w2944 = ~w149 & ~w432;
assign w2945 = w1942 & w2944;
assign w2946 = w2684 & w2941;
assign w2947 = w2942 & w2943;
assign w2948 = w2946 & w2947;
assign w2949 = w2945 & w2948;
assign w2950 = w2099 & w2949;
assign w2951 = ~w217 & ~w266;
assign w2952 = ~w698 & w2951;
assign w2953 = w240 & w628;
assign w2954 = ~w2687 & w2940;
assign w2955 = w2953 & w2954;
assign w2956 = w461 & w2952;
assign w2957 = w1401 & w1740;
assign w2958 = w2926 & w2928;
assign w2959 = w2939 & w2958;
assign w2960 = w2956 & w2957;
assign w2961 = w2955 & w2960;
assign w2962 = w2936 & w2959;
assign w2963 = w2961 & w2962;
assign w2964 = w2950 & w2963;
assign w2965 = ~w181 & ~w260;
assign w2966 = ~w45 & ~w396;
assign w2967 = ~w572 & w1238;
assign w2968 = w2965 & w2966;
assign w2969 = w2967 & w2968;
assign w2970 = ~w94 & ~w1192;
assign w2971 = ~w166 & ~w325;
assign w2972 = w1643 & w2970;
assign w2973 = w2971 & w2972;
assign w2974 = w958 & w2774;
assign w2975 = ~w366 & w1873;
assign w2976 = w1220 & ~w1223;
assign w2977 = w54 & w2976;
assign w2978 = ~w321 & ~w394;
assign w2979 = w1309 & w2978;
assign w2980 = ~w42 & ~w146;
assign w2981 = ~w242 & ~w2134;
assign w2982 = w2980 & w2981;
assign w2983 = w1869 & w2982;
assign w2984 = w2979 & w2983;
assign w2985 = ~w337 & ~w385;
assign w2986 = w1586 & w31567;
assign w2987 = w2984 & w2986;
assign w2988 = ~w178 & ~w907;
assign w2989 = ~w127 & ~w319;
assign w2990 = ~w97 & ~w992;
assign w2991 = ~w619 & ~w671;
assign w2992 = ~w147 & w1422;
assign w2993 = w2988 & w2989;
assign w2994 = w2990 & w2991;
assign w2995 = w2993 & w2994;
assign w2996 = w2992 & w2995;
assign w2997 = ~w878 & ~w2977;
assign w2998 = w1690 & w2997;
assign w2999 = w2974 & w2998;
assign w3000 = w2975 & w2999;
assign w3001 = w1211 & w2969;
assign w3002 = w2973 & w3001;
assign w3003 = w2996 & w3000;
assign w3004 = w3002 & w3003;
assign w3005 = w751 & w2987;
assign w3006 = w3004 & w3005;
assign w3007 = w2964 & w3006;
assign w3008 = ~w207 & w1102;
assign w3009 = ~w238 & ~w393;
assign w3010 = ~w544 & w3009;
assign w3011 = w1102 & w31568;
assign w3012 = w3010 & w3011;
assign w3013 = ~w459 & ~w531;
assign w3014 = ~w312 & ~w1192;
assign w3015 = ~w345 & w986;
assign w3016 = w3014 & w3015;
assign w3017 = ~w547 & w1536;
assign w3018 = w1490 & w3017;
assign w3019 = w853 & w876;
assign w3020 = w1419 & w3019;
assign w3021 = ~w216 & ~w1043;
assign w3022 = w1316 & w2729;
assign w3023 = w3021 & w3022;
assign w3024 = ~w60 & ~w164;
assign w3025 = ~w366 & ~w720;
assign w3026 = w3024 & w3025;
assign w3027 = ~w53 & ~w131;
assign w3028 = ~w396 & w3027;
assign w3029 = w3026 & w3028;
assign w3030 = ~w183 & ~w1040;
assign w3031 = w1044 & w2088;
assign w3032 = w3030 & w3031;
assign w3033 = w740 & w2318;
assign w3034 = w2841 & w3033;
assign w3035 = w3023 & w3032;
assign w3036 = w3029 & w3035;
assign w3037 = w3034 & w3036;
assign w3038 = w280 & w1069;
assign w3039 = w2717 & w2804;
assign w3040 = w3013 & w3039;
assign w3041 = w2887 & w3038;
assign w3042 = w3040 & w3041;
assign w3043 = w1963 & w3016;
assign w3044 = w3018 & w3020;
assign w3045 = w3043 & w3044;
assign w3046 = w3012 & w3042;
assign w3047 = w3045 & w3046;
assign w3048 = w3037 & w3047;
assign w3049 = w2360 & w3048;
assign w3050 = ~w3007 & ~w3049;
assign w3051 = w3007 & w3049;
assign w3052 = ~w3050 & ~w3051;
assign w3053 = w2835 & w2917;
assign w3054 = w2917 & w3007;
assign w3055 = ~w3053 & ~w3054;
assign w3056 = w3052 & w3055;
assign w3057 = ~w2924 & w3056;
assign w3058 = ~w2920 & w3057;
assign w3059 = ~w265 & w2014;
assign w3060 = ~w136 & ~w741;
assign w3061 = w424 & w3060;
assign w3062 = w912 & w3061;
assign w3063 = ~w152 & ~w217;
assign w3064 = w564 & w3063;
assign w3065 = ~w362 & ~w834;
assign w3066 = ~w95 & w3065;
assign w3067 = ~w167 & ~w391;
assign w3068 = ~w671 & w3067;
assign w3069 = w627 & w1534;
assign w3070 = w2093 & w2501;
assign w3071 = w3069 & w3070;
assign w3072 = w1453 & w3068;
assign w3073 = w3059 & w3064;
assign w3074 = w3066 & w3073;
assign w3075 = w3071 & w3072;
assign w3076 = w3062 & w3075;
assign w3077 = w2780 & w3074;
assign w3078 = w3076 & w3077;
assign w3079 = ~w590 & ~w815;
assign w3080 = ~w214 & ~w623;
assign w3081 = ~w60 & ~w312;
assign w3082 = w263 & w3081;
assign w3083 = w324 & w935;
assign w3084 = w1690 & w2942;
assign w3085 = w3079 & w3080;
assign w3086 = w3084 & w3085;
assign w3087 = w3082 & w3083;
assign w3088 = w187 & w3087;
assign w3089 = w3086 & w3088;
assign w3090 = ~w149 & ~w254;
assign w3091 = w346 & w3090;
assign w3092 = ~w166 & ~w315;
assign w3093 = ~w206 & ~w278;
assign w3094 = ~w378 & ~w429;
assign w3095 = ~w541 & ~w1123;
assign w3096 = w3094 & w3095;
assign w3097 = w3092 & w3093;
assign w3098 = w3096 & w3097;
assign w3099 = ~w207 & ~w395;
assign w3100 = ~w128 & ~w732;
assign w3101 = ~w470 & ~w818;
assign w3102 = ~w242 & ~w647;
assign w3103 = ~w342 & w3102;
assign w3104 = ~w127 & ~w321;
assign w3105 = w1052 & w3104;
assign w3106 = w1268 & w1686;
assign w3107 = w1756 & w2087;
assign w3108 = w3099 & w3100;
assign w3109 = w3101 & w3108;
assign w3110 = w3106 & w3107;
assign w3111 = w3091 & w3105;
assign w3112 = w3103 & w3111;
assign w3113 = w3109 & w3110;
assign w3114 = w3098 & w3113;
assign w3115 = w3112 & w3114;
assign w3116 = ~w124 & ~w213;
assign w3117 = ~w389 & ~w597;
assign w3118 = ~w369 & w1413;
assign w3119 = ~w559 & ~w992;
assign w3120 = w338 & ~w356;
assign w3121 = w3119 & w3120;
assign w3122 = ~w540 & ~w776;
assign w3123 = ~w10 & ~w583;
assign w3124 = ~w288 & ~w313;
assign w3125 = ~w89 & ~w153;
assign w3126 = ~w468 & w3125;
assign w3127 = w405 & w1265;
assign w3128 = w3116 & w3117;
assign w3129 = w3122 & w3123;
assign w3130 = w3124 & w3129;
assign w3131 = w3127 & w3128;
assign w3132 = w3118 & w3126;
assign w3133 = w3131 & w3132;
assign w3134 = w725 & w3130;
assign w3135 = w3121 & w3134;
assign w3136 = w3133 & w3135;
assign w3137 = w3089 & w3136;
assign w3138 = w3078 & w3115;
assign w3139 = w3137 & w3138;
assign w3140 = ~w649 & w2494;
assign w3141 = ~w282 & ~w580;
assign w3142 = ~w67 & ~w267;
assign w3143 = ~w337 & w3142;
assign w3144 = ~w138 & ~w741;
assign w3145 = w1661 & w3144;
assign w3146 = w2036 & w2579;
assign w3147 = w2647 & w3141;
assign w3148 = w3146 & w3147;
assign w3149 = w3140 & w3145;
assign w3150 = w3143 & w3149;
assign w3151 = w3148 & w3150;
assign w3152 = w257 & ~w590;
assign w3153 = w1691 & w3152;
assign w3154 = ~w323 & ~w730;
assign w3155 = ~w205 & ~w1051;
assign w3156 = ~w710 & w939;
assign w3157 = w3124 & w3155;
assign w3158 = w3156 & w3157;
assign w3159 = ~w173 & ~w322;
assign w3160 = ~w143 & ~w540;
assign w3161 = ~w94 & w587;
assign w3162 = w604 & w617;
assign w3163 = w1042 & w3162;
assign w3164 = w1642 & w3161;
assign w3165 = w2403 & w3164;
assign w3166 = w3163 & w3165;
assign w3167 = ~w181 & ~w694;
assign w3168 = ~w544 & w1870;
assign w3169 = ~w183 & ~w907;
assign w3170 = ~w147 & w3169;
assign w3171 = ~w186 & w469;
assign w3172 = w1689 & w1720;
assign w3173 = w1988 & w3167;
assign w3174 = w3172 & w3173;
assign w3175 = w2335 & w3171;
assign w3176 = w3008 & w3168;
assign w3177 = w3170 & w3176;
assign w3178 = w3174 & w3175;
assign w3179 = w3177 & w3178;
assign w3180 = w3166 & w3179;
assign w3181 = ~w23 & ~w314;
assign w3182 = ~w559 & ~w732;
assign w3183 = w3181 & w3182;
assign w3184 = w866 & w2182;
assign w3185 = w2398 & w2558;
assign w3186 = w3154 & w3159;
assign w3187 = w3160 & w3186;
assign w3188 = w3184 & w3185;
assign w3189 = w3183 & w3188;
assign w3190 = w1570 & w3187;
assign w3191 = w3153 & w3158;
assign w3192 = w3190 & w3191;
assign w3193 = w3189 & w3192;
assign w3194 = w3151 & w3193;
assign w3195 = w2819 & w3180;
assign w3196 = w3194 & w3195;
assign w3197 = ~w3139 & ~w3196;
assign w3198 = ~w2917 & ~w3007;
assign w3199 = ~w3049 & ~w3139;
assign w3200 = ~w3050 & ~w3199;
assign w3201 = ~w3198 & w3200;
assign w3202 = w3200 & w32658;
assign w3203 = w3049 & w3139;
assign w3204 = w3139 & w3196;
assign w3205 = ~w3203 & ~w3204;
assign w3206 = w1560 & w31569;
assign w3207 = w182 & ~w538;
assign w3208 = ~w39 & ~w208;
assign w3209 = ~w237 & ~w562;
assign w3210 = ~w42 & ~w622;
assign w3211 = ~w18 & ~w1104;
assign w3212 = ~w388 & ~w644;
assign w3213 = ~w186 & w3212;
assign w3214 = ~w541 & ~w597;
assign w3215 = ~w531 & ~w590;
assign w3216 = ~w95 & w3214;
assign w3217 = w3215 & w3216;
assign w3218 = ~w647 & w948;
assign w3219 = w1268 & w1719;
assign w3220 = w3211 & w3219;
assign w3221 = w3213 & w3218;
assign w3222 = w3220 & w3221;
assign w3223 = w3217 & w3222;
assign w3224 = w702 & w1287;
assign w3225 = w2184 & w2929;
assign w3226 = w3208 & w3209;
assign w3227 = w3210 & w3226;
assign w3228 = w3224 & w3225;
assign w3229 = w155 & w3207;
assign w3230 = w3228 & w3229;
assign w3231 = w1602 & w3227;
assign w3232 = w3230 & w3231;
assign w3233 = w3223 & w3232;
assign w3234 = ~w190 & w1152;
assign w3235 = w1273 & w3234;
assign w3236 = w866 & w1860;
assign w3237 = ~w243 & ~w583;
assign w3238 = w1492 & w2402;
assign w3239 = ~w135 & ~w896;
assign w3240 = ~w81 & ~w283;
assign w3241 = w816 & w3240;
assign w3242 = w3237 & w3239;
assign w3243 = w3241 & w3242;
assign w3244 = w3236 & w3238;
assign w3245 = w3243 & w3244;
assign w3246 = ~w290 & w627;
assign w3247 = ~w254 & ~w365;
assign w3248 = ~w65 & ~w623;
assign w3249 = ~w127 & ~w366;
assign w3250 = ~w543 & w3249;
assign w3251 = w2940 & w3247;
assign w3252 = w3248 & w3251;
assign w3253 = w3250 & w3252;
assign w3254 = ~w88 & ~w246;
assign w3255 = w148 & w3254;
assign w3256 = w1281 & w1562;
assign w3257 = w1967 & w2443;
assign w3258 = w2743 & w3159;
assign w3259 = w3257 & w3258;
assign w3260 = w3255 & w3256;
assign w3261 = w478 & w3246;
assign w3262 = w3260 & w3261;
assign w3263 = w3235 & w3259;
assign w3264 = w3262 & w3263;
assign w3265 = w3245 & w3253;
assign w3266 = w3264 & w3265;
assign w3267 = w3233 & w3266;
assign w3268 = w3206 & w3267;
assign w3269 = w3196 & ~w3268;
assign w3270 = ~w3196 & w3268;
assign w3271 = ~w3269 & ~w3270;
assign w3272 = w3205 & ~w3271;
assign w3273 = (w3272 & w3058) | (w3272 & w31570) | (w3058 & w31570);
assign w3274 = ~w147 & ~w463;
assign w3275 = ~w81 & ~w710;
assign w3276 = ~w368 & w3275;
assign w3277 = ~w30 & ~w88;
assign w3278 = ~w115 & ~w314;
assign w3279 = ~w355 & w3278;
assign w3280 = w3277 & w3279;
assign w3281 = w3276 & w3280;
assign w3282 = ~w260 & ~w878;
assign w3283 = ~w144 & ~w151;
assign w3284 = ~w394 & w3283;
assign w3285 = ~w65 & ~w475;
assign w3286 = ~w349 & ~w352;
assign w3287 = ~w251 & w1119;
assign w3288 = ~w149 & ~w458;
assign w3289 = ~w907 & w3288;
assign w3290 = w2008 & w3285;
assign w3291 = w3286 & w3290;
assign w3292 = w3287 & w3289;
assign w3293 = w3291 & w3292;
assign w3294 = ~w140 & ~w206;
assign w3295 = ~w362 & ~w619;
assign w3296 = w3294 & w3295;
assign w3297 = w2796 & w3274;
assign w3298 = w3282 & w3297;
assign w3299 = w951 & w3296;
assign w3300 = w3284 & w3299;
assign w3301 = w3023 & w3298;
assign w3302 = w3300 & w3301;
assign w3303 = w3281 & w3293;
assign w3304 = w3302 & w3303;
assign w3305 = ~w195 & ~w429;
assign w3306 = ~w97 & w1238;
assign w3307 = w3305 & w3306;
assign w3308 = ~w34 & ~w242;
assign w3309 = ~w252 & w1052;
assign w3310 = w2332 & w2717;
assign w3311 = w3308 & w3310;
assign w3312 = w3309 & w3311;
assign w3313 = ~w191 & w3116;
assign w3314 = ~w239 & ~w476;
assign w3315 = w359 & w3314;
assign w3316 = w646 & w2276;
assign w3317 = w3099 & w3316;
assign w3318 = w3010 & w3315;
assign w3319 = w3143 & w3313;
assign w3320 = w3318 & w3319;
assign w3321 = w3029 & w3317;
assign w3322 = w3307 & w3321;
assign w3323 = w2062 & w3320;
assign w3324 = w3312 & w3323;
assign w3325 = w3322 & w3324;
assign w3326 = w3325 & w32659;
assign w3327 = w3268 & w3326;
assign w3328 = (w3058 & w32660) | (w3058 & w32661) | (w32660 & w32661);
assign w3329 = ~w423 & ~w720;
assign w3330 = ~w83 & ~w163;
assign w3331 = ~w94 & ~w216;
assign w3332 = ~w789 & w3331;
assign w3333 = ~w127 & ~w135;
assign w3334 = ~w1117 & w3333;
assign w3335 = w43 & w1436;
assign w3336 = w1524 & w2804;
assign w3337 = w3330 & w3336;
assign w3338 = w3334 & w3335;
assign w3339 = w2287 & w3332;
assign w3340 = w3338 & w3339;
assign w3341 = w3337 & w3340;
assign w3342 = ~w89 & ~w649;
assign w3343 = ~w181 & w3342;
assign w3344 = ~w151 & ~w238;
assign w3345 = ~w217 & ~w369;
assign w3346 = w3344 & w3345;
assign w3347 = ~w352 & ~w396;
assign w3348 = ~w207 & ~w288;
assign w3349 = ~w590 & w3348;
assign w3350 = w2871 & w3347;
assign w3351 = w3349 & w3350;
assign w3352 = w3313 & w3343;
assign w3353 = w3346 & w3352;
assign w3354 = w2803 & w3351;
assign w3355 = w3353 & w3354;
assign w3356 = w1613 & w3355;
assign w3357 = w3341 & w3356;
assign w3358 = w908 & w1550;
assign w3359 = w2255 & w2552;
assign w3360 = w3329 & w3359;
assign w3361 = w2797 & w3358;
assign w3362 = w3360 & w3361;
assign w3363 = w3356 & w32662;
assign w3364 = ~w62 & ~w218;
assign w3365 = ~w237 & ~w468;
assign w3366 = ~w46 & ~w321;
assign w3367 = w3364 & w3366;
assign w3368 = w3365 & w3367;
assign w3369 = ~w281 & ~w583;
assign w3370 = ~w157 & ~w195;
assign w3371 = ~w291 & ~w559;
assign w3372 = w3370 & w3371;
assign w3373 = ~w385 & ~w475;
assign w3374 = ~w541 & ~w645;
assign w3375 = w3373 & w3374;
assign w3376 = w320 & w586;
assign w3377 = w2444 & w3369;
assign w3378 = w3376 & w3377;
assign w3379 = w2363 & w3375;
assign w3380 = w2401 & w3372;
assign w3381 = w3379 & w3380;
assign w3382 = w812 & w3378;
assign w3383 = w1359 & w3382;
assign w3384 = w3381 & w3383;
assign w3385 = ~w399 & w624;
assign w3386 = ~w245 & ~w1040;
assign w3387 = ~w86 & ~w144;
assign w3388 = w960 & w1330;
assign w3389 = w3386 & w3387;
assign w3390 = w3388 & w3389;
assign w3391 = ~w580 & ~w944;
assign w3392 = ~w2706 & w3391;
assign w3393 = w449 & w1770;
assign w3394 = w1895 & w1988;
assign w3395 = w2433 & w3394;
assign w3396 = w3392 & w3393;
assign w3397 = w2928 & w3385;
assign w3398 = w3396 & w3397;
assign w3399 = w3368 & w3395;
assign w3400 = w3390 & w3399;
assign w3401 = w3398 & w3400;
assign w3402 = w3384 & w3401;
assign w3403 = w3363 & w3402;
assign w3404 = ~w238 & ~w734;
assign w3405 = ~w191 & ~w422;
assign w3406 = ~w838 & w3405;
assign w3407 = w1862 & w3406;
assign w3408 = w695 & w790;
assign w3409 = w1424 & w1738;
assign w3410 = w3404 & w3409;
assign w3411 = w1537 & w3408;
assign w3412 = w2608 & w3246;
assign w3413 = w3411 & w3412;
assign w3414 = w3407 & w3410;
assign w3415 = w3413 & w3414;
assign w3416 = w2200 & w3415;
assign w3417 = ~w283 & ~w369;
assign w3418 = ~w1123 & w3417;
assign w3419 = ~w264 & ~w468;
assign w3420 = w289 & w3419;
assign w3421 = ~w18 & ~w142;
assign w3422 = ~w580 & ~w732;
assign w3423 = ~w896 & w3422;
assign w3424 = ~w186 & w3421;
assign w3425 = w3423 & w3424;
assign w3426 = ~w72 & ~w378;
assign w3427 = ~w281 & ~w315;
assign w3428 = ~w89 & ~w172;
assign w3429 = ~w420 & ~w540;
assign w3430 = w1430 & w3429;
assign w3431 = w1435 & w2183;
assign w3432 = w3430 & w3431;
assign w3433 = ~w140 & w2966;
assign w3434 = ~w246 & ~w741;
assign w3435 = ~w10 & ~w1117;
assign w3436 = w293 & w3435;
assign w3437 = w603 & w2089;
assign w3438 = w2871 & w3434;
assign w3439 = w3437 & w3438;
assign w3440 = w3433 & w3436;
assign w3441 = w3439 & w3440;
assign w3442 = ~w144 & ~w696;
assign w3443 = w1151 & w3442;
assign w3444 = ~w126 & ~w432;
assign w3445 = ~w337 & ~w623;
assign w3446 = w3444 & w3445;
assign w3447 = w3426 & w3427;
assign w3448 = w3428 & w3447;
assign w3449 = w3170 & w3443;
assign w3450 = w3446 & w3449;
assign w3451 = w3432 & w3448;
assign w3452 = w3450 & w3451;
assign w3453 = w3441 & w3452;
assign w3454 = w360 & ~w458;
assign w3455 = w3452 & w32663;
assign w3456 = ~w128 & ~w538;
assign w3457 = w77 & ~w355;
assign w3458 = ~w368 & w1026;
assign w3459 = w3364 & w3456;
assign w3460 = w3458 & w3459;
assign w3461 = w1453 & w2133;
assign w3462 = w3457 & w3461;
assign w3463 = w3460 & w3462;
assign w3464 = ~w207 & ~w1077;
assign w3465 = w754 & w857;
assign w3466 = w2708 & w3464;
assign w3467 = w3465 & w3466;
assign w3468 = w1664 & w2178;
assign w3469 = w3418 & w3420;
assign w3470 = w3468 & w3469;
assign w3471 = w1761 & w3467;
assign w3472 = w3425 & w3471;
assign w3473 = w3470 & w3472;
assign w3474 = w3463 & w3473;
assign w3475 = w3474 & w32664;
assign w3476 = ~w3403 & ~w3475;
assign w3477 = ~w134 & ~w776;
assign w3478 = ~w95 & ~w423;
assign w3479 = ~w337 & ~w696;
assign w3480 = ~w737 & w3479;
assign w3481 = ~w142 & ~w217;
assign w3482 = w192 & w3481;
assign w3483 = w962 & w1360;
assign w3484 = w2931 & w3478;
assign w3485 = w3483 & w3484;
assign w3486 = w3480 & w3482;
assign w3487 = w3485 & w3486;
assign w3488 = ~w83 & ~w265;
assign w3489 = ~w188 & ~w255;
assign w3490 = ~w352 & ~w623;
assign w3491 = ~w1192 & w3490;
assign w3492 = w3489 & w3491;
assign w3493 = ~w315 & ~w653;
assign w3494 = w139 & w1288;
assign w3495 = ~w313 & ~w420;
assign w3496 = w1098 & ~w3494;
assign w3497 = w3370 & w3493;
assign w3498 = w3495 & w3497;
assign w3499 = w3496 & w3498;
assign w3500 = ~w124 & ~w177;
assign w3501 = ~w996 & w3500;
assign w3502 = ~w74 & ~w582;
assign w3503 = ~w458 & ~w1040;
assign w3504 = w1080 & w3503;
assign w3505 = w3502 & w3504;
assign w3506 = ~w136 & ~w428;
assign w3507 = w598 & w3506;
assign w3508 = w1571 & w1850;
assign w3509 = w2978 & w3488;
assign w3510 = w3508 & w3509;
assign w3511 = w3501 & w3507;
assign w3512 = w3510 & w3511;
assign w3513 = w3492 & w3505;
assign w3514 = w3512 & w3513;
assign w3515 = w3499 & w3514;
assign w3516 = ~w152 & ~w741;
assign w3517 = ~w16 & ~w166;
assign w3518 = ~w266 & ~w319;
assign w3519 = w715 & w2316;
assign w3520 = ~w30 & ~w164;
assign w3521 = ~w559 & ~w895;
assign w3522 = w3520 & w3521;
assign w3523 = w2416 & w3522;
assign w3524 = ~w349 & w646;
assign w3525 = w858 & w1491;
assign w3526 = w1562 & w1810;
assign w3527 = w3477 & w3516;
assign w3528 = w3517 & w3518;
assign w3529 = w3527 & w3528;
assign w3530 = w3525 & w3526;
assign w3531 = w1682 & w3524;
assign w3532 = w3103 & w3519;
assign w3533 = w3531 & w3532;
assign w3534 = w3529 & w3530;
assign w3535 = w3523 & w3534;
assign w3536 = w3487 & w3533;
assign w3537 = w3535 & w3536;
assign w3538 = w3180 & w3537;
assign w3539 = w3515 & w3538;
assign w3540 = ~w3403 & ~w3539;
assign w3541 = ~w3476 & ~w3540;
assign w3542 = ~w3326 & ~w3475;
assign w3543 = w3269 & w3326;
assign w3544 = (~w3268 & ~w3269) | (~w3268 & w32665) | (~w3269 & w32665);
assign w3545 = ~w3542 & ~w3544;
assign w3546 = w3541 & w3545;
assign w3547 = ~w3328 & w3546;
assign w3548 = w3403 & w3539;
assign w3549 = w3326 & w3475;
assign w3550 = w3403 & w3475;
assign w3551 = ~w3476 & ~w3550;
assign w3552 = ~w3549 & w3551;
assign w3553 = (~w3548 & w3552) | (~w3548 & w32666) | (w3552 & w32666);
assign w3554 = ~w2306 & ~w3539;
assign w3555 = w2306 & w3539;
assign w3556 = w2306 & w2393;
assign w3557 = ~w2394 & ~w3556;
assign w3558 = ~w3555 & w3557;
assign w3559 = (~w3547 & w32668) | (~w3547 & w32669) | (w32668 & w32669);
assign w3560 = ~w173 & ~w944;
assign w3561 = ~w116 & ~w142;
assign w3562 = ~w214 & ~w895;
assign w3563 = w3561 & w3562;
assign w3564 = w539 & ~w653;
assign w3565 = w3560 & w3564;
assign w3566 = w3563 & w3565;
assign w3567 = ~w403 & ~w562;
assign w3568 = ~w177 & ~w339;
assign w3569 = ~w60 & ~w188;
assign w3570 = ~w342 & ~w623;
assign w3571 = w3569 & w3570;
assign w3572 = ~w34 & ~w380;
assign w3573 = w289 & w3572;
assign w3574 = ~w252 & ~w266;
assign w3575 = ~w124 & ~w834;
assign w3576 = ~w212 & ~w290;
assign w3577 = ~w281 & w3574;
assign w3578 = w3575 & w3576;
assign w3579 = w3577 & w3578;
assign w3580 = w912 & w3480;
assign w3581 = w3579 & w3580;
assign w3582 = w2498 & w3581;
assign w3583 = ~w118 & ~w730;
assign w3584 = ~w345 & ~w541;
assign w3585 = ~w10 & ~w53;
assign w3586 = ~w75 & ~w163;
assign w3587 = ~w178 & ~w207;
assign w3588 = ~w1040 & w3587;
assign w3589 = w3585 & w3586;
assign w3590 = w466 & w1273;
assign w3591 = w3583 & w3584;
assign w3592 = w3590 & w3591;
assign w3593 = w3588 & w3589;
assign w3594 = w1642 & w2718;
assign w3595 = w3571 & w3573;
assign w3596 = w3594 & w3595;
assign w3597 = w3592 & w3593;
assign w3598 = w2973 & w3121;
assign w3599 = w3597 & w3598;
assign w3600 = w3596 & w3599;
assign w3601 = w3582 & w3600;
assign w3602 = ~w459 & w1009;
assign w3603 = ~w125 & ~w563;
assign w3604 = w1071 & w3603;
assign w3605 = w1118 & w1291;
assign w3606 = w3567 & w3568;
assign w3607 = w3605 & w3606;
assign w3608 = w872 & w3604;
assign w3609 = w3602 & w3608;
assign w3610 = w2514 & w3607;
assign w3611 = w3609 & w3610;
assign w3612 = w970 & w3566;
assign w3613 = w3611 & w3612;
assign w3614 = w3304 & w3613;
assign w3615 = w3601 & w3614;
assign w3616 = ~w2393 & ~w3615;
assign w3617 = ~w2075 & ~w3615;
assign w3618 = ~w3616 & ~w3617;
assign w3619 = w2148 & w2236;
assign w3620 = w2393 & w3615;
assign w3621 = w2074 & w2148;
assign w3622 = ~w2149 & ~w3621;
assign w3623 = w2075 & w3615;
assign w3624 = ~w3620 & ~w3623;
assign w3625 = w3622 & w3624;
assign w3626 = ~w3619 & w3625;
assign w3627 = ~w126 & ~w256;
assign w3628 = ~w380 & w1436;
assign w3629 = w3627 & w3628;
assign w3630 = ~w181 & ~w907;
assign w3631 = ~w140 & ~w1051;
assign w3632 = ~w118 & ~w123;
assign w3633 = ~w218 & w3632;
assign w3634 = ~w476 & w560;
assign w3635 = ~w283 & ~w385;
assign w3636 = ~w732 & w3635;
assign w3637 = w3274 & w3630;
assign w3638 = w3631 & w3637;
assign w3639 = w2683 & w3636;
assign w3640 = w3633 & w3634;
assign w3641 = w3639 & w3640;
assign w3642 = w881 & w3638;
assign w3643 = w3018 & w3642;
assign w3644 = w3487 & w3641;
assign w3645 = w3643 & w3644;
assign w3646 = w904 & w3645;
assign w3647 = ~w151 & ~w177;
assign w3648 = ~w242 & ~w446;
assign w3649 = ~w470 & ~w653;
assign w3650 = w3648 & w3649;
assign w3651 = w1551 & w3647;
assign w3652 = w3650 & w3651;
assign w3653 = w3238 & w3652;
assign w3654 = w2313 & w3629;
assign w3655 = w3653 & w3654;
assign w3656 = w864 & w3655;
assign w3657 = w2044 & w3656;
assign w3658 = w2526 & w3657;
assign w3659 = w3646 & w3658;
assign w3660 = ~w2006 & ~w3659;
assign w3661 = ~w153 & ~w292;
assign w3662 = ~w473 & w3661;
assign w3663 = ~w309 & ~w366;
assign w3664 = ~w16 & ~w39;
assign w3665 = ~w463 & ~w559;
assign w3666 = ~w597 & w3665;
assign w3667 = w2801 & w3664;
assign w3668 = w3663 & w3667;
assign w3669 = w1542 & w3666;
assign w3670 = w3066 & w3662;
assign w3671 = w3669 & w3670;
assign w3672 = w3668 & w3671;
assign w3673 = ~w337 & w1407;
assign w3674 = ~w156 & ~w531;
assign w3675 = ~w644 & ~w878;
assign w3676 = ~w388 & ~w895;
assign w3677 = ~w248 & ~w572;
assign w3678 = ~w378 & ~w475;
assign w3679 = ~w431 & w3141;
assign w3680 = w3677 & w3678;
assign w3681 = w3679 & w3680;
assign w3682 = ~w146 & ~w422;
assign w3683 = ~w619 & w3682;
assign w3684 = w584 & w3683;
assign w3685 = w1111 & w1205;
assign w3686 = ~w342 & ~w350;
assign w3687 = ~w167 & ~w1123;
assign w3688 = w697 & w3687;
assign w3689 = w754 & w1739;
assign w3690 = w2239 & w3686;
assign w3691 = w3689 & w3690;
assign w3692 = w1849 & w3688;
assign w3693 = w1865 & w2218;
assign w3694 = w3685 & w3693;
assign w3695 = w3691 & w3692;
assign w3696 = w2686 & w3629;
assign w3697 = w3695 & w3696;
assign w3698 = w1429 & w3694;
assign w3699 = w3697 & w3698;
assign w3700 = ~w476 & ~w540;
assign w3701 = ~w818 & w3700;
assign w3702 = w407 & w3674;
assign w3703 = w3675 & w3676;
assign w3704 = w3702 & w3703;
assign w3705 = w618 & w3701;
assign w3706 = w1812 & w3705;
assign w3707 = w3673 & w3704;
assign w3708 = w3681 & w3684;
assign w3709 = w3707 & w3708;
assign w3710 = w2022 & w3706;
assign w3711 = w3709 & w3710;
assign w3712 = w3672 & w3711;
assign w3713 = w3699 & w3712;
assign w3714 = ~w2236 & ~w3713;
assign w3715 = ~w3659 & ~w3713;
assign w3716 = ~w3714 & ~w3715;
assign w3717 = ~w3660 & w3716;
assign w3718 = w2236 & w3713;
assign w3719 = ~w3659 & ~w3718;
assign w3720 = w3659 & w3713;
assign w3721 = (~w2006 & ~w3659) | (~w2006 & w32676) | (~w3659 & w32676);
assign w3722 = ~w3719 & ~w3721;
assign w3723 = (w3559 & w32677) | (w3559 & w32678) | (w32677 & w32678);
assign w3724 = ~w1914 & ~w2006;
assign w3725 = ~w2007 & ~w3724;
assign w3726 = ~w3723 & w3725;
assign w3727 = (w3723 & w32680) | (w3723 & w32681) | (w32680 & w32681);
assign w3728 = ~w1715 & ~w1808;
assign w3729 = ~w1809 & ~w3728;
assign w3730 = ~w1915 & w3729;
assign w3731 = (~w3723 & w32682) | (~w3723 & w32683) | (w32682 & w32683);
assign w3732 = ~w98 & w2216;
assign w3733 = ~w355 & ~w470;
assign w3734 = ~w710 & ~w730;
assign w3735 = w3733 & w3734;
assign w3736 = ~w62 & ~w81;
assign w3737 = ~w896 & w1152;
assign w3738 = w1152 & w32686;
assign w3739 = ~w76 & ~w319;
assign w3740 = ~w146 & ~w191;
assign w3741 = ~w322 & ~w741;
assign w3742 = ~w815 & ~w1192;
assign w3743 = w3741 & w3742;
assign w3744 = w3740 & w3743;
assign w3745 = w651 & w3744;
assign w3746 = ~w323 & ~w389;
assign w3747 = ~w475 & w3746;
assign w3748 = w317 & w646;
assign w3749 = w1989 & w3169;
assign w3750 = w3736 & w3739;
assign w3751 = w3749 & w3750;
assign w3752 = w3747 & w3748;
assign w3753 = w2535 & w3633;
assign w3754 = w3732 & w3735;
assign w3755 = w3753 & w3754;
assign w3756 = w3751 & w3752;
assign w3757 = w3738 & w3756;
assign w3758 = w3745 & w3755;
assign w3759 = w3757 & w3758;
assign w3760 = w715 & w839;
assign w3761 = ~w208 & ~w282;
assign w3762 = w1109 & w3761;
assign w3763 = ~w242 & ~w701;
assign w3764 = ~w363 & ~w653;
assign w3765 = w775 & w3764;
assign w3766 = w3763 & w3765;
assign w3767 = w792 & w994;
assign w3768 = ~w217 & ~w476;
assign w3769 = ~w541 & w3768;
assign w3770 = ~w85 & ~w147;
assign w3771 = w1567 & w1663;
assign w3772 = ~w540 & ~w547;
assign w3773 = ~w56 & ~w708;
assign w3774 = w1418 & w3773;
assign w3775 = w1756 & ~w2885;
assign w3776 = w3772 & w3775;
assign w3777 = w3774 & w3776;
assign w3778 = ~w151 & ~w167;
assign w3779 = ~w252 & ~w288;
assign w3780 = w3778 & w3779;
assign w3781 = w407 & w1645;
assign w3782 = w2645 & w2943;
assign w3783 = w3770 & w3782;
assign w3784 = w3780 & w3781;
assign w3785 = w3771 & w3784;
assign w3786 = w3783 & w3785;
assign w3787 = w1959 & w3777;
assign w3788 = w3786 & w3787;
assign w3789 = ~w126 & ~w720;
assign w3790 = w343 & w3789;
assign w3791 = w1543 & w3790;
assign w3792 = w2799 & w3767;
assign w3793 = w3769 & w3792;
assign w3794 = w3791 & w3793;
assign w3795 = w3788 & w3794;
assign w3796 = ~w134 & ~w589;
assign w3797 = ~w350 & ~w392;
assign w3798 = ~w463 & w3797;
assign w3799 = ~w143 & ~w178;
assign w3800 = ~w278 & ~w992;
assign w3801 = w3799 & w3800;
assign w3802 = w941 & w1720;
assign w3803 = w3796 & w3802;
assign w3804 = w1835 & w3801;
assign w3805 = w2190 & w2770;
assign w3806 = w3760 & w3762;
assign w3807 = w3798 & w3806;
assign w3808 = w3804 & w3805;
assign w3809 = w3766 & w3803;
assign w3810 = w3808 & w3809;
assign w3811 = w3807 & w3810;
assign w3812 = w3759 & w3811;
assign w3813 = w3795 & w3812;
assign w3814 = ~w1808 & ~w3813;
assign w3815 = ~w1629 & ~w3813;
assign w3816 = ~w3814 & ~w3815;
assign w3817 = w1808 & w3813;
assign w3818 = w1629 & w3813;
assign w3819 = ~w3817 & ~w3818;
assign w3820 = w1523 & w1629;
assign w3821 = ~w1630 & ~w3820;
assign w3822 = (w3723 & w32691) | (w3723 & w32692) | (w32691 & w32692);
assign w3823 = ~w1475 & ~w1523;
assign w3824 = w1475 & w1523;
assign w3825 = w1397 & w1475;
assign w3826 = ~w1479 & ~w3825;
assign w3827 = ~w3824 & w3826;
assign w3828 = (w3827 & w3822) | (w3827 & w32694) | (w3822 & w32694);
assign w3829 = ~w1323 & ~w1397;
assign w3830 = w1323 & w1397;
assign w3831 = ~w3829 & ~w3830;
assign w3832 = (w3831 & w3828) | (w3831 & w32695) | (w3828 & w32695);
assign w3833 = ~w3828 & w32696;
assign w3834 = ~w3832 & ~w3833;
assign w3835 = ~w1324 & ~w1398;
assign w3836 = ~w1476 & w3835;
assign w3837 = (w3836 & ~w3834) | (w3836 & w32697) | (~w3834 & w32697);
assign w3838 = w1190 & ~w3837;
assign w3839 = w807 & ~w932;
assign w3840 = ~w933 & ~w3839;
assign w3841 = (~w3837 & w32699) | (~w3837 & w32700) | (w32699 & w32700);
assign w3842 = w574 & ~w710;
assign w3843 = w792 & w837;
assign w3844 = w1865 & w3842;
assign w3845 = w3843 & w3844;
assign w3846 = ~w46 & w728;
assign w3847 = ~w127 & ~w385;
assign w3848 = w3846 & w3847;
assign w3849 = w1372 & w32703;
assign w3850 = w268 & w2216;
assign w3851 = w2337 & w3119;
assign w3852 = w3369 & w3851;
assign w3853 = w3850 & w3852;
assign w3854 = w3845 & w3853;
assign w3855 = w1248 & w3854;
assign w3856 = w3855 & w32704;
assign w3857 = w3849 & w3856;
assign w3858 = ~w815 & w3857;
assign w3859 = ~w932 & ~w3858;
assign w3860 = w932 & w3857;
assign w3861 = (a_29 & w3859) | (a_29 & w32705) | (w3859 & w32705);
assign w3862 = ~w3859 & w32706;
assign w3863 = ~w3861 & ~w3862;
assign w3864 = (w3837 & w32707) | (w3837 & w32708) | (w32707 & w32708);
assign w3865 = (~w3837 & w32709) | (~w3837 & w32710) | (w32709 & w32710);
assign w3866 = ~w3864 & ~w3865;
assign w3867 = ~w127 & w2941;
assign w3868 = ~w316 & w1536;
assign w3869 = ~w593 & w3574;
assign w3870 = ~w400 & w2191;
assign w3871 = w2709 & w3870;
assign w3872 = w1290 & w3842;
assign w3873 = w3867 & w3868;
assign w3874 = w3869 & w3873;
assign w3875 = w3871 & w3872;
assign w3876 = w3874 & w3875;
assign w3877 = w340 & ~w2331;
assign w3878 = ~w138 & ~w365;
assign w3879 = ~w589 & ~w1043;
assign w3880 = w3878 & w3879;
assign w3881 = w1312 & w3880;
assign w3882 = w2123 & w3877;
assign w3883 = w3881 & w3882;
assign w3884 = ~w10 & w2033;
assign w3885 = w1214 & w3884;
assign w3886 = w3883 & w3885;
assign w3887 = w2987 & w3886;
assign w3888 = a_26 & w87;
assign w3889 = ~w4 & ~w21;
assign w3890 = w1222 & w3889;
assign w3891 = w3888 & ~w3890;
assign w3892 = ~w156 & ~w623;
assign w3893 = ~w423 & ~w671;
assign w3894 = ~w56 & w257;
assign w3895 = w986 & w3892;
assign w3896 = w3893 & w3895;
assign w3897 = w716 & w3894;
assign w3898 = w1771 & w3897;
assign w3899 = w3896 & w3898;
assign w3900 = w3898 & w32711;
assign w3901 = w516 & w3843;
assign w3902 = w3900 & w3901;
assign w3903 = w3887 & w3902;
assign w3904 = w3887 & w32712;
assign w3905 = ~w290 & w3876;
assign w3906 = w3904 & w3905;
assign w3907 = (w1327 & ~w3904) | (w1327 & w32713) | (~w3904 & w32713);
assign w3908 = (w1399 & ~w1308) | (w1399 & w32714) | (~w1308 & w32714);
assign w3909 = ~w290 & ~w1228;
assign w3910 = ~w45 & ~w531;
assign w3911 = ~w282 & ~w463;
assign w3912 = ~w907 & w3155;
assign w3913 = w3910 & w3911;
assign w3914 = w3912 & w3913;
assign w3915 = ~w39 & ~w177;
assign w3916 = ~w85 & ~w341;
assign w3917 = ~w46 & w570;
assign w3918 = ~w737 & ~w1336;
assign w3919 = ~w1953 & w3918;
assign w3920 = w3014 & w3456;
assign w3921 = w3916 & w3920;
assign w3922 = w3917 & w3919;
assign w3923 = w3921 & w3922;
assign w3924 = ~w356 & w1464;
assign w3925 = ~w647 & ~w734;
assign w3926 = ~w2049 & w3925;
assign w3927 = w1632 & w3092;
assign w3928 = w3915 & w3927;
assign w3929 = w3924 & w3926;
assign w3930 = w3928 & w3929;
assign w3931 = w3914 & w3930;
assign w3932 = w3923 & w3931;
assign w3933 = w3931 & w32715;
assign w3934 = w3909 & w3933;
assign w3935 = w3904 & w32716;
assign w3936 = w3904 & ~w3935;
assign w3937 = ~w1323 & ~w3906;
assign w3938 = w1323 & w3906;
assign w3939 = ~w3937 & ~w3938;
assign w3940 = (w3828 & w32719) | (w3828 & w32720) | (w32719 & w32720);
assign w3941 = (w3828 & w32723) | (w3828 & w32724) | (w32723 & w32724);
assign w3942 = (~w3828 & w32725) | (~w3828 & w32726) | (w32725 & w32726);
assign w3943 = ~w3941 & ~w3942;
assign w3944 = ~w3907 & ~w3908;
assign w3945 = (w3944 & ~w3943) | (w3944 & w32727) | (~w3943 & w32727);
assign w3946 = w3866 & ~w3945;
assign w3947 = ~w3866 & w3945;
assign w3948 = ~w3946 & ~w3947;
assign w3949 = ~a_28 & a_29;
assign w3950 = a_28 & ~a_29;
assign w3951 = ~w3949 & ~w3950;
assign w3952 = ~a_26 & ~a_27;
assign w3953 = a_26 & a_27;
assign w3954 = ~w3952 & ~w3953;
assign w3955 = ~w7 & ~w31;
assign w3956 = ~w3954 & ~w3955;
assign w3957 = ~w3951 & w3956;
assign w3958 = w3933 & w32728;
assign w3959 = (~a_29 & w3958) | (~a_29 & w32729) | (w3958 & w32729);
assign w3960 = ~w1323 & w1327;
assign w3961 = (w668 & ~w3904) | (w668 & w32730) | (~w3904 & w32730);
assign w3962 = ~w1397 & w1399;
assign w3963 = (~w3828 & w32731) | (~w3828 & w32732) | (w32731 & w32732);
assign w3964 = ~w3940 & ~w3963;
assign w3965 = w1478 & w3964;
assign w3966 = ~w3960 & w32733;
assign w3967 = ~w3965 & w32734;
assign w3968 = (w3837 & w32735) | (w3837 & w32736) | (w32735 & w32736);
assign w3969 = ~w3841 & ~w3968;
assign w3970 = (~w3959 & w3965) | (~w3959 & w32737) | (w3965 & w32737);
assign w3971 = ~w3967 & ~w3970;
assign w3972 = ~w3969 & w3971;
assign w3973 = ~w3967 & ~w3972;
assign w3974 = w3948 & w3973;
assign w3975 = ~w3948 & ~w3973;
assign w3976 = ~w3974 & ~w3975;
assign w3977 = ~w208 & w1966;
assign w3978 = ~w568 & ~w1117;
assign w3979 = ~w195 & ~w356;
assign w3980 = ~w152 & ~w619;
assign w3981 = w792 & w3980;
assign w3982 = w2276 & w2717;
assign w3983 = w3014 & w3978;
assign w3984 = w3979 & w3983;
assign w3985 = w3981 & w3982;
assign w3986 = w1852 & w3977;
assign w3987 = w3985 & w3986;
assign w3988 = w3984 & w3987;
assign w3989 = ~w251 & ~w429;
assign w3990 = w73 & w3989;
assign w3991 = w1251 & w3990;
assign w3992 = w791 & ~w907;
assign w3993 = w171 & ~w191;
assign w3994 = w581 & w1198;
assign w3995 = w2872 & w3102;
assign w3996 = w3994 & w3995;
assign w3997 = w3992 & w3993;
assign w3998 = w3996 & w3997;
assign w3999 = w1940 & w32738;
assign w4000 = ~w531 & w1309;
assign w4001 = w122 & w1288;
assign w4002 = ~w261 & w1074;
assign w4003 = ~w62 & ~w75;
assign w4004 = ~w394 & w4003;
assign w4005 = w739 & w1229;
assign w4006 = w4004 & w4005;
assign w4007 = w70 & w4006;
assign w4008 = ~w278 & ~w389;
assign w4009 = ~w50 & ~w400;
assign w4010 = ~w56 & ~w220;
assign w4011 = ~w365 & ~w369;
assign w4012 = ~w696 & ~w4001;
assign w4013 = w4011 & w4012;
assign w4014 = w743 & w4010;
assign w4015 = w1075 & w1343;
assign w4016 = w1665 & w2485;
assign w4017 = w2871 & w2965;
assign w4018 = w4008 & w4009;
assign w4019 = w4017 & w4018;
assign w4020 = w4015 & w4016;
assign w4021 = w4013 & w4014;
assign w4022 = w2086 & w4000;
assign w4023 = w4002 & w4022;
assign w4024 = w4020 & w4021;
assign w4025 = w955 & w4019;
assign w4026 = w3991 & w4025;
assign w4027 = w4023 & w4024;
assign w4028 = w4007 & w4027;
assign w4029 = w3988 & w4026;
assign w4030 = w4028 & w4029;
assign w4031 = w3999 & w4030;
assign w4032 = w1068 & ~w4031;
assign w4033 = ~w1068 & w4031;
assign w4034 = ~w4032 & ~w4033;
assign w4035 = w668 & ~w1475;
assign w4036 = (w1399 & ~w1628) | (w1399 & w32739) | (~w1628 & w32739);
assign w4037 = (w1327 & ~w643) | (w1327 & w32740) | (~w643 & w32740);
assign w4038 = ~w3823 & ~w3824;
assign w4039 = (w4038 & w3822) | (w4038 & w32741) | (w3822 & w32741);
assign w4040 = ~w3822 & w32742;
assign w4041 = ~w4039 & ~w4040;
assign w4042 = ~w4036 & ~w4037;
assign w4043 = ~w4035 & w4042;
assign w4044 = (w4043 & ~w4041) | (w4043 & w32743) | (~w4041 & w32743);
assign w4045 = w4034 & ~w4044;
assign w4046 = a_26 & ~w1185;
assign w4047 = ~w1186 & ~w4046;
assign w4048 = (~w4044 & w32745) | (~w4044 & w32746) | (w32745 & w32746);
assign w4049 = (w4044 & w32747) | (w4044 & w32748) | (w32747 & w32748);
assign w4050 = ~w4048 & ~w4049;
assign w4051 = w668 & ~w1397;
assign w4052 = w1327 & ~w1475;
assign w4053 = (w1399 & ~w643) | (w1399 & w32749) | (~w643 & w32749);
assign w4054 = ~w3823 & ~w3826;
assign w4055 = (~w3822 & w32750) | (~w3822 & w32751) | (w32750 & w32751);
assign w4056 = ~w3828 & ~w4055;
assign w4057 = ~w4051 & ~w4053;
assign w4058 = ~w4052 & w4057;
assign w4059 = (w4058 & ~w4056) | (w4058 & w32752) | (~w4056 & w32752);
assign w4060 = w4050 & ~w4059;
assign w4061 = (~w4048 & ~w4050) | (~w4048 & w32753) | (~w4050 & w32753);
assign w4062 = (~w3834 & w32754) | (~w3834 & w32755) | (w32754 & w32755);
assign w4063 = ~w3838 & ~w4062;
assign w4064 = ~w4061 & w4063;
assign w4065 = w4061 & ~w4063;
assign w4066 = ~w4064 & ~w4065;
assign w4067 = (w3957 & ~w3904) | (w3957 & w32756) | (~w3904 & w32756);
assign w4068 = ~w3954 & w3955;
assign w4069 = ~w3958 & w4068;
assign w4070 = ~w3951 & w3954;
assign w4071 = (w3828 & w32759) | (w3828 & w32760) | (w32759 & w32760);
assign w4072 = (~w3828 & w32761) | (~w3828 & w32762) | (w32761 & w32762);
assign w4073 = ~w4071 & ~w4072;
assign w4074 = ~w4067 & ~w4069;
assign w4075 = (w4074 & ~w4073) | (w4074 & w32763) | (~w4073 & w32763);
assign w4076 = ~a_29 & w4075;
assign w4077 = (w4073 & w32764) | (w4073 & w32765) | (w32764 & w32765);
assign w4078 = ~w4076 & ~w4077;
assign w4079 = w4066 & w4078;
assign w4080 = (~w4064 & ~w4066) | (~w4064 & w32766) | (~w4066 & w32766);
assign w4081 = w3969 & ~w3971;
assign w4082 = ~w3972 & ~w4081;
assign w4083 = ~w4080 & ~w4082;
assign w4084 = ~w186 & ~w208;
assign w4085 = ~w341 & ~w388;
assign w4086 = ~w112 & w4085;
assign w4087 = w4084 & w4086;
assign w4088 = ~w597 & ~w996;
assign w4089 = ~w279 & ~w538;
assign w4090 = ~w1123 & w3247;
assign w4091 = w4088 & w4089;
assign w4092 = w4090 & w4091;
assign w4093 = ~w197 & ~w626;
assign w4094 = ~w140 & ~w737;
assign w4095 = ~w190 & ~w473;
assign w4096 = ~w895 & w4095;
assign w4097 = w1116 & w1738;
assign w4098 = w1920 & w4093;
assign w4099 = w4094 & w4098;
assign w4100 = w4096 & w4097;
assign w4101 = w2380 & w3735;
assign w4102 = w4100 & w4101;
assign w4103 = w4099 & w4102;
assign w4104 = ~w67 & ~w283;
assign w4105 = ~w71 & ~w447;
assign w4106 = ~w450 & ~w720;
assign w4107 = w4105 & w4106;
assign w4108 = w957 & w3736;
assign w4109 = w4104 & w4108;
assign w4110 = w4107 & w4109;
assign w4111 = ~w10 & ~w671;
assign w4112 = ~w125 & ~w256;
assign w4113 = w1100 & w4112;
assign w4114 = w4111 & w4113;
assign w4115 = w4000 & w4114;
assign w4116 = ~w45 & ~w135;
assign w4117 = ~w350 & ~w468;
assign w4118 = ~w708 & w4117;
assign w4119 = w1640 & w4116;
assign w4120 = w2440 & w3404;
assign w4121 = w4119 & w4120;
assign w4122 = w4118 & w4121;
assign w4123 = w2651 & w4122;
assign w4124 = w4110 & w4115;
assign w4125 = w4123 & w4124;
assign w4126 = w4103 & w4125;
assign w4127 = ~w126 & ~w385;
assign w4128 = ~w701 & ~w789;
assign w4129 = w2250 & w4128;
assign w4130 = ~w776 & w949;
assign w4131 = ~w156 & ~w400;
assign w4132 = ~w562 & w4131;
assign w4133 = w2216 & w2800;
assign w4134 = w3978 & w4127;
assign w4135 = w4133 & w4134;
assign w4136 = w2482 & w4132;
assign w4137 = w4129 & w4130;
assign w4138 = w4136 & w4137;
assign w4139 = w4087 & w4135;
assign w4140 = w4092 & w4139;
assign w4141 = w3293 & w4138;
assign w4142 = w4140 & w4141;
assign w4143 = w4126 & w4142;
assign w4144 = w654 & w673;
assign w4145 = w1431 & w4144;
assign w4146 = ~w128 & ~w392;
assign w4147 = w311 & w4146;
assign w4148 = w836 & w4147;
assign w4149 = w286 & w4148;
assign w4150 = w4145 & w4149;
assign w4151 = ~w115 & ~w143;
assign w4152 = ~w135 & ~w649;
assign w4153 = w733 & w1292;
assign w4154 = w1950 & w2101;
assign w4155 = w4153 & w4154;
assign w4156 = ~w126 & w1680;
assign w4157 = ~w72 & ~w164;
assign w4158 = ~w459 & ~w1117;
assign w4159 = ~w208 & ~w394;
assign w4160 = ~w65 & w4159;
assign w4161 = ~w125 & ~w188;
assign w4162 = ~w710 & w4161;
assign w4163 = ~w16 & ~w127;
assign w4164 = ~w337 & ~w563;
assign w4165 = w421 & w4164;
assign w4166 = w617 & w998;
assign w4167 = w1124 & w2442;
assign w4168 = w4157 & w4158;
assign w4169 = w4163 & w4168;
assign w4170 = w4166 & w4167;
assign w4171 = w1008 & w4165;
assign w4172 = w4160 & w4162;
assign w4173 = w4171 & w4172;
assign w4174 = w4169 & w4170;
assign w4175 = w1570 & w4174;
assign w4176 = w4173 & w4175;
assign w4177 = ~w173 & ~w251;
assign w4178 = w449 & w4177;
assign w4179 = w728 & w1081;
assign w4180 = w1718 & w2502;
assign w4181 = w2579 & w3575;
assign w4182 = w4180 & w4181;
assign w4183 = w4178 & w4179;
assign w4184 = w4156 & w4183;
assign w4185 = w1156 & w4182;
assign w4186 = w1780 & w4155;
assign w4187 = w4185 & w4186;
assign w4188 = w2246 & w4184;
assign w4189 = w4187 & w4188;
assign w4190 = w4176 & w4189;
assign w4191 = ~w423 & ~w541;
assign w4192 = w24 & w4191;
assign w4193 = w735 & w819;
assign w4194 = w3330 & w4193;
assign w4195 = w4192 & w4194;
assign w4196 = ~w183 & ~w248;
assign w4197 = ~w473 & ~w530;
assign w4198 = w4196 & w4197;
assign w4199 = ~w147 & ~w447;
assign w4200 = w1638 & w4199;
assign w4201 = w3123 & w3167;
assign w4202 = w4093 & w4151;
assign w4203 = w4152 & w4202;
assign w4204 = w4200 & w4201;
assign w4205 = w898 & w4198;
assign w4206 = w4204 & w4205;
assign w4207 = w2085 & w4203;
assign w4208 = w4206 & w4207;
assign w4209 = w4195 & w4208;
assign w4210 = w4150 & w4209;
assign w4211 = w4190 & w4210;
assign w4212 = ~w4143 & ~w4211;
assign w4213 = w4143 & w4211;
assign w4214 = ~w4212 & ~w4213;
assign w4215 = ~a_23 & w4214;
assign w4216 = (~w4212 & ~w4214) | (~w4212 & w32767) | (~w4214 & w32767);
assign w4217 = w1068 & ~w4216;
assign w4218 = ~w1068 & w4216;
assign w4219 = ~w4217 & ~w4218;
assign w4220 = w1399 & ~w3813;
assign w4221 = (w668 & ~w643) | (w668 & w32768) | (~w643 & w32768);
assign w4222 = (w1327 & ~w1628) | (w1327 & w32769) | (~w1628 & w32769);
assign w4223 = (~w3723 & w32770) | (~w3723 & w32771) | (w32770 & w32771);
assign w4224 = ~w3822 & ~w4223;
assign w4225 = w1478 & w4224;
assign w4226 = ~w4220 & w32772;
assign w4227 = (w4219 & w4225) | (w4219 & w32773) | (w4225 & w32773);
assign w4228 = (~w4225 & w32774) | (~w4225 & w32775) | (w32774 & w32775);
assign w4229 = (~w4041 & w32776) | (~w4041 & w32777) | (w32776 & w32777);
assign w4230 = ~w4045 & w32778;
assign w4231 = (w4228 & w4045) | (w4228 & w32779) | (w4045 & w32779);
assign w4232 = ~w4230 & ~w4231;
assign w4233 = a_23 & ~w4214;
assign w4234 = ~w4215 & ~w4233;
assign w4235 = w1327 & ~w3813;
assign w4236 = (w668 & ~w1628) | (w668 & w32780) | (~w1628 & w32780);
assign w4237 = (w1399 & ~w1807) | (w1399 & w32781) | (~w1807 & w32781);
assign w4238 = (w3723 & w32782) | (w3723 & w32783) | (w32782 & w32783);
assign w4239 = ~w3814 & ~w3817;
assign w4240 = (w3723 & w32784) | (w3723 & w32785) | (w32784 & w32785);
assign w4241 = ~w3815 & ~w3818;
assign w4242 = ~w3814 & ~w4241;
assign w4243 = (~w3723 & w32786) | (~w3723 & w32787) | (w32786 & w32787);
assign w4244 = ~w4238 & ~w4243;
assign w4245 = w1478 & w4244;
assign w4246 = ~w4235 & w32788;
assign w4247 = (w4234 & w4245) | (w4234 & w32789) | (w4245 & w32789);
assign w4248 = ~w159 & ~w394;
assign w4249 = ~w186 & w4248;
assign w4250 = w2016 & w2439;
assign w4251 = w2495 & w4250;
assign w4252 = w4249 & w4251;
assign w4253 = ~w50 & w3101;
assign w4254 = ~w157 & ~w719;
assign w4255 = ~w350 & ~w429;
assign w4256 = w57 & ~w123;
assign w4257 = ~w279 & ~w626;
assign w4258 = ~w136 & w721;
assign w4259 = w813 & w4257;
assign w4260 = w4258 & w4259;
assign w4261 = w1121 & w4260;
assign w4262 = w448 & w1344;
assign w4263 = w1400 & w2515;
assign w4264 = w4254 & w4255;
assign w4265 = w4263 & w4264;
assign w4266 = w3420 & w4262;
assign w4267 = w4253 & w4256;
assign w4268 = w4266 & w4267;
assign w4269 = w4265 & w4268;
assign w4270 = w4261 & w4269;
assign w4271 = ~w1040 & w1340;
assign w4272 = ~w399 & ~w714;
assign w4273 = w4271 & w4272;
assign w4274 = ~w239 & ~w732;
assign w4275 = ~w143 & ~w256;
assign w4276 = ~w266 & ~w342;
assign w4277 = w1125 & w4276;
assign w4278 = w2332 & w2730;
assign w4279 = w4274 & w4275;
assign w4280 = w4278 & w4279;
assign w4281 = w1110 & w4277;
assign w4282 = w1849 & w4281;
assign w4283 = w4273 & w4280;
assign w4284 = w4282 & w4283;
assign w4285 = w4252 & w4284;
assign w4286 = w3672 & w4285;
assign w4287 = w2901 & w4270;
assign w4288 = w4286 & w4287;
assign w4289 = w4143 & ~w4288;
assign w4290 = ~w16 & ~w178;
assign w4291 = ~w314 & ~w399;
assign w4292 = w4290 & w4291;
assign w4293 = w733 & w2874;
assign w4294 = w3030 & w4293;
assign w4295 = w4130 & w4292;
assign w4296 = w4294 & w4295;
assign w4297 = ~w186 & ~w653;
assign w4298 = ~w166 & ~w246;
assign w4299 = w988 & w1010;
assign w4300 = w1374 & w2280;
assign w4301 = w2420 & w2495;
assign w4302 = w2966 & w3464;
assign w4303 = w4298 & w4302;
assign w4304 = w4300 & w4301;
assign w4305 = w4297 & w4299;
assign w4306 = w4304 & w4305;
assign w4307 = w4303 & w4306;
assign w4308 = w3312 & w4296;
assign w4309 = w4307 & w4308;
assign w4310 = w1153 & w32790;
assign w4311 = ~w95 & w3419;
assign w4312 = ~w85 & ~w169;
assign w4313 = ~w538 & ~w737;
assign w4314 = ~w1104 & w4313;
assign w4315 = ~w194 & w4312;
assign w4316 = w4314 & w4315;
assign w4317 = w148 & ~w385;
assign w4318 = w2121 & w2361;
assign w4319 = w4317 & w4318;
assign w4320 = w793 & w3059;
assign w4321 = w3284 & w4311;
assign w4322 = w4320 & w4321;
assign w4323 = w2435 & w4319;
assign w4324 = w4310 & w4316;
assign w4325 = w4323 & w4324;
assign w4326 = w4322 & w4325;
assign w4327 = w1860 & w3686;
assign w4328 = ~w288 & ~w349;
assign w4329 = w947 & w4328;
assign w4330 = ~w18 & ~w128;
assign w4331 = ~w458 & ~w597;
assign w4332 = w4330 & w4331;
assign w4333 = w817 & w1987;
assign w4334 = w2886 & w4333;
assign w4335 = w1239 & w4332;
assign w4336 = w2580 & w4327;
assign w4337 = w4329 & w4336;
assign w4338 = w4334 & w4335;
assign w4339 = w4337 & w4338;
assign w4340 = w2081 & w4339;
assign w4341 = w2261 & w4340;
assign w4342 = w4309 & w4326;
assign w4343 = w4341 & w4342;
assign w4344 = ~w313 & w1111;
assign w4345 = w911 & w1776;
assign w4346 = ~w83 & ~w124;
assign w4347 = w1361 & w1418;
assign w4348 = w2515 & w2527;
assign w4349 = w3100 & w4346;
assign w4350 = w4348 & w4349;
assign w4351 = w3017 & w4347;
assign w4352 = w4350 & w4351;
assign w4353 = ~w169 & ~w418;
assign w4354 = ~w475 & w4353;
assign w4355 = w1103 & w2873;
assign w4356 = w3154 & w3274;
assign w4357 = w4355 & w4356;
assign w4358 = w4344 & w4345;
assign w4359 = w4354 & w4358;
assign w4360 = w4357 & w4359;
assign w4361 = w2285 & w4352;
assign w4362 = w4360 & w4361;
assign w4363 = ~w221 & ~w238;
assign w4364 = ~w116 & ~w447;
assign w4365 = w876 & w3763;
assign w4366 = ~w369 & w4152;
assign w4367 = w139 & w1952;
assign w4368 = ~w393 & ~w572;
assign w4369 = ~w292 & ~w4367;
assign w4370 = w250 & w4369;
assign w4371 = w4368 & w4370;
assign w4372 = w433 & ~w1965;
assign w4373 = w1125 & w2008;
assign w4374 = w2087 & w3208;
assign w4375 = w3663 & w4328;
assign w4376 = w4363 & w4364;
assign w4377 = w4375 & w4376;
assign w4378 = w4373 & w4374;
assign w4379 = w4271 & w4372;
assign w4380 = w4365 & w4366;
assign w4381 = w4379 & w4380;
assign w4382 = w4377 & w4378;
assign w4383 = w4371 & w4382;
assign w4384 = w4381 & w4383;
assign w4385 = ~w45 & ~w559;
assign w4386 = ~w246 & ~w696;
assign w4387 = ~w278 & w2278;
assign w4388 = ~w191 & w1205;
assign w4389 = w2689 & w4385;
assign w4390 = w4386 & w4389;
assign w4391 = w4387 & w4388;
assign w4392 = w4390 & w4391;
assign w4393 = ~w76 & ~w237;
assign w4394 = ~w113 & ~w161;
assign w4395 = ~w446 & ~w644;
assign w4396 = ~w741 & w4395;
assign w4397 = w219 & w4394;
assign w4398 = w1329 & w2161;
assign w4399 = w3892 & w4393;
assign w4400 = w4398 & w4399;
assign w4401 = w4396 & w4397;
assign w4402 = w4400 & w4401;
assign w4403 = ~w1222 & w1224;
assign w4404 = w9 & w4403;
assign w4405 = w773 & w1562;
assign w4406 = w1689 & w2781;
assign w4407 = w3736 & ~w4404;
assign w4408 = w4406 & w4407;
assign w4409 = w2847 & w4405;
assign w4410 = w4408 & w4409;
assign w4411 = w1486 & w4410;
assign w4412 = w4392 & w4402;
assign w4413 = w4411 & w4412;
assign w4414 = w4362 & w4413;
assign w4415 = w4384 & w4414;
assign w4416 = ~w4343 & ~w4415;
assign w4417 = w4343 & w4415;
assign w4418 = ~w4416 & ~w4417;
assign w4419 = ~a_20 & w4418;
assign w4420 = (~w4416 & ~w4418) | (~w4416 & w32791) | (~w4418 & w32791);
assign w4421 = w4288 & ~w4420;
assign w4422 = ~w4288 & w4420;
assign w4423 = ~w4421 & ~w4422;
assign w4424 = (w1399 & ~w1913) | (w1399 & w32792) | (~w1913 & w32792);
assign w4425 = (w1327 & ~w1714) | (w1327 & w32769) | (~w1714 & w32769);
assign w4426 = (w668 & ~w1807) | (w668 & w32793) | (~w1807 & w32793);
assign w4427 = (w3723 & w32796) | (w3723 & w32797) | (w32796 & w32797);
assign w4428 = ~w3731 & ~w4427;
assign w4429 = ~w4424 & ~w4425;
assign w4430 = ~w4426 & w4429;
assign w4431 = (w4430 & w4428) | (w4430 & w32798) | (w4428 & w32798);
assign w4432 = w4423 & ~w4431;
assign w4433 = ~w4143 & w4288;
assign w4434 = ~w4289 & ~w4433;
assign w4435 = (~w4431 & w32800) | (~w4431 & w32801) | (w32800 & w32801);
assign w4436 = (w4431 & w32802) | (w4431 & w32803) | (w32802 & w32803);
assign w4437 = ~w4245 & w32804;
assign w4438 = ~w4247 & ~w4437;
assign w4439 = ~w4436 & w4438;
assign w4440 = (~w4247 & ~w4438) | (~w4247 & w32805) | (~w4438 & w32805);
assign w4441 = ~w4225 & w32806;
assign w4442 = ~w4227 & ~w4441;
assign w4443 = ~w4440 & w4442;
assign w4444 = w4440 & ~w4442;
assign w4445 = ~w4443 & ~w4444;
assign w4446 = w3951 & w3954;
assign w4447 = (w4446 & ~w1308) | (w4446 & w32807) | (~w1308 & w32807);
assign w4448 = ~w1397 & w4068;
assign w4449 = ~w1475 & w3957;
assign w4450 = ~w4447 & ~w4448;
assign w4451 = ~w4449 & w4450;
assign w4452 = (w4451 & ~w3834) | (w4451 & w32808) | (~w3834 & w32808);
assign w4453 = ~a_29 & w4452;
assign w4454 = (w3834 & w32809) | (w3834 & w32810) | (w32809 & w32810);
assign w4455 = ~w4453 & ~w4454;
assign w4456 = w4445 & w4455;
assign w4457 = (~w4443 & ~w4445) | (~w4443 & w32811) | (~w4445 & w32811);
assign w4458 = w4232 & ~w4457;
assign w4459 = ~w4050 & w4059;
assign w4460 = ~w4060 & ~w4459;
assign w4461 = (~w4457 & w32813) | (~w4457 & w32814) | (w32813 & w32814);
assign w4462 = (w4457 & w32815) | (w4457 & w32816) | (w32815 & w32816);
assign w4463 = ~w4461 & ~w4462;
assign w4464 = (w4068 & ~w3904) | (w4068 & w32817) | (~w3904 & w32817);
assign w4465 = ~w3958 & w4446;
assign w4466 = (w3957 & ~w1308) | (w3957 & w32818) | (~w1308 & w32818);
assign w4467 = ~w4465 & ~w4466;
assign w4468 = ~w4464 & w4467;
assign w4469 = (w4468 & ~w3943) | (w4468 & w32819) | (~w3943 & w32819);
assign w4470 = a_29 & ~w4469;
assign w4471 = (~w3943 & w32820) | (~w3943 & w32821) | (w32820 & w32821);
assign w4472 = ~w4470 & ~w4471;
assign w4473 = w4463 & w4472;
assign w4474 = (~w4461 & ~w4463) | (~w4461 & w32822) | (~w4463 & w32822);
assign w4475 = ~w4066 & ~w4078;
assign w4476 = ~w4079 & ~w4475;
assign w4477 = ~w4474 & w4476;
assign w4478 = (w4068 & ~w1308) | (w4068 & w32823) | (~w1308 & w32823);
assign w4479 = (w4446 & ~w3904) | (w4446 & w32824) | (~w3904 & w32824);
assign w4480 = ~w1397 & w3957;
assign w4481 = ~w4478 & ~w4480;
assign w4482 = ~w4479 & w4481;
assign w4483 = (w4482 & ~w3964) | (w4482 & w32825) | (~w3964 & w32825);
assign w4484 = a_29 & ~w4483;
assign w4485 = (~w3964 & w32826) | (~w3964 & w32827) | (w32826 & w32827);
assign w4486 = (~w3828 & w32830) | (~w3828 & w32831) | (w32830 & w32831);
assign w4487 = ~w4486 & w32832;
assign w4488 = (a_26 & w4486) | (a_26 & w32833) | (w4486 & w32833);
assign w4489 = ~w4487 & ~w4488;
assign w4490 = ~w4484 & w32834;
assign w4491 = ~w4232 & w4457;
assign w4492 = ~w4458 & ~w4491;
assign w4493 = (w4489 & w4484) | (w4489 & w32835) | (w4484 & w32835);
assign w4494 = ~w4490 & ~w4493;
assign w4495 = w4492 & w4494;
assign w4496 = (~w4490 & ~w4492) | (~w4490 & w32836) | (~w4492 & w32836);
assign w4497 = ~w4463 & ~w4472;
assign w4498 = ~w4473 & ~w4497;
assign w4499 = ~w4496 & w4498;
assign w4500 = w4496 & ~w4498;
assign w4501 = ~w4499 & ~w4500;
assign w4502 = (w4431 & w32837) | (w4431 & w32838) | (w32837 & w32838);
assign w4503 = ~w4435 & ~w4502;
assign w4504 = (w1327 & ~w1807) | (w1327 & w32839) | (~w1807 & w32839);
assign w4505 = (w1399 & ~w1714) | (w1399 & w32739) | (~w1714 & w32739);
assign w4506 = w668 & ~w3813;
assign w4507 = (~w3723 & w32840) | (~w3723 & w32841) | (w32840 & w32841);
assign w4508 = ~w4240 & ~w4507;
assign w4509 = ~w4504 & ~w4505;
assign w4510 = ~w4506 & w4509;
assign w4511 = (w4510 & ~w4508) | (w4510 & w32842) | (~w4508 & w32842);
assign w4512 = w4503 & ~w4511;
assign w4513 = ~w582 & w2122;
assign w4514 = w346 & w2087;
assign w4515 = ~w34 & ~w447;
assign w4516 = ~w563 & ~w619;
assign w4517 = ~w992 & w4516;
assign w4518 = w398 & w4515;
assign w4519 = w2419 & w4518;
assign w4520 = w4517 & w4519;
assign w4521 = ~w256 & ~w385;
assign w4522 = ~w446 & ~w473;
assign w4523 = ~w309 & ~w647;
assign w4524 = w2308 & w4523;
assign w4525 = ~w869 & ~w1077;
assign w4526 = w1865 & w4525;
assign w4527 = ~w123 & w424;
assign w4528 = w2193 & w4521;
assign w4529 = w4522 & w4528;
assign w4530 = w558 & w4527;
assign w4531 = w854 & w1728;
assign w4532 = w4514 & w4531;
assign w4533 = w4529 & w4530;
assign w4534 = w4524 & w4526;
assign w4535 = w4533 & w4534;
assign w4536 = w4520 & w4532;
assign w4537 = w4535 & w4536;
assign w4538 = ~w186 & w4537;
assign w4539 = ~w196 & ~w251;
assign w4540 = ~w178 & ~w195;
assign w4541 = w2019 & w4540;
assign w4542 = w3634 & w4541;
assign w4543 = ~w312 & w938;
assign w4544 = ~w151 & ~w815;
assign w4545 = w1861 & w2511;
assign w4546 = w3386 & w4544;
assign w4547 = w4545 & w4546;
assign w4548 = w1810 & w3274;
assign w4549 = ~w1117 & w4539;
assign w4550 = w676 & w4549;
assign w4551 = w2262 & w3685;
assign w4552 = w3762 & w4543;
assign w4553 = w4548 & w4552;
assign w4554 = w4550 & w4551;
assign w4555 = w4542 & w4547;
assign w4556 = w4554 & w4555;
assign w4557 = w4553 & w4556;
assign w4558 = ~w62 & ~w395;
assign w4559 = ~w734 & w4558;
assign w4560 = w317 & w1125;
assign w4561 = w2101 & w4094;
assign w4562 = w4560 & w4561;
assign w4563 = w4513 & w4559;
assign w4564 = w4562 & w4563;
assign w4565 = w1864 & w3217;
assign w4566 = w3673 & w4565;
assign w4567 = w2936 & w4564;
assign w4568 = w4566 & w4567;
assign w4569 = w4557 & w4568;
assign w4570 = w4538 & w4569;
assign w4571 = w4343 & ~w4570;
assign w4572 = ~w4343 & w4570;
assign w4573 = ~w4571 & ~w4572;
assign w4574 = (w1399 & ~w3658) | (w1399 & w32843) | (~w3658 & w32843);
assign w4575 = (w1327 & ~w2005) | (w1327 & w32844) | (~w2005 & w32844);
assign w4576 = (w668 & ~w1913) | (w668 & w32845) | (~w1913 & w32845);
assign w4577 = w3723 & ~w3725;
assign w4578 = ~w3726 & ~w4577;
assign w4579 = ~w4575 & ~w4576;
assign w4580 = ~w4574 & w4579;
assign w4581 = (w4580 & w4578) | (w4580 & w32846) | (w4578 & w32846);
assign w4582 = w4573 & ~w4581;
assign w4583 = a_20 & ~w4418;
assign w4584 = ~w4419 & ~w4583;
assign w4585 = (~w4581 & w32848) | (~w4581 & w32849) | (w32848 & w32849);
assign w4586 = (w4581 & w32850) | (w4581 & w32851) | (w32850 & w32851);
assign w4587 = ~w4585 & ~w4586;
assign w4588 = (w1327 & ~w1913) | (w1327 & w32852) | (~w1913 & w32852);
assign w4589 = (w1399 & ~w2005) | (w1399 & w32853) | (~w2005 & w32853);
assign w4590 = (w668 & ~w1714) | (w668 & w32780) | (~w1714 & w32780);
assign w4591 = (~w3723 & w32854) | (~w3723 & w32855) | (w32854 & w32855);
assign w4592 = ~w3727 & ~w4591;
assign w4593 = ~w4588 & ~w4589;
assign w4594 = ~w4590 & w4593;
assign w4595 = (w4594 & ~w4592) | (w4594 & w32856) | (~w4592 & w32856);
assign w4596 = w4587 & ~w4595;
assign w4597 = (~w4585 & ~w4587) | (~w4585 & w32857) | (~w4587 & w32857);
assign w4598 = (w4428 & w32858) | (w4428 & w32859) | (w32858 & w32859);
assign w4599 = ~w4432 & ~w4598;
assign w4600 = ~w4597 & w4599;
assign w4601 = w4597 & ~w4599;
assign w4602 = ~w4600 & ~w4601;
assign w4603 = ~w3813 & w3957;
assign w4604 = (w4446 & ~w643) | (w4446 & w32860) | (~w643 & w32860);
assign w4605 = (w4068 & ~w1628) | (w4068 & w32861) | (~w1628 & w32861);
assign w4606 = w4070 & w4224;
assign w4607 = ~w4603 & w32862;
assign w4608 = ~w4606 & w32863;
assign w4609 = (~a_29 & w4606) | (~a_29 & w32864) | (w4606 & w32864);
assign w4610 = ~w4608 & ~w4609;
assign w4611 = w4602 & ~w4610;
assign w4612 = (~w4600 & ~w4602) | (~w4600 & w32865) | (~w4602 & w32865);
assign w4613 = ~w4503 & w4511;
assign w4614 = ~w4512 & ~w4613;
assign w4615 = ~w4612 & w4614;
assign w4616 = w4436 & ~w4438;
assign w4617 = ~w4439 & ~w4616;
assign w4618 = (~w4612 & w32867) | (~w4612 & w32868) | (w32867 & w32868);
assign w4619 = (w4612 & w32869) | (w4612 & w32870) | (w32869 & w32870);
assign w4620 = ~w4618 & ~w4619;
assign w4621 = ~w1397 & w4446;
assign w4622 = ~w1475 & w4068;
assign w4623 = (w3957 & ~w643) | (w3957 & w32871) | (~w643 & w32871);
assign w4624 = ~w4621 & ~w4623;
assign w4625 = ~w4622 & w4624;
assign w4626 = (w4625 & ~w4056) | (w4625 & w32872) | (~w4056 & w32872);
assign w4627 = a_29 & ~w4626;
assign w4628 = (~w4056 & w32873) | (~w4056 & w32874) | (w32873 & w32874);
assign w4629 = ~w4627 & ~w4628;
assign w4630 = w4620 & w4629;
assign w4631 = (~w4618 & ~w4620) | (~w4618 & w32875) | (~w4620 & w32875);
assign w4632 = ~w4445 & ~w4455;
assign w4633 = ~w4456 & ~w4632;
assign w4634 = ~w4631 & w4633;
assign w4635 = w4631 & ~w4633;
assign w4636 = ~w4634 & ~w4635;
assign w4637 = (~w518 & ~w3904) | (~w518 & w32876) | (~w3904 & w32876);
assign w4638 = w1222 & ~w3889;
assign w4639 = ~w3958 & w4638;
assign w4640 = ~w4637 & ~w4639;
assign w4641 = (w4640 & ~w4073) | (w4640 & w32877) | (~w4073 & w32877);
assign w4642 = a_26 & w4641;
assign w4643 = (w4073 & w32878) | (w4073 & w32879) | (w32878 & w32879);
assign w4644 = ~w4642 & ~w4643;
assign w4645 = w4636 & ~w4644;
assign w4646 = (~w4634 & ~w4636) | (~w4634 & w32880) | (~w4636 & w32880);
assign w4647 = ~w4492 & ~w4494;
assign w4648 = ~w4495 & ~w4647;
assign w4649 = w4646 & ~w4648;
assign w4650 = ~w4646 & w4648;
assign w4651 = w4612 & ~w4614;
assign w4652 = ~w4615 & ~w4651;
assign w4653 = ~w1475 & w4446;
assign w4654 = (w3957 & ~w1628) | (w3957 & w32881) | (~w1628 & w32881);
assign w4655 = (w4068 & ~w643) | (w4068 & w32882) | (~w643 & w32882);
assign w4656 = ~w4654 & ~w4655;
assign w4657 = ~w4653 & w4656;
assign w4658 = (w4657 & ~w4041) | (w4657 & w32883) | (~w4041 & w32883);
assign w4659 = a_29 & w4658;
assign w4660 = (w4041 & w32884) | (w4041 & w32885) | (w32884 & w32885);
assign w4661 = ~w4659 & ~w4660;
assign w4662 = w4652 & ~w4661;
assign w4663 = ~w4652 & w4661;
assign w4664 = ~w4662 & ~w4663;
assign w4665 = (w4638 & ~w1308) | (w4638 & w32886) | (~w1308 & w32886);
assign w4666 = ~w1222 & w1225;
assign w4667 = (w4666 & ~w3904) | (w4666 & w32887) | (~w3904 & w32887);
assign w4668 = ~w518 & ~w1397;
assign w4669 = ~w4665 & ~w4668;
assign w4670 = ~w4667 & w4669;
assign w4671 = (w4670 & ~w3964) | (w4670 & w32888) | (~w3964 & w32888);
assign w4672 = ~a_26 & w4671;
assign w4673 = (w3964 & w32889) | (w3964 & w32890) | (w32889 & w32890);
assign w4674 = ~w4672 & ~w4673;
assign w4675 = w4664 & w4674;
assign w4676 = (~w4662 & ~w4664) | (~w4662 & w32891) | (~w4664 & w32891);
assign w4677 = (w4638 & ~w3904) | (w4638 & w32892) | (~w3904 & w32892);
assign w4678 = (~w518 & ~w1308) | (~w518 & w32893) | (~w1308 & w32893);
assign w4679 = ~w3958 & w4666;
assign w4680 = ~w4678 & ~w4679;
assign w4681 = ~w4677 & w4680;
assign w4682 = (w4681 & ~w3943) | (w4681 & w32894) | (~w3943 & w32894);
assign w4683 = a_26 & ~w4682;
assign w4684 = (~w3943 & w32895) | (~w3943 & w32896) | (w32895 & w32896);
assign w4685 = ~w4683 & ~w4684;
assign w4686 = ~w4676 & w4685;
assign w4687 = ~w4620 & ~w4629;
assign w4688 = ~w4630 & ~w4687;
assign w4689 = w4676 & ~w4685;
assign w4690 = ~w4686 & ~w4689;
assign w4691 = w4688 & w4690;
assign w4692 = (~w4686 & ~w4690) | (~w4686 & w32897) | (~w4690 & w32897);
assign w4693 = ~w4636 & w4644;
assign w4694 = ~w4645 & ~w4693;
assign w4695 = ~w4692 & w4694;
assign w4696 = w4692 & ~w4694;
assign w4697 = ~w4695 & ~w4696;
assign w4698 = ~w4587 & w4595;
assign w4699 = ~w4596 & ~w4698;
assign w4700 = (w4446 & ~w1628) | (w4446 & w32898) | (~w1628 & w32898);
assign w4701 = (w3957 & ~w1807) | (w3957 & w32899) | (~w1807 & w32899);
assign w4702 = ~w3813 & w4068;
assign w4703 = ~w4700 & ~w4701;
assign w4704 = ~w4702 & w4703;
assign w4705 = (w4704 & ~w4244) | (w4704 & w32900) | (~w4244 & w32900);
assign w4706 = a_29 & ~w4705;
assign w4707 = (~w4244 & w32901) | (~w4244 & w32902) | (w32901 & w32902);
assign w4708 = ~w4706 & ~w4707;
assign w4709 = w4699 & w4708;
assign w4710 = ~w74 & ~w134;
assign w4711 = ~w645 & w2684;
assign w4712 = ~w212 & ~w476;
assign w4713 = ~w475 & ~w698;
assign w4714 = ~w81 & ~w395;
assign w4715 = w650 & w742;
assign w4716 = w866 & w1770;
assign w4717 = w3063 & w4710;
assign w4718 = w4712 & w4713;
assign w4719 = w4714 & w4718;
assign w4720 = w4716 & w4717;
assign w4721 = w4344 & w4715;
assign w4722 = w4711 & w4721;
assign w4723 = w4719 & w4720;
assign w4724 = w1724 & w4723;
assign w4725 = w2996 & w4722;
assign w4726 = w4724 & w4725;
assign w4727 = w1354 & w2753;
assign w4728 = w4726 & w4727;
assign w4729 = w616 & w4728;
assign w4730 = ~w249 & w1758;
assign w4731 = ~w39 & ~w164;
assign w4732 = ~w136 & ~w291;
assign w4733 = ~w220 & ~w996;
assign w4734 = w587 & w4733;
assign w4735 = ~w714 & w2008;
assign w4736 = w4311 & w4735;
assign w4737 = ~w68 & ~w81;
assign w4738 = ~w163 & ~w1051;
assign w4739 = w4737 & w4738;
assign w4740 = w2102 & w2970;
assign w4741 = w4739 & w4740;
assign w4742 = ~w144 & w1423;
assign w4743 = w1861 & w2153;
assign w4744 = w2501 & w3516;
assign w4745 = w4732 & w4744;
assign w4746 = w4742 & w4743;
assign w4747 = w91 & w621;
assign w4748 = w4734 & w4747;
assign w4749 = w4745 & w4746;
assign w4750 = w3121 & w4736;
assign w4751 = w4741 & w4750;
assign w4752 = w4748 & w4749;
assign w4753 = w4751 & w4752;
assign w4754 = ~w130 & ~w180;
assign w4755 = ~w446 & ~w538;
assign w4756 = ~w649 & w4755;
assign w4757 = w17 & ~w544;
assign w4758 = w405 & w672;
assign w4759 = w853 & w952;
assign w4760 = w2183 & w2307;
assign w4761 = w3502 & w4731;
assign w4762 = w4754 & w4761;
assign w4763 = w4759 & w4760;
assign w4764 = w4757 & w4758;
assign w4765 = w1642 & w4730;
assign w4766 = w4756 & w4765;
assign w4767 = w4763 & w4764;
assign w4768 = w566 & w4762;
assign w4769 = w4767 & w4768;
assign w4770 = w4766 & w4769;
assign w4771 = w4753 & w4770;
assign w4772 = w3795 & w4771;
assign w4773 = ~w4729 & ~w4772;
assign w4774 = w4729 & w4772;
assign w4775 = ~w4773 & ~w4774;
assign w4776 = ~a_17 & w4775;
assign w4777 = (~w4773 & ~w4775) | (~w4773 & w32903) | (~w4775 & w32903);
assign w4778 = w4343 & ~w4777;
assign w4779 = ~w4343 & w4777;
assign w4780 = ~w4778 & ~w4779;
assign w4781 = (w1327 & ~w3658) | (w1327 & w32904) | (~w3658 & w32904);
assign w4782 = (w1399 & ~w3712) | (w1399 & w32905) | (~w3712 & w32905);
assign w4783 = (w668 & ~w2005) | (w668 & w32906) | (~w2005 & w32906);
assign w4784 = w2006 & w3659;
assign w4785 = ~w3660 & ~w4784;
assign w4786 = ~w2238 & ~w3718;
assign w4787 = w3625 & w32907;
assign w4788 = (~w3559 & w32909) | (~w3559 & w32910) | (w32909 & w32910);
assign w4789 = (~w3720 & ~w4788) | (~w3720 & w32911) | (~w4788 & w32911);
assign w4790 = w4785 & ~w4789;
assign w4791 = (~w4788 & w32912) | (~w4788 & w32913) | (w32912 & w32913);
assign w4792 = (w1478 & w4790) | (w1478 & w32914) | (w4790 & w32914);
assign w4793 = ~w4782 & ~w4783;
assign w4794 = ~w4781 & w4793;
assign w4795 = (w4780 & w4792) | (w4780 & w32915) | (w4792 & w32915);
assign w4796 = (~w4792 & w32916) | (~w4792 & w32917) | (w32916 & w32917);
assign w4797 = (w4578 & w32918) | (w4578 & w32919) | (w32918 & w32919);
assign w4798 = ~w4582 & ~w4797;
assign w4799 = ~w4796 & w4798;
assign w4800 = w4796 & ~w4798;
assign w4801 = ~w4799 & ~w4800;
assign w4802 = a_17 & ~w4775;
assign w4803 = ~w4776 & ~w4802;
assign w4804 = (w668 & ~w3658) | (w668 & w32920) | (~w3658 & w32920);
assign w4805 = (w1327 & ~w3712) | (w1327 & w32921) | (~w3712 & w32921);
assign w4806 = (w1399 & ~w2235) | (w1399 & w32922) | (~w2235 & w32922);
assign w4807 = ~w3715 & ~w3720;
assign w4808 = (w3559 & w32925) | (w3559 & w32926) | (w32925 & w32926);
assign w4809 = (~w3559 & w32927) | (~w3559 & w32928) | (w32927 & w32928);
assign w4810 = ~w4808 & ~w4809;
assign w4811 = ~w4805 & ~w4806;
assign w4812 = ~w4804 & w4811;
assign w4813 = (w4812 & ~w4810) | (w4812 & w32929) | (~w4810 & w32929);
assign w4814 = w4803 & ~w4813;
assign w4815 = ~w65 & ~w834;
assign w4816 = ~w249 & ~w404;
assign w4817 = ~w653 & w2681;
assign w4818 = ~w245 & ~w256;
assign w4819 = ~w62 & ~w86;
assign w4820 = ~w170 & ~w206;
assign w4821 = ~w341 & ~w4001;
assign w4822 = w4820 & w4821;
assign w4823 = w840 & w4819;
assign w4824 = w877 & w1102;
assign w4825 = w3347 & w4818;
assign w4826 = w4824 & w4825;
assign w4827 = w4822 & w4823;
assign w4828 = w4817 & w4827;
assign w4829 = w3158 & w4826;
assign w4830 = w4828 & w4829;
assign w4831 = ~w319 & ~w907;
assign w4832 = w1041 & w4831;
assign w4833 = w1969 & w2329;
assign w4834 = w2782 & w2925;
assign w4835 = w4815 & w4816;
assign w4836 = w4834 & w4835;
assign w4837 = w4832 & w4833;
assign w4838 = w906 & w4837;
assign w4839 = w1867 & w4836;
assign w4840 = w2844 & w4839;
assign w4841 = w2453 & w4838;
assign w4842 = w4840 & w4841;
assign w4843 = w204 & w4830;
assign w4844 = w4842 & w4843;
assign w4845 = w772 & w4844;
assign w4846 = w4729 & ~w4845;
assign w4847 = ~w288 & ~w357;
assign w4848 = ~w992 & w4847;
assign w4849 = ~w130 & ~w368;
assign w4850 = ~w62 & ~w476;
assign w4851 = w351 & ~w895;
assign w4852 = ~w112 & ~w719;
assign w4853 = ~w593 & ~w647;
assign w4854 = w1124 & w4853;
assign w4855 = w2379 & w2786;
assign w4856 = w4852 & w4855;
assign w4857 = w727 & w4854;
assign w4858 = w1318 & w2217;
assign w4859 = w4851 & w4858;
assign w4860 = w4856 & w4857;
assign w4861 = w2396 & w3766;
assign w4862 = w4860 & w4861;
assign w4863 = w4859 & w4862;
assign w4864 = ~w473 & w1736;
assign w4865 = ~w67 & ~w447;
assign w4866 = w17 & w4865;
assign w4867 = w564 & w4866;
assign w4868 = w4864 & w4867;
assign w4869 = w624 & w840;
assign w4870 = w1199 & w1413;
assign w4871 = w2569 & w4732;
assign w4872 = w4849 & w4850;
assign w4873 = w4871 & w4872;
assign w4874 = w4869 & w4870;
assign w4875 = w2887 & w4848;
assign w4876 = w4874 & w4875;
assign w4877 = w4310 & w4873;
assign w4878 = w4876 & w4877;
assign w4879 = w4868 & w4878;
assign w4880 = w417 & w4879;
assign w4881 = w4863 & w4880;
assign w4882 = w235 & w4881;
assign w4883 = ~w418 & ~w540;
assign w4884 = ~w585 & ~w2331;
assign w4885 = ~w67 & ~w395;
assign w4886 = ~w420 & w4885;
assign w4887 = w950 & w1868;
assign w4888 = w1919 & w2036;
assign w4889 = w2846 & w4883;
assign w4890 = w4884 & w4889;
assign w4891 = w4887 & w4888;
assign w4892 = w1991 & w4886;
assign w4893 = w4891 & w4892;
assign w4894 = w2884 & w4890;
assign w4895 = w4542 & w4894;
assign w4896 = w4893 & w4895;
assign w4897 = ~w423 & ~w1040;
assign w4898 = ~w191 & w1974;
assign w4899 = w4897 & w4898;
assign w4900 = w3332 & w4899;
assign w4901 = w449 & w3567;
assign w4902 = ~w389 & w4731;
assign w4903 = ~w157 & ~w451;
assign w4904 = w1098 & w4903;
assign w4905 = w2549 & w2990;
assign w4906 = w3124 & w3677;
assign w4907 = w4754 & w4906;
assign w4908 = w4904 & w4905;
assign w4909 = w4902 & w4908;
assign w4910 = w4907 & w4909;
assign w4911 = ~w18 & ~w170;
assign w4912 = ~w113 & ~w1192;
assign w4913 = ~w342 & ~w544;
assign w4914 = ~w149 & w735;
assign w4915 = w947 & w3576;
assign w4916 = w3583 & w4911;
assign w4917 = w4912 & w4913;
assign w4918 = w4916 & w4917;
assign w4919 = w4914 & w4915;
assign w4920 = w4817 & w4919;
assign w4921 = w4918 & w4920;
assign w4922 = w1503 & w4921;
assign w4923 = w4910 & w4922;
assign w4924 = ~w590 & ~w671;
assign w4925 = ~w115 & ~w197;
assign w4926 = ~w732 & w4925;
assign w4927 = ~w65 & ~w260;
assign w4928 = ~w356 & w4927;
assign w4929 = w3663 & w4924;
assign w4930 = w4928 & w4929;
assign w4931 = w2018 & w2849;
assign w4932 = w4926 & w4931;
assign w4933 = w4930 & w4932;
assign w4934 = ~w362 & ~w538;
assign w4935 = w810 & w1374;
assign w4936 = w1614 & w3155;
assign w4937 = w4934 & w4936;
assign w4938 = w629 & w4935;
assign w4939 = w2162 & w4256;
assign w4940 = w4901 & w4939;
assign w4941 = w4937 & w4938;
assign w4942 = w4940 & w4941;
assign w4943 = w4900 & w4942;
assign w4944 = w4933 & w4943;
assign w4945 = w4896 & w4944;
assign w4946 = w4923 & w4945;
assign w4947 = ~w4882 & ~w4946;
assign w4948 = w4882 & w4946;
assign w4949 = ~w4947 & ~w4948;
assign w4950 = ~a_14 & w4949;
assign w4951 = (~w4947 & ~w4949) | (~w4947 & w32930) | (~w4949 & w32930);
assign w4952 = w4845 & ~w4951;
assign w4953 = ~w4845 & w4951;
assign w4954 = ~w4952 & ~w4953;
assign w4955 = w1399 & ~w2075;
assign w4956 = (w668 & ~w2235) | (w668 & w32931) | (~w2235 & w32931);
assign w4957 = w1327 & ~w2148;
assign w4958 = (w3625 & w3559) | (w3625 & w32932) | (w3559 & w32932);
assign w4959 = ~w2237 & ~w3619;
assign w4960 = (w4959 & w4958) | (w4959 & w32933) | (w4958 & w32933);
assign w4961 = ~w4958 & w32934;
assign w4962 = ~w4960 & ~w4961;
assign w4963 = ~w4956 & ~w4957;
assign w4964 = ~w4955 & w4963;
assign w4965 = (w4964 & ~w4962) | (w4964 & w32935) | (~w4962 & w32935);
assign w4966 = w4954 & ~w4965;
assign w4967 = ~w4729 & w4845;
assign w4968 = ~w4846 & ~w4967;
assign w4969 = (~w4965 & w32937) | (~w4965 & w32938) | (w32937 & w32938);
assign w4970 = (w4965 & w32939) | (w4965 & w32940) | (w32939 & w32940);
assign w4971 = (~w4810 & w32941) | (~w4810 & w32942) | (w32941 & w32942);
assign w4972 = ~w4814 & ~w4971;
assign w4973 = ~w4970 & w4972;
assign w4974 = ~w4814 & ~w4973;
assign w4975 = ~w4792 & w32943;
assign w4976 = ~w4795 & ~w4975;
assign w4977 = ~w4974 & w4976;
assign w4978 = w4974 & ~w4976;
assign w4979 = ~w4977 & ~w4978;
assign w4980 = (w3957 & ~w1913) | (w3957 & w32944) | (~w1913 & w32944);
assign w4981 = (w4446 & ~w1807) | (w4446 & w32945) | (~w1807 & w32945);
assign w4982 = (w4068 & ~w1714) | (w4068 & w32861) | (~w1714 & w32861);
assign w4983 = ~w4980 & ~w4981;
assign w4984 = ~w4982 & w4983;
assign w4985 = (w4984 & w4428) | (w4984 & w32946) | (w4428 & w32946);
assign w4986 = a_29 & ~w4985;
assign w4987 = (w4428 & w32947) | (w4428 & w32948) | (w32947 & w32948);
assign w4988 = ~w4986 & ~w4987;
assign w4989 = w4979 & w4988;
assign w4990 = (~w4977 & ~w4979) | (~w4977 & w32949) | (~w4979 & w32949);
assign w4991 = w4801 & ~w4990;
assign w4992 = (~w4799 & w4990) | (~w4799 & w32950) | (w4990 & w32950);
assign w4993 = ~w4699 & ~w4708;
assign w4994 = ~w4709 & ~w4993;
assign w4995 = ~w4992 & w4994;
assign w4996 = (~w4709 & w4992) | (~w4709 & w32951) | (w4992 & w32951);
assign w4997 = ~w4602 & w4610;
assign w4998 = ~w4611 & ~w4997;
assign w4999 = ~w4996 & w4998;
assign w5000 = w4996 & ~w4998;
assign w5001 = ~w4999 & ~w5000;
assign w5002 = (w4666 & ~w1308) | (w4666 & w32952) | (~w1308 & w32952);
assign w5003 = ~w1397 & w4638;
assign w5004 = ~w518 & ~w1475;
assign w5005 = ~w5002 & ~w5003;
assign w5006 = ~w5004 & w5005;
assign w5007 = (w5006 & ~w3834) | (w5006 & w32953) | (~w3834 & w32953);
assign w5008 = a_26 & ~w5007;
assign w5009 = (~w3834 & w32954) | (~w3834 & w32955) | (w32954 & w32955);
assign w5010 = ~w5008 & ~w5009;
assign w5011 = w5001 & w5010;
assign w5012 = (~w4999 & ~w5001) | (~w4999 & w32956) | (~w5001 & w32956);
assign w5013 = a_22 & ~a_23;
assign w5014 = ~a_22 & a_23;
assign w5015 = ~w5013 & ~w5014;
assign w5016 = w508 & ~w5015;
assign w5017 = w504 & ~w5015;
assign w5018 = (~w3828 & w32959) | (~w3828 & w32960) | (w32959 & w32960);
assign w5019 = ~w5018 & w32961;
assign w5020 = (a_23 & w5018) | (a_23 & w32962) | (w5018 & w32962);
assign w5021 = ~w5019 & ~w5020;
assign w5022 = ~w5012 & ~w5021;
assign w5023 = ~w4664 & ~w4674;
assign w5024 = ~w4675 & ~w5023;
assign w5025 = w5012 & w5021;
assign w5026 = ~w5022 & ~w5025;
assign w5027 = w5024 & w5026;
assign w5028 = (~w5022 & ~w5026) | (~w5022 & w32963) | (~w5026 & w32963);
assign w5029 = ~w4688 & ~w4690;
assign w5030 = ~w4691 & ~w5029;
assign w5031 = ~w5028 & w5030;
assign w5032 = w5028 & ~w5030;
assign w5033 = ~w5031 & ~w5032;
assign w5034 = w4992 & ~w4994;
assign w5035 = ~w4995 & ~w5034;
assign w5036 = ~w1397 & w4666;
assign w5037 = ~w1475 & w4638;
assign w5038 = (~w518 & ~w643) | (~w518 & w32964) | (~w643 & w32964);
assign w5039 = ~w5036 & ~w5038;
assign w5040 = ~w5037 & w5039;
assign w5041 = (w5040 & ~w4056) | (w5040 & w32965) | (~w4056 & w32965);
assign w5042 = a_26 & ~w5041;
assign w5043 = (~w4056 & w32966) | (~w4056 & w32967) | (w32966 & w32967);
assign w5044 = ~w5042 & ~w5043;
assign w5045 = w5035 & w5044;
assign w5046 = ~w4801 & w4990;
assign w5047 = ~w4991 & ~w5046;
assign w5048 = ~w3813 & w4446;
assign w5049 = (w3957 & ~w1714) | (w3957 & w32881) | (~w1714 & w32881);
assign w5050 = (w4068 & ~w1807) | (w4068 & w32968) | (~w1807 & w32968);
assign w5051 = w4070 & w4508;
assign w5052 = ~w5048 & w32969;
assign w5053 = (a_29 & w5051) | (a_29 & w32970) | (w5051 & w32970);
assign w5054 = ~w5051 & w32971;
assign w5055 = ~w5053 & ~w5054;
assign w5056 = w5047 & w5055;
assign w5057 = ~w5047 & ~w5055;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = ~w1475 & w4666;
assign w5060 = (w4638 & ~w643) | (w4638 & w32972) | (~w643 & w32972);
assign w5061 = (~w518 & ~w1628) | (~w518 & w32973) | (~w1628 & w32973);
assign w5062 = ~w5060 & ~w5061;
assign w5063 = ~w5059 & w5062;
assign w5064 = (w5063 & ~w4041) | (w5063 & w32974) | (~w4041 & w32974);
assign w5065 = a_26 & ~w5064;
assign w5066 = (~w4041 & w32975) | (~w4041 & w32976) | (w32975 & w32976);
assign w5067 = ~w5065 & ~w5066;
assign w5068 = w5058 & w5067;
assign w5069 = (~w5056 & ~w5058) | (~w5056 & w32977) | (~w5058 & w32977);
assign w5070 = ~w5035 & ~w5044;
assign w5071 = ~w5045 & ~w5070;
assign w5072 = ~w5069 & w5071;
assign w5073 = ~w5045 & ~w5072;
assign w5074 = ~w5001 & ~w5010;
assign w5075 = ~w5011 & ~w5074;
assign w5076 = ~w5073 & w5075;
assign w5077 = w5073 & ~w5075;
assign w5078 = ~w5076 & ~w5077;
assign w5079 = (w5016 & ~w3904) | (w5016 & w32978) | (~w3904 & w32978);
assign w5080 = ~w504 & w507;
assign w5081 = ~w3958 & w5080;
assign w5082 = ~w5079 & ~w5081;
assign w5083 = (w5082 & ~w4073) | (w5082 & w32979) | (~w4073 & w32979);
assign w5084 = a_23 & w5083;
assign w5085 = (w4073 & w32980) | (w4073 & w32981) | (w32980 & w32981);
assign w5086 = ~w5084 & ~w5085;
assign w5087 = w5078 & ~w5086;
assign w5088 = (~w5076 & ~w5078) | (~w5076 & w32982) | (~w5078 & w32982);
assign w5089 = ~w5024 & ~w5026;
assign w5090 = ~w5027 & ~w5089;
assign w5091 = ~w5088 & w5090;
assign w5092 = w5033 & w5091;
assign w5093 = ~w4979 & ~w4988;
assign w5094 = ~w4989 & ~w5093;
assign w5095 = (w4965 & w32983) | (w4965 & w32984) | (w32983 & w32984);
assign w5096 = ~w4969 & ~w5095;
assign w5097 = (w668 & ~w3712) | (w668 & w32985) | (~w3712 & w32985);
assign w5098 = w1399 & ~w2148;
assign w5099 = (w1327 & ~w2235) | (w1327 & w32986) | (~w2235 & w32986);
assign w5100 = ~w3714 & ~w3718;
assign w5101 = (w3559 & w32987) | (w3559 & w32988) | (w32987 & w32988);
assign w5102 = (~w3559 & w32989) | (~w3559 & w32990) | (w32989 & w32990);
assign w5103 = ~w5101 & ~w5102;
assign w5104 = w1478 & w5103;
assign w5105 = ~w5098 & w32991;
assign w5106 = ~w5104 & w5105;
assign w5107 = w5096 & ~w5106;
assign w5108 = ~w5096 & w5106;
assign w5109 = ~w5107 & ~w5108;
assign w5110 = (w3957 & ~w3658) | (w3957 & w32992) | (~w3658 & w32992);
assign w5111 = (w4068 & ~w2005) | (w4068 & w32993) | (~w2005 & w32993);
assign w5112 = (w4446 & ~w1913) | (w4446 & w32994) | (~w1913 & w32994);
assign w5113 = ~w5111 & ~w5112;
assign w5114 = ~w5110 & w5113;
assign w5115 = (w5114 & w4578) | (w5114 & w32995) | (w4578 & w32995);
assign w5116 = a_29 & ~w5115;
assign w5117 = (w4578 & w32996) | (w4578 & w32997) | (w32996 & w32997);
assign w5118 = ~w5116 & ~w5117;
assign w5119 = w5109 & w5118;
assign w5120 = (~w5107 & ~w5109) | (~w5107 & w32998) | (~w5109 & w32998);
assign w5121 = w4970 & ~w4972;
assign w5122 = ~w4973 & ~w5121;
assign w5123 = w5120 & ~w5122;
assign w5124 = ~w5120 & w5122;
assign w5125 = ~w5123 & ~w5124;
assign w5126 = (w4068 & ~w1913) | (w4068 & w32999) | (~w1913 & w32999);
assign w5127 = (w3957 & ~w2005) | (w3957 & w33000) | (~w2005 & w33000);
assign w5128 = (w4446 & ~w1714) | (w4446 & w32898) | (~w1714 & w32898);
assign w5129 = ~w5126 & ~w5127;
assign w5130 = ~w5128 & w5129;
assign w5131 = (w5130 & ~w4592) | (w5130 & w33001) | (~w4592 & w33001);
assign w5132 = a_29 & ~w5131;
assign w5133 = (~w4592 & w33002) | (~w4592 & w33003) | (w33002 & w33003);
assign w5134 = ~w5132 & ~w5133;
assign w5135 = w5125 & ~w5134;
assign w5136 = (~w5123 & ~w5125) | (~w5123 & w33004) | (~w5125 & w33004);
assign w5137 = ~w5094 & ~w5136;
assign w5138 = w5094 & w5136;
assign w5139 = ~w5137 & ~w5138;
assign w5140 = ~w518 & ~w3813;
assign w5141 = (w4666 & ~w643) | (w4666 & w33005) | (~w643 & w33005);
assign w5142 = (w4638 & ~w1628) | (w4638 & w33006) | (~w1628 & w33006);
assign w5143 = w1226 & w4224;
assign w5144 = ~w5140 & w33007;
assign w5145 = (a_26 & w5143) | (a_26 & w33008) | (w5143 & w33008);
assign w5146 = ~w5143 & w33009;
assign w5147 = ~w5145 & ~w5146;
assign w5148 = w5139 & ~w5147;
assign w5149 = ~w5139 & w5147;
assign w5150 = ~w5148 & ~w5149;
assign w5151 = ~w5125 & w5134;
assign w5152 = ~w5135 & ~w5151;
assign w5153 = (~w518 & ~w1807) | (~w518 & w33010) | (~w1807 & w33010);
assign w5154 = (w4666 & ~w1628) | (w4666 & w33011) | (~w1628 & w33011);
assign w5155 = ~w3813 & w4638;
assign w5156 = ~w5153 & ~w5154;
assign w5157 = ~w5155 & w5156;
assign w5158 = (w5157 & ~w4244) | (w5157 & w33012) | (~w4244 & w33012);
assign w5159 = a_26 & ~w5158;
assign w5160 = (~w4244 & w33013) | (~w4244 & w33014) | (w33013 & w33014);
assign w5161 = ~w5159 & ~w5160;
assign w5162 = ~w5152 & w5161;
assign w5163 = ~w16 & ~w118;
assign w5164 = ~w180 & ~w1077;
assign w5165 = w5163 & w5164;
assign w5166 = w4254 & w5165;
assign w5167 = w1928 & w5166;
assign w5168 = ~w134 & ~w451;
assign w5169 = ~w365 & ~w737;
assign w5170 = w1266 & w2454;
assign w5171 = ~w188 & w1693;
assign w5172 = ~w249 & ~w530;
assign w5173 = w3770 & w5172;
assign w5174 = w587 & w792;
assign w5175 = w1054 & w3212;
assign w5176 = w4714 & w5168;
assign w5177 = w5169 & w5176;
assign w5178 = w5174 & w5175;
assign w5179 = w3433 & w5170;
assign w5180 = w5171 & w5173;
assign w5181 = w5179 & w5180;
assign w5182 = w5177 & w5178;
assign w5183 = w1637 & w5182;
assign w5184 = w5181 & w5183;
assign w5185 = ~w60 & ~w653;
assign w5186 = ~w356 & ~w547;
assign w5187 = ~w163 & ~w290;
assign w5188 = ~w237 & ~w996;
assign w5189 = ~w671 & ~w896;
assign w5190 = w744 & w5189;
assign w5191 = w757 & w959;
assign w5192 = w5187 & w5188;
assign w5193 = w5191 & w5192;
assign w5194 = w991 & w5190;
assign w5195 = w1159 & w1465;
assign w5196 = w1740 & w4329;
assign w5197 = w5195 & w5196;
assign w5198 = w5193 & w5194;
assign w5199 = w5197 & w5198;
assign w5200 = w4007 & w5199;
assign w5201 = ~w18 & ~w39;
assign w5202 = ~w53 & w5201;
assign w5203 = w430 & w594;
assign w5204 = w2689 & w3013;
assign w5205 = w3169 & w5185;
assign w5206 = w5186 & w5205;
assign w5207 = w5203 & w5204;
assign w5208 = w1601 & w5202;
assign w5209 = w5207 & w5208;
assign w5210 = w3235 & w5206;
assign w5211 = w5209 & w5210;
assign w5212 = w5167 & w5211;
assign w5213 = w336 & w5212;
assign w5214 = w5184 & w5200;
assign w5215 = w5213 & w5214;
assign w5216 = w4882 & ~w5215;
assign w5217 = ~w4882 & w5215;
assign w5218 = ~w5216 & ~w5217;
assign w5219 = w668 & ~w2075;
assign w5220 = w1327 & ~w3615;
assign w5221 = w1399 & ~w2393;
assign w5222 = ~w3617 & ~w3623;
assign w5223 = ~w3616 & ~w3620;
assign w5224 = (w5223 & w3559) | (w5223 & w33015) | (w3559 & w33015);
assign w5225 = (w3559 & w33018) | (w3559 & w33019) | (w33018 & w33019);
assign w5226 = (~w3559 & w33020) | (~w3559 & w33021) | (w33020 & w33021);
assign w5227 = ~w5225 & ~w5226;
assign w5228 = ~w5220 & ~w5221;
assign w5229 = ~w5219 & w5228;
assign w5230 = (w5229 & ~w5227) | (w5229 & w33022) | (~w5227 & w33022);
assign w5231 = w5218 & ~w5230;
assign w5232 = a_14 & ~w4949;
assign w5233 = ~w4950 & ~w5232;
assign w5234 = (~w5230 & w33024) | (~w5230 & w33025) | (w33024 & w33025);
assign w5235 = (w5230 & w33026) | (w5230 & w33027) | (w33026 & w33027);
assign w5236 = ~w5234 & ~w5235;
assign w5237 = w1327 & ~w2075;
assign w5238 = w1399 & ~w3615;
assign w5239 = w668 & ~w2148;
assign w5240 = ~w3617 & ~w3622;
assign w5241 = (~w3559 & w33028) | (~w3559 & w33029) | (w33028 & w33029);
assign w5242 = ~w4958 & ~w5241;
assign w5243 = ~w5238 & ~w5239;
assign w5244 = ~w5237 & w5243;
assign w5245 = (w5244 & ~w5242) | (w5244 & w33030) | (~w5242 & w33030);
assign w5246 = w5236 & ~w5245;
assign w5247 = (~w5234 & ~w5236) | (~w5234 & w33031) | (~w5236 & w33031);
assign w5248 = (~w4962 & w33032) | (~w4962 & w33033) | (w33032 & w33033);
assign w5249 = ~w4966 & ~w5248;
assign w5250 = ~w5247 & w5249;
assign w5251 = w5247 & ~w5249;
assign w5252 = ~w5250 & ~w5251;
assign w5253 = (w4068 & ~w3658) | (w4068 & w33034) | (~w3658 & w33034);
assign w5254 = (w4446 & ~w2005) | (w4446 & w33035) | (~w2005 & w33035);
assign w5255 = (w3957 & ~w3712) | (w3957 & w33036) | (~w3712 & w33036);
assign w5256 = (w4070 & w4790) | (w4070 & w33037) | (w4790 & w33037);
assign w5257 = ~w5254 & ~w5255;
assign w5258 = ~w5253 & w5257;
assign w5259 = (a_29 & w5256) | (a_29 & w33038) | (w5256 & w33038);
assign w5260 = ~w5256 & w33039;
assign w5261 = ~w5259 & ~w5260;
assign w5262 = w5252 & w5261;
assign w5263 = (~w5250 & ~w5252) | (~w5250 & w33040) | (~w5252 & w33040);
assign w5264 = ~w5109 & ~w5118;
assign w5265 = ~w5119 & ~w5264;
assign w5266 = ~w5263 & w5265;
assign w5267 = w5263 & ~w5265;
assign w5268 = ~w5266 & ~w5267;
assign w5269 = ~w3813 & w4666;
assign w5270 = (~w518 & ~w1714) | (~w518 & w32973) | (~w1714 & w32973);
assign w5271 = (w4638 & ~w1807) | (w4638 & w33041) | (~w1807 & w33041);
assign w5272 = w1226 & w4508;
assign w5273 = ~w5269 & w33042;
assign w5274 = (a_26 & w5272) | (a_26 & w33043) | (w5272 & w33043);
assign w5275 = ~w5272 & w33044;
assign w5276 = ~w5274 & ~w5275;
assign w5277 = w5268 & w5276;
assign w5278 = (~w5266 & ~w5268) | (~w5266 & w33045) | (~w5268 & w33045);
assign w5279 = w5152 & ~w5161;
assign w5280 = ~w5162 & ~w5279;
assign w5281 = ~w5278 & w5280;
assign w5282 = (~w5162 & ~w5280) | (~w5162 & w33046) | (~w5280 & w33046);
assign w5283 = w5150 & w5282;
assign w5284 = ~w1397 & w5080;
assign w5285 = ~w1475 & w5016;
assign w5286 = w504 & w5015;
assign w5287 = (w5286 & ~w1308) | (w5286 & w33047) | (~w1308 & w33047);
assign w5288 = ~w5284 & ~w5285;
assign w5289 = ~w5287 & w5288;
assign w5290 = (w5289 & ~w3834) | (w5289 & w33048) | (~w3834 & w33048);
assign w5291 = a_23 & ~w5290;
assign w5292 = (~w3834 & w33049) | (~w3834 & w33050) | (w33049 & w33050);
assign w5293 = ~w5291 & ~w5292;
assign w5294 = ~w5150 & ~w5282;
assign w5295 = ~w5283 & ~w5294;
assign w5296 = ~w5293 & w5295;
assign w5297 = (~w5283 & ~w5295) | (~w5283 & w33051) | (~w5295 & w33051);
assign w5298 = ~a_17 & ~a_18;
assign w5299 = a_17 & a_18;
assign w5300 = ~w5298 & ~w5299;
assign w5301 = ~a_18 & ~a_19;
assign w5302 = a_18 & a_19;
assign w5303 = ~w5301 & ~w5302;
assign w5304 = ~w5300 & ~w5303;
assign w5305 = ~a_19 & a_20;
assign w5306 = a_19 & ~a_20;
assign w5307 = ~w5305 & ~w5306;
assign w5308 = w5304 & ~w5307;
assign w5309 = w5300 & ~w5307;
assign w5310 = (~w3828 & w33054) | (~w3828 & w33055) | (w33054 & w33055);
assign w5311 = ~w5310 & w33056;
assign w5312 = (a_20 & w5310) | (a_20 & w33057) | (w5310 & w33057);
assign w5313 = ~w5311 & ~w5312;
assign w5314 = w5297 & ~w5313;
assign w5315 = ~w5297 & w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = ~w5058 & ~w5067;
assign w5318 = ~w5068 & ~w5317;
assign w5319 = (~w5137 & ~w5139) | (~w5137 & w33058) | (~w5139 & w33058);
assign w5320 = w5318 & w5319;
assign w5321 = ~w5318 & ~w5319;
assign w5322 = ~w5320 & ~w5321;
assign w5323 = ~w1397 & w5016;
assign w5324 = (w5286 & ~w3904) | (w5286 & w33059) | (~w3904 & w33059);
assign w5325 = (w5080 & ~w1308) | (w5080 & w33060) | (~w1308 & w33060);
assign w5326 = ~w5323 & ~w5325;
assign w5327 = ~w5324 & w5326;
assign w5328 = (w5327 & ~w3964) | (w5327 & w33061) | (~w3964 & w33061);
assign w5329 = a_23 & ~w5328;
assign w5330 = (~w3964 & w33062) | (~w3964 & w33063) | (w33062 & w33063);
assign w5331 = ~w5329 & ~w5330;
assign w5332 = w5322 & w5331;
assign w5333 = ~w5322 & ~w5331;
assign w5334 = ~w5332 & ~w5333;
assign w5335 = w5316 & w5334;
assign w5336 = (~w5314 & ~w5316) | (~w5314 & w33064) | (~w5316 & w33064);
assign w5337 = w5069 & ~w5071;
assign w5338 = ~w5072 & ~w5337;
assign w5339 = (~w5320 & ~w5322) | (~w5320 & w33065) | (~w5322 & w33065);
assign w5340 = (w5080 & ~w3904) | (w5080 & w33066) | (~w3904 & w33066);
assign w5341 = ~w3958 & w5286;
assign w5342 = (w5016 & ~w1308) | (w5016 & w33067) | (~w1308 & w33067);
assign w5343 = ~w5341 & ~w5342;
assign w5344 = ~w5340 & w5343;
assign w5345 = (w5344 & ~w3943) | (w5344 & w33068) | (~w3943 & w33068);
assign w5346 = a_23 & ~w5345;
assign w5347 = (~w3943 & w33069) | (~w3943 & w33070) | (w33069 & w33070);
assign w5348 = ~w5346 & ~w5347;
assign w5349 = w5339 & ~w5348;
assign w5350 = ~w5339 & w5348;
assign w5351 = ~w5349 & ~w5350;
assign w5352 = w5338 & w5351;
assign w5353 = ~w5338 & ~w5351;
assign w5354 = ~w5352 & ~w5353;
assign w5355 = ~w5336 & w5354;
assign w5356 = (~w518 & ~w3658) | (~w518 & w33071) | (~w3658 & w33071);
assign w5357 = (w4638 & ~w2005) | (w4638 & w33072) | (~w2005 & w33072);
assign w5358 = (w4666 & ~w1913) | (w4666 & w33073) | (~w1913 & w33073);
assign w5359 = ~w5357 & ~w5358;
assign w5360 = ~w5356 & w5359;
assign w5361 = (w5360 & w4578) | (w5360 & w33074) | (w4578 & w33074);
assign w5362 = a_26 & ~w5361;
assign w5363 = (w4578 & w33075) | (w4578 & w33076) | (w33075 & w33076);
assign w5364 = ~w5362 & ~w5363;
assign w5365 = ~w34 & ~w53;
assign w5366 = ~w349 & w5365;
assign w5367 = ~w559 & ~w741;
assign w5368 = ~w544 & ~w1043;
assign w5369 = ~w65 & ~w572;
assign w5370 = ~w220 & ~w895;
assign w5371 = ~w264 & ~w696;
assign w5372 = ~w166 & w5371;
assign w5373 = ~w337 & ~w431;
assign w5374 = ~w153 & ~w392;
assign w5375 = w2552 & w5374;
assign w5376 = w2807 & w5373;
assign w5377 = w5375 & w5376;
assign w5378 = w605 & w1452;
assign w5379 = w1855 & w2502;
assign w5380 = w4152 & w5370;
assign w5381 = w5379 & w5380;
assign w5382 = w951 & w5378;
assign w5383 = w3418 & w5372;
assign w5384 = w5382 & w5383;
assign w5385 = w5377 & w5381;
assign w5386 = w5384 & w5385;
assign w5387 = ~w159 & ~w170;
assign w5388 = ~w115 & ~w356;
assign w5389 = w132 & w5388;
assign w5390 = ~w71 & ~w180;
assign w5391 = ~w98 & w791;
assign w5392 = w1260 & w1487;
assign w5393 = w3915 & w5387;
assign w5394 = w5390 & w5393;
assign w5395 = w5391 & w5392;
assign w5396 = w2484 & w5389;
assign w5397 = w5395 & w5396;
assign w5398 = w5394 & w5397;
assign w5399 = ~w218 & ~w714;
assign w5400 = w753 & w5399;
assign w5401 = w2501 & w5367;
assign w5402 = w5368 & w5369;
assign w5403 = w5401 & w5402;
assign w5404 = w5366 & w5400;
assign w5405 = w5403 & w5404;
assign w5406 = w259 & w5405;
assign w5407 = w3499 & w4868;
assign w5408 = w5406 & w5407;
assign w5409 = w5386 & w5398;
assign w5410 = w5408 & w5409;
assign w5411 = w1794 & w5410;
assign w5412 = ~w53 & ~w67;
assign w5413 = ~w714 & ~w878;
assign w5414 = w5412 & w5413;
assign w5415 = w2771 & w4088;
assign w5416 = w4852 & w5415;
assign w5417 = w2737 & w5414;
assign w5418 = w5416 & w5417;
assign w5419 = ~w195 & ~w220;
assign w5420 = ~w380 & ~w451;
assign w5421 = w672 & w5420;
assign w5422 = w986 & w1892;
assign w5423 = w2804 & w2871;
assign w5424 = w3119 & w3847;
assign w5425 = w4934 & w5419;
assign w5426 = w5424 & w5425;
assign w5427 = w5422 & w5423;
assign w5428 = w3446 & w5421;
assign w5429 = w5427 & w5428;
assign w5430 = w5426 & w5429;
assign w5431 = w1973 & w5418;
assign w5432 = w5430 & w5431;
assign w5433 = ~w173 & ~w261;
assign w5434 = w165 & w5433;
assign w5435 = w280 & w353;
assign w5436 = w628 & w1152;
assign w5437 = w1423 & w2034;
assign w5438 = w2193 & w2502;
assign w5439 = w3014 & w4710;
assign w5440 = w5438 & w5439;
assign w5441 = w5436 & w5437;
assign w5442 = w5434 & w5435;
assign w5443 = w915 & w5442;
assign w5444 = w5440 & w5441;
assign w5445 = w2124 & w5444;
assign w5446 = w4296 & w5443;
assign w5447 = w5445 & w5446;
assign w5448 = w4103 & w5398;
assign w5449 = w5447 & w5448;
assign w5450 = w5432 & w5449;
assign w5451 = ~w5411 & ~w5450;
assign w5452 = w5411 & w5450;
assign w5453 = ~w5451 & ~w5452;
assign w5454 = ~a_11 & w5453;
assign w5455 = (~w5451 & ~w5453) | (~w5451 & w33077) | (~w5453 & w33077);
assign w5456 = w4882 & ~w5455;
assign w5457 = ~w4882 & w5455;
assign w5458 = ~w5456 & ~w5457;
assign w5459 = w1399 & ~w2306;
assign w5460 = w668 & ~w3615;
assign w5461 = w1327 & ~w2393;
assign w5462 = ~w3559 & w33078;
assign w5463 = ~w5224 & ~w5462;
assign w5464 = ~w5459 & ~w5460;
assign w5465 = ~w5461 & w5464;
assign w5466 = (w5465 & ~w5463) | (w5465 & w33079) | (~w5463 & w33079);
assign w5467 = w5458 & ~w5466;
assign w5468 = (~w5456 & w5466) | (~w5456 & w33080) | (w5466 & w33080);
assign w5469 = (~w5227 & w33081) | (~w5227 & w33082) | (w33081 & w33082);
assign w5470 = ~w5231 & ~w5469;
assign w5471 = ~w5468 & w5470;
assign w5472 = w5468 & ~w5470;
assign w5473 = ~w5471 & ~w5472;
assign w5474 = a_11 & ~w5453;
assign w5475 = ~w5454 & ~w5474;
assign w5476 = w1327 & ~w2306;
assign w5477 = (w1399 & ~w3538) | (w1399 & w33083) | (~w3538 & w33083);
assign w5478 = w668 & ~w2393;
assign w5479 = ~w3554 & ~w3555;
assign w5480 = ~w3547 & w33084;
assign w5481 = ~w3554 & ~w3557;
assign w5482 = (w5481 & w3547) | (w5481 & w33085) | (w3547 & w33085);
assign w5483 = ~w3559 & ~w5482;
assign w5484 = ~w5476 & ~w5477;
assign w5485 = ~w5478 & w5484;
assign w5486 = (w5485 & ~w5483) | (w5485 & w33086) | (~w5483 & w33086);
assign w5487 = w5475 & ~w5486;
assign w5488 = ~w365 & ~w649;
assign w5489 = w950 & w5488;
assign w5490 = ~w88 & ~w216;
assign w5491 = w938 & w5490;
assign w5492 = ~w530 & ~w585;
assign w5493 = ~w206 & ~w282;
assign w5494 = w866 & w5493;
assign w5495 = w5492 & w5494;
assign w5496 = ~w254 & ~w356;
assign w5497 = ~w431 & ~w730;
assign w5498 = w5496 & w5497;
assign w5499 = w517 & w2397;
assign w5500 = w2743 & w2785;
assign w5501 = w5499 & w5500;
assign w5502 = w3662 & w5498;
assign w5503 = w5489 & w5491;
assign w5504 = w5502 & w5503;
assign w5505 = w5495 & w5501;
assign w5506 = w5504 & w5505;
assign w5507 = w4115 & w5506;
assign w5508 = w3166 & w5507;
assign w5509 = w3515 & w5508;
assign w5510 = w3646 & w5509;
assign w5511 = w5411 & ~w5510;
assign w5512 = ~w1104 & w5168;
assign w5513 = ~w74 & ~w313;
assign w5514 = w2715 & w5513;
assign w5515 = w5512 & w5514;
assign w5516 = w648 & w913;
assign w5517 = w1122 & w2093;
assign w5518 = w2620 & w3285;
assign w5519 = w3763 & w5518;
assign w5520 = w5516 & w5517;
assign w5521 = w5519 & w5520;
assign w5522 = ~w178 & ~w339;
assign w5523 = ~w356 & w5522;
assign w5524 = w4816 & w5523;
assign w5525 = w2939 & w5524;
assign w5526 = ~w582 & ~w1123;
assign w5527 = w2405 & w5526;
assign w5528 = w3215 & w3675;
assign w5529 = w5527 & w5528;
assign w5530 = w4162 & w5529;
assign w5531 = ~w10 & ~w83;
assign w5532 = ~w146 & ~w152;
assign w5533 = w5531 & w5532;
assign w5534 = w529 & w758;
assign w5535 = w953 & w2334;
assign w5536 = w3739 & w5535;
assign w5537 = w5533 & w5534;
assign w5538 = w402 & w2011;
assign w5539 = w5537 & w5538;
assign w5540 = w2203 & w5536;
assign w5541 = w5539 & w5540;
assign w5542 = w5525 & w5530;
assign w5543 = w5541 & w5542;
assign w5544 = ~w16 & ~w207;
assign w5545 = w346 & w5544;
assign w5546 = ~w147 & ~w388;
assign w5547 = ~w391 & ~w1192;
assign w5548 = w5546 & w5547;
assign w5549 = w956 & w986;
assign w5550 = w2707 & w3387;
assign w5551 = w4152 & w5550;
assign w5552 = w5548 & w5549;
assign w5553 = w2974 & w4327;
assign w5554 = w5545 & w5553;
assign w5555 = w5551 & w5552;
assign w5556 = w5554 & w5555;
assign w5557 = w4900 & w5556;
assign w5558 = ~w151 & ~w309;
assign w5559 = ~w197 & ~w719;
assign w5560 = w809 & w5559;
assign w5561 = w1265 & w5558;
assign w5562 = w5560 & w5561;
assign w5563 = ~w470 & ~w741;
assign w5564 = ~w337 & ~w544;
assign w5565 = ~w1077 & w5564;
assign w5566 = w464 & w1765;
assign w5567 = w1931 & w2333;
assign w5568 = w3286 & w5419;
assign w5569 = w5563 & w5568;
assign w5570 = w5566 & w5567;
assign w5571 = w5565 & w5570;
assign w5572 = w3425 & w5569;
assign w5573 = w5515 & w5562;
assign w5574 = w5572 & w5573;
assign w5575 = w5521 & w5571;
assign w5576 = w5574 & w5575;
assign w5577 = w5543 & w5576;
assign w5578 = w5557 & w5577;
assign w5579 = w466 & w3495;
assign w5580 = ~w68 & ~w130;
assign w5581 = ~w142 & ~w1965;
assign w5582 = w5580 & w5581;
assign w5583 = w114 & w1079;
assign w5584 = w5582 & w5583;
assign w5585 = w5579 & w5584;
assign w5586 = ~w173 & ~w205;
assign w5587 = w584 & w5586;
assign w5588 = w1157 & w4522;
assign w5589 = w5587 & w5588;
assign w5590 = ~w572 & w1309;
assign w5591 = w129 & ~w152;
assign w5592 = ~w50 & ~w206;
assign w5593 = ~w652 & ~w2716;
assign w5594 = w5592 & w5593;
assign w5595 = w1400 & w3569;
assign w5596 = w4883 & w5595;
assign w5597 = w5591 & w5594;
assign w5598 = w5596 & w5597;
assign w5599 = ~w56 & ~w115;
assign w5600 = ~w135 & w5599;
assign w5601 = w617 & w773;
assign w5602 = w1153 & w1504;
assign w5603 = w3517 & w3739;
assign w5604 = w3916 & w5603;
assign w5605 = w5601 & w5602;
assign w5606 = w4514 & w5600;
assign w5607 = w5590 & w5606;
assign w5608 = w5604 & w5605;
assign w5609 = w1408 & w5589;
assign w5610 = w5608 & w5609;
assign w5611 = w5598 & w5607;
assign w5612 = w5610 & w5611;
assign w5613 = ~w74 & ~w322;
assign w5614 = ~w118 & ~w530;
assign w5615 = w244 & w5614;
assign w5616 = w1273 & w4255;
assign w5617 = w4731 & w5616;
assign w5618 = w5615 & w5617;
assign w5619 = ~w86 & ~w290;
assign w5620 = ~w292 & ~w388;
assign w5621 = ~w585 & ~w776;
assign w5622 = ~w992 & w5621;
assign w5623 = w5619 & w5620;
assign w5624 = w715 & w1028;
assign w5625 = w1639 & w2571;
assign w5626 = w3630 & w4934;
assign w5627 = w5613 & w5626;
assign w5628 = w5624 & w5625;
assign w5629 = w5622 & w5623;
assign w5630 = w5628 & w5629;
assign w5631 = w4526 & w5627;
assign w5632 = w5630 & w5631;
assign w5633 = w5585 & w5618;
assign w5634 = w5632 & w5633;
assign w5635 = w4557 & w5634;
assign w5636 = w5612 & w5635;
assign w5637 = ~w5578 & ~w5636;
assign w5638 = w5578 & w5636;
assign w5639 = ~w5637 & ~w5638;
assign w5640 = ~a_8 & w5639;
assign w5641 = (~w5637 & ~w5639) | (~w5637 & w33087) | (~w5639 & w33087);
assign w5642 = w5411 & ~w5641;
assign w5643 = ~w5411 & w5641;
assign w5644 = ~w5642 & ~w5643;
assign w5645 = w1327 & ~w3403;
assign w5646 = (w668 & ~w3538) | (w668 & w33088) | (~w3538 & w33088);
assign w5647 = w1399 & ~w3475;
assign w5648 = ~w3540 & ~w3548;
assign w5649 = (w3552 & w3328) | (w3552 & w33089) | (w3328 & w33089);
assign w5650 = (w5648 & w5649) | (w5648 & w33090) | (w5649 & w33090);
assign w5651 = ~w5649 & w33091;
assign w5652 = ~w5650 & ~w5651;
assign w5653 = ~w5645 & ~w5646;
assign w5654 = ~w5647 & w5653;
assign w5655 = (w5654 & ~w5652) | (w5654 & w33092) | (~w5652 & w33092);
assign w5656 = w5644 & ~w5655;
assign w5657 = ~w5411 & w5510;
assign w5658 = ~w5511 & ~w5657;
assign w5659 = (~w5655 & w33094) | (~w5655 & w33095) | (w33094 & w33095);
assign w5660 = (w5655 & w33096) | (w5655 & w33097) | (w33096 & w33097);
assign w5661 = (~w5483 & w33098) | (~w5483 & w33099) | (w33098 & w33099);
assign w5662 = ~w5487 & ~w5661;
assign w5663 = ~w5660 & w5662;
assign w5664 = (~w5487 & ~w5662) | (~w5487 & w33100) | (~w5662 & w33100);
assign w5665 = (~w5463 & w33101) | (~w5463 & w33102) | (w33101 & w33102);
assign w5666 = ~w5467 & ~w5665;
assign w5667 = ~w5664 & w5666;
assign w5668 = w5664 & ~w5666;
assign w5669 = ~w5667 & ~w5668;
assign w5670 = ~w2075 & w3957;
assign w5671 = (w4446 & ~w2235) | (w4446 & w33103) | (~w2235 & w33103);
assign w5672 = ~w2148 & w4068;
assign w5673 = ~w5671 & ~w5672;
assign w5674 = ~w5670 & w5673;
assign w5675 = (w5674 & ~w4962) | (w5674 & w33104) | (~w4962 & w33104);
assign w5676 = a_29 & ~w5675;
assign w5677 = (~w4962 & w33105) | (~w4962 & w33106) | (w33105 & w33106);
assign w5678 = ~w5676 & ~w5677;
assign w5679 = w5669 & w5678;
assign w5680 = (~w5667 & ~w5669) | (~w5667 & w33107) | (~w5669 & w33107);
assign w5681 = w5473 & ~w5680;
assign w5682 = ~w5473 & w5680;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = (w4068 & ~w2235) | (w4068 & w33108) | (~w2235 & w33108);
assign w5685 = ~w2148 & w3957;
assign w5686 = (w4446 & ~w3712) | (w4446 & w33109) | (~w3712 & w33109);
assign w5687 = w4070 & w5103;
assign w5688 = ~w5685 & w33110;
assign w5689 = (a_29 & w5687) | (a_29 & w33111) | (w5687 & w33111);
assign w5690 = ~w5687 & w33112;
assign w5691 = ~w5689 & ~w5690;
assign w5692 = w5683 & w5691;
assign w5693 = ~w5683 & ~w5691;
assign w5694 = ~w5692 & ~w5693;
assign w5695 = w5364 & w5694;
assign w5696 = ~w5364 & ~w5694;
assign w5697 = ~w5695 & ~w5696;
assign w5698 = ~w5669 & ~w5678;
assign w5699 = ~w5679 & ~w5698;
assign w5700 = (w5655 & w33113) | (w5655 & w33114) | (w33113 & w33114);
assign w5701 = ~w5659 & ~w5700;
assign w5702 = w1399 & ~w3403;
assign w5703 = w668 & ~w2306;
assign w5704 = (w1327 & ~w3538) | (w1327 & w33115) | (~w3538 & w33115);
assign w5705 = (~w5479 & w3547) | (~w5479 & w33116) | (w3547 & w33116);
assign w5706 = ~w5480 & ~w5705;
assign w5707 = ~w5703 & ~w5704;
assign w5708 = ~w5702 & w5707;
assign w5709 = (w5708 & ~w5706) | (w5708 & w33117) | (~w5706 & w33117);
assign w5710 = w5701 & ~w5709;
assign w5711 = ~w5701 & w5709;
assign w5712 = ~w5710 & ~w5711;
assign w5713 = ~w2075 & w4446;
assign w5714 = ~w2393 & w3957;
assign w5715 = ~w3615 & w4068;
assign w5716 = ~w5714 & ~w5715;
assign w5717 = ~w5713 & w5716;
assign w5718 = (w5717 & ~w5227) | (w5717 & w33118) | (~w5227 & w33118);
assign w5719 = a_29 & w5718;
assign w5720 = (w5227 & w33119) | (w5227 & w33120) | (w33119 & w33120);
assign w5721 = ~w5719 & ~w5720;
assign w5722 = w5712 & ~w5721;
assign w5723 = (~w5710 & ~w5712) | (~w5710 & w33121) | (~w5712 & w33121);
assign w5724 = w5660 & ~w5662;
assign w5725 = ~w5663 & ~w5724;
assign w5726 = w5723 & ~w5725;
assign w5727 = ~w5723 & w5725;
assign w5728 = ~w5726 & ~w5727;
assign w5729 = ~w2075 & w4068;
assign w5730 = ~w2148 & w4446;
assign w5731 = ~w3615 & w3957;
assign w5732 = ~w5730 & ~w5731;
assign w5733 = ~w5729 & w5732;
assign w5734 = (w5733 & ~w5242) | (w5733 & w33122) | (~w5242 & w33122);
assign w5735 = a_29 & ~w5734;
assign w5736 = (~w5242 & w33123) | (~w5242 & w33124) | (w33123 & w33124);
assign w5737 = ~w5735 & ~w5736;
assign w5738 = w5728 & ~w5737;
assign w5739 = (~w5726 & ~w5728) | (~w5726 & w33125) | (~w5728 & w33125);
assign w5740 = ~w5699 & ~w5739;
assign w5741 = (w4638 & ~w3658) | (w4638 & w33126) | (~w3658 & w33126);
assign w5742 = (w4666 & ~w2005) | (w4666 & w33127) | (~w2005 & w33127);
assign w5743 = (~w518 & ~w3712) | (~w518 & w33128) | (~w3712 & w33128);
assign w5744 = (w1226 & w4790) | (w1226 & w33129) | (w4790 & w33129);
assign w5745 = ~w5742 & ~w5743;
assign w5746 = ~w5741 & w5745;
assign w5747 = (a_26 & w5744) | (a_26 & w33130) | (w5744 & w33130);
assign w5748 = ~w5744 & w33131;
assign w5749 = ~w5747 & ~w5748;
assign w5750 = w5699 & w5739;
assign w5751 = ~w5740 & ~w5750;
assign w5752 = ~w5749 & w5751;
assign w5753 = (~w5740 & ~w5751) | (~w5740 & w33132) | (~w5751 & w33132);
assign w5754 = w5697 & w5753;
assign w5755 = ~w5697 & ~w5753;
assign w5756 = ~w5754 & ~w5755;
assign w5757 = ~w3813 & w5286;
assign w5758 = (w5016 & ~w1714) | (w5016 & w33133) | (~w1714 & w33133);
assign w5759 = (w5080 & ~w1807) | (w5080 & w33134) | (~w1807 & w33134);
assign w5760 = w4508 & w5017;
assign w5761 = ~w5757 & w33135;
assign w5762 = ~w5760 & w33136;
assign w5763 = (~a_23 & w5760) | (~a_23 & w33137) | (w5760 & w33137);
assign w5764 = ~w5762 & ~w5763;
assign w5765 = w5756 & ~w5764;
assign w5766 = (~w5754 & ~w5756) | (~w5754 & w33138) | (~w5756 & w33138);
assign w5767 = (~w5692 & ~w5694) | (~w5692 & w33139) | (~w5694 & w33139);
assign w5768 = (~w5471 & w5680) | (~w5471 & w33140) | (w5680 & w33140);
assign w5769 = ~w5236 & w5245;
assign w5770 = ~w5246 & ~w5769;
assign w5771 = (w4446 & ~w3658) | (w4446 & w33141) | (~w3658 & w33141);
assign w5772 = (w4068 & ~w3712) | (w4068 & w33142) | (~w3712 & w33142);
assign w5773 = (w3957 & ~w2235) | (w3957 & w33143) | (~w2235 & w33143);
assign w5774 = ~w5772 & ~w5773;
assign w5775 = ~w5771 & w5774;
assign w5776 = (w5775 & ~w4810) | (w5775 & w33144) | (~w4810 & w33144);
assign w5777 = a_29 & ~w5776;
assign w5778 = (~w4810 & w33145) | (~w4810 & w33146) | (w33145 & w33146);
assign w5779 = ~w5777 & ~w5778;
assign w5780 = w5770 & w5779;
assign w5781 = ~w5770 & ~w5779;
assign w5782 = ~w5780 & ~w5781;
assign w5783 = ~w5768 & w5782;
assign w5784 = w5768 & ~w5782;
assign w5785 = ~w5783 & ~w5784;
assign w5786 = (w4638 & ~w1913) | (w4638 & w33147) | (~w1913 & w33147);
assign w5787 = (~w518 & ~w2005) | (~w518 & w33148) | (~w2005 & w33148);
assign w5788 = (w4666 & ~w1714) | (w4666 & w33011) | (~w1714 & w33011);
assign w5789 = ~w5786 & ~w5787;
assign w5790 = ~w5788 & w5789;
assign w5791 = (w5790 & ~w4592) | (w5790 & w33149) | (~w4592 & w33149);
assign w5792 = a_26 & ~w5791;
assign w5793 = (~w4592 & w33150) | (~w4592 & w33151) | (w33150 & w33151);
assign w5794 = ~w5792 & ~w5793;
assign w5795 = w5785 & w5794;
assign w5796 = ~w5785 & ~w5794;
assign w5797 = ~w5795 & ~w5796;
assign w5798 = ~w5767 & w5797;
assign w5799 = w5767 & ~w5797;
assign w5800 = ~w5798 & ~w5799;
assign w5801 = (w5016 & ~w1807) | (w5016 & w33152) | (~w1807 & w33152);
assign w5802 = (w5286 & ~w1628) | (w5286 & w33153) | (~w1628 & w33153);
assign w5803 = ~w3813 & w5080;
assign w5804 = ~w5801 & ~w5802;
assign w5805 = ~w5803 & w5804;
assign w5806 = (w5805 & ~w4244) | (w5805 & w33154) | (~w4244 & w33154);
assign w5807 = a_23 & ~w5806;
assign w5808 = (~w4244 & w33155) | (~w4244 & w33156) | (w33155 & w33156);
assign w5809 = ~w5807 & ~w5808;
assign w5810 = w5800 & w5809;
assign w5811 = ~w5800 & ~w5809;
assign w5812 = ~w5810 & ~w5811;
assign w5813 = ~w5766 & w5812;
assign w5814 = w5766 & ~w5812;
assign w5815 = ~w5813 & ~w5814;
assign w5816 = w5300 & w5307;
assign w5817 = ~w1397 & w5816;
assign w5818 = ~w5300 & w5303;
assign w5819 = ~w1475 & w5818;
assign w5820 = (w5308 & ~w643) | (w5308 & w33157) | (~w643 & w33157);
assign w5821 = ~w5817 & ~w5820;
assign w5822 = ~w5819 & w5821;
assign w5823 = (w5822 & ~w4056) | (w5822 & w33158) | (~w4056 & w33158);
assign w5824 = a_20 & w5823;
assign w5825 = (w4056 & w33159) | (w4056 & w33160) | (w33159 & w33160);
assign w5826 = ~w5824 & ~w5825;
assign w5827 = w5815 & ~w5826;
assign w5828 = ~w5756 & w5764;
assign w5829 = ~w5765 & ~w5828;
assign w5830 = w5749 & ~w5751;
assign w5831 = ~w5752 & ~w5830;
assign w5832 = ~w5728 & w5737;
assign w5833 = ~w5738 & ~w5832;
assign w5834 = (w4666 & ~w3658) | (w4666 & w33161) | (~w3658 & w33161);
assign w5835 = (w4638 & ~w3712) | (w4638 & w33162) | (~w3712 & w33162);
assign w5836 = (~w518 & ~w2235) | (~w518 & w33163) | (~w2235 & w33163);
assign w5837 = ~w5835 & ~w5836;
assign w5838 = ~w5834 & w5837;
assign w5839 = (w5838 & ~w4810) | (w5838 & w33164) | (~w4810 & w33164);
assign w5840 = a_26 & ~w5839;
assign w5841 = (~w4810 & w33165) | (~w4810 & w33166) | (w33165 & w33166);
assign w5842 = ~w5840 & ~w5841;
assign w5843 = ~w5833 & w5842;
assign w5844 = ~w325 & ~w391;
assign w5845 = ~w468 & ~w896;
assign w5846 = w433 & w5845;
assign w5847 = w2336 & w3517;
assign w5848 = w3569 & w5844;
assign w5849 = w5847 & w5848;
assign w5850 = w1603 & w5846;
assign w5851 = w3207 & w4129;
assign w5852 = w5850 & w5851;
assign w5853 = w295 & w5849;
assign w5854 = w5852 & w5853;
assign w5855 = ~w403 & w1340;
assign w5856 = ~w207 & ~w423;
assign w5857 = ~w652 & w5856;
assign w5858 = ~w206 & w958;
assign w5859 = w1541 & w1686;
assign w5860 = w1967 & w2688;
assign w5861 = w5859 & w5860;
assign w5862 = w318 & w5858;
assign w5863 = w5855 & w5857;
assign w5864 = w5862 & w5863;
assign w5865 = w5562 & w5861;
assign w5866 = w5589 & w5865;
assign w5867 = w5864 & w5866;
assign w5868 = w2509 & w5854;
assign w5869 = w5867 & w5868;
assign w5870 = w4362 & w5869;
assign w5871 = w5578 & ~w5870;
assign w5872 = w2247 & w2275;
assign w5873 = w3796 & w5872;
assign w5874 = w1775 & w5873;
assign w5875 = ~w196 & ~w694;
assign w5876 = w3584 & w5875;
assign w5877 = w3733 & w4386;
assign w5878 = w5876 & w5877;
assign w5879 = w1385 & w1986;
assign w5880 = w3977 & w4156;
assign w5881 = w5879 & w5880;
assign w5882 = w1768 & w5878;
assign w5883 = w5881 & w5882;
assign w5884 = w1735 & w5874;
assign w5885 = w5883 & w5884;
assign w5886 = w1039 & w5885;
assign w5887 = w4923 & w5886;
assign w5888 = ~a_2 & ~w5887;
assign w5889 = a_2 & w5887;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = ~a_5 & w5890;
assign w5892 = (~w5888 & ~w5890) | (~w5888 & w33167) | (~w5890 & w33167);
assign w5893 = w5578 & ~w5892;
assign w5894 = ~w5578 & w5892;
assign w5895 = ~w5893 & ~w5894;
assign w5896 = w668 & ~w3326;
assign w5897 = (w1327 & ~w3267) | (w1327 & w33168) | (~w3267 & w33168);
assign w5898 = w1399 & ~w3196;
assign w5899 = ~w3269 & ~w3326;
assign w5900 = ~w3543 & ~w5899;
assign w5901 = (~w3058 & w33169) | (~w3058 & w33170) | (w33169 & w33170);
assign w5902 = (w3058 & w33171) | (w3058 & w33172) | (w33171 & w33172);
assign w5903 = ~w5901 & ~w5902;
assign w5904 = ~w5897 & ~w5898;
assign w5905 = ~w5896 & w5904;
assign w5906 = (w5905 & w5903) | (w5905 & w33173) | (w5903 & w33173);
assign w5907 = w5895 & ~w5906;
assign w5908 = ~w5578 & w5870;
assign w5909 = ~w5871 & ~w5908;
assign w5910 = (~w5906 & w33175) | (~w5906 & w33176) | (w33175 & w33176);
assign w5911 = (w5906 & w33177) | (w5906 & w33178) | (w33177 & w33178);
assign w5912 = a_8 & ~w5639;
assign w5913 = ~w5640 & ~w5912;
assign w5914 = ~w5911 & w5913;
assign w5915 = w5911 & ~w5913;
assign w5916 = ~w5914 & ~w5915;
assign w5917 = w668 & ~w3403;
assign w5918 = w1327 & ~w3475;
assign w5919 = w1399 & ~w3326;
assign w5920 = w3545 & ~w3551;
assign w5921 = w3326 & w3550;
assign w5922 = (~w5921 & w3328) | (~w5921 & w33179) | (w3328 & w33179);
assign w5923 = ~w5649 & w5922;
assign w5924 = ~w5917 & ~w5918;
assign w5925 = ~w5919 & w5924;
assign w5926 = (w5925 & ~w5923) | (w5925 & w33180) | (~w5923 & w33180);
assign w5927 = w5916 & ~w5926;
assign w5928 = (~w5914 & ~w5916) | (~w5914 & w33181) | (~w5916 & w33181);
assign w5929 = (~w5652 & w33182) | (~w5652 & w33183) | (w33182 & w33183);
assign w5930 = ~w5656 & ~w5929;
assign w5931 = ~w5928 & w5930;
assign w5932 = w5928 & ~w5930;
assign w5933 = ~w5931 & ~w5932;
assign w5934 = ~w2306 & w3957;
assign w5935 = ~w2393 & w4068;
assign w5936 = ~w3615 & w4446;
assign w5937 = ~w5934 & ~w5935;
assign w5938 = ~w5936 & w5937;
assign w5939 = (w5938 & ~w5463) | (w5938 & w33184) | (~w5463 & w33184);
assign w5940 = a_29 & ~w5939;
assign w5941 = (~w5463 & w33185) | (~w5463 & w33186) | (w33185 & w33186);
assign w5942 = ~w5940 & ~w5941;
assign w5943 = w5933 & w5942;
assign w5944 = (~w5931 & ~w5933) | (~w5931 & w33187) | (~w5933 & w33187);
assign w5945 = ~w5712 & w5721;
assign w5946 = ~w5722 & ~w5945;
assign w5947 = ~w5944 & w5946;
assign w5948 = w5944 & ~w5946;
assign w5949 = ~w5947 & ~w5948;
assign w5950 = (w4666 & ~w3712) | (w4666 & w33188) | (~w3712 & w33188);
assign w5951 = (w4638 & ~w2235) | (w4638 & w33189) | (~w2235 & w33189);
assign w5952 = ~w518 & ~w2148;
assign w5953 = ~w5950 & ~w5951;
assign w5954 = ~w5952 & w5953;
assign w5955 = (w5954 & ~w5103) | (w5954 & w33190) | (~w5103 & w33190);
assign w5956 = a_26 & ~w5955;
assign w5957 = (~w5103 & w33191) | (~w5103 & w33192) | (w33191 & w33192);
assign w5958 = ~w5956 & ~w5957;
assign w5959 = w5949 & w5958;
assign w5960 = (~w5947 & ~w5949) | (~w5947 & w33193) | (~w5949 & w33193);
assign w5961 = w5833 & ~w5842;
assign w5962 = ~w5843 & ~w5961;
assign w5963 = ~w5960 & w5962;
assign w5964 = (~w5843 & ~w5962) | (~w5843 & w33194) | (~w5962 & w33194);
assign w5965 = w5831 & w5964;
assign w5966 = ~w5831 & ~w5964;
assign w5967 = ~w5965 & ~w5966;
assign w5968 = (w5016 & ~w1913) | (w5016 & w33195) | (~w1913 & w33195);
assign w5969 = (w5080 & ~w1714) | (w5080 & w33196) | (~w1714 & w33196);
assign w5970 = (w5286 & ~w1807) | (w5286 & w33197) | (~w1807 & w33197);
assign w5971 = ~w5968 & ~w5969;
assign w5972 = ~w5970 & w5971;
assign w5973 = (w5972 & w4428) | (w5972 & w33198) | (w4428 & w33198);
assign w5974 = a_23 & w5973;
assign w5975 = (~w4428 & w33199) | (~w4428 & w33200) | (w33199 & w33200);
assign w5976 = ~w5974 & ~w5975;
assign w5977 = w5967 & w5976;
assign w5978 = (~w5965 & ~w5967) | (~w5965 & w33201) | (~w5967 & w33201);
assign w5979 = w5829 & w5978;
assign w5980 = ~w1475 & w5816;
assign w5981 = (w5308 & ~w1628) | (w5308 & w33202) | (~w1628 & w33202);
assign w5982 = (w5818 & ~w643) | (w5818 & w33203) | (~w643 & w33203);
assign w5983 = ~w5981 & ~w5982;
assign w5984 = ~w5980 & w5983;
assign w5985 = (w5984 & ~w4041) | (w5984 & w33204) | (~w4041 & w33204);
assign w5986 = a_20 & ~w5985;
assign w5987 = (~w4041 & w33205) | (~w4041 & w33206) | (w33205 & w33206);
assign w5988 = ~w5986 & ~w5987;
assign w5989 = ~w5829 & ~w5978;
assign w5990 = ~w5979 & ~w5989;
assign w5991 = w5988 & w5990;
assign w5992 = (~w5979 & ~w5990) | (~w5979 & w33207) | (~w5990 & w33207);
assign w5993 = ~w5815 & w5826;
assign w5994 = ~w5827 & ~w5993;
assign w5995 = ~w5992 & w5994;
assign w5996 = ~w5827 & ~w5995;
assign w5997 = ~w1397 & w5818;
assign w5998 = ~w1475 & w5308;
assign w5999 = (w5816 & ~w1308) | (w5816 & w33208) | (~w1308 & w33208);
assign w6000 = ~w5997 & ~w5998;
assign w6001 = ~w5999 & w6000;
assign w6002 = (w6001 & ~w3834) | (w6001 & w33209) | (~w3834 & w33209);
assign w6003 = a_20 & ~w6002;
assign w6004 = (~w3834 & w33210) | (~w3834 & w33211) | (w33210 & w33211);
assign w6005 = ~w6003 & ~w6004;
assign w6006 = ~w3813 & w5016;
assign w6007 = (w5080 & ~w1628) | (w5080 & w33196) | (~w1628 & w33196);
assign w6008 = (w5286 & ~w643) | (w5286 & w33212) | (~w643 & w33212);
assign w6009 = w4224 & w5017;
assign w6010 = ~w6006 & w33213;
assign w6011 = (a_23 & w6009) | (a_23 & w33214) | (w6009 & w33214);
assign w6012 = ~w6009 & w33215;
assign w6013 = ~w6011 & ~w6012;
assign w6014 = ~w5780 & ~w5783;
assign w6015 = ~w5252 & ~w5261;
assign w6016 = ~w5262 & ~w6015;
assign w6017 = w6014 & ~w6016;
assign w6018 = ~w6014 & w6016;
assign w6019 = ~w6017 & ~w6018;
assign w6020 = (~w518 & ~w1913) | (~w518 & w33216) | (~w1913 & w33216);
assign w6021 = (w4666 & ~w1807) | (w4666 & w33217) | (~w1807 & w33217);
assign w6022 = (w4638 & ~w1714) | (w4638 & w33006) | (~w1714 & w33006);
assign w6023 = ~w6020 & ~w6021;
assign w6024 = ~w6022 & w6023;
assign w6025 = (w6024 & w4428) | (w6024 & w33218) | (w4428 & w33218);
assign w6026 = a_26 & ~w6025;
assign w6027 = (w4428 & w33219) | (w4428 & w33220) | (w33219 & w33220);
assign w6028 = ~w6026 & ~w6027;
assign w6029 = w6019 & ~w6028;
assign w6030 = ~w6019 & w6028;
assign w6031 = ~w6029 & ~w6030;
assign w6032 = ~w5795 & ~w5798;
assign w6033 = w6031 & w6032;
assign w6034 = ~w6031 & ~w6032;
assign w6035 = ~w6033 & ~w6034;
assign w6036 = ~w6013 & w6035;
assign w6037 = w6013 & ~w6035;
assign w6038 = ~w6036 & ~w6037;
assign w6039 = ~w5810 & ~w5813;
assign w6040 = ~w6038 & ~w6039;
assign w6041 = w6038 & w6039;
assign w6042 = ~w6040 & ~w6041;
assign w6043 = w6005 & w6042;
assign w6044 = ~w6005 & ~w6042;
assign w6045 = ~w6043 & ~w6044;
assign w6046 = w5996 & ~w6045;
assign w6047 = ~w5996 & w6045;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = ~a_16 & a_17;
assign w6050 = a_16 & ~a_17;
assign w6051 = ~w6049 & ~w6050;
assign w6052 = ~a_14 & ~a_15;
assign w6053 = a_14 & a_15;
assign w6054 = ~w6052 & ~w6053;
assign w6055 = ~a_15 & ~a_16;
assign w6056 = a_15 & a_16;
assign w6057 = ~w6055 & ~w6056;
assign w6058 = ~w6054 & ~w6057;
assign w6059 = ~w6051 & w6058;
assign w6060 = (w6059 & ~w3904) | (w6059 & w33221) | (~w3904 & w33221);
assign w6061 = ~w6054 & w6057;
assign w6062 = ~w3958 & w6061;
assign w6063 = ~w6051 & w6054;
assign w6064 = ~w6060 & ~w6062;
assign w6065 = (w6064 & ~w4073) | (w6064 & w33222) | (~w4073 & w33222);
assign w6066 = a_17 & ~w6065;
assign w6067 = (~w4073 & w33223) | (~w4073 & w33224) | (w33223 & w33224);
assign w6068 = ~w6066 & ~w6067;
assign w6069 = w6048 & ~w6068;
assign w6070 = ~w6048 & w6068;
assign w6071 = ~w6069 & ~w6070;
assign w6072 = ~w5967 & ~w5976;
assign w6073 = ~w5977 & ~w6072;
assign w6074 = w5960 & ~w5962;
assign w6075 = ~w5963 & ~w6074;
assign w6076 = (w5080 & ~w1913) | (w5080 & w33225) | (~w1913 & w33225);
assign w6077 = (w5016 & ~w2005) | (w5016 & w33226) | (~w2005 & w33226);
assign w6078 = (w5286 & ~w1714) | (w5286 & w33153) | (~w1714 & w33153);
assign w6079 = ~w6076 & ~w6077;
assign w6080 = ~w6078 & w6079;
assign w6081 = (w6080 & ~w4592) | (w6080 & w33227) | (~w4592 & w33227);
assign w6082 = a_23 & w6081;
assign w6083 = (w4592 & w33228) | (w4592 & w33229) | (w33228 & w33229);
assign w6084 = ~w6082 & ~w6083;
assign w6085 = w6075 & ~w6084;
assign w6086 = ~w5949 & ~w5958;
assign w6087 = ~w5959 & ~w6086;
assign w6088 = ~w5916 & w5926;
assign w6089 = ~w5927 & ~w6088;
assign w6090 = ~w2306 & w4068;
assign w6091 = (w3957 & ~w3538) | (w3957 & w33230) | (~w3538 & w33230);
assign w6092 = ~w2393 & w4446;
assign w6093 = ~w6090 & ~w6091;
assign w6094 = ~w6092 & w6093;
assign w6095 = (w6094 & ~w5483) | (w6094 & w33231) | (~w5483 & w33231);
assign w6096 = a_29 & ~w6095;
assign w6097 = (~w5483 & w33232) | (~w5483 & w33233) | (w33232 & w33233);
assign w6098 = ~w6096 & ~w6097;
assign w6099 = w6089 & w6098;
assign w6100 = (w5906 & w33234) | (w5906 & w33235) | (w33234 & w33235);
assign w6101 = ~w5910 & ~w6100;
assign w6102 = w668 & ~w3475;
assign w6103 = (w1399 & ~w3267) | (w1399 & w33236) | (~w3267 & w33236);
assign w6104 = w1327 & ~w3326;
assign w6105 = ~w3542 & ~w3549;
assign w6106 = (w6105 & w3328) | (w6105 & w33237) | (w3328 & w33237);
assign w6107 = ~w3328 & w33238;
assign w6108 = ~w6106 & ~w6107;
assign w6109 = ~w6102 & ~w6103;
assign w6110 = ~w6104 & w6109;
assign w6111 = (w6110 & ~w6108) | (w6110 & w33239) | (~w6108 & w33239);
assign w6112 = w6101 & ~w6111;
assign w6113 = ~w6101 & w6111;
assign w6114 = ~w6112 & ~w6113;
assign w6115 = ~w622 & w1238;
assign w6116 = ~w260 & ~w406;
assign w6117 = ~w88 & ~w125;
assign w6118 = ~w475 & ~w1077;
assign w6119 = w669 & w6118;
assign w6120 = w6116 & w6117;
assign w6121 = w6119 & w6120;
assign w6122 = w1606 & w6121;
assign w6123 = ~w131 & ~w362;
assign w6124 = ~w696 & w6123;
assign w6125 = w2881 & w4850;
assign w6126 = w6124 & w6125;
assign w6127 = w2190 & w5414;
assign w6128 = w5489 & w6115;
assign w6129 = w6127 & w6128;
assign w6130 = w427 & w6126;
assign w6131 = w2092 & w6130;
assign w6132 = w6122 & w6129;
assign w6133 = w6131 & w6132;
assign w6134 = w1599 & w6133;
assign w6135 = w2736 & w3115;
assign w6136 = w6134 & w6135;
assign w6137 = a_2 & ~w6136;
assign w6138 = ~w694 & w1987;
assign w6139 = ~w380 & w4094;
assign w6140 = w6138 & w6139;
assign w6141 = ~w1953 & w2317;
assign w6142 = w3493 & w3569;
assign w6143 = w4393 & w6142;
assign w6144 = w4548 & w6141;
assign w6145 = w4730 & w6144;
assign w6146 = w226 & w6143;
assign w6147 = w1532 & w1780;
assign w6148 = w6140 & w6147;
assign w6149 = w6145 & w6146;
assign w6150 = w1006 & w6149;
assign w6151 = w1678 & w6148;
assign w6152 = w6150 & w6151;
assign w6153 = w2642 & w6152;
assign w6154 = a_2 & ~w6153;
assign w6155 = ~w218 & ~w400;
assign w6156 = ~w156 & ~w251;
assign w6157 = ~w256 & ~w279;
assign w6158 = w6156 & w6157;
assign w6159 = w2332 & w2707;
assign w6160 = w3275 & w6155;
assign w6161 = w6159 & w6160;
assign w6162 = w2164 & w6158;
assign w6163 = w2190 & w2616;
assign w6164 = w5491 & w6163;
assign w6165 = w6161 & w6162;
assign w6166 = w5515 & w6165;
assign w6167 = w6164 & w6166;
assign w6168 = ~w907 & ~w944;
assign w6169 = ~w254 & ~w568;
assign w6170 = w370 & w6169;
assign w6171 = w6168 & w6170;
assign w6172 = w9 & w1952;
assign w6173 = w215 & ~w6172;
assign w6174 = w545 & w990;
assign w6175 = w1693 & w2925;
assign w6176 = w5172 & w6175;
assign w6177 = w6173 & w6174;
assign w6178 = w1099 & w6177;
assign w6179 = w6171 & w6176;
assign w6180 = w6178 & w6179;
assign w6181 = w1086 & w1136;
assign w6182 = w6180 & w6181;
assign w6183 = w6167 & w6182;
assign w6184 = w3601 & w6183;
assign w6185 = a_2 & ~w6184;
assign w6186 = ~a_2 & w6184;
assign w6187 = ~w6185 & ~w6186;
assign w6188 = w3049 & w3198;
assign w6189 = ~w3058 & ~w6188;
assign w6190 = ~w2924 & w3055;
assign w6191 = ~w2920 & w6190;
assign w6192 = ~w3052 & ~w3198;
assign w6193 = ~w6191 & w6192;
assign w6194 = w6189 & ~w6193;
assign w6195 = w1399 & ~w2917;
assign w6196 = w668 & ~w3049;
assign w6197 = w1327 & ~w3007;
assign w6198 = ~w6195 & ~w6196;
assign w6199 = ~w6197 & w6198;
assign w6200 = (w6194 & w32435) | (w6194 & w32436) | (w32435 & w32436);
assign w6201 = ~a_2 & w6153;
assign w6202 = ~w6154 & ~w6201;
assign w6203 = (w6194 & w33242) | (w6194 & w33243) | (w33242 & w33243);
assign w6204 = ~a_2 & w6136;
assign w6205 = ~w6137 & ~w6204;
assign w6206 = (w6205 & w6203) | (w6205 & w33244) | (w6203 & w33244);
assign w6207 = a_5 & ~w5890;
assign w6208 = ~w5891 & ~w6207;
assign w6209 = (w6203 & w33247) | (w6203 & w33248) | (w33247 & w33248);
assign w6210 = (~w6203 & w33249) | (~w6203 & w33250) | (w33249 & w33250);
assign w6211 = ~w6209 & ~w6210;
assign w6212 = (w668 & ~w3267) | (w668 & w33251) | (~w3267 & w33251);
assign w6213 = w1327 & ~w3196;
assign w6214 = w1399 & ~w3139;
assign w6215 = ~w3197 & ~w3204;
assign w6216 = ~w3200 & w6215;
assign w6217 = ~w3197 & w3271;
assign w6218 = ~w6216 & w6217;
assign w6219 = ~w3205 & w6218;
assign w6220 = ~w6188 & w6218;
assign w6221 = ~w3058 & w6220;
assign w6222 = ~w6219 & ~w6221;
assign w6223 = w6222 & w33252;
assign w6224 = ~w6212 & ~w6213;
assign w6225 = ~w6214 & w6224;
assign w6226 = ~w6223 & w6225;
assign w6227 = w6211 & ~w6226;
assign w6228 = (~w6209 & ~w6211) | (~w6209 & w33253) | (~w6211 & w33253);
assign w6229 = (w5903 & w33254) | (w5903 & w33255) | (w33254 & w33255);
assign w6230 = ~w5907 & ~w6229;
assign w6231 = ~w6228 & w6230;
assign w6232 = w6228 & ~w6230;
assign w6233 = ~w6231 & ~w6232;
assign w6234 = ~w3403 & w4068;
assign w6235 = (w4446 & ~w3538) | (w4446 & w33256) | (~w3538 & w33256);
assign w6236 = ~w3475 & w3957;
assign w6237 = ~w6234 & ~w6235;
assign w6238 = ~w6236 & w6237;
assign w6239 = (w6238 & ~w5652) | (w6238 & w33257) | (~w5652 & w33257);
assign w6240 = a_29 & w6239;
assign w6241 = (w5652 & w33258) | (w5652 & w33259) | (w33258 & w33259);
assign w6242 = ~w6240 & ~w6241;
assign w6243 = w6233 & ~w6242;
assign w6244 = (~w6231 & ~w6233) | (~w6231 & w33260) | (~w6233 & w33260);
assign w6245 = w6114 & ~w6244;
assign w6246 = (~w6112 & w6244) | (~w6112 & w33261) | (w6244 & w33261);
assign w6247 = ~w6089 & ~w6098;
assign w6248 = ~w6099 & ~w6247;
assign w6249 = ~w6246 & w6248;
assign w6250 = ~w6099 & ~w6249;
assign w6251 = ~w5933 & ~w5942;
assign w6252 = ~w5943 & ~w6251;
assign w6253 = w6250 & ~w6252;
assign w6254 = ~w6250 & w6252;
assign w6255 = ~w6253 & ~w6254;
assign w6256 = ~w518 & ~w2075;
assign w6257 = (w4666 & ~w2235) | (w4666 & w33262) | (~w2235 & w33262);
assign w6258 = ~w2148 & w4638;
assign w6259 = ~w6257 & ~w6258;
assign w6260 = ~w6256 & w6259;
assign w6261 = (w6260 & ~w4962) | (w6260 & w33263) | (~w4962 & w33263);
assign w6262 = a_26 & ~w6261;
assign w6263 = (~w4962 & w33264) | (~w4962 & w33265) | (w33264 & w33265);
assign w6264 = ~w6262 & ~w6263;
assign w6265 = w6255 & ~w6264;
assign w6266 = (~w6253 & ~w6255) | (~w6253 & w33266) | (~w6255 & w33266);
assign w6267 = w6087 & w6266;
assign w6268 = (w5016 & ~w3658) | (w5016 & w33267) | (~w3658 & w33267);
assign w6269 = (w5080 & ~w2005) | (w5080 & w33268) | (~w2005 & w33268);
assign w6270 = (w5286 & ~w1913) | (w5286 & w33269) | (~w1913 & w33269);
assign w6271 = ~w6269 & ~w6270;
assign w6272 = ~w6268 & w6271;
assign w6273 = (w6272 & w4578) | (w6272 & w33270) | (w4578 & w33270);
assign w6274 = a_23 & ~w6273;
assign w6275 = (w4578 & w33271) | (w4578 & w33272) | (w33271 & w33272);
assign w6276 = ~w6274 & ~w6275;
assign w6277 = ~w6087 & ~w6266;
assign w6278 = ~w6267 & ~w6277;
assign w6279 = w6276 & w6278;
assign w6280 = (~w6267 & ~w6278) | (~w6267 & w33273) | (~w6278 & w33273);
assign w6281 = ~w6075 & w6084;
assign w6282 = ~w6085 & ~w6281;
assign w6283 = ~w6280 & w6282;
assign w6284 = (~w6085 & ~w6282) | (~w6085 & w33274) | (~w6282 & w33274);
assign w6285 = ~w6073 & ~w6284;
assign w6286 = w6073 & w6284;
assign w6287 = ~w6285 & ~w6286;
assign w6288 = ~w3813 & w5308;
assign w6289 = (w5816 & ~w643) | (w5816 & w33275) | (~w643 & w33275);
assign w6290 = (w5818 & ~w1628) | (w5818 & w33276) | (~w1628 & w33276);
assign w6291 = w4224 & w5309;
assign w6292 = ~w6288 & w33277;
assign w6293 = (a_20 & w6291) | (a_20 & w33278) | (w6291 & w33278);
assign w6294 = ~w6291 & w33279;
assign w6295 = ~w6293 & ~w6294;
assign w6296 = w6287 & w6295;
assign w6297 = (~w6285 & ~w6287) | (~w6285 & w33280) | (~w6287 & w33280);
assign w6298 = ~w5988 & ~w5990;
assign w6299 = ~w5991 & ~w6298;
assign w6300 = ~w6297 & w6299;
assign w6301 = w6297 & ~w6299;
assign w6302 = ~w6300 & ~w6301;
assign w6303 = ~w1397 & w6059;
assign w6304 = w6051 & w6054;
assign w6305 = (w6304 & ~w3904) | (w6304 & w33281) | (~w3904 & w33281);
assign w6306 = (w6061 & ~w1308) | (w6061 & w33282) | (~w1308 & w33282);
assign w6307 = ~w6303 & ~w6306;
assign w6308 = ~w6305 & w6307;
assign w6309 = (w6308 & ~w3964) | (w6308 & w33283) | (~w3964 & w33283);
assign w6310 = a_17 & ~w6309;
assign w6311 = (~w3964 & w33284) | (~w3964 & w33285) | (w33284 & w33285);
assign w6312 = ~w6310 & ~w6311;
assign w6313 = w6302 & w6312;
assign w6314 = (~w6300 & ~w6302) | (~w6300 & w33286) | (~w6302 & w33286);
assign w6315 = (w6061 & ~w3904) | (w6061 & w33287) | (~w3904 & w33287);
assign w6316 = ~w3958 & w6304;
assign w6317 = (w6059 & ~w1308) | (w6059 & w33288) | (~w1308 & w33288);
assign w6318 = ~w6316 & ~w6317;
assign w6319 = ~w6315 & w6318;
assign w6320 = (w6319 & ~w3943) | (w6319 & w33289) | (~w3943 & w33289);
assign w6321 = a_17 & ~w6320;
assign w6322 = (~w3943 & w33290) | (~w3943 & w33291) | (w33290 & w33291);
assign w6323 = ~w6321 & ~w6322;
assign w6324 = ~w6314 & w6323;
assign w6325 = w5992 & ~w5994;
assign w6326 = ~w5995 & ~w6325;
assign w6327 = w6314 & ~w6323;
assign w6328 = ~w6324 & ~w6327;
assign w6329 = w6326 & w6328;
assign w6330 = (~w6324 & ~w6328) | (~w6324 & w33292) | (~w6328 & w33292);
assign w6331 = w6071 & w6330;
assign w6332 = w6280 & ~w6282;
assign w6333 = ~w6283 & ~w6332;
assign w6334 = (w5308 & ~w1807) | (w5308 & w33293) | (~w1807 & w33293);
assign w6335 = (w5816 & ~w1628) | (w5816 & w33294) | (~w1628 & w33294);
assign w6336 = ~w3813 & w5818;
assign w6337 = ~w6334 & ~w6335;
assign w6338 = ~w6336 & w6337;
assign w6339 = (w6338 & ~w4244) | (w6338 & w33295) | (~w4244 & w33295);
assign w6340 = a_20 & ~w6339;
assign w6341 = (~w4244 & w33296) | (~w4244 & w33297) | (w33296 & w33297);
assign w6342 = ~w6340 & ~w6341;
assign w6343 = w6333 & w6342;
assign w6344 = ~w6276 & ~w6278;
assign w6345 = ~w6279 & ~w6344;
assign w6346 = ~w6255 & w6264;
assign w6347 = ~w6265 & ~w6346;
assign w6348 = w6246 & ~w6248;
assign w6349 = ~w6249 & ~w6348;
assign w6350 = ~w2075 & w4638;
assign w6351 = ~w518 & ~w3615;
assign w6352 = ~w2148 & w4666;
assign w6353 = ~w6351 & ~w6352;
assign w6354 = ~w6350 & w6353;
assign w6355 = (w6354 & ~w5242) | (w6354 & w33298) | (~w5242 & w33298);
assign w6356 = a_26 & ~w6355;
assign w6357 = (~w5242 & w33299) | (~w5242 & w33300) | (w33299 & w33300);
assign w6358 = ~w6356 & ~w6357;
assign w6359 = w6349 & w6358;
assign w6360 = ~w6114 & w6244;
assign w6361 = ~w6245 & ~w6360;
assign w6362 = ~w3403 & w3957;
assign w6363 = ~w2306 & w4446;
assign w6364 = (w4068 & ~w3538) | (w4068 & w33301) | (~w3538 & w33301);
assign w6365 = ~w6363 & ~w6364;
assign w6366 = ~w6362 & w6365;
assign w6367 = (w6366 & ~w5706) | (w6366 & w33302) | (~w5706 & w33302);
assign w6368 = a_29 & w6367;
assign w6369 = (w5706 & w33303) | (w5706 & w33304) | (w33303 & w33304);
assign w6370 = ~w6368 & ~w6369;
assign w6371 = w6361 & ~w6370;
assign w6372 = ~w2075 & w4666;
assign w6373 = ~w3615 & w4638;
assign w6374 = ~w518 & ~w2393;
assign w6375 = ~w6373 & ~w6374;
assign w6376 = ~w6372 & w6375;
assign w6377 = (w6376 & ~w5227) | (w6376 & w33305) | (~w5227 & w33305);
assign w6378 = a_26 & ~w6377;
assign w6379 = (~w5227 & w33306) | (~w5227 & w33307) | (w33306 & w33307);
assign w6380 = ~w6378 & ~w6379;
assign w6381 = ~w6361 & w6370;
assign w6382 = ~w6371 & ~w6381;
assign w6383 = w6380 & w6382;
assign w6384 = (~w6371 & ~w6382) | (~w6371 & w33308) | (~w6382 & w33308);
assign w6385 = ~w6349 & ~w6358;
assign w6386 = ~w6359 & ~w6385;
assign w6387 = ~w6384 & w6386;
assign w6388 = ~w6359 & ~w6387;
assign w6389 = w6347 & w6388;
assign w6390 = ~w6347 & ~w6388;
assign w6391 = ~w6389 & ~w6390;
assign w6392 = (w5080 & ~w3658) | (w5080 & w33309) | (~w3658 & w33309);
assign w6393 = (w5286 & ~w2005) | (w5286 & w33310) | (~w2005 & w33310);
assign w6394 = (w5016 & ~w3712) | (w5016 & w33311) | (~w3712 & w33311);
assign w6395 = (w5017 & w4790) | (w5017 & w33312) | (w4790 & w33312);
assign w6396 = ~w6393 & ~w6394;
assign w6397 = ~w6392 & w6396;
assign w6398 = (a_23 & w6395) | (a_23 & w33313) | (w6395 & w33313);
assign w6399 = ~w6395 & w33314;
assign w6400 = ~w6398 & ~w6399;
assign w6401 = w6391 & ~w6400;
assign w6402 = (~w6389 & ~w6391) | (~w6389 & w33315) | (~w6391 & w33315);
assign w6403 = w6345 & w6402;
assign w6404 = ~w3813 & w5816;
assign w6405 = (w5818 & ~w1807) | (w5818 & w33316) | (~w1807 & w33316);
assign w6406 = (w5308 & ~w1714) | (w5308 & w33202) | (~w1714 & w33202);
assign w6407 = w4508 & w5309;
assign w6408 = ~w6404 & w33317;
assign w6409 = (a_20 & w6407) | (a_20 & w33318) | (w6407 & w33318);
assign w6410 = ~w6407 & w33319;
assign w6411 = ~w6409 & ~w6410;
assign w6412 = ~w6345 & ~w6402;
assign w6413 = ~w6403 & ~w6412;
assign w6414 = w6411 & w6413;
assign w6415 = (~w6403 & ~w6413) | (~w6403 & w33320) | (~w6413 & w33320);
assign w6416 = ~w6333 & ~w6342;
assign w6417 = ~w6343 & ~w6416;
assign w6418 = ~w6415 & w6417;
assign w6419 = (~w6343 & ~w6417) | (~w6343 & w33321) | (~w6417 & w33321);
assign w6420 = ~w6287 & ~w6295;
assign w6421 = ~w6296 & ~w6420;
assign w6422 = w6419 & ~w6421;
assign w6423 = ~w6419 & w6421;
assign w6424 = ~w6422 & ~w6423;
assign w6425 = ~w1397 & w6061;
assign w6426 = ~w1475 & w6059;
assign w6427 = (w6304 & ~w1308) | (w6304 & w33322) | (~w1308 & w33322);
assign w6428 = ~w6425 & ~w6426;
assign w6429 = ~w6427 & w6428;
assign w6430 = (w6429 & ~w3834) | (w6429 & w33323) | (~w3834 & w33323);
assign w6431 = a_17 & ~w6430;
assign w6432 = (~w3834 & w33324) | (~w3834 & w33325) | (w33324 & w33325);
assign w6433 = ~w6431 & ~w6432;
assign w6434 = w6424 & ~w6433;
assign w6435 = (~w6422 & ~w6424) | (~w6422 & w33326) | (~w6424 & w33326);
assign w6436 = ~a_13 & a_14;
assign w6437 = a_13 & ~a_14;
assign w6438 = ~w6436 & ~w6437;
assign w6439 = ~a_11 & ~a_12;
assign w6440 = a_11 & a_12;
assign w6441 = ~w6439 & ~w6440;
assign w6442 = ~a_12 & ~a_13;
assign w6443 = a_12 & a_13;
assign w6444 = ~w6442 & ~w6443;
assign w6445 = ~w6441 & ~w6444;
assign w6446 = ~w6438 & w6445;
assign w6447 = ~w6438 & w6441;
assign w6448 = (~w3828 & w33329) | (~w3828 & w33330) | (w33329 & w33330);
assign w6449 = ~w6448 & w33331;
assign w6450 = (a_14 & w6448) | (a_14 & w33332) | (w6448 & w33332);
assign w6451 = ~w6449 & ~w6450;
assign w6452 = w6435 & ~w6451;
assign w6453 = ~w6435 & w6451;
assign w6454 = ~w6452 & ~w6453;
assign w6455 = ~w6302 & ~w6312;
assign w6456 = ~w6313 & ~w6455;
assign w6457 = w6454 & w6456;
assign w6458 = (~w6452 & ~w6454) | (~w6452 & w33333) | (~w6454 & w33333);
assign w6459 = ~w6326 & ~w6328;
assign w6460 = ~w6329 & ~w6459;
assign w6461 = ~w6458 & w6460;
assign w6462 = ~w6391 & w6400;
assign w6463 = ~w6401 & ~w6462;
assign w6464 = w6384 & ~w6386;
assign w6465 = ~w6387 & ~w6464;
assign w6466 = (w5286 & ~w3658) | (w5286 & w33334) | (~w3658 & w33334);
assign w6467 = (w5016 & ~w2235) | (w5016 & w33335) | (~w2235 & w33335);
assign w6468 = (w5080 & ~w3712) | (w5080 & w33336) | (~w3712 & w33336);
assign w6469 = ~w6467 & ~w6468;
assign w6470 = ~w6466 & w6469;
assign w6471 = (w6470 & ~w4810) | (w6470 & w33337) | (~w4810 & w33337);
assign w6472 = a_23 & w6471;
assign w6473 = (w4810 & w33338) | (w4810 & w33339) | (w33338 & w33339);
assign w6474 = ~w6472 & ~w6473;
assign w6475 = w6465 & ~w6474;
assign w6476 = ~w6380 & ~w6382;
assign w6477 = ~w6383 & ~w6476;
assign w6478 = ~w6233 & w6242;
assign w6479 = ~w6243 & ~w6478;
assign w6480 = ~w6203 & w33340;
assign w6481 = ~w6206 & ~w6480;
assign w6482 = w668 & ~w3196;
assign w6483 = w1327 & ~w3139;
assign w6484 = w1399 & ~w3049;
assign w6485 = w3201 & ~w6215;
assign w6486 = w3196 & w3203;
assign w6487 = ~w6216 & ~w6486;
assign w6488 = ~w3197 & w3205;
assign w6489 = (w6488 & w3058) | (w6488 & w31572) | (w3058 & w31572);
assign w6490 = (w6487 & w3058) | (w6487 & w31573) | (w3058 & w31573);
assign w6491 = ~w6489 & w6490;
assign w6492 = ~w6482 & ~w6483;
assign w6493 = ~w6484 & w6492;
assign w6494 = (w6493 & ~w6491) | (w6493 & w33341) | (~w6491 & w33341);
assign w6495 = w6481 & ~w6494;
assign w6496 = (~w6194 & w33342) | (~w6194 & w33343) | (w33342 & w33343);
assign w6497 = ~w6203 & ~w6496;
assign w6498 = w668 & ~w3139;
assign w6499 = w1327 & ~w3049;
assign w6500 = w1399 & ~w3007;
assign w6501 = ~w3050 & ~w3198;
assign w6502 = ~w3199 & ~w3203;
assign w6503 = ~w3058 & w31574;
assign w6504 = (~w6502 & w3058) | (~w6502 & w31575) | (w3058 & w31575);
assign w6505 = ~w6503 & ~w6504;
assign w6506 = ~w6498 & ~w6499;
assign w6507 = ~w6500 & w6506;
assign w6508 = (w6507 & w6505) | (w6507 & w33344) | (w6505 & w33344);
assign w6509 = w6497 & ~w6508;
assign w6510 = ~w6497 & w6508;
assign w6511 = ~w6509 & ~w6510;
assign w6512 = ~w237 & ~w322;
assign w6513 = ~w366 & ~w380;
assign w6514 = w6512 & w6513;
assign w6515 = w2008 & w2604;
assign w6516 = w2646 & w3212;
assign w6517 = w4346 & w5185;
assign w6518 = w5388 & w6517;
assign w6519 = w6515 & w6516;
assign w6520 = w1762 & w6514;
assign w6521 = w6519 & w6520;
assign w6522 = w176 & w6518;
assign w6523 = w6521 & w6522;
assign w6524 = w3463 & w6523;
assign w6525 = ~w125 & w1726;
assign w6526 = w5563 & w6525;
assign w6527 = w1947 & w2528;
assign w6528 = w2552 & w3009;
assign w6529 = w3274 & w3796;
assign w6530 = w6528 & w6529;
assign w6531 = ~w519 & w6527;
assign w6532 = w1017 & w2020;
assign w6533 = w6531 & w6532;
assign w6534 = w92 & w6530;
assign w6535 = w6526 & w6534;
assign w6536 = w6533 & w6535;
assign w6537 = w4910 & w6536;
assign w6538 = w4896 & w6524;
assign w6539 = w6537 & w6538;
assign w6540 = w668 & ~w3007;
assign w6541 = w1399 & ~w2835;
assign w6542 = w1327 & ~w2917;
assign w6543 = (~w3053 & w2923) | (~w3053 & w31576) | (w2923 & w31576);
assign w6544 = ~w3054 & ~w3198;
assign w6545 = (w6544 & w2920) | (w6544 & w31577) | (w2920 & w31577);
assign w6546 = ~w2920 & w31578;
assign w6547 = ~w6545 & ~w6546;
assign w6548 = ~w6540 & ~w6541;
assign w6549 = ~w6542 & w6548;
assign w6550 = (w6549 & w6547) | (w6549 & w33345) | (w6547 & w33345);
assign w6551 = w6539 & w6550;
assign w6552 = ~w2837 & ~w2922;
assign w6553 = w2680 & w31579;
assign w6554 = w1478 & ~w6552;
assign w6555 = ~w2680 & w6554;
assign w6556 = (w668 & ~w2766) | (w668 & w33346) | (~w2766 & w33346);
assign w6557 = w1399 & ~w2677;
assign w6558 = w1327 & ~w2546;
assign w6559 = ~w6556 & ~w6557;
assign w6560 = ~w6558 & w6559;
assign w6561 = ~w6555 & w6560;
assign w6562 = ~w16 & ~w86;
assign w6563 = ~w288 & w6562;
assign w6564 = w141 & w222;
assign w6565 = w364 & w3570;
assign w6566 = w6564 & w6565;
assign w6567 = w940 & w6563;
assign w6568 = w4513 & w6567;
assign w6569 = w6566 & w6568;
assign w6570 = ~w146 & ~w281;
assign w6571 = ~w195 & ~w589;
assign w6572 = ~w1953 & w6571;
assign w6573 = w908 & w4818;
assign w6574 = ~w89 & ~w216;
assign w6575 = ~w341 & ~w2331;
assign w6576 = w6574 & w6575;
assign w6577 = ~w4404 & w6576;
assign w6578 = w215 & w709;
assign w6579 = w988 & w1419;
assign w6580 = w2219 & w2371;
assign w6581 = w3154 & w6570;
assign w6582 = w6580 & w6581;
assign w6583 = w6578 & w6579;
assign w6584 = w2403 & w4160;
assign w6585 = w6572 & w6573;
assign w6586 = w6584 & w6585;
assign w6587 = w6582 & w6583;
assign w6588 = w6577 & w6587;
assign w6589 = w6586 & w6588;
assign w6590 = w6569 & w6589;
assign w6591 = w2964 & w6590;
assign w6592 = (~w6591 & ~w6561) | (~w6591 & w31580) | (~w6561 & w31580);
assign w6593 = w6561 & w31581;
assign w6594 = ~w6592 & ~w6593;
assign w6595 = ~w2480 & w2601;
assign w6596 = w1478 & w2677;
assign w6597 = w6595 & w6596;
assign w6598 = w1478 & ~w2677;
assign w6599 = ~w6595 & w6598;
assign w6600 = (w1327 & ~w2479) | (w1327 & w31582) | (~w2479 & w31582);
assign w6601 = (w1399 & ~w2600) | (w1399 & w31583) | (~w2600 & w31583);
assign w6602 = w668 & ~w2677;
assign w6603 = ~w6600 & ~w6601;
assign w6604 = ~w6602 & w6603;
assign w6605 = ~w6597 & ~w6599;
assign w6606 = w962 & w1489;
assign w6607 = ~w580 & w1196;
assign w6608 = w2063 & w4151;
assign w6609 = w6607 & w6608;
assign w6610 = w2738 & w6609;
assign w6611 = ~w357 & w1720;
assign w6612 = ~w30 & ~w473;
assign w6613 = w1482 & w6612;
assign w6614 = ~w363 & ~w396;
assign w6615 = ~w399 & ~w423;
assign w6616 = ~w732 & w6615;
assign w6617 = w1073 & w6614;
assign w6618 = w2804 & w3674;
assign w6619 = w4104 & w6618;
assign w6620 = w6616 & w6617;
assign w6621 = w1773 & w6606;
assign w6622 = w6611 & w6613;
assign w6623 = w6621 & w6622;
assign w6624 = w6619 & w6620;
assign w6625 = w6623 & w6624;
assign w6626 = w6610 & w6625;
assign w6627 = w3089 & w6626;
assign w6628 = w4176 & w4753;
assign w6629 = w6627 & w6628;
assign w6630 = (~w6629 & ~w6605) | (~w6629 & w31584) | (~w6605 & w31584);
assign w6631 = w728 & w33347;
assign w6632 = ~w207 & ~w404;
assign w6633 = w4274 & w6632;
assign w6634 = w1659 & w6633;
assign w6635 = ~w267 & ~w385;
assign w6636 = ~w339 & ~w473;
assign w6637 = ~w476 & ~w590;
assign w6638 = w6636 & w6637;
assign w6639 = w941 & w3488;
assign w6640 = w6638 & w6639;
assign w6641 = w1342 & w6640;
assign w6642 = ~w652 & ~w671;
assign w6643 = w935 & w6642;
assign w6644 = ~w163 & ~w369;
assign w6645 = ~w1965 & w6644;
assign w6646 = w774 & w1078;
assign w6647 = w2276 & w2399;
assign w6648 = w2516 & w2715;
assign w6649 = w3686 & w6635;
assign w6650 = w6648 & w6649;
assign w6651 = w6646 & w6647;
assign w6652 = w546 & w6645;
assign w6653 = w6643 & w6652;
assign w6654 = w6650 & w6651;
assign w6655 = w6653 & w6654;
assign w6656 = w6641 & w6655;
assign w6657 = ~w251 & ~w468;
assign w6658 = ~w714 & w6657;
assign w6659 = w2548 & w6658;
assign w6660 = w712 & w2046;
assign w6661 = w5591 & w6660;
assign w6662 = w3505 & w6659;
assign w6663 = w6631 & w6634;
assign w6664 = w6662 & w6663;
assign w6665 = w2660 & w6661;
assign w6666 = w6664 & w6665;
assign w6667 = w2358 & w6666;
assign w6668 = w6656 & w6667;
assign w6669 = w6630 & ~w6668;
assign w6670 = ~w6630 & w6668;
assign w6671 = w2677 & ~w6595;
assign w6672 = ~w2547 & ~w2678;
assign w6673 = ~w6671 & w6672;
assign w6674 = w6671 & ~w6672;
assign w6675 = ~w6673 & ~w6674;
assign w6676 = w1327 & ~w2677;
assign w6677 = w668 & ~w2546;
assign w6678 = (w1399 & ~w2479) | (w1399 & w33348) | (~w2479 & w33348);
assign w6679 = ~w6676 & ~w6677;
assign w6680 = ~w6678 & w6679;
assign w6681 = (w6680 & ~w6675) | (w6680 & w31585) | (~w6675 & w31585);
assign w6682 = ~w6670 & ~w6681;
assign w6683 = ~w6669 & ~w6682;
assign w6684 = w6594 & ~w6683;
assign w6685 = w1101 & w3065;
assign w6686 = ~w315 & ~w432;
assign w6687 = w669 & w6686;
assign w6688 = w2372 & w3478;
assign w6689 = w4312 & w6688;
assign w6690 = w6685 & w6687;
assign w6691 = w6689 & w6690;
assign w6692 = ~w16 & w1765;
assign w6693 = ~w127 & ~w136;
assign w6694 = ~w218 & w6693;
assign w6695 = w549 & w6694;
assign w6696 = ~w163 & ~w418;
assign w6697 = ~w391 & ~w403;
assign w6698 = w2336 & w6697;
assign w6699 = w2784 & w3308;
assign w6700 = w6696 & w6699;
assign w6701 = w1420 & w6698;
assign w6702 = w3168 & w3501;
assign w6703 = w6692 & w6702;
assign w6704 = w6700 & w6701;
assign w6705 = w5495 & w6695;
assign w6706 = w6704 & w6705;
assign w6707 = w6703 & w6706;
assign w6708 = ~w349 & w5613;
assign w6709 = w2887 & w6708;
assign w6710 = ~w264 & ~w283;
assign w6711 = w959 & w6710;
assign w6712 = w1543 & w2247;
assign w6713 = w4521 & w6712;
assign w6714 = w6711 & w6713;
assign w6715 = w6709 & w6714;
assign w6716 = w1417 & w2880;
assign w6717 = w6691 & w6716;
assign w6718 = w6715 & w6717;
assign w6719 = w5543 & w6707;
assign w6720 = w6718 & w6719;
assign w6721 = w668 & ~w2835;
assign w6722 = w1399 & ~w2546;
assign w6723 = (w1327 & ~w2766) | (w1327 & w33349) | (~w2766 & w33349);
assign w6724 = ~w6721 & ~w6722;
assign w6725 = (~w6720 & ~w6724) | (~w6720 & w33350) | (~w6724 & w33350);
assign w6726 = w2680 & w2838;
assign w6727 = ~w2836 & w2923;
assign w6728 = ~w6726 & w6727;
assign w6729 = ~w2680 & w6552;
assign w6730 = w2546 & w2836;
assign w6731 = ~w2921 & ~w6730;
assign w6732 = ~w6729 & ~w6731;
assign w6733 = ~w6728 & ~w6732;
assign w6734 = w1478 & ~w6720;
assign w6735 = (~w6725 & ~w6733) | (~w6725 & w31586) | (~w6733 & w31586);
assign w6736 = ~w6592 & w6735;
assign w6737 = ~w6684 & w6736;
assign w6738 = w1478 & w6733;
assign w6739 = w6724 & w33351;
assign w6740 = ~w6738 & w6739;
assign w6741 = w477 & ~w789;
assign w6742 = ~w164 & ~w287;
assign w6743 = ~w396 & ~w622;
assign w6744 = ~w391 & w752;
assign w6745 = w1028 & w3456;
assign w6746 = w5492 & w6742;
assign w6747 = w6743 & w6746;
assign w6748 = w6744 & w6745;
assign w6749 = w2496 & w5372;
assign w6750 = w6611 & w6749;
assign w6751 = w6747 & w6748;
assign w6752 = w4741 & w6751;
assign w6753 = w6750 & w6752;
assign w6754 = ~w60 & ~w71;
assign w6755 = ~w149 & ~w393;
assign w6756 = w6754 & w6755;
assign w6757 = w1374 & w6756;
assign w6758 = w738 & w777;
assign w6759 = w1098 & w1464;
assign w6760 = w1813 & w1820;
assign w6761 = w2552 & w2943;
assign w6762 = w3369 & w3428;
assign w6763 = w6761 & w6762;
assign w6764 = w6759 & w6760;
assign w6765 = w348 & w6758;
assign w6766 = w629 & w6741;
assign w6767 = w6765 & w6766;
assign w6768 = w6763 & w6764;
assign w6769 = w6757 & w6768;
assign w6770 = w5418 & w6767;
assign w6771 = w6769 & w6770;
assign w6772 = w1657 & w6771;
assign w6773 = w6753 & w6772;
assign w6774 = w668 & ~w2917;
assign w6775 = (w1399 & ~w2766) | (w1399 & w33352) | (~w2766 & w33352);
assign w6776 = w1327 & ~w2835;
assign w6777 = ~w2918 & ~w3053;
assign w6778 = w2923 & ~w6777;
assign w6779 = ~w6726 & w6778;
assign w6780 = w2838 & w6777;
assign w6781 = w2680 & w6780;
assign w6782 = ~w2923 & w6777;
assign w6783 = ~w6781 & ~w6782;
assign w6784 = ~w6779 & w6783;
assign w6785 = ~w6774 & ~w6775;
assign w6786 = ~w6776 & w6785;
assign w6787 = (~w6784 & w33353) | (~w6784 & w33354) | (w33353 & w33354);
assign w6788 = (w6784 & w33355) | (w6784 & w33356) | (w33355 & w33356);
assign w6789 = ~w6787 & ~w6788;
assign w6790 = ~w6737 & w33357;
assign w6791 = (~w6547 & w33358) | (~w6547 & w33359) | (w33358 & w33359);
assign w6792 = ~w6787 & ~w6791;
assign w6793 = (~w6194 & w33360) | (~w6194 & w33361) | (w33360 & w33361);
assign w6794 = ~w6200 & ~w6793;
assign w6795 = (~w6790 & w33362) | (~w6790 & w33363) | (w33362 & w33363);
assign w6796 = (w6790 & w33364) | (w6790 & w33365) | (w33364 & w33365);
assign w6797 = ~w3268 & w4446;
assign w6798 = ~w3139 & w3957;
assign w6799 = ~w3196 & w4068;
assign w6800 = w6222 & w33366;
assign w6801 = ~w6797 & ~w6798;
assign w6802 = ~w6799 & w6801;
assign w6803 = (a_29 & w6800) | (a_29 & w33367) | (w6800 & w33367);
assign w6804 = ~w6800 & w33368;
assign w6805 = ~w6803 & ~w6804;
assign w6806 = ~w6796 & ~w6805;
assign w6807 = ~w6806 & w33369;
assign w6808 = ~w6481 & w6494;
assign w6809 = ~w6495 & ~w6808;
assign w6810 = (w6809 & w6807) | (w6809 & w33370) | (w6807 & w33370);
assign w6811 = ~w6211 & w6226;
assign w6812 = ~w6227 & ~w6811;
assign w6813 = (w6812 & w6810) | (w6812 & w33371) | (w6810 & w33371);
assign w6814 = ~w3475 & w4068;
assign w6815 = ~w3403 & w4446;
assign w6816 = ~w3326 & w3957;
assign w6817 = ~w6814 & ~w6815;
assign w6818 = ~w6816 & w6817;
assign w6819 = (w6818 & ~w5923) | (w6818 & w33372) | (~w5923 & w33372);
assign w6820 = a_29 & ~w6819;
assign w6821 = (~w5923 & w33373) | (~w5923 & w33374) | (w33373 & w33374);
assign w6822 = ~w6820 & ~w6821;
assign w6823 = ~w6810 & w33375;
assign w6824 = ~w6813 & ~w6823;
assign w6825 = w6822 & w6824;
assign w6826 = (~w6813 & ~w6824) | (~w6813 & w33376) | (~w6824 & w33376);
assign w6827 = ~w6479 & w6826;
assign w6828 = ~w518 & ~w2306;
assign w6829 = ~w3615 & w4666;
assign w6830 = ~w2393 & w4638;
assign w6831 = ~w6828 & ~w6829;
assign w6832 = ~w6830 & w6831;
assign w6833 = (w6832 & ~w5463) | (w6832 & w33377) | (~w5463 & w33377);
assign w6834 = a_26 & ~w6833;
assign w6835 = (~w5463 & w33378) | (~w5463 & w33379) | (w33378 & w33379);
assign w6836 = ~w6834 & ~w6835;
assign w6837 = w6479 & ~w6826;
assign w6838 = ~w6827 & ~w6837;
assign w6839 = ~w6836 & w6838;
assign w6840 = (~w6827 & ~w6838) | (~w6827 & w33380) | (~w6838 & w33380);
assign w6841 = ~w6477 & ~w6840;
assign w6842 = (w5286 & ~w3712) | (w5286 & w33381) | (~w3712 & w33381);
assign w6843 = ~w2148 & w5016;
assign w6844 = (w5080 & ~w2235) | (w5080 & w33382) | (~w2235 & w33382);
assign w6845 = w5017 & w5103;
assign w6846 = ~w6843 & w33383;
assign w6847 = (a_23 & w6845) | (a_23 & w33384) | (w6845 & w33384);
assign w6848 = ~w6845 & w33385;
assign w6849 = ~w6847 & ~w6848;
assign w6850 = w6477 & w6840;
assign w6851 = ~w6841 & ~w6850;
assign w6852 = ~w6849 & w6851;
assign w6853 = (~w6841 & ~w6851) | (~w6841 & w33386) | (~w6851 & w33386);
assign w6854 = ~w6465 & w6474;
assign w6855 = ~w6475 & ~w6854;
assign w6856 = w6853 & w6855;
assign w6857 = ~w6475 & ~w6856;
assign w6858 = ~w6463 & ~w6857;
assign w6859 = (w5308 & ~w1913) | (w5308 & w33387) | (~w1913 & w33387);
assign w6860 = (w5816 & ~w1807) | (w5816 & w33388) | (~w1807 & w33388);
assign w6861 = (w5818 & ~w1714) | (w5818 & w33276) | (~w1714 & w33276);
assign w6862 = ~w6859 & ~w6860;
assign w6863 = ~w6861 & w6862;
assign w6864 = (w6863 & w4428) | (w6863 & w33389) | (w4428 & w33389);
assign w6865 = a_20 & ~w6864;
assign w6866 = (w4428 & w33390) | (w4428 & w33391) | (w33390 & w33391);
assign w6867 = ~w6865 & ~w6866;
assign w6868 = w6463 & w6857;
assign w6869 = ~w6858 & ~w6868;
assign w6870 = w6867 & w6869;
assign w6871 = (~w6858 & ~w6869) | (~w6858 & w33392) | (~w6869 & w33392);
assign w6872 = ~w6411 & ~w6413;
assign w6873 = ~w6414 & ~w6872;
assign w6874 = ~w6871 & w6873;
assign w6875 = w6871 & ~w6873;
assign w6876 = ~w6874 & ~w6875;
assign w6877 = ~w1475 & w6304;
assign w6878 = (w6059 & ~w1628) | (w6059 & w33393) | (~w1628 & w33393);
assign w6879 = (w6061 & ~w643) | (w6061 & w33394) | (~w643 & w33394);
assign w6880 = ~w6878 & ~w6879;
assign w6881 = ~w6877 & w6880;
assign w6882 = (w6881 & ~w4041) | (w6881 & w33395) | (~w4041 & w33395);
assign w6883 = a_17 & w6882;
assign w6884 = (w4041 & w33396) | (w4041 & w33397) | (w33396 & w33397);
assign w6885 = ~w6883 & ~w6884;
assign w6886 = w6876 & ~w6885;
assign w6887 = ~w6876 & w6885;
assign w6888 = ~w6886 & ~w6887;
assign w6889 = ~w6853 & ~w6855;
assign w6890 = ~w6856 & ~w6889;
assign w6891 = (w5818 & ~w1913) | (w5818 & w33398) | (~w1913 & w33398);
assign w6892 = (w5308 & ~w2005) | (w5308 & w33399) | (~w2005 & w33399);
assign w6893 = (w5816 & ~w1714) | (w5816 & w33294) | (~w1714 & w33294);
assign w6894 = ~w6891 & ~w6892;
assign w6895 = ~w6893 & w6894;
assign w6896 = (w6895 & ~w4592) | (w6895 & w33400) | (~w4592 & w33400);
assign w6897 = a_20 & ~w6896;
assign w6898 = (~w4592 & w33401) | (~w4592 & w33402) | (w33401 & w33402);
assign w6899 = ~w6897 & ~w6898;
assign w6900 = w6890 & w6899;
assign w6901 = w6836 & ~w6838;
assign w6902 = ~w6839 & ~w6901;
assign w6903 = ~w2306 & w4638;
assign w6904 = ~w2393 & w4666;
assign w6905 = (~w518 & ~w3538) | (~w518 & w33403) | (~w3538 & w33403);
assign w6906 = ~w6903 & ~w6904;
assign w6907 = ~w6905 & w6906;
assign w6908 = (w6907 & ~w5483) | (w6907 & w33404) | (~w5483 & w33404);
assign w6909 = a_26 & ~w6908;
assign w6910 = (~w5483 & w33405) | (~w5483 & w33406) | (w33405 & w33406);
assign w6911 = ~w6909 & ~w6910;
assign w6912 = ~w6822 & ~w6824;
assign w6913 = ~w6825 & ~w6912;
assign w6914 = ~w6911 & ~w6913;
assign w6915 = w6911 & w6913;
assign w6916 = ~w6807 & w33407;
assign w6917 = ~w6810 & ~w6916;
assign w6918 = ~w3326 & w4068;
assign w6919 = (w3957 & ~w3267) | (w3957 & w33408) | (~w3267 & w33408);
assign w6920 = ~w3475 & w4446;
assign w6921 = ~w6918 & ~w6919;
assign w6922 = ~w6920 & w6921;
assign w6923 = (w6922 & ~w6108) | (w6922 & w33409) | (~w6108 & w33409);
assign w6924 = a_29 & ~w6923;
assign w6925 = (~w6108 & w33410) | (~w6108 & w33411) | (w33410 & w33411);
assign w6926 = ~w6924 & ~w6925;
assign w6927 = ~w6917 & ~w6926;
assign w6928 = ~w518 & ~w3403;
assign w6929 = ~w2306 & w4666;
assign w6930 = (w4638 & ~w3538) | (w4638 & w33412) | (~w3538 & w33412);
assign w6931 = ~w6929 & ~w6930;
assign w6932 = ~w6928 & w6931;
assign w6933 = (w6932 & ~w5706) | (w6932 & w33413) | (~w5706 & w33413);
assign w6934 = a_26 & ~w6933;
assign w6935 = (~w5706 & w33414) | (~w5706 & w33415) | (w33414 & w33415);
assign w6936 = ~w6934 & ~w6935;
assign w6937 = w6917 & w6926;
assign w6938 = ~w6927 & ~w6937;
assign w6939 = ~w6936 & w6938;
assign w6940 = (~w6927 & ~w6938) | (~w6927 & w33416) | (~w6938 & w33416);
assign w6941 = ~w6915 & ~w6940;
assign w6942 = ~w6914 & ~w6941;
assign w6943 = w6902 & ~w6942;
assign w6944 = ~w2075 & w5016;
assign w6945 = (w5286 & ~w2235) | (w5286 & w33417) | (~w2235 & w33417);
assign w6946 = ~w2148 & w5080;
assign w6947 = ~w6945 & ~w6946;
assign w6948 = ~w6944 & w6947;
assign w6949 = (w6948 & ~w4962) | (w6948 & w33418) | (~w4962 & w33418);
assign w6950 = a_23 & ~w6949;
assign w6951 = (~w4962 & w33419) | (~w4962 & w33420) | (w33419 & w33420);
assign w6952 = ~w6950 & ~w6951;
assign w6953 = ~w6902 & w6942;
assign w6954 = ~w6943 & ~w6953;
assign w6955 = ~w6952 & w6954;
assign w6956 = (~w6943 & ~w6954) | (~w6943 & w33421) | (~w6954 & w33421);
assign w6957 = w6849 & ~w6851;
assign w6958 = ~w6852 & ~w6957;
assign w6959 = w6956 & ~w6958;
assign w6960 = (w5308 & ~w3658) | (w5308 & w33422) | (~w3658 & w33422);
assign w6961 = (w5818 & ~w2005) | (w5818 & w33423) | (~w2005 & w33423);
assign w6962 = (w5816 & ~w1913) | (w5816 & w33424) | (~w1913 & w33424);
assign w6963 = ~w6961 & ~w6962;
assign w6964 = ~w6960 & w6963;
assign w6965 = (w6964 & w4578) | (w6964 & w33425) | (w4578 & w33425);
assign w6966 = a_20 & ~w6965;
assign w6967 = (w4578 & w33426) | (w4578 & w33427) | (w33426 & w33427);
assign w6968 = ~w6966 & ~w6967;
assign w6969 = ~w6956 & w6958;
assign w6970 = ~w6959 & ~w6969;
assign w6971 = w6968 & w6970;
assign w6972 = (~w6959 & ~w6970) | (~w6959 & w33428) | (~w6970 & w33428);
assign w6973 = ~w6890 & ~w6899;
assign w6974 = ~w6900 & ~w6973;
assign w6975 = ~w6972 & w6974;
assign w6976 = ~w6900 & ~w6975;
assign w6977 = ~w6867 & ~w6869;
assign w6978 = ~w6870 & ~w6977;
assign w6979 = w6976 & ~w6978;
assign w6980 = ~w6976 & w6978;
assign w6981 = ~w6979 & ~w6980;
assign w6982 = ~w3813 & w6059;
assign w6983 = (w6304 & ~w643) | (w6304 & w33429) | (~w643 & w33429);
assign w6984 = (w6061 & ~w1628) | (w6061 & w33430) | (~w1628 & w33430);
assign w6985 = w4224 & w6063;
assign w6986 = ~w6982 & w33431;
assign w6987 = ~w6985 & w33432;
assign w6988 = (~a_17 & w6985) | (~a_17 & w33433) | (w6985 & w33433);
assign w6989 = ~w6987 & ~w6988;
assign w6990 = w6981 & w6989;
assign w6991 = (~w6979 & ~w6981) | (~w6979 & w33434) | (~w6981 & w33434);
assign w6992 = w6888 & w6991;
assign w6993 = ~w6888 & ~w6991;
assign w6994 = ~w6992 & ~w6993;
assign w6995 = ~w1397 & w6446;
assign w6996 = w6438 & w6441;
assign w6997 = (w6996 & ~w3904) | (w6996 & w33435) | (~w3904 & w33435);
assign w6998 = ~w6441 & w6444;
assign w6999 = (w6998 & ~w1308) | (w6998 & w33436) | (~w1308 & w33436);
assign w7000 = ~w6995 & ~w6999;
assign w7001 = ~w6997 & w7000;
assign w7002 = (w7001 & ~w3964) | (w7001 & w33437) | (~w3964 & w33437);
assign w7003 = a_14 & ~w7002;
assign w7004 = (~w3964 & w33438) | (~w3964 & w33439) | (w33438 & w33439);
assign w7005 = ~w7003 & ~w7004;
assign w7006 = w6994 & w7005;
assign w7007 = (~w6992 & ~w6994) | (~w6992 & w33440) | (~w6994 & w33440);
assign w7008 = (w6998 & ~w3904) | (w6998 & w33441) | (~w3904 & w33441);
assign w7009 = ~w3958 & w6996;
assign w7010 = (w6446 & ~w1308) | (w6446 & w33442) | (~w1308 & w33442);
assign w7011 = ~w7009 & ~w7010;
assign w7012 = ~w7008 & w7011;
assign w7013 = (w7012 & ~w3943) | (w7012 & w33443) | (~w3943 & w33443);
assign w7014 = a_14 & ~w7013;
assign w7015 = (~w3943 & w33444) | (~w3943 & w33445) | (w33444 & w33445);
assign w7016 = ~w7014 & ~w7015;
assign w7017 = ~w7007 & w7016;
assign w7018 = (~w6874 & ~w6876) | (~w6874 & w33446) | (~w6876 & w33446);
assign w7019 = w6415 & ~w6417;
assign w7020 = ~w6418 & ~w7019;
assign w7021 = ~w1397 & w6304;
assign w7022 = ~w1475 & w6061;
assign w7023 = (w6059 & ~w643) | (w6059 & w33447) | (~w643 & w33447);
assign w7024 = ~w7021 & ~w7023;
assign w7025 = ~w7022 & w7024;
assign w7026 = (w7025 & ~w4056) | (w7025 & w33448) | (~w4056 & w33448);
assign w7027 = a_17 & w7026;
assign w7028 = (w4056 & w33449) | (w4056 & w33450) | (w33449 & w33450);
assign w7029 = ~w7027 & ~w7028;
assign w7030 = w7020 & ~w7029;
assign w7031 = ~w7020 & w7029;
assign w7032 = ~w7030 & ~w7031;
assign w7033 = ~w7018 & w7032;
assign w7034 = w7018 & ~w7032;
assign w7035 = ~w7033 & ~w7034;
assign w7036 = w7007 & ~w7016;
assign w7037 = ~w7017 & ~w7036;
assign w7038 = w7035 & w7037;
assign w7039 = (~w7017 & ~w7037) | (~w7017 & w33451) | (~w7037 & w33451);
assign w7040 = ~w6424 & w6433;
assign w7041 = ~w6434 & ~w7040;
assign w7042 = (~w7030 & ~w7032) | (~w7030 & w33452) | (~w7032 & w33452);
assign w7043 = (w6446 & ~w3904) | (w6446 & w33453) | (~w3904 & w33453);
assign w7044 = ~w3958 & w6998;
assign w7045 = ~w7043 & ~w7044;
assign w7046 = (w7045 & ~w4073) | (w7045 & w33454) | (~w4073 & w33454);
assign w7047 = a_14 & ~w7046;
assign w7048 = (~w4073 & w33455) | (~w4073 & w33456) | (w33455 & w33456);
assign w7049 = ~w7047 & ~w7048;
assign w7050 = ~w7042 & w7049;
assign w7051 = w7042 & ~w7049;
assign w7052 = ~w7050 & ~w7051;
assign w7053 = ~w7041 & w7052;
assign w7054 = w7041 & ~w7052;
assign w7055 = ~w7053 & ~w7054;
assign w7056 = w7039 & ~w7055;
assign w7057 = ~w7039 & w7055;
assign w7058 = ~w7056 & ~w7057;
assign w7059 = ~w6981 & ~w6989;
assign w7060 = ~w6990 & ~w7059;
assign w7061 = w6972 & ~w6974;
assign w7062 = ~w6975 & ~w7061;
assign w7063 = (w6059 & ~w1807) | (w6059 & w33457) | (~w1807 & w33457);
assign w7064 = (w6304 & ~w1628) | (w6304 & w33458) | (~w1628 & w33458);
assign w7065 = ~w3813 & w6061;
assign w7066 = ~w7063 & ~w7064;
assign w7067 = ~w7065 & w7066;
assign w7068 = (w7067 & ~w4244) | (w7067 & w33459) | (~w4244 & w33459);
assign w7069 = a_17 & ~w7068;
assign w7070 = (~w4244 & w33460) | (~w4244 & w33461) | (w33460 & w33461);
assign w7071 = ~w7069 & ~w7070;
assign w7072 = w7062 & w7071;
assign w7073 = (~w6511 & w6806) | (~w6511 & w33462) | (w6806 & w33462);
assign w7074 = ~w6807 & ~w7073;
assign w7075 = ~w3326 & w4446;
assign w7076 = ~w3196 & w3957;
assign w7077 = (w4068 & ~w3267) | (w4068 & w33463) | (~w3267 & w33463);
assign w7078 = ~w7076 & ~w7077;
assign w7079 = ~w7075 & w7078;
assign w7080 = (w7079 & w5903) | (w7079 & w33464) | (w5903 & w33464);
assign w7081 = a_29 & w7080;
assign w7082 = (~w5903 & w33465) | (~w5903 & w33466) | (w33465 & w33466);
assign w7083 = ~w7081 & ~w7082;
assign w7084 = w7074 & ~w7083;
assign w7085 = ~w7074 & w7083;
assign w7086 = ~w7084 & ~w7085;
assign w7087 = ~w3403 & w4638;
assign w7088 = (w4666 & ~w3538) | (w4666 & w33467) | (~w3538 & w33467);
assign w7089 = ~w518 & ~w3475;
assign w7090 = ~w7087 & ~w7088;
assign w7091 = ~w7089 & w7090;
assign w7092 = (w7091 & ~w5652) | (w7091 & w33468) | (~w5652 & w33468);
assign w7093 = a_26 & w7092;
assign w7094 = (w5652 & w33469) | (w5652 & w33470) | (w33469 & w33470);
assign w7095 = ~w7093 & ~w7094;
assign w7096 = w7086 & ~w7095;
assign w7097 = (~w7084 & ~w7086) | (~w7084 & w33471) | (~w7086 & w33471);
assign w7098 = ~w2075 & w5286;
assign w7099 = ~w2393 & w5016;
assign w7100 = ~w3615 & w5080;
assign w7101 = ~w7099 & ~w7100;
assign w7102 = ~w7098 & w7101;
assign w7103 = (w7102 & ~w5227) | (w7102 & w33472) | (~w5227 & w33472);
assign w7104 = a_23 & w7103;
assign w7105 = (w5227 & w33473) | (w5227 & w33474) | (w33473 & w33474);
assign w7106 = ~w7104 & ~w7105;
assign w7107 = ~w7097 & ~w7106;
assign w7108 = w6936 & ~w6938;
assign w7109 = ~w6939 & ~w7108;
assign w7110 = w7097 & w7106;
assign w7111 = ~w7107 & ~w7110;
assign w7112 = ~w7109 & w7111;
assign w7113 = ~w7107 & ~w7112;
assign w7114 = ~w6914 & ~w6915;
assign w7115 = ~w2075 & w5080;
assign w7116 = ~w2148 & w5286;
assign w7117 = ~w3615 & w5016;
assign w7118 = ~w7116 & ~w7117;
assign w7119 = ~w7115 & w7118;
assign w7120 = (w7119 & ~w5242) | (w7119 & w33475) | (~w5242 & w33475);
assign w7121 = a_23 & ~w7120;
assign w7122 = (~w5242 & w33476) | (~w5242 & w33477) | (w33476 & w33477);
assign w7123 = ~w7121 & ~w7122;
assign w7124 = w6940 & ~w7123;
assign w7125 = ~w6940 & w7123;
assign w7126 = ~w7124 & ~w7125;
assign w7127 = w7114 & w7126;
assign w7128 = ~w7114 & ~w7126;
assign w7129 = ~w7127 & ~w7128;
assign w7130 = w7113 & ~w7129;
assign w7131 = ~w7123 & w7129;
assign w7132 = ~w7130 & ~w7131;
assign w7133 = (w5818 & ~w3658) | (w5818 & w33478) | (~w3658 & w33478);
assign w7134 = (w5816 & ~w2005) | (w5816 & w33479) | (~w2005 & w33479);
assign w7135 = (w5308 & ~w3712) | (w5308 & w33480) | (~w3712 & w33480);
assign w7136 = (w5309 & w4790) | (w5309 & w33481) | (w4790 & w33481);
assign w7137 = ~w7134 & ~w7135;
assign w7138 = ~w7133 & w7137;
assign w7139 = (a_20 & w7136) | (a_20 & w33482) | (w7136 & w33482);
assign w7140 = ~w7136 & w33483;
assign w7141 = ~w7139 & ~w7140;
assign w7142 = w7132 & w7141;
assign w7143 = w6952 & ~w6954;
assign w7144 = ~w6955 & ~w7143;
assign w7145 = ~w7132 & ~w7141;
assign w7146 = ~w7142 & ~w7145;
assign w7147 = ~w7144 & w7146;
assign w7148 = (~w7142 & ~w7146) | (~w7142 & w33484) | (~w7146 & w33484);
assign w7149 = ~w3813 & w6304;
assign w7150 = (w6061 & ~w1807) | (w6061 & w33485) | (~w1807 & w33485);
assign w7151 = (w6059 & ~w1714) | (w6059 & w33393) | (~w1714 & w33393);
assign w7152 = w4508 & w6063;
assign w7153 = ~w7149 & w33486;
assign w7154 = (a_17 & w7152) | (a_17 & w33487) | (w7152 & w33487);
assign w7155 = ~w7152 & w33488;
assign w7156 = ~w7154 & ~w7155;
assign w7157 = ~w7148 & w7156;
assign w7158 = ~w6968 & ~w6970;
assign w7159 = ~w6971 & ~w7158;
assign w7160 = w7148 & ~w7156;
assign w7161 = ~w7157 & ~w7160;
assign w7162 = w7159 & w7161;
assign w7163 = (~w7157 & ~w7161) | (~w7157 & w33489) | (~w7161 & w33489);
assign w7164 = ~w7062 & ~w7071;
assign w7165 = ~w7072 & ~w7164;
assign w7166 = ~w7163 & w7165;
assign w7167 = (~w7072 & ~w7165) | (~w7072 & w33490) | (~w7165 & w33490);
assign w7168 = ~w7060 & ~w7167;
assign w7169 = ~w1397 & w6998;
assign w7170 = ~w1475 & w6446;
assign w7171 = (w6996 & ~w1308) | (w6996 & w33491) | (~w1308 & w33491);
assign w7172 = ~w7169 & ~w7170;
assign w7173 = ~w7171 & w7172;
assign w7174 = (w7173 & ~w3834) | (w7173 & w33492) | (~w3834 & w33492);
assign w7175 = a_14 & ~w7174;
assign w7176 = (~w3834 & w33493) | (~w3834 & w33494) | (w33493 & w33494);
assign w7177 = ~w7175 & ~w7176;
assign w7178 = w7060 & w7167;
assign w7179 = ~w7168 & ~w7178;
assign w7180 = w7177 & w7179;
assign w7181 = (~w7168 & ~w7179) | (~w7168 & w33495) | (~w7179 & w33495);
assign w7182 = ~a_10 & a_11;
assign w7183 = a_10 & ~a_11;
assign w7184 = ~w7182 & ~w7183;
assign w7185 = ~a_8 & ~a_9;
assign w7186 = a_8 & a_9;
assign w7187 = ~w7185 & ~w7186;
assign w7188 = ~a_9 & ~a_10;
assign w7189 = a_9 & a_10;
assign w7190 = ~w7188 & ~w7189;
assign w7191 = ~w7187 & ~w7190;
assign w7192 = ~w7184 & w7191;
assign w7193 = ~w7184 & w7187;
assign w7194 = (~w3828 & w33498) | (~w3828 & w33499) | (w33498 & w33499);
assign w7195 = ~w7194 & w33500;
assign w7196 = (a_11 & w7194) | (a_11 & w33501) | (w7194 & w33501);
assign w7197 = ~w7195 & ~w7196;
assign w7198 = ~w7181 & ~w7197;
assign w7199 = ~w6994 & ~w7005;
assign w7200 = ~w7006 & ~w7199;
assign w7201 = w7181 & w7197;
assign w7202 = ~w7198 & ~w7201;
assign w7203 = w7200 & w7202;
assign w7204 = (~w7198 & ~w7202) | (~w7198 & w33502) | (~w7202 & w33502);
assign w7205 = ~w7035 & ~w7037;
assign w7206 = ~w7038 & ~w7205;
assign w7207 = ~w7204 & w7206;
assign w7208 = w7163 & ~w7165;
assign w7209 = ~w7166 & ~w7208;
assign w7210 = ~w1397 & w6996;
assign w7211 = ~w1475 & w6998;
assign w7212 = (w6446 & ~w643) | (w6446 & w33503) | (~w643 & w33503);
assign w7213 = ~w7210 & ~w7212;
assign w7214 = ~w7211 & w7213;
assign w7215 = (w7214 & ~w4056) | (w7214 & w33504) | (~w4056 & w33504);
assign w7216 = a_14 & ~w7215;
assign w7217 = (~w4056 & w33505) | (~w4056 & w33506) | (w33505 & w33506);
assign w7218 = ~w7216 & ~w7217;
assign w7219 = w7209 & w7218;
assign w7220 = (w5816 & ~w3658) | (w5816 & w33507) | (~w3658 & w33507);
assign w7221 = (w5308 & ~w2235) | (w5308 & w33508) | (~w2235 & w33508);
assign w7222 = (w5818 & ~w3712) | (w5818 & w33509) | (~w3712 & w33509);
assign w7223 = ~w7221 & ~w7222;
assign w7224 = ~w7220 & w7223;
assign w7225 = (w7224 & ~w4810) | (w7224 & w33510) | (~w4810 & w33510);
assign w7226 = a_20 & w7225;
assign w7227 = (w4810 & w33511) | (w4810 & w33512) | (w33511 & w33512);
assign w7228 = ~w7226 & ~w7227;
assign w7229 = (w5818 & ~w2235) | (w5818 & w33513) | (~w2235 & w33513);
assign w7230 = ~w2148 & w5308;
assign w7231 = (w5816 & ~w3712) | (w5816 & w33514) | (~w3712 & w33514);
assign w7232 = w5103 & w5309;
assign w7233 = ~w7230 & w33515;
assign w7234 = (a_20 & w7232) | (a_20 & w33516) | (w7232 & w33516);
assign w7235 = ~w7232 & w33517;
assign w7236 = ~w7234 & ~w7235;
assign w7237 = ~w7086 & w7095;
assign w7238 = ~w7096 & ~w7237;
assign w7239 = ~w3403 & w4666;
assign w7240 = ~w3475 & w4638;
assign w7241 = ~w518 & ~w3326;
assign w7242 = ~w7239 & ~w7240;
assign w7243 = ~w7241 & w7242;
assign w7244 = (w7243 & ~w5923) | (w7243 & w33518) | (~w5923 & w33518);
assign w7245 = ~a_26 & w7244;
assign w7246 = (w5923 & w33519) | (w5923 & w33520) | (w33519 & w33520);
assign w7247 = ~w7245 & ~w7246;
assign w7248 = ~w6795 & ~w6796;
assign w7249 = w6805 & w7247;
assign w7250 = ~w6805 & ~w7247;
assign w7251 = ~w7249 & ~w7250;
assign w7252 = w7248 & w7251;
assign w7253 = ~w7248 & ~w7251;
assign w7254 = ~w7252 & ~w7253;
assign w7255 = w7247 & ~w7254;
assign w7256 = (~w6789 & w6737) | (~w6789 & w33521) | (w6737 & w33521);
assign w7257 = ~w6790 & ~w7256;
assign w7258 = ~w3007 & w3957;
assign w7259 = ~w3139 & w4446;
assign w7260 = ~w3049 & w4068;
assign w7261 = ~w7258 & ~w7259;
assign w7262 = ~w7260 & w7261;
assign w7263 = (w7262 & w6505) | (w7262 & w33522) | (w6505 & w33522);
assign w7264 = ~a_29 & w7263;
assign w7265 = (~w6505 & w33523) | (~w6505 & w33524) | (w33523 & w33524);
assign w7266 = ~w7264 & ~w7265;
assign w7267 = w7257 & w7266;
assign w7268 = w3949 & w3954;
assign w7269 = ~a_29 & ~w4070;
assign w7270 = ~w2917 & w4446;
assign w7271 = (w3957 & ~w2766) | (w3957 & w33525) | (~w2766 & w33525);
assign w7272 = ~w2835 & w4068;
assign w7273 = ~w7270 & ~w7271;
assign w7274 = w7273 & w33526;
assign w7275 = (a_29 & ~w7273) | (a_29 & w33527) | (~w7273 & w33527);
assign w7276 = w7273 & w33528;
assign w7277 = w6784 & w7276;
assign w7278 = ~w7274 & ~w7275;
assign w7279 = (w7278 & w6784) | (w7278 & w31587) | (w6784 & w31587);
assign w7280 = ~w7277 & w7279;
assign w7281 = ~w6669 & ~w6670;
assign w7282 = ~w6681 & w7281;
assign w7283 = w6681 & ~w7281;
assign w7284 = ~w7282 & ~w7283;
assign w7285 = ~w7280 & ~w7284;
assign w7286 = w2480 & ~w2601;
assign w7287 = ~w6595 & ~w7286;
assign w7288 = w1478 & ~w7287;
assign w7289 = (w668 & ~w2479) | (w668 & w33529) | (~w2479 & w33529);
assign w7290 = (w1327 & ~w2600) | (w1327 & w33530) | (~w2600 & w33530);
assign w7291 = ~w7289 & ~w7290;
assign w7292 = (w7291 & w7287) | (w7291 & w33531) | (w7287 & w33531);
assign w7293 = w2680 & w31588;
assign w7294 = w4070 & ~w6552;
assign w7295 = ~w2680 & w7294;
assign w7296 = ~w2546 & w4068;
assign w7297 = (w4446 & ~w2766) | (w4446 & w33532) | (~w2766 & w33532);
assign w7298 = ~w2677 & w3957;
assign w7299 = ~w7296 & ~w7297;
assign w7300 = ~w7298 & w7299;
assign w7301 = ~w7295 & w7300;
assign w7302 = ~w7293 & w7301;
assign w7303 = (a_29 & w7288) | (a_29 & w31589) | (w7288 & w31589);
assign w7304 = ~w7288 & w31590;
assign w7305 = ~w7303 & ~w7304;
assign w7306 = w7302 & w7305;
assign w7307 = ~w7302 & ~w7305;
assign w7308 = ~w7306 & ~w7307;
assign w7309 = ~w7292 & w7308;
assign w7310 = ~w2546 & w4446;
assign w7311 = (w3957 & ~w2479) | (w3957 & w33533) | (~w2479 & w33533);
assign w7312 = ~w2677 & w4068;
assign w7313 = ~w7310 & ~w7311;
assign w7314 = w7313 & w33534;
assign w7315 = (w7314 & ~w6675) | (w7314 & w33535) | (~w6675 & w33535);
assign w7316 = (a_29 & ~w7313) | (a_29 & w33536) | (~w7313 & w33536);
assign w7317 = (~w7316 & ~w6675) | (~w7316 & w37563) | (~w6675 & w37563);
assign w7318 = ~w7315 & w7317;
assign w7319 = (~w1477 & ~w2600) | (~w1477 & w33537) | (~w2600 & w33537);
assign w7320 = w2677 & w4070;
assign w7321 = w6595 & w7320;
assign w7322 = ~w2677 & w4070;
assign w7323 = ~w6595 & w7322;
assign w7324 = (w4068 & ~w2479) | (w4068 & w31591) | (~w2479 & w31591);
assign w7325 = (w3957 & ~w2600) | (w3957 & w31592) | (~w2600 & w31592);
assign w7326 = ~w2677 & w4446;
assign w7327 = ~w7324 & ~w7325;
assign w7328 = ~w7326 & w7327;
assign w7329 = ~w7321 & ~w7323;
assign w7330 = w7328 & w7329;
assign w7331 = w4070 & ~w7287;
assign w7332 = (w4446 & ~w2479) | (w4446 & w31593) | (~w2479 & w31593);
assign w7333 = (w4068 & ~w2600) | (w4068 & w31594) | (~w2600 & w31594);
assign w7334 = ~w7332 & ~w7333;
assign w7335 = (w3954 & ~w2600) | (w3954 & w31595) | (~w2600 & w31595);
assign w7336 = a_29 & ~w7335;
assign w7337 = w7334 & w7336;
assign w7338 = ~w7331 & w7337;
assign w7339 = w7330 & w7338;
assign w7340 = ~w7319 & ~w7339;
assign w7341 = w7318 & ~w7340;
assign w7342 = ~w7308 & w7341;
assign w7343 = ~w7309 & ~w7342;
assign w7344 = w6605 & w33538;
assign w7345 = ~w6630 & ~w7344;
assign w7346 = ~w2835 & w4446;
assign w7347 = (w4068 & ~w2766) | (w4068 & w31596) | (~w2766 & w31596);
assign w7348 = ~w2546 & w3957;
assign w7349 = ~w7346 & ~w7347;
assign w7350 = (a_29 & ~w7349) | (a_29 & w31597) | (~w7349 & w31597);
assign w7351 = w7349 & w33539;
assign w7352 = ~w7350 & ~w7351;
assign w7353 = ~w6733 & w7352;
assign w7354 = w7349 & w33540;
assign w7355 = ~w7268 & ~w7350;
assign w7356 = ~w7354 & w7355;
assign w7357 = w6733 & w7356;
assign w7358 = ~w7353 & ~w7357;
assign w7359 = w7345 & ~w7358;
assign w7360 = ~w7345 & w7358;
assign w7361 = ~w7359 & ~w7360;
assign w7362 = ~w7343 & w7361;
assign w7363 = w7280 & w7284;
assign w7364 = ~w7359 & ~w7363;
assign w7365 = (~w7285 & w7362) | (~w7285 & w31598) | (w7362 & w31598);
assign w7366 = ~w6594 & w6683;
assign w7367 = ~w6684 & ~w7366;
assign w7368 = w4070 & w6545;
assign w7369 = w4070 & ~w6544;
assign w7370 = ~w2920 & w31599;
assign w7371 = ~w2917 & w4068;
assign w7372 = ~w3007 & w4446;
assign w7373 = ~w2835 & w3957;
assign w7374 = ~w7371 & ~w7372;
assign w7375 = ~w7373 & w7374;
assign w7376 = ~w7370 & w7375;
assign w7377 = ~w7368 & w7376;
assign w7378 = ~a_29 & w7377;
assign w7379 = a_29 & ~w7377;
assign w7380 = ~w7378 & ~w7379;
assign w7381 = w7367 & w7380;
assign w7382 = ~w7367 & ~w7380;
assign w7383 = ~w7381 & ~w7382;
assign w7384 = w7365 & w7383;
assign w7385 = ~w3049 & w4446;
assign w7386 = ~w3007 & w4068;
assign w7387 = ~w2917 & w3957;
assign w7388 = ~w7385 & ~w7386;
assign w7389 = ~w7387 & w7388;
assign w7390 = (w6194 & w33541) | (w6194 & w33542) | (w33541 & w33542);
assign w7391 = (~w6194 & w33543) | (~w6194 & w33544) | (w33543 & w33544);
assign w7392 = ~w7390 & ~w7391;
assign w7393 = w6735 & ~w6740;
assign w7394 = ~w6592 & ~w6684;
assign w7395 = ~w7393 & w7394;
assign w7396 = w7393 & ~w7394;
assign w7397 = ~w7395 & ~w7396;
assign w7398 = (~w7381 & ~w7397) | (~w7381 & w33545) | (~w7397 & w33545);
assign w7399 = ~w7384 & w7398;
assign w7400 = ~w7392 & ~w7397;
assign w7401 = ~w7257 & ~w7266;
assign w7402 = ~w7400 & ~w7401;
assign w7403 = (~w7267 & w7399) | (~w7267 & w33546) | (w7399 & w33546);
assign w7404 = ~w6787 & ~w6790;
assign w7405 = ~w6551 & ~w6791;
assign w7406 = ~w3196 & w4446;
assign w7407 = ~w3139 & w4068;
assign w7408 = ~w3049 & w3957;
assign w7409 = ~w7406 & ~w7407;
assign w7410 = (a_29 & ~w7409) | (a_29 & w33547) | (~w7409 & w33547);
assign w7411 = w4070 & w6491;
assign w7412 = w7409 & w33548;
assign w7413 = ~w7411 & w7412;
assign w7414 = (~w7410 & ~w6491) | (~w7410 & w33549) | (~w6491 & w33549);
assign w7415 = ~w7413 & w7414;
assign w7416 = w7405 & w7415;
assign w7417 = w7404 & w7416;
assign w7418 = ~w7405 & w7415;
assign w7419 = ~w7404 & w7418;
assign w7420 = ~w7417 & ~w7419;
assign w7421 = ~w7405 & ~w7415;
assign w7422 = w7404 & w7421;
assign w7423 = w7405 & ~w7415;
assign w7424 = ~w7404 & w7423;
assign w7425 = ~w7422 & ~w7424;
assign w7426 = (w7425 & ~w7403) | (w7425 & w33550) | (~w7403 & w33550);
assign w7427 = w7254 & w7426;
assign w7428 = ~w7255 & ~w7427;
assign w7429 = w7238 & ~w7428;
assign w7430 = ~w7238 & w7428;
assign w7431 = ~w2306 & w5016;
assign w7432 = ~w3615 & w5286;
assign w7433 = ~w2393 & w5080;
assign w7434 = ~w7431 & ~w7432;
assign w7435 = ~w7433 & w7434;
assign w7436 = (w7435 & ~w5463) | (w7435 & w33551) | (~w5463 & w33551);
assign w7437 = a_23 & ~w7436;
assign w7438 = (~w5463 & w33552) | (~w5463 & w33553) | (w33552 & w33553);
assign w7439 = ~w7437 & ~w7438;
assign w7440 = ~w7430 & w7439;
assign w7441 = (w7236 & w7440) | (w7236 & w33554) | (w7440 & w33554);
assign w7442 = ~w7440 & w33555;
assign w7443 = w7109 & ~w7111;
assign w7444 = ~w7112 & ~w7443;
assign w7445 = ~w7442 & w7444;
assign w7446 = (~w7228 & w7445) | (~w7228 & w33556) | (w7445 & w33556);
assign w7447 = ~w7113 & w7129;
assign w7448 = ~w7130 & ~w7447;
assign w7449 = ~w7445 & w33557;
assign w7450 = ~w7446 & ~w7449;
assign w7451 = ~w7448 & w7450;
assign w7452 = (w6059 & ~w1913) | (w6059 & w33558) | (~w1913 & w33558);
assign w7453 = (w6061 & ~w1714) | (w6061 & w33430) | (~w1714 & w33430);
assign w7454 = (w6304 & ~w1807) | (w6304 & w33559) | (~w1807 & w33559);
assign w7455 = ~w7452 & ~w7453;
assign w7456 = ~w7454 & w7455;
assign w7457 = (w7456 & w4428) | (w7456 & w33560) | (w4428 & w33560);
assign w7458 = a_17 & w7457;
assign w7459 = (~w4428 & w33561) | (~w4428 & w33562) | (w33561 & w33562);
assign w7460 = ~w7458 & ~w7459;
assign w7461 = (~w7460 & w7451) | (~w7460 & w33563) | (w7451 & w33563);
assign w7462 = w7144 & ~w7146;
assign w7463 = ~w7147 & ~w7462;
assign w7464 = ~w7451 & w33564;
assign w7465 = ~w7461 & ~w7464;
assign w7466 = w7463 & w7465;
assign w7467 = (~w7461 & ~w7463) | (~w7461 & w33565) | (~w7463 & w33565);
assign w7468 = ~w7159 & ~w7161;
assign w7469 = ~w7162 & ~w7468;
assign w7470 = ~w7467 & w7469;
assign w7471 = w7467 & ~w7469;
assign w7472 = ~w7470 & ~w7471;
assign w7473 = ~w1475 & w6996;
assign w7474 = (w6446 & ~w1628) | (w6446 & w33566) | (~w1628 & w33566);
assign w7475 = (w6998 & ~w643) | (w6998 & w33567) | (~w643 & w33567);
assign w7476 = ~w7474 & ~w7475;
assign w7477 = ~w7473 & w7476;
assign w7478 = (w7477 & ~w4041) | (w7477 & w33568) | (~w4041 & w33568);
assign w7479 = a_14 & ~w7478;
assign w7480 = (~w4041 & w33569) | (~w4041 & w33570) | (w33569 & w33570);
assign w7481 = ~w7479 & ~w7480;
assign w7482 = w7472 & w7481;
assign w7483 = (~w7470 & ~w7472) | (~w7470 & w33571) | (~w7472 & w33571);
assign w7484 = ~w7209 & ~w7218;
assign w7485 = ~w7219 & ~w7484;
assign w7486 = ~w7483 & w7485;
assign w7487 = (~w7219 & ~w7485) | (~w7219 & w33572) | (~w7485 & w33572);
assign w7488 = (w7192 & ~w3904) | (w7192 & w33573) | (~w3904 & w33573);
assign w7489 = ~w7187 & w7190;
assign w7490 = ~w3958 & w7489;
assign w7491 = ~w7488 & ~w7490;
assign w7492 = (w7491 & ~w4073) | (w7491 & w33574) | (~w4073 & w33574);
assign w7493 = a_11 & ~w7492;
assign w7494 = (~w4073 & w33575) | (~w4073 & w33576) | (w33575 & w33576);
assign w7495 = ~w7493 & ~w7494;
assign w7496 = ~w7487 & w7495;
assign w7497 = ~w7177 & ~w7179;
assign w7498 = ~w7180 & ~w7497;
assign w7499 = w7487 & ~w7495;
assign w7500 = ~w7496 & ~w7499;
assign w7501 = w7498 & w7500;
assign w7502 = (~w7496 & ~w7500) | (~w7496 & w33577) | (~w7500 & w33577);
assign w7503 = ~w7200 & ~w7202;
assign w7504 = ~w7203 & ~w7503;
assign w7505 = w7502 & ~w7504;
assign w7506 = w7204 & ~w7206;
assign w7507 = ~w7207 & ~w7506;
assign w7508 = ~w7505 & w7507;
assign w7509 = ~w7508 & w33578;
assign w7510 = (w7489 & ~w1308) | (w7489 & w33579) | (~w1308 & w33579);
assign w7511 = w7184 & w7187;
assign w7512 = (w7511 & ~w3904) | (w7511 & w33580) | (~w3904 & w33580);
assign w7513 = ~w1397 & w7192;
assign w7514 = ~w7510 & ~w7513;
assign w7515 = ~w7512 & w7514;
assign w7516 = (w7515 & ~w3964) | (w7515 & w33581) | (~w3964 & w33581);
assign w7517 = a_11 & ~w7516;
assign w7518 = (~w3964 & w33582) | (~w3964 & w33583) | (w33582 & w33583);
assign w7519 = ~w7517 & ~w7518;
assign w7520 = ~w7463 & ~w7465;
assign w7521 = ~w7466 & ~w7520;
assign w7522 = ~w3813 & w6446;
assign w7523 = (w6996 & ~w643) | (w6996 & w33584) | (~w643 & w33584);
assign w7524 = (w6998 & ~w1628) | (w6998 & w33585) | (~w1628 & w33585);
assign w7525 = w4224 & w6447;
assign w7526 = ~w7522 & w33586;
assign w7527 = (a_14 & w7525) | (a_14 & w33587) | (w7525 & w33587);
assign w7528 = ~w7525 & w33588;
assign w7529 = ~w7527 & ~w7528;
assign w7530 = w7521 & w7529;
assign w7531 = ~w7521 & ~w7529;
assign w7532 = ~w7530 & ~w7531;
assign w7533 = w7448 & ~w7450;
assign w7534 = ~w7451 & ~w7533;
assign w7535 = ~w7254 & ~w7426;
assign w7536 = ~w7427 & ~w7535;
assign w7537 = ~w2306 & w5080;
assign w7538 = ~w2393 & w5286;
assign w7539 = (w5016 & ~w3538) | (w5016 & w33589) | (~w3538 & w33589);
assign w7540 = ~w7537 & ~w7538;
assign w7541 = ~w7539 & w7540;
assign w7542 = (w7541 & ~w5483) | (w7541 & w33590) | (~w5483 & w33590);
assign w7543 = a_23 & ~w7542;
assign w7544 = (~w5483 & w33591) | (~w5483 & w33592) | (w33591 & w33592);
assign w7545 = ~w7543 & ~w7544;
assign w7546 = w7536 & w7545;
assign w7547 = ~w3326 & w4638;
assign w7548 = (~w518 & ~w3267) | (~w518 & w33593) | (~w3267 & w33593);
assign w7549 = ~w3475 & w4666;
assign w7550 = ~w7547 & ~w7548;
assign w7551 = ~w7549 & w7550;
assign w7552 = (w7551 & ~w6108) | (w7551 & w33594) | (~w6108 & w33594);
assign w7553 = a_26 & ~w7552;
assign w7554 = (~w6108 & w33595) | (~w6108 & w33596) | (w33595 & w33596);
assign w7555 = ~w7553 & ~w7554;
assign w7556 = w7420 & w7425;
assign w7557 = w7555 & ~w7556;
assign w7558 = ~w7555 & w7556;
assign w7559 = ~w7557 & ~w7558;
assign w7560 = w7403 & w7559;
assign w7561 = ~w7403 & ~w7559;
assign w7562 = ~w7560 & ~w7561;
assign w7563 = ~w7555 & ~w7562;
assign w7564 = w7343 & ~w7361;
assign w7565 = ~w7362 & ~w7564;
assign w7566 = ~w3049 & w4666;
assign w7567 = ~w518 & ~w2917;
assign w7568 = ~w3007 & w4638;
assign w7569 = ~w7566 & ~w7567;
assign w7570 = ~w7568 & w7569;
assign w7571 = (w7570 & ~w6194) | (w7570 & w33597) | (~w6194 & w33597);
assign w7572 = a_26 & ~w7571;
assign w7573 = (~w6194 & w33598) | (~w6194 & w33599) | (w33598 & w33599);
assign w7574 = ~w7572 & ~w7573;
assign w7575 = ~w7565 & ~w7574;
assign w7576 = w7308 & ~w7341;
assign w7577 = ~w7342 & ~w7576;
assign w7578 = w1226 & w6545;
assign w7579 = w1226 & ~w6544;
assign w7580 = ~w2920 & w31601;
assign w7581 = ~w2917 & w4638;
assign w7582 = ~w3007 & w4666;
assign w7583 = ~w518 & ~w2835;
assign w7584 = ~w7581 & ~w7582;
assign w7585 = ~w7583 & w7584;
assign w7586 = ~w7580 & w7585;
assign w7587 = ~w7578 & w7586;
assign w7588 = ~a_26 & w7587;
assign w7589 = a_26 & ~w7587;
assign w7590 = ~w7588 & ~w7589;
assign w7591 = w7577 & w7590;
assign w7592 = ~w7577 & ~w7590;
assign w7593 = ~w7591 & ~w7592;
assign w7594 = ~w2677 & w4638;
assign w7595 = (~w518 & ~w2479) | (~w518 & w33600) | (~w2479 & w33600);
assign w7596 = ~w2546 & w4666;
assign w7597 = ~w7594 & ~w7595;
assign w7598 = w7597 & w33601;
assign w7599 = (w7598 & ~w6675) | (w7598 & w33602) | (~w6675 & w33602);
assign w7600 = (a_26 & ~w7597) | (a_26 & w33603) | (~w7597 & w33603);
assign w7601 = (~w7600 & ~w6675) | (~w7600 & w37564) | (~w6675 & w37564);
assign w7602 = ~w7599 & w7601;
assign w7603 = w1226 & w2677;
assign w7604 = w6595 & w7603;
assign w7605 = w1226 & ~w2677;
assign w7606 = ~w6595 & w7605;
assign w7607 = ~w2677 & w4666;
assign w7608 = (~w518 & ~w2600) | (~w518 & w31602) | (~w2600 & w31602);
assign w7609 = (w4638 & ~w2479) | (w4638 & w33604) | (~w2479 & w33604);
assign w7610 = ~w7607 & w33605;
assign w7611 = ~w7604 & ~w7606;
assign w7612 = w7610 & w7611;
assign w7613 = w1226 & ~w7287;
assign w7614 = (w4666 & ~w2479) | (w4666 & w31603) | (~w2479 & w31603);
assign w7615 = (w4638 & ~w2600) | (w4638 & w31604) | (~w2600 & w31604);
assign w7616 = ~w7614 & ~w7615;
assign w7617 = (~w1222 & ~w2600) | (~w1222 & w31605) | (~w2600 & w31605);
assign w7618 = a_26 & ~w7617;
assign w7619 = w7616 & w7618;
assign w7620 = ~w7613 & w7619;
assign w7621 = w7612 & w7620;
assign w7622 = ~w7335 & ~w7621;
assign w7623 = w7602 & ~w7622;
assign w7624 = w2680 & ~w6552;
assign w7625 = ~w6729 & ~w7624;
assign w7626 = (w4666 & ~w2766) | (w4666 & w33606) | (~w2766 & w33606);
assign w7627 = ~w2546 & w4638;
assign w7628 = ~w518 & ~w2677;
assign w7629 = ~w7626 & ~w7627;
assign w7630 = ~w7628 & w7629;
assign w7631 = (w7630 & ~w7625) | (w7630 & w31606) | (~w7625 & w31606);
assign w7632 = a_29 & w7335;
assign w7633 = w7334 & ~w7632;
assign w7634 = ~w7331 & w7633;
assign w7635 = w7268 & w7286;
assign w7636 = ~w7334 & w7632;
assign w7637 = ~w7635 & ~w7636;
assign w7638 = (a_26 & w7634) | (a_26 & w31607) | (w7634 & w31607);
assign w7639 = ~w7634 & w31608;
assign w7640 = ~w7638 & ~w7639;
assign w7641 = w7631 & w7640;
assign w7642 = ~w7631 & ~w7640;
assign w7643 = ~w7641 & ~w7642;
assign w7644 = ~w7623 & w7643;
assign w7645 = (~a_26 & w7634) | (~a_26 & w33607) | (w7634 & w33607);
assign w7646 = w7631 & ~w7645;
assign w7647 = ~w7631 & ~w7638;
assign w7648 = ~w7646 & ~w7647;
assign w7649 = ~w7644 & ~w7648;
assign w7650 = (w1226 & w6781) | (w1226 & w31609) | (w6781 & w31609);
assign w7651 = w1226 & w6778;
assign w7652 = ~w6726 & w7651;
assign w7653 = ~w2835 & w4638;
assign w7654 = ~w2917 & w4666;
assign w7655 = (~w518 & ~w2766) | (~w518 & w33608) | (~w2766 & w33608);
assign w7656 = ~w7653 & ~w7654;
assign w7657 = ~w7655 & w7656;
assign w7658 = ~w7652 & w7657;
assign w7659 = (a_26 & ~w7658) | (a_26 & w31610) | (~w7658 & w31610);
assign w7660 = w7658 & w31611;
assign w7661 = ~w7659 & ~w7660;
assign w7662 = w7319 & w7339;
assign w7663 = ~w7340 & ~w7662;
assign w7664 = w7318 & ~w7663;
assign w7665 = ~w7318 & w7663;
assign w7666 = ~w7664 & ~w7665;
assign w7667 = ~w7661 & w7666;
assign w7668 = (a_29 & w7331) | (a_29 & w33609) | (w7331 & w33609);
assign w7669 = ~w7330 & w7668;
assign w7670 = w7330 & ~w7668;
assign w7671 = ~w7669 & ~w7670;
assign w7672 = ~w2835 & w4666;
assign w7673 = (w4638 & ~w2766) | (w4638 & w31612) | (~w2766 & w31612);
assign w7674 = ~w518 & ~w2546;
assign w7675 = ~w7672 & ~w7673;
assign w7676 = (a_26 & ~w7675) | (a_26 & w31613) | (~w7675 & w31613);
assign w7677 = w7675 & w33610;
assign w7678 = ~w7676 & ~w7677;
assign w7679 = ~w6733 & w7678;
assign w7680 = ~a_26 & ~w1226;
assign w7681 = w7675 & w33611;
assign w7682 = ~w4403 & ~w7676;
assign w7683 = ~w7681 & w7682;
assign w7684 = w6733 & w7683;
assign w7685 = ~w7679 & ~w7684;
assign w7686 = w7671 & ~w7685;
assign w7687 = ~w7671 & w7685;
assign w7688 = ~w7686 & ~w7687;
assign w7689 = ~w7667 & w7688;
assign w7690 = w7649 & w7689;
assign w7691 = w7661 & ~w7666;
assign w7692 = ~w7686 & ~w7691;
assign w7693 = ~w7667 & ~w7692;
assign w7694 = ~w7690 & ~w7693;
assign w7695 = w7593 & ~w7694;
assign w7696 = w7565 & w7574;
assign w7697 = (~w7591 & ~w7565) | (~w7591 & w31614) | (~w7565 & w31614);
assign w7698 = ~w7695 & w7697;
assign w7699 = (~w7575 & w7695) | (~w7575 & w31615) | (w7695 & w31615);
assign w7700 = ~w7359 & ~w7362;
assign w7701 = ~w7285 & ~w7363;
assign w7702 = ~w3058 & w33612;
assign w7703 = w1226 & ~w6502;
assign w7704 = ~w3049 & w4638;
assign w7705 = ~w3139 & w4666;
assign w7706 = ~w518 & ~w3007;
assign w7707 = ~w7704 & ~w7705;
assign w7708 = ~w7706 & w7707;
assign w7709 = (~w3058 & w33613) | (~w3058 & w33614) | (w33613 & w33614);
assign w7710 = ~w7702 & w7709;
assign w7711 = ~a_26 & w7710;
assign w7712 = a_26 & ~w7710;
assign w7713 = ~w7711 & ~w7712;
assign w7714 = w7701 & w7713;
assign w7715 = w7700 & w7714;
assign w7716 = ~w7701 & w7713;
assign w7717 = ~w7700 & w7716;
assign w7718 = ~w7715 & ~w7717;
assign w7719 = ~w7699 & w7718;
assign w7720 = ~w7701 & ~w7713;
assign w7721 = w7700 & w7720;
assign w7722 = w7701 & ~w7713;
assign w7723 = ~w7700 & w7722;
assign w7724 = ~w7721 & ~w7723;
assign w7725 = ~w3139 & w4638;
assign w7726 = ~w518 & ~w3049;
assign w7727 = ~w3196 & w4666;
assign w7728 = ~w7725 & ~w7726;
assign w7729 = (a_26 & ~w7728) | (a_26 & w33615) | (~w7728 & w33615);
assign w7730 = w1226 & w6491;
assign w7731 = w7728 & w33616;
assign w7732 = ~w7730 & w7731;
assign w7733 = (~w7729 & ~w6491) | (~w7729 & w33617) | (~w6491 & w33617);
assign w7734 = ~w7732 & w7733;
assign w7735 = w7383 & ~w7734;
assign w7736 = ~w7383 & w7734;
assign w7737 = ~w7735 & ~w7736;
assign w7738 = w7365 & w7737;
assign w7739 = ~w7365 & ~w7737;
assign w7740 = ~w7738 & ~w7739;
assign w7741 = w7724 & ~w7740;
assign w7742 = ~w7719 & w7741;
assign w7743 = w7734 & w7740;
assign w7744 = (~w7381 & ~w7365) | (~w7381 & w33618) | (~w7365 & w33618);
assign w7745 = ~w3196 & w4638;
assign w7746 = ~w518 & ~w3139;
assign w7747 = (w4666 & ~w3267) | (w4666 & w33619) | (~w3267 & w33619);
assign w7748 = ~w7745 & ~w7746;
assign w7749 = w7748 & w33620;
assign w7750 = (w7749 & ~w6222) | (w7749 & w31617) | (~w6222 & w31617);
assign w7751 = w6222 & w33621;
assign w7752 = w7748 & w33622;
assign w7753 = (a_26 & ~w7748) | (a_26 & w33623) | (~w7748 & w33623);
assign w7754 = ~w7752 & ~w7753;
assign w7755 = ~w7750 & w7754;
assign w7756 = ~w7751 & w7755;
assign w7757 = w7392 & ~w7756;
assign w7758 = ~w7392 & w7756;
assign w7759 = ~w7757 & ~w7758;
assign w7760 = w7397 & ~w7759;
assign w7761 = ~w7397 & w7759;
assign w7762 = ~w7760 & ~w7761;
assign w7763 = w7744 & w7762;
assign w7764 = ~w7744 & ~w7762;
assign w7765 = ~w7763 & ~w7764;
assign w7766 = ~w7743 & ~w7765;
assign w7767 = ~w7742 & w7766;
assign w7768 = ~w7756 & w7765;
assign w7769 = ~w7767 & ~w7768;
assign w7770 = (~w7400 & w7384) | (~w7400 & w33624) | (w7384 & w33624);
assign w7771 = w1226 & w5902;
assign w7772 = w1226 & ~w5900;
assign w7773 = (~w3058 & w33625) | (~w3058 & w33626) | (w33625 & w33626);
assign w7774 = (w4638 & ~w3267) | (w4638 & w33627) | (~w3267 & w33627);
assign w7775 = ~w518 & ~w3196;
assign w7776 = ~w3326 & w4666;
assign w7777 = ~w7774 & ~w7775;
assign w7778 = ~w7776 & w7777;
assign w7779 = ~w7773 & w7778;
assign w7780 = ~w7771 & w7779;
assign w7781 = ~a_26 & w7780;
assign w7782 = a_26 & ~w7780;
assign w7783 = ~w7781 & ~w7782;
assign w7784 = w7266 & ~w7783;
assign w7785 = ~w7266 & w7783;
assign w7786 = ~w7784 & ~w7785;
assign w7787 = w7257 & ~w7786;
assign w7788 = ~w7257 & w7786;
assign w7789 = ~w7787 & ~w7788;
assign w7790 = w7770 & w7789;
assign w7791 = ~w7770 & ~w7789;
assign w7792 = ~w7790 & ~w7791;
assign w7793 = ~w7767 & w33628;
assign w7794 = w7783 & ~w7792;
assign w7795 = w7562 & ~w7794;
assign w7796 = ~w7793 & w7795;
assign w7797 = ~w7563 & ~w7796;
assign w7798 = ~w7536 & ~w7545;
assign w7799 = ~w7546 & ~w7798;
assign w7800 = w7797 & w7799;
assign w7801 = (~w7546 & ~w7797) | (~w7546 & w33629) | (~w7797 & w33629);
assign w7802 = ~w7429 & ~w7430;
assign w7803 = w7439 & w7802;
assign w7804 = ~w7439 & ~w7802;
assign w7805 = ~w7803 & ~w7804;
assign w7806 = w7801 & ~w7805;
assign w7807 = ~w2075 & w5308;
assign w7808 = (w5816 & ~w2235) | (w5816 & w33630) | (~w2235 & w33630);
assign w7809 = ~w2148 & w5818;
assign w7810 = ~w7808 & ~w7809;
assign w7811 = ~w7807 & w7810;
assign w7812 = (w7811 & ~w4962) | (w7811 & w33631) | (~w4962 & w33631);
assign w7813 = a_20 & ~w7812;
assign w7814 = (~w4962 & w33632) | (~w4962 & w33633) | (w33632 & w33633);
assign w7815 = ~w7813 & ~w7814;
assign w7816 = ~w7801 & w7805;
assign w7817 = ~w7806 & ~w7816;
assign w7818 = ~w7815 & w7817;
assign w7819 = (~w7806 & ~w7817) | (~w7806 & w33634) | (~w7817 & w33634);
assign w7820 = ~w7441 & ~w7442;
assign w7821 = w7444 & w7820;
assign w7822 = ~w7444 & ~w7820;
assign w7823 = ~w7821 & ~w7822;
assign w7824 = w7819 & w7823;
assign w7825 = (w6059 & ~w3658) | (w6059 & w33635) | (~w3658 & w33635);
assign w7826 = (w6061 & ~w2005) | (w6061 & w33636) | (~w2005 & w33636);
assign w7827 = (w6304 & ~w1913) | (w6304 & w33637) | (~w1913 & w33637);
assign w7828 = ~w7826 & ~w7827;
assign w7829 = ~w7825 & w7828;
assign w7830 = (w7829 & w4578) | (w7829 & w33638) | (w4578 & w33638);
assign w7831 = a_17 & ~w7830;
assign w7832 = (w4578 & w33639) | (w4578 & w33640) | (w33639 & w33640);
assign w7833 = ~w7831 & ~w7832;
assign w7834 = ~w7819 & ~w7823;
assign w7835 = ~w7824 & ~w7834;
assign w7836 = w7833 & w7835;
assign w7837 = (~w7824 & ~w7835) | (~w7824 & w33641) | (~w7835 & w33641);
assign w7838 = w7534 & ~w7837;
assign w7839 = ~w7534 & w7837;
assign w7840 = ~w7838 & ~w7839;
assign w7841 = (w6061 & ~w1913) | (w6061 & w33642) | (~w1913 & w33642);
assign w7842 = (w6059 & ~w2005) | (w6059 & w33643) | (~w2005 & w33643);
assign w7843 = (w6304 & ~w1714) | (w6304 & w33458) | (~w1714 & w33458);
assign w7844 = ~w7841 & ~w7842;
assign w7845 = ~w7843 & w7844;
assign w7846 = (w7845 & ~w4592) | (w7845 & w33644) | (~w4592 & w33644);
assign w7847 = a_17 & ~w7846;
assign w7848 = (~w4592 & w33645) | (~w4592 & w33646) | (w33645 & w33646);
assign w7849 = ~w7847 & ~w7848;
assign w7850 = w7840 & w7849;
assign w7851 = (~w7838 & ~w7840) | (~w7838 & w33647) | (~w7840 & w33647);
assign w7852 = w7532 & ~w7851;
assign w7853 = (~w7530 & ~w7532) | (~w7530 & w33648) | (~w7532 & w33648);
assign w7854 = ~w7519 & w7853;
assign w7855 = ~w7472 & ~w7481;
assign w7856 = ~w7482 & ~w7855;
assign w7857 = w7519 & ~w7853;
assign w7858 = ~w7854 & ~w7857;
assign w7859 = ~w7856 & w7858;
assign w7860 = (w7489 & ~w3904) | (w7489 & w33649) | (~w3904 & w33649);
assign w7861 = ~w3958 & w7511;
assign w7862 = (w7192 & ~w1308) | (w7192 & w33650) | (~w1308 & w33650);
assign w7863 = ~w7861 & ~w7862;
assign w7864 = ~w7860 & w7863;
assign w7865 = (w7864 & ~w3943) | (w7864 & w33651) | (~w3943 & w33651);
assign w7866 = a_11 & ~w7865;
assign w7867 = (~w3943 & w33652) | (~w3943 & w33653) | (w33652 & w33653);
assign w7868 = ~w7866 & ~w7867;
assign w7869 = ~w7859 & w33654;
assign w7870 = w7483 & ~w7485;
assign w7871 = ~w7486 & ~w7870;
assign w7872 = (~w7868 & w7859) | (~w7868 & w33655) | (w7859 & w33655);
assign w7873 = ~w7869 & ~w7872;
assign w7874 = w7871 & w7873;
assign w7875 = (~w7869 & ~w7873) | (~w7869 & w33656) | (~w7873 & w33656);
assign w7876 = ~w7498 & ~w7500;
assign w7877 = ~w7501 & ~w7876;
assign w7878 = w7875 & ~w7877;
assign w7879 = ~w7871 & ~w7873;
assign w7880 = ~w7874 & ~w7879;
assign w7881 = ~w7532 & w7851;
assign w7882 = ~w7852 & ~w7881;
assign w7883 = (w6446 & ~w1807) | (w6446 & w33657) | (~w1807 & w33657);
assign w7884 = (w6996 & ~w1628) | (w6996 & w33658) | (~w1628 & w33658);
assign w7885 = ~w3813 & w6998;
assign w7886 = ~w7883 & ~w7884;
assign w7887 = ~w7885 & w7886;
assign w7888 = (w7887 & ~w4244) | (w7887 & w33659) | (~w4244 & w33659);
assign w7889 = a_14 & ~w7888;
assign w7890 = (~w4244 & w33660) | (~w4244 & w33661) | (w33660 & w33661);
assign w7891 = ~w7889 & ~w7890;
assign w7892 = ~w7833 & ~w7835;
assign w7893 = ~w7836 & ~w7892;
assign w7894 = ~w7797 & ~w7799;
assign w7895 = ~w7800 & ~w7894;
assign w7896 = ~w2075 & w5818;
assign w7897 = ~w2148 & w5816;
assign w7898 = ~w3615 & w5308;
assign w7899 = ~w7897 & ~w7898;
assign w7900 = ~w7896 & w7899;
assign w7901 = (w7900 & ~w5242) | (w7900 & w33662) | (~w5242 & w33662);
assign w7902 = a_20 & ~w7901;
assign w7903 = (~w5242 & w33663) | (~w5242 & w33664) | (w33663 & w33664);
assign w7904 = ~w7902 & ~w7903;
assign w7905 = w7895 & w7904;
assign w7906 = ~w7895 & ~w7904;
assign w7907 = ~w7905 & ~w7906;
assign w7908 = (~w7591 & w7694) | (~w7591 & w31618) | (w7694 & w31618);
assign w7909 = ~w7575 & ~w7696;
assign w7910 = ~w3196 & w5080;
assign w7911 = (w5286 & ~w3267) | (w5286 & w33665) | (~w3267 & w33665);
assign w7912 = ~w3139 & w5016;
assign w7913 = w6222 & w33666;
assign w7914 = ~w7910 & ~w7911;
assign w7915 = ~w7912 & w7914;
assign w7916 = (a_23 & w7913) | (a_23 & w33667) | (w7913 & w33667);
assign w7917 = ~w7913 & w33668;
assign w7918 = ~w7916 & ~w7917;
assign w7919 = ~w7909 & w7918;
assign w7920 = ~w7908 & w7919;
assign w7921 = w7909 & w7918;
assign w7922 = w7908 & w7921;
assign w7923 = ~w7920 & ~w7922;
assign w7924 = ~w7909 & ~w7918;
assign w7925 = ~w7921 & ~w7924;
assign w7926 = w7908 & w7925;
assign w7927 = ~w7908 & ~w7925;
assign w7928 = ~w7926 & ~w7927;
assign w7929 = w7923 & w7928;
assign w7930 = w7623 & ~w7643;
assign w7931 = ~w7644 & ~w7930;
assign w7932 = w5017 & w6545;
assign w7933 = w5017 & ~w6544;
assign w7934 = ~w2920 & w31619;
assign w7935 = ~w2835 & w5016;
assign w7936 = ~w3007 & w5286;
assign w7937 = ~w2917 & w5080;
assign w7938 = ~w7935 & ~w7936;
assign w7939 = ~w7937 & w7938;
assign w7940 = ~w7934 & w7939;
assign w7941 = ~w7932 & w7940;
assign w7942 = ~a_23 & w7941;
assign w7943 = a_23 & ~w7941;
assign w7944 = ~w7942 & ~w7943;
assign w7945 = w7931 & ~w7944;
assign w7946 = a_26 & w7617;
assign w7947 = w7616 & ~w7946;
assign w7948 = ~w7613 & w7947;
assign w7949 = (a_26 & w7613) | (a_26 & w33669) | (w7613 & w33669);
assign w7950 = ~w7612 & w7949;
assign w7951 = w7612 & ~w7949;
assign w7952 = ~w7950 & ~w7951;
assign w7953 = ~w2835 & w5286;
assign w7954 = ~w2546 & w5016;
assign w7955 = (w5080 & ~w2766) | (w5080 & w33670) | (~w2766 & w33670);
assign w7956 = ~w7953 & ~w7954;
assign w7957 = (a_23 & ~w7956) | (a_23 & w31620) | (~w7956 & w31620);
assign w7958 = w7956 & w33671;
assign w7959 = ~w7957 & ~w7958;
assign w7960 = ~w6733 & w7959;
assign w7961 = w504 & w5014;
assign w7962 = ~a_23 & ~w5017;
assign w7963 = w7956 & w33672;
assign w7964 = ~w7957 & ~w7961;
assign w7965 = ~w7963 & w7964;
assign w7966 = w6733 & w7965;
assign w7967 = ~w7960 & ~w7966;
assign w7968 = ~w7952 & w7967;
assign w7969 = ~w2677 & w6595;
assign w7970 = ~w6671 & ~w7969;
assign w7971 = w5017 & w7970;
assign w7972 = (w5080 & ~w2479) | (w5080 & w33673) | (~w2479 & w33673);
assign w7973 = ~w2677 & w5286;
assign w7974 = (w5016 & ~w2600) | (w5016 & w33674) | (~w2600 & w33674);
assign w7975 = ~w7973 & w33675;
assign w7976 = ~w7971 & w7975;
assign w7977 = w5017 & ~w7287;
assign w7978 = (w5286 & ~w2479) | (w5286 & w31621) | (~w2479 & w31621);
assign w7979 = (w5080 & ~w2600) | (w5080 & w31622) | (~w2600 & w31622);
assign w7980 = ~w7978 & ~w7979;
assign w7981 = (w504 & ~w2600) | (w504 & w31623) | (~w2600 & w31623);
assign w7982 = a_23 & w7981;
assign w7983 = w7980 & ~w7982;
assign w7984 = ~w7977 & w7983;
assign w7985 = ~w7977 & w31624;
assign w7986 = (~w7617 & ~w7976) | (~w7617 & w31625) | (~w7976 & w31625);
assign w7987 = ~w2546 & w5286;
assign w7988 = (w5016 & ~w2479) | (w5016 & w33676) | (~w2479 & w33676);
assign w7989 = ~w2677 & w5080;
assign w7990 = ~w7987 & ~w7988;
assign w7991 = (a_23 & ~w7990) | (a_23 & w33677) | (~w7990 & w33677);
assign w7992 = w5017 & w6675;
assign w7993 = w7990 & w33678;
assign w7994 = ~w7992 & w7993;
assign w7995 = (~w7991 & ~w6675) | (~w7991 & w33679) | (~w6675 & w33679);
assign w7996 = ~w7994 & w7995;
assign w7997 = ~w7986 & w7996;
assign w7998 = (w5286 & ~w2766) | (w5286 & w33680) | (~w2766 & w33680);
assign w7999 = ~w2677 & w5016;
assign w8000 = ~w2546 & w5080;
assign w8001 = ~w7998 & ~w7999;
assign w8002 = ~w8000 & w8001;
assign w8003 = (w8002 & ~w7625) | (w8002 & w31626) | (~w7625 & w31626);
assign w8004 = w4403 & w7286;
assign w8005 = ~w7616 & w7946;
assign w8006 = ~w8004 & ~w8005;
assign w8007 = ~w7948 & w31627;
assign w8008 = (a_23 & w7948) | (a_23 & w31628) | (w7948 & w31628);
assign w8009 = ~w8007 & ~w8008;
assign w8010 = w8003 & w8009;
assign w8011 = ~w8003 & ~w8009;
assign w8012 = ~w8010 & ~w8011;
assign w8013 = w7997 & w8012;
assign w8014 = w7952 & ~w7967;
assign w8015 = ~w7948 & w33681;
assign w8016 = w8003 & ~w8015;
assign w8017 = ~w8003 & ~w8007;
assign w8018 = ~w8016 & ~w8017;
assign w8019 = ~w8014 & ~w8018;
assign w8020 = (~w7968 & ~w8019) | (~w7968 & w31629) | (~w8019 & w31629);
assign w8021 = (w5017 & w6781) | (w5017 & w32439) | (w6781 & w32439);
assign w8022 = w5017 & w6778;
assign w8023 = ~w6726 & w8022;
assign w8024 = ~w2835 & w5080;
assign w8025 = ~w2917 & w5286;
assign w8026 = (w5016 & ~w2766) | (w5016 & w33682) | (~w2766 & w33682);
assign w8027 = ~w8024 & ~w8025;
assign w8028 = ~w8026 & w8027;
assign w8029 = ~w8023 & w8028;
assign w8030 = w8029 & w32440;
assign w8031 = (a_23 & ~w8029) | (a_23 & w32441) | (~w8029 & w32441);
assign w8032 = ~w8030 & ~w8031;
assign w8033 = w7335 & w7621;
assign w8034 = ~w7622 & ~w8033;
assign w8035 = w7602 & ~w8034;
assign w8036 = ~w7602 & w8034;
assign w8037 = ~w8035 & ~w8036;
assign w8038 = w8032 & ~w8037;
assign w8039 = ~w8032 & w8037;
assign w8040 = ~w8038 & ~w8039;
assign w8041 = w8020 & w8040;
assign w8042 = ~w7931 & w7944;
assign w8043 = ~w8038 & ~w8042;
assign w8044 = ~w8041 & w8043;
assign w8045 = ~w7945 & ~w8044;
assign w8046 = ~w7648 & ~w7687;
assign w8047 = (~w7686 & ~w8046) | (~w7686 & w31630) | (~w8046 & w31630);
assign w8048 = ~w7667 & ~w7691;
assign w8049 = ~w3058 & w33683;
assign w8050 = w5017 & ~w6502;
assign w8051 = ~w3007 & w5016;
assign w8052 = ~w3139 & w5286;
assign w8053 = ~w3049 & w5080;
assign w8054 = ~w8051 & ~w8052;
assign w8055 = ~w8053 & w8054;
assign w8056 = (~w3058 & w33684) | (~w3058 & w33685) | (w33684 & w33685);
assign w8057 = ~w8049 & w8056;
assign w8058 = ~a_23 & w8057;
assign w8059 = a_23 & ~w8057;
assign w8060 = ~w8058 & ~w8059;
assign w8061 = ~w8048 & ~w8060;
assign w8062 = w8047 & w8061;
assign w8063 = w8048 & ~w8060;
assign w8064 = ~w8047 & w8063;
assign w8065 = ~w8062 & ~w8064;
assign w8066 = ~w3049 & w5286;
assign w8067 = ~w2917 & w5016;
assign w8068 = ~w3007 & w5080;
assign w8069 = ~w8066 & ~w8067;
assign w8070 = w8069 & w33686;
assign w8071 = w6194 & w7961;
assign w8072 = w8069 & w33687;
assign w8073 = (a_23 & ~w8069) | (a_23 & w33688) | (~w8069 & w33688);
assign w8074 = ~w8072 & ~w8073;
assign w8075 = (w8074 & w6194) | (w8074 & w31632) | (w6194 & w31632);
assign w8076 = ~w8071 & w8075;
assign w8077 = w7688 & w8076;
assign w8078 = ~w7688 & ~w8076;
assign w8079 = ~w8077 & ~w8078;
assign w8080 = w7649 & w8079;
assign w8081 = ~w7649 & ~w8079;
assign w8082 = ~w8080 & ~w8081;
assign w8083 = w8065 & w8082;
assign w8084 = w8045 & w8083;
assign w8085 = w8048 & w8060;
assign w8086 = w8047 & w8085;
assign w8087 = ~w8048 & w8060;
assign w8088 = ~w8047 & w8087;
assign w8089 = ~w8086 & ~w8088;
assign w8090 = w7649 & ~w7688;
assign w8091 = ~w7649 & w7688;
assign w8092 = ~w8090 & ~w8091;
assign w8093 = w8076 & ~w8092;
assign w8094 = w8089 & ~w8093;
assign w8095 = w8065 & ~w8094;
assign w8096 = ~w8084 & ~w8095;
assign w8097 = ~w3196 & w5286;
assign w8098 = ~w3049 & w5016;
assign w8099 = ~w3139 & w5080;
assign w8100 = ~w8097 & ~w8098;
assign w8101 = (a_23 & ~w8100) | (a_23 & w33689) | (~w8100 & w33689);
assign w8102 = w5017 & w6491;
assign w8103 = w8100 & w33690;
assign w8104 = ~w8102 & w8103;
assign w8105 = (~w8101 & ~w6491) | (~w8101 & w33691) | (~w6491 & w33691);
assign w8106 = ~w8104 & w8105;
assign w8107 = w7593 & ~w8106;
assign w8108 = ~w7593 & w8106;
assign w8109 = ~w8107 & ~w8108;
assign w8110 = w7694 & w8109;
assign w8111 = ~w7694 & ~w8109;
assign w8112 = ~w8110 & ~w8111;
assign w8113 = ~w8096 & w8112;
assign w8114 = w8106 & ~w8112;
assign w8115 = w7923 & ~w8114;
assign w8116 = ~w8113 & w8115;
assign w8117 = ~w7929 & ~w8116;
assign w8118 = w7718 & w7724;
assign w8119 = ~w3326 & w5286;
assign w8120 = (w5080 & ~w3267) | (w5080 & w33692) | (~w3267 & w33692);
assign w8121 = ~w3196 & w5016;
assign w8122 = ~w8120 & ~w8121;
assign w8123 = ~w8119 & w8122;
assign w8124 = (w8123 & w5903) | (w8123 & w33693) | (w5903 & w33693);
assign w8125 = a_23 & ~w8124;
assign w8126 = (w5903 & w33694) | (w5903 & w33695) | (w33694 & w33695);
assign w8127 = ~w8125 & ~w8126;
assign w8128 = w8118 & ~w8127;
assign w8129 = ~w8118 & w8127;
assign w8130 = ~w8128 & ~w8129;
assign w8131 = w7699 & w8130;
assign w8132 = ~w7699 & ~w8130;
assign w8133 = ~w8131 & ~w8132;
assign w8134 = w8117 & ~w8133;
assign w8135 = w8127 & w8133;
assign w8136 = ~w7575 & w7724;
assign w8137 = ~w7698 & w8136;
assign w8138 = w7718 & ~w8137;
assign w8139 = ~w8137 & w31633;
assign w8140 = ~w3326 & w5080;
assign w8141 = (w5016 & ~w3267) | (w5016 & w33696) | (~w3267 & w33696);
assign w8142 = ~w3475 & w5286;
assign w8143 = ~w8140 & ~w8141;
assign w8144 = ~w8142 & w8143;
assign w8145 = (w8144 & ~w6108) | (w8144 & w33697) | (~w6108 & w33697);
assign w8146 = ~a_23 & w8145;
assign w8147 = (w6108 & w33698) | (w6108 & w33699) | (w33698 & w33699);
assign w8148 = ~w8146 & ~w8147;
assign w8149 = ~w7742 & w8148;
assign w8150 = ~w8139 & w8149;
assign w8151 = ~w8135 & ~w8150;
assign w8152 = ~w8134 & w8151;
assign w8153 = w7724 & ~w8148;
assign w8154 = ~w7740 & w8153;
assign w8155 = ~w7719 & w8154;
assign w8156 = w7740 & ~w8148;
assign w8157 = w8138 & w8156;
assign w8158 = ~w8155 & ~w8157;
assign w8159 = ~w7742 & ~w7743;
assign w8160 = ~w3475 & w5080;
assign w8161 = ~w3403 & w5286;
assign w8162 = ~w3326 & w5016;
assign w8163 = ~w8160 & ~w8161;
assign w8164 = ~w8162 & w8163;
assign w8165 = (w8164 & ~w5923) | (w8164 & w33700) | (~w5923 & w33700);
assign w8166 = a_23 & ~w8165;
assign w8167 = (~w5923 & w33701) | (~w5923 & w33702) | (w33701 & w33702);
assign w8168 = ~w8166 & ~w8167;
assign w8169 = w7765 & w8168;
assign w8170 = ~w7765 & ~w8168;
assign w8171 = ~w8169 & ~w8170;
assign w8172 = ~w8159 & w8171;
assign w8173 = ~w7767 & ~w8168;
assign w8174 = ~w8172 & w8173;
assign w8175 = w8158 & ~w8174;
assign w8176 = ~w8152 & w8175;
assign w8177 = w8159 & ~w8171;
assign w8178 = ~w8172 & ~w8177;
assign w8179 = w8168 & w8178;
assign w8180 = ~w3403 & w5080;
assign w8181 = (w5286 & ~w3538) | (w5286 & w33703) | (~w3538 & w33703);
assign w8182 = ~w3475 & w5016;
assign w8183 = ~w8180 & ~w8181;
assign w8184 = ~w8182 & w8183;
assign w8185 = (w8184 & ~w5652) | (w8184 & w33704) | (~w5652 & w33704);
assign w8186 = a_23 & ~w8185;
assign w8187 = (~w5652 & w33705) | (~w5652 & w33706) | (w33705 & w33706);
assign w8188 = ~w8186 & ~w8187;
assign w8189 = ~w7792 & w8188;
assign w8190 = w7792 & ~w8188;
assign w8191 = ~w8189 & ~w8190;
assign w8192 = w7769 & w8191;
assign w8193 = ~w7769 & ~w8191;
assign w8194 = ~w8192 & ~w8193;
assign w8195 = ~w8179 & ~w8194;
assign w8196 = ~w8176 & w8195;
assign w8197 = ~w8188 & w8194;
assign w8198 = (~w8197 & w8176) | (~w8197 & w31634) | (w8176 & w31634);
assign w8199 = ~w7793 & ~w7794;
assign w8200 = ~w3403 & w5016;
assign w8201 = ~w2306 & w5286;
assign w8202 = (w5080 & ~w3538) | (w5080 & w33707) | (~w3538 & w33707);
assign w8203 = ~w8201 & ~w8202;
assign w8204 = ~w8200 & w8203;
assign w8205 = (w8204 & ~w5706) | (w8204 & w33708) | (~w5706 & w33708);
assign w8206 = a_23 & w8205;
assign w8207 = (w5706 & w33709) | (w5706 & w33710) | (w33709 & w33710);
assign w8208 = ~w8206 & ~w8207;
assign w8209 = ~w7562 & w8208;
assign w8210 = w7562 & ~w8208;
assign w8211 = ~w8209 & ~w8210;
assign w8212 = w8199 & w8211;
assign w8213 = ~w8199 & ~w8211;
assign w8214 = ~w8212 & ~w8213;
assign w8215 = w8208 & w8214;
assign w8216 = (~w8215 & w8198) | (~w8215 & w33711) | (w8198 & w33711);
assign w8217 = w7907 & w8216;
assign w8218 = ~w7905 & ~w8217;
assign w8219 = w7815 & ~w7817;
assign w8220 = ~w7818 & ~w8219;
assign w8221 = ~w8218 & ~w8220;
assign w8222 = w8218 & w8220;
assign w8223 = ~w8221 & ~w8222;
assign w8224 = (w6061 & ~w3658) | (w6061 & w33712) | (~w3658 & w33712);
assign w8225 = (w6059 & ~w3712) | (w6059 & w33713) | (~w3712 & w33713);
assign w8226 = (w6304 & ~w2005) | (w6304 & w33714) | (~w2005 & w33714);
assign w8227 = (w6063 & w4790) | (w6063 & w33715) | (w4790 & w33715);
assign w8228 = ~w8225 & ~w8226;
assign w8229 = ~w8224 & w8228;
assign w8230 = ~w8227 & w33716;
assign w8231 = (~a_17 & w8227) | (~a_17 & w33717) | (w8227 & w33717);
assign w8232 = ~w8230 & ~w8231;
assign w8233 = w8223 & ~w8232;
assign w8234 = (~w8221 & ~w8223) | (~w8221 & w33718) | (~w8223 & w33718);
assign w8235 = w7893 & ~w8234;
assign w8236 = ~w7893 & w8234;
assign w8237 = ~w3813 & w6996;
assign w8238 = (w6998 & ~w1807) | (w6998 & w33719) | (~w1807 & w33719);
assign w8239 = (w6446 & ~w1714) | (w6446 & w33566) | (~w1714 & w33566);
assign w8240 = w4508 & w6447;
assign w8241 = ~w8237 & w33720;
assign w8242 = (a_14 & w8240) | (a_14 & w33721) | (w8240 & w33721);
assign w8243 = ~w8240 & w33722;
assign w8244 = ~w8242 & ~w8243;
assign w8245 = (w8244 & ~w8234) | (w8244 & w33723) | (~w8234 & w33723);
assign w8246 = ~w8235 & ~w8245;
assign w8247 = w7891 & ~w8246;
assign w8248 = ~w7891 & w8246;
assign w8249 = ~w7840 & ~w7849;
assign w8250 = ~w7850 & ~w8249;
assign w8251 = ~w8248 & w8250;
assign w8252 = ~w8247 & ~w8251;
assign w8253 = w7882 & ~w8252;
assign w8254 = ~w7882 & w8252;
assign w8255 = ~w8253 & ~w8254;
assign w8256 = (w7511 & ~w1308) | (w7511 & w33724) | (~w1308 & w33724);
assign w8257 = ~w1397 & w7489;
assign w8258 = ~w1475 & w7192;
assign w8259 = ~w8256 & ~w8257;
assign w8260 = ~w8258 & w8259;
assign w8261 = (w8260 & ~w3834) | (w8260 & w33725) | (~w3834 & w33725);
assign w8262 = a_11 & ~w8261;
assign w8263 = (~w3834 & w33726) | (~w3834 & w33727) | (w33726 & w33727);
assign w8264 = ~w8262 & ~w8263;
assign w8265 = w8255 & w8264;
assign w8266 = (~w8253 & ~w8255) | (~w8253 & w33728) | (~w8255 & w33728);
assign w8267 = a_7 & ~a_8;
assign w8268 = ~a_7 & a_8;
assign w8269 = ~w8267 & ~w8268;
assign w8270 = a_5 & ~a_6;
assign w8271 = ~a_5 & a_6;
assign w8272 = ~w8270 & ~w8271;
assign w8273 = ~a_6 & ~a_7;
assign w8274 = a_6 & a_7;
assign w8275 = ~w8273 & ~w8274;
assign w8276 = w8272 & ~w8275;
assign w8277 = ~w8269 & w8276;
assign w8278 = ~w8269 & ~w8272;
assign w8279 = (~w3828 & w33731) | (~w3828 & w33732) | (w33731 & w33732);
assign w8280 = ~w8279 & w33733;
assign w8281 = (a_8 & w8279) | (a_8 & w33734) | (w8279 & w33734);
assign w8282 = ~w8280 & ~w8281;
assign w8283 = w8266 & w8282;
assign w8284 = w7856 & ~w7858;
assign w8285 = ~w7859 & ~w8284;
assign w8286 = ~w8266 & ~w8282;
assign w8287 = ~w8283 & ~w8286;
assign w8288 = w8285 & w8287;
assign w8289 = (~w8283 & ~w8287) | (~w8283 & w33735) | (~w8287 & w33735);
assign w8290 = w7880 & w8289;
assign w8291 = ~w7875 & w7877;
assign w8292 = ~w7878 & ~w8291;
assign w8293 = ~w8290 & w8292;
assign w8294 = ~w7878 & ~w8293;
assign w8295 = w8269 & ~w8272;
assign w8296 = (w8295 & ~w3712) | (w8295 & w33736) | (~w3712 & w33736);
assign w8297 = ~w2148 & w8277;
assign w8298 = w8272 & w8275;
assign w8299 = (w8298 & ~w2235) | (w8298 & w33737) | (~w2235 & w33737);
assign w8300 = w5103 & w8278;
assign w8301 = ~w8297 & w33738;
assign w8302 = (a_8 & w8300) | (a_8 & w33739) | (w8300 & w33739);
assign w8303 = ~w8300 & w33740;
assign w8304 = ~w8302 & ~w8303;
assign w8305 = ~w2835 & w5816;
assign w8306 = ~w2546 & w5308;
assign w8307 = (w5818 & ~w2766) | (w5818 & w33741) | (~w2766 & w33741);
assign w8308 = ~w8305 & ~w8306;
assign w8309 = w8308 & w33742;
assign w8310 = (w8309 & ~w6733) | (w8309 & w31635) | (~w6733 & w31635);
assign w8311 = w5300 & w5305;
assign w8312 = (a_20 & ~w8308) | (a_20 & w33743) | (~w8308 & w33743);
assign w8313 = (~w8312 & ~w6733) | (~w8312 & w31636) | (~w6733 & w31636);
assign w8314 = ~w8310 & w8313;
assign w8315 = (a_23 & w7977) | (a_23 & w33744) | (w7977 & w33744);
assign w8316 = ~w7976 & w8315;
assign w8317 = w7976 & ~w8315;
assign w8318 = ~w8316 & ~w8317;
assign w8319 = w8314 & w8318;
assign w8320 = ~w8314 & ~w8318;
assign w8321 = ~w8319 & ~w8320;
assign w8322 = w5309 & w7970;
assign w8323 = (w5818 & ~w2479) | (w5818 & w33745) | (~w2479 & w33745);
assign w8324 = ~w2677 & w5816;
assign w8325 = (w5308 & ~w2600) | (w5308 & w33746) | (~w2600 & w33746);
assign w8326 = ~w8324 & w33747;
assign w8327 = ~w8322 & w8326;
assign w8328 = w5309 & ~w7287;
assign w8329 = (w5816 & ~w2479) | (w5816 & w31637) | (~w2479 & w31637);
assign w8330 = (w5818 & ~w2600) | (w5818 & w31638) | (~w2600 & w31638);
assign w8331 = ~w8329 & ~w8330;
assign w8332 = (w5300 & ~w2600) | (w5300 & w31639) | (~w2600 & w31639);
assign w8333 = a_20 & w8332;
assign w8334 = w8331 & ~w8333;
assign w8335 = ~w8328 & w8334;
assign w8336 = ~w8328 & w31640;
assign w8337 = (~w7981 & ~w8327) | (~w7981 & w31641) | (~w8327 & w31641);
assign w8338 = w6675 & w8311;
assign w8339 = w5300 & w5306;
assign w8340 = w6675 & w8339;
assign w8341 = ~w2677 & w5818;
assign w8342 = (w5308 & ~w2479) | (w5308 & w33748) | (~w2479 & w33748);
assign w8343 = ~w2546 & w5816;
assign w8344 = ~w8341 & ~w8342;
assign w8345 = w8344 & w33749;
assign w8346 = (~a_20 & ~w8344) | (~a_20 & w33750) | (~w8344 & w33750);
assign w8347 = ~w8345 & ~w8346;
assign w8348 = ~w8340 & w8347;
assign w8349 = ~w8338 & ~w8348;
assign w8350 = ~w8337 & w8349;
assign w8351 = (w5816 & ~w2766) | (w5816 & w33751) | (~w2766 & w33751);
assign w8352 = ~w2677 & w5308;
assign w8353 = ~w2546 & w5818;
assign w8354 = ~w8351 & ~w8352;
assign w8355 = ~w8353 & w8354;
assign w8356 = (w8355 & ~w7625) | (w8355 & w31642) | (~w7625 & w31642);
assign w8357 = w7286 & w7961;
assign w8358 = ~w7980 & w7982;
assign w8359 = ~w8357 & ~w8358;
assign w8360 = ~w7984 & w8359;
assign w8361 = (a_20 & w7984) | (a_20 & w31643) | (w7984 & w31643);
assign w8362 = ~w7984 & w31644;
assign w8363 = ~w8361 & ~w8362;
assign w8364 = w8356 & w8363;
assign w8365 = ~w8356 & ~w8363;
assign w8366 = ~w8364 & ~w8365;
assign w8367 = ~w8350 & w8366;
assign w8368 = ~w8360 & ~w8366;
assign w8369 = ~w8367 & ~w8368;
assign w8370 = w8321 & w8369;
assign w8371 = ~w8321 & ~w8369;
assign w8372 = ~w8370 & ~w8371;
assign w8373 = ~w3049 & w6304;
assign w8374 = ~w3007 & w6061;
assign w8375 = ~w2917 & w6059;
assign w8376 = ~w8373 & ~w8374;
assign w8377 = ~w8375 & w8376;
assign w8378 = (w8377 & ~w6194) | (w8377 & w33752) | (~w6194 & w33752);
assign w8379 = a_17 & w8378;
assign w8380 = (w6194 & w33753) | (w6194 & w33754) | (w33753 & w33754);
assign w8381 = ~w8379 & ~w8380;
assign w8382 = w8372 & ~w8381;
assign w8383 = ~w8372 & w8381;
assign w8384 = ~w8382 & ~w8383;
assign w8385 = ~w2835 & w6304;
assign w8386 = ~w2546 & w6059;
assign w8387 = (w6061 & ~w2766) | (w6061 & w33755) | (~w2766 & w33755);
assign w8388 = ~w8385 & ~w8386;
assign w8389 = w8388 & w33756;
assign w8390 = (w8389 & ~w6733) | (w8389 & w31645) | (~w6733 & w31645);
assign w8391 = w6049 & w6054;
assign w8392 = (a_17 & ~w8388) | (a_17 & w33757) | (~w8388 & w33757);
assign w8393 = (~w8392 & ~w6733) | (~w8392 & w31646) | (~w6733 & w31646);
assign w8394 = ~w8390 & w8393;
assign w8395 = (a_20 & w8328) | (a_20 & w33758) | (w8328 & w33758);
assign w8396 = ~w8327 & w8395;
assign w8397 = w8327 & ~w8395;
assign w8398 = ~w8396 & ~w8397;
assign w8399 = w8394 & w8398;
assign w8400 = ~w8394 & ~w8398;
assign w8401 = ~w8399 & ~w8400;
assign w8402 = w6063 & w7970;
assign w8403 = (w6061 & ~w2479) | (w6061 & w33759) | (~w2479 & w33759);
assign w8404 = ~w2677 & w6304;
assign w8405 = (w6059 & ~w2600) | (w6059 & w33760) | (~w2600 & w33760);
assign w8406 = ~w8404 & w33761;
assign w8407 = ~w8402 & w8406;
assign w8408 = w6063 & ~w7287;
assign w8409 = (w6304 & ~w2479) | (w6304 & w31647) | (~w2479 & w31647);
assign w8410 = (w6061 & ~w2600) | (w6061 & w31648) | (~w2600 & w31648);
assign w8411 = ~w8409 & ~w8410;
assign w8412 = (w6054 & ~w2600) | (w6054 & w31649) | (~w2600 & w31649);
assign w8413 = a_17 & w8412;
assign w8414 = w8411 & ~w8413;
assign w8415 = ~w8408 & w8414;
assign w8416 = ~w8408 & w31650;
assign w8417 = (~w8332 & ~w8407) | (~w8332 & w31651) | (~w8407 & w31651);
assign w8418 = w6675 & w8391;
assign w8419 = w6050 & w6054;
assign w8420 = w6675 & w8419;
assign w8421 = ~w2677 & w6061;
assign w8422 = (w6059 & ~w2479) | (w6059 & w33762) | (~w2479 & w33762);
assign w8423 = ~w2546 & w6304;
assign w8424 = ~w8421 & ~w8422;
assign w8425 = w8424 & w33763;
assign w8426 = (~a_17 & ~w8424) | (~a_17 & w33764) | (~w8424 & w33764);
assign w8427 = ~w8425 & ~w8426;
assign w8428 = ~w8420 & w8427;
assign w8429 = ~w8418 & ~w8428;
assign w8430 = ~w8417 & w8429;
assign w8431 = (w6304 & ~w2766) | (w6304 & w33765) | (~w2766 & w33765);
assign w8432 = ~w2677 & w6059;
assign w8433 = ~w2546 & w6061;
assign w8434 = ~w8431 & ~w8432;
assign w8435 = ~w8433 & w8434;
assign w8436 = (w8435 & ~w7625) | (w8435 & w31652) | (~w7625 & w31652);
assign w8437 = w7286 & w8311;
assign w8438 = ~w8331 & w8333;
assign w8439 = ~w8437 & ~w8438;
assign w8440 = ~w8335 & w8439;
assign w8441 = (a_17 & w8335) | (a_17 & w31653) | (w8335 & w31653);
assign w8442 = ~w8335 & w31654;
assign w8443 = ~w8441 & ~w8442;
assign w8444 = w8436 & w8443;
assign w8445 = ~w8436 & ~w8443;
assign w8446 = ~w8444 & ~w8445;
assign w8447 = ~w8430 & w8446;
assign w8448 = ~w8440 & ~w8446;
assign w8449 = ~w8447 & ~w8448;
assign w8450 = w8401 & w8449;
assign w8451 = ~w8399 & ~w8450;
assign w8452 = ~w2917 & w6304;
assign w8453 = ~w2835 & w6061;
assign w8454 = (w6059 & ~w2766) | (w6059 & w33766) | (~w2766 & w33766);
assign w8455 = ~w8452 & ~w8453;
assign w8456 = ~w8454 & w8455;
assign w8457 = (~w6784 & w33767) | (~w6784 & w33768) | (w33767 & w33768);
assign w8458 = (w6784 & w33769) | (w6784 & w33770) | (w33769 & w33770);
assign w8459 = ~w8457 & ~w8458;
assign w8460 = w8327 & w31656;
assign w8461 = ~w8337 & ~w8460;
assign w8462 = w8349 & ~w8461;
assign w8463 = ~w8349 & w8461;
assign w8464 = ~w8462 & ~w8463;
assign w8465 = w8459 & ~w8464;
assign w8466 = ~w8459 & w8464;
assign w8467 = ~w8465 & ~w8466;
assign w8468 = w8350 & ~w8366;
assign w8469 = ~w8367 & ~w8468;
assign w8470 = w6063 & w6545;
assign w8471 = w6063 & ~w6544;
assign w8472 = ~w2920 & w31657;
assign w8473 = ~w2917 & w6061;
assign w8474 = ~w3007 & w6304;
assign w8475 = ~w2835 & w6059;
assign w8476 = ~w8473 & ~w8474;
assign w8477 = ~w8475 & w8476;
assign w8478 = ~w8472 & w8477;
assign w8479 = ~w8470 & w8478;
assign w8480 = a_17 & ~w8479;
assign w8481 = ~a_17 & w8479;
assign w8482 = ~w8480 & ~w8481;
assign w8483 = w8469 & ~w8482;
assign w8484 = w8467 & ~w8483;
assign w8485 = ~w8451 & w8484;
assign w8486 = ~w8469 & w8482;
assign w8487 = ~w8465 & ~w8486;
assign w8488 = ~w8483 & ~w8487;
assign w8489 = ~w8485 & ~w8488;
assign w8490 = w8384 & ~w8489;
assign w8491 = ~w8382 & ~w8490;
assign w8492 = ~w3326 & w6996;
assign w8493 = (w6998 & ~w3267) | (w6998 & w33771) | (~w3267 & w33771);
assign w8494 = ~w3196 & w6446;
assign w8495 = ~w8493 & ~w8494;
assign w8496 = ~w8492 & w8495;
assign w8497 = (w8496 & w5903) | (w8496 & w33772) | (w5903 & w33772);
assign w8498 = a_14 & ~w8497;
assign w8499 = (w5903 & w33773) | (w5903 & w33774) | (w33773 & w33774);
assign w8500 = ~w8498 & ~w8499;
assign w8501 = ~w8319 & ~w8370;
assign w8502 = ~w2835 & w5818;
assign w8503 = ~w2917 & w5816;
assign w8504 = (w5308 & ~w2766) | (w5308 & w33775) | (~w2766 & w33775);
assign w8505 = ~w8502 & ~w8503;
assign w8506 = ~w8504 & w8505;
assign w8507 = (~w6784 & w33776) | (~w6784 & w33777) | (w33776 & w33777);
assign w8508 = (w6784 & w33778) | (w6784 & w33779) | (w33778 & w33779);
assign w8509 = ~w8507 & ~w8508;
assign w8510 = w7976 & w31659;
assign w8511 = ~w7986 & ~w8510;
assign w8512 = w7996 & ~w8511;
assign w8513 = ~w7996 & w8511;
assign w8514 = ~w8512 & ~w8513;
assign w8515 = ~w8509 & w8514;
assign w8516 = w8509 & ~w8514;
assign w8517 = ~w8515 & ~w8516;
assign w8518 = ~w3007 & w6059;
assign w8519 = ~w3139 & w6304;
assign w8520 = ~w3049 & w6061;
assign w8521 = ~w8518 & ~w8519;
assign w8522 = ~w8520 & w8521;
assign w8523 = (w8522 & w6505) | (w8522 & w33780) | (w6505 & w33780);
assign w8524 = ~a_17 & w8523;
assign w8525 = (~w6505 & w33781) | (~w6505 & w33782) | (w33781 & w33782);
assign w8526 = ~w8524 & ~w8525;
assign w8527 = ~w8517 & ~w8526;
assign w8528 = w8501 & w8527;
assign w8529 = w8517 & ~w8526;
assign w8530 = ~w8501 & w8529;
assign w8531 = ~w8528 & ~w8530;
assign w8532 = w8517 & w8526;
assign w8533 = w8501 & w8532;
assign w8534 = ~w8517 & w8526;
assign w8535 = ~w8501 & w8534;
assign w8536 = ~w8533 & ~w8535;
assign w8537 = w8531 & w8536;
assign w8538 = w8500 & ~w8537;
assign w8539 = ~w8500 & w8537;
assign w8540 = ~w8538 & ~w8539;
assign w8541 = ~w8491 & w8540;
assign w8542 = w8491 & ~w8540;
assign w8543 = ~w8541 & ~w8542;
assign w8544 = ~w8401 & ~w8449;
assign w8545 = ~w8450 & ~w8544;
assign w8546 = ~w3049 & w6996;
assign w8547 = ~w3007 & w6998;
assign w8548 = ~w2917 & w6446;
assign w8549 = ~w8546 & ~w8547;
assign w8550 = ~w8548 & w8549;
assign w8551 = (w8550 & ~w6194) | (w8550 & w33783) | (~w6194 & w33783);
assign w8552 = a_14 & ~w8551;
assign w8553 = (~w6194 & w33784) | (~w6194 & w33785) | (w33784 & w33785);
assign w8554 = ~w8552 & ~w8553;
assign w8555 = w8545 & w8554;
assign w8556 = ~w8545 & ~w8554;
assign w8557 = ~w8555 & ~w8556;
assign w8558 = ~w2835 & w6996;
assign w8559 = ~w2546 & w6446;
assign w8560 = (w6998 & ~w2766) | (w6998 & w33786) | (~w2766 & w33786);
assign w8561 = ~w8558 & ~w8559;
assign w8562 = w8561 & w33787;
assign w8563 = (w8562 & ~w6733) | (w8562 & w31660) | (~w6733 & w31660);
assign w8564 = w6436 & w6441;
assign w8565 = (a_14 & ~w8561) | (a_14 & w33788) | (~w8561 & w33788);
assign w8566 = (~w8565 & ~w6733) | (~w8565 & w31661) | (~w6733 & w31661);
assign w8567 = ~w8563 & w8566;
assign w8568 = (a_17 & w8408) | (a_17 & w33789) | (w8408 & w33789);
assign w8569 = ~w8407 & w8568;
assign w8570 = w8407 & ~w8568;
assign w8571 = ~w8569 & ~w8570;
assign w8572 = w8567 & w8571;
assign w8573 = ~w8567 & ~w8571;
assign w8574 = ~w8572 & ~w8573;
assign w8575 = w6447 & w7970;
assign w8576 = (w6998 & ~w2479) | (w6998 & w33790) | (~w2479 & w33790);
assign w8577 = ~w2677 & w6996;
assign w8578 = (w6446 & ~w2600) | (w6446 & w33791) | (~w2600 & w33791);
assign w8579 = ~w8577 & w33792;
assign w8580 = ~w8575 & w8579;
assign w8581 = w6447 & ~w7287;
assign w8582 = (w6996 & ~w2479) | (w6996 & w31662) | (~w2479 & w31662);
assign w8583 = (w6998 & ~w2600) | (w6998 & w31663) | (~w2600 & w31663);
assign w8584 = ~w8582 & ~w8583;
assign w8585 = (w6441 & ~w2600) | (w6441 & w31664) | (~w2600 & w31664);
assign w8586 = a_14 & w8585;
assign w8587 = w8584 & ~w8586;
assign w8588 = ~w8581 & w8587;
assign w8589 = ~w8581 & w31665;
assign w8590 = (~w8412 & ~w8580) | (~w8412 & w31666) | (~w8580 & w31666);
assign w8591 = w6675 & w8564;
assign w8592 = w6437 & w6441;
assign w8593 = w6675 & w8592;
assign w8594 = ~w2677 & w6998;
assign w8595 = (w6446 & ~w2479) | (w6446 & w33793) | (~w2479 & w33793);
assign w8596 = ~w2546 & w6996;
assign w8597 = ~w8594 & ~w8595;
assign w8598 = w8597 & w33794;
assign w8599 = (~a_14 & ~w8597) | (~a_14 & w33795) | (~w8597 & w33795);
assign w8600 = ~w8598 & ~w8599;
assign w8601 = ~w8593 & w8600;
assign w8602 = ~w8591 & ~w8601;
assign w8603 = ~w8590 & w8602;
assign w8604 = (w6996 & ~w2766) | (w6996 & w33796) | (~w2766 & w33796);
assign w8605 = ~w2677 & w6446;
assign w8606 = ~w2546 & w6998;
assign w8607 = ~w8604 & ~w8605;
assign w8608 = ~w8606 & w8607;
assign w8609 = (w8608 & ~w7625) | (w8608 & w31667) | (~w7625 & w31667);
assign w8610 = w7286 & w8391;
assign w8611 = ~w8411 & w8413;
assign w8612 = ~w8610 & ~w8611;
assign w8613 = ~w8415 & w8612;
assign w8614 = (a_14 & w8415) | (a_14 & w31668) | (w8415 & w31668);
assign w8615 = ~w8415 & w31669;
assign w8616 = ~w8614 & ~w8615;
assign w8617 = w8609 & w8616;
assign w8618 = ~w8609 & ~w8616;
assign w8619 = ~w8617 & ~w8618;
assign w8620 = ~w8603 & w8619;
assign w8621 = ~w8613 & ~w8619;
assign w8622 = ~w8620 & ~w8621;
assign w8623 = w8574 & w8622;
assign w8624 = ~w8572 & ~w8623;
assign w8625 = w8430 & ~w8446;
assign w8626 = ~w8447 & ~w8625;
assign w8627 = w6447 & w6545;
assign w8628 = w6447 & ~w6544;
assign w8629 = ~w2920 & w31670;
assign w8630 = ~w3007 & w6996;
assign w8631 = ~w2917 & w6998;
assign w8632 = ~w2835 & w6446;
assign w8633 = ~w8630 & ~w8631;
assign w8634 = ~w8632 & w8633;
assign w8635 = ~w8629 & w8634;
assign w8636 = ~w8627 & w8635;
assign w8637 = a_14 & ~w8636;
assign w8638 = ~a_14 & w8636;
assign w8639 = ~w8637 & ~w8638;
assign w8640 = w8626 & ~w8639;
assign w8641 = ~w2835 & w6998;
assign w8642 = ~w2917 & w6996;
assign w8643 = (w6446 & ~w2766) | (w6446 & w33797) | (~w2766 & w33797);
assign w8644 = ~w8641 & ~w8642;
assign w8645 = ~w8643 & w8644;
assign w8646 = (~w6784 & w33798) | (~w6784 & w33799) | (w33798 & w33799);
assign w8647 = (w6784 & w33800) | (w6784 & w33801) | (w33800 & w33801);
assign w8648 = ~w8646 & ~w8647;
assign w8649 = w8407 & w31672;
assign w8650 = ~w8417 & ~w8649;
assign w8651 = w8429 & ~w8650;
assign w8652 = ~w8429 & w8650;
assign w8653 = ~w8651 & ~w8652;
assign w8654 = w8648 & ~w8653;
assign w8655 = ~w8648 & w8653;
assign w8656 = ~w8654 & ~w8655;
assign w8657 = ~w8640 & w8656;
assign w8658 = ~w8624 & w8657;
assign w8659 = ~w8626 & w8639;
assign w8660 = ~w8640 & w8654;
assign w8661 = ~w8659 & ~w8660;
assign w8662 = ~w8658 & w8661;
assign w8663 = w8557 & ~w8662;
assign w8664 = ~w3007 & w6446;
assign w8665 = ~w3139 & w6996;
assign w8666 = ~w3049 & w6998;
assign w8667 = ~w8664 & ~w8665;
assign w8668 = ~w8666 & w8667;
assign w8669 = (w8668 & w6505) | (w8668 & w33802) | (w6505 & w33802);
assign w8670 = a_14 & ~w8669;
assign w8671 = (w6505 & w33803) | (w6505 & w33804) | (w33803 & w33804);
assign w8672 = ~w8670 & ~w8671;
assign w8673 = w8467 & w8672;
assign w8674 = w8451 & w8673;
assign w8675 = ~w8467 & w8672;
assign w8676 = ~w8451 & w8675;
assign w8677 = ~w8674 & ~w8676;
assign w8678 = ~w8555 & w8677;
assign w8679 = ~w8663 & w8678;
assign w8680 = ~w8467 & ~w8672;
assign w8681 = w8451 & w8680;
assign w8682 = w8467 & ~w8672;
assign w8683 = ~w8451 & w8682;
assign w8684 = ~w8681 & ~w8683;
assign w8685 = ~w8399 & ~w8465;
assign w8686 = ~w8450 & w8685;
assign w8687 = ~w8466 & ~w8686;
assign w8688 = w6491 & w8564;
assign w8689 = ~w6216 & w33805;
assign w8690 = (w8689 & w3058) | (w8689 & w33806) | (w3058 & w33806);
assign w8691 = ~w3196 & w6996;
assign w8692 = ~w3049 & w6446;
assign w8693 = ~w3139 & w6998;
assign w8694 = ~w8691 & ~w8692;
assign w8695 = (~a_14 & ~w8694) | (~a_14 & w33807) | (~w8694 & w33807);
assign w8696 = w8694 & w33808;
assign w8697 = ~w8695 & ~w8696;
assign w8698 = (w8697 & ~w8690) | (w8697 & w31673) | (~w8690 & w31673);
assign w8699 = ~w8688 & ~w8698;
assign w8700 = w8482 & ~w8699;
assign w8701 = ~w8482 & w8699;
assign w8702 = ~w8700 & ~w8701;
assign w8703 = w8469 & ~w8702;
assign w8704 = ~w8469 & w8702;
assign w8705 = ~w8703 & ~w8704;
assign w8706 = w8687 & w8705;
assign w8707 = ~w8687 & ~w8705;
assign w8708 = ~w8706 & ~w8707;
assign w8709 = w8684 & ~w8708;
assign w8710 = ~w8679 & w8709;
assign w8711 = w8699 & w8708;
assign w8712 = ~w8710 & ~w8711;
assign w8713 = ~w8384 & w8489;
assign w8714 = ~w8490 & ~w8713;
assign w8715 = (w6996 & ~w3267) | (w6996 & w33809) | (~w3267 & w33809);
assign w8716 = ~w3196 & w6998;
assign w8717 = ~w3139 & w6446;
assign w8718 = w6222 & w33810;
assign w8719 = ~w8715 & ~w8716;
assign w8720 = ~w8717 & w8719;
assign w8721 = (a_14 & w8718) | (a_14 & w33811) | (w8718 & w33811);
assign w8722 = ~w8718 & w33812;
assign w8723 = ~w8721 & ~w8722;
assign w8724 = w8714 & w8723;
assign w8725 = w8712 & ~w8724;
assign w8726 = ~w8714 & ~w8723;
assign w8727 = (~w8726 & ~w8712) | (~w8726 & w33813) | (~w8712 & w33813);
assign w8728 = ~w8543 & w8727;
assign w8729 = ~w8382 & w8536;
assign w8730 = ~w8490 & w8729;
assign w8731 = ~w8319 & ~w8516;
assign w8732 = ~w8370 & w8731;
assign w8733 = ~w8515 & ~w8732;
assign w8734 = ~w7997 & ~w8012;
assign w8735 = ~w8013 & ~w8734;
assign w8736 = w5309 & w6545;
assign w8737 = w5309 & ~w6544;
assign w8738 = ~w2920 & w31674;
assign w8739 = ~w3007 & w5816;
assign w8740 = ~w2917 & w5818;
assign w8741 = ~w2835 & w5308;
assign w8742 = ~w8739 & ~w8740;
assign w8743 = ~w8741 & w8742;
assign w8744 = ~w8738 & w8743;
assign w8745 = ~w8736 & w8744;
assign w8746 = a_20 & ~w8745;
assign w8747 = ~a_20 & w8745;
assign w8748 = ~w8746 & ~w8747;
assign w8749 = w6491 & w8391;
assign w8750 = ~w6216 & w33814;
assign w8751 = (w8750 & w3058) | (w8750 & w33815) | (w3058 & w33815);
assign w8752 = ~w3196 & w6304;
assign w8753 = ~w3049 & w6059;
assign w8754 = ~w3139 & w6061;
assign w8755 = ~w8752 & ~w8753;
assign w8756 = (~a_17 & ~w8755) | (~a_17 & w33816) | (~w8755 & w33816);
assign w8757 = w8755 & w33817;
assign w8758 = ~w8756 & ~w8757;
assign w8759 = (w8758 & ~w8751) | (w8758 & w31675) | (~w8751 & w31675);
assign w8760 = ~w8749 & ~w8759;
assign w8761 = w8748 & ~w8760;
assign w8762 = ~w8748 & w8760;
assign w8763 = ~w8761 & ~w8762;
assign w8764 = w8735 & ~w8763;
assign w8765 = ~w8735 & w8763;
assign w8766 = ~w8764 & ~w8765;
assign w8767 = w8733 & w8766;
assign w8768 = ~w8733 & ~w8766;
assign w8769 = ~w8767 & ~w8768;
assign w8770 = w8531 & w8769;
assign w8771 = ~w8730 & w8770;
assign w8772 = w8760 & ~w8769;
assign w8773 = ~w8771 & ~w8772;
assign w8774 = ~w3475 & w6998;
assign w8775 = ~w3403 & w6996;
assign w8776 = ~w3326 & w6446;
assign w8777 = ~w8774 & ~w8775;
assign w8778 = ~w8776 & w8777;
assign w8779 = (w8778 & ~w5923) | (w8778 & w33818) | (~w5923 & w33818);
assign w8780 = a_14 & w8779;
assign w8781 = (w5923 & w33819) | (w5923 & w33820) | (w33819 & w33820);
assign w8782 = ~w8780 & ~w8781;
assign w8783 = ~w8735 & ~w8748;
assign w8784 = ~w8515 & ~w8783;
assign w8785 = ~w8732 & w8784;
assign w8786 = w8735 & w8748;
assign w8787 = ~w8785 & ~w8786;
assign w8788 = ~w8013 & ~w8018;
assign w8789 = ~w7968 & ~w8014;
assign w8790 = w6194 & w8311;
assign w8791 = ~w3007 & w5818;
assign w8792 = ~w2917 & w5308;
assign w8793 = ~w3049 & w5816;
assign w8794 = ~w8791 & ~w8792;
assign w8795 = (~a_20 & ~w8794) | (~a_20 & w33821) | (~w8794 & w33821);
assign w8796 = w8794 & w33822;
assign w8797 = ~w8795 & ~w8796;
assign w8798 = (w8797 & ~w6194) | (w8797 & w31676) | (~w6194 & w31676);
assign w8799 = ~w8790 & ~w8798;
assign w8800 = w8789 & w8799;
assign w8801 = w8788 & w8800;
assign w8802 = ~w8789 & w8799;
assign w8803 = ~w8788 & w8802;
assign w8804 = ~w8801 & ~w8803;
assign w8805 = ~w8789 & ~w8799;
assign w8806 = w8788 & w8805;
assign w8807 = w8789 & ~w8799;
assign w8808 = ~w8788 & w8807;
assign w8809 = ~w8806 & ~w8808;
assign w8810 = w8804 & w8809;
assign w8811 = w6222 & w33823;
assign w8812 = (w6304 & ~w3267) | (w6304 & w33824) | (~w3267 & w33824);
assign w8813 = ~w3139 & w6059;
assign w8814 = ~w3196 & w6061;
assign w8815 = ~w8812 & ~w8813;
assign w8816 = (a_17 & ~w8815) | (a_17 & w33825) | (~w8815 & w33825);
assign w8817 = w6222 & w33826;
assign w8818 = w8815 & w33827;
assign w8819 = ~w8817 & w8818;
assign w8820 = ~w8811 & ~w8816;
assign w8821 = ~w8819 & w8820;
assign w8822 = ~w8810 & w8821;
assign w8823 = w8810 & ~w8821;
assign w8824 = ~w8822 & ~w8823;
assign w8825 = w8787 & ~w8824;
assign w8826 = ~w8787 & w8824;
assign w8827 = ~w8825 & ~w8826;
assign w8828 = ~w8782 & ~w8827;
assign w8829 = w8773 & w8828;
assign w8830 = ~w8782 & w8827;
assign w8831 = ~w8773 & w8830;
assign w8832 = ~w8829 & ~w8831;
assign w8833 = (w8500 & ~w8491) | (w8500 & w33828) | (~w8491 & w33828);
assign w8834 = ~w8541 & w8833;
assign w8835 = w8531 & ~w8730;
assign w8836 = (~w8769 & w8730) | (~w8769 & w33829) | (w8730 & w33829);
assign w8837 = ~w3475 & w6996;
assign w8838 = (w6446 & ~w3267) | (w6446 & w33830) | (~w3267 & w33830);
assign w8839 = ~w3326 & w6998;
assign w8840 = ~w8837 & ~w8838;
assign w8841 = ~w8839 & w8840;
assign w8842 = (w8841 & ~w6108) | (w8841 & w33831) | (~w6108 & w33831);
assign w8843 = a_14 & ~w8842;
assign w8844 = (~w6108 & w33832) | (~w6108 & w33833) | (w33832 & w33833);
assign w8845 = ~w8843 & ~w8844;
assign w8846 = ~w8771 & w8845;
assign w8847 = ~w8836 & w8846;
assign w8848 = ~w8834 & ~w8847;
assign w8849 = w8832 & w33834;
assign w8850 = w8771 & ~w8845;
assign w8851 = ~w8769 & ~w8845;
assign w8852 = ~w8835 & w8851;
assign w8853 = ~w8850 & ~w8852;
assign w8854 = w8782 & w8827;
assign w8855 = w8773 & w8854;
assign w8856 = w8782 & ~w8827;
assign w8857 = ~w8773 & w8856;
assign w8858 = ~w8855 & ~w8857;
assign w8859 = w8853 & w8858;
assign w8860 = w8832 & ~w8859;
assign w8861 = ~w8849 & ~w8860;
assign w8862 = ~w2306 & w7192;
assign w8863 = ~w3615 & w7511;
assign w8864 = ~w2393 & w7489;
assign w8865 = ~w8862 & ~w8863;
assign w8866 = ~w8864 & w8865;
assign w8867 = (w8866 & ~w5463) | (w8866 & w33835) | (~w5463 & w33835);
assign w8868 = a_11 & ~w8867;
assign w8869 = (~w5463 & w33836) | (~w5463 & w33837) | (w33836 & w33837);
assign w8870 = ~w8868 & ~w8869;
assign w8871 = ~w8787 & w8822;
assign w8872 = w8810 & w8821;
assign w8873 = w8787 & w8872;
assign w8874 = ~w8871 & ~w8873;
assign w8875 = w8827 & w8874;
assign w8876 = ~w8772 & w8874;
assign w8877 = ~w8771 & w8876;
assign w8878 = ~w8875 & ~w8877;
assign w8879 = ~w8786 & w8804;
assign w8880 = (w8809 & ~w8879) | (w8809 & w31677) | (~w8879 & w31677);
assign w8881 = ~w3058 & w33838;
assign w8882 = w5309 & ~w6502;
assign w8883 = ~w3007 & w5308;
assign w8884 = ~w3139 & w5816;
assign w8885 = ~w3049 & w5818;
assign w8886 = ~w8883 & ~w8884;
assign w8887 = ~w8885 & w8886;
assign w8888 = (~w3058 & w33839) | (~w3058 & w33840) | (w33839 & w33840);
assign w8889 = ~w8881 & w8888;
assign w8890 = a_20 & ~w8889;
assign w8891 = ~a_20 & w8889;
assign w8892 = ~w8890 & ~w8891;
assign w8893 = w8040 & ~w8892;
assign w8894 = w8020 & w8893;
assign w8895 = ~w8040 & ~w8892;
assign w8896 = ~w8020 & w8895;
assign w8897 = ~w8894 & ~w8896;
assign w8898 = ~w8040 & w8892;
assign w8899 = w8020 & w8898;
assign w8900 = w8040 & w8892;
assign w8901 = ~w8020 & w8900;
assign w8902 = ~w8899 & ~w8901;
assign w8903 = w8897 & w8902;
assign w8904 = ~w3326 & w6304;
assign w8905 = ~w3196 & w6059;
assign w8906 = (w6061 & ~w3267) | (w6061 & w33841) | (~w3267 & w33841);
assign w8907 = ~w8905 & ~w8906;
assign w8908 = ~w8904 & w8907;
assign w8909 = (w8908 & w5903) | (w8908 & w33842) | (w5903 & w33842);
assign w8910 = a_17 & w8909;
assign w8911 = (~w5903 & w33843) | (~w5903 & w33844) | (w33843 & w33844);
assign w8912 = ~w8910 & ~w8911;
assign w8913 = w8903 & ~w8912;
assign w8914 = ~w8903 & w8912;
assign w8915 = ~w8913 & ~w8914;
assign w8916 = w8880 & w8915;
assign w8917 = ~w8880 & ~w8915;
assign w8918 = ~w8916 & ~w8917;
assign w8919 = ~w3403 & w6998;
assign w8920 = (w6996 & ~w3538) | (w6996 & w33845) | (~w3538 & w33845);
assign w8921 = ~w3475 & w6446;
assign w8922 = ~w8919 & ~w8920;
assign w8923 = ~w8921 & w8922;
assign w8924 = (w8923 & ~w5652) | (w8923 & w33846) | (~w5652 & w33846);
assign w8925 = a_14 & ~w8924;
assign w8926 = (~w5652 & w33847) | (~w5652 & w33848) | (w33847 & w33848);
assign w8927 = ~w8925 & ~w8926;
assign w8928 = w8918 & ~w8927;
assign w8929 = ~w8918 & w8927;
assign w8930 = ~w8928 & ~w8929;
assign w8931 = w8878 & w8930;
assign w8932 = ~w8878 & ~w8930;
assign w8933 = ~w8931 & ~w8932;
assign w8934 = w8870 & w8933;
assign w8935 = ~w8870 & ~w8933;
assign w8936 = ~w8934 & ~w8935;
assign w8937 = w8861 & w8936;
assign w8938 = ~w8861 & ~w8936;
assign w8939 = ~w8937 & ~w8938;
assign w8940 = ~w8848 & w8853;
assign w8941 = ~w8543 & w8853;
assign w8942 = w8727 & w8941;
assign w8943 = ~w8940 & ~w8942;
assign w8944 = w8832 & w8858;
assign w8945 = ~w2306 & w7489;
assign w8946 = (w7192 & ~w3538) | (w7192 & w33849) | (~w3538 & w33849);
assign w8947 = ~w2393 & w7511;
assign w8948 = ~w8945 & ~w8946;
assign w8949 = ~w8947 & w8948;
assign w8950 = (w8949 & ~w5483) | (w8949 & w33850) | (~w5483 & w33850);
assign w8951 = a_11 & w8950;
assign w8952 = (w5483 & w33851) | (w5483 & w33852) | (w33851 & w33852);
assign w8953 = ~w8951 & ~w8952;
assign w8954 = w8944 & w8953;
assign w8955 = ~w8943 & ~w8954;
assign w8956 = ~w8944 & w8953;
assign w8957 = w8943 & ~w8956;
assign w8958 = ~w8955 & ~w8957;
assign w8959 = w8491 & w33853;
assign w8960 = ~w8491 & w8539;
assign w8961 = ~w8726 & ~w8960;
assign w8962 = ~w8959 & w8961;
assign w8963 = ~w8725 & w8962;
assign w8964 = ~w8834 & ~w8963;
assign w8965 = ~w8847 & w8853;
assign w8966 = ~w3403 & w7192;
assign w8967 = ~w2306 & w7511;
assign w8968 = (w7489 & ~w3538) | (w7489 & w33854) | (~w3538 & w33854);
assign w8969 = ~w8967 & ~w8968;
assign w8970 = ~w8966 & w8969;
assign w8971 = (w8970 & ~w5706) | (w8970 & w33855) | (~w5706 & w33855);
assign w8972 = a_11 & w8971;
assign w8973 = (w5706 & w33856) | (w5706 & w33857) | (w33856 & w33857);
assign w8974 = ~w8972 & ~w8973;
assign w8975 = ~w8965 & w8974;
assign w8976 = w8965 & ~w8974;
assign w8977 = ~w8975 & ~w8976;
assign w8978 = w8964 & w8977;
assign w8979 = (~w8974 & w8964) | (~w8974 & w33858) | (w8964 & w33858);
assign w8980 = ~w8978 & w8979;
assign w8981 = ~w8944 & ~w8953;
assign w8982 = ~w8943 & ~w8981;
assign w8983 = w8944 & ~w8953;
assign w8984 = w8943 & ~w8983;
assign w8985 = ~w8982 & ~w8984;
assign w8986 = ~w8980 & ~w8985;
assign w8987 = ~w8958 & ~w8986;
assign w8988 = ~w3326 & w7489;
assign w8989 = (w7192 & ~w3267) | (w7192 & w33859) | (~w3267 & w33859);
assign w8990 = ~w3475 & w7511;
assign w8991 = ~w8988 & ~w8989;
assign w8992 = ~w8990 & w8991;
assign w8993 = (w8992 & ~w6108) | (w8992 & w33860) | (~w6108 & w33860);
assign w8994 = a_11 & ~w8993;
assign w8995 = (~w6108 & w33861) | (~w6108 & w33862) | (w33861 & w33862);
assign w8996 = ~w8994 & ~w8995;
assign w8997 = w8710 & ~w8996;
assign w8998 = ~w8679 & w8684;
assign w8999 = w8708 & ~w8996;
assign w9000 = ~w8998 & w8999;
assign w9001 = ~w8997 & ~w9000;
assign w9002 = (w8708 & w8679) | (w8708 & w33863) | (w8679 & w33863);
assign w9003 = ~w8710 & w8996;
assign w9004 = ~w9002 & w9003;
assign w9005 = ~w3326 & w7511;
assign w9006 = ~w3196 & w7192;
assign w9007 = (w7489 & ~w3267) | (w7489 & w33864) | (~w3267 & w33864);
assign w9008 = ~w9006 & ~w9007;
assign w9009 = ~w9005 & w9008;
assign w9010 = (w9009 & w5903) | (w9009 & w33865) | (w5903 & w33865);
assign w9011 = a_11 & w9010;
assign w9012 = (~w5903 & w33866) | (~w5903 & w33867) | (w33866 & w33867);
assign w9013 = ~w9011 & ~w9012;
assign w9014 = w8677 & w8684;
assign w9015 = ~w8555 & ~w8663;
assign w9016 = ~w9014 & ~w9015;
assign w9017 = w9014 & w9015;
assign w9018 = ~w9016 & ~w9017;
assign w9019 = ~w9013 & ~w9018;
assign w9020 = ~w9004 & ~w9019;
assign w9021 = w9001 & ~w9020;
assign w9022 = ~w9013 & w9014;
assign w9023 = w9013 & ~w9014;
assign w9024 = ~w9022 & ~w9023;
assign w9025 = w9015 & w9024;
assign w9026 = ~w9015 & ~w9024;
assign w9027 = ~w9025 & ~w9026;
assign w9028 = ~w8557 & w8662;
assign w9029 = ~w8663 & ~w9028;
assign w9030 = ~w3139 & w7192;
assign w9031 = (w7511 & ~w3267) | (w7511 & w33868) | (~w3267 & w33868);
assign w9032 = ~w3196 & w7489;
assign w9033 = w6222 & w33869;
assign w9034 = ~w9030 & ~w9031;
assign w9035 = ~w9032 & w9034;
assign w9036 = (a_11 & w9033) | (a_11 & w33870) | (w9033 & w33870);
assign w9037 = ~w9033 & w33871;
assign w9038 = ~w9036 & ~w9037;
assign w9039 = w9029 & w9038;
assign w9040 = ~w9029 & ~w9038;
assign w9041 = ~w8574 & ~w8622;
assign w9042 = ~w8623 & ~w9041;
assign w9043 = ~w2917 & w7192;
assign w9044 = ~w3049 & w7511;
assign w9045 = ~w3007 & w7489;
assign w9046 = ~w9043 & ~w9044;
assign w9047 = ~w9045 & w9046;
assign w9048 = (w9047 & ~w6194) | (w9047 & w33872) | (~w6194 & w33872);
assign w9049 = a_11 & ~w9048;
assign w9050 = (~w6194 & w33873) | (~w6194 & w33874) | (w33873 & w33874);
assign w9051 = ~w9049 & ~w9050;
assign w9052 = w9042 & w9051;
assign w9053 = ~w9042 & ~w9051;
assign w9054 = ~w9052 & ~w9053;
assign w9055 = ~w2835 & w7511;
assign w9056 = ~w2546 & w7192;
assign w9057 = (w7489 & ~w2766) | (w7489 & w33875) | (~w2766 & w33875);
assign w9058 = ~w9055 & ~w9056;
assign w9059 = w9058 & w33876;
assign w9060 = (w9059 & ~w6733) | (w9059 & w31679) | (~w6733 & w31679);
assign w9061 = w7182 & w7187;
assign w9062 = (a_11 & ~w9058) | (a_11 & w33877) | (~w9058 & w33877);
assign w9063 = (~w9062 & ~w6733) | (~w9062 & w31680) | (~w6733 & w31680);
assign w9064 = ~w9060 & w9063;
assign w9065 = (a_14 & w8581) | (a_14 & w33878) | (w8581 & w33878);
assign w9066 = ~w8580 & w9065;
assign w9067 = w8580 & ~w9065;
assign w9068 = ~w9066 & ~w9067;
assign w9069 = w9064 & w9068;
assign w9070 = ~w9064 & ~w9068;
assign w9071 = ~w9069 & ~w9070;
assign w9072 = w7193 & w7970;
assign w9073 = (w7489 & ~w2479) | (w7489 & w33879) | (~w2479 & w33879);
assign w9074 = ~w2677 & w7511;
assign w9075 = (w7192 & ~w2600) | (w7192 & w33880) | (~w2600 & w33880);
assign w9076 = ~w9074 & w33881;
assign w9077 = ~w9072 & w9076;
assign w9078 = w7193 & ~w7287;
assign w9079 = (w7511 & ~w2479) | (w7511 & w31681) | (~w2479 & w31681);
assign w9080 = (w7489 & ~w2600) | (w7489 & w31682) | (~w2600 & w31682);
assign w9081 = ~w9079 & ~w9080;
assign w9082 = (w7187 & ~w2600) | (w7187 & w31683) | (~w2600 & w31683);
assign w9083 = a_11 & w9082;
assign w9084 = w9081 & ~w9083;
assign w9085 = ~w9078 & w9084;
assign w9086 = ~w9078 & w31684;
assign w9087 = (~w8585 & ~w9077) | (~w8585 & w31685) | (~w9077 & w31685);
assign w9088 = w6675 & w9061;
assign w9089 = w7183 & w7187;
assign w9090 = w6675 & w9089;
assign w9091 = ~w2546 & w7511;
assign w9092 = (w7192 & ~w2479) | (w7192 & w33882) | (~w2479 & w33882);
assign w9093 = ~w2677 & w7489;
assign w9094 = ~w9091 & ~w9092;
assign w9095 = w9094 & w33883;
assign w9096 = (~a_11 & ~w9094) | (~a_11 & w33884) | (~w9094 & w33884);
assign w9097 = ~w9095 & ~w9096;
assign w9098 = ~w9090 & w9097;
assign w9099 = ~w9088 & ~w9098;
assign w9100 = ~w9087 & w9099;
assign w9101 = (w7511 & ~w2766) | (w7511 & w33885) | (~w2766 & w33885);
assign w9102 = ~w2677 & w7192;
assign w9103 = ~w2546 & w7489;
assign w9104 = ~w9101 & ~w9102;
assign w9105 = ~w9103 & w9104;
assign w9106 = (w9105 & ~w7625) | (w9105 & w31686) | (~w7625 & w31686);
assign w9107 = w7286 & w8564;
assign w9108 = ~w8584 & w8586;
assign w9109 = ~w9107 & ~w9108;
assign w9110 = ~w8588 & w9109;
assign w9111 = (a_11 & w8588) | (a_11 & w31687) | (w8588 & w31687);
assign w9112 = ~w8588 & w31688;
assign w9113 = ~w9111 & ~w9112;
assign w9114 = w9106 & w9113;
assign w9115 = ~w9106 & ~w9113;
assign w9116 = ~w9114 & ~w9115;
assign w9117 = ~w9100 & w9116;
assign w9118 = ~w9110 & ~w9116;
assign w9119 = ~w9117 & ~w9118;
assign w9120 = w9071 & w9119;
assign w9121 = ~w9069 & ~w9120;
assign w9122 = w8603 & ~w8619;
assign w9123 = ~w8620 & ~w9122;
assign w9124 = w6545 & w7193;
assign w9125 = ~w6544 & w7193;
assign w9126 = ~w2920 & w31689;
assign w9127 = ~w3007 & w7511;
assign w9128 = ~w2917 & w7489;
assign w9129 = ~w2835 & w7192;
assign w9130 = ~w9127 & ~w9128;
assign w9131 = ~w9129 & w9130;
assign w9132 = ~w9126 & w9131;
assign w9133 = ~w9124 & w9132;
assign w9134 = a_11 & ~w9133;
assign w9135 = ~a_11 & w9133;
assign w9136 = ~w9134 & ~w9135;
assign w9137 = w9123 & ~w9136;
assign w9138 = ~w2835 & w7489;
assign w9139 = ~w2917 & w7511;
assign w9140 = (w7192 & ~w2766) | (w7192 & w33886) | (~w2766 & w33886);
assign w9141 = ~w9138 & ~w9139;
assign w9142 = ~w9140 & w9141;
assign w9143 = (~w6784 & w33887) | (~w6784 & w33888) | (w33887 & w33888);
assign w9144 = (w6784 & w33889) | (w6784 & w33890) | (w33889 & w33890);
assign w9145 = ~w9143 & ~w9144;
assign w9146 = w8580 & w31691;
assign w9147 = ~w8590 & ~w9146;
assign w9148 = w8602 & ~w9147;
assign w9149 = ~w8602 & w9147;
assign w9150 = ~w9148 & ~w9149;
assign w9151 = w9145 & ~w9150;
assign w9152 = ~w9145 & w9150;
assign w9153 = ~w9151 & ~w9152;
assign w9154 = ~w9137 & w9153;
assign w9155 = ~w9121 & w9154;
assign w9156 = ~w9123 & w9136;
assign w9157 = ~w9137 & w9151;
assign w9158 = ~w9156 & ~w9157;
assign w9159 = ~w9155 & w9158;
assign w9160 = w9054 & ~w9159;
assign w9161 = ~w3007 & w7192;
assign w9162 = ~w3139 & w7511;
assign w9163 = ~w3049 & w7489;
assign w9164 = ~w9161 & ~w9162;
assign w9165 = ~w9163 & w9164;
assign w9166 = (w9165 & w6505) | (w9165 & w33891) | (w6505 & w33891);
assign w9167 = a_11 & ~w9166;
assign w9168 = (w6505 & w33892) | (w6505 & w33893) | (w33892 & w33893);
assign w9169 = ~w9167 & ~w9168;
assign w9170 = ~w8656 & w9169;
assign w9171 = ~w8624 & w9170;
assign w9172 = w8656 & w9169;
assign w9173 = w8624 & w9172;
assign w9174 = ~w9171 & ~w9173;
assign w9175 = ~w9052 & w9174;
assign w9176 = ~w9160 & w9175;
assign w9177 = ~w8656 & ~w9169;
assign w9178 = w8624 & w9177;
assign w9179 = w8656 & ~w9169;
assign w9180 = ~w8624 & w9179;
assign w9181 = ~w9178 & ~w9180;
assign w9182 = ~w8572 & ~w8654;
assign w9183 = ~w8623 & w9182;
assign w9184 = ~w8655 & ~w9183;
assign w9185 = w6491 & w9061;
assign w9186 = ~w6216 & w33894;
assign w9187 = (w9186 & w3058) | (w9186 & w33895) | (w3058 & w33895);
assign w9188 = ~w3196 & w7511;
assign w9189 = ~w3049 & w7192;
assign w9190 = ~w3139 & w7489;
assign w9191 = ~w9188 & ~w9189;
assign w9192 = (~a_11 & ~w9191) | (~a_11 & w33896) | (~w9191 & w33896);
assign w9193 = w9191 & w33897;
assign w9194 = ~w9192 & ~w9193;
assign w9195 = (w9194 & ~w9187) | (w9194 & w31692) | (~w9187 & w31692);
assign w9196 = ~w9185 & ~w9195;
assign w9197 = w8639 & ~w9196;
assign w9198 = ~w8639 & w9196;
assign w9199 = ~w9197 & ~w9198;
assign w9200 = w8626 & ~w9199;
assign w9201 = ~w8626 & w9199;
assign w9202 = ~w9200 & ~w9201;
assign w9203 = w9184 & w9202;
assign w9204 = ~w9184 & ~w9202;
assign w9205 = ~w9203 & ~w9204;
assign w9206 = w9181 & ~w9205;
assign w9207 = ~w9176 & w9206;
assign w9208 = w9196 & w9205;
assign w9209 = ~w9207 & ~w9208;
assign w9210 = (~w9039 & w9209) | (~w9039 & w33898) | (w9209 & w33898);
assign w9211 = w9001 & ~w9027;
assign w9212 = ~w9210 & w9211;
assign w9213 = ~w9021 & ~w9212;
assign w9214 = ~w3403 & w7511;
assign w9215 = ~w3475 & w7489;
assign w9216 = ~w3326 & w7192;
assign w9217 = ~w9214 & ~w9215;
assign w9218 = ~w9216 & w9217;
assign w9219 = (w9218 & ~w5923) | (w9218 & w33899) | (~w5923 & w33899);
assign w9220 = a_11 & w9219;
assign w9221 = (w5923 & w33900) | (w5923 & w33901) | (w33900 & w33901);
assign w9222 = ~w9220 & ~w9221;
assign w9223 = w8723 & ~w9222;
assign w9224 = ~w8723 & w9222;
assign w9225 = ~w9223 & ~w9224;
assign w9226 = w8714 & ~w9225;
assign w9227 = ~w8714 & w9225;
assign w9228 = ~w9226 & ~w9227;
assign w9229 = w8712 & w9228;
assign w9230 = ~w8712 & ~w9228;
assign w9231 = ~w9229 & ~w9230;
assign w9232 = ~w9213 & w9231;
assign w9233 = ~w9222 & ~w9231;
assign w9234 = ~w3403 & w7489;
assign w9235 = (w7511 & ~w3538) | (w7511 & w33902) | (~w3538 & w33902);
assign w9236 = ~w3475 & w7192;
assign w9237 = ~w9234 & ~w9235;
assign w9238 = ~w9236 & w9237;
assign w9239 = (w9238 & ~w5652) | (w9238 & w33903) | (~w5652 & w33903);
assign w9240 = a_11 & ~w9239;
assign w9241 = (~w5652 & w33904) | (~w5652 & w33905) | (w33904 & w33905);
assign w9242 = ~w9240 & ~w9241;
assign w9243 = ~w8543 & w9242;
assign w9244 = ~w8727 & w9243;
assign w9245 = w8543 & w9242;
assign w9246 = w8727 & w9245;
assign w9247 = ~w9244 & ~w9246;
assign w9248 = ~w9233 & w9247;
assign w9249 = ~w9232 & w9248;
assign w9250 = w8543 & ~w9242;
assign w9251 = ~w8727 & w9250;
assign w9252 = ~w8543 & ~w9242;
assign w9253 = w8727 & w9252;
assign w9254 = ~w9251 & ~w9253;
assign w9255 = ~w9249 & w9254;
assign w9256 = ~w8964 & ~w8977;
assign w9257 = ~w8978 & ~w9256;
assign w9258 = ~w8958 & ~w9257;
assign w9259 = w9255 & w9258;
assign w9260 = ~w8987 & ~w9259;
assign w9261 = ~w8939 & ~w9260;
assign w9262 = w8861 & ~w8933;
assign w9263 = (w8870 & ~w8861) | (w8870 & w8934) | (~w8861 & w8934);
assign w9264 = ~w8938 & w9263;
assign w9265 = (~w9264 & w9260) | (~w9264 & w31693) | (w9260 & w31693);
assign w9266 = w8927 & w8933;
assign w9267 = ~w9262 & ~w9266;
assign w9268 = w8804 & w8902;
assign w9269 = ~w8880 & w9268;
assign w9270 = ~w8038 & ~w8041;
assign w9271 = w6491 & w8311;
assign w9272 = ~w6216 & w33906;
assign w9273 = (w9272 & w3058) | (w9272 & w33907) | (w3058 & w33907);
assign w9274 = ~w3139 & w5818;
assign w9275 = ~w3049 & w5308;
assign w9276 = ~w3196 & w5816;
assign w9277 = ~w9274 & ~w9275;
assign w9278 = (~a_20 & ~w9277) | (~a_20 & w33908) | (~w9277 & w33908);
assign w9279 = w9277 & w33909;
assign w9280 = ~w9278 & ~w9279;
assign w9281 = (w9280 & ~w9273) | (w9280 & w31694) | (~w9273 & w31694);
assign w9282 = ~w9271 & ~w9281;
assign w9283 = w7944 & ~w9282;
assign w9284 = ~w7944 & w9282;
assign w9285 = ~w9283 & ~w9284;
assign w9286 = w7931 & ~w9285;
assign w9287 = ~w7931 & w9285;
assign w9288 = ~w9286 & ~w9287;
assign w9289 = w9270 & w9288;
assign w9290 = ~w9270 & ~w9288;
assign w9291 = ~w9289 & ~w9290;
assign w9292 = w8897 & w9291;
assign w9293 = ~w9269 & w9292;
assign w9294 = ~w3475 & w6304;
assign w9295 = (w6059 & ~w3267) | (w6059 & w33910) | (~w3267 & w33910);
assign w9296 = ~w3326 & w6061;
assign w9297 = ~w9294 & ~w9295;
assign w9298 = ~w9296 & w9297;
assign w9299 = (w9298 & ~w6108) | (w9298 & w33911) | (~w6108 & w33911);
assign w9300 = a_17 & ~w9299;
assign w9301 = (~w6108 & w33912) | (~w6108 & w33913) | (w33912 & w33913);
assign w9302 = ~w9300 & ~w9301;
assign w9303 = w9293 & ~w9302;
assign w9304 = w8897 & ~w9269;
assign w9305 = ~w9291 & ~w9302;
assign w9306 = ~w9304 & w9305;
assign w9307 = ~w9303 & ~w9306;
assign w9308 = (~w9291 & w9269) | (~w9291 & w33914) | (w9269 & w33914);
assign w9309 = ~w9293 & w9302;
assign w9310 = ~w9308 & w9309;
assign w9311 = w9307 & ~w9310;
assign w9312 = ~w3403 & w6446;
assign w9313 = ~w2306 & w6996;
assign w9314 = (w6998 & ~w3538) | (w6998 & w33915) | (~w3538 & w33915);
assign w9315 = ~w9313 & ~w9314;
assign w9316 = ~w9312 & w9315;
assign w9317 = (w9316 & ~w5706) | (w9316 & w33916) | (~w5706 & w33916);
assign w9318 = a_14 & w9317;
assign w9319 = (w5706 & w33917) | (w5706 & w33918) | (w33917 & w33918);
assign w9320 = ~w9318 & ~w9319;
assign w9321 = w9311 & ~w9320;
assign w9322 = ~w9311 & w9320;
assign w9323 = ~w9321 & ~w9322;
assign w9324 = w8878 & w8918;
assign w9325 = ~w8912 & ~w8918;
assign w9326 = ~w9324 & ~w9325;
assign w9327 = ~w2075 & w7511;
assign w9328 = ~w2393 & w7192;
assign w9329 = ~w3615 & w7489;
assign w9330 = ~w9328 & ~w9329;
assign w9331 = ~w9327 & w9330;
assign w9332 = (w9331 & ~w5227) | (w9331 & w33919) | (~w5227 & w33919);
assign w9333 = a_11 & ~w9332;
assign w9334 = (~w5227 & w33920) | (~w5227 & w33921) | (w33920 & w33921);
assign w9335 = ~w9333 & ~w9334;
assign w9336 = ~w9324 & w31695;
assign w9337 = (w9335 & w9324) | (w9335 & w31696) | (w9324 & w31696);
assign w9338 = ~w9336 & ~w9337;
assign w9339 = w9323 & ~w9338;
assign w9340 = ~w9323 & w9338;
assign w9341 = ~w9339 & ~w9340;
assign w9342 = w9267 & w9341;
assign w9343 = ~w9267 & ~w9341;
assign w9344 = ~w9342 & ~w9343;
assign w9345 = ~w8304 & w9344;
assign w9346 = w8304 & ~w9344;
assign w9347 = ~w9345 & ~w9346;
assign w9348 = w9265 & ~w9347;
assign w9349 = ~w9265 & w9347;
assign w9350 = ~w9348 & ~w9349;
assign w9351 = w8304 & w9350;
assign w9352 = ~w2306 & w8298;
assign w9353 = ~w2393 & w8295;
assign w9354 = (w8277 & ~w3538) | (w8277 & w33922) | (~w3538 & w33922);
assign w9355 = ~w9352 & ~w9353;
assign w9356 = ~w9354 & w9355;
assign w9357 = (w9356 & ~w5483) | (w9356 & w33923) | (~w5483 & w33923);
assign w9358 = a_8 & ~w9357;
assign w9359 = (~w5483 & w33924) | (~w5483 & w33925) | (w33924 & w33925);
assign w9360 = ~w9358 & ~w9359;
assign w9361 = w9231 & w9360;
assign w9362 = w9213 & w9361;
assign w9363 = ~w9231 & w9360;
assign w9364 = ~w9213 & w9363;
assign w9365 = ~w9362 & ~w9364;
assign w9366 = ~w9027 & ~w9210;
assign w9367 = ~w9019 & ~w9366;
assign w9368 = w9001 & ~w9004;
assign w9369 = ~w3403 & w8277;
assign w9370 = ~w2306 & w8295;
assign w9371 = (w8298 & ~w3538) | (w8298 & w33926) | (~w3538 & w33926);
assign w9372 = ~w9370 & ~w9371;
assign w9373 = ~w9369 & w9372;
assign w9374 = (w9373 & ~w5706) | (w9373 & w33927) | (~w5706 & w33927);
assign w9375 = a_8 & ~w9374;
assign w9376 = (~w5706 & w33928) | (~w5706 & w33929) | (w33928 & w33929);
assign w9377 = ~w9375 & ~w9376;
assign w9378 = ~w9368 & w9377;
assign w9379 = ~w9367 & w9378;
assign w9380 = w9368 & w9377;
assign w9381 = w9367 & w9380;
assign w9382 = ~w9379 & ~w9381;
assign w9383 = w9365 & w9382;
assign w9384 = ~w9231 & ~w9360;
assign w9385 = w9213 & w9384;
assign w9386 = w9231 & ~w9360;
assign w9387 = ~w9213 & w9386;
assign w9388 = ~w9385 & ~w9387;
assign w9389 = ~w9383 & w9388;
assign w9390 = ~w3475 & w8295;
assign w9391 = (w8277 & ~w3267) | (w8277 & w33930) | (~w3267 & w33930);
assign w9392 = ~w3326 & w8298;
assign w9393 = ~w9390 & ~w9391;
assign w9394 = ~w9392 & w9393;
assign w9395 = (w9394 & ~w6108) | (w9394 & w33931) | (~w6108 & w33931);
assign w9396 = a_8 & ~w9395;
assign w9397 = (~w6108 & w33932) | (~w6108 & w33933) | (w33932 & w33933);
assign w9398 = ~w9396 & ~w9397;
assign w9399 = w9207 & ~w9398;
assign w9400 = ~w9176 & w9181;
assign w9401 = w9205 & ~w9398;
assign w9402 = ~w9400 & w9401;
assign w9403 = ~w9399 & ~w9402;
assign w9404 = (w9205 & w9176) | (w9205 & w33934) | (w9176 & w33934);
assign w9405 = ~w9207 & w9398;
assign w9406 = ~w9404 & w9405;
assign w9407 = ~w3326 & w8295;
assign w9408 = (w8298 & ~w3267) | (w8298 & w33935) | (~w3267 & w33935);
assign w9409 = ~w3196 & w8277;
assign w9410 = ~w9408 & ~w9409;
assign w9411 = ~w9407 & w9410;
assign w9412 = (w9411 & w5903) | (w9411 & w33936) | (w5903 & w33936);
assign w9413 = a_8 & ~w9412;
assign w9414 = (w5903 & w33937) | (w5903 & w33938) | (w33937 & w33938);
assign w9415 = ~w9413 & ~w9414;
assign w9416 = ~w9052 & ~w9160;
assign w9417 = w9174 & w9181;
assign w9418 = ~w9416 & ~w9417;
assign w9419 = w9416 & w9417;
assign w9420 = ~w9418 & ~w9419;
assign w9421 = w9415 & ~w9420;
assign w9422 = ~w9406 & ~w9421;
assign w9423 = w9403 & ~w9422;
assign w9424 = ~w9054 & w9159;
assign w9425 = ~w9160 & ~w9424;
assign w9426 = ~w3196 & w8298;
assign w9427 = (w8295 & ~w3267) | (w8295 & w33939) | (~w3267 & w33939);
assign w9428 = ~w3139 & w8277;
assign w9429 = w6222 & w33940;
assign w9430 = ~w9426 & ~w9427;
assign w9431 = ~w9428 & w9430;
assign w9432 = ~w9429 & w33941;
assign w9433 = (~a_8 & w9429) | (~a_8 & w33942) | (w9429 & w33942);
assign w9434 = ~w9432 & ~w9433;
assign w9435 = w9425 & ~w9434;
assign w9436 = ~w9071 & ~w9119;
assign w9437 = ~w9120 & ~w9436;
assign w9438 = ~w3007 & w8298;
assign w9439 = ~w3049 & w8295;
assign w9440 = ~w2917 & w8277;
assign w9441 = ~w9438 & ~w9439;
assign w9442 = ~w9440 & w9441;
assign w9443 = (w9442 & ~w6194) | (w9442 & w33943) | (~w6194 & w33943);
assign w9444 = a_8 & ~w9443;
assign w9445 = (~w6194 & w33944) | (~w6194 & w33945) | (w33944 & w33945);
assign w9446 = ~w9444 & ~w9445;
assign w9447 = w9437 & w9446;
assign w9448 = ~w9437 & ~w9446;
assign w9449 = ~w9447 & ~w9448;
assign w9450 = (w8298 & ~w2766) | (w8298 & w33946) | (~w2766 & w33946);
assign w9451 = ~w2546 & w8277;
assign w9452 = ~w2835 & w8295;
assign w9453 = ~w9450 & ~w9451;
assign w9454 = w9453 & w33947;
assign w9455 = (w9454 & ~w6733) | (w9454 & w31697) | (~w6733 & w31697);
assign w9456 = w8268 & ~w8272;
assign w9457 = (a_8 & ~w9453) | (a_8 & w33948) | (~w9453 & w33948);
assign w9458 = (~w9457 & ~w6733) | (~w9457 & w31698) | (~w6733 & w31698);
assign w9459 = ~w9455 & w9458;
assign w9460 = (a_11 & w9078) | (a_11 & w33949) | (w9078 & w33949);
assign w9461 = ~w9077 & w9460;
assign w9462 = w9077 & ~w9460;
assign w9463 = ~w9461 & ~w9462;
assign w9464 = w9459 & w9463;
assign w9465 = ~w9459 & ~w9463;
assign w9466 = ~w9464 & ~w9465;
assign w9467 = w7970 & w8278;
assign w9468 = (w8298 & ~w2479) | (w8298 & w33950) | (~w2479 & w33950);
assign w9469 = ~w2677 & w8295;
assign w9470 = (w8277 & ~w2600) | (w8277 & w33951) | (~w2600 & w33951);
assign w9471 = ~w9469 & w33952;
assign w9472 = ~w9467 & w9471;
assign w9473 = ~w7287 & w8278;
assign w9474 = (w8295 & ~w2479) | (w8295 & w31699) | (~w2479 & w31699);
assign w9475 = (w8298 & ~w2600) | (w8298 & w31700) | (~w2600 & w31700);
assign w9476 = ~w9474 & ~w9475;
assign w9477 = (~w8272 & ~w2600) | (~w8272 & w31701) | (~w2600 & w31701);
assign w9478 = a_8 & w9477;
assign w9479 = w9476 & ~w9478;
assign w9480 = ~w9473 & w9479;
assign w9481 = ~w9473 & w31702;
assign w9482 = (~w9082 & ~w9472) | (~w9082 & w31703) | (~w9472 & w31703);
assign w9483 = w6675 & w9456;
assign w9484 = w8267 & ~w8272;
assign w9485 = w6675 & w9484;
assign w9486 = ~w2677 & w8298;
assign w9487 = ~w2546 & w8295;
assign w9488 = (w8277 & ~w2479) | (w8277 & w33953) | (~w2479 & w33953);
assign w9489 = ~w9486 & ~w9487;
assign w9490 = w9489 & w33954;
assign w9491 = (~a_8 & ~w9489) | (~a_8 & w33955) | (~w9489 & w33955);
assign w9492 = ~w9490 & ~w9491;
assign w9493 = ~w9485 & w9492;
assign w9494 = ~w9483 & ~w9493;
assign w9495 = ~w9482 & w9494;
assign w9496 = (w8295 & ~w2766) | (w8295 & w33956) | (~w2766 & w33956);
assign w9497 = ~w2677 & w8277;
assign w9498 = ~w2546 & w8298;
assign w9499 = ~w9496 & ~w9497;
assign w9500 = ~w9498 & w9499;
assign w9501 = (w9500 & ~w7625) | (w9500 & w31704) | (~w7625 & w31704);
assign w9502 = w7286 & w9061;
assign w9503 = ~w9081 & w9083;
assign w9504 = ~w9502 & ~w9503;
assign w9505 = ~w9085 & w9504;
assign w9506 = (a_8 & w9085) | (a_8 & w31705) | (w9085 & w31705);
assign w9507 = ~w9085 & w31706;
assign w9508 = ~w9506 & ~w9507;
assign w9509 = w9501 & w9508;
assign w9510 = ~w9501 & ~w9508;
assign w9511 = ~w9509 & ~w9510;
assign w9512 = ~w9495 & w9511;
assign w9513 = ~w9505 & ~w9511;
assign w9514 = ~w9512 & ~w9513;
assign w9515 = w9466 & w9514;
assign w9516 = ~w9464 & ~w9515;
assign w9517 = w9100 & ~w9116;
assign w9518 = ~w9117 & ~w9517;
assign w9519 = w6545 & w8278;
assign w9520 = ~w6544 & w8278;
assign w9521 = ~w2920 & w31707;
assign w9522 = ~w3007 & w8295;
assign w9523 = ~w2917 & w8298;
assign w9524 = ~w2835 & w8277;
assign w9525 = ~w9522 & ~w9523;
assign w9526 = ~w9524 & w9525;
assign w9527 = ~w9521 & w9526;
assign w9528 = ~w9519 & w9527;
assign w9529 = a_8 & ~w9528;
assign w9530 = ~a_8 & w9528;
assign w9531 = ~w9529 & ~w9530;
assign w9532 = w9518 & ~w9531;
assign w9533 = ~w2917 & w8295;
assign w9534 = ~w2835 & w8298;
assign w9535 = (w8277 & ~w2766) | (w8277 & w33957) | (~w2766 & w33957);
assign w9536 = ~w9533 & ~w9534;
assign w9537 = ~w9535 & w9536;
assign w9538 = (~w6784 & w33958) | (~w6784 & w33959) | (w33958 & w33959);
assign w9539 = (w6784 & w33960) | (w6784 & w33961) | (w33960 & w33961);
assign w9540 = ~w9538 & ~w9539;
assign w9541 = w9077 & w31709;
assign w9542 = ~w9087 & ~w9541;
assign w9543 = w9099 & ~w9542;
assign w9544 = ~w9099 & w9542;
assign w9545 = ~w9543 & ~w9544;
assign w9546 = w9540 & ~w9545;
assign w9547 = ~w9540 & w9545;
assign w9548 = ~w9546 & ~w9547;
assign w9549 = ~w9532 & w9548;
assign w9550 = ~w9516 & w9549;
assign w9551 = ~w9518 & w9531;
assign w9552 = ~w9532 & w9546;
assign w9553 = ~w9551 & ~w9552;
assign w9554 = ~w9550 & w9553;
assign w9555 = w9449 & ~w9554;
assign w9556 = ~w3007 & w8277;
assign w9557 = ~w3139 & w8295;
assign w9558 = ~w3049 & w8298;
assign w9559 = ~w9556 & ~w9557;
assign w9560 = ~w9558 & w9559;
assign w9561 = (w9560 & w6505) | (w9560 & w33962) | (w6505 & w33962);
assign w9562 = a_8 & ~w9561;
assign w9563 = (w6505 & w33963) | (w6505 & w33964) | (w33963 & w33964);
assign w9564 = ~w9562 & ~w9563;
assign w9565 = w9153 & w9564;
assign w9566 = w9121 & w9565;
assign w9567 = ~w9153 & w9564;
assign w9568 = ~w9121 & w9567;
assign w9569 = ~w9566 & ~w9568;
assign w9570 = ~w9447 & w9569;
assign w9571 = ~w9555 & w9570;
assign w9572 = ~w9153 & ~w9564;
assign w9573 = w9121 & w9572;
assign w9574 = w9153 & ~w9564;
assign w9575 = ~w9121 & w9574;
assign w9576 = ~w9573 & ~w9575;
assign w9577 = ~w9069 & ~w9151;
assign w9578 = ~w9120 & w9577;
assign w9579 = ~w9152 & ~w9578;
assign w9580 = w6491 & w9456;
assign w9581 = ~w6216 & w33965;
assign w9582 = (w9581 & w3058) | (w9581 & w33966) | (w3058 & w33966);
assign w9583 = ~w3196 & w8295;
assign w9584 = ~w3139 & w8298;
assign w9585 = ~w3049 & w8277;
assign w9586 = ~w9583 & ~w9584;
assign w9587 = (~a_8 & ~w9586) | (~a_8 & w33967) | (~w9586 & w33967);
assign w9588 = w9586 & w33968;
assign w9589 = ~w9587 & ~w9588;
assign w9590 = (w9589 & ~w9582) | (w9589 & w31710) | (~w9582 & w31710);
assign w9591 = ~w9580 & ~w9590;
assign w9592 = w9136 & ~w9591;
assign w9593 = ~w9136 & w9591;
assign w9594 = ~w9592 & ~w9593;
assign w9595 = w9123 & ~w9594;
assign w9596 = ~w9123 & w9594;
assign w9597 = ~w9595 & ~w9596;
assign w9598 = w9579 & w9597;
assign w9599 = ~w9579 & ~w9597;
assign w9600 = ~w9598 & ~w9599;
assign w9601 = w9576 & ~w9600;
assign w9602 = ~w9571 & w9601;
assign w9603 = w9591 & w9600;
assign w9604 = ~w9602 & ~w9603;
assign w9605 = ~w9425 & w9434;
assign w9606 = ~w9435 & ~w9605;
assign w9607 = ~w9604 & w9606;
assign w9608 = ~w9435 & ~w9607;
assign w9609 = w9415 & w9417;
assign w9610 = ~w9415 & ~w9417;
assign w9611 = ~w9609 & ~w9610;
assign w9612 = w9416 & w9611;
assign w9613 = ~w9416 & ~w9611;
assign w9614 = ~w9612 & ~w9613;
assign w9615 = w9403 & ~w9614;
assign w9616 = ~w9608 & w9615;
assign w9617 = ~w9423 & ~w9616;
assign w9618 = ~w3475 & w8298;
assign w9619 = ~w3403 & w8295;
assign w9620 = ~w3326 & w8277;
assign w9621 = ~w9618 & ~w9619;
assign w9622 = ~w9620 & w9621;
assign w9623 = (w9622 & ~w5923) | (w9622 & w33969) | (~w5923 & w33969);
assign w9624 = a_8 & ~w9623;
assign w9625 = (~w5923 & w33970) | (~w5923 & w33971) | (w33970 & w33971);
assign w9626 = ~w9624 & ~w9625;
assign w9627 = ~w9038 & w9626;
assign w9628 = w9038 & ~w9626;
assign w9629 = ~w9627 & ~w9628;
assign w9630 = w9029 & ~w9629;
assign w9631 = ~w9029 & w9629;
assign w9632 = ~w9630 & ~w9631;
assign w9633 = w9209 & w9632;
assign w9634 = ~w9209 & ~w9632;
assign w9635 = ~w9633 & ~w9634;
assign w9636 = ~w9617 & ~w9635;
assign w9637 = w9626 & w9635;
assign w9638 = ~w3403 & w8298;
assign w9639 = (w8295 & ~w3538) | (w8295 & w33972) | (~w3538 & w33972);
assign w9640 = ~w3475 & w8277;
assign w9641 = ~w9638 & ~w9639;
assign w9642 = ~w9640 & w9641;
assign w9643 = (w9642 & ~w5652) | (w9642 & w33973) | (~w5652 & w33973);
assign w9644 = a_8 & ~w9643;
assign w9645 = (~w5652 & w33974) | (~w5652 & w33975) | (w33974 & w33975);
assign w9646 = ~w9644 & ~w9645;
assign w9647 = w9027 & w9646;
assign w9648 = ~w9210 & w9647;
assign w9649 = ~w9027 & w9646;
assign w9650 = w9210 & w9649;
assign w9651 = ~w9648 & ~w9650;
assign w9652 = ~w9637 & w9651;
assign w9653 = ~w9636 & w9652;
assign w9654 = ~w9027 & ~w9646;
assign w9655 = ~w9210 & w9654;
assign w9656 = w9027 & ~w9646;
assign w9657 = w9210 & w9656;
assign w9658 = ~w9655 & ~w9657;
assign w9659 = ~w9653 & w9658;
assign w9660 = ~w9368 & ~w9377;
assign w9661 = ~w9380 & ~w9660;
assign w9662 = w9367 & w9661;
assign w9663 = ~w9367 & ~w9661;
assign w9664 = ~w9662 & ~w9663;
assign w9665 = w9388 & ~w9664;
assign w9666 = w9659 & w9665;
assign w9667 = ~w9389 & ~w9666;
assign w9668 = (~w9233 & w9213) | (~w9233 & w33976) | (w9213 & w33976);
assign w9669 = ~w9243 & ~w9250;
assign w9670 = ~w3615 & w8295;
assign w9671 = ~w2393 & w8298;
assign w9672 = ~w2306 & w8277;
assign w9673 = ~w9670 & ~w9671;
assign w9674 = (a_8 & ~w9673) | (a_8 & w33977) | (~w9673 & w33977);
assign w9675 = w5463 & w8278;
assign w9676 = w9673 & w33978;
assign w9677 = ~w9675 & w9676;
assign w9678 = (~w9674 & ~w5463) | (~w9674 & w33979) | (~w5463 & w33979);
assign w9679 = ~w9677 & w9678;
assign w9680 = w8727 & ~w9679;
assign w9681 = ~w8727 & w9679;
assign w9682 = ~w9680 & ~w9681;
assign w9683 = w9669 & ~w9682;
assign w9684 = ~w9669 & w9682;
assign w9685 = ~w9683 & ~w9684;
assign w9686 = w9668 & w9685;
assign w9687 = ~w9668 & ~w9685;
assign w9688 = ~w9686 & ~w9687;
assign w9689 = ~w9667 & ~w9688;
assign w9690 = ~w2075 & w8295;
assign w9691 = ~w3615 & w8298;
assign w9692 = ~w2393 & w8277;
assign w9693 = ~w9691 & ~w9692;
assign w9694 = ~w9690 & w9693;
assign w9695 = (w9694 & ~w5227) | (w9694 & w33980) | (~w5227 & w33980);
assign w9696 = a_8 & ~w9695;
assign w9697 = (~w5227 & w33981) | (~w5227 & w33982) | (w33981 & w33982);
assign w9698 = ~w9696 & ~w9697;
assign w9699 = w9257 & w9698;
assign w9700 = w9255 & w9699;
assign w9701 = ~w9257 & w9698;
assign w9702 = ~w9255 & w9701;
assign w9703 = ~w9700 & ~w9702;
assign w9704 = w9247 & w9254;
assign w9705 = ~w9668 & ~w9704;
assign w9706 = w9668 & w9704;
assign w9707 = ~w9705 & ~w9706;
assign w9708 = w9679 & ~w9707;
assign w9709 = w9703 & ~w9708;
assign w9710 = ~w9689 & w9709;
assign w9711 = ~w9257 & ~w9698;
assign w9712 = w9255 & w9711;
assign w9713 = w9257 & ~w9698;
assign w9714 = ~w9255 & w9713;
assign w9715 = ~w9712 & ~w9714;
assign w9716 = ~w8964 & w33983;
assign w9717 = w8964 & w8975;
assign w9718 = w9254 & ~w9717;
assign w9719 = ~w9716 & w9718;
assign w9720 = ~w9249 & w9719;
assign w9721 = ~w8980 & ~w9720;
assign w9722 = ~w2148 & w8295;
assign w9723 = ~w3615 & w8277;
assign w9724 = ~w2075 & w8298;
assign w9725 = ~w9722 & ~w9723;
assign w9726 = (a_8 & ~w9725) | (a_8 & w33984) | (~w9725 & w33984);
assign w9727 = w5242 & w8278;
assign w9728 = w9725 & w33985;
assign w9729 = ~w9727 & w9728;
assign w9730 = (~w9726 & ~w5242) | (~w9726 & w33986) | (~w5242 & w33986);
assign w9731 = ~w9729 & w9730;
assign w9732 = ~w8943 & ~w9731;
assign w9733 = w8943 & w9731;
assign w9734 = ~w9732 & ~w9733;
assign w9735 = ~w8956 & ~w8983;
assign w9736 = ~w9734 & w9735;
assign w9737 = w9734 & ~w9735;
assign w9738 = ~w9736 & ~w9737;
assign w9739 = w9721 & w9738;
assign w9740 = ~w9721 & ~w9738;
assign w9741 = ~w9739 & ~w9740;
assign w9742 = w9715 & ~w9741;
assign w9743 = ~w9710 & w9742;
assign w9744 = w9731 & w9741;
assign w9745 = ~w2075 & w8277;
assign w9746 = (w8295 & ~w2235) | (w8295 & w33987) | (~w2235 & w33987);
assign w9747 = ~w2148 & w8298;
assign w9748 = ~w9746 & ~w9747;
assign w9749 = ~w9745 & w9748;
assign w9750 = (w9749 & ~w4962) | (w9749 & w33988) | (~w4962 & w33988);
assign w9751 = a_8 & ~w9750;
assign w9752 = (~w4962 & w33989) | (~w4962 & w33990) | (w33989 & w33990);
assign w9753 = ~w9751 & ~w9752;
assign w9754 = ~w8939 & w9753;
assign w9755 = w9260 & ~w9754;
assign w9756 = w8939 & w9753;
assign w9757 = ~w9260 & ~w9756;
assign w9758 = ~w9755 & ~w9757;
assign w9759 = ~w9744 & ~w9758;
assign w9760 = ~w9743 & w9759;
assign w9761 = ~w9265 & w9345;
assign w9762 = w8939 & ~w9753;
assign w9763 = w9260 & ~w9762;
assign w9764 = ~w8939 & ~w9753;
assign w9765 = ~w9260 & ~w9764;
assign w9766 = ~w9763 & ~w9765;
assign w9767 = (~w8304 & w8938) | (~w8304 & w31711) | (w8938 & w31711);
assign w9768 = ~w9344 & w9767;
assign w9769 = ~w9261 & w9768;
assign w9770 = ~w9766 & ~w9769;
assign w9771 = ~w9761 & w9770;
assign w9772 = ~w9760 & w9771;
assign w9773 = ~w9351 & ~w9772;
assign w9774 = ~a_2 & ~a_3;
assign w9775 = a_2 & a_3;
assign w9776 = ~w9774 & ~w9775;
assign w9777 = ~a_3 & ~a_4;
assign w9778 = a_3 & a_4;
assign w9779 = ~w9777 & ~w9778;
assign w9780 = ~w9776 & w9779;
assign w9781 = (w9780 & ~w1913) | (w9780 & w33991) | (~w1913 & w33991);
assign w9782 = ~a_4 & a_5;
assign w9783 = a_4 & ~a_5;
assign w9784 = ~w9782 & ~w9783;
assign w9785 = ~w9776 & ~w9779;
assign w9786 = ~w9784 & w9785;
assign w9787 = (w9786 & ~w2005) | (w9786 & w33992) | (~w2005 & w33992);
assign w9788 = w9776 & w9784;
assign w9789 = (w9788 & ~w1714) | (w9788 & w33993) | (~w1714 & w33993);
assign w9790 = w9776 & ~w9784;
assign w9791 = ~w9781 & ~w9787;
assign w9792 = ~w9789 & w9791;
assign w9793 = (w9792 & ~w4592) | (w9792 & w33994) | (~w4592 & w33994);
assign w9794 = a_5 & w9793;
assign w9795 = (w4592 & w33995) | (w4592 & w33996) | (w33995 & w33996);
assign w9796 = ~w9794 & ~w9795;
assign w9797 = ~w9323 & w9326;
assign w9798 = w9323 & ~w9326;
assign w9799 = ~w9797 & ~w9798;
assign w9800 = w9335 & w9799;
assign w9801 = w9267 & w9800;
assign w9802 = w9335 & ~w9799;
assign w9803 = ~w9267 & w9802;
assign w9804 = ~w9801 & ~w9803;
assign w9805 = ~w9264 & w9804;
assign w9806 = ~w9261 & w9805;
assign w9807 = ~w9344 & w9804;
assign w9808 = ~w9806 & ~w9807;
assign w9809 = w4810 & w9456;
assign w9810 = (w8277 & ~w2235) | (w8277 & w33997) | (~w2235 & w33997);
assign w9811 = (w8298 & ~w3712) | (w8298 & w33998) | (~w3712 & w33998);
assign w9812 = (w8295 & ~w3658) | (w8295 & w33999) | (~w3658 & w33999);
assign w9813 = ~w9810 & ~w9811;
assign w9814 = ~w9812 & w9813;
assign w9815 = a_8 & ~w9814;
assign w9816 = ~a_8 & w9814;
assign w9817 = (w9816 & ~w4810) | (w9816 & w34000) | (~w4810 & w34000);
assign w9818 = ~w9809 & ~w9815;
assign w9819 = ~w9817 & w9818;
assign w9820 = w9321 & w9326;
assign w9821 = ~w9311 & ~w9320;
assign w9822 = ~w9326 & w9821;
assign w9823 = ~w9820 & ~w9822;
assign w9824 = ~w9799 & w9823;
assign w9825 = ~w9266 & w9823;
assign w9826 = ~w9262 & w9825;
assign w9827 = ~w9824 & ~w9826;
assign w9828 = ~w9310 & ~w9325;
assign w9829 = ~w9324 & w9828;
assign w9830 = w9307 & ~w9829;
assign w9831 = w9282 & ~w9291;
assign w9832 = ~w9293 & ~w9831;
assign w9833 = ~w3475 & w6061;
assign w9834 = ~w3403 & w6304;
assign w9835 = ~w3326 & w6059;
assign w9836 = ~w9833 & ~w9834;
assign w9837 = ~w9835 & w9836;
assign w9838 = (w9837 & ~w5923) | (w9837 & w34001) | (~w5923 & w34001);
assign w9839 = a_17 & w9838;
assign w9840 = (w5923 & w34002) | (w5923 & w34003) | (w34002 & w34003);
assign w9841 = ~w9839 & ~w9840;
assign w9842 = (w5816 & ~w3267) | (w5816 & w34004) | (~w3267 & w34004);
assign w9843 = ~w3196 & w5818;
assign w9844 = ~w3139 & w5308;
assign w9845 = w6222 & w34005;
assign w9846 = ~w9842 & ~w9843;
assign w9847 = ~w9844 & w9846;
assign w9848 = (a_20 & w9845) | (a_20 & w34006) | (w9845 & w34006);
assign w9849 = ~w9845 & w34007;
assign w9850 = ~w9848 & ~w9849;
assign w9851 = w8082 & ~w9850;
assign w9852 = w8045 & w9851;
assign w9853 = ~w8082 & ~w9850;
assign w9854 = ~w8045 & w9853;
assign w9855 = ~w9852 & ~w9854;
assign w9856 = ~w8082 & w9850;
assign w9857 = w8045 & w9856;
assign w9858 = w8082 & w9850;
assign w9859 = ~w8045 & w9858;
assign w9860 = ~w9857 & ~w9859;
assign w9861 = w9855 & w9860;
assign w9862 = w9841 & w9861;
assign w9863 = ~w9841 & ~w9861;
assign w9864 = ~w9862 & ~w9863;
assign w9865 = ~w9832 & w9864;
assign w9866 = w9832 & ~w9864;
assign w9867 = ~w9865 & ~w9866;
assign w9868 = ~w9830 & w9867;
assign w9869 = w9830 & ~w9867;
assign w9870 = ~w9868 & ~w9869;
assign w9871 = ~w2306 & w6998;
assign w9872 = ~w2393 & w6996;
assign w9873 = (w6446 & ~w3538) | (w6446 & w34008) | (~w3538 & w34008);
assign w9874 = ~w9871 & ~w9872;
assign w9875 = ~w9873 & w9874;
assign w9876 = (w9875 & ~w5483) | (w9875 & w34009) | (~w5483 & w34009);
assign w9877 = a_14 & ~w9876;
assign w9878 = (~w5483 & w34010) | (~w5483 & w34011) | (w34010 & w34011);
assign w9879 = ~w9877 & ~w9878;
assign w9880 = ~w2148 & w7511;
assign w9881 = ~w3615 & w7192;
assign w9882 = ~w2075 & w7489;
assign w9883 = ~w9880 & ~w9881;
assign w9884 = (a_11 & ~w9883) | (a_11 & w34012) | (~w9883 & w34012);
assign w9885 = w5242 & w7193;
assign w9886 = w9883 & w34013;
assign w9887 = ~w9885 & w9886;
assign w9888 = (~w9884 & ~w5242) | (~w9884 & w34014) | (~w5242 & w34014);
assign w9889 = ~w9887 & w9888;
assign w9890 = w9879 & ~w9889;
assign w9891 = ~w9879 & w9889;
assign w9892 = ~w9890 & ~w9891;
assign w9893 = w9870 & ~w9892;
assign w9894 = ~w9870 & w9892;
assign w9895 = ~w9893 & ~w9894;
assign w9896 = w9827 & w9895;
assign w9897 = ~w9827 & ~w9895;
assign w9898 = ~w9896 & ~w9897;
assign w9899 = w9819 & ~w9898;
assign w9900 = ~w9819 & w9898;
assign w9901 = ~w9899 & ~w9900;
assign w9902 = w9808 & w9901;
assign w9903 = ~w9808 & ~w9901;
assign w9904 = ~w9902 & ~w9903;
assign w9905 = ~w9796 & ~w9904;
assign w9906 = w9773 & w9905;
assign w9907 = ~w9796 & w9904;
assign w9908 = ~w9773 & w9907;
assign w9909 = ~w9906 & ~w9908;
assign w9910 = ~w2306 & w9780;
assign w9911 = ~w2393 & w9788;
assign w9912 = (w9786 & ~w3538) | (w9786 & w34015) | (~w3538 & w34015);
assign w9913 = ~w9910 & ~w9911;
assign w9914 = ~w9912 & w9913;
assign w9915 = (w9914 & ~w5483) | (w9914 & w34016) | (~w5483 & w34016);
assign w9916 = a_5 & ~w9915;
assign w9917 = (~w5483 & w34017) | (~w5483 & w34018) | (w34017 & w34018);
assign w9918 = ~w9916 & ~w9917;
assign w9919 = ~w9635 & w9918;
assign w9920 = w9617 & w9919;
assign w9921 = w9635 & w9918;
assign w9922 = ~w9617 & w9921;
assign w9923 = ~w9920 & ~w9922;
assign w9924 = (~w9421 & w9608) | (~w9421 & w34019) | (w9608 & w34019);
assign w9925 = w9403 & ~w9406;
assign w9926 = ~w3403 & w9786;
assign w9927 = ~w2306 & w9788;
assign w9928 = (w9780 & ~w3538) | (w9780 & w34020) | (~w3538 & w34020);
assign w9929 = ~w9927 & ~w9928;
assign w9930 = ~w9926 & w9929;
assign w9931 = (w9930 & ~w5706) | (w9930 & w34021) | (~w5706 & w34021);
assign w9932 = a_5 & ~w9931;
assign w9933 = (~w5706 & w34022) | (~w5706 & w34023) | (w34022 & w34023);
assign w9934 = ~w9932 & ~w9933;
assign w9935 = ~w9925 & w9934;
assign w9936 = ~w9924 & w9935;
assign w9937 = w9925 & w9934;
assign w9938 = w9924 & w9937;
assign w9939 = ~w9936 & ~w9938;
assign w9940 = w9923 & w9939;
assign w9941 = w9635 & ~w9918;
assign w9942 = w9617 & w9941;
assign w9943 = ~w9635 & ~w9918;
assign w9944 = ~w9617 & w9943;
assign w9945 = ~w9942 & ~w9944;
assign w9946 = ~w9940 & w9945;
assign w9947 = ~w3403 & w9780;
assign w9948 = (w9788 & ~w3538) | (w9788 & w34024) | (~w3538 & w34024);
assign w9949 = ~w3475 & w9786;
assign w9950 = ~w9947 & ~w9948;
assign w9951 = ~w9949 & w9950;
assign w9952 = (w9951 & ~w5652) | (w9951 & w34025) | (~w5652 & w34025);
assign w9953 = a_5 & ~w9952;
assign w9954 = (~w5652 & w34026) | (~w5652 & w34027) | (w34026 & w34027);
assign w9955 = ~w9953 & ~w9954;
assign w9956 = w9614 & w9955;
assign w9957 = ~w9608 & w9956;
assign w9958 = ~w9614 & w9955;
assign w9959 = w9608 & w9958;
assign w9960 = ~w9957 & ~w9959;
assign w9961 = w9614 & ~w9955;
assign w9962 = ~w9958 & ~w9961;
assign w9963 = w9608 & w9962;
assign w9964 = ~w9608 & ~w9962;
assign w9965 = ~w9963 & ~w9964;
assign w9966 = w9960 & w9965;
assign w9967 = ~w3326 & w9780;
assign w9968 = (w9786 & ~w3267) | (w9786 & w34028) | (~w3267 & w34028);
assign w9969 = ~w3475 & w9788;
assign w9970 = ~w9967 & ~w9968;
assign w9971 = ~w9969 & w9970;
assign w9972 = (w9971 & ~w6108) | (w9971 & w34029) | (~w6108 & w34029);
assign w9973 = a_5 & ~w9972;
assign w9974 = (~w6108 & w34030) | (~w6108 & w34031) | (w34030 & w34031);
assign w9975 = ~w9973 & ~w9974;
assign w9976 = w9602 & ~w9975;
assign w9977 = ~w9571 & w9576;
assign w9978 = w9600 & ~w9975;
assign w9979 = ~w9977 & w9978;
assign w9980 = ~w9976 & ~w9979;
assign w9981 = (w9600 & w9571) | (w9600 & w34032) | (w9571 & w34032);
assign w9982 = ~w9602 & w9975;
assign w9983 = ~w9981 & w9982;
assign w9984 = ~w3326 & w9788;
assign w9985 = ~w3196 & w9786;
assign w9986 = (w9780 & ~w3267) | (w9780 & w34033) | (~w3267 & w34033);
assign w9987 = ~w9985 & ~w9986;
assign w9988 = ~w9984 & w9987;
assign w9989 = (w9988 & w5903) | (w9988 & w34034) | (w5903 & w34034);
assign w9990 = a_5 & ~w9989;
assign w9991 = (w5903 & w34035) | (w5903 & w34036) | (w34035 & w34036);
assign w9992 = ~w9990 & ~w9991;
assign w9993 = ~w9447 & ~w9555;
assign w9994 = w9569 & w9576;
assign w9995 = ~w9993 & ~w9994;
assign w9996 = w9993 & w9994;
assign w9997 = ~w9995 & ~w9996;
assign w9998 = w9992 & ~w9997;
assign w9999 = ~w9983 & ~w9998;
assign w10000 = w9980 & ~w9999;
assign w10001 = ~w9449 & w9554;
assign w10002 = ~w9555 & ~w10001;
assign w10003 = (w9788 & ~w3267) | (w9788 & w34037) | (~w3267 & w34037);
assign w10004 = ~w3196 & w9780;
assign w10005 = ~w3139 & w9786;
assign w10006 = w6222 & w34038;
assign w10007 = ~w10003 & ~w10004;
assign w10008 = ~w10005 & w10007;
assign w10009 = ~w10006 & w34039;
assign w10010 = (~a_5 & w10006) | (~a_5 & w34040) | (w10006 & w34040);
assign w10011 = ~w10009 & ~w10010;
assign w10012 = w10002 & ~w10011;
assign w10013 = ~w9466 & ~w9514;
assign w10014 = ~w9515 & ~w10013;
assign w10015 = ~w3049 & w9788;
assign w10016 = ~w3007 & w9780;
assign w10017 = ~w2917 & w9786;
assign w10018 = ~w10015 & ~w10016;
assign w10019 = ~w10017 & w10018;
assign w10020 = (w10019 & ~w6194) | (w10019 & w34041) | (~w6194 & w34041);
assign w10021 = a_5 & w10020;
assign w10022 = (w6194 & w34042) | (w6194 & w34043) | (w34042 & w34043);
assign w10023 = ~w10021 & ~w10022;
assign w10024 = w10014 & ~w10023;
assign w10025 = ~w10014 & w10023;
assign w10026 = ~w10024 & ~w10025;
assign w10027 = ~w2835 & w9788;
assign w10028 = (w9780 & ~w2766) | (w9780 & w34044) | (~w2766 & w34044);
assign w10029 = ~w2546 & w9786;
assign w10030 = ~w10027 & ~w10028;
assign w10031 = w10030 & w34045;
assign w10032 = (w10031 & ~w6733) | (w10031 & w31712) | (~w6733 & w31712);
assign w10033 = w9776 & w9782;
assign w10034 = (a_5 & ~w10030) | (a_5 & w34046) | (~w10030 & w34046);
assign w10035 = (~w10034 & ~w6733) | (~w10034 & w31713) | (~w6733 & w31713);
assign w10036 = ~w10032 & w10035;
assign w10037 = (a_8 & w9473) | (a_8 & w34047) | (w9473 & w34047);
assign w10038 = ~w9472 & w10037;
assign w10039 = w9472 & ~w10037;
assign w10040 = ~w10038 & ~w10039;
assign w10041 = w10036 & w10040;
assign w10042 = ~w10036 & ~w10040;
assign w10043 = ~w10041 & ~w10042;
assign w10044 = (w9776 & ~w2600) | (w9776 & w34048) | (~w2600 & w34048);
assign w10045 = a_5 & w10044;
assign w10046 = ~w7287 & w9790;
assign w10047 = (w9780 & ~w2600) | (w9780 & w34049) | (~w2600 & w34049);
assign w10048 = (w9788 & ~w2479) | (w9788 & w34050) | (~w2479 & w34050);
assign w10049 = ~w10047 & ~w10048;
assign w10050 = (w10049 & w7287) | (w10049 & w34051) | (w7287 & w34051);
assign w10051 = ~w10046 & w31714;
assign w10052 = ~w2677 & w9788;
assign w10053 = (w9786 & ~w2600) | (w9786 & w34052) | (~w2600 & w34052);
assign w10054 = (w9780 & ~w2479) | (w9780 & w34053) | (~w2479 & w34053);
assign w10055 = w7970 & w9790;
assign w10056 = ~w10052 & w34054;
assign w10057 = ~w10055 & w10056;
assign w10058 = ~w10046 & w34055;
assign w10059 = (~w9477 & ~w10057) | (~w9477 & w34056) | (~w10057 & w34056);
assign w10060 = w6675 & w10033;
assign w10061 = w9776 & w9783;
assign w10062 = w6675 & w10061;
assign w10063 = ~w2677 & w9780;
assign w10064 = ~w2546 & w9788;
assign w10065 = (w9786 & ~w2479) | (w9786 & w34057) | (~w2479 & w34057);
assign w10066 = ~w10063 & ~w10064;
assign w10067 = w10066 & w34058;
assign w10068 = (~a_5 & ~w10066) | (~a_5 & w34059) | (~w10066 & w34059);
assign w10069 = ~w10067 & ~w10068;
assign w10070 = ~w10062 & w10069;
assign w10071 = ~w10060 & ~w10070;
assign w10072 = ~w10059 & w10071;
assign w10073 = ~w2546 & w9780;
assign w10074 = (w9788 & ~w2766) | (w9788 & w34060) | (~w2766 & w34060);
assign w10075 = ~w2677 & w9786;
assign w10076 = ~w10073 & ~w10074;
assign w10077 = ~w10075 & w10076;
assign w10078 = (w10077 & ~w7625) | (w10077 & w31715) | (~w7625 & w31715);
assign w10079 = w7286 & w9456;
assign w10080 = ~w9476 & w9478;
assign w10081 = ~w10079 & ~w10080;
assign w10082 = ~w9480 & w10081;
assign w10083 = (a_5 & w9480) | (a_5 & w31716) | (w9480 & w31716);
assign w10084 = ~w9480 & w31717;
assign w10085 = ~w10083 & ~w10084;
assign w10086 = w10078 & w10085;
assign w10087 = ~w10078 & ~w10085;
assign w10088 = ~w10086 & ~w10087;
assign w10089 = ~w10072 & w10088;
assign w10090 = ~w10082 & ~w10088;
assign w10091 = ~w10089 & ~w10090;
assign w10092 = w10043 & w10091;
assign w10093 = ~w10041 & ~w10092;
assign w10094 = w9495 & ~w9511;
assign w10095 = ~w9512 & ~w10094;
assign w10096 = ~w2917 & w9780;
assign w10097 = ~w3007 & w9788;
assign w10098 = ~w2835 & w9786;
assign w10099 = ~w10096 & ~w10097;
assign w10100 = ~w10098 & w10099;
assign w10101 = (w10100 & w6547) | (w10100 & w34061) | (w6547 & w34061);
assign w10102 = a_5 & ~w10101;
assign w10103 = (w6547 & w34062) | (w6547 & w34063) | (w34062 & w34063);
assign w10104 = ~w10102 & ~w10103;
assign w10105 = w10095 & ~w10104;
assign w10106 = ~w2917 & w9788;
assign w10107 = ~w2835 & w9780;
assign w10108 = (w9786 & ~w2766) | (w9786 & w34064) | (~w2766 & w34064);
assign w10109 = ~w10106 & ~w10107;
assign w10110 = ~w10108 & w10109;
assign w10111 = (w6784 & w34065) | (w6784 & w34066) | (w34065 & w34066);
assign w10112 = (~w6784 & w34067) | (~w6784 & w34068) | (w34067 & w34068);
assign w10113 = ~w10111 & ~w10112;
assign w10114 = w9472 & w31719;
assign w10115 = ~w9482 & ~w10114;
assign w10116 = w9494 & ~w10115;
assign w10117 = ~w9494 & w10115;
assign w10118 = ~w10116 & ~w10117;
assign w10119 = w10113 & ~w10118;
assign w10120 = ~w10113 & w10118;
assign w10121 = ~w10119 & ~w10120;
assign w10122 = ~w10105 & w10121;
assign w10123 = ~w10093 & w10122;
assign w10124 = ~w10095 & w10104;
assign w10125 = ~w10105 & w10119;
assign w10126 = ~w10124 & ~w10125;
assign w10127 = ~w10123 & w10126;
assign w10128 = w10026 & ~w10127;
assign w10129 = ~w3007 & w9786;
assign w10130 = ~w3139 & w9788;
assign w10131 = ~w3049 & w9780;
assign w10132 = ~w10129 & ~w10130;
assign w10133 = ~w10131 & w10132;
assign w10134 = (w10133 & w6505) | (w10133 & w34069) | (w6505 & w34069);
assign w10135 = ~a_5 & w10134;
assign w10136 = (~w6505 & w34070) | (~w6505 & w34071) | (w34070 & w34071);
assign w10137 = ~w10135 & ~w10136;
assign w10138 = w9548 & w10137;
assign w10139 = w9516 & w10138;
assign w10140 = ~w9548 & w10137;
assign w10141 = ~w9516 & w10140;
assign w10142 = ~w10139 & ~w10141;
assign w10143 = ~w10024 & w10142;
assign w10144 = ~w10128 & w10143;
assign w10145 = ~w9464 & ~w9546;
assign w10146 = ~w9515 & w10145;
assign w10147 = ~w9547 & ~w10146;
assign w10148 = w6491 & w10033;
assign w10149 = ~w6216 & w34072;
assign w10150 = (w10149 & w3058) | (w10149 & w34073) | (w3058 & w34073);
assign w10151 = ~w3196 & w9788;
assign w10152 = ~w3139 & w9780;
assign w10153 = ~w3049 & w9786;
assign w10154 = ~w10151 & ~w10152;
assign w10155 = (~a_5 & ~w10154) | (~a_5 & w34074) | (~w10154 & w34074);
assign w10156 = w10154 & w34075;
assign w10157 = ~w10155 & ~w10156;
assign w10158 = (w10157 & ~w10150) | (w10157 & w31720) | (~w10150 & w31720);
assign w10159 = ~w10148 & ~w10158;
assign w10160 = w9531 & ~w10159;
assign w10161 = ~w9531 & w10159;
assign w10162 = ~w10160 & ~w10161;
assign w10163 = w9518 & ~w10162;
assign w10164 = ~w9518 & w10162;
assign w10165 = ~w10163 & ~w10164;
assign w10166 = w10147 & w10165;
assign w10167 = ~w10147 & ~w10165;
assign w10168 = ~w10166 & ~w10167;
assign w10169 = w9516 & ~w9548;
assign w10170 = ~w9516 & w9548;
assign w10171 = ~w10169 & ~w10170;
assign w10172 = ~w10137 & ~w10171;
assign w10173 = ~w10168 & ~w10172;
assign w10174 = ~w10144 & w10173;
assign w10175 = w10159 & w10168;
assign w10176 = ~w10174 & ~w10175;
assign w10177 = ~w10002 & w10011;
assign w10178 = ~w10012 & ~w10177;
assign w10179 = ~w10176 & w10178;
assign w10180 = ~w10012 & ~w10179;
assign w10181 = w9992 & w9994;
assign w10182 = ~w9992 & ~w9994;
assign w10183 = ~w10181 & ~w10182;
assign w10184 = w9993 & w10183;
assign w10185 = ~w9993 & ~w10183;
assign w10186 = ~w10184 & ~w10185;
assign w10187 = w9980 & ~w10186;
assign w10188 = ~w10180 & w10187;
assign w10189 = ~w10000 & ~w10188;
assign w10190 = w9604 & ~w9606;
assign w10191 = ~w9607 & ~w10190;
assign w10192 = ~w3475 & w9780;
assign w10193 = ~w3403 & w9788;
assign w10194 = ~w3326 & w9786;
assign w10195 = ~w10192 & ~w10193;
assign w10196 = ~w10194 & w10195;
assign w10197 = (w10196 & ~w5923) | (w10196 & w34076) | (~w5923 & w34076);
assign w10198 = a_5 & w10197;
assign w10199 = (w5923 & w34077) | (w5923 & w34078) | (w34077 & w34078);
assign w10200 = ~w10198 & ~w10199;
assign w10201 = ~w10191 & w10200;
assign w10202 = ~w10189 & ~w10201;
assign w10203 = w10191 & ~w10200;
assign w10204 = w9960 & ~w10203;
assign w10205 = ~w10202 & w10204;
assign w10206 = ~w9966 & ~w10205;
assign w10207 = ~w9925 & ~w9934;
assign w10208 = ~w9937 & ~w10207;
assign w10209 = w9924 & w10208;
assign w10210 = ~w9924 & ~w10208;
assign w10211 = ~w10209 & ~w10210;
assign w10212 = w9945 & ~w10211;
assign w10213 = w10206 & w10212;
assign w10214 = ~w9946 & ~w10213;
assign w10215 = (~w9637 & w9617) | (~w9637 & w34079) | (w9617 & w34079);
assign w10216 = w9651 & w9658;
assign w10217 = ~w2306 & w9786;
assign w10218 = ~w2393 & w9780;
assign w10219 = ~w3615 & w9788;
assign w10220 = ~w10217 & ~w10218;
assign w10221 = ~w10219 & w10220;
assign w10222 = (w10221 & ~w5463) | (w10221 & w34080) | (~w5463 & w34080);
assign w10223 = a_5 & ~w10222;
assign w10224 = (~w5463 & w34081) | (~w5463 & w34082) | (w34081 & w34082);
assign w10225 = ~w10223 & ~w10224;
assign w10226 = w10216 & ~w10225;
assign w10227 = ~w10216 & w10225;
assign w10228 = ~w10226 & ~w10227;
assign w10229 = w10215 & ~w10228;
assign w10230 = ~w10215 & w10228;
assign w10231 = ~w10229 & ~w10230;
assign w10232 = ~w10214 & ~w10231;
assign w10233 = ~w2075 & w9788;
assign w10234 = ~w3615 & w9780;
assign w10235 = ~w2393 & w9786;
assign w10236 = ~w10234 & ~w10235;
assign w10237 = ~w10233 & w10236;
assign w10238 = (w10237 & ~w5227) | (w10237 & w34083) | (~w5227 & w34083);
assign w10239 = a_5 & ~w10238;
assign w10240 = (~w5227 & w34084) | (~w5227 & w34085) | (w34084 & w34085);
assign w10241 = ~w10239 & ~w10240;
assign w10242 = w9664 & w10241;
assign w10243 = w9659 & w10242;
assign w10244 = ~w9664 & w10241;
assign w10245 = ~w9659 & w10244;
assign w10246 = ~w10243 & ~w10245;
assign w10247 = ~w10215 & w10227;
assign w10248 = w9658 & w10225;
assign w10249 = w9653 & w10248;
assign w10250 = ~w10247 & ~w10249;
assign w10251 = w10246 & w10250;
assign w10252 = ~w10232 & w10251;
assign w10253 = ~w9664 & ~w10241;
assign w10254 = w9659 & w10253;
assign w10255 = w9664 & ~w10241;
assign w10256 = ~w9659 & w10255;
assign w10257 = ~w10254 & ~w10256;
assign w10258 = ~w10252 & w10257;
assign w10259 = ~w2075 & w9786;
assign w10260 = (w9788 & ~w2235) | (w9788 & w34086) | (~w2235 & w34086);
assign w10261 = ~w2148 & w9780;
assign w10262 = ~w10260 & ~w10261;
assign w10263 = ~w10259 & w10262;
assign w10264 = (w10263 & ~w4962) | (w10263 & w34087) | (~w4962 & w34087);
assign w10265 = a_5 & ~w10264;
assign w10266 = (~w4962 & w34088) | (~w4962 & w34089) | (w34088 & w34089);
assign w10267 = ~w10265 & ~w10266;
assign w10268 = w9688 & ~w10267;
assign w10269 = w9667 & w10268;
assign w10270 = ~w9688 & ~w10267;
assign w10271 = ~w9667 & w10270;
assign w10272 = ~w10269 & ~w10271;
assign w10273 = (w9382 & ~w9659) | (w9382 & w34090) | (~w9659 & w34090);
assign w10274 = w9365 & w9388;
assign w10275 = ~w2075 & w9780;
assign w10276 = ~w2148 & w9788;
assign w10277 = ~w3615 & w9786;
assign w10278 = ~w10276 & ~w10277;
assign w10279 = ~w10275 & w10278;
assign w10280 = (w10279 & ~w5242) | (w10279 & w34091) | (~w5242 & w34091);
assign w10281 = a_5 & w10280;
assign w10282 = (w5242 & w34092) | (w5242 & w34093) | (w34092 & w34093);
assign w10283 = ~w10281 & ~w10282;
assign w10284 = w10274 & ~w10283;
assign w10285 = ~w10274 & w10283;
assign w10286 = ~w10284 & ~w10285;
assign w10287 = w10273 & w10286;
assign w10288 = ~w10273 & ~w10286;
assign w10289 = ~w10287 & ~w10288;
assign w10290 = w10272 & ~w10289;
assign w10291 = w10258 & w10290;
assign w10292 = ~w9688 & w10267;
assign w10293 = w9667 & w10292;
assign w10294 = w9688 & w10267;
assign w10295 = ~w9667 & w10294;
assign w10296 = ~w10293 & ~w10295;
assign w10297 = ~w10274 & ~w10283;
assign w10298 = ~w10273 & w10297;
assign w10299 = w10273 & w10284;
assign w10300 = ~w10298 & ~w10299;
assign w10301 = w10296 & w10300;
assign w10302 = w10272 & ~w10301;
assign w10303 = ~w10291 & ~w10302;
assign w10304 = (~w9708 & w9667) | (~w9708 & w34094) | (w9667 & w34094);
assign w10305 = w9703 & w9715;
assign w10306 = (w9788 & ~w3712) | (w9788 & w34095) | (~w3712 & w34095);
assign w10307 = ~w2148 & w9786;
assign w10308 = (w9780 & ~w2235) | (w9780 & w34096) | (~w2235 & w34096);
assign w10309 = w5103 & w9790;
assign w10310 = ~w10307 & w34097;
assign w10311 = (a_5 & w10309) | (a_5 & w34098) | (w10309 & w34098);
assign w10312 = ~w10309 & w34099;
assign w10313 = ~w10311 & ~w10312;
assign w10314 = w10305 & ~w10313;
assign w10315 = ~w10305 & w10313;
assign w10316 = ~w10314 & ~w10315;
assign w10317 = w10304 & w10316;
assign w10318 = ~w10304 & ~w10316;
assign w10319 = ~w10317 & ~w10318;
assign w10320 = ~w10303 & w10319;
assign w10321 = ~w9710 & w9715;
assign w10322 = (w9788 & ~w3658) | (w9788 & w34100) | (~w3658 & w34100);
assign w10323 = (w9780 & ~w3712) | (w9780 & w34101) | (~w3712 & w34101);
assign w10324 = (w9786 & ~w2235) | (w9786 & w34102) | (~w2235 & w34102);
assign w10325 = ~w10323 & ~w10324;
assign w10326 = ~w10322 & w10325;
assign w10327 = (w10326 & ~w4810) | (w10326 & w34103) | (~w4810 & w34103);
assign w10328 = a_5 & ~w10327;
assign w10329 = (~w4810 & w34104) | (~w4810 & w34105) | (w34104 & w34105);
assign w10330 = ~w10328 & ~w10329;
assign w10331 = w9741 & w10330;
assign w10332 = w10321 & w10331;
assign w10333 = ~w9741 & w10330;
assign w10334 = ~w10321 & w10333;
assign w10335 = ~w10332 & ~w10334;
assign w10336 = ~w10304 & ~w10305;
assign w10337 = w10304 & w10305;
assign w10338 = ~w10336 & ~w10337;
assign w10339 = w10313 & ~w10338;
assign w10340 = w10335 & ~w10339;
assign w10341 = ~w10320 & w10340;
assign w10342 = w9743 & ~w10330;
assign w10343 = w9741 & ~w10330;
assign w10344 = ~w10321 & w10343;
assign w10345 = ~w10342 & ~w10344;
assign w10346 = ~w8958 & ~w8985;
assign w10347 = ~w9731 & ~w10346;
assign w10348 = w9721 & w10347;
assign w10349 = ~w9731 & w10346;
assign w10350 = ~w9721 & w10349;
assign w10351 = w9715 & ~w10348;
assign w10352 = ~w10350 & w10351;
assign w10353 = (~w9744 & ~w10352) | (~w9744 & w31721) | (~w10352 & w31721);
assign w10354 = (w9780 & ~w3658) | (w9780 & w34106) | (~w3658 & w34106);
assign w10355 = (w9788 & ~w2005) | (w9788 & w34107) | (~w2005 & w34107);
assign w10356 = (w9786 & ~w3712) | (w9786 & w34108) | (~w3712 & w34108);
assign w10357 = (w9790 & w4790) | (w9790 & w34109) | (w4790 & w34109);
assign w10358 = ~w10355 & ~w10356;
assign w10359 = ~w10354 & w10358;
assign w10360 = (a_5 & w10357) | (a_5 & w34110) | (w10357 & w34110);
assign w10361 = ~w10357 & w34111;
assign w10362 = ~w10360 & ~w10361;
assign w10363 = ~w9260 & ~w10362;
assign w10364 = w9260 & w10362;
assign w10365 = ~w10363 & ~w10364;
assign w10366 = ~w9754 & ~w9762;
assign w10367 = w10365 & w10366;
assign w10368 = ~w10365 & ~w10366;
assign w10369 = ~w10367 & ~w10368;
assign w10370 = w10353 & w10369;
assign w10371 = ~w10353 & ~w10369;
assign w10372 = ~w10370 & ~w10371;
assign w10373 = w10345 & w10372;
assign w10374 = ~w10341 & w10373;
assign w10375 = (~w9766 & ~w9759) | (~w9766 & w31722) | (~w9759 & w31722);
assign w10376 = (w9786 & ~w3658) | (w9786 & w34112) | (~w3658 & w34112);
assign w10377 = (w9780 & ~w2005) | (w9780 & w34113) | (~w2005 & w34113);
assign w10378 = (w9788 & ~w1913) | (w9788 & w34114) | (~w1913 & w34114);
assign w10379 = ~w10377 & ~w10378;
assign w10380 = ~w10376 & w10379;
assign w10381 = (w10380 & w4578) | (w10380 & w34115) | (w4578 & w34115);
assign w10382 = a_5 & ~w10381;
assign w10383 = (w4578 & w34116) | (w4578 & w34117) | (w34116 & w34117);
assign w10384 = ~w10382 & ~w10383;
assign w10385 = w9350 & w10384;
assign w10386 = w10375 & w10385;
assign w10387 = ~w9350 & w10384;
assign w10388 = ~w10375 & w10387;
assign w10389 = ~w10386 & ~w10388;
assign w10390 = ~w9758 & ~w9766;
assign w10391 = ~w10353 & ~w10390;
assign w10392 = w10353 & w10390;
assign w10393 = ~w10391 & ~w10392;
assign w10394 = w10362 & ~w10393;
assign w10395 = w10389 & ~w10394;
assign w10396 = ~w10374 & w10395;
assign w10397 = ~w9350 & ~w10384;
assign w10398 = w10375 & w10397;
assign w10399 = w9350 & ~w10384;
assign w10400 = ~w10375 & w10399;
assign w10401 = ~w10398 & ~w10400;
assign w10402 = w9796 & w9904;
assign w10403 = w9773 & w10402;
assign w10404 = w9796 & ~w9904;
assign w10405 = ~w9773 & w10404;
assign w10406 = ~w10403 & ~w10405;
assign w10407 = w10401 & w10406;
assign w10408 = ~w10396 & w10407;
assign w10409 = w9909 & ~w10408;
assign w10410 = ~w9350 & w10375;
assign w10411 = w9808 & ~w9899;
assign w10412 = w9819 & w9898;
assign w10413 = ~w9808 & ~w10412;
assign w10414 = ~w10411 & ~w10413;
assign w10415 = ~w9351 & ~w10414;
assign w10416 = ~w10410 & w10415;
assign w10417 = ~w9819 & w9904;
assign w10418 = ~w10416 & ~w10417;
assign w10419 = (w9786 & ~w1913) | (w9786 & w34118) | (~w1913 & w34118);
assign w10420 = (w9780 & ~w1714) | (w9780 & w34119) | (~w1714 & w34119);
assign w10421 = (w9788 & ~w1807) | (w9788 & w34120) | (~w1807 & w34120);
assign w10422 = ~w10419 & ~w10420;
assign w10423 = ~w10421 & w10422;
assign w10424 = (w10423 & w4428) | (w10423 & w34121) | (w4428 & w34121);
assign w10425 = a_5 & w10424;
assign w10426 = (~w4428 & w34122) | (~w4428 & w34123) | (w34122 & w34123);
assign w10427 = ~w10425 & ~w10426;
assign w10428 = ~w9807 & w9898;
assign w10429 = ~w9806 & w10428;
assign w10430 = w9889 & ~w9898;
assign w10431 = ~w10429 & ~w10430;
assign w10432 = ~w2075 & w7192;
assign w10433 = (w7511 & ~w2235) | (w7511 & w34124) | (~w2235 & w34124);
assign w10434 = ~w2148 & w7489;
assign w10435 = ~w10433 & ~w10434;
assign w10436 = ~w10432 & w10435;
assign w10437 = (w10436 & ~w4962) | (w10436 & w34125) | (~w4962 & w34125);
assign w10438 = a_11 & ~w10437;
assign w10439 = (~w4962 & w34126) | (~w4962 & w34127) | (w34126 & w34127);
assign w10440 = ~w10438 & ~w10439;
assign w10441 = w9832 & ~w9861;
assign w10442 = ~w9841 & ~w10441;
assign w10443 = ~w9865 & w10442;
assign w10444 = w9841 & w10441;
assign w10445 = ~w9832 & w9862;
assign w10446 = w9307 & ~w10445;
assign w10447 = ~w10444 & w10446;
assign w10448 = ~w9829 & w10447;
assign w10449 = ~w10443 & ~w10448;
assign w10450 = ~w9831 & w9860;
assign w10451 = (w9855 & ~w10450) | (w9855 & w31723) | (~w10450 & w31723);
assign w10452 = ~w3403 & w6061;
assign w10453 = (w6304 & ~w3538) | (w6304 & w34128) | (~w3538 & w34128);
assign w10454 = ~w3475 & w6059;
assign w10455 = ~w10452 & ~w10453;
assign w10456 = ~w10454 & w10455;
assign w10457 = (w10456 & ~w5652) | (w10456 & w34129) | (~w5652 & w34129);
assign w10458 = a_17 & w10457;
assign w10459 = (w5652 & w34130) | (w5652 & w34131) | (w34130 & w34131);
assign w10460 = ~w10458 & ~w10459;
assign w10461 = w8045 & w8082;
assign w10462 = ~w8093 & ~w10461;
assign w10463 = w8065 & w8089;
assign w10464 = ~w3326 & w5816;
assign w10465 = ~w3196 & w5308;
assign w10466 = (w5818 & ~w3267) | (w5818 & w34132) | (~w3267 & w34132);
assign w10467 = ~w10465 & ~w10466;
assign w10468 = ~w10464 & w10467;
assign w10469 = (w10468 & w5903) | (w10468 & w34133) | (w5903 & w34133);
assign w10470 = a_20 & w10469;
assign w10471 = (~w5903 & w34134) | (~w5903 & w34135) | (w34134 & w34135);
assign w10472 = ~w10470 & ~w10471;
assign w10473 = w10463 & ~w10472;
assign w10474 = ~w10463 & w10472;
assign w10475 = ~w10473 & ~w10474;
assign w10476 = w10462 & w10475;
assign w10477 = ~w10462 & ~w10475;
assign w10478 = ~w10476 & ~w10477;
assign w10479 = w10460 & ~w10478;
assign w10480 = w10451 & w10479;
assign w10481 = w10460 & w10478;
assign w10482 = ~w10451 & w10481;
assign w10483 = ~w10480 & ~w10482;
assign w10484 = ~w10460 & w10478;
assign w10485 = w10451 & w10484;
assign w10486 = ~w10460 & ~w10478;
assign w10487 = ~w10451 & w10486;
assign w10488 = ~w10485 & ~w10487;
assign w10489 = w10483 & w10488;
assign w10490 = ~w2306 & w6446;
assign w10491 = ~w2393 & w6998;
assign w10492 = ~w3615 & w6996;
assign w10493 = ~w10490 & ~w10491;
assign w10494 = ~w10492 & w10493;
assign w10495 = (w10494 & ~w5463) | (w10494 & w34136) | (~w5463 & w34136);
assign w10496 = a_14 & ~w10495;
assign w10497 = (~w5463 & w34137) | (~w5463 & w34138) | (w34137 & w34138);
assign w10498 = ~w10496 & ~w10497;
assign w10499 = w10489 & w10498;
assign w10500 = ~w10489 & ~w10498;
assign w10501 = ~w10499 & ~w10500;
assign w10502 = w10449 & w10501;
assign w10503 = ~w10449 & ~w10501;
assign w10504 = ~w10502 & ~w10503;
assign w10505 = w10440 & w10504;
assign w10506 = ~w10440 & ~w10504;
assign w10507 = ~w10505 & ~w10506;
assign w10508 = (w8298 & ~w3658) | (w8298 & w34139) | (~w3658 & w34139);
assign w10509 = (w8277 & ~w3712) | (w8277 & w34140) | (~w3712 & w34140);
assign w10510 = (w8295 & ~w2005) | (w8295 & w34141) | (~w2005 & w34141);
assign w10511 = (w8278 & w4790) | (w8278 & w34142) | (w4790 & w34142);
assign w10512 = ~w10509 & ~w10510;
assign w10513 = ~w10508 & w10512;
assign w10514 = ~w10511 & w34143;
assign w10515 = (~a_8 & w10511) | (~a_8 & w34144) | (w10511 & w34144);
assign w10516 = ~w10514 & ~w10515;
assign w10517 = ~w9867 & ~w9879;
assign w10518 = w9830 & ~w10517;
assign w10519 = w9867 & ~w9879;
assign w10520 = ~w9830 & ~w10519;
assign w10521 = ~w10518 & ~w10520;
assign w10522 = w9799 & ~w10521;
assign w10523 = ~w9267 & w10522;
assign w10524 = w9823 & ~w9879;
assign w10525 = ~w9823 & w9879;
assign w10526 = ~w9870 & ~w10525;
assign w10527 = ~w10524 & ~w10526;
assign w10528 = ~w10523 & ~w10527;
assign w10529 = w10516 & ~w10528;
assign w10530 = ~w10516 & w10528;
assign w10531 = ~w10529 & ~w10530;
assign w10532 = w10507 & ~w10531;
assign w10533 = ~w10507 & w10531;
assign w10534 = ~w10532 & ~w10533;
assign w10535 = w10431 & w10534;
assign w10536 = ~w10431 & ~w10534;
assign w10537 = ~w10535 & ~w10536;
assign w10538 = ~w10427 & w10537;
assign w10539 = w10427 & ~w10537;
assign w10540 = ~w10538 & ~w10539;
assign w10541 = w10418 & ~w10540;
assign w10542 = ~w10418 & w10540;
assign w10543 = ~w10541 & ~w10542;
assign w10544 = w10409 & ~w10543;
assign w10545 = ~w10417 & w10537;
assign w10546 = ~w10416 & w10545;
assign w10547 = ~w10539 & ~w10546;
assign w10548 = ~w10541 & ~w10547;
assign w10549 = ~w10516 & ~w10537;
assign w10550 = ~w10546 & ~w10549;
assign w10551 = w10440 & ~w10504;
assign w10552 = w10528 & ~w10551;
assign w10553 = ~w10505 & ~w10528;
assign w10554 = ~w10552 & ~w10553;
assign w10555 = ~w10430 & ~w10554;
assign w10556 = ~w10429 & w10555;
assign w10557 = ~w10506 & ~w10528;
assign w10558 = ~w10440 & w10504;
assign w10559 = w10528 & ~w10558;
assign w10560 = ~w10557 & ~w10559;
assign w10561 = ~w10504 & ~w10528;
assign w10562 = ~w10489 & w10498;
assign w10563 = ~w10449 & w10562;
assign w10564 = w10449 & w10499;
assign w10565 = ~w10563 & ~w10564;
assign w10566 = (w10565 & w10528) | (w10565 & w31724) | (w10528 & w31724);
assign w10567 = (w8277 & ~w3658) | (w8277 & w34145) | (~w3658 & w34145);
assign w10568 = (w8298 & ~w2005) | (w8298 & w34146) | (~w2005 & w34146);
assign w10569 = (w8295 & ~w1913) | (w8295 & w34147) | (~w1913 & w34147);
assign w10570 = ~w10568 & ~w10569;
assign w10571 = ~w10567 & w10570;
assign w10572 = (w10571 & w4578) | (w10571 & w34148) | (w4578 & w34148);
assign w10573 = a_8 & ~w10572;
assign w10574 = (w4578 & w34149) | (w4578 & w34150) | (w34149 & w34150);
assign w10575 = ~w10573 & ~w10574;
assign w10576 = ~w10443 & w10488;
assign w10577 = w10483 & ~w10576;
assign w10578 = ~w9867 & w10483;
assign w10579 = w9830 & w10578;
assign w10580 = ~w10577 & ~w10579;
assign w10581 = w10451 & ~w10478;
assign w10582 = ~w10463 & ~w10472;
assign w10583 = ~w10462 & w10582;
assign w10584 = w10462 & w10473;
assign w10585 = ~w10583 & ~w10584;
assign w10586 = ~w10581 & w10585;
assign w10587 = ~w3403 & w6059;
assign w10588 = ~w2306 & w6304;
assign w10589 = (w6061 & ~w3538) | (w6061 & w34151) | (~w3538 & w34151);
assign w10590 = ~w10588 & ~w10589;
assign w10591 = ~w10587 & w10590;
assign w10592 = (w10591 & ~w5706) | (w10591 & w34152) | (~w5706 & w34152);
assign w10593 = a_17 & w10592;
assign w10594 = (w5706 & w34153) | (w5706 & w34154) | (w34153 & w34154);
assign w10595 = ~w10593 & ~w10594;
assign w10596 = ~w8096 & ~w10595;
assign w10597 = w8096 & w10595;
assign w10598 = ~w10596 & ~w10597;
assign w10599 = ~w3326 & w5818;
assign w10600 = (w5308 & ~w3267) | (w5308 & w34155) | (~w3267 & w34155);
assign w10601 = ~w3475 & w5816;
assign w10602 = ~w10599 & ~w10600;
assign w10603 = ~w10601 & w10602;
assign w10604 = (w10603 & ~w6108) | (w10603 & w34156) | (~w6108 & w34156);
assign w10605 = a_20 & w10604;
assign w10606 = (w6108 & w34157) | (w6108 & w34158) | (w34157 & w34158);
assign w10607 = ~w10605 & ~w10606;
assign w10608 = ~w8112 & w10607;
assign w10609 = w8112 & ~w10607;
assign w10610 = ~w10608 & ~w10609;
assign w10611 = w10598 & w10610;
assign w10612 = ~w10598 & ~w10610;
assign w10613 = ~w10611 & ~w10612;
assign w10614 = w10586 & w10613;
assign w10615 = ~w10586 & ~w10613;
assign w10616 = ~w10614 & ~w10615;
assign w10617 = ~w2075 & w6996;
assign w10618 = ~w2393 & w6446;
assign w10619 = ~w3615 & w6998;
assign w10620 = ~w10618 & ~w10619;
assign w10621 = ~w10617 & w10620;
assign w10622 = (w10621 & ~w5227) | (w10621 & w34159) | (~w5227 & w34159);
assign w10623 = a_14 & w10622;
assign w10624 = (w5227 & w34160) | (w5227 & w34161) | (w34160 & w34161);
assign w10625 = ~w10623 & ~w10624;
assign w10626 = w5103 & w9061;
assign w10627 = (w7511 & ~w3712) | (w7511 & w34162) | (~w3712 & w34162);
assign w10628 = ~w2148 & w7192;
assign w10629 = (w7489 & ~w2235) | (w7489 & w34163) | (~w2235 & w34163);
assign w10630 = ~w10628 & w34164;
assign w10631 = a_11 & w10630;
assign w10632 = ~a_11 & ~w10630;
assign w10633 = ~w10631 & ~w10632;
assign w10634 = (w10633 & ~w5103) | (w10633 & w34165) | (~w5103 & w34165);
assign w10635 = ~w10626 & ~w10634;
assign w10636 = w10625 & ~w10635;
assign w10637 = ~w10625 & w10635;
assign w10638 = ~w10636 & ~w10637;
assign w10639 = w10616 & ~w10638;
assign w10640 = ~w10616 & w10638;
assign w10641 = ~w10639 & ~w10640;
assign w10642 = w10580 & w10641;
assign w10643 = ~w10580 & ~w10641;
assign w10644 = ~w10642 & ~w10643;
assign w10645 = w10575 & ~w10644;
assign w10646 = ~w10575 & w10644;
assign w10647 = ~w10645 & ~w10646;
assign w10648 = w10566 & w10647;
assign w10649 = ~w10566 & ~w10647;
assign w10650 = ~w10648 & ~w10649;
assign w10651 = (~w10650 & w10556) | (~w10650 & w31725) | (w10556 & w31725);
assign w10652 = ~w10556 & w31726;
assign w10653 = ~w10651 & ~w10652;
assign w10654 = ~w3813 & w9788;
assign w10655 = (w9786 & ~w1714) | (w9786 & w34166) | (~w1714 & w34166);
assign w10656 = (w9780 & ~w1807) | (w9780 & w34167) | (~w1807 & w34167);
assign w10657 = w4508 & w9790;
assign w10658 = ~w10654 & w34168;
assign w10659 = ~w10657 & w34169;
assign w10660 = (~a_5 & w10657) | (~a_5 & w34170) | (w10657 & w34170);
assign w10661 = ~w10659 & ~w10660;
assign w10662 = w10653 & ~w10661;
assign w10663 = ~w10653 & w10661;
assign w10664 = ~w10662 & ~w10663;
assign w10665 = w10550 & w10664;
assign w10666 = ~w10550 & ~w10664;
assign w10667 = ~w10665 & ~w10666;
assign w10668 = ~w10548 & w10667;
assign w10669 = ~w10544 & w10668;
assign w10670 = ~w10661 & ~w10667;
assign w10671 = ~w10669 & ~w10670;
assign w10672 = ~w10566 & ~w10644;
assign w10673 = w10565 & w10644;
assign w10674 = ~w10561 & w10673;
assign w10675 = ~w10560 & ~w10674;
assign w10676 = ~w10672 & w10675;
assign w10677 = ~w10556 & w10676;
assign w10678 = w10575 & ~w10677;
assign w10679 = ~w10651 & w10678;
assign w10680 = ~w10549 & ~w10679;
assign w10681 = ~w10546 & w10680;
assign w10682 = w10653 & ~w10678;
assign w10683 = ~w10561 & w31727;
assign w10684 = w10635 & ~w10644;
assign w10685 = ~w10566 & w10684;
assign w10686 = ~w10683 & ~w10685;
assign w10687 = ~w10677 & w10686;
assign w10688 = w10616 & w10625;
assign w10689 = w10580 & w10688;
assign w10690 = ~w10616 & w10625;
assign w10691 = ~w10580 & w10690;
assign w10692 = ~w10689 & ~w10691;
assign w10693 = ~w10504 & w10692;
assign w10694 = ~w10528 & w10693;
assign w10695 = ~w10565 & ~w10625;
assign w10696 = w10565 & w10625;
assign w10697 = ~w10580 & ~w10616;
assign w10698 = w10580 & w10616;
assign w10699 = ~w10697 & ~w10698;
assign w10700 = ~w10696 & w10699;
assign w10701 = ~w10695 & ~w10700;
assign w10702 = ~w10694 & w10701;
assign w10703 = w4592 & w9456;
assign w10704 = (w8298 & ~w1913) | (w8298 & w34171) | (~w1913 & w34171);
assign w10705 = (w8277 & ~w2005) | (w8277 & w34172) | (~w2005 & w34172);
assign w10706 = (w8295 & ~w1714) | (w8295 & w34173) | (~w1714 & w34173);
assign w10707 = ~w10704 & ~w10705;
assign w10708 = w10707 & w34174;
assign w10709 = (~a_8 & ~w10707) | (~a_8 & w34175) | (~w10707 & w34175);
assign w10710 = ~w10708 & ~w10709;
assign w10711 = (w10710 & ~w4592) | (w10710 & w34176) | (~w4592 & w34176);
assign w10712 = ~w10703 & ~w10711;
assign w10713 = w10702 & ~w10712;
assign w10714 = ~w10702 & w10712;
assign w10715 = ~w10713 & ~w10714;
assign w10716 = (w7511 & ~w3658) | (w7511 & w34177) | (~w3658 & w34177);
assign w10717 = (w7192 & ~w2235) | (w7192 & w34178) | (~w2235 & w34178);
assign w10718 = (w7489 & ~w3712) | (w7489 & w34179) | (~w3712 & w34179);
assign w10719 = ~w10717 & ~w10718;
assign w10720 = ~w10716 & w10719;
assign w10721 = (w10720 & ~w4810) | (w10720 & w34180) | (~w4810 & w34180);
assign w10722 = a_11 & ~w10721;
assign w10723 = (~w4810 & w34181) | (~w4810 & w34182) | (w34181 & w34182);
assign w10724 = ~w10722 & ~w10723;
assign w10725 = ~w10595 & ~w10613;
assign w10726 = w10586 & w10725;
assign w10727 = ~w10595 & w10613;
assign w10728 = ~w10586 & w10727;
assign w10729 = ~w10726 & ~w10728;
assign w10730 = (w10729 & w10580) | (w10729 & w31728) | (w10580 & w31728);
assign w10731 = ~w8113 & ~w8114;
assign w10732 = ~w3475 & w5818;
assign w10733 = ~w3403 & w5816;
assign w10734 = ~w3326 & w5308;
assign w10735 = ~w10732 & ~w10733;
assign w10736 = ~w10734 & w10735;
assign w10737 = (w10736 & ~w5923) | (w10736 & w34183) | (~w5923 & w34183);
assign w10738 = a_20 & ~w10737;
assign w10739 = (~w5923 & w34184) | (~w5923 & w34185) | (w34184 & w34185);
assign w10740 = ~w10738 & ~w10739;
assign w10741 = (w6059 & ~w3538) | (w6059 & w34186) | (~w3538 & w34186);
assign w10742 = ~w2393 & w6304;
assign w10743 = ~w2306 & w6061;
assign w10744 = ~w10741 & ~w10742;
assign w10745 = ~w10743 & w10744;
assign w10746 = (w10745 & ~w5483) | (w10745 & w34187) | (~w5483 & w34187);
assign w10747 = a_17 & ~w10746;
assign w10748 = (~w5483 & w34188) | (~w5483 & w34189) | (w34188 & w34189);
assign w10749 = ~w10747 & ~w10748;
assign w10750 = ~w10740 & ~w10749;
assign w10751 = w7928 & w10750;
assign w10752 = w10740 & ~w10749;
assign w10753 = ~w7928 & w10752;
assign w10754 = ~w10751 & ~w10753;
assign w10755 = w10731 & ~w10754;
assign w10756 = w7928 & w10752;
assign w10757 = ~w7928 & w10750;
assign w10758 = ~w10756 & ~w10757;
assign w10759 = ~w10731 & ~w10758;
assign w10760 = ~w10755 & ~w10759;
assign w10761 = w10740 & w10749;
assign w10762 = w7928 & w10761;
assign w10763 = ~w10740 & w10749;
assign w10764 = ~w7928 & w10763;
assign w10765 = ~w10762 & ~w10764;
assign w10766 = w10731 & ~w10765;
assign w10767 = w7928 & w10763;
assign w10768 = ~w7928 & w10761;
assign w10769 = ~w10767 & ~w10768;
assign w10770 = ~w10731 & ~w10769;
assign w10771 = ~w10766 & ~w10770;
assign w10772 = w10760 & w10771;
assign w10773 = w8096 & ~w10608;
assign w10774 = w8112 & w10607;
assign w10775 = ~w8096 & ~w10774;
assign w10776 = ~w10773 & ~w10775;
assign w10777 = w8096 & ~w10609;
assign w10778 = ~w8112 & ~w10607;
assign w10779 = ~w8096 & ~w10778;
assign w10780 = ~w10777 & ~w10779;
assign w10781 = w10585 & ~w10780;
assign w10782 = ~w10776 & ~w10781;
assign w10783 = ~w10478 & ~w10776;
assign w10784 = w10451 & w10783;
assign w10785 = ~w10782 & ~w10784;
assign w10786 = w10772 & ~w10785;
assign w10787 = ~w10772 & w10785;
assign w10788 = ~w10786 & ~w10787;
assign w10789 = w5242 & w8564;
assign w10790 = ~w2148 & w6996;
assign w10791 = ~w3615 & w6446;
assign w10792 = ~w2075 & w6998;
assign w10793 = ~w10790 & ~w10791;
assign w10794 = w10793 & w34190;
assign w10795 = (~a_14 & ~w10793) | (~a_14 & w34191) | (~w10793 & w34191);
assign w10796 = ~w10794 & ~w10795;
assign w10797 = (w10796 & ~w5242) | (w10796 & w34192) | (~w5242 & w34192);
assign w10798 = ~w10789 & ~w10797;
assign w10799 = w10788 & ~w10798;
assign w10800 = ~w10788 & w10798;
assign w10801 = ~w10799 & ~w10800;
assign w10802 = w10730 & w10801;
assign w10803 = ~w10730 & ~w10801;
assign w10804 = ~w10802 & ~w10803;
assign w10805 = ~w10724 & w10804;
assign w10806 = w10724 & ~w10804;
assign w10807 = ~w10805 & ~w10806;
assign w10808 = w10715 & ~w10807;
assign w10809 = ~w10715 & w10807;
assign w10810 = ~w10808 & ~w10809;
assign w10811 = w10687 & w10810;
assign w10812 = ~w10687 & ~w10810;
assign w10813 = ~w10811 & ~w10812;
assign w10814 = ~w10682 & ~w10813;
assign w10815 = ~w10681 & w10814;
assign w10816 = (w9786 & ~w1807) | (w9786 & w34193) | (~w1807 & w34193);
assign w10817 = (w9788 & ~w1628) | (w9788 & w33993) | (~w1628 & w33993);
assign w10818 = ~w3813 & w9780;
assign w10819 = ~w10816 & ~w10817;
assign w10820 = ~w10818 & w10819;
assign w10821 = (w10820 & ~w4244) | (w10820 & w34194) | (~w4244 & w34194);
assign w10822 = a_5 & ~w10821;
assign w10823 = (~w4244 & w34195) | (~w4244 & w34196) | (w34195 & w34196);
assign w10824 = ~w10822 & ~w10823;
assign w10825 = w10815 & ~w10824;
assign w10826 = ~w10681 & ~w10682;
assign w10827 = w10813 & ~w10824;
assign w10828 = ~w10826 & w10827;
assign w10829 = ~w10825 & ~w10828;
assign w10830 = (w10813 & w10681) | (w10813 & w31729) | (w10681 & w31729);
assign w10831 = ~w10815 & w10824;
assign w10832 = ~w10830 & w10831;
assign w10833 = w10829 & ~w10832;
assign w10834 = w3 & ~w1397;
assign w10835 = ~a_0 & a_1;
assign w10836 = ~w1475 & w10835;
assign w10837 = a_0 & w2;
assign w10838 = ~w10834 & ~w10836;
assign w10839 = ~a_0 & ~a_1;
assign w10840 = (w10839 & ~w643) | (w10839 & w34198) | (~w643 & w34198);
assign w10841 = a_2 & ~w10840;
assign w10842 = (~w4056 & w34199) | (~w4056 & w34200) | (w34199 & w34200);
assign w10843 = (w4056 & w34201) | (w4056 & w34202) | (w34201 & w34202);
assign w10844 = ~w10842 & ~w10843;
assign w10845 = w10833 & w10844;
assign w10846 = w10671 & w10845;
assign w10847 = ~w10833 & w10844;
assign w10848 = ~w10671 & w10847;
assign w10849 = ~w10846 & ~w10848;
assign w10850 = w10272 & w10296;
assign w10851 = (w10300 & ~w10258) | (w10300 & w34203) | (~w10258 & w34203);
assign w10852 = ~w10850 & w10851;
assign w10853 = w10850 & ~w10851;
assign w10854 = ~w10852 & ~w10853;
assign w10855 = (w10835 & ~w3658) | (w10835 & w34204) | (~w3658 & w34204);
assign w10856 = (w3 & ~w2005) | (w3 & w34205) | (~w2005 & w34205);
assign w10857 = (w10837 & w4790) | (w10837 & w34206) | (w4790 & w34206);
assign w10858 = ~w10855 & ~w10856;
assign w10859 = (w10839 & ~w3712) | (w10839 & w34207) | (~w3712 & w34207);
assign w10860 = a_2 & ~w10859;
assign w10861 = ~w10857 & w34208;
assign w10862 = (a_2 & w10857) | (a_2 & w34209) | (w10857 & w34209);
assign w10863 = ~w10861 & ~w10862;
assign w10864 = w10854 & w10863;
assign w10865 = w10206 & ~w10211;
assign w10866 = ~w10206 & w10211;
assign w10867 = ~w10865 & ~w10866;
assign w10868 = w3 & ~w2075;
assign w10869 = ~w3615 & w10835;
assign w10870 = ~w10868 & ~w10869;
assign w10871 = (w10870 & ~w5227) | (w10870 & w34210) | (~w5227 & w34210);
assign w10872 = (a_2 & w2393) | (a_2 & w34211) | (w2393 & w34211);
assign w10873 = w10871 & ~w10872;
assign w10874 = (w5227 & w34212) | (w5227 & w34213) | (w34212 & w34213);
assign w10875 = ~w10873 & ~w10874;
assign w10876 = ~w10867 & ~w10875;
assign w10877 = w9980 & ~w9983;
assign w10878 = ~w10180 & ~w10186;
assign w10879 = (~w9998 & w10180) | (~w9998 & w34214) | (w10180 & w34214);
assign w10880 = ~w10877 & w10879;
assign w10881 = w10877 & ~w10879;
assign w10882 = ~w10880 & ~w10881;
assign w10883 = w3 & ~w2306;
assign w10884 = (w10835 & ~w3538) | (w10835 & w34215) | (~w3538 & w34215);
assign w10885 = ~w10883 & ~w10884;
assign w10886 = (w10885 & ~w5706) | (w10885 & w34216) | (~w5706 & w34216);
assign w10887 = (a_2 & w3403) | (a_2 & w34211) | (w3403 & w34211);
assign w10888 = w10886 & ~w10887;
assign w10889 = (w5706 & w34217) | (w5706 & w34218) | (w34217 & w34218);
assign w10890 = ~w10888 & ~w10889;
assign w10891 = ~w10882 & ~w10890;
assign w10892 = (a_5 & w10046) | (a_5 & w34219) | (w10046 & w34219);
assign w10893 = ~w10057 & w10892;
assign w10894 = w10057 & ~w10892;
assign w10895 = ~w10893 & ~w10894;
assign w10896 = (w10835 & ~w2766) | (w10835 & w34220) | (~w2766 & w34220);
assign w10897 = w3 & ~w2835;
assign w10898 = ~w10896 & ~w10897;
assign w10899 = (w10898 & ~w6733) | (w10898 & w31730) | (~w6733 & w31730);
assign w10900 = (w6733 & w34221) | (w6733 & w34222) | (w34221 & w34222);
assign w10901 = (a_2 & w2546) | (a_2 & w34211) | (w2546 & w34211);
assign w10902 = w10899 & ~w10901;
assign w10903 = ~w10902 & w34223;
assign w10904 = w10057 & w34224;
assign w10905 = ~w10059 & ~w10904;
assign w10906 = w10071 & ~w10905;
assign w10907 = ~w10071 & w10905;
assign w10908 = ~w10906 & ~w10907;
assign w10909 = a_2 & w10839;
assign w10910 = (w10909 & ~w2766) | (w10909 & w34225) | (~w2766 & w34225);
assign w10911 = w3 & ~w2917;
assign w10912 = ~w2835 & w10835;
assign w10913 = ~w10911 & ~w10912;
assign w10914 = (~w6784 & w34226) | (~w6784 & w34227) | (w34226 & w34227);
assign w10915 = (w6784 & w34228) | (w6784 & w34229) | (w34228 & w34229);
assign w10916 = ~w10914 & ~w10915;
assign w10917 = ~w10910 & ~w10916;
assign w10918 = ~w10908 & w10917;
assign w10919 = w10045 & ~w10050;
assign w10920 = ~w10051 & ~w10919;
assign w10921 = w3 & ~w2546;
assign w10922 = ~w2677 & w10835;
assign w10923 = ~w10921 & ~w10922;
assign w10924 = (w10923 & ~w6675) | (w10923 & w34230) | (~w6675 & w34230);
assign w10925 = a_2 & ~w10924;
assign w10926 = (w10839 & ~w2479) | (w10839 & w34231) | (~w2479 & w34231);
assign w10927 = a_2 & ~w10926;
assign w10928 = (~w6675 & w34232) | (~w6675 & w34233) | (w34232 & w34233);
assign w10929 = w3 & ~w2677;
assign w10930 = (~w10839 & ~w2479) | (~w10839 & w34234) | (~w2479 & w34234);
assign w10931 = w7970 & w10837;
assign w10932 = w2600 & w34235;
assign w10933 = ~w10929 & w34236;
assign w10934 = (~w10044 & w10931) | (~w10044 & w34237) | (w10931 & w34237);
assign w10935 = ~w10925 & w34238;
assign w10936 = ~w10920 & ~w10935;
assign w10937 = (~w10895 & w10902) | (~w10895 & w34239) | (w10902 & w34239);
assign w10938 = w10920 & w10935;
assign w10939 = ~w2677 & w10909;
assign w10940 = ~w2546 & w10835;
assign w10941 = (w3 & ~w2766) | (w3 & w34240) | (~w2766 & w34240);
assign w10942 = ~w10940 & ~w10941;
assign w10943 = (w10942 & ~w7625) | (w10942 & w34241) | (~w7625 & w34241);
assign w10944 = (~w7625 & w34242) | (~w7625 & w34243) | (w34242 & w34243);
assign w10945 = (~w10939 & w10943) | (~w10939 & w34244) | (w10943 & w34244);
assign w10946 = ~w10944 & w10945;
assign w10947 = ~w10938 & ~w10946;
assign w10948 = ~w10936 & ~w10937;
assign w10949 = ~w10947 & w10948;
assign w10950 = ~w10903 & ~w10918;
assign w10951 = ~w10949 & w10950;
assign w10952 = w10908 & ~w10917;
assign w10953 = w10072 & ~w10088;
assign w10954 = ~w10089 & ~w10953;
assign w10955 = ~w2835 & w10909;
assign w10956 = w3 & ~w3007;
assign w10957 = ~w2917 & w10835;
assign w10958 = ~w10956 & ~w10957;
assign w10959 = (w10958 & w6547) | (w10958 & w34245) | (w6547 & w34245);
assign w10960 = ~a_2 & ~w10959;
assign w10961 = (w6547 & w34246) | (w6547 & w34247) | (w34246 & w34247);
assign w10962 = (~w10955 & w10960) | (~w10955 & w34248) | (w10960 & w34248);
assign w10963 = w10954 & ~w10962;
assign w10964 = ~w10952 & ~w10963;
assign w10965 = ~w10951 & w10964;
assign w10966 = ~w10954 & w10962;
assign w10967 = ~w10965 & ~w10966;
assign w10968 = ~w10043 & ~w10091;
assign w10969 = ~w10092 & ~w10968;
assign w10970 = w3 & ~w3049;
assign w10971 = ~w3007 & w10835;
assign w10972 = ~w10970 & ~w10971;
assign w10973 = (w10972 & ~w6194) | (w10972 & w34249) | (~w6194 & w34249);
assign w10974 = (a_2 & w2917) | (a_2 & w34211) | (w2917 & w34211);
assign w10975 = w10973 & ~w10974;
assign w10976 = (w6194 & w34250) | (w6194 & w34251) | (w34250 & w34251);
assign w10977 = ~w10975 & ~w10976;
assign w10978 = ~w10969 & ~w10977;
assign w10979 = ~w10967 & ~w10978;
assign w10980 = w10969 & w10977;
assign w10981 = ~w10093 & w10121;
assign w10982 = w10093 & ~w10121;
assign w10983 = ~w10981 & ~w10982;
assign w10984 = w3 & ~w3139;
assign w10985 = ~w3049 & w10835;
assign w10986 = ~w10984 & ~w10985;
assign w10987 = (w10986 & w6505) | (w10986 & w34252) | (w6505 & w34252);
assign w10988 = (a_2 & w3007) | (a_2 & w34211) | (w3007 & w34211);
assign w10989 = w10987 & ~w10988;
assign w10990 = (~w6505 & w34253) | (~w6505 & w34254) | (w34253 & w34254);
assign w10991 = ~w10989 & ~w10990;
assign w10992 = (~w10980 & ~w10983) | (~w10980 & w34255) | (~w10983 & w34255);
assign w10993 = ~w10979 & w10992;
assign w10994 = ~w10983 & ~w10991;
assign w10995 = w3 & ~w3196;
assign w10996 = ~w3139 & w10835;
assign w10997 = ~w10995 & ~w10996;
assign w10998 = (w10997 & ~w6491) | (w10997 & w34256) | (~w6491 & w34256);
assign w10999 = (a_2 & w3049) | (a_2 & w34211) | (w3049 & w34211);
assign w11000 = w10998 & ~w10999;
assign w11001 = (w6491 & w34257) | (w6491 & w34258) | (w34257 & w34258);
assign w11002 = ~w11000 & ~w11001;
assign w11003 = (~w10119 & w10093) | (~w10119 & w34259) | (w10093 & w34259);
assign w11004 = ~w10105 & ~w10124;
assign w11005 = ~w11003 & w11004;
assign w11006 = w11003 & ~w11004;
assign w11007 = ~w11005 & ~w11006;
assign w11008 = ~w11002 & ~w11007;
assign w11009 = ~w10993 & ~w10994;
assign w11010 = ~w11008 & w11009;
assign w11011 = w11002 & w11007;
assign w11012 = ~w10026 & w10127;
assign w11013 = ~w10128 & ~w11012;
assign w11014 = (w3 & ~w3267) | (w3 & w34260) | (~w3267 & w34260);
assign w11015 = ~w3196 & w10835;
assign w11016 = w6222 & w34261;
assign w11017 = ~w11014 & ~w11015;
assign w11018 = ~w11016 & w11017;
assign w11019 = (a_2 & w3139) | (a_2 & w34211) | (w3139 & w34211);
assign w11020 = w11018 & ~w11019;
assign w11021 = (a_2 & w11016) | (a_2 & w34262) | (w11016 & w34262);
assign w11022 = ~w11020 & ~w11021;
assign w11023 = w11013 & w11022;
assign w11024 = ~w11011 & ~w11023;
assign w11025 = ~w11010 & w11024;
assign w11026 = ~w11013 & ~w11022;
assign w11027 = ~w10024 & ~w10128;
assign w11028 = w10142 & ~w10172;
assign w11029 = w11027 & ~w11028;
assign w11030 = ~w11027 & w11028;
assign w11031 = ~w11029 & ~w11030;
assign w11032 = w3 & ~w3326;
assign w11033 = (w10835 & ~w3267) | (w10835 & w34263) | (~w3267 & w34263);
assign w11034 = ~w11032 & ~w11033;
assign w11035 = (w11034 & w5903) | (w11034 & w34264) | (w5903 & w34264);
assign w11036 = (a_2 & w3196) | (a_2 & w34211) | (w3196 & w34211);
assign w11037 = w11035 & ~w11036;
assign w11038 = (~w5903 & w34265) | (~w5903 & w34266) | (w34265 & w34266);
assign w11039 = ~w11037 & ~w11038;
assign w11040 = (~w11026 & w11031) | (~w11026 & w34267) | (w11031 & w34267);
assign w11041 = ~w11025 & w11040;
assign w11042 = w11031 & w11039;
assign w11043 = (w10168 & w10144) | (w10168 & w34268) | (w10144 & w34268);
assign w11044 = ~w10174 & ~w11043;
assign w11045 = w3 & ~w3475;
assign w11046 = ~w3326 & w10835;
assign w11047 = ~w11045 & ~w11046;
assign w11048 = (w11047 & ~w6108) | (w11047 & w34269) | (~w6108 & w34269);
assign w11049 = (a_2 & w3268) | (a_2 & w34211) | (w3268 & w34211);
assign w11050 = w11048 & ~w11049;
assign w11051 = (w6108 & w34270) | (w6108 & w34271) | (w34270 & w34271);
assign w11052 = ~w11050 & ~w11051;
assign w11053 = w11044 & w11052;
assign w11054 = ~w11042 & ~w11053;
assign w11055 = ~w11041 & w11054;
assign w11056 = ~w11044 & ~w11052;
assign w11057 = w10176 & ~w10178;
assign w11058 = ~w10179 & ~w11057;
assign w11059 = w3 & ~w3403;
assign w11060 = ~w3475 & w10835;
assign w11061 = ~w11059 & ~w11060;
assign w11062 = (w11061 & ~w5923) | (w11061 & w34272) | (~w5923 & w34272);
assign w11063 = (a_2 & w3326) | (a_2 & w34211) | (w3326 & w34211);
assign w11064 = w11062 & ~w11063;
assign w11065 = (w5923 & w34273) | (w5923 & w34274) | (w34273 & w34274);
assign w11066 = ~w11064 & ~w11065;
assign w11067 = (~w11056 & w11058) | (~w11056 & w34275) | (w11058 & w34275);
assign w11068 = ~w11055 & w11067;
assign w11069 = ~w3403 & w10835;
assign w11070 = (w3 & ~w3538) | (w3 & w34276) | (~w3538 & w34276);
assign w11071 = ~w11069 & ~w11070;
assign w11072 = (w11071 & ~w5652) | (w11071 & w34277) | (~w5652 & w34277);
assign w11073 = (a_2 & w3475) | (a_2 & w34211) | (w3475 & w34211);
assign w11074 = w11072 & ~w11073;
assign w11075 = (w5652 & w34278) | (w5652 & w34279) | (w34278 & w34279);
assign w11076 = ~w11074 & ~w11075;
assign w11077 = w10186 & w11076;
assign w11078 = ~w10180 & w11077;
assign w11079 = w11058 & w11066;
assign w11080 = ~w10186 & w11076;
assign w11081 = w10180 & w11080;
assign w11082 = ~w11078 & ~w11079;
assign w11083 = ~w11081 & w11082;
assign w11084 = ~w11068 & w11083;
assign w11085 = w10180 & w10186;
assign w11086 = ~w10878 & ~w11085;
assign w11087 = ~w11076 & ~w11086;
assign w11088 = ~w11084 & ~w11087;
assign w11089 = ~w10891 & w11088;
assign w11090 = w10882 & w10890;
assign w11091 = ~w2306 & w10835;
assign w11092 = w3 & ~w2393;
assign w11093 = ~w11091 & ~w11092;
assign w11094 = (w11093 & ~w5483) | (w11093 & w34280) | (~w5483 & w34280);
assign w11095 = (a_2 & w3539) | (a_2 & w34211) | (w3539 & w34211);
assign w11096 = w11094 & ~w11095;
assign w11097 = (w5483 & w34281) | (w5483 & w34282) | (w34281 & w34282);
assign w11098 = ~w11096 & ~w11097;
assign w11099 = ~w10201 & ~w10203;
assign w11100 = w10189 & ~w11099;
assign w11101 = ~w10189 & w11099;
assign w11102 = ~w11100 & ~w11101;
assign w11103 = w11098 & w11102;
assign w11104 = ~w11090 & ~w11103;
assign w11105 = ~w11089 & w11104;
assign w11106 = (~w10203 & w10189) | (~w10203 & w34283) | (w10189 & w34283);
assign w11107 = ~w9965 & ~w11106;
assign w11108 = w3 & ~w3615;
assign w11109 = ~w2393 & w10835;
assign w11110 = ~w11108 & ~w11109;
assign w11111 = (w11110 & ~w5463) | (w11110 & w34284) | (~w5463 & w34284);
assign w11112 = (a_2 & w2306) | (a_2 & w34211) | (w2306 & w34211);
assign w11113 = w11111 & ~w11112;
assign w11114 = (w5463 & w34285) | (w5463 & w34286) | (w34285 & w34286);
assign w11115 = ~w11113 & ~w11114;
assign w11116 = w11107 & ~w11115;
assign w11117 = w9965 & ~w11115;
assign w11118 = w11106 & w11117;
assign w11119 = ~w11098 & ~w11102;
assign w11120 = ~w11118 & ~w11119;
assign w11121 = ~w11116 & w11120;
assign w11122 = ~w11105 & w11121;
assign w11123 = w9965 & w11106;
assign w11124 = ~w11107 & w11115;
assign w11125 = ~w11123 & w11124;
assign w11126 = ~w11122 & ~w11125;
assign w11127 = ~w10876 & ~w11126;
assign w11128 = (w9939 & ~w10206) | (w9939 & w34287) | (~w10206 & w34287);
assign w11129 = w9923 & w9945;
assign w11130 = ~w2075 & w10835;
assign w11131 = w3 & ~w2148;
assign w11132 = ~w11130 & ~w11131;
assign w11133 = (w11132 & ~w5242) | (w11132 & w34288) | (~w5242 & w34288);
assign w11134 = (a_2 & w3615) | (a_2 & w34211) | (w3615 & w34211);
assign w11135 = w11133 & ~w11134;
assign w11136 = (w5242 & w34289) | (w5242 & w34290) | (w34289 & w34290);
assign w11137 = ~w11135 & ~w11136;
assign w11138 = ~w11128 & w34291;
assign w11139 = w11129 & w11137;
assign w11140 = w11128 & w11139;
assign w11141 = w10867 & w10875;
assign w11142 = ~w11141 & w34292;
assign w11143 = ~w11127 & w11142;
assign w11144 = w10214 & w10231;
assign w11145 = ~w10232 & ~w11144;
assign w11146 = (w3 & ~w2235) | (w3 & w34293) | (~w2235 & w34293);
assign w11147 = ~w2148 & w10835;
assign w11148 = ~w11146 & ~w11147;
assign w11149 = (w11148 & ~w4962) | (w11148 & w34294) | (~w4962 & w34294);
assign w11150 = (a_2 & w2075) | (a_2 & w34211) | (w2075 & w34211);
assign w11151 = w11149 & ~w11150;
assign w11152 = (w4962 & w34295) | (w4962 & w34296) | (w34295 & w34296);
assign w11153 = ~w11151 & ~w11152;
assign w11154 = w11128 & w11129;
assign w11155 = (~w11137 & w11128) | (~w11137 & w34297) | (w11128 & w34297);
assign w11156 = ~w11154 & w11155;
assign w11157 = (~w11156 & w11145) | (~w11156 & w34298) | (w11145 & w34298);
assign w11158 = ~w11143 & w11157;
assign w11159 = ~w10232 & w10250;
assign w11160 = w10246 & w10257;
assign w11161 = (w3 & ~w3712) | (w3 & w34299) | (~w3712 & w34299);
assign w11162 = (w10835 & ~w2235) | (w10835 & w34300) | (~w2235 & w34300);
assign w11163 = ~w11161 & ~w11162;
assign w11164 = (w11163 & ~w5103) | (w11163 & w34301) | (~w5103 & w34301);
assign w11165 = (a_2 & w2148) | (a_2 & w34211) | (w2148 & w34211);
assign w11166 = w11164 & ~w11165;
assign w11167 = (w5103 & w34302) | (w5103 & w34303) | (w34302 & w34303);
assign w11168 = ~w11166 & ~w11167;
assign w11169 = ~w11159 & w34304;
assign w11170 = w11160 & w11168;
assign w11171 = w11159 & w11170;
assign w11172 = w11145 & w11153;
assign w11173 = ~w11171 & ~w11172;
assign w11174 = ~w11169 & w11173;
assign w11175 = ~w11158 & w11174;
assign w11176 = (w3 & ~w3658) | (w3 & w34305) | (~w3658 & w34305);
assign w11177 = (w10835 & ~w3712) | (w10835 & w34306) | (~w3712 & w34306);
assign w11178 = ~w11176 & ~w11177;
assign w11179 = (w11178 & ~w4810) | (w11178 & w34307) | (~w4810 & w34307);
assign w11180 = (a_2 & w2236) | (a_2 & w34211) | (w2236 & w34211);
assign w11181 = w11179 & ~w11180;
assign w11182 = (w4810 & w34308) | (w4810 & w34309) | (w34308 & w34309);
assign w11183 = ~w11181 & ~w11182;
assign w11184 = ~w10289 & ~w11183;
assign w11185 = w10258 & w11184;
assign w11186 = w10289 & ~w11183;
assign w11187 = ~w10258 & w11186;
assign w11188 = w10252 & w10257;
assign w11189 = (~w11168 & w11159) | (~w11168 & w34310) | (w11159 & w34310);
assign w11190 = ~w11188 & w11189;
assign w11191 = ~w11185 & ~w11187;
assign w11192 = ~w11190 & w11191;
assign w11193 = ~w11175 & w11192;
assign w11194 = ~w10258 & w10289;
assign w11195 = (w11183 & ~w10258) | (w11183 & w34311) | (~w10258 & w34311);
assign w11196 = ~w11194 & w11195;
assign w11197 = ~w11193 & ~w11196;
assign w11198 = ~w10864 & w11197;
assign w11199 = ~w10854 & ~w10863;
assign w11200 = w10303 & ~w10319;
assign w11201 = ~w10320 & ~w11200;
assign w11202 = (w3 & ~w1913) | (w3 & w34312) | (~w1913 & w34312);
assign w11203 = (w10835 & ~w2005) | (w10835 & w34313) | (~w2005 & w34313);
assign w11204 = ~w11202 & ~w11203;
assign w11205 = (w11204 & w4578) | (w11204 & w34314) | (w4578 & w34314);
assign w11206 = (a_2 & w3659) | (a_2 & w34211) | (w3659 & w34211);
assign w11207 = w11205 & ~w11206;
assign w11208 = (~w4578 & w34315) | (~w4578 & w34316) | (w34315 & w34316);
assign w11209 = ~w11207 & ~w11208;
assign w11210 = ~w11201 & ~w11209;
assign w11211 = ~w11199 & ~w11210;
assign w11212 = ~w11198 & w11211;
assign w11213 = ~w10320 & ~w10339;
assign w11214 = w10335 & w10345;
assign w11215 = (w10835 & ~w1913) | (w10835 & w34317) | (~w1913 & w34317);
assign w11216 = (w3 & ~w1714) | (w3 & w34318) | (~w1714 & w34318);
assign w11217 = ~w11215 & ~w11216;
assign w11218 = (w11217 & ~w4592) | (w11217 & w34319) | (~w4592 & w34319);
assign w11219 = (a_2 & w2006) | (a_2 & w34211) | (w2006 & w34211);
assign w11220 = w11218 & ~w11219;
assign w11221 = (w4592 & w34320) | (w4592 & w34321) | (w34320 & w34321);
assign w11222 = ~w11220 & ~w11221;
assign w11223 = ~w11213 & w34322;
assign w11224 = w11214 & w11222;
assign w11225 = w11213 & w11224;
assign w11226 = w11201 & w11209;
assign w11227 = ~w11225 & ~w11226;
assign w11228 = ~w11223 & w11227;
assign w11229 = ~w11212 & w11228;
assign w11230 = (w3 & ~w1807) | (w3 & w34323) | (~w1807 & w34323);
assign w11231 = (w10835 & ~w1714) | (w10835 & w34324) | (~w1714 & w34324);
assign w11232 = ~w11230 & ~w11231;
assign w11233 = (w11232 & w4428) | (w11232 & w34325) | (w4428 & w34325);
assign w11234 = (a_2 & w1914) | (a_2 & w34211) | (w1914 & w34211);
assign w11235 = w11233 & ~w11234;
assign w11236 = (~w4428 & w34326) | (~w4428 & w34327) | (w34326 & w34327);
assign w11237 = ~w11235 & ~w11236;
assign w11238 = w10373 & w31732;
assign w11239 = ~w10341 & w10345;
assign w11240 = ~w10372 & ~w11237;
assign w11241 = ~w11239 & w11240;
assign w11242 = w11213 & w11214;
assign w11243 = (~w11222 & w11213) | (~w11222 & w34328) | (w11213 & w34328);
assign w11244 = ~w11242 & w11243;
assign w11245 = ~w11238 & ~w11241;
assign w11246 = ~w11244 & w11245;
assign w11247 = ~w11229 & w11246;
assign w11248 = (~w10394 & ~w10373) | (~w10394 & w31733) | (~w10373 & w31733);
assign w11249 = w10389 & w10401;
assign w11250 = w3 & ~w3813;
assign w11251 = (w10835 & ~w1807) | (w10835 & w34329) | (~w1807 & w34329);
assign w11252 = ~w11250 & ~w11251;
assign w11253 = (w11252 & ~w4508) | (w11252 & w34330) | (~w4508 & w34330);
assign w11254 = (a_2 & w1715) | (a_2 & w34211) | (w1715 & w34211);
assign w11255 = w11253 & ~w11254;
assign w11256 = (w4508 & w34331) | (w4508 & w34332) | (w34331 & w34332);
assign w11257 = ~w11255 & ~w11256;
assign w11258 = w11249 & w11257;
assign w11259 = w11248 & w11258;
assign w11260 = ~w11249 & w11257;
assign w11261 = ~w11248 & w11260;
assign w11262 = ~w10372 & ~w11239;
assign w11263 = (w11237 & ~w10373) | (w11237 & w34333) | (~w10373 & w34333);
assign w11264 = ~w11262 & w11263;
assign w11265 = ~w11259 & ~w11261;
assign w11266 = ~w11264 & w11265;
assign w11267 = ~w11247 & w11266;
assign w11268 = ~w10396 & w10401;
assign w11269 = w9909 & w10406;
assign w11270 = ~w3813 & w10835;
assign w11271 = (w3 & ~w1628) | (w3 & w34318) | (~w1628 & w34318);
assign w11272 = ~w11270 & ~w11271;
assign w11273 = (w11272 & ~w4244) | (w11272 & w34334) | (~w4244 & w34334);
assign w11274 = (a_2 & w1808) | (a_2 & w34211) | (w1808 & w34211);
assign w11275 = w11273 & ~w11274;
assign w11276 = (w4244 & w34335) | (w4244 & w34336) | (w34335 & w34336);
assign w11277 = ~w11275 & ~w11276;
assign w11278 = ~w11268 & w31734;
assign w11279 = w11269 & ~w11277;
assign w11280 = w11268 & w11279;
assign w11281 = w11249 & ~w11257;
assign w11282 = ~w11248 & w11281;
assign w11283 = ~w11249 & ~w11257;
assign w11284 = w11248 & w11283;
assign w11285 = ~w11282 & ~w11284;
assign w11286 = ~w11280 & w11285;
assign w11287 = ~w11278 & w11286;
assign w11288 = ~w11267 & w11287;
assign w11289 = (w10835 & ~w1628) | (w10835 & w34324) | (~w1628 & w34324);
assign w11290 = (w3 & ~w643) | (w3 & w34337) | (~w643 & w34337);
assign w11291 = ~w11289 & ~w11290;
assign w11292 = (w11291 & ~w4224) | (w11291 & w34338) | (~w4224 & w34338);
assign w11293 = (a_2 & w3813) | (a_2 & w34211) | (w3813 & w34211);
assign w11294 = w11292 & ~w11293;
assign w11295 = (w4224 & w34339) | (w4224 & w34340) | (w34339 & w34340);
assign w11296 = ~w11294 & ~w11295;
assign w11297 = ~w10543 & w11296;
assign w11298 = w10409 & w11297;
assign w11299 = w10543 & w11296;
assign w11300 = ~w10409 & w11299;
assign w11301 = w11268 & w11269;
assign w11302 = (w11277 & w11268) | (w11277 & w31735) | (w11268 & w31735);
assign w11303 = ~w11301 & w11302;
assign w11304 = ~w11298 & ~w11300;
assign w11305 = ~w11303 & w11304;
assign w11306 = ~w11288 & w11305;
assign w11307 = (~w10548 & ~w10409) | (~w10548 & w31736) | (~w10409 & w31736);
assign w11308 = w3 & ~w1475;
assign w11309 = (w10835 & ~w643) | (w10835 & w34341) | (~w643 & w34341);
assign w11310 = ~w11308 & ~w11309;
assign w11311 = (w11310 & ~w4041) | (w11310 & w34342) | (~w4041 & w34342);
assign w11312 = (a_2 & w1629) | (a_2 & w34211) | (w1629 & w34211);
assign w11313 = w11311 & ~w11312;
assign w11314 = (w4041 & w34343) | (w4041 & w34344) | (w34343 & w34344);
assign w11315 = ~w11313 & ~w11314;
assign w11316 = ~w10667 & ~w11315;
assign w11317 = ~w11307 & w11316;
assign w11318 = ~w10548 & ~w11315;
assign w11319 = w10667 & w11318;
assign w11320 = ~w10544 & w11319;
assign w11321 = w10543 & ~w11296;
assign w11322 = w10409 & w11321;
assign w11323 = ~w10543 & ~w11296;
assign w11324 = ~w10409 & w11323;
assign w11325 = ~w11322 & ~w11324;
assign w11326 = ~w11320 & w11325;
assign w11327 = ~w11317 & w11326;
assign w11328 = ~w11306 & w11327;
assign w11329 = ~w10667 & ~w11307;
assign w11330 = ~w10669 & w11315;
assign w11331 = ~w11329 & w11330;
assign w11332 = ~w11328 & ~w11331;
assign w11333 = w10849 & w11332;
assign w11334 = ~w10833 & ~w10844;
assign w11335 = w10671 & w11334;
assign w11336 = w10833 & ~w10844;
assign w11337 = ~w10671 & w11336;
assign w11338 = ~w11335 & ~w11337;
assign w11339 = ~w10670 & ~w10832;
assign w11340 = ~w10669 & w11339;
assign w11341 = w10829 & ~w11340;
assign w11342 = ~w10724 & ~w10804;
assign w11343 = w10702 & ~w11342;
assign w11344 = ~w10702 & ~w10805;
assign w11345 = ~w11343 & ~w11344;
assign w11346 = w10724 & w10804;
assign w11347 = w10702 & ~w11346;
assign w11348 = ~w10702 & ~w10806;
assign w11349 = ~w11347 & ~w11348;
assign w11350 = ~w11345 & ~w11349;
assign w11351 = ~w10687 & ~w11350;
assign w11352 = w10687 & w11350;
assign w11353 = ~w11351 & ~w11352;
assign w11354 = w10712 & ~w11353;
assign w11355 = ~w10815 & ~w11354;
assign w11356 = ~w3813 & w9786;
assign w11357 = (w9788 & ~w643) | (w9788 & w34345) | (~w643 & w34345);
assign w11358 = (w9780 & ~w1628) | (w9780 & w34119) | (~w1628 & w34119);
assign w11359 = w4224 & w9790;
assign w11360 = ~w11356 & w34346;
assign w11361 = ~w11359 & w34347;
assign w11362 = (~a_5 & w11359) | (~a_5 & w34348) | (w11359 & w34348);
assign w11363 = ~w11361 & ~w11362;
assign w11364 = w10686 & ~w11349;
assign w11365 = ~w10677 & w11364;
assign w11366 = ~w11345 & ~w11365;
assign w11367 = w10760 & w10785;
assign w11368 = w10731 & w10758;
assign w11369 = ~w10731 & w10754;
assign w11370 = ~w11368 & ~w11369;
assign w11371 = ~w10785 & ~w11370;
assign w11372 = ~w11367 & ~w11371;
assign w11373 = w10771 & w10785;
assign w11374 = w10731 & w10769;
assign w11375 = ~w10731 & w10765;
assign w11376 = ~w11374 & ~w11375;
assign w11377 = ~w10785 & ~w11376;
assign w11378 = ~w11373 & ~w11377;
assign w11379 = ~w11372 & ~w11378;
assign w11380 = w10798 & w11379;
assign w11381 = w10730 & w11380;
assign w11382 = w10798 & ~w11379;
assign w11383 = ~w10730 & w11382;
assign w11384 = ~w11381 & ~w11383;
assign w11385 = ~w10702 & w10804;
assign w11386 = (w11384 & w10702) | (w11384 & w31737) | (w10702 & w31737);
assign w11387 = (w8277 & ~w1913) | (w8277 & w34349) | (~w1913 & w34349);
assign w11388 = (w8298 & ~w1714) | (w8298 & w34350) | (~w1714 & w34350);
assign w11389 = (w8295 & ~w1807) | (w8295 & w34351) | (~w1807 & w34351);
assign w11390 = ~w11387 & ~w11388;
assign w11391 = ~w11389 & w11390;
assign w11392 = (w11391 & w4428) | (w11391 & w34352) | (w4428 & w34352);
assign w11393 = a_8 & w11392;
assign w11394 = (~w4428 & w34353) | (~w4428 & w34354) | (w34353 & w34354);
assign w11395 = ~w11393 & ~w11394;
assign w11396 = w10729 & ~w11378;
assign w11397 = ~w11372 & ~w11396;
assign w11398 = ~w10616 & ~w11372;
assign w11399 = ~w10580 & w11398;
assign w11400 = ~w11397 & ~w11399;
assign w11401 = ~w7928 & w10731;
assign w11402 = w7928 & ~w10731;
assign w11403 = ~w11401 & ~w11402;
assign w11404 = ~w10740 & w11403;
assign w11405 = ~w10785 & ~w11404;
assign w11406 = w10740 & ~w11403;
assign w11407 = ~w11405 & ~w11406;
assign w11408 = ~w2306 & w6059;
assign w11409 = ~w2393 & w6061;
assign w11410 = ~w3615 & w6304;
assign w11411 = ~w11408 & ~w11409;
assign w11412 = ~w11410 & w11411;
assign w11413 = (w11412 & ~w5463) | (w11412 & w34355) | (~w5463 & w34355);
assign w11414 = a_17 & ~w11413;
assign w11415 = (~w5463 & w34356) | (~w5463 & w34357) | (w34356 & w34357);
assign w11416 = ~w11414 & ~w11415;
assign w11417 = (~a_20 & ~w5300) | (~a_20 & w34358) | (~w5300 & w34358);
assign w11418 = ~w3403 & w5818;
assign w11419 = (w5816 & ~w3538) | (w5816 & w34359) | (~w3538 & w34359);
assign w11420 = ~w3475 & w5308;
assign w11421 = ~w11418 & ~w11419;
assign w11422 = w11421 & w34360;
assign w11423 = (~a_20 & ~w11421) | (~a_20 & w34361) | (~w11421 & w34361);
assign w11424 = ~w11422 & ~w11423;
assign w11425 = w11421 & w34362;
assign w11426 = w5652 & w8311;
assign w11427 = (~w11424 & w5652) | (~w11424 & w34363) | (w5652 & w34363);
assign w11428 = ~w11426 & w11427;
assign w11429 = w7699 & ~w11428;
assign w11430 = ~w7699 & w11428;
assign w11431 = ~w11429 & ~w11430;
assign w11432 = ~w8130 & w11431;
assign w11433 = w8130 & ~w11431;
assign w11434 = ~w11432 & ~w11433;
assign w11435 = w8117 & w11434;
assign w11436 = ~w8117 & ~w11434;
assign w11437 = ~w11435 & ~w11436;
assign w11438 = w11416 & ~w11437;
assign w11439 = ~w11416 & w11437;
assign w11440 = ~w11438 & ~w11439;
assign w11441 = w11407 & w11440;
assign w11442 = ~w11407 & ~w11440;
assign w11443 = ~w11441 & ~w11442;
assign w11444 = ~w2075 & w6446;
assign w11445 = (w6996 & ~w2235) | (w6996 & w34364) | (~w2235 & w34364);
assign w11446 = ~w2148 & w6998;
assign w11447 = ~w11445 & ~w11446;
assign w11448 = ~w11444 & w11447;
assign w11449 = (w11448 & ~w4962) | (w11448 & w34365) | (~w4962 & w34365);
assign w11450 = a_14 & ~w11449;
assign w11451 = (~w4962 & w34366) | (~w4962 & w34367) | (w34366 & w34367);
assign w11452 = ~w11450 & ~w11451;
assign w11453 = (w7193 & w4790) | (w7193 & w34368) | (w4790 & w34368);
assign w11454 = (w7511 & ~w2005) | (w7511 & w34369) | (~w2005 & w34369);
assign w11455 = (w7192 & ~w3712) | (w7192 & w34370) | (~w3712 & w34370);
assign w11456 = (w7489 & ~w3658) | (w7489 & w34371) | (~w3658 & w34371);
assign w11457 = ~w11454 & ~w11455;
assign w11458 = ~w11456 & w11457;
assign w11459 = (a_11 & w11453) | (a_11 & w34372) | (w11453 & w34372);
assign w11460 = ~w11453 & w34373;
assign w11461 = ~w11459 & ~w11460;
assign w11462 = w11452 & w11461;
assign w11463 = ~w11452 & ~w11461;
assign w11464 = ~w11462 & ~w11463;
assign w11465 = w11443 & ~w11464;
assign w11466 = ~w11443 & w11464;
assign w11467 = ~w11465 & ~w11466;
assign w11468 = w11400 & w11467;
assign w11469 = ~w11400 & ~w11467;
assign w11470 = ~w11468 & ~w11469;
assign w11471 = w11395 & ~w11470;
assign w11472 = ~w11395 & w11470;
assign w11473 = ~w11471 & ~w11472;
assign w11474 = w11386 & ~w11473;
assign w11475 = ~w11386 & w11473;
assign w11476 = ~w11474 & ~w11475;
assign w11477 = w11366 & w11476;
assign w11478 = ~w11366 & ~w11476;
assign w11479 = ~w11477 & ~w11478;
assign w11480 = w11363 & ~w11479;
assign w11481 = ~w11363 & w11479;
assign w11482 = ~w11480 & ~w11481;
assign w11483 = w11355 & w11482;
assign w11484 = ~w11355 & ~w11482;
assign w11485 = ~w11483 & ~w11484;
assign w11486 = ~w1397 & w10835;
assign w11487 = (w3 & ~w1308) | (w3 & w34374) | (~w1308 & w34374);
assign w11488 = ~w11486 & ~w11487;
assign w11489 = (w11488 & ~w3834) | (w11488 & w34375) | (~w3834 & w34375);
assign w11490 = (a_2 & w1475) | (a_2 & w34211) | (w1475 & w34211);
assign w11491 = w11489 & ~w11490;
assign w11492 = (w3834 & w34376) | (w3834 & w34377) | (w34376 & w34377);
assign w11493 = ~w11491 & ~w11492;
assign w11494 = w11485 & ~w11493;
assign w11495 = ~w11485 & w11493;
assign w11496 = ~w11494 & ~w11495;
assign w11497 = ~w11341 & w11496;
assign w11498 = w11341 & ~w11496;
assign w11499 = ~w11497 & ~w11498;
assign w11500 = w11338 & w11499;
assign w11501 = ~w11333 & w11500;
assign w11502 = w11493 & ~w11499;
assign w11503 = ~w11363 & ~w11485;
assign w11504 = w11363 & w11483;
assign w11505 = ~w11355 & w11480;
assign w11506 = w10829 & ~w11505;
assign w11507 = ~w11504 & w11506;
assign w11508 = ~w11340 & w11507;
assign w11509 = ~w11503 & ~w11508;
assign w11510 = ~w11386 & ~w11470;
assign w11511 = w11384 & w11470;
assign w11512 = ~w11385 & w11511;
assign w11513 = ~w11510 & ~w11512;
assign w11514 = ~w11395 & ~w11513;
assign w11515 = w11366 & w11514;
assign w11516 = ~w11395 & w11513;
assign w11517 = ~w11366 & w11516;
assign w11518 = ~w11515 & ~w11517;
assign w11519 = ~w11354 & w11518;
assign w11520 = ~w10815 & w11519;
assign w11521 = w11395 & w11479;
assign w11522 = ~w11345 & ~w11512;
assign w11523 = ~w11510 & w11522;
assign w11524 = ~w11365 & w11523;
assign w11525 = w11461 & w11512;
assign w11526 = w11461 & ~w11470;
assign w11527 = ~w11386 & w11526;
assign w11528 = ~w11525 & ~w11527;
assign w11529 = ~w11524 & w11528;
assign w11530 = w11384 & ~w11452;
assign w11531 = ~w11400 & ~w11443;
assign w11532 = w11400 & w11443;
assign w11533 = ~w11531 & ~w11532;
assign w11534 = ~w11450 & w34378;
assign w11535 = w11379 & w11534;
assign w11536 = w10730 & w11535;
assign w11537 = ~w11379 & w11534;
assign w11538 = ~w10730 & w11537;
assign w11539 = ~w11536 & ~w11538;
assign w11540 = ~w11533 & w11539;
assign w11541 = ~w11530 & ~w11540;
assign w11542 = w11443 & ~w11452;
assign w11543 = w11400 & w11542;
assign w11544 = ~w11443 & ~w11452;
assign w11545 = ~w11400 & w11544;
assign w11546 = ~w11543 & ~w11545;
assign w11547 = w10804 & w11546;
assign w11548 = ~w10702 & w11547;
assign w11549 = ~w11541 & ~w11548;
assign w11550 = w11416 & w11443;
assign w11551 = ~w11531 & ~w11550;
assign w11552 = w8133 & w11428;
assign w11553 = w8117 & w11552;
assign w11554 = ~w8133 & w11428;
assign w11555 = ~w8117 & w11554;
assign w11556 = ~w11553 & ~w11555;
assign w11557 = w11437 & w11556;
assign w11558 = ~w11406 & w11556;
assign w11559 = ~w11405 & w11558;
assign w11560 = ~w11557 & ~w11559;
assign w11561 = (w6998 & ~w2235) | (w6998 & w34379) | (~w2235 & w34379);
assign w11562 = ~w2148 & w6446;
assign w11563 = (w6996 & ~w3712) | (w6996 & w34380) | (~w3712 & w34380);
assign w11564 = w5103 & w6447;
assign w11565 = ~w11562 & w34381;
assign w11566 = (a_14 & w11564) | (a_14 & w34382) | (w11564 & w34382);
assign w11567 = ~w11564 & w34383;
assign w11568 = ~w11566 & ~w11567;
assign w11569 = ~w11559 & w31738;
assign w11570 = (~w11568 & w11559) | (~w11568 & w31739) | (w11559 & w31739);
assign w11571 = ~w11569 & ~w11570;
assign w11572 = ~w8134 & ~w8135;
assign w11573 = ~w3403 & w5308;
assign w11574 = ~w2306 & w5816;
assign w11575 = (w5818 & ~w3538) | (w5818 & w34384) | (~w3538 & w34384);
assign w11576 = ~w11574 & ~w11575;
assign w11577 = ~w11573 & w11576;
assign w11578 = (w11577 & ~w5706) | (w11577 & w34385) | (~w5706 & w34385);
assign w11579 = a_20 & w11578;
assign w11580 = (w5706 & w34386) | (w5706 & w34387) | (w34386 & w34387);
assign w11581 = ~w11579 & ~w11580;
assign w11582 = ~w8157 & w31740;
assign w11583 = ~w8150 & w11582;
assign w11584 = ~w8139 & w11581;
assign w11585 = w8149 & w11584;
assign w11586 = (w11581 & w8157) | (w11581 & w31741) | (w8157 & w31741);
assign w11587 = ~w11585 & ~w11586;
assign w11588 = ~w11583 & w11587;
assign w11589 = ~w11572 & w11588;
assign w11590 = w11572 & ~w11588;
assign w11591 = ~w11589 & ~w11590;
assign w11592 = ~w2075 & w6304;
assign w11593 = ~w3615 & w6061;
assign w11594 = ~w2393 & w6059;
assign w11595 = ~w11593 & ~w11594;
assign w11596 = ~w11592 & w11595;
assign w11597 = (w11596 & ~w5227) | (w11596 & w34388) | (~w5227 & w34388);
assign w11598 = a_17 & ~w11597;
assign w11599 = (~w5227 & w34389) | (~w5227 & w34390) | (w34389 & w34390);
assign w11600 = ~w11598 & ~w11599;
assign w11601 = w11591 & ~w11600;
assign w11602 = ~w11591 & w11600;
assign w11603 = ~w11601 & ~w11602;
assign w11604 = w11571 & ~w11603;
assign w11605 = ~w11571 & w11603;
assign w11606 = ~w11604 & ~w11605;
assign w11607 = w11551 & w11606;
assign w11608 = ~w11551 & ~w11606;
assign w11609 = ~w11607 & ~w11608;
assign w11610 = ~w11549 & ~w11609;
assign w11611 = w11549 & w11609;
assign w11612 = ~w11610 & ~w11611;
assign w11613 = (w7192 & ~w3658) | (w7192 & w34391) | (~w3658 & w34391);
assign w11614 = (w7489 & ~w2005) | (w7489 & w34392) | (~w2005 & w34392);
assign w11615 = (w7511 & ~w1913) | (w7511 & w34393) | (~w1913 & w34393);
assign w11616 = ~w11614 & ~w11615;
assign w11617 = ~w11613 & w11616;
assign w11618 = (w11617 & w4578) | (w11617 & w34394) | (w4578 & w34394);
assign w11619 = a_11 & ~w11618;
assign w11620 = (w4578 & w34395) | (w4578 & w34396) | (w34395 & w34396);
assign w11621 = ~w11619 & ~w11620;
assign w11622 = w4508 & w9456;
assign w11623 = (w8298 & ~w1807) | (w8298 & w34397) | (~w1807 & w34397);
assign w11624 = (w8277 & ~w1714) | (w8277 & w34398) | (~w1714 & w34398);
assign w11625 = ~w3813 & w8295;
assign w11626 = ~w11623 & ~w11624;
assign w11627 = ~w11625 & w11626;
assign w11628 = a_8 & w11627;
assign w11629 = ~a_8 & ~w11627;
assign w11630 = ~w11628 & ~w11629;
assign w11631 = (w11630 & ~w4508) | (w11630 & w34399) | (~w4508 & w34399);
assign w11632 = ~w11622 & ~w11631;
assign w11633 = w11621 & ~w11632;
assign w11634 = ~w11621 & w11632;
assign w11635 = ~w11633 & ~w11634;
assign w11636 = w11612 & ~w11635;
assign w11637 = ~w11612 & w11635;
assign w11638 = ~w11636 & ~w11637;
assign w11639 = w11529 & w11638;
assign w11640 = ~w11529 & ~w11638;
assign w11641 = ~w11639 & ~w11640;
assign w11642 = ~w11521 & ~w11641;
assign w11643 = ~w11520 & w11642;
assign w11644 = ~w1475 & w9788;
assign w11645 = (w9786 & ~w1628) | (w9786 & w34166) | (~w1628 & w34166);
assign w11646 = (w9780 & ~w643) | (w9780 & w34400) | (~w643 & w34400);
assign w11647 = ~w11645 & ~w11646;
assign w11648 = ~w11644 & w11647;
assign w11649 = (w11648 & ~w4041) | (w11648 & w34401) | (~w4041 & w34401);
assign w11650 = a_5 & w11649;
assign w11651 = (w4041 & w34402) | (w4041 & w34403) | (w34402 & w34403);
assign w11652 = ~w11650 & ~w11651;
assign w11653 = w11643 & w11652;
assign w11654 = ~w11520 & ~w11521;
assign w11655 = w11641 & w11652;
assign w11656 = ~w11654 & w11655;
assign w11657 = ~w11653 & ~w11656;
assign w11658 = w11641 & ~w11652;
assign w11659 = w11654 & w11658;
assign w11660 = ~w11641 & ~w11652;
assign w11661 = ~w11654 & w11660;
assign w11662 = ~w11659 & ~w11661;
assign w11663 = w11657 & w11662;
assign w11664 = (w3 & ~w3904) | (w3 & w34404) | (~w3904 & w34404);
assign w11665 = (w10835 & ~w1308) | (w10835 & w34405) | (~w1308 & w34405);
assign w11666 = ~w11664 & ~w11665;
assign w11667 = (w11666 & ~w3964) | (w11666 & w34406) | (~w3964 & w34406);
assign w11668 = (a_2 & w1397) | (a_2 & w34211) | (w1397 & w34211);
assign w11669 = w11667 & ~w11668;
assign w11670 = (w3964 & w34407) | (w3964 & w34408) | (w34407 & w34408);
assign w11671 = ~w11669 & ~w11670;
assign w11672 = w11663 & w11671;
assign w11673 = w11509 & w11672;
assign w11674 = ~w11663 & w11671;
assign w11675 = ~w11509 & w11674;
assign w11676 = ~w11673 & ~w11675;
assign w11677 = ~w11502 & w11676;
assign w11678 = ~w11501 & w11677;
assign w11679 = ~w11663 & ~w11671;
assign w11680 = w11509 & w11679;
assign w11681 = w11663 & ~w11671;
assign w11682 = ~w11509 & w11681;
assign w11683 = ~w11680 & ~w11682;
assign w11684 = w11485 & w11657;
assign w11685 = w11341 & w11684;
assign w11686 = ~w11503 & w11662;
assign w11687 = w11657 & ~w11686;
assign w11688 = ~w11685 & ~w11687;
assign w11689 = (w10835 & ~w3904) | (w10835 & w34409) | (~w3904 & w34409);
assign w11690 = w3 & ~w3958;
assign w11691 = ~w11689 & ~w11690;
assign w11692 = (w11691 & ~w3943) | (w11691 & w34410) | (~w3943 & w34410);
assign w11693 = (a_2 & w1323) | (a_2 & w34211) | (w1323 & w34211);
assign w11694 = w11692 & ~w11693;
assign w11695 = (w3943 & w34411) | (w3943 & w34412) | (w34411 & w34412);
assign w11696 = ~w11694 & ~w11695;
assign w11697 = w11632 & w11641;
assign w11698 = ~w11643 & ~w11697;
assign w11699 = ~w1397 & w9788;
assign w11700 = (w9786 & ~w643) | (w9786 & w34413) | (~w643 & w34413);
assign w11701 = ~w1475 & w9780;
assign w11702 = ~w11699 & ~w11700;
assign w11703 = (a_5 & ~w11702) | (a_5 & w34414) | (~w11702 & w34414);
assign w11704 = w4056 & w9790;
assign w11705 = w11702 & w34415;
assign w11706 = ~w11704 & w11705;
assign w11707 = (~w11703 & ~w4056) | (~w11703 & w34416) | (~w4056 & w34416);
assign w11708 = ~w11706 & w11707;
assign w11709 = ~w11612 & ~w11621;
assign w11710 = ~w11609 & w11621;
assign w11711 = w11549 & w11710;
assign w11712 = w11609 & w11621;
assign w11713 = ~w11549 & w11712;
assign w11714 = ~w11711 & ~w11713;
assign w11715 = w11528 & w11714;
assign w11716 = ~w11524 & w11715;
assign w11717 = ~w11709 & ~w11716;
assign w11718 = w11560 & ~w11601;
assign w11719 = ~w11591 & ~w11600;
assign w11720 = ~w11560 & ~w11719;
assign w11721 = ~w11718 & ~w11720;
assign w11722 = w11560 & ~w11602;
assign w11723 = w11591 & w11600;
assign w11724 = ~w11560 & ~w11723;
assign w11725 = ~w11722 & ~w11724;
assign w11726 = ~w11721 & ~w11725;
assign w11727 = w11568 & w11726;
assign w11728 = w11551 & w11727;
assign w11729 = w11568 & ~w11726;
assign w11730 = ~w11551 & w11729;
assign w11731 = ~w11728 & ~w11730;
assign w11732 = (w11731 & w11549) | (w11731 & w31742) | (w11549 & w31742);
assign w11733 = ~w11550 & ~w11725;
assign w11734 = ~w11531 & w11733;
assign w11735 = ~w11721 & ~w11734;
assign w11736 = (w7489 & ~w1913) | (w7489 & w34417) | (~w1913 & w34417);
assign w11737 = (w7192 & ~w2005) | (w7192 & w34418) | (~w2005 & w34418);
assign w11738 = (w7511 & ~w1714) | (w7511 & w34419) | (~w1714 & w34419);
assign w11739 = ~w11736 & ~w11737;
assign w11740 = ~w11738 & w11739;
assign w11741 = (w11740 & ~w4592) | (w11740 & w34420) | (~w4592 & w34420);
assign w11742 = a_11 & w11741;
assign w11743 = (w4592 & w34421) | (w4592 & w34422) | (w34421 & w34422);
assign w11744 = ~w11742 & ~w11743;
assign w11745 = ~w11734 & w31743;
assign w11746 = (w11744 & w11734) | (w11744 & w31744) | (w11734 & w31744);
assign w11747 = ~w11745 & ~w11746;
assign w11748 = (w6996 & ~w3658) | (w6996 & w34423) | (~w3658 & w34423);
assign w11749 = (w6998 & ~w3712) | (w6998 & w34424) | (~w3712 & w34424);
assign w11750 = (w6446 & ~w2235) | (w6446 & w34425) | (~w2235 & w34425);
assign w11751 = ~w11749 & ~w11750;
assign w11752 = ~w11748 & w11751;
assign w11753 = (w11752 & ~w4810) | (w11752 & w34426) | (~w4810 & w34426);
assign w11754 = a_14 & ~w11753;
assign w11755 = (~w4810 & w34427) | (~w4810 & w34428) | (w34427 & w34428);
assign w11756 = ~w11754 & ~w11755;
assign w11757 = ~w11560 & w11591;
assign w11758 = w11581 & ~w11591;
assign w11759 = ~w11757 & ~w11758;
assign w11760 = ~w2306 & w5818;
assign w11761 = ~w2393 & w5816;
assign w11762 = (w5308 & ~w3538) | (w5308 & w34429) | (~w3538 & w34429);
assign w11763 = ~w11760 & ~w11761;
assign w11764 = ~w11762 & w11763;
assign w11765 = (w11764 & ~w5483) | (w11764 & w34430) | (~w5483 & w34430);
assign w11766 = a_20 & ~w11765;
assign w11767 = (~w5483 & w34431) | (~w5483 & w34432) | (w34431 & w34432);
assign w11768 = ~w11766 & ~w11767;
assign w11769 = w5242 & w8391;
assign w11770 = ~w3615 & w6059;
assign w11771 = ~w2148 & w6304;
assign w11772 = ~w2075 & w6061;
assign w11773 = ~w11770 & ~w11771;
assign w11774 = w11773 & w34433;
assign w11775 = (~a_17 & ~w11773) | (~a_17 & w34434) | (~w11773 & w34434);
assign w11776 = ~w11774 & ~w11775;
assign w11777 = (w11776 & ~w5242) | (w11776 & w34435) | (~w5242 & w34435);
assign w11778 = ~w11769 & ~w11777;
assign w11779 = ~w11768 & ~w11778;
assign w11780 = w11768 & w11778;
assign w11781 = ~w11779 & ~w11780;
assign w11782 = (w8178 & w8152) | (w8178 & w31745) | (w8152 & w31745);
assign w11783 = ~w8152 & w31746;
assign w11784 = ~w11782 & ~w11783;
assign w11785 = w11781 & ~w11784;
assign w11786 = ~w11781 & w11784;
assign w11787 = ~w11785 & ~w11786;
assign w11788 = w11759 & w11787;
assign w11789 = ~w11759 & ~w11787;
assign w11790 = ~w11788 & ~w11789;
assign w11791 = w11756 & w11790;
assign w11792 = ~w11756 & ~w11790;
assign w11793 = ~w11791 & ~w11792;
assign w11794 = w4244 & w8278;
assign w11795 = ~w3813 & w8298;
assign w11796 = (w8277 & ~w1807) | (w8277 & w34436) | (~w1807 & w34436);
assign w11797 = (w8295 & ~w1628) | (w8295 & w34173) | (~w1628 & w34173);
assign w11798 = ~w11795 & w34437;
assign w11799 = ~w11794 & w34438;
assign w11800 = (a_8 & w11794) | (a_8 & w34439) | (w11794 & w34439);
assign w11801 = ~w11799 & ~w11800;
assign w11802 = w11793 & ~w11801;
assign w11803 = ~w11793 & w11801;
assign w11804 = ~w11802 & ~w11803;
assign w11805 = w11747 & ~w11804;
assign w11806 = ~w11747 & w11804;
assign w11807 = ~w11805 & ~w11806;
assign w11808 = w11732 & ~w11807;
assign w11809 = ~w11732 & w11807;
assign w11810 = ~w11808 & ~w11809;
assign w11811 = w11717 & w11810;
assign w11812 = ~w11717 & ~w11810;
assign w11813 = ~w11811 & ~w11812;
assign w11814 = w11708 & ~w11813;
assign w11815 = ~w11708 & w11813;
assign w11816 = ~w11814 & ~w11815;
assign w11817 = w11698 & w11816;
assign w11818 = ~w11698 & ~w11816;
assign w11819 = ~w11817 & ~w11818;
assign w11820 = w11696 & ~w11819;
assign w11821 = ~w11696 & w11819;
assign w11822 = ~w11820 & ~w11821;
assign w11823 = w11688 & w11822;
assign w11824 = ~w11688 & ~w11822;
assign w11825 = ~w11823 & ~w11824;
assign w11826 = w11683 & ~w11825;
assign w11827 = ~w11678 & w11826;
assign w11828 = w11688 & ~w11819;
assign w11829 = ~w11708 & w11819;
assign w11830 = (~w11829 & ~w11688) | (~w11829 & w31747) | (~w11688 & w31747);
assign w11831 = ~w3958 & w10835;
assign w11832 = (~w11831 & ~w4073) | (~w11831 & w34440) | (~w4073 & w34440);
assign w11833 = (a_2 & w3906) | (a_2 & w34211) | (w3906 & w34211);
assign w11834 = w11832 & ~w11833;
assign w11835 = (w4073 & w34441) | (w4073 & w34442) | (w34441 & w34442);
assign w11836 = ~w11834 & ~w11835;
assign w11837 = w11747 & ~w11793;
assign w11838 = ~w11747 & w11793;
assign w11839 = ~w11837 & ~w11838;
assign w11840 = w11732 & w11839;
assign w11841 = ~w11732 & ~w11839;
assign w11842 = ~w11840 & ~w11841;
assign w11843 = w11801 & w11842;
assign w11844 = w11717 & w11843;
assign w11845 = w11801 & ~w11842;
assign w11846 = ~w11717 & w11845;
assign w11847 = ~w11844 & ~w11846;
assign w11848 = w11813 & w11847;
assign w11849 = ~w11697 & w11847;
assign w11850 = ~w11643 & w11849;
assign w11851 = ~w11848 & ~w11850;
assign w11852 = ~w1397 & w9780;
assign w11853 = ~w1475 & w9786;
assign w11854 = (w9788 & ~w1308) | (w9788 & w34443) | (~w1308 & w34443);
assign w11855 = ~w11852 & ~w11853;
assign w11856 = ~w11854 & w11855;
assign w11857 = (w11856 & ~w3834) | (w11856 & w34444) | (~w3834 & w34444);
assign w11858 = a_5 & ~w11857;
assign w11859 = (~w3834 & w34445) | (~w3834 & w34446) | (w34445 & w34446);
assign w11860 = ~w11858 & ~w11859;
assign w11861 = ~w11716 & w31748;
assign w11862 = ~w11744 & w11842;
assign w11863 = ~w11861 & ~w11862;
assign w11864 = ~w11735 & ~w11790;
assign w11865 = ~w11735 & w31749;
assign w11866 = w11735 & w11791;
assign w11867 = w11731 & ~w11866;
assign w11868 = ~w11865 & w11867;
assign w11869 = ~w11610 & w11868;
assign w11870 = w11735 & w11790;
assign w11871 = (~w11756 & w11735) | (~w11756 & w34447) | (w11735 & w34447);
assign w11872 = ~w11870 & w11871;
assign w11873 = ~w11869 & ~w11872;
assign w11874 = ~w11778 & w11790;
assign w11875 = ~w11864 & ~w11874;
assign w11876 = ~w11768 & ~w11784;
assign w11877 = w11768 & w11784;
assign w11878 = (~w11877 & w11757) | (~w11877 & w31750) | (w11757 & w31750);
assign w11879 = ~w11876 & ~w11878;
assign w11880 = (~w8179 & w8152) | (~w8179 & w31751) | (w8152 & w31751);
assign w11881 = w8194 & ~w11880;
assign w11882 = ~w8196 & ~w11881;
assign w11883 = ~w2306 & w5308;
assign w11884 = ~w2393 & w5818;
assign w11885 = ~w3615 & w5816;
assign w11886 = ~w11883 & ~w11884;
assign w11887 = ~w11885 & w11886;
assign w11888 = (w11887 & ~w5463) | (w11887 & w34448) | (~w5463 & w34448);
assign w11889 = a_20 & ~w11888;
assign w11890 = (~w5463 & w34449) | (~w5463 & w34450) | (w34449 & w34450);
assign w11891 = ~w11889 & ~w11890;
assign w11892 = ~w11882 & w11891;
assign w11893 = w11882 & ~w11891;
assign w11894 = ~w11892 & ~w11893;
assign w11895 = ~w2075 & w6059;
assign w11896 = (w6304 & ~w2235) | (w6304 & w34451) | (~w2235 & w34451);
assign w11897 = ~w2148 & w6061;
assign w11898 = ~w11896 & ~w11897;
assign w11899 = ~w11895 & w11898;
assign w11900 = (w11899 & ~w4962) | (w11899 & w34452) | (~w4962 & w34452);
assign w11901 = a_17 & ~w11900;
assign w11902 = (~w4962 & w34453) | (~w4962 & w34454) | (w34453 & w34454);
assign w11903 = ~w11901 & ~w11902;
assign w11904 = (w6998 & ~w3658) | (w6998 & w34455) | (~w3658 & w34455);
assign w11905 = (w6996 & ~w2005) | (w6996 & w34456) | (~w2005 & w34456);
assign w11906 = (w6446 & ~w3712) | (w6446 & w34457) | (~w3712 & w34457);
assign w11907 = (w6447 & w4790) | (w6447 & w34458) | (w4790 & w34458);
assign w11908 = ~w11905 & ~w11906;
assign w11909 = ~w11904 & w11908;
assign w11910 = (a_14 & w11907) | (a_14 & w34459) | (w11907 & w34459);
assign w11911 = ~w11907 & w34460;
assign w11912 = ~w11910 & ~w11911;
assign w11913 = w11903 & ~w11912;
assign w11914 = ~w11903 & w11912;
assign w11915 = ~w11913 & ~w11914;
assign w11916 = w11894 & ~w11915;
assign w11917 = ~w11894 & w11915;
assign w11918 = ~w11916 & ~w11917;
assign w11919 = w11879 & ~w11918;
assign w11920 = ~w11879 & w11918;
assign w11921 = ~w11919 & ~w11920;
assign w11922 = w11875 & w11921;
assign w11923 = ~w11875 & ~w11921;
assign w11924 = ~w11922 & ~w11923;
assign w11925 = w11873 & ~w11924;
assign w11926 = ~w11873 & w11924;
assign w11927 = ~w11925 & ~w11926;
assign w11928 = (w7511 & ~w1807) | (w7511 & w34461) | (~w1807 & w34461);
assign w11929 = (w7489 & ~w1714) | (w7489 & w34462) | (~w1714 & w34462);
assign w11930 = (w7192 & ~w1913) | (w7192 & w34463) | (~w1913 & w34463);
assign w11931 = ~w11928 & ~w11929;
assign w11932 = ~w11930 & w11931;
assign w11933 = (w11932 & w4428) | (w11932 & w34464) | (w4428 & w34464);
assign w11934 = a_11 & ~w11933;
assign w11935 = (w4428 & w34465) | (w4428 & w34466) | (w34465 & w34466);
assign w11936 = ~w11934 & ~w11935;
assign w11937 = ~w3813 & w8277;
assign w11938 = (w8298 & ~w1628) | (w8298 & w34350) | (~w1628 & w34350);
assign w11939 = (w8295 & ~w643) | (w8295 & w34467) | (~w643 & w34467);
assign w11940 = w4224 & w8278;
assign w11941 = ~w11937 & w34468;
assign w11942 = (a_8 & w11940) | (a_8 & w34469) | (w11940 & w34469);
assign w11943 = ~w11940 & w34470;
assign w11944 = ~w11942 & ~w11943;
assign w11945 = ~w11936 & w11944;
assign w11946 = w11936 & ~w11944;
assign w11947 = ~w11945 & ~w11946;
assign w11948 = w11927 & ~w11947;
assign w11949 = ~w11927 & w11947;
assign w11950 = ~w11948 & ~w11949;
assign w11951 = w11863 & w11950;
assign w11952 = ~w11863 & ~w11950;
assign w11953 = ~w11951 & ~w11952;
assign w11954 = w11860 & ~w11953;
assign w11955 = ~w11860 & w11953;
assign w11956 = ~w11954 & ~w11955;
assign w11957 = w11851 & w11956;
assign w11958 = ~w11851 & ~w11956;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = w11836 & w11959;
assign w11961 = ~w11830 & w11960;
assign w11962 = (w11836 & ~w11819) | (w11836 & w31752) | (~w11819 & w31752);
assign w11963 = ~w11959 & w11962;
assign w11964 = ~w11828 & w11963;
assign w11965 = w11688 & ~w11820;
assign w11966 = w11696 & w11819;
assign w11967 = ~w11688 & ~w11966;
assign w11968 = ~w11965 & ~w11967;
assign w11969 = ~w11964 & ~w11968;
assign w11970 = ~w11961 & w11969;
assign w11971 = ~w11827 & w11970;
assign w11972 = ~w11836 & w11959;
assign w11973 = w11830 & ~w11972;
assign w11974 = ~w11836 & ~w11959;
assign w11975 = ~w11830 & ~w11974;
assign w11976 = ~w11973 & ~w11975;
assign w11977 = ~w11971 & ~w11976;
assign w11978 = w11851 & ~w11953;
assign w11979 = ~w11851 & w11953;
assign w11980 = ~w11978 & ~w11979;
assign w11981 = w11860 & w11980;
assign w11982 = ~w11860 & ~w11980;
assign w11983 = ~w11829 & ~w11982;
assign w11984 = ~w11828 & w11983;
assign w11985 = w11944 & w11953;
assign w11986 = ~w11978 & ~w11985;
assign w11987 = (w9780 & ~w1308) | (w9780 & w34471) | (~w1308 & w34471);
assign w11988 = (w9788 & ~w3904) | (w9788 & w34472) | (~w3904 & w34472);
assign w11989 = ~w1397 & w9786;
assign w11990 = ~w11987 & ~w11989;
assign w11991 = ~w11988 & w11990;
assign w11992 = (w11991 & ~w3964) | (w11991 & w34473) | (~w3964 & w34473);
assign w11993 = a_5 & ~w11992;
assign w11994 = (~w3964 & w34474) | (~w3964 & w34475) | (w34474 & w34475);
assign w11995 = (w3828 & w34476) | (w3828 & w34477) | (w34476 & w34477);
assign w11996 = (a_2 & w3958) | (a_2 & w34211) | (w3958 & w34211);
assign w11997 = ~w11995 & w11996;
assign w11998 = a_1 & w11995;
assign w11999 = ~w11997 & ~w11998;
assign w12000 = ~w11993 & w34478;
assign w12001 = (w11999 & w11993) | (w11999 & w34479) | (w11993 & w34479);
assign w12002 = ~w12000 & ~w12001;
assign w12003 = ~w11927 & ~w11936;
assign w12004 = w11924 & w11936;
assign w12005 = w11873 & ~w12004;
assign w12006 = ~w11924 & w11936;
assign w12007 = ~w11873 & ~w12006;
assign w12008 = ~w12005 & ~w12007;
assign w12009 = ~w11862 & ~w12008;
assign w12010 = ~w11861 & w12009;
assign w12011 = ~w12003 & ~w12010;
assign w12012 = w11912 & w11924;
assign w12013 = ~w11925 & ~w12012;
assign w12014 = ~w1475 & w8295;
assign w12015 = (w8277 & ~w1628) | (w8277 & w34398) | (~w1628 & w34398);
assign w12016 = (w8298 & ~w643) | (w8298 & w34480) | (~w643 & w34480);
assign w12017 = ~w12015 & ~w12016;
assign w12018 = ~w12014 & w12017;
assign w12019 = (w12018 & ~w4041) | (w12018 & w34481) | (~w4041 & w34481);
assign w12020 = a_8 & w12019;
assign w12021 = (w4041 & w34482) | (w4041 & w34483) | (w34482 & w34483);
assign w12022 = ~w12020 & ~w12021;
assign w12023 = w11879 & w11894;
assign w12024 = ~w11879 & ~w11894;
assign w12025 = ~w12023 & ~w12024;
assign w12026 = ~w11903 & ~w12025;
assign w12027 = w11903 & w12025;
assign w12028 = (~w12026 & w11875) | (~w12026 & w31753) | (w11875 & w31753);
assign w12029 = (~w11892 & ~w11879) | (~w11892 & w32442) | (~w11879 & w32442);
assign w12030 = ~w3813 & w7511;
assign w12031 = (w7192 & ~w1714) | (w7192 & w34484) | (~w1714 & w34484);
assign w12032 = (w7489 & ~w1807) | (w7489 & w34485) | (~w1807 & w34485);
assign w12033 = w4508 & w7193;
assign w12034 = ~w12030 & w34486;
assign w12035 = (a_11 & w12033) | (a_11 & w34487) | (w12033 & w34487);
assign w12036 = ~w12033 & w34488;
assign w12037 = ~w12035 & ~w12036;
assign w12038 = ~w2075 & w5816;
assign w12039 = ~w3615 & w5818;
assign w12040 = ~w2393 & w5308;
assign w12041 = ~w12039 & ~w12040;
assign w12042 = ~w12038 & w12041;
assign w12043 = (w12042 & ~w5227) | (w12042 & w34489) | (~w5227 & w34489);
assign w12044 = a_20 & ~w12043;
assign w12045 = (~w5227 & w34490) | (~w5227 & w34491) | (w34490 & w34491);
assign w12046 = ~w12044 & ~w12045;
assign w12047 = ~w8214 & w12046;
assign w12048 = w8214 & ~w12046;
assign w12049 = ~w12047 & ~w12048;
assign w12050 = w8198 & w12049;
assign w12051 = ~w8198 & ~w12049;
assign w12052 = ~w12050 & ~w12051;
assign w12053 = (w6061 & ~w2235) | (w6061 & w34492) | (~w2235 & w34492);
assign w12054 = ~w2148 & w6059;
assign w12055 = (w6304 & ~w3712) | (w6304 & w34493) | (~w3712 & w34493);
assign w12056 = w5103 & w6063;
assign w12057 = ~w12054 & w34494;
assign w12058 = (a_17 & w12056) | (a_17 & w34495) | (w12056 & w34495);
assign w12059 = ~w12056 & w34496;
assign w12060 = ~w12058 & ~w12059;
assign w12061 = (w6446 & ~w3658) | (w6446 & w34497) | (~w3658 & w34497);
assign w12062 = (w6998 & ~w2005) | (w6998 & w34498) | (~w2005 & w34498);
assign w12063 = (w6996 & ~w1913) | (w6996 & w34499) | (~w1913 & w34499);
assign w12064 = ~w12062 & ~w12063;
assign w12065 = ~w12061 & w12064;
assign w12066 = (w12065 & w4578) | (w12065 & w34500) | (w4578 & w34500);
assign w12067 = a_14 & ~w12066;
assign w12068 = (w4578 & w34501) | (w4578 & w34502) | (w34501 & w34502);
assign w12069 = ~w12067 & ~w12068;
assign w12070 = w12060 & w12069;
assign w12071 = ~w12060 & ~w12069;
assign w12072 = ~w12070 & ~w12071;
assign w12073 = w12052 & w12072;
assign w12074 = ~w12052 & ~w12072;
assign w12075 = ~w12073 & ~w12074;
assign w12076 = w12037 & ~w12075;
assign w12077 = ~w12037 & w12075;
assign w12078 = ~w12076 & ~w12077;
assign w12079 = w12029 & ~w12078;
assign w12080 = ~w12029 & w12078;
assign w12081 = ~w12079 & ~w12080;
assign w12082 = w12028 & w12081;
assign w12083 = ~w12028 & ~w12081;
assign w12084 = ~w12082 & ~w12083;
assign w12085 = w12022 & ~w12084;
assign w12086 = ~w12022 & w12084;
assign w12087 = ~w12085 & ~w12086;
assign w12088 = w12013 & ~w12087;
assign w12089 = ~w12013 & w12087;
assign w12090 = ~w12088 & ~w12089;
assign w12091 = w12011 & w12090;
assign w12092 = ~w12011 & ~w12090;
assign w12093 = ~w12091 & ~w12092;
assign w12094 = w12002 & w12093;
assign w12095 = ~w12002 & ~w12093;
assign w12096 = ~w12094 & ~w12095;
assign w12097 = w11986 & w12096;
assign w12098 = ~w11986 & ~w12096;
assign w12099 = ~w12097 & ~w12098;
assign w12100 = (w12099 & w11984) | (w12099 & w31754) | (w11984 & w31754);
assign w12101 = ~w11985 & ~w12093;
assign w12102 = ~w11978 & w12101;
assign w12103 = w12022 & w12093;
assign w12104 = ~w12102 & ~w12103;
assign w12105 = ~w12029 & w12075;
assign w12106 = w12029 & ~w12075;
assign w12107 = ~w12105 & ~w12106;
assign w12108 = w12028 & w12107;
assign w12109 = ~w12028 & ~w12107;
assign w12110 = ~w12108 & ~w12109;
assign w12111 = (w12110 & w11925) | (w12110 & w31755) | (w11925 & w31755);
assign w12112 = ~w11925 & w31756;
assign w12113 = ~w12111 & ~w12112;
assign w12114 = ~w12037 & ~w12113;
assign w12115 = w12011 & ~w12114;
assign w12116 = ~w11925 & w34503;
assign w12117 = (w12084 & w11925) | (w12084 & w34504) | (w11925 & w34504);
assign w12118 = w12037 & ~w12116;
assign w12119 = ~w12117 & w12118;
assign w12120 = (~w12119 & ~w12011) | (~w12119 & w34505) | (~w12011 & w34505);
assign w12121 = (w9780 & ~w3904) | (w9780 & w34506) | (~w3904 & w34506);
assign w12122 = (w9786 & ~w1308) | (w9786 & w34507) | (~w1308 & w34507);
assign w12123 = ~w3958 & w9788;
assign w12124 = ~w12122 & ~w12123;
assign w12125 = ~w12121 & w12124;
assign w12126 = (w12125 & ~w3943) | (w12125 & w34508) | (~w3943 & w34508);
assign w12127 = a_5 & w12126;
assign w12128 = (w3943 & w34509) | (w3943 & w34510) | (w34509 & w34510);
assign w12129 = ~w12127 & ~w12128;
assign w12130 = ~w12052 & w12060;
assign w12131 = w12052 & ~w12060;
assign w12132 = ~w12130 & ~w12131;
assign w12133 = w12029 & w12132;
assign w12134 = ~w12029 & ~w12132;
assign w12135 = ~w12133 & ~w12134;
assign w12136 = ~w12028 & w12135;
assign w12137 = w12028 & ~w12135;
assign w12138 = ~w12136 & ~w12137;
assign w12139 = w12069 & ~w12138;
assign w12140 = ~w12111 & ~w12139;
assign w12141 = ~w12060 & ~w12135;
assign w12142 = (~w12141 & w12028) | (~w12141 & w34511) | (w12028 & w34511);
assign w12143 = ~w1397 & w8295;
assign w12144 = ~w1475 & w8298;
assign w12145 = (w8277 & ~w643) | (w8277 & w34512) | (~w643 & w34512);
assign w12146 = ~w12143 & ~w12145;
assign w12147 = ~w12144 & w12146;
assign w12148 = (w12147 & ~w4056) | (w12147 & w34513) | (~w4056 & w34513);
assign w12149 = ~a_8 & w12148;
assign w12150 = (w4056 & w34514) | (w4056 & w34515) | (w34514 & w34515);
assign w12151 = ~w12149 & ~w12150;
assign w12152 = ~w12046 & ~w12052;
assign w12153 = ~w11892 & w12052;
assign w12154 = (~w12152 & w12023) | (~w12152 & w32443) | (w12023 & w32443);
assign w12155 = w4244 & w7193;
assign w12156 = ~w3813 & w7489;
assign w12157 = (w7192 & ~w1807) | (w7192 & w34516) | (~w1807 & w34516);
assign w12158 = (w7511 & ~w1628) | (w7511 & w34419) | (~w1628 & w34419);
assign w12159 = ~w12156 & w34517;
assign w12160 = (a_11 & w12155) | (a_11 & w34518) | (w12155 & w34518);
assign w12161 = ~w12155 & w34519;
assign w12162 = ~w12160 & ~w12161;
assign w12163 = ~w7907 & ~w8216;
assign w12164 = ~w8217 & ~w12163;
assign w12165 = (w6304 & ~w3658) | (w6304 & w34520) | (~w3658 & w34520);
assign w12166 = (w6061 & ~w3712) | (w6061 & w34521) | (~w3712 & w34521);
assign w12167 = (w6059 & ~w2235) | (w6059 & w34522) | (~w2235 & w34522);
assign w12168 = ~w12166 & ~w12167;
assign w12169 = ~w12165 & w12168;
assign w12170 = (w12169 & ~w4810) | (w12169 & w34523) | (~w4810 & w34523);
assign w12171 = a_17 & ~w12170;
assign w12172 = (~w4810 & w34524) | (~w4810 & w34525) | (w34524 & w34525);
assign w12173 = ~w12171 & ~w12172;
assign w12174 = w4592 & w8564;
assign w12175 = (w6998 & ~w1913) | (w6998 & w34526) | (~w1913 & w34526);
assign w12176 = (w6446 & ~w2005) | (w6446 & w34527) | (~w2005 & w34527);
assign w12177 = (w6996 & ~w1714) | (w6996 & w33658) | (~w1714 & w33658);
assign w12178 = ~w12175 & ~w12176;
assign w12179 = w12178 & w34528;
assign w12180 = (~a_14 & ~w12178) | (~a_14 & w34529) | (~w12178 & w34529);
assign w12181 = ~w12179 & ~w12180;
assign w12182 = (w12181 & ~w4592) | (w12181 & w34530) | (~w4592 & w34530);
assign w12183 = ~w12174 & ~w12182;
assign w12184 = w12173 & ~w12183;
assign w12185 = ~w12173 & w12183;
assign w12186 = ~w12184 & ~w12185;
assign w12187 = w12164 & w12186;
assign w12188 = ~w12164 & ~w12186;
assign w12189 = ~w12187 & ~w12188;
assign w12190 = w12162 & ~w12189;
assign w12191 = ~w12162 & w12189;
assign w12192 = ~w12190 & ~w12191;
assign w12193 = w12154 & w12192;
assign w12194 = ~w12154 & ~w12192;
assign w12195 = ~w12193 & ~w12194;
assign w12196 = w12151 & ~w12195;
assign w12197 = ~w12151 & w12195;
assign w12198 = ~w12196 & ~w12197;
assign w12199 = w12142 & ~w12198;
assign w12200 = ~w12142 & w12198;
assign w12201 = ~w12199 & ~w12200;
assign w12202 = w12140 & w12201;
assign w12203 = ~w12140 & ~w12201;
assign w12204 = ~w12202 & ~w12203;
assign w12205 = w12129 & ~w12204;
assign w12206 = ~w12129 & w12204;
assign w12207 = ~w12205 & ~w12206;
assign w12208 = w12120 & w12207;
assign w12209 = ~w12120 & ~w12207;
assign w12210 = ~w12208 & ~w12209;
assign w12211 = w12104 & w12210;
assign w12212 = ~w12104 & ~w12210;
assign w12213 = ~w12211 & ~w12212;
assign w12214 = ~w11986 & w12094;
assign w12215 = (~w12000 & ~w12102) | (~w12000 & w31757) | (~w12102 & w31757);
assign w12216 = ~w12214 & w12215;
assign w12217 = w12213 & ~w12216;
assign w12218 = ~w12129 & ~w12210;
assign w12219 = ~w12211 & ~w12218;
assign w12220 = ~w12115 & w31758;
assign w12221 = (w9786 & ~w3904) | (w9786 & w34531) | (~w3904 & w34531);
assign w12222 = ~w3958 & w9780;
assign w12223 = ~w12221 & ~w12222;
assign w12224 = (w12223 & ~w4073) | (w12223 & w34532) | (~w4073 & w34532);
assign w12225 = a_5 & ~w12224;
assign w12226 = (~w4073 & w34533) | (~w4073 & w34534) | (w34533 & w34534);
assign w12227 = ~w12225 & ~w12226;
assign w12228 = (~w12227 & ~w12204) | (~w12227 & w34535) | (~w12204 & w34535);
assign w12229 = ~w12220 & w12228;
assign w12230 = (~w12204 & w12115) | (~w12204 & w31759) | (w12115 & w31759);
assign w12231 = (w12227 & ~w12204) | (w12227 & w34536) | (~w12204 & w34536);
assign w12232 = ~w12230 & w12231;
assign w12233 = ~w12229 & ~w12232;
assign w12234 = ~w1397 & w8298;
assign w12235 = ~w1475 & w8277;
assign w12236 = (w8295 & ~w1308) | (w8295 & w34537) | (~w1308 & w34537);
assign w12237 = ~w12234 & ~w12235;
assign w12238 = ~w12236 & w12237;
assign w12239 = (w12238 & ~w3834) | (w12238 & w34538) | (~w3834 & w34538);
assign w12240 = a_8 & ~w12239;
assign w12241 = (~w3834 & w34539) | (~w3834 & w34540) | (w34539 & w34540);
assign w12242 = ~w12240 & ~w12241;
assign w12243 = ~w8223 & w8232;
assign w12244 = ~w8233 & ~w12243;
assign w12245 = (~w12023 & w34541) | (~w12023 & w34542) | (w34541 & w34542);
assign w12246 = (w12023 & w34543) | (w12023 & w34544) | (w34543 & w34544);
assign w12247 = ~w12173 & ~w12246;
assign w12248 = ~w12245 & ~w12247;
assign w12249 = w12244 & w12248;
assign w12250 = ~w12244 & ~w12248;
assign w12251 = ~w12249 & ~w12250;
assign w12252 = (w6446 & ~w1913) | (w6446 & w34545) | (~w1913 & w34545);
assign w12253 = (w6998 & ~w1714) | (w6998 & w33585) | (~w1714 & w33585);
assign w12254 = (w6996 & ~w1807) | (w6996 & w34546) | (~w1807 & w34546);
assign w12255 = ~w12252 & ~w12253;
assign w12256 = ~w12254 & w12255;
assign w12257 = (w12256 & w4428) | (w12256 & w34547) | (w4428 & w34547);
assign w12258 = a_14 & w12257;
assign w12259 = (~w4428 & w34548) | (~w4428 & w34549) | (w34548 & w34549);
assign w12260 = ~w12258 & ~w12259;
assign w12261 = w12251 & ~w12260;
assign w12262 = ~w12251 & w12260;
assign w12263 = ~w12261 & ~w12262;
assign w12264 = w12154 & w12189;
assign w12265 = ~w12154 & ~w12189;
assign w12266 = ~w12264 & ~w12265;
assign w12267 = w12183 & w12266;
assign w12268 = ~w12141 & ~w12266;
assign w12269 = (~w12267 & w12136) | (~w12267 & w32444) | (w12136 & w32444);
assign w12270 = ~w3813 & w7192;
assign w12271 = (w7489 & ~w1628) | (w7489 & w34462) | (~w1628 & w34462);
assign w12272 = (w7511 & ~w643) | (w7511 & w34550) | (~w643 & w34550);
assign w12273 = w4224 & w7193;
assign w12274 = ~w12270 & w34551;
assign w12275 = (a_11 & w12273) | (a_11 & w34552) | (w12273 & w34552);
assign w12276 = ~w12273 & w34553;
assign w12277 = ~w12275 & ~w12276;
assign w12278 = ~w12269 & w12277;
assign w12279 = w12269 & ~w12277;
assign w12280 = ~w12278 & ~w12279;
assign w12281 = w12263 & w12280;
assign w12282 = ~w12263 & ~w12280;
assign w12283 = ~w12281 & ~w12282;
assign w12284 = w12142 & ~w12195;
assign w12285 = ~w12142 & w12195;
assign w12286 = ~w12284 & ~w12285;
assign w12287 = ~w12111 & w34554;
assign w12288 = ~w12162 & w12286;
assign w12289 = ~w12287 & ~w12288;
assign w12290 = w12283 & w12289;
assign w12291 = ~w12283 & ~w12289;
assign w12292 = ~w12290 & ~w12291;
assign w12293 = w12242 & ~w12292;
assign w12294 = ~w12242 & w12292;
assign w12295 = ~w12293 & ~w12294;
assign w12296 = w12233 & w12295;
assign w12297 = ~w12233 & ~w12295;
assign w12298 = ~w12296 & ~w12297;
assign w12299 = ~w12219 & w12298;
assign w12300 = ~w12217 & ~w12299;
assign w12301 = ~w12100 & w12300;
assign w12302 = ~w11977 & w12301;
assign w12303 = ~w1397 & w7511;
assign w12304 = ~w1475 & w7489;
assign w12305 = (w7192 & ~w643) | (w7192 & w34555) | (~w643 & w34555);
assign w12306 = ~w12303 & ~w12305;
assign w12307 = ~w12304 & w12306;
assign w12308 = (w12307 & ~w4056) | (w12307 & w34556) | (~w4056 & w34556);
assign w12309 = a_11 & ~w12308;
assign w12310 = (~w4056 & w34557) | (~w4056 & w34558) | (w34557 & w34558);
assign w12311 = ~w12309 & ~w12310;
assign w12312 = (~w12249 & ~w12251) | (~w12249 & w34559) | (~w12251 & w34559);
assign w12313 = ~w8235 & ~w8236;
assign w12314 = w8244 & w12313;
assign w12315 = ~w8244 & ~w12313;
assign w12316 = ~w12314 & ~w12315;
assign w12317 = ~w12312 & w12316;
assign w12318 = w12312 & ~w12316;
assign w12319 = ~w12317 & ~w12318;
assign w12320 = ~w1475 & w7511;
assign w12321 = (w7192 & ~w1628) | (w7192 & w34484) | (~w1628 & w34484);
assign w12322 = (w7489 & ~w643) | (w7489 & w34560) | (~w643 & w34560);
assign w12323 = ~w12321 & ~w12322;
assign w12324 = ~w12320 & w12323;
assign w12325 = (w12324 & ~w4041) | (w12324 & w34561) | (~w4041 & w34561);
assign w12326 = a_11 & w12325;
assign w12327 = (w4041 & w34562) | (w4041 & w34563) | (w34562 & w34563);
assign w12328 = ~w12326 & ~w12327;
assign w12329 = w12319 & ~w12328;
assign w12330 = (~w12317 & ~w12319) | (~w12317 & w34564) | (~w12319 & w34564);
assign w12331 = ~w12311 & w12330;
assign w12332 = w12311 & ~w12330;
assign w12333 = ~w12331 & ~w12332;
assign w12334 = ~w8247 & ~w8248;
assign w12335 = w8250 & w12334;
assign w12336 = ~w8250 & ~w12334;
assign w12337 = ~w12335 & ~w12336;
assign w12338 = w12333 & w12337;
assign w12339 = ~w12333 & ~w12337;
assign w12340 = ~w12338 & ~w12339;
assign w12341 = (~w12278 & ~w12280) | (~w12278 & w34565) | (~w12280 & w34565);
assign w12342 = ~w1397 & w8277;
assign w12343 = (w8295 & ~w3904) | (w8295 & w34566) | (~w3904 & w34566);
assign w12344 = (w8298 & ~w1308) | (w8298 & w34567) | (~w1308 & w34567);
assign w12345 = ~w12342 & ~w12344;
assign w12346 = ~w12343 & w12345;
assign w12347 = (w12346 & ~w3964) | (w12346 & w34568) | (~w3964 & w34568);
assign w12348 = a_8 & ~w12347;
assign w12349 = (~w3964 & w34569) | (~w3964 & w34570) | (w34569 & w34570);
assign w12350 = ~w12348 & ~w12349;
assign w12351 = w12341 & ~w12350;
assign w12352 = ~w12341 & w12350;
assign w12353 = ~w12351 & ~w12352;
assign w12354 = ~w12319 & w12328;
assign w12355 = ~w12329 & ~w12354;
assign w12356 = w12353 & ~w12355;
assign w12357 = (~w12351 & ~w12353) | (~w12351 & w34571) | (~w12353 & w34571);
assign w12358 = (w8298 & ~w3904) | (w8298 & w34572) | (~w3904 & w34572);
assign w12359 = (w8277 & ~w1308) | (w8277 & w34573) | (~w1308 & w34573);
assign w12360 = ~w3958 & w8295;
assign w12361 = ~w12359 & ~w12360;
assign w12362 = ~w12358 & w12361;
assign w12363 = (w12362 & ~w3943) | (w12362 & w34574) | (~w3943 & w34574);
assign w12364 = a_8 & w12363;
assign w12365 = (w3943 & w34575) | (w3943 & w34576) | (w34575 & w34576);
assign w12366 = ~w12364 & ~w12365;
assign w12367 = w12357 & ~w12366;
assign w12368 = ~w12357 & w12366;
assign w12369 = ~w12367 & ~w12368;
assign w12370 = w12340 & w12369;
assign w12371 = ~w12340 & ~w12369;
assign w12372 = ~w12370 & ~w12371;
assign w12373 = (~w3828 & w34579) | (~w3828 & w34580) | (w34579 & w34580);
assign w12374 = ~w12373 & w34581;
assign w12375 = (a_5 & w12373) | (a_5 & w34582) | (w12373 & w34582);
assign w12376 = ~w12374 & ~w12375;
assign w12377 = w12242 & ~w12291;
assign w12378 = ~w12290 & ~w12376;
assign w12379 = ~w12377 & w12378;
assign w12380 = ~w12376 & ~w12379;
assign w12381 = ~w12242 & ~w12290;
assign w12382 = ~w12291 & w12376;
assign w12383 = ~w12381 & w12382;
assign w12384 = ~w12379 & ~w12383;
assign w12385 = ~w12353 & w12355;
assign w12386 = ~w12356 & ~w12385;
assign w12387 = ~w12384 & ~w12386;
assign w12388 = ~w12380 & ~w12387;
assign w12389 = w12372 & ~w12388;
assign w12390 = ~w12372 & w12388;
assign w12391 = ~w12389 & ~w12390;
assign w12392 = ~w12213 & w12216;
assign w12393 = ~w11981 & ~w12099;
assign w12394 = ~w11984 & w12393;
assign w12395 = ~w12392 & ~w12394;
assign w12396 = w12300 & ~w12395;
assign w12397 = w12219 & ~w12298;
assign w12398 = (w12227 & w12230) | (w12227 & w34583) | (w12230 & w34583);
assign w12399 = (~w12398 & w12233) | (~w12398 & w34584) | (w12233 & w34584);
assign w12400 = w12384 & w12386;
assign w12401 = ~w12387 & ~w12400;
assign w12402 = w12399 & ~w12401;
assign w12403 = (~w12402 & ~w12219) | (~w12402 & w34585) | (~w12219 & w34585);
assign w12404 = ~w12396 & w12403;
assign w12405 = ~w12396 & w32445;
assign w12406 = ~w12399 & w12401;
assign w12407 = w12391 & w12406;
assign w12408 = ~w8285 & ~w8287;
assign w12409 = ~w8288 & ~w12408;
assign w12410 = (w8277 & ~w3904) | (w8277 & w34586) | (~w3904 & w34586);
assign w12411 = ~w3958 & w8298;
assign w12412 = ~w12410 & ~w12411;
assign w12413 = (w12412 & ~w4073) | (w12412 & w34587) | (~w4073 & w34587);
assign w12414 = a_8 & ~w12413;
assign w12415 = (~w4073 & w34588) | (~w4073 & w34589) | (w34588 & w34589);
assign w12416 = ~w12414 & ~w12415;
assign w12417 = ~w8255 & ~w8264;
assign w12418 = ~w8265 & ~w12417;
assign w12419 = ~w12416 & ~w12418;
assign w12420 = (~w12332 & ~w12333) | (~w12332 & w34590) | (~w12333 & w34590);
assign w12421 = w12416 & w12418;
assign w12422 = ~w12419 & ~w12421;
assign w12423 = w12420 & w12422;
assign w12424 = ~w12419 & ~w12423;
assign w12425 = ~w12409 & w12424;
assign w12426 = (~w12367 & ~w12369) | (~w12367 & w34591) | (~w12369 & w34591);
assign w12427 = ~w12420 & ~w12422;
assign w12428 = ~w12423 & ~w12427;
assign w12429 = ~w12426 & ~w12428;
assign w12430 = ~w12389 & w34592;
assign w12431 = ~w12407 & w12430;
assign w12432 = (w12431 & w12302) | (w12431 & w34593) | (w12302 & w34593);
assign w12433 = w12426 & w12428;
assign w12434 = ~w7880 & ~w8289;
assign w12435 = ~w8290 & ~w12434;
assign w12436 = w12409 & ~w12424;
assign w12437 = (~w12436 & ~w12433) | (~w12436 & w34594) | (~w12433 & w34594);
assign w12438 = w12435 & w12437;
assign w12439 = w12437 & w34595;
assign w12440 = ~w7502 & w7504;
assign w12441 = ~w7057 & ~w7207;
assign w12442 = ~w12440 & w12441;
assign w12443 = (~w7056 & w7508) | (~w7056 & w34597) | (w7508 & w34597);
assign w12444 = ~w7050 & ~w7053;
assign w12445 = ~w6454 & ~w6456;
assign w12446 = ~w6457 & ~w12445;
assign w12447 = ~w12444 & w12446;
assign w12448 = w12444 & ~w12446;
assign w12449 = w6458 & ~w6460;
assign w12450 = ~w6461 & ~w12449;
assign w12451 = ~w12448 & w12450;
assign w12452 = (~w12432 & w34602) | (~w12432 & w34603) | (w34602 & w34603);
assign w12453 = ~w6461 & ~w12452;
assign w12454 = ~w6071 & ~w6330;
assign w12455 = ~w1475 & w5286;
assign w12456 = (w5080 & ~w643) | (w5080 & w34605) | (~w643 & w34605);
assign w12457 = (w5016 & ~w1628) | (w5016 & w33133) | (~w1628 & w33133);
assign w12458 = ~w12456 & ~w12457;
assign w12459 = ~w12455 & w12458;
assign w12460 = (w12459 & ~w4041) | (w12459 & w34606) | (~w4041 & w34606);
assign w12461 = a_23 & ~w12460;
assign w12462 = (~w4041 & w34607) | (~w4041 & w34608) | (w34607 & w34608);
assign w12463 = ~w12461 & ~w12462;
assign w12464 = ~w5268 & ~w5276;
assign w12465 = ~w5277 & ~w12464;
assign w12466 = (~w6017 & ~w6019) | (~w6017 & w34609) | (~w6019 & w34609);
assign w12467 = w12465 & w12466;
assign w12468 = ~w12465 & ~w12466;
assign w12469 = ~w12467 & ~w12468;
assign w12470 = w12463 & w12469;
assign w12471 = ~w12463 & ~w12469;
assign w12472 = ~w12470 & ~w12471;
assign w12473 = (~w6033 & ~w6035) | (~w6033 & w34610) | (~w6035 & w34610);
assign w12474 = w12472 & w12473;
assign w12475 = ~w12472 & ~w12473;
assign w12476 = ~w12474 & ~w12475;
assign w12477 = ~w1397 & w5308;
assign w12478 = (w5816 & ~w3904) | (w5816 & w34611) | (~w3904 & w34611);
assign w12479 = (w5818 & ~w1308) | (w5818 & w34612) | (~w1308 & w34612);
assign w12480 = ~w12477 & ~w12479;
assign w12481 = ~w12478 & w12480;
assign w12482 = (w12481 & ~w3964) | (w12481 & w34613) | (~w3964 & w34613);
assign w12483 = a_20 & ~w12482;
assign w12484 = (~w3964 & w34614) | (~w3964 & w34615) | (w34614 & w34615);
assign w12485 = ~w12483 & ~w12484;
assign w12486 = w12476 & w12485;
assign w12487 = ~w12476 & ~w12485;
assign w12488 = ~w12486 & ~w12487;
assign w12489 = (~w6040 & ~w6042) | (~w6040 & w34616) | (~w6042 & w34616);
assign w12490 = (w3828 & w34617) | (w3828 & w34618) | (w34617 & w34618);
assign w12491 = (~w3958 & w12490) | (~w3958 & w34619) | (w12490 & w34619);
assign w12492 = ~a_17 & w12491;
assign w12493 = (~w12490 & w34620) | (~w12490 & w34621) | (w34620 & w34621);
assign w12494 = ~w12492 & ~w12493;
assign w12495 = ~w12489 & ~w12494;
assign w12496 = w12489 & w12494;
assign w12497 = ~w12495 & ~w12496;
assign w12498 = w12488 & w12497;
assign w12499 = ~w12488 & ~w12497;
assign w12500 = ~w12498 & ~w12499;
assign w12501 = (~w6046 & ~w6048) | (~w6046 & w34622) | (~w6048 & w34622);
assign w12502 = w12500 & w12501;
assign w12503 = (~w12502 & w6330) | (~w12502 & w34623) | (w6330 & w34623);
assign w12504 = ~w12500 & ~w12501;
assign w12505 = (~w12495 & ~w12497) | (~w12495 & w34626) | (~w12497 & w34626);
assign w12506 = (~w12467 & ~w12469) | (~w12467 & w34627) | (~w12469 & w34627);
assign w12507 = w5278 & ~w5280;
assign w12508 = ~w5281 & ~w12507;
assign w12509 = ~w1397 & w5286;
assign w12510 = ~w1475 & w5080;
assign w12511 = (w5016 & ~w643) | (w5016 & w34628) | (~w643 & w34628);
assign w12512 = ~w12509 & ~w12511;
assign w12513 = ~w12510 & w12512;
assign w12514 = (w12513 & ~w4056) | (w12513 & w34629) | (~w4056 & w34629);
assign w12515 = a_23 & ~w12514;
assign w12516 = (~w4056 & w34630) | (~w4056 & w34631) | (w34630 & w34631);
assign w12517 = ~w12515 & ~w12516;
assign w12518 = w12508 & w12517;
assign w12519 = ~w12508 & ~w12517;
assign w12520 = ~w12518 & ~w12519;
assign w12521 = ~w12506 & w12520;
assign w12522 = w12506 & ~w12520;
assign w12523 = ~w12521 & ~w12522;
assign w12524 = (~w12474 & ~w12476) | (~w12474 & w34632) | (~w12476 & w34632);
assign w12525 = (w5818 & ~w3904) | (w5818 & w34633) | (~w3904 & w34633);
assign w12526 = (w5308 & ~w1308) | (w5308 & w34634) | (~w1308 & w34634);
assign w12527 = ~w3958 & w5816;
assign w12528 = ~w12526 & ~w12527;
assign w12529 = ~w12525 & w12528;
assign w12530 = (w12529 & ~w3943) | (w12529 & w34635) | (~w3943 & w34635);
assign w12531 = a_20 & w12530;
assign w12532 = (w3943 & w34636) | (w3943 & w34637) | (w34636 & w34637);
assign w12533 = ~w12531 & ~w12532;
assign w12534 = ~w12524 & ~w12533;
assign w12535 = w12524 & w12533;
assign w12536 = ~w12534 & ~w12535;
assign w12537 = w12523 & w12536;
assign w12538 = ~w12523 & ~w12536;
assign w12539 = ~w12537 & ~w12538;
assign w12540 = ~w12505 & w12539;
assign w12541 = w12505 & ~w12539;
assign w12542 = ~w12540 & ~w12541;
assign w12543 = ~w12504 & w12542;
assign w12544 = (~w12534 & ~w12536) | (~w12534 & w34638) | (~w12536 & w34638);
assign w12545 = w5293 & ~w5295;
assign w12546 = ~w5296 & ~w12545;
assign w12547 = (~w12518 & ~w12520) | (~w12518 & w34639) | (~w12520 & w34639);
assign w12548 = ~w12546 & ~w12547;
assign w12549 = w12546 & w12547;
assign w12550 = ~w12548 & ~w12549;
assign w12551 = (w5308 & ~w3904) | (w5308 & w34640) | (~w3904 & w34640);
assign w12552 = ~w3958 & w5818;
assign w12553 = ~w12551 & ~w12552;
assign w12554 = (w12553 & ~w4073) | (w12553 & w34641) | (~w4073 & w34641);
assign w12555 = a_20 & w12554;
assign w12556 = (w4073 & w34642) | (w4073 & w34643) | (w34642 & w34643);
assign w12557 = ~w12555 & ~w12556;
assign w12558 = w12550 & ~w12557;
assign w12559 = ~w12550 & w12557;
assign w12560 = ~w12558 & ~w12559;
assign w12561 = w12544 & ~w12560;
assign w12562 = w5336 & ~w5354;
assign w12563 = ~w5355 & ~w12562;
assign w12564 = (~w12548 & ~w12550) | (~w12548 & w34644) | (~w12550 & w34644);
assign w12565 = ~w5316 & ~w5334;
assign w12566 = ~w5335 & ~w12565;
assign w12567 = w12564 & ~w12566;
assign w12568 = ~w12561 & ~w12567;
assign w12569 = w12563 & w12568;
assign w12570 = w12543 & w12569;
assign w12571 = ~w12564 & w12566;
assign w12572 = w12563 & w12571;
assign w12573 = ~w12544 & w12560;
assign w12574 = ~w12540 & ~w12573;
assign w12575 = w12569 & ~w12574;
assign w12576 = ~w12572 & ~w12575;
assign w12577 = (~w12452 & w34647) | (~w12452 & w34648) | (w34647 & w34648);
assign w12578 = (~w5350 & ~w5351) | (~w5350 & w34649) | (~w5351 & w34649);
assign w12579 = ~w5078 & w5086;
assign w12580 = ~w5087 & ~w12579;
assign w12581 = ~w12578 & w12580;
assign w12582 = w12578 & ~w12580;
assign w12583 = w5088 & ~w5090;
assign w12584 = (~w12583 & ~w12578) | (~w12583 & w34651) | (~w12578 & w34651);
assign w12585 = w5033 & w12584;
assign w12586 = ~w5031 & ~w5092;
assign w12587 = (~w12577 & w34655) | (~w12577 & w34656) | (w34655 & w34656);
assign w12588 = (~w4649 & w12587) | (~w4649 & w34658) | (w12587 & w34658);
assign w12589 = w4501 & w12588;
assign w12590 = w4474 & ~w4476;
assign w12591 = ~w4477 & ~w12590;
assign w12592 = (w12588 & w34660) | (w12588 & w34661) | (w34660 & w34661);
assign w12593 = w4080 & w4082;
assign w12594 = ~w4083 & ~w12593;
assign w12595 = (w12588 & w34664) | (w12588 & w34665) | (w34664 & w34665);
assign w12596 = (w12588 & w34668) | (w12588 & w34669) | (w34668 & w34669);
assign w12597 = (~w12588 & w34670) | (~w12588 & w34671) | (w34670 & w34671);
assign w12598 = ~w12596 & ~w12597;
assign w12599 = w668 & w12598;
assign w12600 = (~w12588 & w34672) | (~w12588 & w34673) | (w34672 & w34673);
assign w12601 = ~w12595 & ~w12600;
assign w12602 = w1327 & w12601;
assign w12603 = (~w12588 & w34674) | (~w12588 & w34675) | (w34674 & w34675);
assign w12604 = ~w12592 & ~w12603;
assign w12605 = w1399 & w12604;
assign w12606 = (~w12587 & w34676) | (~w12587 & w34677) | (w34676 & w34677);
assign w12607 = ~w12589 & ~w12606;
assign w12608 = ~w12604 & ~w12607;
assign w12609 = ~w4697 & ~w5031;
assign w12610 = (w12577 & w34678) | (w12577 & w34679) | (w34678 & w34679);
assign w12611 = (w12577 & w34680) | (w12577 & w34681) | (w34680 & w34681);
assign w12612 = ~w4697 & ~w12611;
assign w12613 = ~w12610 & ~w12612;
assign w12614 = (w4650 & w12587) | (w4650 & w34682) | (w12587 & w34682);
assign w12615 = ~w12587 & w34683;
assign w12616 = ~w12588 & ~w12615;
assign w12617 = ~w12614 & ~w12616;
assign w12618 = ~w12613 & ~w12617;
assign w12619 = ~w12447 & ~w12448;
assign w12620 = (w12432 & w34684) | (w12432 & w34685) | (w34684 & w34685);
assign w12621 = (~w12432 & w34686) | (~w12432 & w34687) | (w34686 & w34687);
assign w12622 = ~w12620 & ~w12621;
assign w12623 = ~w7505 & ~w12440;
assign w12624 = (w31761 & w12432) | (w31761 & w34688) | (w12432 & w34688);
assign w12625 = (w12432 & w34689) | (w12432 & w34690) | (w34689 & w34690);
assign w12626 = (~w7058 & w7508) | (~w7058 & w34691) | (w7508 & w34691);
assign w12627 = ~w7509 & ~w12626;
assign w12628 = (~w12432 & w34692) | (~w12432 & w34693) | (w34692 & w34693);
assign w12629 = (w12432 & w34694) | (w12432 & w34695) | (w34694 & w34695);
assign w12630 = ~w12628 & ~w12629;
assign w12631 = ~w12622 & w12630;
assign w12632 = (~w12302 & w34696) | (~w12302 & w34697) | (w34696 & w34697);
assign w12633 = w8290 & ~w8292;
assign w12634 = ~w8293 & ~w12633;
assign w12635 = w12632 & w12634;
assign w12636 = ~w12632 & ~w12634;
assign w12637 = ~w12635 & ~w12636;
assign w12638 = ~w12429 & ~w12433;
assign w12639 = ~w12389 & w12638;
assign w12640 = ~w12407 & w12639;
assign w12641 = ~w12425 & ~w12436;
assign w12642 = ~w12433 & w12641;
assign w12643 = (~w12302 & w34698) | (~w12302 & w34699) | (w34698 & w34699);
assign w12644 = ~w12425 & ~w12435;
assign w12645 = (w12302 & w34700) | (w12302 & w34701) | (w34700 & w34701);
assign w12646 = ~w12632 & ~w12645;
assign w12647 = w12637 & ~w12646;
assign w12648 = ~w12634 & w12646;
assign w12649 = ~w12647 & ~w12648;
assign w12650 = (w12302 & w34702) | (w12302 & w34703) | (w34702 & w34703);
assign w12651 = ~w12643 & ~w12650;
assign w12652 = w12646 & w12651;
assign w12653 = w12425 & w12435;
assign w12654 = ~w12644 & ~w12653;
assign w12655 = ~w12650 & ~w12654;
assign w12656 = w12650 & w12654;
assign w12657 = ~w12655 & ~w12656;
assign w12658 = ~w12652 & w12657;
assign w12659 = w12649 & ~w12658;
assign w12660 = (~w12432 & w34704) | (~w12432 & w34705) | (w34704 & w34705);
assign w12661 = ~w12624 & ~w12660;
assign w12662 = ~w12637 & ~w12661;
assign w12663 = ~w12648 & ~w12662;
assign w12664 = ~w12659 & w12663;
assign w12665 = w7505 & ~w7507;
assign w12666 = ~w7508 & ~w12665;
assign w12667 = (~w12432 & w34706) | (~w12432 & w34707) | (w34706 & w34707);
assign w12668 = ~w12625 & ~w12667;
assign w12669 = w12627 & w12668;
assign w12670 = w12637 & w12661;
assign w12671 = (~w12432 & w34708) | (~w12432 & w34709) | (w34708 & w34709);
assign w12672 = (w12432 & w34710) | (w12432 & w34711) | (w34710 & w34711);
assign w12673 = ~w12671 & ~w12672;
assign w12674 = ~w11501 & ~w11502;
assign w12675 = w11676 & w11683;
assign w12676 = w10849 & w11338;
assign w12677 = w11332 & ~w12676;
assign w12678 = ~w11332 & w12676;
assign w12679 = ~w12677 & ~w12678;
assign w12680 = w12675 & ~w12679;
assign w12681 = ~w12674 & w12680;
assign w12682 = ~w11338 & ~w11499;
assign w12683 = w11333 & ~w11499;
assign w12684 = ~w12682 & ~w12683;
assign w12685 = ~w11501 & w12684;
assign w12686 = ~w11502 & ~w12675;
assign w12687 = ~w12679 & w12686;
assign w12688 = w12685 & ~w12687;
assign w12689 = ~w12681 & w12688;
assign w12690 = ~w12674 & w12675;
assign w12691 = ~w12674 & w31766;
assign w12692 = w11676 & w11825;
assign w12693 = ~w11676 & ~w11825;
assign w12694 = ~w12692 & ~w12693;
assign w12695 = w12674 & ~w12675;
assign w12696 = ~w12694 & w12695;
assign w12697 = ~w12691 & ~w12696;
assign w12698 = w12689 & w12697;
assign w12699 = ~w11678 & w11683;
assign w12700 = (w11825 & w11678) | (w11825 & w31767) | (w11678 & w31767);
assign w12701 = ~w11827 & ~w12700;
assign w12702 = ~w12690 & ~w12695;
assign w12703 = w12701 & w12702;
assign w12704 = ~w12698 & ~w12703;
assign w12705 = ~w11960 & ~w11974;
assign w12706 = w11830 & ~w12705;
assign w12707 = ~w11830 & w12705;
assign w12708 = ~w12706 & ~w12707;
assign w12709 = ~w11968 & w12708;
assign w12710 = w11968 & ~w12708;
assign w12711 = ~w12709 & ~w12710;
assign w12712 = w12700 & w12711;
assign w12713 = ~w12700 & ~w12711;
assign w12714 = ~w12712 & ~w12713;
assign w12715 = w12704 & ~w12714;
assign w12716 = ~w12701 & w12714;
assign w12717 = ~w12715 & ~w12716;
assign w12718 = ~w12100 & ~w12394;
assign w12719 = ~w11827 & ~w11968;
assign w12720 = ~w11961 & ~w11964;
assign w12721 = (~w12720 & w11827) | (~w12720 & w31768) | (w11827 & w31768);
assign w12722 = ~w11827 & w31769;
assign w12723 = ~w12721 & ~w12722;
assign w12724 = ~w12718 & ~w12723;
assign w12725 = ~w12708 & w12718;
assign w12726 = ~w11971 & w12718;
assign w12727 = (~w12725 & ~w12726) | (~w12725 & w31770) | (~w12726 & w31770);
assign w12728 = ~w12724 & w12727;
assign w12729 = w12717 & w12728;
assign w12730 = (~w12718 & w11971) | (~w12718 & w31771) | (w11971 & w31771);
assign w12731 = ~w11971 & w31772;
assign w12732 = ~w12730 & ~w12731;
assign w12733 = ~w12217 & ~w12392;
assign w12734 = w12100 & ~w12733;
assign w12735 = ~w12100 & w12733;
assign w12736 = ~w12734 & ~w12735;
assign w12737 = w12708 & w12719;
assign w12738 = ~w12708 & ~w12719;
assign w12739 = ~w12737 & ~w12738;
assign w12740 = w12736 & ~w12739;
assign w12741 = w12732 & ~w12740;
assign w12742 = (~w12741 & ~w12717) | (~w12741 & w31773) | (~w12717 & w31773);
assign w12743 = w12730 & w12736;
assign w12744 = w12718 & w12733;
assign w12745 = w11977 & w12744;
assign w12746 = ~w12743 & ~w12745;
assign w12747 = ~w11976 & ~w12394;
assign w12748 = ~w11971 & w12747;
assign w12749 = (~w12100 & w11971) | (~w12100 & w31774) | (w11971 & w31774);
assign w12750 = ~w12299 & ~w12397;
assign w12751 = ~w12392 & ~w12750;
assign w12752 = w12392 & w12750;
assign w12753 = ~w12751 & ~w12752;
assign w12754 = w12749 & ~w12753;
assign w12755 = w12217 & ~w12750;
assign w12756 = ~w12217 & w12750;
assign w12757 = ~w12755 & ~w12756;
assign w12758 = ~w12749 & w12757;
assign w12759 = ~w12754 & ~w12758;
assign w12760 = w12746 & ~w12759;
assign w12761 = ~w12742 & w12760;
assign w12762 = ~w12100 & ~w12217;
assign w12763 = ~w12750 & w12762;
assign w12764 = ~w11977 & w12763;
assign w12765 = ~w11977 & w12744;
assign w12766 = ~w12217 & ~w12395;
assign w12767 = ~w12750 & w12766;
assign w12768 = w12750 & ~w12766;
assign w12769 = ~w12767 & ~w12768;
assign w12770 = ~w12765 & ~w12769;
assign w12771 = ~w12764 & ~w12770;
assign w12772 = w12735 & ~w12748;
assign w12773 = ~w12733 & ~w12749;
assign w12774 = ~w12772 & ~w12773;
assign w12775 = w12771 & ~w12774;
assign w12776 = ~w12402 & ~w12406;
assign w12777 = w12299 & ~w12776;
assign w12778 = ~w12299 & w12776;
assign w12779 = ~w12777 & ~w12778;
assign w12780 = ~w12770 & w31775;
assign w12781 = ~w12775 & ~w12780;
assign w12782 = (~w12776 & w12396) | (~w12776 & w31776) | (w12396 & w31776);
assign w12783 = w12300 & w32450;
assign w12784 = ~w11977 & w12783;
assign w12785 = ~w12396 & w12776;
assign w12786 = ~w12396 & w31777;
assign w12787 = ~w12302 & w12786;
assign w12788 = ~w12782 & ~w12784;
assign w12789 = ~w12787 & w12788;
assign w12790 = ~w12391 & ~w12406;
assign w12791 = (w12790 & w12302) | (w12790 & w31778) | (w12302 & w31778);
assign w12792 = (~w12407 & w12302) | (~w12407 & w32451) | (w12302 & w32451);
assign w12793 = ~w12791 & w12792;
assign w12794 = w12789 & w12793;
assign w12795 = w12389 & ~w12638;
assign w12796 = ~w12639 & ~w12795;
assign w12797 = w12792 & w31779;
assign w12798 = ~w12794 & ~w12797;
assign w12799 = w12781 & w12798;
assign w12800 = ~w12761 & w12799;
assign w12801 = (w12762 & w11971) | (w12762 & w31780) | (w11971 & w31780);
assign w12802 = (w12299 & w12395) | (w12299 & w34712) | (w12395 & w34712);
assign w12803 = ~w12801 & w12802;
assign w12804 = ~w12302 & w12785;
assign w12805 = ~w12803 & w12804;
assign w12806 = ~w12766 & w12777;
assign w12807 = w12750 & w12776;
assign w12808 = ~w12806 & ~w12807;
assign w12809 = w12762 & ~w12807;
assign w12810 = ~w11977 & w12809;
assign w12811 = ~w12808 & ~w12810;
assign w12812 = ~w12750 & ~w12776;
assign w12813 = w12396 & w12812;
assign w12814 = w12301 & w12812;
assign w12815 = ~w11977 & w12814;
assign w12816 = ~w12813 & ~w12815;
assign w12817 = ~w12811 & w12816;
assign w12818 = ~w12805 & w12817;
assign w12819 = ~w12780 & ~w12818;
assign w12820 = ~w12789 & ~w12793;
assign w12821 = ~w12819 & ~w12820;
assign w12822 = w12798 & ~w12821;
assign w12823 = ~w12390 & w12638;
assign w12824 = w12390 & ~w12638;
assign w12825 = ~w12823 & ~w12824;
assign w12826 = ~w12793 & ~w12825;
assign w12827 = (~w12826 & w12821) | (~w12826 & w32452) | (w12821 & w32452);
assign w12828 = ~w12800 & w12827;
assign w12829 = (w12825 & ~w12792) | (w12825 & w31781) | (~w12792 & w31781);
assign w12830 = ~w12797 & ~w12829;
assign w12831 = w12651 & ~w12830;
assign w12832 = ~w12651 & w12830;
assign w12833 = ~w12831 & ~w12832;
assign w12834 = w12828 & w12833;
assign w12835 = (~w12652 & w12830) | (~w12652 & w34713) | (w12830 & w34713);
assign w12836 = ~w12831 & w32453;
assign w12837 = ~w12831 & w34714;
assign w12838 = (w12837 & ~w12828) | (w12837 & w34715) | (~w12828 & w34715);
assign w12839 = ~w12670 & w12673;
assign w12840 = ~w12669 & w12839;
assign w12841 = ~w12664 & w12840;
assign w12842 = ~w12838 & w12841;
assign w12843 = w12622 & ~w12630;
assign w12844 = ~w12661 & ~w12668;
assign w12845 = ~w12630 & ~w12668;
assign w12846 = ~w12844 & ~w12845;
assign w12847 = ~w12843 & w12846;
assign w12848 = ~w12447 & ~w12450;
assign w12849 = w12447 & w12450;
assign w12850 = ~w12848 & ~w12849;
assign w12851 = (w12432 & w34716) | (w12432 & w34717) | (w34716 & w34717);
assign w12852 = (~w12432 & w34718) | (~w12432 & w34719) | (w34718 & w34719);
assign w12853 = ~w12851 & ~w12852;
assign w12854 = (w12842 & w34720) | (w12842 & w34721) | (w34720 & w34721);
assign w12855 = (w12432 & w34722) | (w12432 & w34723) | (w34722 & w34723);
assign w12856 = ~w12452 & ~w12855;
assign w12857 = (~w12452 & w34724) | (~w12452 & w34725) | (w34724 & w34725);
assign w12858 = w6331 & w12453;
assign w12859 = (w12454 & w12452) | (w12454 & w34726) | (w12452 & w34726);
assign w12860 = (~w12859 & w12858) | (~w12859 & w34727) | (w12858 & w34727);
assign w12861 = ~w12856 & w12860;
assign w12862 = (w12842 & w34728) | (w12842 & w34729) | (w34728 & w34729);
assign w12863 = w12622 & w12856;
assign w12864 = w12856 & ~w12860;
assign w12865 = (~w12863 & w12860) | (~w12863 & w34730) | (w12860 & w34730);
assign w12866 = ~w12502 & ~w12504;
assign w12867 = (w12452 & w34731) | (w12452 & w34732) | (w34731 & w34732);
assign w12868 = (~w12452 & w34733) | (~w12452 & w34734) | (w34733 & w34734);
assign w12869 = ~w12867 & ~w12868;
assign w12870 = ~w12860 & w12869;
assign w12871 = (w12452 & w34736) | (w12452 & w34737) | (w34736 & w34737);
assign w12872 = ~w12502 & ~w12542;
assign w12873 = (~w12452 & w34738) | (~w12452 & w34739) | (w34738 & w34739);
assign w12874 = ~w12871 & ~w12873;
assign w12875 = ~w12561 & ~w12573;
assign w12876 = (~w12452 & w34742) | (~w12452 & w34743) | (w34742 & w34743);
assign w12877 = (w12452 & w34744) | (w12452 & w34745) | (w34744 & w34745);
assign w12878 = ~w12876 & ~w12877;
assign w12879 = ~w12874 & w12878;
assign w12880 = w12502 & w12542;
assign w12881 = ~w12872 & ~w12880;
assign w12882 = (~w12452 & w34746) | (~w12452 & w34747) | (w34746 & w34747);
assign w12883 = (w12452 & w34748) | (w12452 & w34749) | (w34748 & w34749);
assign w12884 = ~w12882 & ~w12883;
assign w12885 = (~w12884 & ~w12860) | (~w12884 & w34750) | (~w12860 & w34750);
assign w12886 = ~w12879 & w12885;
assign w12887 = w12874 & ~w12878;
assign w12888 = w12869 & w12874;
assign w12889 = ~w12887 & ~w12888;
assign w12890 = ~w12567 & ~w12571;
assign w12891 = (w12452 & w34754) | (w12452 & w34755) | (w34754 & w34755);
assign w12892 = w12890 & w12891;
assign w12893 = (~w12452 & w34756) | (~w12452 & w34757) | (w34756 & w34757);
assign w12894 = ~w12892 & ~w12893;
assign w12895 = ~w12878 & w12894;
assign w12896 = w12889 & ~w12895;
assign w12897 = w12878 & ~w12894;
assign w12898 = ~w12563 & ~w12571;
assign w12899 = ~w12572 & ~w12898;
assign w12900 = (~w12452 & w34760) | (~w12452 & w34761) | (w34760 & w34761);
assign w12901 = (w12452 & w34762) | (w12452 & w34763) | (w34762 & w34763);
assign w12902 = ~w12900 & ~w12901;
assign w12903 = (~w12902 & w12894) | (~w12902 & w34764) | (w12894 & w34764);
assign w12904 = (w12862 & w34765) | (w12862 & w34766) | (w34765 & w34766);
assign w12905 = (w12898 & ~w12891) | (w12898 & w34767) | (~w12891 & w34767);
assign w12906 = w12577 & ~w12905;
assign w12907 = ~w12581 & ~w12582;
assign w12908 = (~w12907 & ~w12577) | (~w12907 & w34768) | (~w12577 & w34768);
assign w12909 = w12577 & w34769;
assign w12910 = ~w12908 & ~w12909;
assign w12911 = ~w12906 & w12910;
assign w12912 = ~w5091 & ~w12583;
assign w12913 = (~w12582 & ~w12577) | (~w12582 & w34770) | (~w12577 & w34770);
assign w12914 = w12912 & w12913;
assign w12915 = (w12577 & w34771) | (w12577 & w34772) | (w34771 & w34772);
assign w12916 = ~w12914 & ~w12915;
assign w12917 = ~w12910 & w12916;
assign w12918 = w12906 & ~w12910;
assign w12919 = w12894 & w12906;
assign w12920 = ~w12918 & ~w12919;
assign w12921 = ~w12917 & w12920;
assign w12922 = w12910 & ~w12916;
assign w12923 = ~w5033 & ~w5091;
assign w12924 = ~w5092 & ~w12923;
assign w12925 = (w12577 & w34774) | (w12577 & w34775) | (w34774 & w34775);
assign w12926 = (~w12577 & w34776) | (~w12577 & w34777) | (w34776 & w34777);
assign w12927 = ~w12925 & ~w12926;
assign w12928 = (~w12927 & w12916) | (~w12927 & w34778) | (w12916 & w34778);
assign w12929 = (w12904 & w34779) | (w12904 & w34780) | (w34779 & w34780);
assign w12930 = (w12923 & ~w12913) | (w12923 & w34781) | (~w12913 & w34781);
assign w12931 = w12611 & ~w12930;
assign w12932 = w12613 & ~w12931;
assign w12933 = (w12904 & w34782) | (w12904 & w34783) | (w34782 & w34783);
assign w12934 = w12916 & w12931;
assign w12935 = ~w12930 & w34784;
assign w12936 = ~w12934 & ~w12935;
assign w12937 = w12613 & w12617;
assign w12938 = ~w12618 & ~w12937;
assign w12939 = (w12938 & w12933) | (w12938 & w34785) | (w12933 & w34785);
assign w12940 = ~w12614 & ~w12615;
assign w12941 = w4501 & ~w12940;
assign w12942 = ~w4501 & w12940;
assign w12943 = ~w12941 & ~w12942;
assign w12944 = (w12933 & w34788) | (w12933 & w34789) | (w34788 & w34789);
assign w12945 = w12607 & ~w12617;
assign w12946 = w12604 & w12607;
assign w12947 = ~w12945 & ~w12946;
assign w12948 = ~w12601 & ~w12604;
assign w12949 = w12601 & w12604;
assign w12950 = ~w12948 & ~w12949;
assign w12951 = (~w12944 & w34791) | (~w12944 & w34792) | (w34791 & w34792);
assign w12952 = (w12588 & w34793) | (w12588 & w34794) | (w34793 & w34794);
assign w12953 = (~w12588 & w34795) | (~w12588 & w34796) | (w34795 & w34796);
assign w12954 = ~w12952 & ~w12953;
assign w12955 = w3976 & w12954;
assign w12956 = ~w3976 & ~w12954;
assign w12957 = ~w12955 & ~w12956;
assign w12958 = ~w12948 & w12957;
assign w12959 = (w12944 & w34797) | (w12944 & w34798) | (w34797 & w34798);
assign w12960 = (~w12944 & w34801) | (~w12944 & w34802) | (w34801 & w34802);
assign w12961 = ~w12959 & ~w12960;
assign w12962 = ~w12602 & ~w12605;
assign w12963 = ~w12599 & w12962;
assign w12964 = (w12963 & ~w12961) | (w12963 & w34803) | (~w12961 & w34803);
assign w12965 = w666 & ~w12964;
assign w12966 = (~w664 & w12964) | (~w664 & w34804) | (w12964 & w34804);
assign w12967 = ~w252 & ~w265;
assign w12968 = w340 & w3014;
assign w12969 = ~w290 & w1377;
assign w12970 = w1814 & w2159;
assign w12971 = w12967 & w12970;
assign w12972 = w2217 & w12969;
assign w12973 = w12968 & w12972;
assign w12974 = w1359 & w12971;
assign w12975 = w12973 & w12974;
assign w12976 = w1315 & w12975;
assign w12977 = w1451 & w34805;
assign w12978 = w663 & ~w12977;
assign w12979 = w527 & ~w663;
assign w12980 = w12977 & w12979;
assign w12981 = ~w12978 & ~w12980;
assign w12982 = (~w3865 & ~w3866) | (~w3865 & w34806) | (~w3866 & w34806);
assign w12983 = ~w130 & w3883;
assign w12984 = ~w89 & w2454;
assign w12985 = w1237 & w12984;
assign w12986 = w1335 & w2979;
assign w12987 = w12985 & w12986;
assign w12988 = w3923 & w12987;
assign w12989 = w5521 & w12988;
assign w12990 = w1599 & w12983;
assign w12991 = w12989 & w12990;
assign w12992 = w528 & w12991;
assign w12993 = w1306 & w12992;
assign w12994 = ~w3862 & w34807;
assign w12995 = (w12993 & w3862) | (w12993 & w34808) | (w3862 & w34808);
assign w12996 = ~w12994 & ~w12995;
assign w12997 = w1327 & ~w3958;
assign w12998 = (~w12997 & ~w4073) | (~w12997 & w34809) | (~w4073 & w34809);
assign w12999 = w12996 & ~w12998;
assign w13000 = (~w4073 & w34810) | (~w4073 & w34811) | (w34810 & w34811);
assign w13001 = ~w12999 & ~w13000;
assign w13002 = ~w12982 & w13001;
assign w13003 = w12982 & ~w13001;
assign w13004 = ~w13002 & ~w13003;
assign w13005 = w3974 & ~w13004;
assign w13006 = ~w3974 & w13004;
assign w13007 = ~w13005 & ~w13006;
assign w13008 = (~w12588 & w34812) | (~w12588 & w34813) | (w34812 & w34813);
assign w13009 = (w12588 & w34814) | (w12588 & w34815) | (w34814 & w34815);
assign w13010 = ~w13008 & ~w13009;
assign w13011 = ~w12598 & ~w13010;
assign w13012 = (~w12588 & w34816) | (~w12588 & w34817) | (w34816 & w34817);
assign w13013 = ~w13011 & ~w13012;
assign w13014 = ~w13011 & w34818;
assign w13015 = w1327 & w12598;
assign w13016 = w1399 & w12601;
assign w13017 = w12598 & w12601;
assign w13018 = (~w12944 & w34819) | (~w12944 & w34820) | (w34819 & w34820);
assign w13019 = w13010 & w13018;
assign w13020 = ~w13010 & ~w13018;
assign w13021 = ~w13019 & ~w13020;
assign w13022 = ~w13015 & ~w13016;
assign w13023 = ~w13014 & w13022;
assign w13024 = (w13023 & w13021) | (w13023 & w34821) | (w13021 & w34821);
assign w13025 = w12981 & ~w13024;
assign w13026 = (w13021 & w34822) | (w13021 & w34823) | (w34822 & w34823);
assign w13027 = ~w13025 & w34824;
assign w13028 = (w12966 & w13025) | (w12966 & w34825) | (w13025 & w34825);
assign w13029 = ~w13027 & ~w13028;
assign w13030 = ~w404 & w3627;
assign w13031 = ~w167 & ~w368;
assign w13032 = ~w789 & w13031;
assign w13033 = ~w451 & ~w583;
assign w13034 = ~w730 & w13033;
assign w13035 = w871 & w13034;
assign w13036 = ~w112 & ~w206;
assign w13037 = ~w428 & w13036;
assign w13038 = w1041 & w1273;
assign w13039 = w2370 & w2839;
assign w13040 = w2966 & w3344;
assign w13041 = w13039 & w13040;
assign w13042 = w13037 & w13038;
assign w13043 = w13030 & w13032;
assign w13044 = w13042 & w13043;
assign w13045 = w2568 & w13041;
assign w13046 = w13035 & w13045;
assign w13047 = w13044 & w13046;
assign w13048 = w2273 & w34826;
assign w13049 = w308 & ~w13048;
assign w13050 = ~w429 & ~w543;
assign w13051 = ~w157 & ~w169;
assign w13052 = ~w459 & ~w710;
assign w13053 = w13051 & w13052;
assign w13054 = w1604 & w13050;
assign w13055 = w13053 & w13054;
assign w13056 = w695 & w1009;
assign w13057 = w2192 & w3160;
assign w13058 = w13056 & w13057;
assign w13059 = ~w213 & w995;
assign w13060 = ~w170 & ~w352;
assign w13061 = w1641 & w4085;
assign w13062 = ~w152 & ~w220;
assign w13063 = ~w446 & w13062;
assign w13064 = w13060 & w13063;
assign w13065 = w4864 & w13059;
assign w13066 = w13061 & w13065;
assign w13067 = w13064 & w13066;
assign w13068 = ~w147 & ~w363;
assign w13069 = ~w428 & w13068;
assign w13070 = w2438 & w2681;
assign w13071 = w3119 & w4713;
assign w13072 = w13070 & w13071;
assign w13073 = w2015 & w13069;
assign w13074 = w4851 & w13073;
assign w13075 = w13055 & w13072;
assign w13076 = w13058 & w13075;
assign w13077 = w13074 & w13076;
assign w13078 = w102 & w277;
assign w13079 = w13067 & w13078;
assign w13080 = w13077 & w13079;
assign w13081 = w2642 & w13080;
assign w13082 = ~w242 & ~w1123;
assign w13083 = w911 & w1640;
assign w13084 = ~w197 & w1691;
assign w13085 = w2151 & w2398;
assign w13086 = w3305 & w5390;
assign w13087 = w13082 & w13086;
assign w13088 = w13084 & w13085;
assign w13089 = w13083 & w13088;
assign w13090 = w1508 & w13087;
assign w13091 = w2618 & w13090;
assign w13092 = w3566 & w13089;
assign w13093 = w13091 & w13092;
assign w13094 = ~w309 & ~w580;
assign w13095 = w731 & w1988;
assign w13096 = w2337 & w3489;
assign w13097 = w3674 & w4111;
assign w13098 = w4911 & w5169;
assign w13099 = w13094 & w13098;
assign w13100 = w13096 & w13097;
assign w13101 = w4344 & w13095;
assign w13102 = w13100 & w13101;
assign w13103 = w13099 & w13102;
assign w13104 = w2158 & w13103;
assign w13105 = w2566 & w13104;
assign w13106 = w13093 & w13105;
assign w13107 = w3357 & w13106;
assign w13108 = ~w13081 & ~w13107;
assign w13109 = a_20 & ~w5304;
assign w13110 = ~a_19 & w5298;
assign w13111 = (~w13110 & w5304) | (~w13110 & w34827) | (w5304 & w34827);
assign w13112 = w13081 & w13107;
assign w13113 = ~w13108 & ~w13112;
assign w13114 = ~w13111 & w13113;
assign w13115 = (~w13108 & ~w13113) | (~w13108 & w34828) | (~w13113 & w34828);
assign w13116 = w13048 & ~w13115;
assign w13117 = ~w13048 & w13115;
assign w13118 = ~w13116 & ~w13117;
assign w13119 = (w1327 & w12616) | (w1327 & w34829) | (w12616 & w34829);
assign w13120 = (w1399 & w12612) | (w1399 & w34830) | (w12612 & w34830);
assign w13121 = ~w12589 & w34831;
assign w13122 = (~w12933 & w34832) | (~w12933 & w34833) | (w34832 & w34833);
assign w13123 = ~w12944 & ~w13122;
assign w13124 = ~w13119 & ~w13120;
assign w13125 = ~w13121 & w13124;
assign w13126 = (w13125 & ~w13123) | (w13125 & w34834) | (~w13123 & w34834);
assign w13127 = w13118 & ~w13126;
assign w13128 = ~w308 & w13048;
assign w13129 = ~w13049 & ~w13128;
assign w13130 = (~w13126 & w34836) | (~w13126 & w34837) | (w34836 & w34837);
assign w13131 = w511 & ~w513;
assign w13132 = ~w514 & ~w13131;
assign w13133 = (~w13126 & w34840) | (~w13126 & w34841) | (w34840 & w34841);
assign w13134 = (w13126 & w34842) | (w13126 & w34843) | (w34842 & w34843);
assign w13135 = ~w13133 & ~w13134;
assign w13136 = w668 & w12601;
assign w13137 = w1327 & w12604;
assign w13138 = ~w12589 & w34844;
assign w13139 = (w12944 & w34845) | (w12944 & w34846) | (w34845 & w34846);
assign w13140 = ~w12951 & ~w13139;
assign w13141 = ~w13137 & ~w13138;
assign w13142 = ~w13136 & w13141;
assign w13143 = (w13142 & w13140) | (w13142 & w34847) | (w13140 & w34847);
assign w13144 = w13135 & ~w13143;
assign w13145 = (~w13133 & ~w13135) | (~w13133 & w34848) | (~w13135 & w34848);
assign w13146 = (~w12961 & w34849) | (~w12961 & w34850) | (w34849 & w34850);
assign w13147 = ~w12965 & ~w13146;
assign w13148 = ~w13145 & w13147;
assign w13149 = w13145 & ~w13147;
assign w13150 = ~w13148 & ~w13149;
assign w13151 = ~w1965 & w12967;
assign w13152 = w3924 & w13151;
assign w13153 = w1328 & w13152;
assign w13154 = w3914 & w13153;
assign w13155 = w3845 & w13154;
assign w13156 = w3887 & w13155;
assign w13157 = w12993 & ~w13156;
assign w13158 = w574 & w1694;
assign w13159 = w1335 & w13158;
assign w13160 = w3869 & w13159;
assign w13161 = w1590 & w13160;
assign w13162 = w3900 & w13161;
assign w13163 = w1308 & w13162;
assign w13164 = ~w12993 & w13163;
assign w13165 = w12993 & ~w13163;
assign w13166 = ~w13164 & ~w13165;
assign w13167 = ~w13157 & w13166;
assign w13168 = ~w12993 & w13156;
assign w13169 = ~w13157 & ~w13168;
assign w13170 = (~w12998 & w34852) | (~w12998 & w34853) | (w34852 & w34853);
assign w13171 = (w12998 & w34854) | (w12998 & w34855) | (w34854 & w34855);
assign w13172 = ~w13170 & ~w13171;
assign w13173 = (w12588 & w34860) | (w12588 & w34861) | (w34860 & w34861);
assign w13174 = w13172 & w13173;
assign w13175 = (w13173 & w34863) | (w13173 & w34864) | (w34863 & w34864);
assign w13176 = (~w13173 & w13188) | (~w13173 & w34865) | (w13188 & w34865);
assign w13177 = ~w13175 & ~w13176;
assign w13178 = w4446 & w13177;
assign w13179 = (~w12588 & w34866) | (~w12588 & w34867) | (w34866 & w34867);
assign w13180 = ~w13174 & ~w13179;
assign w13181 = ~w13174 & w34868;
assign w13182 = ~w13011 & w34869;
assign w13183 = (~w12998 & w34870) | (~w12998 & w34871) | (w34870 & w34871);
assign w13184 = (w12998 & w34872) | (w12998 & w34873) | (w34872 & w34873);
assign w13185 = ~w13183 & ~w13184;
assign w13186 = (~w12588 & w34874) | (~w12588 & w34875) | (w34874 & w34875);
assign w13187 = (~w12998 & w34876) | (~w12998 & w34877) | (w34876 & w34877);
assign w13188 = (w12998 & w34878) | (w12998 & w34879) | (w34878 & w34879);
assign w13189 = ~w13187 & ~w13188;
assign w13190 = (w12588 & w34880) | (w12588 & w34881) | (w34880 & w34881);
assign w13191 = ~w13186 & ~w13190;
assign w13192 = w13013 & w34882;
assign w13193 = (~w12588 & w34883) | (~w12588 & w34884) | (w34883 & w34884);
assign w13194 = (w12588 & w34885) | (w12588 & w34886) | (w34885 & w34886);
assign w13195 = ~w13193 & ~w13194;
assign w13196 = w13172 & w13195;
assign w13197 = ~w13172 & ~w13195;
assign w13198 = ~w13196 & ~w13197;
assign w13199 = ~w12601 & w13007;
assign w13200 = w12598 & ~w13199;
assign w13201 = (w12944 & w34887) | (w12944 & w34888) | (w34887 & w34888);
assign w13202 = ~w13200 & ~w13201;
assign w13203 = w13191 & ~w13198;
assign w13204 = (~w13201 & w34890) | (~w13201 & w34891) | (w34890 & w34891);
assign w13205 = ~w13198 & ~w13202;
assign w13206 = (~w13191 & ~w13013) | (~w13191 & w34892) | (~w13013 & w34892);
assign w13207 = (w13204 & w13205) | (w13204 & w34893) | (w13205 & w34893);
assign w13208 = ~w13181 & ~w13182;
assign w13209 = ~w13178 & w13208;
assign w13210 = (w13209 & ~w13207) | (w13209 & w34894) | (~w13207 & w34894);
assign w13211 = a_29 & ~w13210;
assign w13212 = (~w13207 & w34895) | (~w13207 & w34896) | (w34895 & w34896);
assign w13213 = ~w13211 & ~w13212;
assign w13214 = w13150 & w13213;
assign w13215 = (w13029 & w13214) | (w13029 & w34897) | (w13214 & w34897);
assign w13216 = ~w13027 & ~w13215;
assign w13217 = ~a_26 & ~w15;
assign w13218 = ~w49 & ~w13217;
assign w13219 = w3900 & w34899;
assign w13220 = ~w16 & ~w85;
assign w13221 = ~w265 & w13220;
assign w13222 = w840 & w13221;
assign w13223 = w1217 & w34900;
assign w13224 = w1306 & w34901;
assign w13225 = ~w663 & ~w13224;
assign w13226 = w663 & w13224;
assign w13227 = ~w13225 & ~w13226;
assign w13228 = w13218 & w13227;
assign w13229 = ~w13218 & ~w13227;
assign w13230 = ~w13228 & ~w13229;
assign w13231 = (w13024 & w34902) | (w13024 & w34903) | (w34902 & w34903);
assign w13232 = (~w13024 & w34904) | (~w13024 & w34905) | (w34904 & w34905);
assign w13233 = ~w13231 & ~w13232;
assign w13234 = ~w13174 & w34906;
assign w13235 = ~w13011 & w34907;
assign w13236 = w1399 & w12598;
assign w13237 = ~w13201 & w34908;
assign w13238 = ~w13205 & w34909;
assign w13239 = ~w13235 & w34910;
assign w13240 = ~w13238 & w13239;
assign w13241 = w13233 & ~w13240;
assign w13242 = ~w13233 & w13240;
assign w13243 = ~w13241 & ~w13242;
assign w13244 = w13177 & ~w13183;
assign w13245 = (w13201 & w34913) | (w13201 & w34914) | (w34913 & w34914);
assign w13246 = ~w4068 & ~w4446;
assign w13247 = (w13246 & ~w13177) | (w13246 & w34915) | (~w13177 & w34915);
assign w13248 = ~w13245 & w34916;
assign w13249 = (a_29 & w13245) | (a_29 & w34917) | (w13245 & w34917);
assign w13250 = ~w13248 & ~w13249;
assign w13251 = w13243 & w13250;
assign w13252 = ~w13243 & ~w13250;
assign w13253 = ~w13251 & ~w13252;
assign w13254 = w13216 & ~w13253;
assign w13255 = ~w13216 & w13253;
assign w13256 = ~w13254 & ~w13255;
assign w13257 = w4068 & w13177;
assign w13258 = ~w13174 & w34918;
assign w13259 = (~w13173 & w34919) | (~w13173 & w34920) | (w34919 & w34920);
assign w13260 = w4446 & ~w13259;
assign w13261 = w13177 & w13180;
assign w13262 = (w13201 & w34923) | (w13201 & w34924) | (w34923 & w34924);
assign w13263 = (~w13201 & w34925) | (~w13201 & w34926) | (w34925 & w34926);
assign w13264 = ~w13262 & ~w13263;
assign w13265 = ~w13258 & ~w13260;
assign w13266 = ~w13257 & w13265;
assign w13267 = (w13266 & w13264) | (w13266 & w34927) | (w13264 & w34927);
assign w13268 = ~a_29 & w13267;
assign w13269 = (~w13264 & w34928) | (~w13264 & w34929) | (w34928 & w34929);
assign w13270 = ~w13268 & w34930;
assign w13271 = ~w13214 & w34931;
assign w13272 = ~w13215 & ~w13271;
assign w13273 = (w13218 & w13268) | (w13218 & w34932) | (w13268 & w34932);
assign w13274 = ~w13270 & ~w13273;
assign w13275 = w13272 & w13274;
assign w13276 = (~w13270 & ~w13272) | (~w13270 & w34933) | (~w13272 & w34933);
assign w13277 = w13256 & ~w13276;
assign w13278 = ~w13256 & w13276;
assign w13279 = ~w13277 & ~w13278;
assign w13280 = (w13126 & w34934) | (w13126 & w34935) | (w34934 & w34935);
assign w13281 = ~w13130 & ~w13280;
assign w13282 = w668 & w12604;
assign w13283 = ~w12589 & w34936;
assign w13284 = (w1399 & w12616) | (w1399 & w34937) | (w12616 & w34937);
assign w13285 = ~w12608 & ~w12946;
assign w13286 = ~w12944 & w34938;
assign w13287 = (~w13285 & w12944) | (~w13285 & w34939) | (w12944 & w34939);
assign w13288 = ~w13286 & ~w13287;
assign w13289 = ~w13283 & ~w13284;
assign w13290 = ~w13282 & w13289;
assign w13291 = (w13290 & w13288) | (w13290 & w34940) | (w13288 & w34940);
assign w13292 = w13281 & ~w13291;
assign w13293 = ~w13281 & w13291;
assign w13294 = ~w13292 & ~w13293;
assign w13295 = ~w13011 & w34941;
assign w13296 = w4068 & w12598;
assign w13297 = w3957 & w12601;
assign w13298 = ~w13296 & ~w13297;
assign w13299 = ~w13295 & w13298;
assign w13300 = (w13299 & w13021) | (w13299 & w34942) | (w13021 & w34942);
assign w13301 = a_29 & ~w13300;
assign w13302 = (w13021 & w34943) | (w13021 & w34944) | (w34943 & w34944);
assign w13303 = ~w13301 & ~w13302;
assign w13304 = w13294 & w13303;
assign w13305 = ~w13135 & w13143;
assign w13306 = ~w13144 & ~w13305;
assign w13307 = (w13306 & w13304) | (w13306 & w34945) | (w13304 & w34945);
assign w13308 = ~w13304 & w34946;
assign w13309 = ~w13307 & ~w13308;
assign w13310 = ~w13174 & w34947;
assign w13311 = ~w13011 & w34948;
assign w13312 = w3957 & w12598;
assign w13313 = ~w13205 & w34949;
assign w13314 = ~w13311 & w34950;
assign w13315 = (a_29 & w13313) | (a_29 & w34951) | (w13313 & w34951);
assign w13316 = ~w13313 & w34952;
assign w13317 = ~w13315 & ~w13316;
assign w13318 = w13309 & w13317;
assign w13319 = (~w13307 & ~w13309) | (~w13307 & w34953) | (~w13309 & w34953);
assign w13320 = ~w13150 & ~w13213;
assign w13321 = ~w13214 & ~w13320;
assign w13322 = ~w13319 & w13321;
assign w13323 = w13319 & ~w13321;
assign w13324 = ~w13322 & ~w13323;
assign w13325 = (~w13173 & w34956) | (~w13173 & w34957) | (w34956 & w34957);
assign w13326 = ~a_26 & w13325;
assign w13327 = (w13173 & w34958) | (w13173 & w34959) | (w34958 & w34959);
assign w13328 = ~w13326 & ~w13327;
assign w13329 = w13324 & w13328;
assign w13330 = (~w13322 & ~w13324) | (~w13322 & w34960) | (~w13324 & w34960);
assign w13331 = ~w13272 & ~w13274;
assign w13332 = ~w13275 & ~w13331;
assign w13333 = ~w13330 & w13332;
assign w13334 = (~w13123 & w34961) | (~w13123 & w34962) | (w34961 & w34962);
assign w13335 = ~w13127 & ~w13334;
assign w13336 = ~w94 & ~w589;
assign w13337 = ~w180 & ~w213;
assign w13338 = ~w563 & w13337;
assign w13339 = w908 & w2034;
assign w13340 = w2481 & w2966;
assign w13341 = w4127 & w13336;
assign w13342 = w13340 & w13341;
assign w13343 = w13338 & w13339;
assign w13344 = w3760 & w13343;
assign w13345 = w211 & w13342;
assign w13346 = w13344 & w13345;
assign w13347 = w3253 & w13346;
assign w13348 = ~w68 & ~w95;
assign w13349 = ~w75 & ~w196;
assign w13350 = ~w619 & w13349;
assign w13351 = w3214 & w13350;
assign w13352 = w711 & w1293;
assign w13353 = w2786 & w3427;
assign w13354 = w3772 & w13348;
assign w13355 = w13353 & w13354;
assign w13356 = w4345 & w13352;
assign w13357 = w4543 & w4848;
assign w13358 = w13356 & w13357;
assign w13359 = w2056 & w13355;
assign w13360 = w13351 & w13359;
assign w13361 = w3245 & w13358;
assign w13362 = w13360 & w13361;
assign w13363 = w5543 & w13362;
assign w13364 = w13347 & w13363;
assign w13365 = w13081 & ~w13364;
assign w13366 = ~w13081 & w13364;
assign w13367 = ~w13365 & ~w13366;
assign w13368 = (w668 & w12612) | (w668 & w34963) | (w12612 & w34963);
assign w13369 = ~w12914 & w34964;
assign w13370 = ~w12930 & w34965;
assign w13371 = (~w12904 & w34966) | (~w12904 & w34967) | (w34966 & w34967);
assign w13372 = ~w12932 & ~w12935;
assign w13373 = ~w13371 & w13372;
assign w13374 = w13371 & ~w13372;
assign w13375 = ~w13373 & ~w13374;
assign w13376 = ~w13369 & ~w13370;
assign w13377 = ~w13368 & w13376;
assign w13378 = (w13377 & ~w13375) | (w13377 & w34968) | (~w13375 & w34968);
assign w13379 = w13367 & ~w13378;
assign w13380 = w13111 & ~w13113;
assign w13381 = ~w13114 & ~w13380;
assign w13382 = (w13378 & w34970) | (w13378 & w34971) | (w34970 & w34971);
assign w13383 = (~w13378 & w34972) | (~w13378 & w34973) | (w34972 & w34973);
assign w13384 = ~w13382 & ~w13383;
assign w13385 = (w668 & w12616) | (w668 & w34974) | (w12616 & w34974);
assign w13386 = (w1327 & w12612) | (w1327 & w34975) | (w12612 & w34975);
assign w13387 = ~w12930 & w34976;
assign w13388 = ~w12933 & w34977;
assign w13389 = ~w12939 & ~w13388;
assign w13390 = ~w13386 & ~w13387;
assign w13391 = ~w13385 & w13390;
assign w13392 = (w13391 & ~w13389) | (w13391 & w34978) | (~w13389 & w34978);
assign w13393 = w13384 & w13392;
assign w13394 = (~w13382 & ~w13384) | (~w13382 & w34979) | (~w13384 & w34979);
assign w13395 = w13335 & w13394;
assign w13396 = ~w13335 & ~w13394;
assign w13397 = ~w13395 & ~w13396;
assign w13398 = w4446 & w12598;
assign w13399 = w4068 & w12601;
assign w13400 = w3957 & w12604;
assign w13401 = ~w13399 & ~w13400;
assign w13402 = ~w13398 & w13401;
assign w13403 = (w13402 & ~w12961) | (w13402 & w34980) | (~w12961 & w34980);
assign w13404 = ~a_29 & w13403;
assign w13405 = (w12961 & w34981) | (w12961 & w34982) | (w34981 & w34982);
assign w13406 = ~w13404 & ~w13405;
assign w13407 = w13397 & w13406;
assign w13408 = (~w13395 & ~w13397) | (~w13395 & w34983) | (~w13397 & w34983);
assign w13409 = ~w13294 & ~w13303;
assign w13410 = ~w13304 & ~w13409;
assign w13411 = ~w13408 & w13410;
assign w13412 = w13408 & ~w13410;
assign w13413 = ~w13411 & ~w13412;
assign w13414 = w4638 & w13177;
assign w13415 = ~w13174 & w34984;
assign w13416 = (w13173 & w34985) | (w13173 & w34986) | (w34985 & w34986);
assign w13417 = ~w13415 & ~w13416;
assign w13418 = ~w13414 & w13417;
assign w13419 = (w13418 & w13264) | (w13418 & w34987) | (w13264 & w34987);
assign w13420 = a_26 & ~w13419;
assign w13421 = (w13264 & w34988) | (w13264 & w34989) | (w34988 & w34989);
assign w13422 = ~w13420 & ~w13421;
assign w13423 = w13413 & w13422;
assign w13424 = (~w13411 & ~w13413) | (~w13411 & w34990) | (~w13413 & w34990);
assign w13425 = ~w518 & w13177;
assign w13426 = (w13201 & w34993) | (w13201 & w34994) | (w34993 & w34994);
assign w13427 = (~w13173 & w34995) | (~w13173 & w34996) | (w34995 & w34996);
assign w13428 = ~w13425 & w13427;
assign w13429 = (a_26 & w13426) | (a_26 & w34997) | (w13426 & w34997);
assign w13430 = ~w13426 & w34998;
assign w13431 = ~w13429 & ~w13430;
assign w13432 = ~w13424 & w13431;
assign w13433 = ~w13309 & ~w13317;
assign w13434 = ~w13318 & ~w13433;
assign w13435 = w13424 & ~w13431;
assign w13436 = ~w13432 & ~w13435;
assign w13437 = w13434 & w13436;
assign w13438 = (~w13432 & ~w13436) | (~w13432 & w34999) | (~w13436 & w34999);
assign w13439 = ~w13324 & ~w13328;
assign w13440 = ~w13329 & ~w13439;
assign w13441 = ~w13438 & w13440;
assign w13442 = w13438 & ~w13440;
assign w13443 = ~w13441 & ~w13442;
assign w13444 = ~w13397 & ~w13406;
assign w13445 = ~w13407 & ~w13444;
assign w13446 = ~w13384 & ~w13392;
assign w13447 = ~w13393 & ~w13446;
assign w13448 = ~w116 & ~w282;
assign w13449 = w1725 & w13448;
assign w13450 = w2177 & w2555;
assign w13451 = w13449 & w13450;
assign w13452 = ~w422 & ~w475;
assign w13453 = ~w23 & ~w94;
assign w13454 = ~w447 & ~w544;
assign w13455 = w13453 & w13454;
assign w13456 = w549 & w990;
assign w13457 = w1772 & w1853;
assign w13458 = w2402 & w2454;
assign w13459 = w2943 & w13452;
assign w13460 = w13458 & w13459;
assign w13461 = w13456 & w13457;
assign w13462 = w2330 & w13455;
assign w13463 = w2741 & w13462;
assign w13464 = w13460 & w13461;
assign w13465 = w13451 & w13464;
assign w13466 = w5598 & w13463;
assign w13467 = w13465 & w13466;
assign w13468 = w2859 & w13467;
assign w13469 = w4309 & w13468;
assign w13470 = w2576 & w2772;
assign w13471 = ~w88 & ~w238;
assign w13472 = ~w251 & ~w312;
assign w13473 = w13471 & w13472;
assign w13474 = w1103 & w1309;
assign w13475 = w2250 & w3517;
assign w13476 = w13474 & w13475;
assign w13477 = w361 & w13473;
assign w13478 = w1108 & w6572;
assign w13479 = w13470 & w13478;
assign w13480 = w13476 & w13477;
assign w13481 = w13479 & w13480;
assign w13482 = w2629 & w13481;
assign w13483 = w13067 & w13482;
assign w13484 = w852 & w5200;
assign w13485 = w13483 & w13484;
assign w13486 = ~w13469 & ~w13485;
assign w13487 = a_17 & ~w6058;
assign w13488 = ~a_16 & w6052;
assign w13489 = (~w13488 & w6058) | (~w13488 & w35000) | (w6058 & w35000);
assign w13490 = w13469 & w13485;
assign w13491 = ~w13486 & ~w13490;
assign w13492 = ~w13489 & w13491;
assign w13493 = (~w13486 & ~w13491) | (~w13486 & w35001) | (~w13491 & w35001);
assign w13494 = w13081 & ~w13493;
assign w13495 = ~w13081 & w13493;
assign w13496 = ~w13494 & ~w13495;
assign w13497 = ~w12930 & w35002;
assign w13498 = w1399 & ~w12910;
assign w13499 = ~w12914 & w35003;
assign w13500 = (w12904 & w35004) | (w12904 & w35005) | (w35004 & w35005);
assign w13501 = w12927 & ~w13500;
assign w13502 = ~w13501 & w35006;
assign w13503 = ~w13498 & ~w13499;
assign w13504 = ~w13497 & w13503;
assign w13505 = (w13496 & w13502) | (w13496 & w35007) | (w13502 & w35007);
assign w13506 = (~w13502 & w35008) | (~w13502 & w35009) | (w35008 & w35009);
assign w13507 = (~w13375 & w35010) | (~w13375 & w35011) | (w35010 & w35011);
assign w13508 = ~w13379 & w35012;
assign w13509 = (w13506 & w13379) | (w13506 & w35013) | (w13379 & w35013);
assign w13510 = ~w13508 & ~w13509;
assign w13511 = w13489 & ~w13491;
assign w13512 = ~w13492 & ~w13511;
assign w13513 = ~w12914 & w35014;
assign w13514 = w1327 & ~w12910;
assign w13515 = ~w12905 & w35015;
assign w13516 = ~w12917 & ~w12922;
assign w13517 = (w12920 & ~w12904) | (w12920 & w35016) | (~w12904 & w35016);
assign w13518 = w13516 & w13517;
assign w13519 = (w12904 & w35017) | (w12904 & w35018) | (w35017 & w35018);
assign w13520 = (w1478 & w13518) | (w1478 & w35019) | (w13518 & w35019);
assign w13521 = ~w13514 & ~w13515;
assign w13522 = ~w13513 & w13521;
assign w13523 = (w13512 & w13520) | (w13512 & w35020) | (w13520 & w35020);
assign w13524 = ~w260 & ~w447;
assign w13525 = ~w547 & w13524;
assign w13526 = w1199 & w1691;
assign w13527 = w1822 & w2438;
assign w13528 = w3575 & w13527;
assign w13529 = w13525 & w13526;
assign w13530 = w187 & w13529;
assign w13531 = w13528 & w13530;
assign w13532 = w2397 & w3517;
assign w13533 = w209 & ~w649;
assign w13534 = w444 & w13533;
assign w13535 = ~w266 & w1533;
assign w13536 = w3248 & w13082;
assign w13537 = w13535 & w13536;
assign w13538 = w2930 & w3276;
assign w13539 = w6573 & w13532;
assign w13540 = w13538 & w13539;
assign w13541 = w1013 & w13537;
assign w13542 = w13540 & w13541;
assign w13543 = w13531 & w13542;
assign w13544 = w2588 & w13543;
assign w13545 = w13534 & w13544;
assign w13546 = w13469 & ~w13545;
assign w13547 = ~w72 & ~w530;
assign w13548 = w865 & w5432;
assign w13549 = ~w89 & ~w356;
assign w13550 = ~w149 & ~w216;
assign w13551 = w1098 & w13550;
assign w13552 = w1344 & w1425;
assign w13553 = w2796 & w13547;
assign w13554 = w13549 & w13553;
assign w13555 = w13551 & w13552;
assign w13556 = w5590 & w13555;
assign w13557 = w13554 & w13556;
assign w13558 = w2107 & w2429;
assign w13559 = w13557 & w13558;
assign w13560 = w3759 & w13559;
assign w13561 = w13548 & w13560;
assign w13562 = w853 & w941;
assign w13563 = ~w98 & ~w563;
assign w13564 = ~w265 & ~w325;
assign w13565 = ~w68 & ~w776;
assign w13566 = ~w208 & ~w385;
assign w13567 = w1810 & w13566;
assign w13568 = w13564 & w13565;
assign w13569 = w13567 & w13568;
assign w13570 = ~w181 & ~w319;
assign w13571 = w2240 & w13570;
assign w13572 = w2773 & w13563;
assign w13573 = w13571 & w13572;
assign w13574 = w1318 & w1825;
assign w13575 = w4901 & w13562;
assign w13576 = w13574 & w13575;
assign w13577 = w4273 & w13573;
assign w13578 = w13569 & w13577;
assign w13579 = w3441 & w13576;
assign w13580 = w13578 & w13579;
assign w13581 = w3416 & w13580;
assign w13582 = w6524 & w13581;
assign w13583 = ~w13561 & ~w13582;
assign w13584 = a_14 & ~w6445;
assign w13585 = ~a_13 & w6439;
assign w13586 = (~w13585 & w6445) | (~w13585 & w35021) | (w6445 & w35021);
assign w13587 = w13561 & w13582;
assign w13588 = ~w13583 & ~w13587;
assign w13589 = ~w13586 & w13588;
assign w13590 = (~w13583 & ~w13588) | (~w13583 & w35022) | (~w13588 & w35022);
assign w13591 = w13545 & ~w13590;
assign w13592 = ~w13545 & w13590;
assign w13593 = ~w13591 & ~w13592;
assign w13594 = ~w12905 & w35023;
assign w13595 = ~w12892 & w35024;
assign w13596 = w1399 & ~w12878;
assign w13597 = (w12862 & w35025) | (w12862 & w35026) | (w35025 & w35026);
assign w13598 = w12902 & ~w13597;
assign w13599 = ~w13598 & w35027;
assign w13600 = ~w13595 & ~w13596;
assign w13601 = ~w13594 & w13600;
assign w13602 = (w13593 & w13599) | (w13593 & w35028) | (w13599 & w35028);
assign w13603 = ~w13469 & w13545;
assign w13604 = ~w13546 & ~w13603;
assign w13605 = (w13599 & w35031) | (w13599 & w35032) | (w35031 & w35032);
assign w13606 = (~w13599 & w35033) | (~w13599 & w35034) | (w35033 & w35034);
assign w13607 = ~w13520 & w35035;
assign w13608 = ~w13523 & ~w13607;
assign w13609 = ~w13606 & w13608;
assign w13610 = (~w13523 & ~w13608) | (~w13523 & w35036) | (~w13608 & w35036);
assign w13611 = ~w13502 & w35037;
assign w13612 = ~w13505 & ~w13611;
assign w13613 = ~w13610 & w13612;
assign w13614 = w13610 & ~w13612;
assign w13615 = ~w13613 & ~w13614;
assign w13616 = (w4068 & w12616) | (w4068 & w35038) | (w12616 & w35038);
assign w13617 = (w3957 & w12612) | (w3957 & w35039) | (w12612 & w35039);
assign w13618 = ~w12589 & w35040;
assign w13619 = ~w13616 & ~w13617;
assign w13620 = ~w13618 & w13619;
assign w13621 = (w13620 & ~w13123) | (w13620 & w35041) | (~w13123 & w35041);
assign w13622 = a_29 & ~w13621;
assign w13623 = (~w13123 & w35042) | (~w13123 & w35043) | (w35042 & w35043);
assign w13624 = ~w13622 & ~w13623;
assign w13625 = w13615 & w13624;
assign w13626 = (~w13613 & ~w13615) | (~w13613 & w35044) | (~w13615 & w35044);
assign w13627 = w13510 & ~w13626;
assign w13628 = (w13626 & w35046) | (w13626 & w35047) | (w35046 & w35047);
assign w13629 = (~w13626 & w35048) | (~w13626 & w35049) | (w35048 & w35049);
assign w13630 = ~w13628 & ~w13629;
assign w13631 = w4446 & w12601;
assign w13632 = w4068 & w12604;
assign w13633 = ~w12589 & w35050;
assign w13634 = ~w13632 & ~w13633;
assign w13635 = ~w13631 & w13634;
assign w13636 = (w13635 & w13140) | (w13635 & w35051) | (w13140 & w35051);
assign w13637 = ~a_29 & w13636;
assign w13638 = (~w13140 & w35052) | (~w13140 & w35053) | (w35052 & w35053);
assign w13639 = ~w13637 & ~w13638;
assign w13640 = w13630 & ~w13639;
assign w13641 = (~w13628 & ~w13630) | (~w13628 & w35054) | (~w13630 & w35054);
assign w13642 = ~w13445 & ~w13641;
assign w13643 = w13445 & w13641;
assign w13644 = ~w13642 & ~w13643;
assign w13645 = w4666 & w13177;
assign w13646 = ~w13011 & w35055;
assign w13647 = ~w13174 & w35056;
assign w13648 = ~w13646 & ~w13647;
assign w13649 = ~w13645 & w13648;
assign w13650 = (w13649 & ~w13207) | (w13649 & w35057) | (~w13207 & w35057);
assign w13651 = ~a_26 & w13650;
assign w13652 = (w13207 & w35058) | (w13207 & w35059) | (w35058 & w35059);
assign w13653 = ~w13651 & ~w13652;
assign w13654 = w13644 & ~w13653;
assign w13655 = (~w13642 & ~w13644) | (~w13642 & w35060) | (~w13644 & w35060);
assign w13656 = w511 & w13655;
assign w13657 = ~w13413 & ~w13422;
assign w13658 = ~w13423 & ~w13657;
assign w13659 = ~w511 & ~w13655;
assign w13660 = ~w13656 & ~w13659;
assign w13661 = w13658 & w13660;
assign w13662 = (~w13656 & ~w13660) | (~w13656 & w35061) | (~w13660 & w35061);
assign w13663 = ~w13434 & ~w13436;
assign w13664 = ~w13437 & ~w13663;
assign w13665 = ~w13662 & w13664;
assign w13666 = w13662 & ~w13664;
assign w13667 = ~w13665 & ~w13666;
assign w13668 = ~w13658 & ~w13660;
assign w13669 = ~w13661 & ~w13668;
assign w13670 = ~w13644 & w13653;
assign w13671 = ~w13654 & ~w13670;
assign w13672 = ~w13630 & w13639;
assign w13673 = ~w13640 & ~w13672;
assign w13674 = ~w13174 & w35062;
assign w13675 = ~w518 & w12598;
assign w13676 = ~w13011 & w35063;
assign w13677 = ~w13205 & w35064;
assign w13678 = ~w13676 & w35065;
assign w13679 = ~w13677 & w35066;
assign w13680 = (~a_26 & w13677) | (~a_26 & w35067) | (w13677 & w35067);
assign w13681 = ~w13679 & ~w13680;
assign w13682 = ~w13673 & ~w13681;
assign w13683 = ~w13510 & w13626;
assign w13684 = ~w13627 & ~w13683;
assign w13685 = w4446 & w12604;
assign w13686 = ~w12589 & w35068;
assign w13687 = (w3957 & w12616) | (w3957 & w35069) | (w12616 & w35069);
assign w13688 = ~w13686 & ~w13687;
assign w13689 = ~w13685 & w13688;
assign w13690 = (w13689 & w13288) | (w13689 & w35070) | (w13288 & w35070);
assign w13691 = ~a_29 & w13690;
assign w13692 = (~w13288 & w35071) | (~w13288 & w35072) | (w35071 & w35072);
assign w13693 = ~w13691 & ~w13692;
assign w13694 = w13684 & w13693;
assign w13695 = ~w13684 & ~w13693;
assign w13696 = ~w13694 & ~w13695;
assign w13697 = ~w13011 & w35073;
assign w13698 = ~w518 & w12601;
assign w13699 = w4638 & w12598;
assign w13700 = ~w13698 & ~w13699;
assign w13701 = ~w13697 & w13700;
assign w13702 = (w13701 & w13021) | (w13701 & w35074) | (w13021 & w35074);
assign w13703 = ~a_26 & w13702;
assign w13704 = (~w13021 & w35075) | (~w13021 & w35076) | (w35075 & w35076);
assign w13705 = ~w13703 & ~w13704;
assign w13706 = w13696 & w13705;
assign w13707 = (~w13694 & ~w13696) | (~w13694 & w35077) | (~w13696 & w35077);
assign w13708 = w13673 & w13681;
assign w13709 = ~w13682 & ~w13708;
assign w13710 = ~w13707 & w13709;
assign w13711 = (~w13682 & ~w13709) | (~w13682 & w35078) | (~w13709 & w35078);
assign w13712 = w13671 & w13711;
assign w13713 = ~w13671 & ~w13711;
assign w13714 = ~w13712 & ~w13713;
assign w13715 = (~w13173 & w35081) | (~w13173 & w35082) | (w35081 & w35082);
assign w13716 = (~w13173 & w35083) | (~w13173 & w35084) | (w35083 & w35084);
assign w13717 = ~w13715 & w13716;
assign w13718 = ~w509 & ~w13717;
assign w13719 = w13714 & ~w13718;
assign w13720 = (~w13712 & ~w13714) | (~w13712 & w35085) | (~w13714 & w35085);
assign w13721 = w13669 & w13720;
assign w13722 = ~w13669 & ~w13720;
assign w13723 = ~w13599 & w35086;
assign w13724 = ~w13602 & ~w13723;
assign w13725 = w934 & w4714;
assign w13726 = ~w261 & ~w589;
assign w13727 = w1191 & w13726;
assign w13728 = w2191 & w13727;
assign w13729 = w986 & w2035;
assign w13730 = ~w394 & ~w468;
assign w13731 = w449 & w13730;
assign w13732 = w817 & w2798;
assign w13733 = w3212 & w13732;
assign w13734 = w1015 & w13731;
assign w13735 = w1407 & w2120;
assign w13736 = w3798 & w13729;
assign w13737 = w13735 & w13736;
assign w13738 = w13733 & w13734;
assign w13739 = w13728 & w13738;
assign w13740 = w13737 & w13739;
assign w13741 = ~w313 & ~w458;
assign w13742 = w43 & ~w543;
assign w13743 = w13741 & w13742;
assign w13744 = w1345 & w3457;
assign w13745 = w4084 & w4366;
assign w13746 = w13744 & w13745;
assign w13747 = w13743 & w13746;
assign w13748 = ~w71 & ~w337;
assign w13749 = w584 & w13748;
assign w13750 = w1813 & w4363;
assign w13751 = w5368 & w13750;
assign w13752 = w2806 & w13749;
assign w13753 = w3732 & w13725;
assign w13754 = w13752 & w13753;
assign w13755 = w2884 & w13751;
assign w13756 = w4092 & w13755;
assign w13757 = w13754 & w13756;
assign w13758 = w13747 & w13757;
assign w13759 = w3078 & w13740;
assign w13760 = w13758 & w13759;
assign w13761 = w13561 & ~w13760;
assign w13762 = ~w13561 & w13760;
assign w13763 = ~w13761 & ~w13762;
assign w13764 = w668 & ~w12878;
assign w13765 = w1327 & w12874;
assign w13766 = w1399 & w12869;
assign w13767 = ~w12879 & ~w12887;
assign w13768 = (w12885 & w12862) | (w12885 & w35087) | (w12862 & w35087);
assign w13769 = (w13767 & w13768) | (w13767 & w35088) | (w13768 & w35088);
assign w13770 = ~w13768 & w35089;
assign w13771 = ~w13769 & ~w13770;
assign w13772 = ~w13765 & ~w13766;
assign w13773 = ~w13764 & w13772;
assign w13774 = (w13773 & ~w13771) | (w13773 & w35090) | (~w13771 & w35090);
assign w13775 = w13763 & ~w13774;
assign w13776 = w13586 & ~w13588;
assign w13777 = ~w13589 & ~w13776;
assign w13778 = (w13774 & w35092) | (w13774 & w35093) | (w35092 & w35093);
assign w13779 = (~w13774 & w35094) | (~w13774 & w35095) | (w35094 & w35095);
assign w13780 = ~w13778 & ~w13779;
assign w13781 = ~w12892 & w35096;
assign w13782 = w1327 & ~w12878;
assign w13783 = w1399 & w12874;
assign w13784 = ~w12895 & ~w12897;
assign w13785 = (w12862 & w35099) | (w12862 & w35100) | (w35099 & w35100);
assign w13786 = (~w12862 & w35101) | (~w12862 & w35102) | (w35101 & w35102);
assign w13787 = ~w13785 & ~w13786;
assign w13788 = ~w13782 & ~w13783;
assign w13789 = ~w13781 & w13788;
assign w13790 = (w13789 & ~w13787) | (w13789 & w35103) | (~w13787 & w35103);
assign w13791 = w13780 & w13790;
assign w13792 = (~w13778 & ~w13780) | (~w13778 & w35104) | (~w13780 & w35104);
assign w13793 = w13724 & w13792;
assign w13794 = ~w13724 & ~w13792;
assign w13795 = ~w13793 & ~w13794;
assign w13796 = ~w12930 & w35105;
assign w13797 = w3957 & ~w12910;
assign w13798 = ~w12914 & w35106;
assign w13799 = ~w13501 & w35107;
assign w13800 = ~w13797 & ~w13798;
assign w13801 = ~w13796 & w13800;
assign w13802 = ~w13799 & w35108;
assign w13803 = (a_29 & w13799) | (a_29 & w35109) | (w13799 & w35109);
assign w13804 = ~w13802 & ~w13803;
assign w13805 = w13795 & w13804;
assign w13806 = (~w13793 & ~w13795) | (~w13793 & w35110) | (~w13795 & w35110);
assign w13807 = (~w13599 & w35111) | (~w13599 & w35112) | (w35111 & w35112);
assign w13808 = ~w13605 & ~w13807;
assign w13809 = ~w12905 & w35113;
assign w13810 = w668 & ~w12910;
assign w13811 = ~w12892 & w35114;
assign w13812 = ~w12911 & ~w12918;
assign w13813 = (w13812 & w12904) | (w13812 & w35115) | (w12904 & w35115);
assign w13814 = ~w12904 & w35116;
assign w13815 = ~w13813 & ~w13814;
assign w13816 = w1478 & w13815;
assign w13817 = ~w13810 & w35117;
assign w13818 = ~w13816 & w13817;
assign w13819 = w13808 & ~w13818;
assign w13820 = ~w13808 & w13818;
assign w13821 = ~w13819 & ~w13820;
assign w13822 = (w4446 & w12612) | (w4446 & w35118) | (w12612 & w35118);
assign w13823 = ~w12914 & w35119;
assign w13824 = ~w12930 & w35120;
assign w13825 = ~w13823 & ~w13824;
assign w13826 = ~w13822 & w13825;
assign w13827 = (w13826 & ~w13375) | (w13826 & w35121) | (~w13375 & w35121);
assign w13828 = ~a_29 & w13827;
assign w13829 = (w13375 & w35122) | (w13375 & w35123) | (w35122 & w35123);
assign w13830 = ~w13828 & ~w13829;
assign w13831 = w13821 & w13830;
assign w13832 = ~w13821 & ~w13830;
assign w13833 = ~w13831 & ~w13832;
assign w13834 = ~w13806 & w13833;
assign w13835 = w13806 & ~w13833;
assign w13836 = ~w13834 & ~w13835;
assign w13837 = w4666 & w12604;
assign w13838 = (~w518 & w12616) | (~w518 & w35124) | (w12616 & w35124);
assign w13839 = ~w12589 & w35125;
assign w13840 = ~w13838 & ~w13839;
assign w13841 = ~w13837 & w13840;
assign w13842 = (w13841 & w13288) | (w13841 & w35126) | (w13288 & w35126);
assign w13843 = a_26 & ~w13842;
assign w13844 = (w13288 & w35127) | (w13288 & w35128) | (w35127 & w35128);
assign w13845 = ~w13843 & ~w13844;
assign w13846 = w13836 & w13845;
assign w13847 = (~w13834 & ~w13836) | (~w13834 & w35129) | (~w13836 & w35129);
assign w13848 = ~w13819 & ~w13831;
assign w13849 = w13606 & ~w13608;
assign w13850 = ~w13609 & ~w13849;
assign w13851 = w13848 & ~w13850;
assign w13852 = ~w13848 & w13850;
assign w13853 = ~w13851 & ~w13852;
assign w13854 = (w4446 & w12616) | (w4446 & w35130) | (w12616 & w35130);
assign w13855 = (w4068 & w12612) | (w4068 & w35131) | (w12612 & w35131);
assign w13856 = ~w12930 & w35132;
assign w13857 = ~w13855 & ~w13856;
assign w13858 = ~w13854 & w13857;
assign w13859 = (w13858 & ~w13389) | (w13858 & w35133) | (~w13389 & w35133);
assign w13860 = ~a_29 & w13859;
assign w13861 = (w13389 & w35134) | (w13389 & w35135) | (w35134 & w35135);
assign w13862 = ~w13860 & ~w13861;
assign w13863 = w13853 & w13862;
assign w13864 = ~w13853 & ~w13862;
assign w13865 = ~w13863 & ~w13864;
assign w13866 = w4666 & w12601;
assign w13867 = ~w12589 & w35136;
assign w13868 = w4638 & w12604;
assign w13869 = ~w13867 & ~w13868;
assign w13870 = ~w13866 & w13869;
assign w13871 = (w13870 & w13140) | (w13870 & w35137) | (w13140 & w35137);
assign w13872 = a_26 & w13871;
assign w13873 = (~w13140 & w35138) | (~w13140 & w35139) | (w35138 & w35139);
assign w13874 = ~w13872 & ~w13873;
assign w13875 = w13865 & ~w13874;
assign w13876 = ~w13865 & w13874;
assign w13877 = ~w13875 & ~w13876;
assign w13878 = ~w13847 & w13877;
assign w13879 = w13847 & ~w13877;
assign w13880 = ~w13878 & ~w13879;
assign w13881 = ~w13174 & w35140;
assign w13882 = w5016 & w12598;
assign w13883 = ~w13011 & w35141;
assign w13884 = ~w13205 & w35142;
assign w13885 = ~w13883 & w35143;
assign w13886 = ~w13884 & w35144;
assign w13887 = (~a_23 & w13884) | (~a_23 & w35145) | (w13884 & w35145);
assign w13888 = ~w13886 & ~w13887;
assign w13889 = w13880 & ~w13888;
assign w13890 = ~w13780 & ~w13790;
assign w13891 = ~w13791 & ~w13890;
assign w13892 = ~w12914 & w35146;
assign w13893 = w4068 & ~w12910;
assign w13894 = ~w12905 & w35147;
assign w13895 = (w4070 & w13518) | (w4070 & w35148) | (w13518 & w35148);
assign w13896 = ~w13893 & ~w13894;
assign w13897 = ~w13892 & w13896;
assign w13898 = (a_29 & w13895) | (a_29 & w35149) | (w13895 & w35149);
assign w13899 = ~w13895 & w35150;
assign w13900 = ~w13898 & ~w13899;
assign w13901 = ~w13891 & w13900;
assign w13902 = ~w339 & w736;
assign w13903 = w1921 & w3847;
assign w13904 = w13902 & w13903;
assign w13905 = ~w147 & w573;
assign w13906 = w1374 & ~w1891;
assign w13907 = w4924 & w13906;
assign w13908 = w2560 & w13905;
assign w13909 = w3571 & w13908;
assign w13910 = w13907 & w13909;
assign w13911 = ~w113 & ~w619;
assign w13912 = ~w321 & w648;
assign w13913 = w820 & w1493;
assign w13914 = w2798 & w3676;
assign w13915 = w4151 & w13911;
assign w13916 = w13914 & w13915;
assign w13917 = w13912 & w13913;
assign w13918 = w3140 & w5170;
assign w13919 = w13917 & w13918;
assign w13920 = w4736 & w13916;
assign w13921 = w13904 & w13920;
assign w13922 = w13919 & w13921;
assign w13923 = w13910 & w13922;
assign w13924 = w1150 & w6167;
assign w13925 = w13923 & w13924;
assign w13926 = ~w30 & ~w85;
assign w13927 = w2008 & w2990;
assign w13928 = w13547 & w13926;
assign w13929 = w13927 & w13928;
assign w13930 = ~w568 & ~w818;
assign w13931 = ~w463 & w814;
assign w13932 = w2093 & w2404;
assign w13933 = w2873 & w3342;
assign w13934 = w13930 & w13933;
assign w13935 = w13931 & w13932;
assign w13936 = w1426 & w3735;
assign w13937 = w4851 & w13936;
assign w13938 = w13934 & w13935;
assign w13939 = w13929 & w13938;
assign w13940 = w13937 & w13939;
assign w13941 = w1657 & w2132;
assign w13942 = w5854 & w13941;
assign w13943 = w616 & w13940;
assign w13944 = w13942 & w13943;
assign w13945 = ~w13925 & ~w13944;
assign w13946 = a_11 & ~w7191;
assign w13947 = ~a_10 & w7185;
assign w13948 = (~w13947 & w7191) | (~w13947 & w35151) | (w7191 & w35151);
assign w13949 = w13925 & w13944;
assign w13950 = ~w13945 & ~w13949;
assign w13951 = ~w13948 & w13950;
assign w13952 = (~w13945 & ~w13950) | (~w13945 & w35152) | (~w13950 & w35152);
assign w13953 = w13561 & ~w13952;
assign w13954 = ~w13561 & w13952;
assign w13955 = ~w13953 & ~w13954;
assign w13956 = w668 & w12874;
assign w13957 = w1399 & ~w12860;
assign w13958 = w1327 & w12869;
assign w13959 = ~w12858 & w35153;
assign w13960 = (w12866 & w12858) | (w12866 & w35154) | (w12858 & w35154);
assign w13961 = ~w13959 & ~w13960;
assign w13962 = (~w13961 & w12862) | (~w13961 & w35155) | (w12862 & w35155);
assign w13963 = (w12884 & w12860) | (w12884 & w35156) | (w12860 & w35156);
assign w13964 = (~w12862 & w35157) | (~w12862 & w35158) | (w35157 & w35158);
assign w13965 = ~w13768 & ~w13964;
assign w13966 = w1478 & w13965;
assign w13967 = ~w13957 & w35159;
assign w13968 = (w13955 & w13966) | (w13955 & w35160) | (w13966 & w35160);
assign w13969 = (~w13966 & w35161) | (~w13966 & w35162) | (w35161 & w35162);
assign w13970 = (~w13771 & w35163) | (~w13771 & w35164) | (w35163 & w35164);
assign w13971 = ~w13775 & w35165;
assign w13972 = (w13969 & w13775) | (w13969 & w35166) | (w13775 & w35166);
assign w13973 = ~w13971 & ~w13972;
assign w13974 = w13948 & ~w13950;
assign w13975 = ~w13951 & ~w13974;
assign w13976 = w1399 & w12856;
assign w13977 = w668 & w12869;
assign w13978 = ~w12862 & w35167;
assign w13979 = ~w13962 & ~w13978;
assign w13980 = (~w13976 & w12860) | (~w13976 & w35168) | (w12860 & w35168);
assign w13981 = ~w13977 & w13980;
assign w13982 = (w13981 & ~w13979) | (w13981 & w35169) | (~w13979 & w35169);
assign w13983 = w13975 & ~w13982;
assign w13984 = w2417 & w5367;
assign w13985 = ~w159 & ~w1040;
assign w13986 = ~w173 & ~w316;
assign w13987 = w2975 & w13986;
assign w13988 = w343 & w756;
assign w13989 = w1071 & w1206;
assign w13990 = w2337 & w2707;
assign w13991 = w4157 & w13985;
assign w13992 = w13990 & w13991;
assign w13993 = w13988 & w13989;
assign w13994 = w2783 & w13984;
assign w13995 = w13993 & w13994;
assign w13996 = w1540 & w13992;
assign w13997 = w2662 & w13987;
assign w13998 = w13996 & w13997;
assign w13999 = w13995 & w13998;
assign w14000 = w3223 & w13999;
assign w14001 = w452 & w739;
assign w14002 = w1193 & w2083;
assign w14003 = w5370 & w13050;
assign w14004 = w14002 & w14003;
assign w14005 = w14001 & w14004;
assign w14006 = ~w217 & ~w1123;
assign w14007 = ~w447 & ~w996;
assign w14008 = w1293 & w14007;
assign w14009 = w1572 & w2499;
assign w14010 = w5186 & w14006;
assign w14011 = w14009 & w14010;
assign w14012 = w1535 & w14008;
assign w14013 = w3519 & w13729;
assign w14014 = w14012 & w14013;
assign w14015 = w14011 & w14014;
assign w14016 = w14005 & w14015;
assign w14017 = w4830 & w14016;
assign w14018 = w14000 & w14017;
assign w14019 = w13925 & ~w14018;
assign w14020 = ~w208 & ~w582;
assign w14021 = ~w341 & ~w432;
assign w14022 = ~w547 & w14021;
assign w14023 = w742 & w755;
assign w14024 = w1813 & w1854;
assign w14025 = w3117 & w14024;
assign w14026 = w14022 & w14023;
assign w14027 = w3287 & w4734;
assign w14028 = w14026 & w14027;
assign w14029 = w14025 & w14028;
assign w14030 = w1052 & w35170;
assign w14031 = ~w88 & w2249;
assign w14032 = w2861 & w14031;
assign w14033 = w14032 & w35171;
assign w14034 = ~w278 & ~w292;
assign w14035 = ~w540 & ~w559;
assign w14036 = w14034 & w14035;
assign w14037 = w2052 & w2150;
assign w14038 = w14020 & w14037;
assign w14039 = w1114 & w14036;
assign w14040 = w3769 & w5855;
assign w14041 = w14039 & w14040;
assign w14042 = w1763 & w14038;
assign w14043 = w4316 & w14042;
assign w14044 = w14041 & w14043;
assign w14045 = w377 & w14029;
assign w14046 = w14033 & w14045;
assign w14047 = w2901 & w14044;
assign w14048 = w14046 & w14047;
assign w14049 = ~w388 & ~w653;
assign w14050 = w1489 & w14049;
assign w14051 = w2559 & w3477;
assign w14052 = w14050 & w14051;
assign w14053 = w3346 & w14052;
assign w14054 = w3153 & w14053;
assign w14055 = ~w355 & ~w395;
assign w14056 = ~w719 & w2078;
assign w14057 = w4897 & w14055;
assign w14058 = w14056 & w14057;
assign w14059 = ~w89 & ~w159;
assign w14060 = ~w181 & ~w342;
assign w14061 = ~w559 & ~w568;
assign w14062 = w14060 & w14061;
assign w14063 = w1583 & w14059;
assign w14064 = w2154 & w2643;
assign w14065 = w2881 & w3237;
assign w14066 = w4298 & w5369;
assign w14067 = w14065 & w14066;
assign w14068 = w14063 & w14064;
assign w14069 = w14062 & w14068;
assign w14070 = w3307 & w14067;
assign w14071 = w14058 & w14070;
assign w14072 = w14069 & w14071;
assign w14073 = w14054 & w14072;
assign w14074 = w1097 & w2118;
assign w14075 = w14073 & w14074;
assign w14076 = ~w14048 & ~w14075;
assign w14077 = a_8 & ~w8276;
assign w14078 = ~a_5 & w8273;
assign w14079 = (~w14078 & w8276) | (~w14078 & w35172) | (w8276 & w35172);
assign w14080 = w14048 & w14075;
assign w14081 = ~w14076 & ~w14080;
assign w14082 = ~w14079 & w14081;
assign w14083 = (~w14076 & ~w14081) | (~w14076 & w35173) | (~w14081 & w35173);
assign w14084 = w13925 & ~w14083;
assign w14085 = ~w13925 & w14083;
assign w14086 = ~w14084 & ~w14085;
assign w14087 = w668 & w12856;
assign w14088 = w1327 & w12622;
assign w14089 = w1399 & ~w12630;
assign w14090 = (~w12842 & w35174) | (~w12842 & w35175) | (w35174 & w35175);
assign w14091 = ~w12854 & ~w14090;
assign w14092 = ~w14088 & ~w14089;
assign w14093 = ~w14087 & w14092;
assign w14094 = (w14093 & ~w14091) | (w14093 & w35176) | (~w14091 & w35176);
assign w14095 = w14086 & ~w14094;
assign w14096 = ~w13925 & w14018;
assign w14097 = ~w14019 & ~w14096;
assign w14098 = (~w14094 & w35178) | (~w14094 & w35179) | (w35178 & w35179);
assign w14099 = (w14094 & w35180) | (w14094 & w35181) | (w35180 & w35181);
assign w14100 = (~w13979 & w35182) | (~w13979 & w35183) | (w35182 & w35183);
assign w14101 = ~w13983 & w35184;
assign w14102 = ~w13983 & ~w14101;
assign w14103 = ~w13966 & w35185;
assign w14104 = ~w13968 & ~w14103;
assign w14105 = ~w14102 & w14104;
assign w14106 = w14102 & ~w14104;
assign w14107 = ~w14105 & ~w14106;
assign w14108 = ~w12905 & w35186;
assign w14109 = w3957 & ~w12878;
assign w14110 = ~w12892 & w35187;
assign w14111 = ~w13598 & w35188;
assign w14112 = ~w14109 & ~w14110;
assign w14113 = ~w14108 & w14112;
assign w14114 = ~w14111 & w35189;
assign w14115 = (a_29 & w14111) | (a_29 & w35190) | (w14111 & w35190);
assign w14116 = ~w14114 & ~w14115;
assign w14117 = w14107 & w14116;
assign w14118 = (~w14105 & ~w14107) | (~w14105 & w35191) | (~w14107 & w35191);
assign w14119 = w13973 & ~w14118;
assign w14120 = (~w13971 & w14118) | (~w13971 & w35192) | (w14118 & w35192);
assign w14121 = w13891 & ~w13900;
assign w14122 = ~w13901 & ~w14121;
assign w14123 = ~w14120 & w14122;
assign w14124 = ~w13901 & ~w14123;
assign w14125 = ~w13795 & ~w13804;
assign w14126 = ~w13805 & ~w14125;
assign w14127 = ~w14124 & w14126;
assign w14128 = w14124 & ~w14126;
assign w14129 = ~w14127 & ~w14128;
assign w14130 = ~w12589 & w35193;
assign w14131 = (~w518 & w12612) | (~w518 & w35194) | (w12612 & w35194);
assign w14132 = (w4638 & w12616) | (w4638 & w35195) | (w12616 & w35195);
assign w14133 = ~w14130 & ~w14131;
assign w14134 = ~w14132 & w14133;
assign w14135 = (w14134 & ~w13123) | (w14134 & w35196) | (~w13123 & w35196);
assign w14136 = a_26 & ~w14135;
assign w14137 = (~w13123 & w35197) | (~w13123 & w35198) | (w35197 & w35198);
assign w14138 = ~w14136 & ~w14137;
assign w14139 = w14129 & w14138;
assign w14140 = (~w14127 & ~w14129) | (~w14127 & w35199) | (~w14129 & w35199);
assign w14141 = ~w13836 & ~w13845;
assign w14142 = ~w13846 & ~w14141;
assign w14143 = ~w14140 & w14142;
assign w14144 = w14140 & ~w14142;
assign w14145 = ~w14143 & ~w14144;
assign w14146 = ~w13011 & w35200;
assign w14147 = w5016 & w12601;
assign w14148 = w5080 & w12598;
assign w14149 = ~w14147 & ~w14148;
assign w14150 = ~w14146 & w14149;
assign w14151 = (w14150 & w13021) | (w14150 & w35201) | (w13021 & w35201);
assign w14152 = ~a_23 & w14151;
assign w14153 = (~w13021 & w35202) | (~w13021 & w35203) | (w35202 & w35203);
assign w14154 = ~w14152 & ~w14153;
assign w14155 = w14145 & w14154;
assign w14156 = (~w14143 & ~w14145) | (~w14143 & w35204) | (~w14145 & w35204);
assign w14157 = ~w13880 & w13888;
assign w14158 = ~w13889 & ~w14157;
assign w14159 = ~w14156 & w14158;
assign w14160 = (~w13889 & ~w14158) | (~w13889 & w35205) | (~w14158 & w35205);
assign w14161 = (~w13875 & ~w13877) | (~w13875 & w35206) | (~w13877 & w35206);
assign w14162 = (~w13852 & ~w13853) | (~w13852 & w35207) | (~w13853 & w35207);
assign w14163 = ~w13615 & ~w13624;
assign w14164 = ~w13625 & ~w14163;
assign w14165 = w14162 & ~w14164;
assign w14166 = ~w14162 & w14164;
assign w14167 = ~w14165 & ~w14166;
assign w14168 = w4666 & w12598;
assign w14169 = ~w518 & w12604;
assign w14170 = w4638 & w12601;
assign w14171 = ~w14169 & ~w14170;
assign w14172 = ~w14168 & w14171;
assign w14173 = (w14172 & ~w12961) | (w14172 & w35208) | (~w12961 & w35208);
assign w14174 = ~a_26 & w14173;
assign w14175 = (w12961 & w35209) | (w12961 & w35210) | (w35209 & w35210);
assign w14176 = ~w14174 & ~w14175;
assign w14177 = w14167 & w14176;
assign w14178 = ~w14167 & ~w14176;
assign w14179 = ~w14177 & ~w14178;
assign w14180 = ~w14161 & w14179;
assign w14181 = w14161 & ~w14179;
assign w14182 = ~w14180 & ~w14181;
assign w14183 = w5286 & w13177;
assign w14184 = ~w13011 & w35211;
assign w14185 = ~w13174 & w35212;
assign w14186 = ~w14184 & ~w14185;
assign w14187 = ~w14183 & w14186;
assign w14188 = (w14187 & ~w13207) | (w14187 & w35213) | (~w13207 & w35213);
assign w14189 = ~a_23 & w14188;
assign w14190 = (w13207 & w35214) | (w13207 & w35215) | (w35214 & w35215);
assign w14191 = ~w14189 & ~w14190;
assign w14192 = w14182 & w14191;
assign w14193 = ~w14182 & ~w14191;
assign w14194 = ~w14192 & ~w14193;
assign w14195 = ~w14160 & w14194;
assign w14196 = w14160 & ~w14194;
assign w14197 = ~w14195 & ~w14196;
assign w14198 = (~w13173 & w35218) | (~w13173 & w35219) | (w35218 & w35219);
assign w14199 = (~w13173 & w35220) | (~w13173 & w35221) | (w35220 & w35221);
assign w14200 = ~w14198 & w14199;
assign w14201 = ~w13109 & ~w14200;
assign w14202 = w14197 & w14201;
assign w14203 = (~w14195 & ~w14197) | (~w14195 & w35222) | (~w14197 & w35222);
assign w14204 = (~w14180 & ~w14182) | (~w14180 & w35223) | (~w14182 & w35223);
assign w14205 = w13111 & ~w14204;
assign w14206 = ~w13111 & w14204;
assign w14207 = ~w14205 & ~w14206;
assign w14208 = (~w14166 & ~w14167) | (~w14166 & w35224) | (~w14167 & w35224);
assign w14209 = ~w13696 & ~w13705;
assign w14210 = ~w13706 & ~w14209;
assign w14211 = w14208 & ~w14210;
assign w14212 = ~w14208 & w14210;
assign w14213 = ~w14211 & ~w14212;
assign w14214 = w5080 & w13177;
assign w14215 = ~w13174 & w35225;
assign w14216 = (w13173 & w35226) | (w13173 & w35227) | (w35226 & w35227);
assign w14217 = ~w14215 & ~w14216;
assign w14218 = ~w14214 & w14217;
assign w14219 = (w14218 & w13264) | (w14218 & w35228) | (w13264 & w35228);
assign w14220 = ~a_23 & w14219;
assign w14221 = (~w13264 & w35229) | (~w13264 & w35230) | (w35229 & w35230);
assign w14222 = ~w14220 & ~w14221;
assign w14223 = w14213 & w14222;
assign w14224 = ~w14213 & ~w14222;
assign w14225 = ~w14223 & ~w14224;
assign w14226 = w14207 & w14225;
assign w14227 = ~w14207 & ~w14225;
assign w14228 = ~w14226 & ~w14227;
assign w14229 = w14203 & ~w14228;
assign w14230 = w14120 & ~w14122;
assign w14231 = ~w14123 & ~w14230;
assign w14232 = (w4666 & w12616) | (w4666 & w35231) | (w12616 & w35231);
assign w14233 = ~w12930 & w35232;
assign w14234 = (w4638 & w12612) | (w4638 & w35233) | (w12612 & w35233);
assign w14235 = ~w14233 & ~w14234;
assign w14236 = ~w14232 & w14235;
assign w14237 = (w14236 & ~w13389) | (w14236 & w35234) | (~w13389 & w35234);
assign w14238 = a_26 & ~w14237;
assign w14239 = (~w13389 & w35235) | (~w13389 & w35236) | (w35235 & w35236);
assign w14240 = ~w14238 & ~w14239;
assign w14241 = w14231 & w14240;
assign w14242 = ~w13973 & w14118;
assign w14243 = ~w14119 & ~w14242;
assign w14244 = ~w12905 & w35237;
assign w14245 = w4446 & ~w12910;
assign w14246 = ~w12892 & w35238;
assign w14247 = w4070 & w13815;
assign w14248 = ~w14245 & w35239;
assign w14249 = ~w14247 & w35240;
assign w14250 = (a_29 & w14247) | (a_29 & w35241) | (w14247 & w35241);
assign w14251 = ~w14249 & ~w14250;
assign w14252 = w14243 & w14251;
assign w14253 = ~w14243 & ~w14251;
assign w14254 = ~w14252 & ~w14253;
assign w14255 = (w4666 & w12612) | (w4666 & w35242) | (w12612 & w35242);
assign w14256 = ~w12914 & w35243;
assign w14257 = ~w12930 & w35244;
assign w14258 = ~w14256 & ~w14257;
assign w14259 = ~w14255 & w14258;
assign w14260 = (w14259 & ~w13375) | (w14259 & w35245) | (~w13375 & w35245);
assign w14261 = a_26 & ~w14260;
assign w14262 = (~w13375 & w35246) | (~w13375 & w35247) | (w35246 & w35247);
assign w14263 = ~w14261 & ~w14262;
assign w14264 = w14254 & w14263;
assign w14265 = (~w14252 & ~w14254) | (~w14252 & w35248) | (~w14254 & w35248);
assign w14266 = ~w14231 & ~w14240;
assign w14267 = ~w14241 & ~w14266;
assign w14268 = ~w14265 & w14267;
assign w14269 = ~w14241 & ~w14268;
assign w14270 = ~w14129 & ~w14138;
assign w14271 = ~w14139 & ~w14270;
assign w14272 = ~w14269 & w14271;
assign w14273 = w14269 & ~w14271;
assign w14274 = ~w14272 & ~w14273;
assign w14275 = w5286 & w12598;
assign w14276 = w5016 & w12604;
assign w14277 = w5080 & w12601;
assign w14278 = ~w14276 & ~w14277;
assign w14279 = ~w14275 & w14278;
assign w14280 = (w14279 & ~w12961) | (w14279 & w35249) | (~w12961 & w35249);
assign w14281 = ~a_23 & w14280;
assign w14282 = (w12961 & w35250) | (w12961 & w35251) | (w35250 & w35251);
assign w14283 = ~w14281 & ~w14282;
assign w14284 = w14274 & w14283;
assign w14285 = (~w14272 & ~w14274) | (~w14272 & w35252) | (~w14274 & w35252);
assign w14286 = ~w14145 & ~w14154;
assign w14287 = ~w14155 & ~w14286;
assign w14288 = ~w14285 & w14287;
assign w14289 = w14285 & ~w14287;
assign w14290 = ~w14288 & ~w14289;
assign w14291 = w5818 & w13177;
assign w14292 = ~w13174 & w35253;
assign w14293 = (w13173 & w35254) | (w13173 & w35255) | (w35254 & w35255);
assign w14294 = ~w14292 & ~w14293;
assign w14295 = ~w14291 & w14294;
assign w14296 = (w14295 & w13264) | (w14295 & w35256) | (w13264 & w35256);
assign w14297 = a_20 & ~w14296;
assign w14298 = (w13264 & w35257) | (w13264 & w35258) | (w35257 & w35258);
assign w14299 = ~w14297 & ~w14298;
assign w14300 = w14290 & w14299;
assign w14301 = (~w14288 & ~w14290) | (~w14288 & w35259) | (~w14290 & w35259);
assign w14302 = w5308 & w13177;
assign w14303 = (w13201 & w35262) | (w13201 & w35263) | (w35262 & w35263);
assign w14304 = (~w13173 & w35264) | (~w13173 & w35265) | (w35264 & w35265);
assign w14305 = ~w14302 & w14304;
assign w14306 = (a_20 & w14303) | (a_20 & w35266) | (w14303 & w35266);
assign w14307 = ~w14303 & w35267;
assign w14308 = ~w14306 & ~w14307;
assign w14309 = ~w14301 & w14308;
assign w14310 = w14156 & ~w14158;
assign w14311 = ~w14159 & ~w14310;
assign w14312 = w14301 & ~w14308;
assign w14313 = ~w14309 & ~w14312;
assign w14314 = w14311 & w14313;
assign w14315 = (~w14309 & ~w14313) | (~w14309 & w35268) | (~w14313 & w35268);
assign w14316 = ~w14197 & ~w14201;
assign w14317 = ~w14202 & ~w14316;
assign w14318 = ~w14315 & w14317;
assign w14319 = ~w14203 & w14228;
assign w14320 = ~w14229 & ~w14319;
assign w14321 = ~w14318 & w14320;
assign w14322 = (~w14229 & w14318) | (~w14229 & w35269) | (w14318 & w35269);
assign w14323 = ~w429 & w2008;
assign w14324 = w2008 & w35270;
assign w14325 = ~w547 & w1124;
assign w14326 = w1644 & w2942;
assign w14327 = w3893 & w4913;
assign w14328 = w13911 & w14327;
assign w14329 = w14325 & w14326;
assign w14330 = w5545 & w12968;
assign w14331 = w14329 & w14330;
assign w14332 = w1531 & w14328;
assign w14333 = w14324 & w14332;
assign w14334 = w1549 & w14331;
assign w14335 = w14333 & w14334;
assign w14336 = w3233 & w14335;
assign w14337 = w3453 & w14336;
assign w14338 = w14048 & ~w14337;
assign w14339 = ~a_2 & ~w10839;
assign w14340 = ~w136 & ~w166;
assign w14341 = ~w220 & w14340;
assign w14342 = w280 & w947;
assign w14343 = w1018 & w1100;
assign w14344 = w2100 & w2400;
assign w14345 = w2742 & w14344;
assign w14346 = w14342 & w14343;
assign w14347 = w14341 & w14346;
assign w14348 = w1566 & w14345;
assign w14349 = w14347 & w14348;
assign w14350 = ~w248 & ~w1123;
assign w14351 = w5367 & w14350;
assign w14352 = w1109 & w2417;
assign w14353 = w14351 & w14352;
assign w14354 = w779 & w1679;
assign w14355 = w2151 & w3419;
assign w14356 = w14354 & w14355;
assign w14357 = w2926 & w4354;
assign w14358 = w13562 & w14357;
assign w14359 = w3991 & w14356;
assign w14360 = w14353 & w14359;
assign w14361 = w2614 & w14358;
assign w14362 = w14360 & w14361;
assign w14363 = w14349 & w14362;
assign w14364 = ~w255 & ~w287;
assign w14365 = w938 & w14364;
assign w14366 = w1631 & w1639;
assign w14367 = w2603 & w4094;
assign w14368 = w14366 & w14367;
assign w14369 = w4344 & w14365;
assign w14370 = w14368 & w14369;
assign w14371 = w6171 & w6577;
assign w14372 = w14370 & w14371;
assign w14373 = w4195 & w14372;
assign w14374 = w13910 & w14373;
assign w14375 = w14363 & w14374;
assign w14376 = ~w14339 & ~w14375;
assign w14377 = a_5 & ~w9785;
assign w14378 = ~a_4 & w9774;
assign w14379 = (~w14378 & w9785) | (~w14378 & w35271) | (w9785 & w35271);
assign w14380 = w14339 & w14375;
assign w14381 = ~w14376 & ~w14380;
assign w14382 = ~w14379 & w14381;
assign w14383 = (~w14376 & ~w14381) | (~w14376 & w35272) | (~w14381 & w35272);
assign w14384 = w14048 & ~w14383;
assign w14385 = ~w14048 & w14383;
assign w14386 = ~w14384 & ~w14385;
assign w14387 = w668 & ~w12668;
assign w14388 = w1327 & ~w12661;
assign w14389 = w1399 & ~w12637;
assign w14390 = (~w12670 & w12659) | (~w12670 & w35273) | (w12659 & w35273);
assign w14391 = ~w12838 & w31783;
assign w14392 = (~w12673 & w12838) | (~w12673 & w35274) | (w12838 & w35274);
assign w14393 = ~w14391 & ~w14392;
assign w14394 = ~w14388 & ~w14389;
assign w14395 = ~w14387 & w14394;
assign w14396 = (w14395 & ~w14393) | (w14395 & w35275) | (~w14393 & w35275);
assign w14397 = w14386 & ~w14396;
assign w14398 = ~w14048 & w14337;
assign w14399 = ~w14338 & ~w14398;
assign w14400 = (~w14396 & w35277) | (~w14396 & w35278) | (w35277 & w35278);
assign w14401 = w14079 & ~w14081;
assign w14402 = ~w14082 & ~w14401;
assign w14403 = (~w14396 & w35281) | (~w14396 & w35282) | (w35281 & w35282);
assign w14404 = (w14396 & w35283) | (w14396 & w35284) | (w35283 & w35284);
assign w14405 = ~w14403 & ~w14404;
assign w14406 = w1327 & ~w12630;
assign w14407 = w1399 & ~w12668;
assign w14408 = w668 & w12622;
assign w14409 = ~w12631 & ~w12843;
assign w14410 = ~w12842 & w35285;
assign w14411 = (~w14409 & w12842) | (~w14409 & w35286) | (w12842 & w35286);
assign w14412 = ~w14410 & ~w14411;
assign w14413 = ~w14406 & ~w14407;
assign w14414 = ~w14408 & w14413;
assign w14415 = (w14414 & w14412) | (w14414 & w35287) | (w14412 & w35287);
assign w14416 = w14405 & ~w14415;
assign w14417 = (~w14403 & ~w14405) | (~w14403 & w35288) | (~w14405 & w35288);
assign w14418 = (~w14091 & w35289) | (~w14091 & w35290) | (w35289 & w35290);
assign w14419 = ~w14095 & ~w14418;
assign w14420 = ~w14417 & w14419;
assign w14421 = w14417 & ~w14419;
assign w14422 = ~w14420 & ~w14421;
assign w14423 = w4446 & w12874;
assign w14424 = w3957 & ~w12860;
assign w14425 = w4068 & w12869;
assign w14426 = w4070 & w13965;
assign w14427 = ~w14424 & w35291;
assign w14428 = ~w14426 & w35292;
assign w14429 = (a_29 & w14426) | (a_29 & w35293) | (w14426 & w35293);
assign w14430 = ~w14428 & ~w14429;
assign w14431 = w14422 & w14430;
assign w14432 = (~w14420 & ~w14422) | (~w14420 & w35294) | (~w14422 & w35294);
assign w14433 = (w14094 & w35295) | (w14094 & w35296) | (w35295 & w35296);
assign w14434 = ~w14098 & ~w14433;
assign w14435 = w668 & ~w12860;
assign w14436 = w1327 & w12856;
assign w14437 = w1399 & w12622;
assign w14438 = (~w12842 & w35297) | (~w12842 & w35298) | (w35297 & w35298);
assign w14439 = ~w12861 & ~w12864;
assign w14440 = w14438 & ~w14439;
assign w14441 = ~w14438 & w14439;
assign w14442 = ~w14440 & ~w14441;
assign w14443 = ~w14436 & ~w14437;
assign w14444 = ~w14435 & w14443;
assign w14445 = (w14444 & ~w14442) | (w14444 & w35299) | (~w14442 & w35299);
assign w14446 = w14434 & ~w14445;
assign w14447 = ~w14434 & w14445;
assign w14448 = ~w14446 & ~w14447;
assign w14449 = w4446 & ~w12878;
assign w14450 = w4068 & w12874;
assign w14451 = w3957 & w12869;
assign w14452 = ~w14450 & ~w14451;
assign w14453 = ~w14449 & w14452;
assign w14454 = (w14453 & ~w13771) | (w14453 & w35300) | (~w13771 & w35300);
assign w14455 = a_29 & ~w14454;
assign w14456 = (~w13771 & w35301) | (~w13771 & w35302) | (w35301 & w35302);
assign w14457 = ~w14455 & ~w14456;
assign w14458 = w14448 & w14457;
assign w14459 = ~w14448 & ~w14457;
assign w14460 = ~w14458 & ~w14459;
assign w14461 = ~w14432 & w14460;
assign w14462 = w14432 & ~w14460;
assign w14463 = ~w14461 & ~w14462;
assign w14464 = ~w12905 & w35303;
assign w14465 = w4666 & ~w12910;
assign w14466 = ~w12892 & w35304;
assign w14467 = w1226 & w13815;
assign w14468 = ~w14465 & w35305;
assign w14469 = ~w14467 & w35306;
assign w14470 = (a_26 & w14467) | (a_26 & w35307) | (w14467 & w35307);
assign w14471 = ~w14469 & ~w14470;
assign w14472 = w14463 & w14471;
assign w14473 = (~w14461 & ~w14463) | (~w14461 & w35308) | (~w14463 & w35308);
assign w14474 = (w14099 & w13983) | (w14099 & w35309) | (w13983 & w35309);
assign w14475 = ~w14101 & ~w14474;
assign w14476 = (w14475 & w14458) | (w14475 & w35310) | (w14458 & w35310);
assign w14477 = ~w14458 & w35311;
assign w14478 = ~w14476 & ~w14477;
assign w14479 = ~w12892 & w35312;
assign w14480 = w4068 & ~w12878;
assign w14481 = w3957 & w12874;
assign w14482 = ~w14480 & ~w14481;
assign w14483 = ~w14479 & w14482;
assign w14484 = (w14483 & ~w13787) | (w14483 & w35313) | (~w13787 & w35313);
assign w14485 = ~a_29 & w14484;
assign w14486 = (w13787 & w35314) | (w13787 & w35315) | (w35314 & w35315);
assign w14487 = ~w14485 & ~w14486;
assign w14488 = w14478 & w14487;
assign w14489 = ~w14478 & ~w14487;
assign w14490 = ~w14488 & ~w14489;
assign w14491 = ~w12914 & w35316;
assign w14492 = w4638 & ~w12910;
assign w14493 = ~w12905 & w35317;
assign w14494 = (w1226 & w13518) | (w1226 & w35318) | (w13518 & w35318);
assign w14495 = ~w14492 & ~w14493;
assign w14496 = ~w14491 & w14495;
assign w14497 = ~w14494 & w35319;
assign w14498 = (a_26 & w14494) | (a_26 & w35320) | (w14494 & w35320);
assign w14499 = ~w14497 & ~w14498;
assign w14500 = w14490 & w14499;
assign w14501 = ~w14490 & ~w14499;
assign w14502 = ~w14500 & ~w14501;
assign w14503 = ~w14473 & w14502;
assign w14504 = w14473 & ~w14502;
assign w14505 = ~w14503 & ~w14504;
assign w14506 = (w5286 & w12616) | (w5286 & w35321) | (w12616 & w35321);
assign w14507 = (w5080 & w12612) | (w5080 & w35322) | (w12612 & w35322);
assign w14508 = ~w12930 & w35323;
assign w14509 = ~w14507 & ~w14508;
assign w14510 = ~w14506 & w14509;
assign w14511 = (w14510 & ~w13389) | (w14510 & w35324) | (~w13389 & w35324);
assign w14512 = a_23 & ~w14511;
assign w14513 = (~w13389 & w35325) | (~w13389 & w35326) | (w35325 & w35326);
assign w14514 = ~w14512 & ~w14513;
assign w14515 = w14505 & w14514;
assign w14516 = ~w14405 & w14415;
assign w14517 = ~w14416 & ~w14516;
assign w14518 = w3957 & w12856;
assign w14519 = w4446 & w12869;
assign w14520 = (~w14518 & w12860) | (~w14518 & w35327) | (w12860 & w35327);
assign w14521 = ~w14519 & w14520;
assign w14522 = (w14521 & ~w13979) | (w14521 & w35328) | (~w13979 & w35328);
assign w14523 = a_29 & ~w14522;
assign w14524 = (~w13979 & w35329) | (~w13979 & w35330) | (w35329 & w35330);
assign w14525 = ~w14523 & ~w14524;
assign w14526 = w14517 & w14525;
assign w14527 = (w14396 & w35331) | (w14396 & w35332) | (w35331 & w35332);
assign w14528 = ~w14400 & ~w14527;
assign w14529 = w668 & ~w12630;
assign w14530 = w1399 & ~w12661;
assign w14531 = w1327 & ~w12668;
assign w14532 = ~w12669 & ~w12845;
assign w14533 = (~w14532 & w14391) | (~w14532 & w35333) | (w14391 & w35333);
assign w14534 = ~w14391 & w35334;
assign w14535 = ~w14533 & ~w14534;
assign w14536 = ~w14530 & ~w14531;
assign w14537 = ~w14529 & w14536;
assign w14538 = (w14537 & w14535) | (w14537 & w35335) | (w14535 & w35335);
assign w14539 = w14528 & ~w14538;
assign w14540 = ~w14528 & w14538;
assign w14541 = ~w14539 & ~w14540;
assign w14542 = (~w14393 & w35336) | (~w14393 & w35337) | (w35336 & w35337);
assign w14543 = ~w14397 & ~w14542;
assign w14544 = ~w76 & ~w85;
assign w14545 = ~w896 & w14544;
assign w14546 = w2619 & w3079;
assign w14547 = w3305 & w3516;
assign w14548 = w4368 & w14547;
assign w14549 = w14545 & w14546;
assign w14550 = w2053 & w14549;
assign w14551 = w873 & w14548;
assign w14552 = w2574 & w14551;
assign w14553 = w1024 & w14550;
assign w14554 = w14552 & w14553;
assign w14555 = w1434 & w14554;
assign w14556 = w4126 & w14555;
assign w14557 = w14339 & ~w14556;
assign w14558 = ~w14339 & w14556;
assign w14559 = ~w14557 & ~w14558;
assign w14560 = w1309 & w2743;
assign w14561 = w387 & w6692;
assign w14562 = ~w53 & w2990;
assign w14563 = w3282 & w4714;
assign w14564 = w13060 & w14563;
assign w14565 = w1302 & w14562;
assign w14566 = w2554 & w3236;
assign w14567 = w14560 & w14566;
assign w14568 = w14564 & w14565;
assign w14569 = w13035 & w14561;
assign w14570 = w14568 & w14569;
assign w14571 = w903 & w14567;
assign w14572 = w1859 & w14571;
assign w14573 = w14570 & w14572;
assign w14574 = w14363 & w14573;
assign w14575 = ~w14339 & w14574;
assign w14576 = ~w134 & ~w214;
assign w14577 = w595 & w6696;
assign w14578 = w4926 & w14577;
assign w14579 = ~w10 & w2988;
assign w14580 = ~w113 & w3211;
assign w14581 = w4902 & w14580;
assign w14582 = w14579 & w14581;
assign w14583 = ~w582 & ~w652;
assign w14584 = w1153 & w14583;
assign w14585 = w2681 & w2796;
assign w14586 = w3122 & w3740;
assign w14587 = w4089 & w14586;
assign w14588 = w14584 & w14585;
assign w14589 = w915 & w4198;
assign w14590 = w14588 & w14589;
assign w14591 = w3390 & w14587;
assign w14592 = w14590 & w14591;
assign w14593 = w14582 & w14592;
assign w14594 = ~w152 & ~w287;
assign w14595 = w2252 & w14594;
assign w14596 = w3343 & w14595;
assign w14597 = w14592 & w35338;
assign w14598 = ~w585 & ~w720;
assign w14599 = w467 & w879;
assign w14600 = w1009 & w2555;
assign w14601 = w14576 & w14598;
assign w14602 = w14600 & w14601;
assign w14603 = w943 & w14599;
assign w14604 = w3118 & w13984;
assign w14605 = w14603 & w14604;
assign w14606 = w3368 & w14602;
assign w14607 = w14605 & w14606;
assign w14608 = w14578 & w14607;
assign w14609 = w13347 & w14608;
assign w14610 = w14609 & w35339;
assign w14611 = (w14339 & ~w14609) | (w14339 & w35340) | (~w14609 & w35340);
assign w14612 = ~w14610 & ~w14611;
assign w14613 = ~w12828 & ~w12833;
assign w14614 = ~w12834 & ~w14613;
assign w14615 = w668 & w12651;
assign w14616 = w1399 & w12793;
assign w14617 = w1327 & ~w12830;
assign w14618 = ~w14615 & ~w14616;
assign w14619 = ~w14617 & w14618;
assign w14620 = (~w14614 & w35341) | (~w14614 & w35342) | (w35341 & w35342);
assign w14621 = (w14614 & w35343) | (w14614 & w35344) | (w35343 & w35344);
assign w14622 = w14339 & ~w14574;
assign w14623 = ~w14575 & ~w14622;
assign w14624 = ~w14621 & w14623;
assign w14625 = (w14621 & w35346) | (w14621 & w35347) | (w35346 & w35347);
assign w14626 = w14379 & ~w14381;
assign w14627 = ~w14382 & ~w14626;
assign w14628 = (w14621 & w35350) | (w14621 & w35351) | (w35350 & w35351);
assign w14629 = (~w14621 & w35352) | (~w14621 & w35353) | (w35352 & w35353);
assign w14630 = w668 & ~w12661;
assign w14631 = w1327 & ~w12637;
assign w14632 = w1399 & w12646;
assign w14633 = (w12836 & ~w12828) | (w12836 & w31785) | (~w12828 & w31785);
assign w14634 = ~w12662 & ~w12670;
assign w14635 = (~w12648 & ~w12649) | (~w12648 & w32454) | (~w12649 & w32454);
assign w14636 = ~w14634 & ~w14635;
assign w14637 = ~w14633 & w14636;
assign w14638 = w12836 & w14634;
assign w14639 = w14634 & w14635;
assign w14640 = (~w14639 & w12834) | (~w14639 & w35354) | (w12834 & w35354);
assign w14641 = ~w14637 & w14640;
assign w14642 = ~w14631 & ~w14632;
assign w14643 = ~w14630 & w14642;
assign w14644 = (w14643 & w14641) | (w14643 & w35355) | (w14641 & w35355);
assign w14645 = ~w14629 & ~w14644;
assign w14646 = ~w14628 & ~w14645;
assign w14647 = w14543 & ~w14646;
assign w14648 = ~w14543 & w14646;
assign w14649 = w4446 & w12856;
assign w14650 = w4068 & w12622;
assign w14651 = w3957 & ~w12630;
assign w14652 = ~w14650 & ~w14651;
assign w14653 = ~w14649 & w14652;
assign w14654 = (w14653 & ~w14091) | (w14653 & w35356) | (~w14091 & w35356);
assign w14655 = ~a_29 & w14654;
assign w14656 = (w14091 & w35357) | (w14091 & w35358) | (w35357 & w35358);
assign w14657 = ~w14655 & ~w14656;
assign w14658 = ~w14648 & w14657;
assign w14659 = ~w14647 & ~w14658;
assign w14660 = w14541 & ~w14659;
assign w14661 = (~w14539 & w14659) | (~w14539 & w35359) | (w14659 & w35359);
assign w14662 = ~w14517 & ~w14525;
assign w14663 = ~w14526 & ~w14662;
assign w14664 = ~w14661 & w14663;
assign w14665 = ~w14526 & ~w14664;
assign w14666 = ~w14422 & ~w14430;
assign w14667 = ~w14431 & ~w14666;
assign w14668 = ~w14665 & w14667;
assign w14669 = w14665 & ~w14667;
assign w14670 = ~w14668 & ~w14669;
assign w14671 = ~w12905 & w35360;
assign w14672 = ~w518 & ~w12878;
assign w14673 = ~w12892 & w35361;
assign w14674 = ~w13598 & w35362;
assign w14675 = ~w14672 & ~w14673;
assign w14676 = ~w14671 & w14675;
assign w14677 = ~w14674 & w35363;
assign w14678 = (a_26 & w14674) | (a_26 & w35364) | (w14674 & w35364);
assign w14679 = ~w14677 & ~w14678;
assign w14680 = w14670 & w14679;
assign w14681 = (~w14668 & ~w14670) | (~w14668 & w35365) | (~w14670 & w35365);
assign w14682 = ~w14463 & ~w14471;
assign w14683 = ~w14472 & ~w14682;
assign w14684 = ~w14681 & w14683;
assign w14685 = w14681 & ~w14683;
assign w14686 = ~w14684 & ~w14685;
assign w14687 = (w5286 & w12612) | (w5286 & w35366) | (w12612 & w35366);
assign w14688 = ~w12914 & w35367;
assign w14689 = ~w12930 & w35368;
assign w14690 = ~w14688 & ~w14689;
assign w14691 = ~w14687 & w14690;
assign w14692 = (w14691 & ~w13375) | (w14691 & w35369) | (~w13375 & w35369);
assign w14693 = a_23 & w14692;
assign w14694 = (w13375 & w35370) | (w13375 & w35371) | (w35370 & w35371);
assign w14695 = ~w14693 & ~w14694;
assign w14696 = w14686 & ~w14695;
assign w14697 = (~w14684 & ~w14686) | (~w14684 & w35372) | (~w14686 & w35372);
assign w14698 = ~w14505 & ~w14514;
assign w14699 = ~w14515 & ~w14698;
assign w14700 = ~w14697 & w14699;
assign w14701 = (~w14515 & ~w14699) | (~w14515 & w35373) | (~w14699 & w35373);
assign w14702 = (~w14500 & ~w14502) | (~w14500 & w35374) | (~w14502 & w35374);
assign w14703 = (~w14476 & ~w14478) | (~w14476 & w35375) | (~w14478 & w35375);
assign w14704 = ~w14107 & ~w14116;
assign w14705 = ~w14117 & ~w14704;
assign w14706 = ~w14703 & w14705;
assign w14707 = w14703 & ~w14705;
assign w14708 = ~w14706 & ~w14707;
assign w14709 = ~w12930 & w35376;
assign w14710 = ~w12914 & w35377;
assign w14711 = ~w518 & ~w12910;
assign w14712 = ~w13501 & w35378;
assign w14713 = ~w14710 & ~w14711;
assign w14714 = ~w14709 & w14713;
assign w14715 = (a_26 & w14712) | (a_26 & w35379) | (w14712 & w35379);
assign w14716 = ~w14712 & w35380;
assign w14717 = ~w14715 & ~w14716;
assign w14718 = w14708 & w14717;
assign w14719 = ~w14708 & ~w14717;
assign w14720 = ~w14718 & ~w14719;
assign w14721 = w14702 & ~w14720;
assign w14722 = ~w14702 & w14720;
assign w14723 = ~w14721 & ~w14722;
assign w14724 = (w5080 & w12616) | (w5080 & w35381) | (w12616 & w35381);
assign w14725 = (w5016 & w12612) | (w5016 & w35382) | (w12612 & w35382);
assign w14726 = ~w12589 & w35383;
assign w14727 = ~w14724 & ~w14725;
assign w14728 = ~w14726 & w14727;
assign w14729 = (w14728 & ~w13123) | (w14728 & w35384) | (~w13123 & w35384);
assign w14730 = ~a_23 & w14729;
assign w14731 = (w13123 & w35385) | (w13123 & w35386) | (w35385 & w35386);
assign w14732 = ~w14730 & ~w14731;
assign w14733 = w14723 & w14732;
assign w14734 = ~w14723 & ~w14732;
assign w14735 = ~w14733 & ~w14734;
assign w14736 = ~w14701 & w14735;
assign w14737 = w14701 & ~w14735;
assign w14738 = ~w14736 & ~w14737;
assign w14739 = w5816 & w12598;
assign w14740 = w5818 & w12601;
assign w14741 = w5308 & w12604;
assign w14742 = ~w14740 & ~w14741;
assign w14743 = ~w14739 & w14742;
assign w14744 = (w14743 & ~w12961) | (w14743 & w35387) | (~w12961 & w35387);
assign w14745 = a_20 & ~w14744;
assign w14746 = (~w12961 & w35388) | (~w12961 & w35389) | (w35388 & w35389);
assign w14747 = ~w14745 & ~w14746;
assign w14748 = w14738 & w14747;
assign w14749 = (~w14736 & ~w14738) | (~w14736 & w35390) | (~w14738 & w35390);
assign w14750 = (~w14722 & ~w14723) | (~w14722 & w35391) | (~w14723 & w35391);
assign w14751 = (~w14706 & ~w14708) | (~w14706 & w35392) | (~w14708 & w35392);
assign w14752 = ~w14254 & ~w14263;
assign w14753 = ~w14264 & ~w14752;
assign w14754 = ~w14751 & w14753;
assign w14755 = w14751 & ~w14753;
assign w14756 = ~w14754 & ~w14755;
assign w14757 = w5286 & w12604;
assign w14758 = (w5016 & w12616) | (w5016 & w35393) | (w12616 & w35393);
assign w14759 = ~w12589 & w35394;
assign w14760 = ~w14758 & ~w14759;
assign w14761 = ~w14757 & w14760;
assign w14762 = (w14761 & w13288) | (w14761 & w35395) | (w13288 & w35395);
assign w14763 = ~a_23 & w14762;
assign w14764 = (~w13288 & w35396) | (~w13288 & w35397) | (w35396 & w35397);
assign w14765 = ~w14763 & ~w14764;
assign w14766 = w14756 & w14765;
assign w14767 = ~w14756 & ~w14765;
assign w14768 = ~w14766 & ~w14767;
assign w14769 = w14750 & ~w14768;
assign w14770 = ~w14750 & w14768;
assign w14771 = ~w14769 & ~w14770;
assign w14772 = ~w13011 & w35398;
assign w14773 = w5818 & w12598;
assign w14774 = w5308 & w12601;
assign w14775 = ~w14773 & ~w14774;
assign w14776 = ~w14772 & w14775;
assign w14777 = (w14776 & w13021) | (w14776 & w35399) | (w13021 & w35399);
assign w14778 = ~a_20 & w14777;
assign w14779 = (~w13021 & w35400) | (~w13021 & w35401) | (w35400 & w35401);
assign w14780 = ~w14778 & ~w14779;
assign w14781 = w14771 & w14780;
assign w14782 = ~w14771 & ~w14780;
assign w14783 = ~w14781 & ~w14782;
assign w14784 = ~w14749 & w14783;
assign w14785 = w14749 & ~w14783;
assign w14786 = ~w14784 & ~w14785;
assign w14787 = w6061 & w13177;
assign w14788 = ~w13174 & w35402;
assign w14789 = (w13173 & w35403) | (w13173 & w35404) | (w35403 & w35404);
assign w14790 = ~w14788 & ~w14789;
assign w14791 = ~w14787 & w14790;
assign w14792 = (w14791 & w13264) | (w14791 & w35405) | (w13264 & w35405);
assign w14793 = ~a_17 & w14792;
assign w14794 = (~w13264 & w35406) | (~w13264 & w35407) | (w35406 & w35407);
assign w14795 = ~w14793 & ~w14794;
assign w14796 = w14786 & w14795;
assign w14797 = (~w14784 & ~w14786) | (~w14784 & w35408) | (~w14786 & w35408);
assign w14798 = w6059 & w13177;
assign w14799 = (w13201 & w35411) | (w13201 & w35412) | (w35411 & w35412);
assign w14800 = (~w13173 & w35413) | (~w13173 & w35414) | (w35413 & w35414);
assign w14801 = ~w14798 & w14800;
assign w14802 = (a_17 & w14799) | (a_17 & w35415) | (w14799 & w35415);
assign w14803 = ~w14799 & w35416;
assign w14804 = ~w14802 & ~w14803;
assign w14805 = ~w14797 & w14804;
assign w14806 = (~w14770 & ~w14771) | (~w14770 & w35417) | (~w14771 & w35417);
assign w14807 = (~w14754 & ~w14756) | (~w14754 & w35418) | (~w14756 & w35418);
assign w14808 = w14265 & ~w14267;
assign w14809 = ~w14268 & ~w14808;
assign w14810 = w5286 & w12601;
assign w14811 = ~w12589 & w35419;
assign w14812 = w5080 & w12604;
assign w14813 = ~w14811 & ~w14812;
assign w14814 = ~w14810 & w14813;
assign w14815 = (w14814 & w13140) | (w14814 & w35420) | (w13140 & w35420);
assign w14816 = a_23 & w14815;
assign w14817 = (~w13140 & w35421) | (~w13140 & w35422) | (w35421 & w35422);
assign w14818 = ~w14816 & ~w14817;
assign w14819 = w14809 & ~w14818;
assign w14820 = ~w14809 & w14818;
assign w14821 = ~w14819 & ~w14820;
assign w14822 = ~w14807 & w14821;
assign w14823 = w14807 & ~w14821;
assign w14824 = ~w14822 & ~w14823;
assign w14825 = ~w13174 & w35423;
assign w14826 = ~w13011 & w35424;
assign w14827 = w5308 & w12598;
assign w14828 = ~w13205 & w35425;
assign w14829 = ~w14826 & w35426;
assign w14830 = (a_20 & w14828) | (a_20 & w35427) | (w14828 & w35427);
assign w14831 = ~w14828 & w35428;
assign w14832 = ~w14830 & ~w14831;
assign w14833 = w14824 & w14832;
assign w14834 = ~w14824 & ~w14832;
assign w14835 = ~w14833 & ~w14834;
assign w14836 = ~w14806 & w14835;
assign w14837 = w14806 & ~w14835;
assign w14838 = ~w14836 & ~w14837;
assign w14839 = w14797 & ~w14804;
assign w14840 = ~w14805 & ~w14839;
assign w14841 = w14838 & w14840;
assign w14842 = (~w14805 & ~w14840) | (~w14805 & w35429) | (~w14840 & w35429);
assign w14843 = ~w14833 & ~w14836;
assign w14844 = ~w14819 & ~w14822;
assign w14845 = ~w14274 & ~w14283;
assign w14846 = ~w14284 & ~w14845;
assign w14847 = ~w14844 & w14846;
assign w14848 = w14844 & ~w14846;
assign w14849 = ~w14847 & ~w14848;
assign w14850 = w5816 & w13177;
assign w14851 = ~w13174 & w35430;
assign w14852 = ~w13011 & w35431;
assign w14853 = ~w14851 & ~w14852;
assign w14854 = ~w14850 & w14853;
assign w14855 = (w14854 & ~w13207) | (w14854 & w35432) | (~w13207 & w35432);
assign w14856 = a_20 & ~w14855;
assign w14857 = (~w13207 & w35433) | (~w13207 & w35434) | (w35433 & w35434);
assign w14858 = ~w14856 & ~w14857;
assign w14859 = w14849 & w14858;
assign w14860 = ~w14849 & ~w14858;
assign w14861 = ~w14859 & ~w14860;
assign w14862 = ~w14843 & w14861;
assign w14863 = w14843 & ~w14861;
assign w14864 = ~w14862 & ~w14863;
assign w14865 = (~w13173 & w35437) | (~w13173 & w35438) | (w35437 & w35438);
assign w14866 = (~w13173 & w35439) | (~w13173 & w35440) | (w35439 & w35440);
assign w14867 = ~w14865 & w14866;
assign w14868 = ~w13487 & ~w14867;
assign w14869 = w14864 & w14868;
assign w14870 = ~w14864 & ~w14868;
assign w14871 = ~w14869 & ~w14870;
assign w14872 = w14842 & ~w14871;
assign w14873 = (~w14847 & ~w14849) | (~w14847 & w35441) | (~w14849 & w35441);
assign w14874 = w13489 & ~w14873;
assign w14875 = ~w13489 & w14873;
assign w14876 = ~w14874 & ~w14875;
assign w14877 = ~w14290 & ~w14299;
assign w14878 = ~w14300 & ~w14877;
assign w14879 = w14876 & w14878;
assign w14880 = (~w14874 & ~w14876) | (~w14874 & w35442) | (~w14876 & w35442);
assign w14881 = ~w14311 & ~w14313;
assign w14882 = ~w14314 & ~w14881;
assign w14883 = ~w14880 & w14882;
assign w14884 = ~w14842 & w14871;
assign w14885 = (~w14862 & ~w14864) | (~w14862 & w35443) | (~w14864 & w35443);
assign w14886 = ~w14876 & ~w14878;
assign w14887 = ~w14879 & ~w14886;
assign w14888 = ~w14885 & w14887;
assign w14889 = ~w14883 & ~w14888;
assign w14890 = ~w14884 & w14889;
assign w14891 = w14872 & w14890;
assign w14892 = w14661 & ~w14663;
assign w14893 = ~w14664 & ~w14892;
assign w14894 = ~w12892 & w35444;
assign w14895 = ~w518 & w12874;
assign w14896 = w4638 & ~w12878;
assign w14897 = ~w14895 & ~w14896;
assign w14898 = ~w14894 & w14897;
assign w14899 = (w14898 & ~w13787) | (w14898 & w35445) | (~w13787 & w35445);
assign w14900 = a_26 & ~w14899;
assign w14901 = (~w13787 & w35446) | (~w13787 & w35447) | (w35446 & w35447);
assign w14902 = ~w14900 & ~w14901;
assign w14903 = w14893 & w14902;
assign w14904 = ~w14541 & w14659;
assign w14905 = ~w14660 & ~w14904;
assign w14906 = w4446 & ~w12860;
assign w14907 = w4068 & w12856;
assign w14908 = w3957 & w12622;
assign w14909 = ~w14907 & ~w14908;
assign w14910 = ~w14906 & w14909;
assign w14911 = (w14910 & ~w14442) | (w14910 & w35448) | (~w14442 & w35448);
assign w14912 = a_29 & ~w14911;
assign w14913 = (~w14442 & w35449) | (~w14442 & w35450) | (w35449 & w35450);
assign w14914 = ~w14912 & ~w14913;
assign w14915 = w14905 & w14914;
assign w14916 = ~w14905 & ~w14914;
assign w14917 = ~w14915 & ~w14916;
assign w14918 = w4666 & ~w12878;
assign w14919 = ~w518 & w12869;
assign w14920 = w4638 & w12874;
assign w14921 = ~w14919 & ~w14920;
assign w14922 = ~w14918 & w14921;
assign w14923 = (w14922 & ~w13771) | (w14922 & w35451) | (~w13771 & w35451);
assign w14924 = ~a_26 & w14923;
assign w14925 = (w13771 & w35452) | (w13771 & w35453) | (w35452 & w35453);
assign w14926 = ~w14924 & ~w14925;
assign w14927 = w14917 & w14926;
assign w14928 = (~w14915 & ~w14917) | (~w14915 & w35454) | (~w14917 & w35454);
assign w14929 = ~w14893 & ~w14902;
assign w14930 = ~w14903 & ~w14929;
assign w14931 = ~w14928 & w14930;
assign w14932 = ~w14903 & ~w14931;
assign w14933 = ~w14670 & ~w14679;
assign w14934 = ~w14680 & ~w14933;
assign w14935 = ~w14932 & w14934;
assign w14936 = w14932 & ~w14934;
assign w14937 = ~w14935 & ~w14936;
assign w14938 = ~w12930 & w35455;
assign w14939 = w5016 & ~w12910;
assign w14940 = ~w12914 & w35456;
assign w14941 = ~w13501 & w35457;
assign w14942 = ~w14939 & ~w14940;
assign w14943 = ~w14938 & w14942;
assign w14944 = ~w14941 & w35458;
assign w14945 = (~a_23 & w14941) | (~a_23 & w35459) | (w14941 & w35459);
assign w14946 = ~w14944 & ~w14945;
assign w14947 = w14937 & ~w14946;
assign w14948 = (~w14935 & ~w14937) | (~w14935 & w35460) | (~w14937 & w35460);
assign w14949 = ~w14686 & w14695;
assign w14950 = ~w14696 & ~w14949;
assign w14951 = ~w14948 & w14950;
assign w14952 = w14948 & ~w14950;
assign w14953 = ~w14951 & ~w14952;
assign w14954 = w5816 & w12604;
assign w14955 = ~w12589 & w35461;
assign w14956 = (w5308 & w12616) | (w5308 & w35462) | (w12616 & w35462);
assign w14957 = ~w14955 & ~w14956;
assign w14958 = ~w14954 & w14957;
assign w14959 = (w14958 & w13288) | (w14958 & w35463) | (w13288 & w35463);
assign w14960 = a_20 & ~w14959;
assign w14961 = (w13288 & w35464) | (w13288 & w35465) | (w35464 & w35465);
assign w14962 = ~w14960 & ~w14961;
assign w14963 = w14953 & w14962;
assign w14964 = (~w14951 & ~w14953) | (~w14951 & w35466) | (~w14953 & w35466);
assign w14965 = w14697 & ~w14699;
assign w14966 = ~w14700 & ~w14965;
assign w14967 = w5816 & w12601;
assign w14968 = w5818 & w12604;
assign w14969 = ~w12589 & w35467;
assign w14970 = ~w14968 & ~w14969;
assign w14971 = ~w14967 & w14970;
assign w14972 = (w14971 & w13140) | (w14971 & w35468) | (w13140 & w35468);
assign w14973 = ~a_20 & w14972;
assign w14974 = (~w13140 & w35469) | (~w13140 & w35470) | (w35469 & w35470);
assign w14975 = ~w14973 & ~w14974;
assign w14976 = w14966 & w14975;
assign w14977 = ~w14966 & ~w14975;
assign w14978 = ~w14976 & ~w14977;
assign w14979 = ~w14964 & w14978;
assign w14980 = w14964 & ~w14978;
assign w14981 = ~w14979 & ~w14980;
assign w14982 = ~w13174 & w35471;
assign w14983 = ~w13011 & w35472;
assign w14984 = w6059 & w12598;
assign w14985 = ~w13205 & w35473;
assign w14986 = ~w14983 & w35474;
assign w14987 = (a_17 & w14985) | (a_17 & w35475) | (w14985 & w35475);
assign w14988 = ~w14985 & w35476;
assign w14989 = ~w14987 & ~w14988;
assign w14990 = w14981 & w14989;
assign w14991 = w14928 & ~w14930;
assign w14992 = ~w14931 & ~w14991;
assign w14993 = ~w12914 & w35477;
assign w14994 = w5080 & ~w12910;
assign w14995 = ~w12905 & w35478;
assign w14996 = (w5017 & w13518) | (w5017 & w35479) | (w13518 & w35479);
assign w14997 = ~w14994 & ~w14995;
assign w14998 = ~w14993 & w14997;
assign w14999 = (a_23 & w14996) | (a_23 & w35480) | (w14996 & w35480);
assign w15000 = ~w14996 & w35481;
assign w15001 = ~w14999 & ~w15000;
assign w15002 = w14992 & w15001;
assign w15003 = ~w14917 & ~w14926;
assign w15004 = ~w14927 & ~w15003;
assign w15005 = w4068 & ~w12630;
assign w15006 = w3957 & ~w12668;
assign w15007 = w4446 & w12622;
assign w15008 = ~w15005 & ~w15006;
assign w15009 = ~w15007 & w15008;
assign w15010 = (w15009 & w14412) | (w15009 & w35482) | (w14412 & w35482);
assign w15011 = a_29 & ~w15010;
assign w15012 = (w14412 & w35483) | (w14412 & w35484) | (w35483 & w35484);
assign w15013 = ~w15011 & ~w15012;
assign w15014 = ~w14628 & ~w14629;
assign w15015 = ~w14644 & w15014;
assign w15016 = w14644 & ~w15014;
assign w15017 = ~w15015 & ~w15016;
assign w15018 = w15013 & w15017;
assign w15019 = (~w14621 & w35485) | (~w14621 & w35486) | (w35485 & w35486);
assign w15020 = ~w14625 & ~w15019;
assign w15021 = w1327 & w12646;
assign w15022 = w668 & ~w12637;
assign w15023 = w1399 & w12651;
assign w15024 = (w12835 & ~w12828) | (w12835 & w31786) | (~w12828 & w31786);
assign w15025 = ~w15024 & w35487;
assign w15026 = (w12649 & w15024) | (w12649 & w35488) | (w15024 & w35488);
assign w15027 = ~w15025 & ~w15026;
assign w15028 = w1478 & ~w15027;
assign w15029 = ~w15022 & w35489;
assign w15030 = ~w15028 & w15029;
assign w15031 = w15020 & ~w15030;
assign w15032 = ~w15020 & w15030;
assign w15033 = ~w15031 & ~w15032;
assign w15034 = w14621 & ~w14623;
assign w15035 = ~w14624 & ~w15034;
assign w15036 = w1327 & w12651;
assign w15037 = w668 & w12646;
assign w15038 = (~w12831 & w12800) | (~w12831 & w31787) | (w12800 & w31787);
assign w15039 = (w31787 & w35490) | (w31787 & w35491) | (w35490 & w35491);
assign w15040 = (~w12826 & ~w12830) | (~w12826 & w35492) | (~w12830 & w35492);
assign w15041 = ~w12657 & ~w15040;
assign w15042 = w12657 & w15040;
assign w15043 = ~w15041 & ~w15042;
assign w15044 = ~w15038 & w15043;
assign w15045 = ~w15039 & ~w15044;
assign w15046 = ~w15044 & w35493;
assign w15047 = (~w15036 & w12830) | (~w15036 & w35494) | (w12830 & w35494);
assign w15048 = ~w15037 & w15047;
assign w15049 = ~w15046 & w15048;
assign w15050 = w15035 & w15049;
assign w15051 = ~w15035 & ~w15049;
assign w15052 = (w14614 & w35495) | (w14614 & w35496) | (w35495 & w35496);
assign w15053 = ~w14620 & ~w15052;
assign w15054 = w4068 & ~w12637;
assign w15055 = w3957 & w12646;
assign w15056 = w4446 & ~w12661;
assign w15057 = ~w15054 & ~w15055;
assign w15058 = ~w15056 & w15057;
assign w15059 = (~w31788 & w35497) | (~w31788 & w35498) | (w35497 & w35498);
assign w15060 = a_29 & ~w15059;
assign w15061 = ~a_29 & w15059;
assign w15062 = ~w15060 & ~w15061;
assign w15063 = w15053 & ~w15062;
assign w15064 = ~w12797 & ~w12826;
assign w15065 = (w12760 & w12818) | (w12760 & w31789) | (w12818 & w31789);
assign w15066 = ~w12742 & w15065;
assign w15067 = w12781 & ~w15066;
assign w15068 = (~w12820 & w15066) | (~w12820 & w35499) | (w15066 & w35499);
assign w15069 = ~w15068 & w35500;
assign w15070 = (w15064 & w15068) | (w15064 & w35501) | (w15068 & w35501);
assign w15071 = ~w15069 & ~w15070;
assign w15072 = w1327 & w12793;
assign w15073 = w1399 & w12789;
assign w15074 = w668 & ~w12830;
assign w15075 = ~w15072 & ~w15073;
assign w15076 = ~w15074 & w15075;
assign w15077 = (w15076 & ~w15071) | (w15076 & w35502) | (~w15071 & w35502);
assign w15078 = ~w81 & ~w88;
assign w15079 = ~w341 & ~w423;
assign w15080 = w15078 & w15079;
assign w15081 = w4008 & w5169;
assign w15082 = w15080 & w15081;
assign w15083 = ~w262 & ~w391;
assign w15084 = ~w547 & w15083;
assign w15085 = w673 & w1722;
assign w15086 = w2549 & w2886;
assign w15087 = w15085 & w15086;
assign w15088 = w987 & w15084;
assign w15089 = w2578 & w4365;
assign w15090 = w15088 & w15089;
assign w15091 = w2969 & w15087;
assign w15092 = w13904 & w15082;
assign w15093 = w15091 & w15092;
assign w15094 = w15090 & w15093;
assign w15095 = w1985 & w15094;
assign w15096 = w5200 & w15095;
assign w15097 = (~w15071 & w35503) | (~w15071 & w35504) | (w35503 & w35504);
assign w15098 = ~w12794 & ~w12820;
assign w15099 = (~w15098 & w15066) | (~w15098 & w35505) | (w15066 & w35505);
assign w15100 = ~w15066 & w35506;
assign w15101 = ~w15099 & ~w15100;
assign w15102 = w1327 & w12789;
assign w15103 = ~w12770 & w35507;
assign w15104 = w668 & w12793;
assign w15105 = ~w15102 & ~w15103;
assign w15106 = ~w15104 & w15105;
assign w15107 = ~w94 & ~w580;
assign w15108 = w448 & w15107;
assign w15109 = w1820 & w2102;
assign w15110 = w2989 & w12967;
assign w15111 = w15109 & w15110;
assign w15112 = w4730 & w15108;
assign w15113 = w14351 & w15112;
assign w15114 = w2714 & w15111;
assign w15115 = w15113 & w15114;
assign w15116 = w787 & w6122;
assign w15117 = w15115 & w15116;
assign w15118 = w1887 & w15117;
assign w15119 = w2214 & w15118;
assign w15120 = (w15101 & w35509) | (w15101 & w35510) | (w35509 & w35510);
assign w15121 = ~w12775 & w12818;
assign w15122 = ~w12761 & w15121;
assign w15123 = ~w12741 & ~w12775;
assign w15124 = ~w12729 & w15123;
assign w15125 = ~w12760 & ~w12775;
assign w15126 = ~w12818 & ~w15125;
assign w15127 = ~w15124 & w15126;
assign w15128 = ~w15122 & ~w15127;
assign w15129 = w1478 & ~w15128;
assign w15130 = w668 & w12789;
assign w15131 = w1399 & ~w12774;
assign w15132 = ~w12770 & w35511;
assign w15133 = ~w15130 & w35512;
assign w15134 = ~w166 & ~w1043;
assign w15135 = w2991 & w15134;
assign w15136 = w3495 & w4815;
assign w15137 = w15135 & w15136;
assign w15138 = w1294 & w2287;
assign w15139 = w2606 & w3213;
assign w15140 = w4851 & w15139;
assign w15141 = w15137 & w15138;
assign w15142 = w15140 & w15141;
assign w15143 = w2493 & w15142;
assign w15144 = w3384 & w15143;
assign w15145 = w14597 & w15144;
assign w15146 = (~w15145 & w15129) | (~w15145 & w35513) | (w15129 & w35513);
assign w15147 = ~w15129 & w35514;
assign w15148 = ~w15146 & ~w15147;
assign w15149 = ~w12730 & ~w12736;
assign w15150 = ~w12743 & ~w15149;
assign w15151 = w12728 & ~w15150;
assign w15152 = w12732 & w12739;
assign w15153 = ~w12736 & w15152;
assign w15154 = (~w15153 & ~w12717) | (~w15153 & w31790) | (~w12717 & w31790);
assign w15155 = w15150 & ~w15152;
assign w15156 = (w15155 & ~w12717) | (w15155 & w31791) | (~w12717 & w31791);
assign w15157 = w15154 & ~w15156;
assign w15158 = w1327 & w12732;
assign w15159 = w1399 & w12739;
assign w15160 = w668 & ~w12774;
assign w15161 = ~w15158 & ~w15159;
assign w15162 = ~w15160 & w15161;
assign w15163 = w984 & w6743;
assign w15164 = ~w246 & ~w538;
assign w15165 = ~w895 & w15164;
assign w15166 = ~w378 & w1329;
assign w15167 = w1987 & w4712;
assign w15168 = w6116 & w15167;
assign w15169 = w2315 & w15166;
assign w15170 = w13725 & w15165;
assign w15171 = w15169 & w15170;
assign w15172 = w4371 & w15168;
assign w15173 = w15171 & w15172;
assign w15174 = w6691 & w15173;
assign w15175 = w550 & ~w582;
assign w15176 = w13549 & w15175;
assign w15177 = w712 & w989;
assign w15178 = w3868 & w5512;
assign w15179 = w14579 & w15178;
assign w15180 = w15176 & w15177;
assign w15181 = w1297 & w14030;
assign w15182 = w15180 & w15181;
assign w15183 = w15179 & w15182;
assign w15184 = ~w152 & ~w357;
assign w15185 = w935 & w15184;
assign w15186 = w4275 & w6570;
assign w15187 = w13565 & w15186;
assign w15188 = w1127 & w15185;
assign w15189 = w1263 & w3573;
assign w15190 = w14560 & w15163;
assign w15191 = w15189 & w15190;
assign w15192 = w15187 & w15188;
assign w15193 = w1272 & w6526;
assign w15194 = w15192 & w15193;
assign w15195 = w15191 & w15194;
assign w15196 = w13747 & w15195;
assign w15197 = w15174 & w15183;
assign w15198 = w15196 & w15197;
assign w15199 = (w15157 & w35516) | (w15157 & w35517) | (w35516 & w35517);
assign w15200 = w1478 & ~w12728;
assign w15201 = w1399 & w12701;
assign w15202 = w668 & w12732;
assign w15203 = ~w12717 & w12728;
assign w15204 = ~w12717 & w31792;
assign w15205 = (~w15201 & ~w12739) | (~w15201 & w35518) | (~w12739 & w35518);
assign w15206 = ~w15202 & w15205;
assign w15207 = (w15206 & ~w12717) | (w15206 & w35519) | (~w12717 & w35519);
assign w15208 = w1464 & w2689;
assign w15209 = ~w180 & ~w264;
assign w15210 = ~w540 & w15209;
assign w15211 = w474 & w866;
assign w15212 = w1639 & w2035;
assign w15213 = w2087 & w3365;
assign w15214 = w15212 & w15213;
assign w15215 = w15210 & w15211;
assign w15216 = w1070 & w4002;
assign w15217 = w15208 & w15216;
assign w15218 = w15214 & w15215;
assign w15219 = w15217 & w15218;
assign w15220 = w3582 & w15219;
assign w15221 = w14054 & w15220;
assign w15222 = ~w378 & ~w1040;
assign w15223 = w293 & ~w1051;
assign w15224 = w808 & w822;
assign w15225 = w993 & w1113;
assign w15226 = w1206 & w1721;
assign w15227 = w2700 & w2971;
assign w15228 = w3274 & w3675;
assign w15229 = w3686 & w4364;
assign w15230 = w15222 & w15229;
assign w15231 = w15227 & w15228;
assign w15232 = w15225 & w15226;
assign w15233 = w15223 & w15224;
assign w15234 = w4756 & w15233;
assign w15235 = w15231 & w15232;
assign w15236 = w3407 & w15230;
assign w15237 = w15235 & w15236;
assign w15238 = w15234 & w15237;
assign w15239 = w3988 & w15238;
assign w15240 = w15221 & w15239;
assign w15241 = (~w15240 & ~w15207) | (~w15240 & w31793) | (~w15207 & w31793);
assign w15242 = w15207 & w31794;
assign w15243 = ~w737 & w2512;
assign w15244 = w13452 & w15243;
assign w15245 = w433 & ~w649;
assign w15246 = w13741 & w15245;
assign w15247 = w592 & w15246;
assign w15248 = ~w734 & ~w878;
assign w15249 = ~w45 & w398;
assign w15250 = w1113 & w1764;
assign w15251 = w3740 & w13563;
assign w15252 = w15248 & w15251;
assign w15253 = w15249 & w15250;
assign w15254 = w3877 & w15253;
assign w15255 = w15244 & w15252;
assign w15256 = w15254 & w15255;
assign w15257 = w14005 & w15247;
assign w15258 = w15256 & w15257;
assign w15259 = ~w399 & w3575;
assign w15260 = ~w116 & ~w741;
assign w15261 = ~w907 & w15260;
assign w15262 = w3344 & w15261;
assign w15263 = w2011 & w3917;
assign w15264 = w4297 & w15259;
assign w15265 = w15263 & w15264;
assign w15266 = w328 & w15262;
assign w15267 = w1818 & w15266;
assign w15268 = w15265 & w15267;
assign w15269 = w2870 & w15268;
assign w15270 = w983 & w15258;
assign w15271 = w15269 & w15270;
assign w15272 = w1327 & w12701;
assign w15273 = w1399 & w12702;
assign w15274 = w668 & w12739;
assign w15275 = ~w15272 & ~w15273;
assign w15276 = (~w15271 & w15274) | (~w15271 & w35520) | (w15274 & w35520);
assign w15277 = ~w12704 & w12714;
assign w15278 = ~w12715 & ~w15277;
assign w15279 = w1478 & ~w15271;
assign w15280 = (~w15276 & w15278) | (~w15276 & w35521) | (w15278 & w35521);
assign w15281 = w12694 & ~w12695;
assign w15282 = ~w12696 & ~w15281;
assign w15283 = ~w12689 & w15282;
assign w15284 = w1478 & w15283;
assign w15285 = w1478 & ~w12681;
assign w15286 = w12688 & w15285;
assign w15287 = ~w15282 & w15286;
assign w15288 = w668 & ~w11825;
assign w15289 = ~w12699 & w15288;
assign w15290 = w1327 & ~w12675;
assign w15291 = ~w12674 & w15290;
assign w15292 = w1327 & ~w11501;
assign w15293 = w11677 & w11683;
assign w15294 = w15292 & w15293;
assign w15295 = w668 & w11825;
assign w15296 = w12699 & w15295;
assign w15297 = w12684 & w31795;
assign w15298 = ~w15291 & ~w15294;
assign w15299 = ~w15289 & w15298;
assign w15300 = ~w15296 & ~w15297;
assign w15301 = w15299 & w15300;
assign w15302 = ~w15287 & w15301;
assign w15303 = ~w15284 & w15302;
assign w15304 = ~w123 & ~w127;
assign w15305 = ~w177 & ~w214;
assign w15306 = ~w282 & w15305;
assign w15307 = w564 & w15304;
assign w15308 = w15306 & w15307;
assign w15309 = w1282 & w4387;
assign w15310 = w15308 & w15309;
assign w15311 = w1234 & w2653;
assign w15312 = w6757 & w15311;
assign w15313 = w5618 & w15310;
assign w15314 = w15312 & w15313;
assign w15315 = w692 & w850;
assign w15316 = w15314 & w15315;
assign w15317 = w4362 & w15316;
assign w15318 = ~w15303 & ~w15317;
assign w15319 = w11332 & ~w11338;
assign w15320 = ~w10849 & ~w11332;
assign w15321 = ~w15319 & ~w15320;
assign w15322 = w11499 & ~w15321;
assign w15323 = ~w11499 & w15321;
assign w15324 = ~w15322 & ~w15323;
assign w15325 = w1478 & ~w15324;
assign w15326 = w668 & ~w11501;
assign w15327 = w12684 & w15326;
assign w15328 = w1327 & w12679;
assign w15329 = ~w15327 & ~w15328;
assign w15330 = ~w15325 & w15329;
assign w15331 = ~w81 & ~w572;
assign w15332 = w1260 & w15331;
assign w15333 = w1505 & w1872;
assign w15334 = w2809 & w4163;
assign w15335 = w15248 & w15334;
assign w15336 = w15332 & w15333;
assign w15337 = w915 & w1242;
assign w15338 = w1968 & w3737;
assign w15339 = w3992 & w15338;
assign w15340 = w15336 & w15337;
assign w15341 = w15335 & w15340;
assign w15342 = w14578 & w15339;
assign w15343 = w15341 & w15342;
assign w15344 = w486 & w15343;
assign w15345 = w14000 & w15344;
assign w15346 = w15330 & ~w15345;
assign w15347 = ~w652 & w1076;
assign w15348 = w1309 & w15347;
assign w15349 = w6741 & w15348;
assign w15350 = ~w149 & ~w394;
assign w15351 = w821 & w2082;
assign w15352 = w4312 & w6155;
assign w15353 = w15350 & w15352;
assign w15354 = w15351 & w15353;
assign w15355 = ~w404 & w620;
assign w15356 = w1524 & w1567;
assign w15357 = w1607 & w4884;
assign w15358 = w15356 & w15357;
assign w15359 = w1168 & w15355;
assign w15360 = w1339 & w6115;
assign w15361 = w15359 & w15360;
assign w15362 = w15358 & w15361;
assign w15363 = w15349 & w15354;
assign w15364 = w15362 & w15363;
assign w15365 = w474 & w1081;
assign w15366 = w1153 & w2445;
assign w15367 = w15365 & w15366;
assign w15368 = w2160 & w15367;
assign w15369 = w1411 & w3016;
assign w15370 = w3062 & w3098;
assign w15371 = w15369 & w15370;
assign w15372 = w15368 & w15371;
assign w15373 = w6569 & w15372;
assign w15374 = w2769 & w15364;
assign w15375 = w15373 & w15374;
assign w15376 = (~w15375 & ~w12679) | (~w15375 & w31796) | (~w12679 & w31796);
assign w15377 = ~w15327 & w15376;
assign w15378 = ~w15325 & w15377;
assign w15379 = ~w15345 & ~w15375;
assign w15380 = w15345 & w15375;
assign w15381 = ~w15379 & ~w15380;
assign w15382 = ~w15378 & w15381;
assign w15383 = ~w15346 & ~w15382;
assign w15384 = ~w11500 & ~w12682;
assign w15385 = ~w12679 & w15384;
assign w15386 = w12702 & ~w15385;
assign w15387 = w12702 & w31797;
assign w15388 = w1478 & w15385;
assign w15389 = ~w12702 & w15388;
assign w15390 = w1399 & w12679;
assign w15391 = w668 & ~w12675;
assign w15392 = ~w12674 & w15391;
assign w15393 = w15293 & w15326;
assign w15394 = w12684 & w15292;
assign w15395 = ~w15390 & ~w15392;
assign w15396 = ~w15393 & ~w15394;
assign w15397 = w15395 & w15396;
assign w15398 = ~w15389 & w15397;
assign w15399 = ~w15387 & w15398;
assign w15400 = ~w15383 & ~w15399;
assign w15401 = ~w15330 & w15379;
assign w15402 = ~w15400 & ~w15401;
assign w15403 = w15303 & w15317;
assign w15404 = ~w15402 & ~w15403;
assign w15405 = ~w15318 & ~w15404;
assign w15406 = w1478 & ~w15278;
assign w15407 = ~w15274 & w35522;
assign w15408 = ~w15406 & w15407;
assign w15409 = ~w15405 & ~w15408;
assign w15410 = w15280 & ~w15409;
assign w15411 = (~w15241 & w15410) | (~w15241 & w31798) | (w15410 & w31798);
assign w15412 = ~w15199 & ~w15411;
assign w15413 = (~w15157 & w35523) | (~w15157 & w35524) | (w35523 & w35524);
assign w15414 = ~w252 & ~w708;
assign w15415 = ~w422 & ~w597;
assign w15416 = w1281 & w15415;
assign w15417 = w3583 & w4849;
assign w15418 = w15414 & w15417;
assign w15419 = w712 & w15416;
assign w15420 = w2287 & w6611;
assign w15421 = w15419 & w15420;
assign w15422 = w15418 & w15421;
assign w15423 = w579 & w4402;
assign w15424 = w15349 & w15423;
assign w15425 = w15422 & w15424;
assign w15426 = w4190 & w15425;
assign w15427 = ~w12770 & w35525;
assign w15428 = w1399 & w12732;
assign w15429 = w1327 & ~w12774;
assign w15430 = ~w15427 & ~w15428;
assign w15431 = (~w15426 & ~w15430) | (~w15426 & w35526) | (~w15430 & w35526);
assign w15432 = ~w12746 & w12759;
assign w15433 = ~w12741 & w12759;
assign w15434 = (~w15432 & w12729) | (~w15432 & w31799) | (w12729 & w31799);
assign w15435 = ~w12761 & w15434;
assign w15436 = w1478 & ~w15426;
assign w15437 = (~w15431 & ~w15435) | (~w15431 & w35527) | (~w15435 & w35527);
assign w15438 = ~w15413 & w15437;
assign w15439 = w1478 & w15435;
assign w15440 = w15430 & w35528;
assign w15441 = ~w15439 & w15440;
assign w15442 = (~w15441 & w15412) | (~w15441 & w35529) | (w15412 & w35529);
assign w15443 = w15148 & w15442;
assign w15444 = (~w15101 & w35530) | (~w15101 & w35531) | (w35530 & w35531);
assign w15445 = ~w15146 & ~w15444;
assign w15446 = (~w15120 & w15443) | (~w15120 & w35532) | (w15443 & w35532);
assign w15447 = ~w15077 & ~w15096;
assign w15448 = ~w15097 & ~w15447;
assign w15449 = ~w15446 & w15448;
assign w15450 = (~w15097 & w15446) | (~w15097 & w35533) | (w15446 & w35533);
assign w15451 = ~w15053 & w15062;
assign w15452 = ~w15063 & ~w15451;
assign w15453 = ~w15450 & w15452;
assign w15454 = (~w15063 & ~w15452) | (~w15063 & w35534) | (~w15452 & w35534);
assign w15455 = (~w15050 & w15454) | (~w15050 & w35535) | (w15454 & w35535);
assign w15456 = w15033 & w15455;
assign w15457 = ~w15013 & ~w15017;
assign w15458 = ~w15018 & ~w15457;
assign w15459 = (w15455 & w35537) | (w15455 & w35538) | (w35537 & w35538);
assign w15460 = ~w14647 & ~w14648;
assign w15461 = w14657 & w15460;
assign w15462 = ~w14657 & ~w15460;
assign w15463 = ~w15461 & ~w15462;
assign w15464 = ~w15459 & w35539;
assign w15465 = (w15463 & w15459) | (w15463 & w35540) | (w15459 & w35540);
assign w15466 = ~w15464 & ~w15465;
assign w15467 = w4666 & w12874;
assign w15468 = w4638 & w12869;
assign w15469 = ~w518 & ~w12860;
assign w15470 = w1226 & w13965;
assign w15471 = ~w15469 & w35541;
assign w15472 = ~w15470 & w35542;
assign w15473 = (~a_26 & w15470) | (~a_26 & w35543) | (w15470 & w35543);
assign w15474 = ~w15472 & ~w15473;
assign w15475 = w15466 & w15474;
assign w15476 = (~w15464 & ~w15466) | (~w15464 & w35544) | (~w15466 & w35544);
assign w15477 = w15004 & w15476;
assign w15478 = ~w15004 & ~w15476;
assign w15479 = ~w15477 & ~w15478;
assign w15480 = ~w12905 & w35545;
assign w15481 = ~w12892 & w35546;
assign w15482 = w5286 & ~w12910;
assign w15483 = w5017 & w13815;
assign w15484 = ~w15482 & w35547;
assign w15485 = ~w15483 & w35548;
assign w15486 = (a_23 & w15483) | (a_23 & w35549) | (w15483 & w35549);
assign w15487 = ~w15485 & ~w15486;
assign w15488 = w15479 & w15487;
assign w15489 = (~w15477 & ~w15479) | (~w15477 & w35550) | (~w15479 & w35550);
assign w15490 = ~w14992 & ~w15001;
assign w15491 = ~w15002 & ~w15490;
assign w15492 = ~w15489 & w15491;
assign w15493 = ~w15002 & ~w15492;
assign w15494 = ~w14937 & w14946;
assign w15495 = ~w14947 & ~w15494;
assign w15496 = ~w15493 & w15495;
assign w15497 = w15493 & ~w15495;
assign w15498 = ~w15496 & ~w15497;
assign w15499 = ~w12589 & w35551;
assign w15500 = (w5308 & w12612) | (w5308 & w35552) | (w12612 & w35552);
assign w15501 = (w5818 & w12616) | (w5818 & w35553) | (w12616 & w35553);
assign w15502 = ~w15499 & ~w15500;
assign w15503 = ~w15501 & w15502;
assign w15504 = (w15503 & ~w13123) | (w15503 & w35554) | (~w13123 & w35554);
assign w15505 = a_20 & ~w15504;
assign w15506 = (~w13123 & w35555) | (~w13123 & w35556) | (w35555 & w35556);
assign w15507 = ~w15505 & ~w15506;
assign w15508 = w15498 & w15507;
assign w15509 = (~w15496 & ~w15498) | (~w15496 & w35557) | (~w15498 & w35557);
assign w15510 = ~w14953 & ~w14962;
assign w15511 = ~w14963 & ~w15510;
assign w15512 = ~w15509 & w15511;
assign w15513 = w15509 & ~w15511;
assign w15514 = ~w15512 & ~w15513;
assign w15515 = ~w13011 & w35558;
assign w15516 = w6061 & w12598;
assign w15517 = w6059 & w12601;
assign w15518 = ~w15516 & ~w15517;
assign w15519 = ~w15515 & w15518;
assign w15520 = (w15519 & w13021) | (w15519 & w35559) | (w13021 & w35559);
assign w15521 = ~a_17 & w15520;
assign w15522 = (~w13021 & w35560) | (~w13021 & w35561) | (w35560 & w35561);
assign w15523 = ~w15521 & ~w15522;
assign w15524 = w15514 & w15523;
assign w15525 = (~w15512 & ~w15514) | (~w15512 & w35562) | (~w15514 & w35562);
assign w15526 = ~w14981 & ~w14989;
assign w15527 = ~w14990 & ~w15526;
assign w15528 = ~w15525 & w15527;
assign w15529 = (~w14990 & ~w15527) | (~w14990 & w35563) | (~w15527 & w35563);
assign w15530 = (~w14976 & ~w14978) | (~w14976 & w35564) | (~w14978 & w35564);
assign w15531 = ~w14738 & ~w14747;
assign w15532 = ~w14748 & ~w15531;
assign w15533 = ~w15530 & w15532;
assign w15534 = w15530 & ~w15532;
assign w15535 = ~w15533 & ~w15534;
assign w15536 = w6304 & w13177;
assign w15537 = ~w13174 & w35565;
assign w15538 = ~w13011 & w35566;
assign w15539 = ~w15537 & ~w15538;
assign w15540 = ~w15536 & w15539;
assign w15541 = (w15540 & ~w13207) | (w15540 & w35567) | (~w13207 & w35567);
assign w15542 = a_17 & ~w15541;
assign w15543 = (~w13207 & w35568) | (~w13207 & w35569) | (w35568 & w35569);
assign w15544 = ~w15542 & ~w15543;
assign w15545 = w15535 & w15544;
assign w15546 = ~w15535 & ~w15544;
assign w15547 = ~w15545 & ~w15546;
assign w15548 = ~w15529 & w15547;
assign w15549 = w15529 & ~w15547;
assign w15550 = ~w15548 & ~w15549;
assign w15551 = (~w13173 & w35572) | (~w13173 & w35573) | (w35572 & w35573);
assign w15552 = (~w13173 & w35574) | (~w13173 & w35575) | (w35574 & w35575);
assign w15553 = ~w15551 & w15552;
assign w15554 = ~w13584 & ~w15553;
assign w15555 = w15550 & w15554;
assign w15556 = (~w15548 & ~w15550) | (~w15548 & w35576) | (~w15550 & w35576);
assign w15557 = (~w15533 & ~w15535) | (~w15533 & w35577) | (~w15535 & w35577);
assign w15558 = w13586 & ~w15557;
assign w15559 = ~w13586 & w15557;
assign w15560 = ~w15558 & ~w15559;
assign w15561 = ~w14786 & ~w14795;
assign w15562 = ~w14796 & ~w15561;
assign w15563 = w15560 & w15562;
assign w15564 = ~w15560 & ~w15562;
assign w15565 = ~w15563 & ~w15564;
assign w15566 = ~w15556 & w15565;
assign w15567 = w15489 & ~w15491;
assign w15568 = ~w15492 & ~w15567;
assign w15569 = (w5816 & w12616) | (w5816 & w35578) | (w12616 & w35578);
assign w15570 = (w5818 & w12612) | (w5818 & w35579) | (w12612 & w35579);
assign w15571 = ~w12930 & w35580;
assign w15572 = ~w15570 & ~w15571;
assign w15573 = ~w15569 & w15572;
assign w15574 = (w15573 & ~w13389) | (w15573 & w35581) | (~w13389 & w35581);
assign w15575 = a_20 & ~w15574;
assign w15576 = (~w13389 & w35582) | (~w13389 & w35583) | (w35582 & w35583);
assign w15577 = ~w15575 & ~w15576;
assign w15578 = w15568 & w15577;
assign w15579 = ~w15479 & ~w15487;
assign w15580 = ~w15488 & ~w15579;
assign w15581 = (~w15455 & w35584) | (~w15455 & w35585) | (w35584 & w35585);
assign w15582 = ~w15459 & ~w15581;
assign w15583 = ~w518 & w12856;
assign w15584 = w4666 & w12869;
assign w15585 = (~w15583 & w12860) | (~w15583 & w35586) | (w12860 & w35586);
assign w15586 = ~w15584 & w15585;
assign w15587 = (w15586 & ~w13979) | (w15586 & w35587) | (~w13979 & w35587);
assign w15588 = ~a_26 & w15587;
assign w15589 = (w13979 & w35588) | (w13979 & w35589) | (w35588 & w35589);
assign w15590 = ~w15588 & ~w15589;
assign w15591 = ~w15582 & ~w15590;
assign w15592 = (~w15454 & w35590) | (~w15454 & w35591) | (w35590 & w35591);
assign w15593 = w4446 & ~w12630;
assign w15594 = w3957 & ~w12661;
assign w15595 = w4068 & ~w12668;
assign w15596 = ~w15594 & ~w15595;
assign w15597 = ~w15593 & w15596;
assign w15598 = (w15597 & w14535) | (w15597 & w35592) | (w14535 & w35592);
assign w15599 = a_29 & w15598;
assign w15600 = (~w14535 & w35593) | (~w14535 & w35594) | (w35593 & w35594);
assign w15601 = ~w15599 & ~w15600;
assign w15602 = ~w15456 & w35595;
assign w15603 = (w15601 & w15456) | (w15601 & w35596) | (w15456 & w35596);
assign w15604 = ~w15602 & ~w15603;
assign w15605 = w4666 & ~w12860;
assign w15606 = ~w518 & w12622;
assign w15607 = w4638 & w12856;
assign w15608 = ~w15606 & ~w15607;
assign w15609 = ~w15605 & w15608;
assign w15610 = (w15609 & ~w14442) | (w15609 & w35597) | (~w14442 & w35597);
assign w15611 = ~a_26 & w15610;
assign w15612 = (w14442 & w35598) | (w14442 & w35599) | (w35598 & w35599);
assign w15613 = ~w15611 & ~w15612;
assign w15614 = w15604 & w15613;
assign w15615 = (~w15602 & ~w15604) | (~w15602 & w35600) | (~w15604 & w35600);
assign w15616 = w15582 & w15590;
assign w15617 = ~w15591 & ~w15616;
assign w15618 = w15615 & w15617;
assign w15619 = ~w15591 & ~w15618;
assign w15620 = ~w15466 & ~w15474;
assign w15621 = ~w15475 & ~w15620;
assign w15622 = w15619 & ~w15621;
assign w15623 = ~w15619 & w15621;
assign w15624 = ~w15622 & ~w15623;
assign w15625 = ~w12905 & w35601;
assign w15626 = w5016 & ~w12878;
assign w15627 = ~w12892 & w35602;
assign w15628 = ~w13598 & w35603;
assign w15629 = ~w15626 & ~w15627;
assign w15630 = ~w15625 & w15629;
assign w15631 = ~w15628 & w35604;
assign w15632 = (a_23 & w15628) | (a_23 & w35605) | (w15628 & w35605);
assign w15633 = ~w15631 & ~w15632;
assign w15634 = w15624 & w15633;
assign w15635 = (~w15622 & ~w15624) | (~w15622 & w35606) | (~w15624 & w35606);
assign w15636 = w15580 & ~w15635;
assign w15637 = ~w15580 & w15635;
assign w15638 = ~w15636 & ~w15637;
assign w15639 = (w5816 & w12612) | (w5816 & w35607) | (w12612 & w35607);
assign w15640 = ~w12914 & w35608;
assign w15641 = ~w12930 & w35609;
assign w15642 = ~w15640 & ~w15641;
assign w15643 = ~w15639 & w15642;
assign w15644 = (w15643 & ~w13375) | (w15643 & w35610) | (~w13375 & w35610);
assign w15645 = ~a_20 & w15644;
assign w15646 = (w13375 & w35611) | (w13375 & w35612) | (w35611 & w35612);
assign w15647 = ~w15645 & ~w15646;
assign w15648 = w15638 & w15647;
assign w15649 = (~w15636 & ~w15638) | (~w15636 & w35613) | (~w15638 & w35613);
assign w15650 = ~w15568 & ~w15577;
assign w15651 = ~w15578 & ~w15650;
assign w15652 = ~w15649 & w15651;
assign w15653 = ~w15578 & ~w15652;
assign w15654 = ~w15498 & ~w15507;
assign w15655 = ~w15508 & ~w15654;
assign w15656 = ~w15653 & w15655;
assign w15657 = w15653 & ~w15655;
assign w15658 = ~w15656 & ~w15657;
assign w15659 = w6304 & w12598;
assign w15660 = w6061 & w12601;
assign w15661 = w6059 & w12604;
assign w15662 = ~w15660 & ~w15661;
assign w15663 = ~w15659 & w15662;
assign w15664 = (w15663 & ~w12961) | (w15663 & w35614) | (~w12961 & w35614);
assign w15665 = ~a_17 & w15664;
assign w15666 = (w12961 & w35615) | (w12961 & w35616) | (w35615 & w35616);
assign w15667 = ~w15665 & ~w15666;
assign w15668 = w15658 & w15667;
assign w15669 = (~w15656 & ~w15658) | (~w15656 & w35617) | (~w15658 & w35617);
assign w15670 = ~w15514 & ~w15523;
assign w15671 = ~w15524 & ~w15670;
assign w15672 = ~w15669 & w15671;
assign w15673 = w15669 & ~w15671;
assign w15674 = ~w15672 & ~w15673;
assign w15675 = w6998 & w13177;
assign w15676 = ~w13174 & w35618;
assign w15677 = (w13173 & w35619) | (w13173 & w35620) | (w35619 & w35620);
assign w15678 = ~w15676 & ~w15677;
assign w15679 = ~w15675 & w15678;
assign w15680 = (w15679 & w13264) | (w15679 & w35621) | (w13264 & w35621);
assign w15681 = ~a_14 & w15680;
assign w15682 = (~w13264 & w35622) | (~w13264 & w35623) | (w35622 & w35623);
assign w15683 = ~w15681 & ~w15682;
assign w15684 = w15674 & w15683;
assign w15685 = (~w15672 & ~w15674) | (~w15672 & w35624) | (~w15674 & w35624);
assign w15686 = w6446 & w13177;
assign w15687 = (w13201 & w35627) | (w13201 & w35628) | (w35627 & w35628);
assign w15688 = (~w13173 & w35629) | (~w13173 & w35630) | (w35629 & w35630);
assign w15689 = ~w15686 & w15688;
assign w15690 = (a_14 & w15687) | (a_14 & w35631) | (w15687 & w35631);
assign w15691 = ~w15687 & w35632;
assign w15692 = ~w15690 & ~w15691;
assign w15693 = ~w15685 & w15692;
assign w15694 = w15525 & ~w15527;
assign w15695 = ~w15528 & ~w15694;
assign w15696 = w15685 & ~w15692;
assign w15697 = ~w15693 & ~w15696;
assign w15698 = w15695 & w15697;
assign w15699 = (~w15693 & ~w15697) | (~w15693 & w35633) | (~w15697 & w35633);
assign w15700 = ~w15550 & ~w15554;
assign w15701 = ~w15555 & ~w15700;
assign w15702 = ~w15699 & w15701;
assign w15703 = ~w15566 & ~w15702;
assign w15704 = w15649 & ~w15651;
assign w15705 = ~w15652 & ~w15704;
assign w15706 = w6304 & w12601;
assign w15707 = w6061 & w12604;
assign w15708 = ~w12589 & w35634;
assign w15709 = ~w15707 & ~w15708;
assign w15710 = ~w15706 & w15709;
assign w15711 = (w15710 & w13140) | (w15710 & w35635) | (w13140 & w35635);
assign w15712 = ~a_17 & w15711;
assign w15713 = (~w13140 & w35636) | (~w13140 & w35637) | (w35636 & w35637);
assign w15714 = ~w15712 & ~w15713;
assign w15715 = w15705 & w15714;
assign w15716 = ~w15638 & ~w15647;
assign w15717 = ~w15648 & ~w15716;
assign w15718 = ~w12930 & w35638;
assign w15719 = w5308 & ~w12910;
assign w15720 = ~w12914 & w35639;
assign w15721 = ~w13501 & w35640;
assign w15722 = ~w15719 & ~w15720;
assign w15723 = ~w15718 & w15722;
assign w15724 = ~w15721 & w35641;
assign w15725 = (a_20 & w15721) | (a_20 & w35642) | (w15721 & w35642);
assign w15726 = ~w15724 & ~w15725;
assign w15727 = ~w15615 & ~w15617;
assign w15728 = ~w15618 & ~w15727;
assign w15729 = ~w12892 & w35643;
assign w15730 = w5016 & w12874;
assign w15731 = w5080 & ~w12878;
assign w15732 = ~w15730 & ~w15731;
assign w15733 = ~w15729 & w15732;
assign w15734 = (w15733 & ~w13787) | (w15733 & w35644) | (~w13787 & w35644);
assign w15735 = a_23 & w15734;
assign w15736 = (w13787 & w35645) | (w13787 & w35646) | (w35645 & w35646);
assign w15737 = ~w15735 & ~w15736;
assign w15738 = ~w15728 & ~w15737;
assign w15739 = w15728 & w15737;
assign w15740 = w4666 & w12856;
assign w15741 = ~w518 & ~w12630;
assign w15742 = w4638 & w12622;
assign w15743 = ~w15741 & ~w15742;
assign w15744 = ~w15740 & w15743;
assign w15745 = (w15744 & ~w14091) | (w15744 & w35647) | (~w14091 & w35647);
assign w15746 = ~a_26 & w15745;
assign w15747 = (w14091 & w35648) | (w14091 & w35649) | (w35648 & w35649);
assign w15748 = ~w15746 & ~w15747;
assign w15749 = ~w15050 & ~w15051;
assign w15750 = w4446 & ~w12668;
assign w15751 = w3957 & ~w12637;
assign w15752 = w4068 & ~w12661;
assign w15753 = ~w15751 & ~w15752;
assign w15754 = ~w15750 & w15753;
assign w15755 = (w15754 & ~w14393) | (w15754 & w35650) | (~w14393 & w35650);
assign w15756 = ~a_29 & w15755;
assign w15757 = (w14393 & w35651) | (w14393 & w35652) | (w35651 & w35652);
assign w15758 = ~w15756 & ~w15757;
assign w15759 = w15749 & ~w15758;
assign w15760 = ~w15749 & w15758;
assign w15761 = ~w15759 & ~w15760;
assign w15762 = w15454 & w15761;
assign w15763 = ~w15454 & ~w15761;
assign w15764 = ~w15762 & ~w15763;
assign w15765 = w15748 & ~w15764;
assign w15766 = w15758 & w15764;
assign w15767 = ~w15765 & ~w15766;
assign w15768 = w5286 & ~w12878;
assign w15769 = w5016 & w12869;
assign w15770 = w5080 & w12874;
assign w15771 = ~w15769 & ~w15770;
assign w15772 = ~w15768 & w15771;
assign w15773 = (w15772 & ~w13771) | (w15772 & w35653) | (~w13771 & w35653);
assign w15774 = a_23 & w15773;
assign w15775 = (w13771 & w35654) | (w13771 & w35655) | (w35654 & w35655);
assign w15776 = ~w15774 & ~w15775;
assign w15777 = w15767 & w15776;
assign w15778 = ~w15604 & ~w15613;
assign w15779 = ~w15614 & ~w15778;
assign w15780 = ~w15767 & ~w15776;
assign w15781 = ~w15777 & ~w15780;
assign w15782 = ~w15779 & w15781;
assign w15783 = ~w15777 & ~w15782;
assign w15784 = ~w15739 & w15783;
assign w15785 = (w15726 & w15784) | (w15726 & w35656) | (w15784 & w35656);
assign w15786 = ~w15624 & ~w15633;
assign w15787 = ~w15634 & ~w15786;
assign w15788 = ~w15784 & w35657;
assign w15789 = ~w15785 & ~w15788;
assign w15790 = w15787 & w15789;
assign w15791 = ~w15785 & ~w15790;
assign w15792 = ~w15717 & w15791;
assign w15793 = w15717 & ~w15791;
assign w15794 = ~w15792 & ~w15793;
assign w15795 = w6304 & w12604;
assign w15796 = ~w12589 & w35658;
assign w15797 = (w6059 & w12616) | (w6059 & w35659) | (w12616 & w35659);
assign w15798 = ~w15796 & ~w15797;
assign w15799 = ~w15795 & w15798;
assign w15800 = (w15799 & w13288) | (w15799 & w35660) | (w13288 & w35660);
assign w15801 = a_17 & ~w15800;
assign w15802 = (w13288 & w35661) | (w13288 & w35662) | (w35661 & w35662);
assign w15803 = ~w15801 & ~w15802;
assign w15804 = w15794 & ~w15803;
assign w15805 = (~w15792 & ~w15794) | (~w15792 & w35663) | (~w15794 & w35663);
assign w15806 = ~w15705 & ~w15714;
assign w15807 = ~w15715 & ~w15806;
assign w15808 = w15805 & w15807;
assign w15809 = ~w15715 & ~w15808;
assign w15810 = ~w15658 & ~w15667;
assign w15811 = ~w15668 & ~w15810;
assign w15812 = ~w15809 & w15811;
assign w15813 = w15809 & ~w15811;
assign w15814 = ~w15812 & ~w15813;
assign w15815 = w6996 & w13177;
assign w15816 = ~w13174 & w35664;
assign w15817 = ~w13011 & w35665;
assign w15818 = ~w15816 & ~w15817;
assign w15819 = ~w15815 & w15818;
assign w15820 = (w15819 & ~w13207) | (w15819 & w35666) | (~w13207 & w35666);
assign w15821 = a_14 & ~w15820;
assign w15822 = (~w13207 & w35667) | (~w13207 & w35668) | (w35667 & w35668);
assign w15823 = ~w15821 & ~w15822;
assign w15824 = w15814 & w15823;
assign w15825 = (~w15812 & ~w15814) | (~w15812 & w35669) | (~w15814 & w35669);
assign w15826 = w13948 & ~w15825;
assign w15827 = ~w13948 & w15825;
assign w15828 = ~w15826 & ~w15827;
assign w15829 = ~w15674 & ~w15683;
assign w15830 = ~w15684 & ~w15829;
assign w15831 = w15828 & w15830;
assign w15832 = (~w15826 & ~w15828) | (~w15826 & w35670) | (~w15828 & w35670);
assign w15833 = ~w15695 & ~w15697;
assign w15834 = ~w15698 & ~w15833;
assign w15835 = w15832 & ~w15834;
assign w15836 = w15699 & ~w15701;
assign w15837 = ~w15702 & ~w15836;
assign w15838 = ~w15835 & w15837;
assign w15839 = w15703 & ~w15838;
assign w15840 = w15556 & ~w15565;
assign w15841 = ~w15558 & ~w15563;
assign w15842 = ~w14838 & ~w14840;
assign w15843 = ~w14841 & ~w15842;
assign w15844 = ~w15841 & w15843;
assign w15845 = w15841 & ~w15843;
assign w15846 = ~w15844 & ~w15845;
assign w15847 = ~w15840 & w15846;
assign w15848 = ~w15839 & w15847;
assign w15849 = ~w15787 & ~w15789;
assign w15850 = ~w15790 & ~w15849;
assign w15851 = ~w15748 & w15764;
assign w15852 = ~w15765 & ~w15851;
assign w15853 = w15450 & ~w15452;
assign w15854 = ~w15453 & ~w15853;
assign w15855 = w4638 & ~w12630;
assign w15856 = ~w518 & ~w12668;
assign w15857 = w4666 & w12622;
assign w15858 = ~w15855 & ~w15856;
assign w15859 = ~w15857 & w15858;
assign w15860 = (w15859 & w14412) | (w15859 & w35671) | (w14412 & w35671);
assign w15861 = a_26 & ~w15860;
assign w15862 = (w14412 & w35672) | (w14412 & w35673) | (w35672 & w35673);
assign w15863 = ~w15861 & ~w15862;
assign w15864 = w15854 & ~w15863;
assign w15865 = ~w15854 & w15863;
assign w15866 = ~w15864 & ~w15865;
assign w15867 = w15446 & ~w15448;
assign w15868 = ~w15449 & ~w15867;
assign w15869 = w4070 & ~w15027;
assign w15870 = w3957 & w12651;
assign w15871 = w4446 & ~w12637;
assign w15872 = w4068 & w12646;
assign w15873 = ~w15871 & w35674;
assign w15874 = ~w15869 & w35675;
assign w15875 = (a_29 & w15869) | (a_29 & w35676) | (w15869 & w35676);
assign w15876 = ~w15874 & ~w15875;
assign w15877 = w15868 & ~w15876;
assign w15878 = w4446 & w12646;
assign w15879 = w4068 & w12651;
assign w15880 = ~w15044 & w35677;
assign w15881 = (~w15878 & w12830) | (~w15878 & w35678) | (w12830 & w35678);
assign w15882 = ~w15879 & w15881;
assign w15883 = ~w15880 & w35679;
assign w15884 = (a_29 & w15880) | (a_29 & w35680) | (w15880 & w35680);
assign w15885 = ~w15883 & ~w15884;
assign w15886 = ~w15120 & ~w15444;
assign w15887 = ~w15443 & w35681;
assign w15888 = (w15886 & w15443) | (w15886 & w35682) | (w15443 & w35682);
assign w15889 = ~w15887 & ~w15888;
assign w15890 = ~w15885 & ~w15889;
assign w15891 = ~w15148 & ~w15442;
assign w15892 = ~w15443 & ~w15891;
assign w15893 = w4446 & w12651;
assign w15894 = w3957 & w12793;
assign w15895 = w4068 & ~w12830;
assign w15896 = ~w15893 & ~w15894;
assign w15897 = (a_29 & w15895) | (a_29 & w35683) | (w15895 & w35683);
assign w15898 = w4070 & w14614;
assign w15899 = ~w15895 & w35684;
assign w15900 = ~w15898 & w15899;
assign w15901 = (~w15897 & ~w14614) | (~w15897 & w35685) | (~w14614 & w35685);
assign w15902 = ~w15900 & w15901;
assign w15903 = ~w15892 & ~w15902;
assign w15904 = w4070 & w15099;
assign w15905 = w4070 & w15098;
assign w15906 = w4068 & w12789;
assign w15907 = ~w12770 & w35686;
assign w15908 = w4446 & w12793;
assign w15909 = ~w15906 & ~w15907;
assign w15910 = ~w15908 & w15909;
assign w15911 = (w15910 & ~w15067) | (w15910 & w35687) | (~w15067 & w35687);
assign w15912 = ~w15904 & w15911;
assign w15913 = a_29 & w15912;
assign w15914 = ~a_29 & ~w15912;
assign w15915 = ~w15913 & ~w15914;
assign w15916 = ~w15199 & ~w15413;
assign w15917 = w15411 & ~w15916;
assign w15918 = ~w15411 & w15916;
assign w15919 = ~w15917 & ~w15918;
assign w15920 = ~w15915 & w15919;
assign w15921 = w4446 & w12789;
assign w15922 = (w4068 & w11977) | (w4068 & w31800) | (w11977 & w31800);
assign w15923 = ~w12770 & w15922;
assign w15924 = w3957 & ~w12733;
assign w15925 = ~w12749 & w15924;
assign w15926 = ~w12748 & w31801;
assign w15927 = ~w15925 & ~w15926;
assign w15928 = ~w15923 & w15927;
assign w15929 = ~w15921 & w15928;
assign w15930 = ~w15121 & w15929;
assign w15931 = (w4070 & w12740) | (w4070 & w31802) | (w12740 & w31802);
assign w15932 = (w15931 & ~w12717) | (w15931 & w31803) | (~w12717 & w31803);
assign w15933 = w4070 & ~w12760;
assign w15934 = w15929 & ~w15933;
assign w15935 = ~w15932 & w15934;
assign w15936 = ~w15930 & ~w15935;
assign w15937 = w4070 & w15127;
assign w15938 = ~w15936 & ~w15937;
assign w15939 = ~a_29 & w15938;
assign w15940 = a_29 & ~w15938;
assign w15941 = ~w15939 & ~w15940;
assign w15942 = ~w15241 & ~w15242;
assign w15943 = w15410 & ~w15942;
assign w15944 = ~w15410 & w15942;
assign w15945 = ~w15943 & ~w15944;
assign w15946 = w15941 & w15945;
assign w15947 = w4070 & ~w15154;
assign w15948 = w15150 & w15931;
assign w15949 = ~w12729 & w15948;
assign w15950 = w4446 & ~w12774;
assign w15951 = w4068 & w12732;
assign w15952 = w3957 & w12739;
assign w15953 = ~w15951 & ~w15952;
assign w15954 = ~w15950 & w15953;
assign w15955 = (w15954 & w12729) | (w15954 & w31804) | (w12729 & w31804);
assign w15956 = ~w15947 & w15955;
assign w15957 = a_29 & ~w15956;
assign w15958 = ~a_29 & w15954;
assign w15959 = ~w15949 & w15958;
assign w15960 = ~w15947 & w15959;
assign w15961 = ~w15318 & ~w15403;
assign w15962 = w15402 & ~w15961;
assign w15963 = ~w15318 & w15404;
assign w15964 = ~w15962 & ~w15963;
assign w15965 = ~w15960 & w15964;
assign w15966 = ~w15957 & w15965;
assign w15967 = w15960 & ~w15964;
assign w15968 = a_29 & ~w15964;
assign w15969 = ~w15956 & w15968;
assign w15970 = ~w15967 & ~w15969;
assign w15971 = ~w15966 & w15970;
assign w15972 = w4446 & w12732;
assign w15973 = w3957 & w12701;
assign w15974 = (~w15973 & ~w12739) | (~w15973 & w31805) | (~w12739 & w31805);
assign w15975 = ~w15972 & w15974;
assign w15976 = w12717 & ~w12728;
assign w15977 = ~w15203 & ~w15976;
assign w15978 = ~a_29 & w15975;
assign w15979 = w15977 & w15978;
assign w15980 = w7268 & ~w12728;
assign w15981 = w12717 & w15980;
assign w15982 = w7268 & w12728;
assign w15983 = ~w12717 & w15982;
assign w15984 = w7269 & w15975;
assign w15985 = a_29 & ~w15975;
assign w15986 = ~w15981 & ~w15983;
assign w15987 = ~w15984 & ~w15985;
assign w15988 = w15986 & w15987;
assign w15989 = ~w15979 & w15988;
assign w15990 = w15383 & w15399;
assign w15991 = ~w15400 & ~w15990;
assign w15992 = ~w15989 & ~w15991;
assign w15993 = ~w15330 & w15375;
assign w15994 = ~w15378 & ~w15993;
assign w15995 = ~w1477 & w12679;
assign w15996 = w12702 & w31806;
assign w15997 = w4070 & w15385;
assign w15998 = ~w12702 & w15997;
assign w15999 = w3957 & w12679;
assign w16000 = w4446 & w11683;
assign w16001 = w11678 & w16000;
assign w16002 = w4446 & ~w12675;
assign w16003 = ~w12674 & w16002;
assign w16004 = w4068 & ~w11501;
assign w16005 = w12684 & w16004;
assign w16006 = ~w15999 & ~w16001;
assign w16007 = ~w16003 & ~w16005;
assign w16008 = w16006 & w16007;
assign w16009 = ~w15998 & w16008;
assign w16010 = ~w15996 & w16009;
assign w16011 = w3954 & w12679;
assign w16012 = w4068 & w12679;
assign w16013 = w12684 & w35688;
assign w16014 = (~w16012 & w15324) | (~w16012 & w31807) | (w15324 & w31807);
assign w16015 = (a_29 & ~w12679) | (a_29 & w35689) | (~w12679 & w35689);
assign w16016 = w16014 & w35690;
assign w16017 = w16010 & w31808;
assign w16018 = (~w15995 & ~w16010) | (~w15995 & w31809) | (~w16010 & w31809);
assign w16019 = ~w16017 & ~w16018;
assign w16020 = w4070 & w15283;
assign w16021 = w4070 & ~w12681;
assign w16022 = w12688 & w16021;
assign w16023 = ~w15282 & w16022;
assign w16024 = w4446 & ~w11825;
assign w16025 = ~w12699 & w16024;
assign w16026 = w11825 & w16000;
assign w16027 = ~w11678 & w16026;
assign w16028 = w15293 & w16004;
assign w16029 = ~w12674 & w31810;
assign w16030 = w12684 & w31811;
assign w16031 = ~w16027 & ~w16028;
assign w16032 = ~w16025 & w16031;
assign w16033 = ~w16029 & ~w16030;
assign w16034 = w16032 & w16033;
assign w16035 = ~w16023 & w16034;
assign w16036 = ~w16020 & w16035;
assign w16037 = a_29 & ~w16036;
assign w16038 = ~a_29 & w16036;
assign w16039 = ~w16037 & ~w16038;
assign w16040 = w16019 & w16039;
assign w16041 = (~w16017 & ~w16039) | (~w16017 & w31812) | (~w16039 & w31812);
assign w16042 = ~w15994 & ~w16041;
assign w16043 = w15994 & ~w16017;
assign w16044 = (w16043 & ~w16039) | (w16043 & w31813) | (~w16039 & w31813);
assign w16045 = w7268 & ~w15278;
assign w16046 = w4446 & w12739;
assign w16047 = w3957 & w12702;
assign w16048 = w4068 & w12701;
assign w16049 = ~w16047 & ~w16048;
assign w16050 = ~w16046 & w31814;
assign w16051 = (a_29 & w16046) | (a_29 & w31815) | (w16046 & w31815);
assign w16052 = ~w16046 & w35691;
assign w16053 = w15278 & w16052;
assign w16054 = ~w16050 & ~w16051;
assign w16055 = ~w16045 & w16054;
assign w16056 = ~w16053 & w16055;
assign w16057 = ~w16044 & w16056;
assign w16058 = ~w16042 & ~w16057;
assign w16059 = w15989 & w15991;
assign w16060 = w16058 & ~w16059;
assign w16061 = ~w15992 & ~w16060;
assign w16062 = w15971 & w16061;
assign w16063 = ~w15932 & ~w15933;
assign w16064 = w15434 & ~w16063;
assign w16065 = ~w12770 & w35692;
assign w16066 = w3957 & w12732;
assign w16067 = w4068 & ~w12774;
assign w16068 = ~w16065 & ~w16066;
assign w16069 = ~w16067 & w16068;
assign w16070 = (a_29 & w16064) | (a_29 & w35693) | (w16064 & w35693);
assign w16071 = ~a_29 & w16069;
assign w16072 = ~w16064 & w16071;
assign w16073 = w15280 & ~w15408;
assign w16074 = w15405 & ~w16073;
assign w16075 = w15280 & w15409;
assign w16076 = ~w16074 & ~w16075;
assign w16077 = w16076 & w16080;
assign w16078 = ~w15966 & ~w16077;
assign w16079 = ~w16062 & w16078;
assign w16080 = ~w16070 & ~w16072;
assign w16081 = ~w16076 & ~w16080;
assign w16082 = ~w15941 & ~w15945;
assign w16083 = (~w16081 & w15941) | (~w16081 & w35694) | (w15941 & w35694);
assign w16084 = (~w15946 & w16079) | (~w15946 & w35695) | (w16079 & w35695);
assign w16085 = w15915 & ~w15919;
assign w16086 = ~w15920 & ~w16085;
assign w16087 = ~w16084 & w16086;
assign w16088 = (~w15920 & w16084) | (~w15920 & w31816) | (w16084 & w31816);
assign w16089 = w15437 & ~w15441;
assign w16090 = (~w15413 & w15411) | (~w15413 & w35696) | (w15411 & w35696);
assign w16091 = ~w16089 & w16090;
assign w16092 = w16089 & ~w16090;
assign w16093 = ~w16091 & ~w16092;
assign w16094 = w4068 & w12793;
assign w16095 = w3957 & w12789;
assign w16096 = w4446 & ~w12830;
assign w16097 = ~w16094 & ~w16095;
assign w16098 = (a_29 & w16096) | (a_29 & w35697) | (w16096 & w35697);
assign w16099 = ~w16096 & w35698;
assign w16100 = ~w16098 & ~w16099;
assign w16101 = ~w15071 & w16100;
assign w16102 = ~w16096 & w35699;
assign w16103 = ~w7268 & ~w16098;
assign w16104 = ~w16102 & w16103;
assign w16105 = w15071 & w16104;
assign w16106 = ~w16101 & ~w16105;
assign w16107 = ~w16093 & w16106;
assign w16108 = ~w16088 & ~w16107;
assign w16109 = w16093 & ~w16106;
assign w16110 = w15892 & w15902;
assign w16111 = ~w16109 & ~w16110;
assign w16112 = (~w15903 & w16108) | (~w15903 & w35700) | (w16108 & w35700);
assign w16113 = w15885 & w15889;
assign w16114 = ~w15890 & ~w16113;
assign w16115 = ~w16112 & w16114;
assign w16116 = (~w15890 & w16112) | (~w15890 & w35701) | (w16112 & w35701);
assign w16117 = ~w15868 & w15876;
assign w16118 = (~w15877 & w16116) | (~w15877 & w35702) | (w16116 & w35702);
assign w16119 = w15866 & ~w16118;
assign w16120 = (~w15864 & ~w15866) | (~w15864 & w35703) | (~w15866 & w35703);
assign w16121 = w15852 & w16120;
assign w16122 = ~w15852 & ~w16120;
assign w16123 = ~w16121 & ~w16122;
assign w16124 = w5286 & w12874;
assign w16125 = w5016 & ~w12860;
assign w16126 = w5080 & w12869;
assign w16127 = w5017 & w13965;
assign w16128 = ~w16125 & w35704;
assign w16129 = ~w16127 & w35705;
assign w16130 = (a_23 & w16127) | (a_23 & w35706) | (w16127 & w35706);
assign w16131 = ~w16129 & ~w16130;
assign w16132 = w16123 & w16131;
assign w16133 = (~w16121 & ~w16123) | (~w16121 & w35707) | (~w16123 & w35707);
assign w16134 = w8311 & w13815;
assign w16135 = ~w12892 & w35708;
assign w16136 = w5816 & ~w12910;
assign w16137 = ~w12905 & w35709;
assign w16138 = ~w16136 & w35710;
assign w16139 = a_20 & ~w16138;
assign w16140 = ~a_20 & w16138;
assign w16141 = (w16140 & ~w13815) | (w16140 & w35711) | (~w13815 & w35711);
assign w16142 = ~w16134 & ~w16139;
assign w16143 = ~w16141 & w16142;
assign w16144 = ~w16133 & w16143;
assign w16145 = w15779 & ~w15781;
assign w16146 = ~w15782 & ~w16145;
assign w16147 = w16133 & ~w16143;
assign w16148 = ~w16144 & ~w16147;
assign w16149 = ~w16146 & w16148;
assign w16150 = (~w16144 & ~w16148) | (~w16144 & w35712) | (~w16148 & w35712);
assign w16151 = ~w15738 & ~w15739;
assign w16152 = ~w12914 & w35713;
assign w16153 = w5818 & ~w12910;
assign w16154 = ~w12905 & w35714;
assign w16155 = (w5309 & w13518) | (w5309 & w35715) | (w13518 & w35715);
assign w16156 = ~w16153 & ~w16154;
assign w16157 = ~w16152 & w16156;
assign w16158 = (a_20 & w16155) | (a_20 & w35716) | (w16155 & w35716);
assign w16159 = ~w16155 & w35717;
assign w16160 = ~w16158 & ~w16159;
assign w16161 = ~w15782 & w35718;
assign w16162 = (w16160 & w15782) | (w16160 & w35719) | (w15782 & w35719);
assign w16163 = ~w16161 & ~w16162;
assign w16164 = w16151 & w16163;
assign w16165 = ~w16151 & ~w16163;
assign w16166 = ~w16164 & ~w16165;
assign w16167 = ~w16150 & ~w16166;
assign w16168 = w16160 & w16166;
assign w16169 = ~w16167 & ~w16168;
assign w16170 = ~w12589 & w35720;
assign w16171 = (w6059 & w12612) | (w6059 & w35721) | (w12612 & w35721);
assign w16172 = (w6061 & w12616) | (w6061 & w35722) | (w12616 & w35722);
assign w16173 = ~w16170 & ~w16171;
assign w16174 = ~w16172 & w16173;
assign w16175 = (w16174 & ~w13123) | (w16174 & w35723) | (~w13123 & w35723);
assign w16176 = a_17 & ~w16175;
assign w16177 = (~w13123 & w35724) | (~w13123 & w35725) | (w35724 & w35725);
assign w16178 = ~w16176 & ~w16177;
assign w16179 = ~w16169 & w16178;
assign w16180 = w16169 & ~w16178;
assign w16181 = ~w16179 & ~w16180;
assign w16182 = w15850 & w16181;
assign w16183 = ~w15850 & ~w16181;
assign w16184 = ~w16182 & ~w16183;
assign w16185 = w6998 & w12601;
assign w16186 = w6446 & w12604;
assign w16187 = w6996 & w12598;
assign w16188 = ~w16185 & ~w16186;
assign w16189 = (a_14 & ~w16188) | (a_14 & w35726) | (~w16188 & w35726);
assign w16190 = w8592 & w12961;
assign w16191 = w16188 & w35727;
assign w16192 = ~w16190 & w16191;
assign w16193 = (~w16189 & ~w12961) | (~w16189 & w35728) | (~w12961 & w35728);
assign w16194 = ~w16192 & w16193;
assign w16195 = w16150 & w16166;
assign w16196 = ~w16167 & ~w16195;
assign w16197 = (w6304 & w12616) | (w6304 & w35729) | (w12616 & w35729);
assign w16198 = (w6061 & w12612) | (w6061 & w35730) | (w12612 & w35730);
assign w16199 = ~w12930 & w35731;
assign w16200 = ~w16198 & ~w16199;
assign w16201 = ~w16197 & w16200;
assign w16202 = (w16201 & ~w13389) | (w16201 & w35732) | (~w13389 & w35732);
assign w16203 = a_17 & w16202;
assign w16204 = (w13389 & w35733) | (w13389 & w35734) | (w35733 & w35734);
assign w16205 = ~w16203 & ~w16204;
assign w16206 = ~w16196 & w16205;
assign w16207 = w16196 & ~w16205;
assign w16208 = w16146 & ~w16148;
assign w16209 = ~w16149 & ~w16208;
assign w16210 = (w6304 & w12612) | (w6304 & w35735) | (w12612 & w35735);
assign w16211 = ~w12914 & w35736;
assign w16212 = ~w12930 & w35737;
assign w16213 = ~w16211 & ~w16212;
assign w16214 = ~w16210 & w16213;
assign w16215 = (w16214 & ~w13375) | (w16214 & w35738) | (~w13375 & w35738);
assign w16216 = a_17 & ~w16215;
assign w16217 = (~w13375 & w35739) | (~w13375 & w35740) | (w35739 & w35740);
assign w16218 = ~w16216 & ~w16217;
assign w16219 = ~w16209 & ~w16218;
assign w16220 = ~w16123 & ~w16131;
assign w16221 = ~w16132 & ~w16220;
assign w16222 = ~w12905 & w35741;
assign w16223 = ~w12892 & w35742;
assign w16224 = w5308 & ~w12878;
assign w16225 = ~w13598 & w35743;
assign w16226 = ~w16223 & ~w16224;
assign w16227 = ~w16222 & w16226;
assign w16228 = ~w16225 & w35744;
assign w16229 = (a_20 & w16225) | (a_20 & w35745) | (w16225 & w35745);
assign w16230 = ~w16228 & ~w16229;
assign w16231 = ~w16221 & ~w16230;
assign w16232 = w16221 & w16230;
assign w16233 = ~w16231 & ~w16232;
assign w16234 = ~w15866 & w16118;
assign w16235 = ~w16119 & ~w16234;
assign w16236 = w16112 & ~w16114;
assign w16237 = ~w16115 & ~w16236;
assign w16238 = w4666 & ~w12668;
assign w16239 = ~w518 & ~w12637;
assign w16240 = w4638 & ~w12661;
assign w16241 = ~w16239 & ~w16240;
assign w16242 = ~w16238 & w16241;
assign w16243 = (w16242 & ~w14393) | (w16242 & w35746) | (~w14393 & w35746);
assign w16244 = ~a_26 & w16243;
assign w16245 = (w14393 & w35747) | (w14393 & w35748) | (w35747 & w35748);
assign w16246 = ~w16244 & ~w16245;
assign w16247 = w16237 & ~w16246;
assign w16248 = ~w16237 & w16246;
assign w16249 = ~w518 & w12646;
assign w16250 = w4638 & ~w12637;
assign w16251 = w4666 & ~w12661;
assign w16252 = ~w16249 & ~w16250;
assign w16253 = ~w16251 & w16252;
assign w16254 = (~w31817 & w35749) | (~w31817 & w35750) | (w35749 & w35750);
assign w16255 = a_26 & ~w16254;
assign w16256 = ~a_26 & w16254;
assign w16257 = ~w16255 & ~w16256;
assign w16258 = (~w16109 & w16088) | (~w16109 & w35751) | (w16088 & w35751);
assign w16259 = ~w15903 & ~w16110;
assign w16260 = w16257 & ~w16259;
assign w16261 = ~w16257 & w16259;
assign w16262 = ~w16260 & ~w16261;
assign w16263 = w16258 & w16262;
assign w16264 = ~w16258 & ~w16262;
assign w16265 = ~w16263 & ~w16264;
assign w16266 = ~w16257 & ~w16265;
assign w16267 = w4666 & w12651;
assign w16268 = ~w518 & w12793;
assign w16269 = w4638 & ~w12830;
assign w16270 = ~w16267 & ~w16268;
assign w16271 = ~w16269 & w16270;
assign w16272 = (~w14614 & w35752) | (~w14614 & w35753) | (w35752 & w35753);
assign w16273 = (w14614 & w35754) | (w14614 & w35755) | (w35754 & w35755);
assign w16274 = ~w16272 & ~w16273;
assign w16275 = ~w15946 & ~w16082;
assign w16276 = (~w16081 & w16062) | (~w16081 & w35756) | (w16062 & w35756);
assign w16277 = w16275 & ~w16276;
assign w16278 = ~w16275 & w16276;
assign w16279 = ~w16277 & ~w16278;
assign w16280 = ~w16274 & w16279;
assign w16281 = ~w15971 & ~w16061;
assign w16282 = ~w16062 & ~w16281;
assign w16283 = w1226 & w15099;
assign w16284 = w1226 & w15098;
assign w16285 = ~w12770 & w35757;
assign w16286 = w4638 & w12789;
assign w16287 = w4666 & w12793;
assign w16288 = ~w16285 & ~w16286;
assign w16289 = ~w16287 & w16288;
assign w16290 = (w16289 & ~w15067) | (w16289 & w35758) | (~w15067 & w35758);
assign w16291 = ~w16283 & w16290;
assign w16292 = a_26 & ~w16291;
assign w16293 = ~a_26 & w16291;
assign w16294 = ~w16292 & ~w16293;
assign w16295 = w16282 & w16294;
assign w16296 = (w1226 & w12740) | (w1226 & w35759) | (w12740 & w35759);
assign w16297 = w1226 & ~w12760;
assign w16298 = (~w16297 & w12729) | (~w16297 & w31819) | (w12729 & w31819);
assign w16299 = w15434 & ~w16298;
assign w16300 = ~w12770 & w35760;
assign w16301 = ~w518 & w12732;
assign w16302 = w4638 & ~w12774;
assign w16303 = ~w16300 & ~w16301;
assign w16304 = ~w16302 & w16303;
assign w16305 = (a_26 & w16299) | (a_26 & w35761) | (w16299 & w35761);
assign w16306 = ~w16299 & w35762;
assign w16307 = ~w16305 & ~w16306;
assign w16308 = ~w16042 & ~w16044;
assign w16309 = ~w16056 & w16308;
assign w16310 = w16056 & ~w16308;
assign w16311 = ~w16309 & ~w16310;
assign w16312 = w16307 & ~w16311;
assign w16313 = ~w16307 & w16311;
assign w16314 = ~w16312 & ~w16313;
assign w16315 = w4666 & w12732;
assign w16316 = ~w518 & w12701;
assign w16317 = (~w16316 & ~w12739) | (~w16316 & w31820) | (~w12739 & w31820);
assign w16318 = ~w16315 & w16317;
assign w16319 = ~a_26 & w16318;
assign w16320 = w15977 & w16319;
assign w16321 = w4403 & ~w12728;
assign w16322 = w12717 & w16321;
assign w16323 = w4403 & w12728;
assign w16324 = ~w12717 & w16323;
assign w16325 = w7680 & w16318;
assign w16326 = a_26 & ~w16318;
assign w16327 = ~w16322 & ~w16324;
assign w16328 = ~w16325 & ~w16326;
assign w16329 = w16327 & w16328;
assign w16330 = ~w16320 & w16329;
assign w16331 = w12679 & w35763;
assign w16332 = w16014 & w35764;
assign w16333 = a_29 & ~w16332;
assign w16334 = ~w16010 & w16333;
assign w16335 = w16010 & ~w16333;
assign w16336 = ~w16334 & ~w16335;
assign w16337 = ~w16330 & ~w16336;
assign w16338 = (w16331 & ~w16014) | (w16331 & w35765) | (~w16014 & w35765);
assign w16339 = ~w16332 & ~w16338;
assign w16340 = w1226 & w15283;
assign w16341 = w1226 & ~w12681;
assign w16342 = w12688 & w16341;
assign w16343 = ~w15282 & w16342;
assign w16344 = w4666 & ~w11825;
assign w16345 = ~w12699 & w16344;
assign w16346 = w4666 & w11683;
assign w16347 = w11825 & w16346;
assign w16348 = ~w11678 & w16347;
assign w16349 = w4638 & ~w11501;
assign w16350 = w15293 & w16349;
assign w16351 = w12684 & w31821;
assign w16352 = ~w12674 & w31822;
assign w16353 = ~w16348 & ~w16350;
assign w16354 = ~w16345 & w16353;
assign w16355 = ~w16351 & ~w16352;
assign w16356 = w16354 & w16355;
assign w16357 = ~w16343 & w16356;
assign w16358 = ~w16340 & w16357;
assign w16359 = a_26 & ~w16358;
assign w16360 = ~a_26 & w16358;
assign w16361 = ~w16359 & ~w16360;
assign w16362 = w12702 & w31823;
assign w16363 = w1226 & w15385;
assign w16364 = ~w12702 & w16363;
assign w16365 = ~w518 & w12679;
assign w16366 = w4666 & ~w12675;
assign w16367 = ~w12674 & w16366;
assign w16368 = w11678 & w16346;
assign w16369 = w12684 & w16349;
assign w16370 = ~w16365 & ~w16367;
assign w16371 = ~w16368 & ~w16369;
assign w16372 = w16370 & w16371;
assign w16373 = ~w16364 & w16372;
assign w16374 = ~w16362 & w16373;
assign w16375 = w1226 & w12679;
assign w16376 = ~w12685 & ~w16375;
assign w16377 = w12684 & w31824;
assign w16378 = ~w16376 & ~w16377;
assign w16379 = ~w1222 & w12679;
assign w16380 = w12679 & w35766;
assign w16381 = w4638 & w12679;
assign w16382 = ~w16363 & w35767;
assign w16383 = ~w16378 & w16382;
assign w16384 = ~w16378 & w35768;
assign w16385 = (~w16011 & ~w16374) | (~w16011 & w35769) | (~w16374 & w35769);
assign w16386 = (~w16339 & ~w16361) | (~w16339 & w31825) | (~w16361 & w31825);
assign w16387 = w16361 & w31826;
assign w16388 = w4403 & ~w15278;
assign w16389 = w4666 & w12739;
assign w16390 = w4638 & w12701;
assign w16391 = ~w518 & w12702;
assign w16392 = ~w16390 & ~w16391;
assign w16393 = ~w16389 & w31827;
assign w16394 = (a_26 & w16389) | (a_26 & w31828) | (w16389 & w31828);
assign w16395 = ~w16389 & w35770;
assign w16396 = w15278 & w16395;
assign w16397 = ~w16393 & ~w16394;
assign w16398 = ~w16388 & w16397;
assign w16399 = ~w16396 & w16398;
assign w16400 = (~w16386 & w16399) | (~w16386 & w31829) | (w16399 & w31829);
assign w16401 = w16330 & w16336;
assign w16402 = ~w16400 & ~w16401;
assign w16403 = ~w16337 & ~w16402;
assign w16404 = w4638 & w12732;
assign w16405 = ~w518 & w12739;
assign w16406 = w4666 & ~w12774;
assign w16407 = ~w16404 & ~w16405;
assign w16408 = ~w16406 & w16407;
assign w16409 = (w16408 & w15157) | (w16408 & w35771) | (w15157 & w35771);
assign w16410 = ~w16019 & ~w16039;
assign w16411 = ~w16040 & ~w16410;
assign w16412 = a_26 & ~w16411;
assign w16413 = ~a_26 & w16411;
assign w16414 = ~w16412 & ~w16413;
assign w16415 = w16409 & w16414;
assign w16416 = ~w16409 & ~w16414;
assign w16417 = ~w16415 & ~w16416;
assign w16418 = w16403 & w16417;
assign w16419 = w16411 & ~w16417;
assign w16420 = ~w16418 & ~w16419;
assign w16421 = w16314 & ~w16420;
assign w16422 = w15121 & ~w16298;
assign w16423 = w1226 & w15127;
assign w16424 = w4666 & w12789;
assign w16425 = ~w518 & ~w12774;
assign w16426 = ~w12770 & w35772;
assign w16427 = ~w16424 & w35773;
assign w16428 = ~w16422 & w16427;
assign w16429 = ~w16423 & w16428;
assign w16430 = a_26 & ~w16429;
assign w16431 = ~a_26 & w16429;
assign w16432 = ~w16430 & ~w16431;
assign w16433 = ~w15992 & ~w16059;
assign w16434 = w16058 & ~w16433;
assign w16435 = ~w16058 & w16433;
assign w16436 = ~w16434 & ~w16435;
assign w16437 = w16432 & w16436;
assign w16438 = (~w16312 & ~w16436) | (~w16312 & w31830) | (~w16436 & w31830);
assign w16439 = ~w16421 & w16438;
assign w16440 = ~w16432 & ~w16436;
assign w16441 = ~w16282 & ~w16294;
assign w16442 = ~w16440 & ~w16441;
assign w16443 = ~w16439 & w16442;
assign w16444 = ~w16295 & ~w16443;
assign w16445 = ~w16077 & ~w16081;
assign w16446 = ~w16062 & w35774;
assign w16447 = (w16445 & w16062) | (w16445 & w35775) | (w16062 & w35775);
assign w16448 = ~w16446 & ~w16447;
assign w16449 = w4638 & w12793;
assign w16450 = ~w518 & w12789;
assign w16451 = w4666 & ~w12830;
assign w16452 = ~w16449 & ~w16450;
assign w16453 = ~w16451 & w35776;
assign w16454 = w4403 & w15071;
assign w16455 = ~w16451 & w35777;
assign w16456 = (a_26 & w16451) | (a_26 & w35778) | (w16451 & w35778);
assign w16457 = ~w16455 & ~w16456;
assign w16458 = (w16457 & w15071) | (w16457 & w35779) | (w15071 & w35779);
assign w16459 = ~w16454 & w16458;
assign w16460 = w16448 & w16459;
assign w16461 = ~w16448 & ~w16459;
assign w16462 = ~w16460 & ~w16461;
assign w16463 = ~w16444 & w16462;
assign w16464 = w16274 & ~w16279;
assign w16465 = ~w16460 & ~w16464;
assign w16466 = ~w16463 & w16465;
assign w16467 = (~w16280 & w16463) | (~w16280 & w35780) | (w16463 & w35780);
assign w16468 = w16084 & ~w16086;
assign w16469 = ~w16087 & ~w16468;
assign w16470 = w4666 & w12646;
assign w16471 = w4638 & w12651;
assign w16472 = ~w518 & ~w12830;
assign w16473 = ~w15044 & w35781;
assign w16474 = ~w16470 & ~w16471;
assign w16475 = ~w16472 & w16474;
assign w16476 = ~w16473 & w35782;
assign w16477 = (a_26 & w16473) | (a_26 & w35783) | (w16473 & w35783);
assign w16478 = ~w16476 & ~w16477;
assign w16479 = w16469 & w16478;
assign w16480 = ~w16469 & ~w16478;
assign w16481 = ~w16479 & ~w16480;
assign w16482 = ~w16107 & ~w16109;
assign w16483 = w4666 & ~w12637;
assign w16484 = ~w518 & w12651;
assign w16485 = w4638 & w12646;
assign w16486 = ~w16483 & w35784;
assign w16487 = a_26 & ~w16486;
assign w16488 = ~a_26 & w16486;
assign w16489 = ~w16487 & ~w16488;
assign w16490 = w15027 & w16489;
assign w16491 = w7680 & w16486;
assign w16492 = (~w4403 & w16486) | (~w4403 & w32424) | (w16486 & w32424);
assign w16493 = ~w16491 & w16492;
assign w16494 = ~w15027 & w16493;
assign w16495 = ~w16490 & ~w16494;
assign w16496 = ~w16482 & w16495;
assign w16497 = w16088 & w16496;
assign w16498 = w16482 & w16495;
assign w16499 = ~w16088 & w16498;
assign w16500 = ~w16497 & ~w16499;
assign w16501 = w16481 & w16500;
assign w16502 = w16467 & w16501;
assign w16503 = w16482 & ~w16495;
assign w16504 = w16088 & w16503;
assign w16505 = ~w16482 & ~w16495;
assign w16506 = ~w16088 & w16505;
assign w16507 = ~w16504 & ~w16506;
assign w16508 = ~w16479 & w16507;
assign w16509 = w16500 & ~w16508;
assign w16510 = ~w16502 & ~w16509;
assign w16511 = ~w16502 & w31831;
assign w16512 = ~w16266 & ~w16511;
assign w16513 = (~w16248 & w16511) | (~w16248 & w35785) | (w16511 & w35785);
assign w16514 = ~w16247 & ~w16513;
assign w16515 = ~w15877 & ~w16117;
assign w16516 = w4638 & ~w12668;
assign w16517 = ~w518 & ~w12661;
assign w16518 = w4666 & ~w12630;
assign w16519 = ~w16516 & ~w16517;
assign w16520 = ~w16518 & w16519;
assign w16521 = (w16520 & w14535) | (w16520 & w35786) | (w14535 & w35786);
assign w16522 = ~a_26 & w16521;
assign w16523 = (~w14535 & w35787) | (~w14535 & w35788) | (w35787 & w35788);
assign w16524 = ~w16522 & ~w16523;
assign w16525 = w16515 & ~w16524;
assign w16526 = ~w16515 & w16524;
assign w16527 = ~w16525 & ~w16526;
assign w16528 = w16116 & w16527;
assign w16529 = ~w16116 & ~w16527;
assign w16530 = ~w16528 & ~w16529;
assign w16531 = (~w16530 & w16513) | (~w16530 & w35789) | (w16513 & w35789);
assign w16532 = ~w16524 & w16530;
assign w16533 = (w16235 & w16531) | (w16235 & w35790) | (w16531 & w35790);
assign w16534 = ~w16531 & w35791;
assign w16535 = w5016 & w12856;
assign w16536 = w5286 & w12869;
assign w16537 = (~w16535 & w12860) | (~w16535 & w35792) | (w12860 & w35792);
assign w16538 = ~w16536 & w16537;
assign w16539 = (w16538 & ~w13979) | (w16538 & w35793) | (~w13979 & w35793);
assign w16540 = a_23 & w16539;
assign w16541 = (w13979 & w35794) | (w13979 & w35795) | (w35794 & w35795);
assign w16542 = ~w16540 & ~w16541;
assign w16543 = ~w16534 & w16542;
assign w16544 = ~w16533 & ~w16543;
assign w16545 = w16233 & ~w16544;
assign w16546 = (~w16231 & ~w16233) | (~w16231 & w35796) | (~w16233 & w35796);
assign w16547 = w16209 & w16218;
assign w16548 = ~w16219 & ~w16547;
assign w16549 = ~w16546 & w16548;
assign w16550 = (~w16219 & ~w16548) | (~w16219 & w35797) | (~w16548 & w35797);
assign w16551 = ~w16207 & ~w16550;
assign w16552 = (~w16194 & w16551) | (~w16194 & w35798) | (w16551 & w35798);
assign w16553 = ~w16551 & w35799;
assign w16554 = ~w16552 & ~w16553;
assign w16555 = ~w16184 & w16554;
assign w16556 = w16184 & ~w16554;
assign w16557 = ~w16555 & ~w16556;
assign w16558 = w6996 & w12601;
assign w16559 = w6998 & w12604;
assign w16560 = ~w12589 & w35800;
assign w16561 = ~w16559 & ~w16560;
assign w16562 = ~w16558 & w16561;
assign w16563 = (w16562 & w13140) | (w16562 & w35801) | (w13140 & w35801);
assign w16564 = ~a_14 & w16563;
assign w16565 = (~w13140 & w35802) | (~w13140 & w35803) | (w35802 & w35803);
assign w16566 = ~w16564 & ~w16565;
assign w16567 = ~w16206 & ~w16207;
assign w16568 = w16550 & ~w16567;
assign w16569 = ~w16550 & w16567;
assign w16570 = ~w16568 & ~w16569;
assign w16571 = w16566 & ~w16570;
assign w16572 = ~w16566 & w16570;
assign w16573 = w16546 & ~w16548;
assign w16574 = ~w16549 & ~w16573;
assign w16575 = ~w16233 & w16544;
assign w16576 = ~w16545 & ~w16575;
assign w16577 = ~w16533 & ~w16534;
assign w16578 = ~w12892 & w35804;
assign w16579 = w5818 & ~w12878;
assign w16580 = w5308 & w12874;
assign w16581 = ~w16579 & ~w16580;
assign w16582 = ~w16578 & w16581;
assign w16583 = (w16582 & ~w13787) | (w16582 & w35805) | (~w13787 & w35805);
assign w16584 = a_20 & ~w16583;
assign w16585 = (~w13787 & w35806) | (~w13787 & w35807) | (w35806 & w35807);
assign w16586 = ~w16584 & ~w16585;
assign w16587 = w16542 & ~w16586;
assign w16588 = ~w16542 & w16586;
assign w16589 = ~w16587 & ~w16588;
assign w16590 = w16577 & w16589;
assign w16591 = ~w16577 & ~w16589;
assign w16592 = ~w16590 & ~w16591;
assign w16593 = w5080 & ~w12630;
assign w16594 = w5016 & ~w12668;
assign w16595 = w5286 & w12622;
assign w16596 = ~w16593 & ~w16594;
assign w16597 = ~w16595 & w16596;
assign w16598 = (w16597 & w14412) | (w16597 & w35808) | (w14412 & w35808);
assign w16599 = a_23 & ~w16598;
assign w16600 = (w14412 & w35809) | (w14412 & w35810) | (w35809 & w35810);
assign w16601 = ~w16599 & ~w16600;
assign w16602 = w16265 & w16601;
assign w16603 = w16510 & ~w16602;
assign w16604 = ~w16265 & w16601;
assign w16605 = ~w16510 & ~w16604;
assign w16606 = ~w16603 & ~w16605;
assign w16607 = w16265 & ~w16601;
assign w16608 = ~w16604 & ~w16607;
assign w16609 = w16510 & w16608;
assign w16610 = ~w16510 & ~w16608;
assign w16611 = ~w16609 & ~w16610;
assign w16612 = ~w16606 & ~w16611;
assign w16613 = ~w16314 & w16420;
assign w16614 = ~w16421 & ~w16613;
assign w16615 = w5080 & w12793;
assign w16616 = w5016 & w12789;
assign w16617 = w5286 & ~w12830;
assign w16618 = ~w16615 & ~w16616;
assign w16619 = ~w16617 & w35811;
assign w16620 = w7961 & w15071;
assign w16621 = ~w16617 & w35812;
assign w16622 = (a_23 & w16617) | (a_23 & w35813) | (w16617 & w35813);
assign w16623 = ~w16621 & ~w16622;
assign w16624 = (w16623 & w15071) | (w16623 & w35814) | (w15071 & w35814);
assign w16625 = ~w16620 & w16624;
assign w16626 = ~w16614 & ~w16625;
assign w16627 = ~w16403 & ~w16417;
assign w16628 = ~w16418 & ~w16627;
assign w16629 = w5017 & w15099;
assign w16630 = w5017 & w15098;
assign w16631 = ~w12770 & w35815;
assign w16632 = w5080 & w12789;
assign w16633 = w5286 & w12793;
assign w16634 = ~w16631 & ~w16632;
assign w16635 = ~w16633 & w16634;
assign w16636 = (w16635 & ~w15067) | (w16635 & w35816) | (~w15067 & w35816);
assign w16637 = ~w16629 & w16636;
assign w16638 = a_23 & w16637;
assign w16639 = ~a_23 & ~w16637;
assign w16640 = ~w16638 & ~w16639;
assign w16641 = ~w16628 & w16640;
assign w16642 = ~w16386 & ~w16387;
assign w16643 = w16399 & ~w16642;
assign w16644 = ~w16399 & w16642;
assign w16645 = ~w16643 & ~w16644;
assign w16646 = (w5017 & w12740) | (w5017 & w35817) | (w12740 & w35817);
assign w16647 = w5017 & ~w12760;
assign w16648 = (~w16647 & w12729) | (~w16647 & w31832) | (w12729 & w31832);
assign w16649 = w15434 & ~w16648;
assign w16650 = ~w12770 & w31833;
assign w16651 = w5016 & w12732;
assign w16652 = w5080 & ~w12774;
assign w16653 = ~w16650 & ~w16651;
assign w16654 = w16653 & w35818;
assign w16655 = (a_23 & ~w16653) | (a_23 & w35819) | (~w16653 & w35819);
assign w16656 = ~w16654 & ~w16655;
assign w16657 = ~w16649 & w16656;
assign w16658 = w16649 & ~w16656;
assign w16659 = ~w16657 & ~w16658;
assign w16660 = w16645 & w16659;
assign w16661 = (a_26 & w16378) | (a_26 & w35820) | (w16378 & w35820);
assign w16662 = ~w16374 & w16661;
assign w16663 = w16374 & ~w16661;
assign w16664 = ~w16662 & ~w16663;
assign w16665 = w5016 & w12701;
assign w16666 = w5286 & w12732;
assign w16667 = (~w16665 & ~w12739) | (~w16665 & w35821) | (~w12739 & w35821);
assign w16668 = ~w16666 & w16667;
assign w16669 = w16664 & w35822;
assign w16670 = w16664 & w31834;
assign w16671 = w16664 & w35823;
assign w16672 = (w16671 & w15977) | (w16671 & w37565) | (w15977 & w37565);
assign w16673 = (~w16669 & w15977) | (~w16669 & w35824) | (w15977 & w35824);
assign w16674 = ~w16672 & w16673;
assign w16675 = ~w16664 & w35825;
assign w16676 = (w16675 & w15977) | (w16675 & w37566) | (w15977 & w37566);
assign w16677 = w7961 & ~w16664;
assign w16678 = ~w16664 & w35826;
assign w16679 = (~w16678 & w15977) | (~w16678 & w37567) | (w15977 & w37567);
assign w16680 = ~w16676 & w16679;
assign w16681 = ~w16376 & w35827;
assign w16682 = ~w16383 & ~w16681;
assign w16683 = w12702 & w31835;
assign w16684 = w5017 & w15385;
assign w16685 = ~w12702 & w16684;
assign w16686 = w5286 & ~w12675;
assign w16687 = ~w12674 & w16686;
assign w16688 = w5016 & w12679;
assign w16689 = w5080 & ~w11501;
assign w16690 = w12684 & w16689;
assign w16691 = w5286 & w11683;
assign w16692 = w11678 & w16691;
assign w16693 = ~w16687 & ~w16688;
assign w16694 = ~w16690 & ~w16692;
assign w16695 = w16693 & w16694;
assign w16696 = ~w16685 & w16695;
assign w16697 = ~w16683 & w16696;
assign w16698 = w504 & w12679;
assign w16699 = w12684 & w31836;
assign w16700 = w5080 & w12679;
assign w16701 = w5017 & ~w15324;
assign w16702 = ~w16699 & ~w16700;
assign w16703 = ~w16701 & w16702;
assign w16704 = (a_23 & ~w12679) | (a_23 & w35828) | (~w12679 & w35828);
assign w16705 = w16703 & w16704;
assign w16706 = (~w16379 & ~w16697) | (~w16379 & w31837) | (~w16697 & w31837);
assign w16707 = w5017 & w15283;
assign w16708 = w5017 & ~w12681;
assign w16709 = w12688 & w16708;
assign w16710 = ~w15282 & w16709;
assign w16711 = w5286 & ~w11825;
assign w16712 = ~w12699 & w16711;
assign w16713 = w11825 & w16691;
assign w16714 = ~w11678 & w16713;
assign w16715 = w15293 & w16689;
assign w16716 = ~w12674 & w31838;
assign w16717 = w12684 & w31839;
assign w16718 = ~w16714 & ~w16715;
assign w16719 = ~w16712 & w16718;
assign w16720 = ~w16716 & ~w16717;
assign w16721 = w16719 & w16720;
assign w16722 = ~w16710 & w16721;
assign w16723 = ~w16707 & w16722;
assign w16724 = a_23 & ~w16723;
assign w16725 = ~a_23 & w16723;
assign w16726 = ~w16724 & ~w16725;
assign w16727 = (~w16682 & ~w16726) | (~w16682 & w31840) | (~w16726 & w31840);
assign w16728 = w5017 & w12715;
assign w16729 = w5286 & w12739;
assign w16730 = w5080 & w12701;
assign w16731 = w5016 & w12702;
assign w16732 = w5017 & ~w12700;
assign w16733 = w12711 & ~w16732;
assign w16734 = w5017 & w12700;
assign w16735 = ~w12711 & ~w16734;
assign w16736 = ~w16733 & ~w16735;
assign w16737 = ~w12704 & w16736;
assign w16738 = ~w16730 & ~w16731;
assign w16739 = ~w16729 & w16738;
assign w16740 = ~w16737 & w16739;
assign w16741 = ~w16728 & w16740;
assign w16742 = a_23 & ~w16741;
assign w16743 = ~a_23 & w16741;
assign w16744 = ~w16742 & ~w16743;
assign w16745 = w16726 & w31841;
assign w16746 = (~w16727 & w16744) | (~w16727 & w31842) | (w16744 & w31842);
assign w16747 = w16680 & w16746;
assign w16748 = w16674 & ~w16747;
assign w16749 = w5080 & w12732;
assign w16750 = w5016 & w12739;
assign w16751 = w5286 & ~w12774;
assign w16752 = ~w16749 & ~w16750;
assign w16753 = ~w16751 & w16752;
assign w16754 = (w16753 & w15157) | (w16753 & w35829) | (w15157 & w35829);
assign w16755 = w16374 & w37568;
assign w16756 = ~w16385 & ~w16755;
assign w16757 = w16361 & w16756;
assign w16758 = ~w16361 & ~w16756;
assign w16759 = ~w16757 & ~w16758;
assign w16760 = ~a_23 & w16759;
assign w16761 = a_23 & ~w16759;
assign w16762 = ~w16760 & ~w16761;
assign w16763 = w16754 & w16762;
assign w16764 = ~w16754 & ~w16762;
assign w16765 = ~w16763 & ~w16764;
assign w16766 = ~w16748 & w16765;
assign w16767 = ~w16754 & ~w16760;
assign w16768 = a_23 & w16759;
assign w16769 = w16754 & ~w16768;
assign w16770 = ~w16767 & ~w16769;
assign w16771 = ~w16645 & ~w16659;
assign w16772 = ~w16770 & ~w16771;
assign w16773 = (~w16660 & w16766) | (~w16660 & w31843) | (w16766 & w31843);
assign w16774 = w15121 & ~w16648;
assign w16775 = w5286 & w12789;
assign w16776 = w5016 & ~w12774;
assign w16777 = ~w12770 & w35830;
assign w16778 = ~w16775 & w35831;
assign w16779 = (w16778 & ~w15127) | (w16778 & w31844) | (~w15127 & w31844);
assign w16780 = (a_23 & ~w16779) | (a_23 & w35832) | (~w16779 & w35832);
assign w16781 = w16779 & w35833;
assign w16782 = ~w16780 & ~w16781;
assign w16783 = ~w16337 & ~w16401;
assign w16784 = w16400 & w16783;
assign w16785 = ~w16400 & ~w16783;
assign w16786 = ~w16784 & ~w16785;
assign w16787 = w16782 & w16786;
assign w16788 = ~w16782 & ~w16786;
assign w16789 = ~w16787 & ~w16788;
assign w16790 = w16773 & w16789;
assign w16791 = w16628 & ~w16640;
assign w16792 = ~w16787 & ~w16791;
assign w16793 = ~w16790 & w16792;
assign w16794 = ~w16641 & ~w16793;
assign w16795 = w16614 & w16625;
assign w16796 = ~w16626 & ~w16795;
assign w16797 = ~w16794 & w16796;
assign w16798 = ~w16626 & ~w16797;
assign w16799 = (~w16312 & w16420) | (~w16312 & w31845) | (w16420 & w31845);
assign w16800 = ~w16437 & ~w16440;
assign w16801 = w5286 & w12651;
assign w16802 = w5016 & w12793;
assign w16803 = w5080 & ~w12830;
assign w16804 = ~w16801 & ~w16802;
assign w16805 = ~w16803 & w35834;
assign w16806 = (a_23 & w16803) | (a_23 & w35835) | (w16803 & w35835);
assign w16807 = ~w16803 & w35836;
assign w16808 = ~w14614 & w16807;
assign w16809 = ~w16805 & ~w16806;
assign w16810 = (w16809 & ~w14614) | (w16809 & w31846) | (~w14614 & w31846);
assign w16811 = ~w16808 & w16810;
assign w16812 = w16800 & w16811;
assign w16813 = w16799 & w16812;
assign w16814 = ~w16800 & w16811;
assign w16815 = ~w16799 & w16814;
assign w16816 = ~w16813 & ~w16815;
assign w16817 = (~w16440 & w16421) | (~w16440 & w31847) | (w16421 & w31847);
assign w16818 = ~w16295 & ~w16441;
assign w16819 = ~w15044 & w35837;
assign w16820 = w5286 & w12646;
assign w16821 = w5080 & w12651;
assign w16822 = (~w16820 & w12830) | (~w16820 & w35838) | (w12830 & w35838);
assign w16823 = w16822 & w35839;
assign w16824 = (a_23 & ~w16822) | (a_23 & w35840) | (~w16822 & w35840);
assign w16825 = w16822 & w35841;
assign w16826 = ~w15045 & w16825;
assign w16827 = ~w16823 & ~w16824;
assign w16828 = ~w16819 & w16827;
assign w16829 = ~w16826 & w16828;
assign w16830 = ~w16818 & w16829;
assign w16831 = w16817 & w16830;
assign w16832 = w16818 & w16829;
assign w16833 = ~w16817 & w16832;
assign w16834 = ~w16831 & ~w16833;
assign w16835 = w16816 & w16834;
assign w16836 = ~w16798 & w16835;
assign w16837 = ~w16800 & ~w16811;
assign w16838 = w16799 & w16837;
assign w16839 = w16800 & ~w16811;
assign w16840 = ~w16799 & w16839;
assign w16841 = ~w16838 & ~w16840;
assign w16842 = w16818 & ~w16829;
assign w16843 = w16817 & w16842;
assign w16844 = ~w16818 & ~w16829;
assign w16845 = ~w16817 & w16844;
assign w16846 = ~w16843 & ~w16845;
assign w16847 = w16841 & w16846;
assign w16848 = w16834 & ~w16847;
assign w16849 = ~w16836 & ~w16848;
assign w16850 = w16444 & ~w16462;
assign w16851 = ~w16463 & ~w16850;
assign w16852 = w7961 & ~w15027;
assign w16853 = w5286 & ~w12637;
assign w16854 = w5016 & w12651;
assign w16855 = w5080 & w12646;
assign w16856 = ~w16853 & w35842;
assign w16857 = a_23 & ~w16856;
assign w16858 = ~a_23 & w16856;
assign w16859 = (w16858 & w15027) | (w16858 & w35843) | (w15027 & w35843);
assign w16860 = ~w16852 & ~w16857;
assign w16861 = ~w16859 & w16860;
assign w16862 = w16851 & w16861;
assign w16863 = ~w16849 & ~w16862;
assign w16864 = ~w16851 & ~w16861;
assign w16865 = (~w16460 & w16444) | (~w16460 & w35844) | (w16444 & w35844);
assign w16866 = w5080 & ~w12637;
assign w16867 = w5016 & w12646;
assign w16868 = w5286 & ~w12661;
assign w16869 = ~w16866 & ~w16867;
assign w16870 = (a_23 & ~w16869) | (a_23 & w35845) | (~w16869 & w35845);
assign w16871 = w16869 & w35846;
assign w16872 = ~w16870 & ~w16871;
assign w16873 = w14640 & w31848;
assign w16874 = w16869 & w35847;
assign w16875 = ~w7961 & ~w16870;
assign w16876 = ~w16874 & w16875;
assign w16877 = (w16876 & ~w14640) | (w16876 & w31849) | (~w14640 & w31849);
assign w16878 = ~w16873 & ~w16877;
assign w16879 = w16274 & ~w16878;
assign w16880 = ~w16274 & w16878;
assign w16881 = ~w16879 & ~w16880;
assign w16882 = w16279 & ~w16881;
assign w16883 = ~w16279 & w16881;
assign w16884 = ~w16882 & ~w16883;
assign w16885 = w16865 & w16884;
assign w16886 = ~w16865 & ~w16884;
assign w16887 = ~w16885 & ~w16886;
assign w16888 = ~w16864 & ~w16887;
assign w16889 = ~w16863 & w16888;
assign w16890 = ~w16878 & w16887;
assign w16891 = w5286 & ~w12668;
assign w16892 = w5016 & ~w12637;
assign w16893 = w5080 & ~w12661;
assign w16894 = ~w16892 & ~w16893;
assign w16895 = ~w16891 & w16894;
assign w16896 = (w16895 & ~w14393) | (w16895 & w35848) | (~w14393 & w35848);
assign w16897 = a_23 & w16896;
assign w16898 = (w14393 & w35849) | (w14393 & w35850) | (w35849 & w35850);
assign w16899 = ~w16897 & ~w16898;
assign w16900 = w16481 & ~w16899;
assign w16901 = ~w16467 & w16900;
assign w16902 = ~w16481 & ~w16899;
assign w16903 = w16467 & w16902;
assign w16904 = ~w16901 & ~w16903;
assign w16905 = ~w16890 & w16904;
assign w16906 = ~w16889 & w16905;
assign w16907 = ~w16280 & ~w16480;
assign w16908 = ~w16466 & w16907;
assign w16909 = (~w16479 & w16466) | (~w16479 & w35851) | (w16466 & w35851);
assign w16910 = w16500 & w16507;
assign w16911 = w5080 & ~w12668;
assign w16912 = w5016 & ~w12661;
assign w16913 = w5286 & ~w12630;
assign w16914 = ~w16911 & ~w16912;
assign w16915 = (a_23 & ~w16914) | (a_23 & w35852) | (~w16914 & w35852);
assign w16916 = w5017 & ~w14535;
assign w16917 = w16914 & w35853;
assign w16918 = ~w16916 & w16917;
assign w16919 = (~w16915 & w14535) | (~w16915 & w35854) | (w14535 & w35854);
assign w16920 = ~w16918 & w16919;
assign w16921 = ~w16908 & w35855;
assign w16922 = ~w16481 & w16899;
assign w16923 = ~w16467 & w16922;
assign w16924 = w16481 & w16899;
assign w16925 = w16467 & w16924;
assign w16926 = ~w16923 & ~w16925;
assign w16927 = w16910 & ~w16920;
assign w16928 = ~w16909 & w16927;
assign w16929 = w16926 & ~w16928;
assign w16930 = ~w16921 & w16929;
assign w16931 = ~w16906 & w16930;
assign w16932 = ~w16909 & w16910;
assign w16933 = (w16920 & w16908) | (w16920 & w35856) | (w16908 & w35856);
assign w16934 = ~w16932 & w16933;
assign w16935 = ~w16606 & ~w16934;
assign w16936 = (~w16612 & w16931) | (~w16612 & w35857) | (w16931 & w35857);
assign w16937 = w5016 & ~w12630;
assign w16938 = w5080 & w12622;
assign w16939 = w5286 & w12856;
assign w16940 = ~w16937 & ~w16938;
assign w16941 = ~w16939 & w16940;
assign w16942 = (w16941 & ~w14091) | (w16941 & w35858) | (~w14091 & w35858);
assign w16943 = ~a_23 & w16942;
assign w16944 = (w14091 & w35859) | (w14091 & w35860) | (w35859 & w35860);
assign w16945 = ~w16943 & ~w16944;
assign w16946 = w16246 & ~w16945;
assign w16947 = ~w16246 & w16945;
assign w16948 = ~w16946 & ~w16947;
assign w16949 = w16237 & ~w16948;
assign w16950 = ~w16237 & w16948;
assign w16951 = ~w16949 & ~w16950;
assign w16952 = w16512 & w16951;
assign w16953 = ~w16512 & ~w16951;
assign w16954 = ~w16952 & ~w16953;
assign w16955 = ~w16945 & w16954;
assign w16956 = (~w16955 & w16936) | (~w16955 & w35861) | (w16936 & w35861);
assign w16957 = w5286 & ~w12860;
assign w16958 = w5016 & w12622;
assign w16959 = w5080 & w12856;
assign w16960 = ~w16958 & ~w16959;
assign w16961 = ~w16957 & w16960;
assign w16962 = (w16961 & ~w14442) | (w16961 & w35862) | (~w14442 & w35862);
assign w16963 = ~a_23 & w16962;
assign w16964 = (w14442 & w35863) | (w14442 & w35864) | (w35863 & w35864);
assign w16965 = ~w16963 & ~w16964;
assign w16966 = ~w16530 & w16965;
assign w16967 = w16530 & ~w16965;
assign w16968 = ~w16966 & ~w16967;
assign w16969 = w16514 & w16968;
assign w16970 = ~w16514 & ~w16968;
assign w16971 = ~w16969 & ~w16970;
assign w16972 = ~w16965 & ~w16971;
assign w16973 = (~w16972 & w16956) | (~w16972 & w35865) | (w16956 & w35865);
assign w16974 = w16592 & w16973;
assign w16975 = w16586 & ~w16592;
assign w16976 = ~w16974 & ~w16975;
assign w16977 = ~w16576 & ~w16976;
assign w16978 = w16576 & w16976;
assign w16979 = ~w16977 & ~w16978;
assign w16980 = ~w12930 & w35866;
assign w16981 = w6059 & ~w12910;
assign w16982 = ~w12914 & w35867;
assign w16983 = ~w13501 & w35868;
assign w16984 = ~w16981 & ~w16982;
assign w16985 = ~w16980 & w16984;
assign w16986 = ~w16983 & w35869;
assign w16987 = (a_17 & w16983) | (a_17 & w35870) | (w16983 & w35870);
assign w16988 = ~w16986 & ~w16987;
assign w16989 = w16979 & w16988;
assign w16990 = (~w16977 & ~w16979) | (~w16977 & w35871) | (~w16979 & w35871);
assign w16991 = w16574 & w16990;
assign w16992 = ~w16574 & ~w16990;
assign w16993 = ~w16991 & ~w16992;
assign w16994 = w6996 & w12604;
assign w16995 = ~w12589 & w35872;
assign w16996 = (w6446 & w12616) | (w6446 & w35873) | (w12616 & w35873);
assign w16997 = ~w16995 & ~w16996;
assign w16998 = ~w16994 & w16997;
assign w16999 = (w16998 & w13288) | (w16998 & w35874) | (w13288 & w35874);
assign w17000 = a_14 & ~w16999;
assign w17001 = (w13288 & w35875) | (w13288 & w35876) | (w35875 & w35876);
assign w17002 = ~w17000 & ~w17001;
assign w17003 = w16993 & ~w17002;
assign w17004 = (~w16991 & ~w16993) | (~w16991 & w35877) | (~w16993 & w35877);
assign w17005 = (~w16571 & ~w17004) | (~w16571 & w35878) | (~w17004 & w35878);
assign w17006 = ~w16557 & ~w17005;
assign w17007 = w16557 & w17005;
assign w17008 = ~w17006 & ~w17007;
assign w17009 = w7511 & w13177;
assign w17010 = ~w13174 & w35879;
assign w17011 = ~w13011 & w35880;
assign w17012 = ~w17010 & ~w17011;
assign w17013 = ~w17009 & w17012;
assign w17014 = (w17013 & ~w13207) | (w17013 & w35881) | (~w13207 & w35881);
assign w17015 = a_11 & w17014;
assign w17016 = (w13207 & w35882) | (w13207 & w35883) | (w35882 & w35883);
assign w17017 = ~w17015 & ~w17016;
assign w17018 = w17008 & ~w17017;
assign w17019 = (~w17006 & ~w17008) | (~w17006 & w35884) | (~w17008 & w35884);
assign w17020 = w14079 & ~w17019;
assign w17021 = ~w14079 & w17019;
assign w17022 = ~w17020 & ~w17021;
assign w17023 = (~w16179 & ~w16181) | (~w16179 & w35885) | (~w16181 & w35885);
assign w17024 = ~w15794 & w15803;
assign w17025 = ~w15804 & ~w17024;
assign w17026 = ~w17023 & ~w17025;
assign w17027 = w17023 & w17025;
assign w17028 = ~w17026 & ~w17027;
assign w17029 = ~w13011 & w35886;
assign w17030 = w6998 & w12598;
assign w17031 = w6446 & w12601;
assign w17032 = ~w17030 & ~w17031;
assign w17033 = ~w17029 & w17032;
assign w17034 = (w17033 & w13021) | (w17033 & w35887) | (w13021 & w35887);
assign w17035 = ~a_14 & w17034;
assign w17036 = (~w13021 & w35888) | (~w13021 & w35889) | (w35888 & w35889);
assign w17037 = ~w17035 & ~w17036;
assign w17038 = w17028 & w17037;
assign w17039 = ~w17028 & ~w17037;
assign w17040 = ~w17038 & ~w17039;
assign w17041 = ~w16552 & ~w16555;
assign w17042 = w17040 & w17041;
assign w17043 = ~w17040 & ~w17041;
assign w17044 = ~w17042 & ~w17043;
assign w17045 = w7489 & w13177;
assign w17046 = ~w13174 & w35890;
assign w17047 = (w13173 & w35891) | (w13173 & w35892) | (w35891 & w35892);
assign w17048 = ~w17046 & ~w17047;
assign w17049 = ~w17045 & w17048;
assign w17050 = (w17049 & w13264) | (w17049 & w35893) | (w13264 & w35893);
assign w17051 = ~a_11 & w17050;
assign w17052 = (~w13264 & w35894) | (~w13264 & w35895) | (w35894 & w35895);
assign w17053 = ~w17051 & ~w17052;
assign w17054 = w17044 & ~w17053;
assign w17055 = ~w17044 & w17053;
assign w17056 = ~w17054 & ~w17055;
assign w17057 = w17022 & ~w17056;
assign w17058 = (~w17020 & w17056) | (~w17020 & w35896) | (w17056 & w35896);
assign w17059 = (~w17026 & ~w17028) | (~w17026 & w35897) | (~w17028 & w35897);
assign w17060 = ~w15805 & ~w15807;
assign w17061 = ~w15808 & ~w17060;
assign w17062 = ~w13174 & w35898;
assign w17063 = ~w13011 & w35899;
assign w17064 = w6446 & w12598;
assign w17065 = ~w13205 & w35900;
assign w17066 = ~w17063 & w35901;
assign w17067 = (a_14 & w17065) | (a_14 & w35902) | (w17065 & w35902);
assign w17068 = ~w17065 & w35903;
assign w17069 = ~w17067 & ~w17068;
assign w17070 = w17061 & w17069;
assign w17071 = ~w17061 & ~w17069;
assign w17072 = ~w17070 & ~w17071;
assign w17073 = ~w17059 & w17072;
assign w17074 = w17059 & ~w17072;
assign w17075 = ~w17073 & ~w17074;
assign w17076 = (~w17043 & ~w17044) | (~w17043 & w35904) | (~w17044 & w35904);
assign w17077 = w7192 & w13177;
assign w17078 = (w13201 & w35907) | (w13201 & w35908) | (w35907 & w35908);
assign w17079 = (~w13173 & w35909) | (~w13173 & w35910) | (w35909 & w35910);
assign w17080 = ~w17077 & w17079;
assign w17081 = (a_11 & w17078) | (a_11 & w35911) | (w17078 & w35911);
assign w17082 = ~w17078 & w35912;
assign w17083 = ~w17081 & ~w17082;
assign w17084 = w17076 & w17083;
assign w17085 = ~w17076 & ~w17083;
assign w17086 = ~w17084 & ~w17085;
assign w17087 = w17075 & w17086;
assign w17088 = ~w17075 & ~w17086;
assign w17089 = ~w17087 & ~w17088;
assign w17090 = ~w17058 & w17089;
assign w17091 = ~w17008 & w17017;
assign w17092 = ~w17018 & ~w17091;
assign w17093 = ~w13174 & w35913;
assign w17094 = ~w13011 & w35914;
assign w17095 = w7192 & w12598;
assign w17096 = ~w13205 & w35915;
assign w17097 = ~w17094 & w35916;
assign w17098 = (a_11 & w17096) | (a_11 & w35917) | (w17096 & w35917);
assign w17099 = ~w17096 & w35918;
assign w17100 = ~w17098 & ~w17099;
assign w17101 = ~w16571 & ~w16572;
assign w17102 = w17004 & w17101;
assign w17103 = ~w17004 & ~w17101;
assign w17104 = ~w17102 & ~w17103;
assign w17105 = ~w17100 & ~w17104;
assign w17106 = w17100 & w17104;
assign w17107 = ~w16592 & ~w16973;
assign w17108 = ~w16974 & ~w17107;
assign w17109 = ~w12914 & w35919;
assign w17110 = w6061 & ~w12910;
assign w17111 = ~w12905 & w35920;
assign w17112 = (w6063 & w13518) | (w6063 & w35921) | (w13518 & w35921);
assign w17113 = ~w17110 & ~w17111;
assign w17114 = ~w17109 & w17113;
assign w17115 = (a_17 & w17112) | (a_17 & w35922) | (w17112 & w35922);
assign w17116 = ~w17112 & w35923;
assign w17117 = ~w17115 & ~w17116;
assign w17118 = w17108 & w17117;
assign w17119 = ~w17108 & ~w17117;
assign w17120 = ~w17118 & ~w17119;
assign w17121 = w5816 & w12874;
assign w17122 = w5308 & ~w12860;
assign w17123 = w5818 & w12869;
assign w17124 = w5309 & w13965;
assign w17125 = ~w17122 & w35924;
assign w17126 = (a_20 & w17124) | (a_20 & w35925) | (w17124 & w35925);
assign w17127 = ~w17124 & w35926;
assign w17128 = ~w17126 & ~w17127;
assign w17129 = ~w16954 & ~w17128;
assign w17130 = w16936 & w17129;
assign w17131 = w16954 & ~w17128;
assign w17132 = ~w16936 & w17131;
assign w17133 = ~w17130 & ~w17132;
assign w17134 = w16954 & w17128;
assign w17135 = w16936 & w17134;
assign w17136 = ~w16954 & w17128;
assign w17137 = ~w16936 & w17136;
assign w17138 = ~w17135 & ~w17137;
assign w17139 = w5308 & w12856;
assign w17140 = w5816 & w12869;
assign w17141 = (~w17139 & w12860) | (~w17139 & w35927) | (w12860 & w35927);
assign w17142 = ~w17140 & w17141;
assign w17143 = (w17142 & ~w13979) | (w17142 & w35928) | (~w13979 & w35928);
assign w17144 = ~a_20 & w17143;
assign w17145 = (w13979 & w35929) | (w13979 & w35930) | (w35929 & w35930);
assign w17146 = ~w17144 & ~w17145;
assign w17147 = (~w16934 & w16906) | (~w16934 & w35931) | (w16906 & w35931);
assign w17148 = ~w16611 & w17146;
assign w17149 = w16611 & ~w17146;
assign w17150 = ~w17148 & ~w17149;
assign w17151 = w17147 & w17150;
assign w17152 = ~w17147 & ~w17150;
assign w17153 = ~w17151 & ~w17152;
assign w17154 = ~w17146 & ~w17153;
assign w17155 = (w16926 & w16889) | (w16926 & w35932) | (w16889 & w35932);
assign w17156 = w8311 & w14442;
assign w17157 = w5818 & w12856;
assign w17158 = w5308 & w12622;
assign w17159 = w5816 & ~w12860;
assign w17160 = ~w17157 & ~w17158;
assign w17161 = ~w17159 & w35933;
assign w17162 = (~a_20 & w17159) | (~a_20 & w35934) | (w17159 & w35934);
assign w17163 = ~w17161 & ~w17162;
assign w17164 = (w17163 & ~w14442) | (w17163 & w35935) | (~w14442 & w35935);
assign w17165 = ~w17156 & ~w17164;
assign w17166 = ~w16910 & w16920;
assign w17167 = ~w16927 & ~w17166;
assign w17168 = w16909 & ~w17167;
assign w17169 = ~w16909 & w17167;
assign w17170 = ~w17168 & ~w17169;
assign w17171 = ~w17165 & ~w17170;
assign w17172 = w17155 & w17171;
assign w17173 = ~w17165 & w17170;
assign w17174 = ~w17155 & w17173;
assign w17175 = ~w17172 & ~w17174;
assign w17176 = w17165 & w17170;
assign w17177 = w17155 & w17176;
assign w17178 = w17165 & ~w17170;
assign w17179 = ~w17155 & w17178;
assign w17180 = ~w17177 & ~w17179;
assign w17181 = (~w16890 & w16863) | (~w16890 & w35936) | (w16863 & w35936);
assign w17182 = ~w16902 & ~w16924;
assign w17183 = w5818 & w12622;
assign w17184 = w5308 & ~w12630;
assign w17185 = w5816 & w12856;
assign w17186 = ~w17183 & ~w17184;
assign w17187 = ~w17185 & w17186;
assign w17188 = (w17187 & ~w14091) | (w17187 & w35937) | (~w14091 & w35937);
assign w17189 = ~a_20 & w17188;
assign w17190 = (w14091 & w35938) | (w14091 & w35939) | (w35938 & w35939);
assign w17191 = ~w17189 & ~w17190;
assign w17192 = w16467 & ~w17191;
assign w17193 = ~w16467 & w17191;
assign w17194 = ~w17192 & ~w17193;
assign w17195 = w17182 & w17194;
assign w17196 = ~w17182 & ~w17194;
assign w17197 = ~w17195 & ~w17196;
assign w17198 = ~w17181 & ~w17197;
assign w17199 = w16904 & w16926;
assign w17200 = w17181 & ~w17199;
assign w17201 = w17191 & ~w17198;
assign w17202 = ~w17200 & w17201;
assign w17203 = w17180 & ~w17202;
assign w17204 = w17175 & ~w17203;
assign w17205 = w5818 & ~w12630;
assign w17206 = w5308 & ~w12668;
assign w17207 = w5816 & w12622;
assign w17208 = ~w17205 & ~w17206;
assign w17209 = ~w17207 & w17208;
assign w17210 = (w17209 & w14412) | (w17209 & w35940) | (w14412 & w35940);
assign w17211 = a_20 & ~w17210;
assign w17212 = (w14412 & w35941) | (w14412 & w35942) | (w35941 & w35942);
assign w17213 = ~w17211 & ~w17212;
assign w17214 = ~w16863 & w35943;
assign w17215 = (~w16864 & w16849) | (~w16864 & w31851) | (w16849 & w31851);
assign w17216 = w16887 & ~w17213;
assign w17217 = ~w17215 & w17216;
assign w17218 = ~w17214 & ~w17217;
assign w17219 = ~w16626 & w16841;
assign w17220 = ~w16797 & w17219;
assign w17221 = w16816 & ~w17220;
assign w17222 = w16834 & w16846;
assign w17223 = w5816 & ~w12668;
assign w17224 = w5308 & ~w12637;
assign w17225 = w5818 & ~w12661;
assign w17226 = ~w17224 & ~w17225;
assign w17227 = ~w17223 & w17226;
assign w17228 = (w17227 & ~w14393) | (w17227 & w35944) | (~w14393 & w35944);
assign w17229 = ~a_20 & w17228;
assign w17230 = (w14393 & w35945) | (w14393 & w35946) | (w35945 & w35946);
assign w17231 = ~w17229 & ~w17230;
assign w17232 = ~w17222 & ~w17231;
assign w17233 = w17221 & w17232;
assign w17234 = w17222 & ~w17231;
assign w17235 = ~w17221 & w17234;
assign w17236 = ~w17233 & ~w17235;
assign w17237 = w16816 & w16841;
assign w17238 = w5816 & ~w12661;
assign w17239 = w5818 & ~w12637;
assign w17240 = w5308 & w12646;
assign w17241 = ~w17239 & ~w17240;
assign w17242 = ~w17238 & w17241;
assign w17243 = (w17242 & w14641) | (w17242 & w35947) | (w14641 & w35947);
assign w17244 = a_20 & w17243;
assign w17245 = (~w14641 & w35948) | (~w14641 & w35949) | (w35948 & w35949);
assign w17246 = ~w17244 & ~w17245;
assign w17247 = w17237 & w17246;
assign w17248 = ~w17237 & ~w17246;
assign w17249 = ~w17247 & ~w17248;
assign w17250 = w16798 & w17249;
assign w17251 = (~w17246 & w16798) | (~w17246 & w31852) | (w16798 & w31852);
assign w17252 = ~w17250 & w17251;
assign w17253 = w17222 & w17231;
assign w17254 = w17221 & w17253;
assign w17255 = ~w17222 & w17231;
assign w17256 = ~w17221 & w17255;
assign w17257 = ~w17254 & ~w17256;
assign w17258 = ~w17252 & w17257;
assign w17259 = w17236 & ~w17258;
assign w17260 = ~w16773 & ~w16789;
assign w17261 = ~w16790 & ~w17260;
assign w17262 = w8311 & w14614;
assign w17263 = w5816 & w12651;
assign w17264 = w5308 & w12793;
assign w17265 = w5818 & ~w12830;
assign w17266 = ~w17263 & ~w17264;
assign w17267 = ~w17265 & w35950;
assign w17268 = (~a_20 & w17265) | (~a_20 & w35951) | (w17265 & w35951);
assign w17269 = ~w17267 & ~w17268;
assign w17270 = (w17269 & ~w14614) | (w17269 & w35952) | (~w14614 & w35952);
assign w17271 = ~w17262 & ~w17270;
assign w17272 = ~w17261 & ~w17271;
assign w17273 = w16748 & ~w16765;
assign w17274 = ~w16766 & ~w17273;
assign w17275 = w8311 & ~w15101;
assign w17276 = w5818 & w12789;
assign w17277 = ~w12770 & w35953;
assign w17278 = w5816 & w12793;
assign w17279 = ~w17276 & ~w17277;
assign w17280 = (~a_20 & ~w17279) | (~a_20 & w35954) | (~w17279 & w35954);
assign w17281 = w17279 & w35955;
assign w17282 = ~w17280 & ~w17281;
assign w17283 = (w17282 & w15101) | (w17282 & w35956) | (w15101 & w35956);
assign w17284 = ~w17275 & ~w17283;
assign w17285 = ~w17274 & ~w17284;
assign w17286 = ~w12770 & w31853;
assign w17287 = w5308 & w12732;
assign w17288 = w5818 & ~w12774;
assign w17289 = ~w17286 & ~w17287;
assign w17290 = (~a_20 & ~w17289) | (~a_20 & w35957) | (~w17289 & w35957);
assign w17291 = w17289 & w35958;
assign w17292 = ~w17290 & ~w17291;
assign w17293 = ~w15435 & w17292;
assign w17294 = ~w8311 & ~w11417;
assign w17295 = w17289 & w35959;
assign w17296 = ~w17290 & ~w17295;
assign w17297 = w15435 & w17296;
assign w17298 = ~w17293 & ~w17297;
assign w17299 = ~w16727 & ~w16745;
assign w17300 = w16744 & ~w17299;
assign w17301 = ~w16744 & w17299;
assign w17302 = ~w17300 & ~w17301;
assign w17303 = ~w17298 & w17302;
assign w17304 = w12679 & w35960;
assign w17305 = w16703 & ~w17304;
assign w17306 = (a_23 & ~w16703) | (a_23 & w35961) | (~w16703 & w35961);
assign w17307 = ~w16697 & w17306;
assign w17308 = w16697 & ~w17306;
assign w17309 = ~w17307 & ~w17308;
assign w17310 = w5308 & w12701;
assign w17311 = w5816 & w12732;
assign w17312 = (~w17310 & ~w12739) | (~w17310 & w35962) | (~w12739 & w35962);
assign w17313 = ~w17311 & w17312;
assign w17314 = a_20 & w17313;
assign w17315 = w17309 & w17314;
assign w17316 = (w17315 & w15977) | (w17315 & w35963) | (w15977 & w35963);
assign w17317 = w8339 & w17309;
assign w17318 = ~a_20 & ~w17313;
assign w17319 = w17309 & w17318;
assign w17320 = (~w17319 & w15977) | (~w17319 & w35964) | (w15977 & w35964);
assign w17321 = ~w17316 & w17320;
assign w17322 = ~a_20 & w17313;
assign w17323 = ~w17309 & w17322;
assign w17324 = (w17323 & w15977) | (w17323 & w35965) | (w15977 & w35965);
assign w17325 = w8311 & ~w17309;
assign w17326 = a_20 & ~w17313;
assign w17327 = ~w17309 & w17326;
assign w17328 = (~w17327 & w15977) | (~w17327 & w35966) | (w15977 & w35966);
assign w17329 = ~w17324 & w17328;
assign w17330 = ~w16703 & w17304;
assign w17331 = ~w17305 & ~w17330;
assign w17332 = w12702 & w31854;
assign w17333 = w5309 & w15385;
assign w17334 = ~w12702 & w17333;
assign w17335 = w5308 & w12679;
assign w17336 = w5816 & w11683;
assign w17337 = w11678 & w17336;
assign w17338 = w5816 & ~w12675;
assign w17339 = ~w12674 & w17338;
assign w17340 = w5818 & ~w11501;
assign w17341 = w12684 & w17340;
assign w17342 = ~w17335 & ~w17337;
assign w17343 = ~w17339 & ~w17341;
assign w17344 = w17342 & w17343;
assign w17345 = ~w17334 & w17344;
assign w17346 = ~w17332 & w17345;
assign w17347 = w5300 & w12679;
assign w17348 = w12684 & w31855;
assign w17349 = w5818 & w12679;
assign w17350 = w5309 & ~w15324;
assign w17351 = ~w17348 & ~w17349;
assign w17352 = ~w17350 & w17351;
assign w17353 = (a_20 & ~w12679) | (a_20 & w35967) | (~w12679 & w35967);
assign w17354 = w17352 & w17353;
assign w17355 = (~w16698 & ~w17346) | (~w16698 & w31856) | (~w17346 & w31856);
assign w17356 = w5309 & w15283;
assign w17357 = w5309 & ~w12681;
assign w17358 = w12688 & w17357;
assign w17359 = ~w15282 & w17358;
assign w17360 = w5816 & ~w11825;
assign w17361 = ~w12699 & w17360;
assign w17362 = w11825 & w17336;
assign w17363 = ~w11678 & w17362;
assign w17364 = w15293 & w17340;
assign w17365 = ~w12674 & w31857;
assign w17366 = w12684 & w31858;
assign w17367 = ~w17363 & ~w17364;
assign w17368 = ~w17361 & w17367;
assign w17369 = ~w17365 & ~w17366;
assign w17370 = w17368 & w17369;
assign w17371 = ~w17359 & w17370;
assign w17372 = ~w17356 & w17371;
assign w17373 = a_20 & ~w17372;
assign w17374 = ~a_20 & w17372;
assign w17375 = ~w17373 & ~w17374;
assign w17376 = (~w17331 & ~w17375) | (~w17331 & w31859) | (~w17375 & w31859);
assign w17377 = w17375 & w31860;
assign w17378 = w5309 & w12715;
assign w17379 = w5816 & w12739;
assign w17380 = w5308 & w12702;
assign w17381 = w5818 & w12701;
assign w17382 = w5309 & ~w12700;
assign w17383 = w12711 & ~w17382;
assign w17384 = w5309 & w12700;
assign w17385 = ~w12711 & ~w17384;
assign w17386 = ~w17383 & ~w17385;
assign w17387 = ~w12704 & w17386;
assign w17388 = ~w17380 & ~w17381;
assign w17389 = ~w17379 & w17388;
assign w17390 = ~w17387 & w17389;
assign w17391 = ~w17378 & w17390;
assign w17392 = a_20 & ~w17391;
assign w17393 = ~a_20 & w17391;
assign w17394 = ~w17392 & ~w17393;
assign w17395 = (~w17376 & w17394) | (~w17376 & w31861) | (w17394 & w31861);
assign w17396 = w17329 & w17395;
assign w17397 = w17321 & ~w17396;
assign w17398 = w5818 & w12732;
assign w17399 = w5308 & w12739;
assign w17400 = w5816 & ~w12774;
assign w17401 = ~w17398 & ~w17399;
assign w17402 = ~w17400 & w17401;
assign w17403 = (w17402 & w15157) | (w17402 & w35968) | (w15157 & w35968);
assign w17404 = w16697 & w31862;
assign w17405 = ~w16706 & ~w17404;
assign w17406 = w16726 & w17405;
assign w17407 = ~w16726 & ~w17405;
assign w17408 = ~w17406 & ~w17407;
assign w17409 = ~a_20 & w17408;
assign w17410 = a_20 & ~w17408;
assign w17411 = ~w17409 & ~w17410;
assign w17412 = w17403 & w17411;
assign w17413 = ~w17403 & ~w17411;
assign w17414 = ~w17412 & ~w17413;
assign w17415 = ~w17397 & w17414;
assign w17416 = w17298 & ~w17302;
assign w17417 = ~w17403 & ~w17409;
assign w17418 = a_20 & w17408;
assign w17419 = w17403 & ~w17418;
assign w17420 = ~w17417 & ~w17419;
assign w17421 = ~w17416 & ~w17420;
assign w17422 = (~w17303 & w17415) | (~w17303 & w31863) | (w17415 & w31863);
assign w17423 = w5308 & ~w12774;
assign w17424 = w5816 & w12789;
assign w17425 = ~w12770 & w35969;
assign w17426 = ~w17424 & w35970;
assign w17427 = ~w5309 & w17426;
assign w17428 = ~w15127 & w17426;
assign w17429 = (~w17427 & ~w17428) | (~w17427 & w31864) | (~w17428 & w31864);
assign w17430 = ~a_20 & w17429;
assign w17431 = a_20 & ~w17429;
assign w17432 = ~w17430 & ~w17431;
assign w17433 = w16674 & w16680;
assign w17434 = ~w16746 & w17433;
assign w17435 = w16746 & ~w17433;
assign w17436 = ~w17434 & ~w17435;
assign w17437 = ~w17432 & ~w17436;
assign w17438 = w17432 & w17436;
assign w17439 = ~w17437 & ~w17438;
assign w17440 = w17422 & w17439;
assign w17441 = w17274 & w17284;
assign w17442 = (~w17437 & ~w17274) | (~w17437 & w37569) | (~w17274 & w37569);
assign w17443 = ~w17440 & w17442;
assign w17444 = ~w17285 & ~w17443;
assign w17445 = w8311 & w15071;
assign w17446 = w5818 & w12793;
assign w17447 = w5308 & w12789;
assign w17448 = w5816 & ~w12830;
assign w17449 = ~w17446 & ~w17447;
assign w17450 = (~a_20 & w17448) | (~a_20 & w35971) | (w17448 & w35971);
assign w17451 = ~w17448 & w35972;
assign w17452 = ~w17450 & ~w17451;
assign w17453 = (w17452 & ~w15071) | (w17452 & w35973) | (~w15071 & w35973);
assign w17454 = ~w17445 & ~w17453;
assign w17455 = ~w16660 & ~w16771;
assign w17456 = ~w16766 & w31865;
assign w17457 = (~w17455 & w16766) | (~w17455 & w31866) | (w16766 & w31866);
assign w17458 = ~w17456 & ~w17457;
assign w17459 = w17454 & ~w17458;
assign w17460 = ~w17454 & w17458;
assign w17461 = ~w17459 & ~w17460;
assign w17462 = w17444 & w17461;
assign w17463 = w17261 & w17271;
assign w17464 = (~w17459 & ~w17261) | (~w17459 & w31867) | (~w17261 & w31867);
assign w17465 = ~w17462 & w17464;
assign w17466 = (~w17272 & w17462) | (~w17272 & w31868) | (w17462 & w31868);
assign w17467 = (~w16787 & ~w16789) | (~w16787 & w31869) | (~w16789 & w31869);
assign w17468 = ~w16641 & ~w16791;
assign w17469 = ~w15044 & w35974;
assign w17470 = ~w15044 & w35975;
assign w17471 = w5816 & w12646;
assign w17472 = w5818 & w12651;
assign w17473 = (~w17471 & w12830) | (~w17471 & w35976) | (w12830 & w35976);
assign w17474 = (~a_20 & ~w17473) | (~a_20 & w35977) | (~w17473 & w35977);
assign w17475 = w17473 & w35978;
assign w17476 = ~w17474 & ~w17475;
assign w17477 = ~w17470 & w17476;
assign w17478 = ~w17469 & ~w17477;
assign w17479 = ~w17468 & ~w17478;
assign w17480 = w17468 & w17478;
assign w17481 = ~w17479 & ~w17480;
assign w17482 = w17467 & w17481;
assign w17483 = ~w17467 & ~w17481;
assign w17484 = ~w17482 & ~w17483;
assign w17485 = w17466 & ~w17484;
assign w17486 = w17478 & w17484;
assign w17487 = w16794 & ~w16796;
assign w17488 = ~w16797 & ~w17487;
assign w17489 = w8311 & ~w15027;
assign w17490 = w5816 & ~w12637;
assign w17491 = w5308 & w12651;
assign w17492 = w5818 & w12646;
assign w17493 = ~w17490 & w35979;
assign w17494 = a_20 & ~w17493;
assign w17495 = ~a_20 & w17493;
assign w17496 = (w17495 & w15027) | (w17495 & w35980) | (w15027 & w35980);
assign w17497 = ~w17489 & ~w17494;
assign w17498 = ~w17496 & w17497;
assign w17499 = ~w17488 & w17498;
assign w17500 = ~w17486 & ~w17499;
assign w17501 = ~w17485 & w17500;
assign w17502 = w17488 & ~w17498;
assign w17503 = (~w17502 & ~w17500) | (~w17502 & w31870) | (~w17500 & w31870);
assign w17504 = ~w16798 & ~w17249;
assign w17505 = ~w17250 & ~w17504;
assign w17506 = w17236 & ~w17505;
assign w17507 = w17503 & w17506;
assign w17508 = ~w17259 & ~w17507;
assign w17509 = w8311 & ~w14535;
assign w17510 = ~w14391 & w35981;
assign w17511 = w8339 & ~w14532;
assign w17512 = w5818 & ~w12668;
assign w17513 = w5308 & ~w12661;
assign w17514 = w5816 & ~w12630;
assign w17515 = ~w17512 & ~w17513;
assign w17516 = (a_20 & ~w17515) | (a_20 & w35983) | (~w17515 & w35983);
assign w17517 = w17515 & w35984;
assign w17518 = ~w17516 & ~w17517;
assign w17519 = (~w14391 & w35985) | (~w14391 & w35986) | (w35985 & w35986);
assign w17520 = ~w17510 & w17519;
assign w17521 = ~w17509 & ~w17520;
assign w17522 = ~w16861 & w17521;
assign w17523 = w16861 & ~w17521;
assign w17524 = ~w17522 & ~w17523;
assign w17525 = w16851 & ~w17524;
assign w17526 = ~w16851 & w17524;
assign w17527 = ~w17525 & ~w17526;
assign w17528 = w16849 & w17527;
assign w17529 = ~w16849 & ~w17527;
assign w17530 = ~w17528 & ~w17529;
assign w17531 = ~w17508 & w17530;
assign w17532 = w17521 & ~w17530;
assign w17533 = w16887 & w17213;
assign w17534 = w17215 & w17533;
assign w17535 = ~w16887 & w17213;
assign w17536 = ~w17215 & w17535;
assign w17537 = ~w17534 & ~w17536;
assign w17538 = ~w17532 & w17537;
assign w17539 = (w17218 & w17531) | (w17218 & w31871) | (w17531 & w31871);
assign w17540 = w17181 & w17197;
assign w17541 = ~w17198 & ~w17540;
assign w17542 = w17175 & ~w17541;
assign w17543 = w17539 & w17542;
assign w17544 = ~w17204 & ~w17543;
assign w17545 = (~w17154 & ~w17544) | (~w17154 & w31872) | (~w17544 & w31872);
assign w17546 = (w17133 & w17545) | (w17133 & w35987) | (w17545 & w35987);
assign w17547 = w5816 & ~w12878;
assign w17548 = w5818 & w12874;
assign w17549 = w5308 & w12869;
assign w17550 = ~w17548 & ~w17549;
assign w17551 = ~w17547 & w17550;
assign w17552 = (w17551 & ~w13771) | (w17551 & w35988) | (~w13771 & w35988);
assign w17553 = a_20 & ~w17552;
assign w17554 = (~w13771 & w35989) | (~w13771 & w35990) | (w35989 & w35990);
assign w17555 = ~w17553 & ~w17554;
assign w17556 = ~w16971 & w17555;
assign w17557 = w16971 & ~w17555;
assign w17558 = ~w17556 & ~w17557;
assign w17559 = w16956 & w17558;
assign w17560 = ~w16956 & ~w17558;
assign w17561 = ~w17559 & ~w17560;
assign w17562 = (~w17545 & w35991) | (~w17545 & w35992) | (w35991 & w35992);
assign w17563 = ~w17555 & w17561;
assign w17564 = ~w17562 & ~w17563;
assign w17565 = w17120 & w17564;
assign w17566 = ~w17118 & ~w17565;
assign w17567 = ~w16979 & ~w16988;
assign w17568 = ~w16989 & ~w17567;
assign w17569 = w17566 & ~w17568;
assign w17570 = ~w17566 & w17568;
assign w17571 = ~w17569 & ~w17570;
assign w17572 = (w6998 & w12616) | (w6998 & w35993) | (w12616 & w35993);
assign w17573 = (w6446 & w12612) | (w6446 & w35994) | (w12612 & w35994);
assign w17574 = ~w12589 & w35995;
assign w17575 = ~w17572 & ~w17573;
assign w17576 = ~w17574 & w17575;
assign w17577 = (w17576 & ~w13123) | (w17576 & w35996) | (~w13123 & w35996);
assign w17578 = a_14 & w17577;
assign w17579 = (w13123 & w35997) | (w13123 & w35998) | (w35997 & w35998);
assign w17580 = ~w17578 & ~w17579;
assign w17581 = w17571 & w17580;
assign w17582 = (~w17569 & ~w17571) | (~w17569 & w35999) | (~w17571 & w35999);
assign w17583 = ~w16993 & w17002;
assign w17584 = ~w17003 & ~w17583;
assign w17585 = ~w17582 & w17584;
assign w17586 = w17582 & ~w17584;
assign w17587 = ~w17585 & ~w17586;
assign w17588 = ~w13011 & w36000;
assign w17589 = w7489 & w12598;
assign w17590 = w7192 & w12601;
assign w17591 = ~w17589 & ~w17590;
assign w17592 = ~w17588 & w17591;
assign w17593 = (w17592 & w13021) | (w17592 & w36001) | (w13021 & w36001);
assign w17594 = ~a_11 & w17593;
assign w17595 = (~w13021 & w36002) | (~w13021 & w36003) | (w36002 & w36003);
assign w17596 = ~w17594 & ~w17595;
assign w17597 = w17587 & ~w17596;
assign w17598 = (~w17585 & ~w17587) | (~w17585 & w36004) | (~w17587 & w36004);
assign w17599 = (~w17105 & w17598) | (~w17105 & w36005) | (w17598 & w36005);
assign w17600 = w17092 & w17599;
assign w17601 = ~w17092 & ~w17599;
assign w17602 = ~w17600 & ~w17601;
assign w17603 = (~w13173 & w36008) | (~w13173 & w36009) | (w36008 & w36009);
assign w17604 = (~w13173 & w36010) | (~w13173 & w36011) | (w36010 & w36011);
assign w17605 = ~w17603 & w17604;
assign w17606 = ~w14077 & ~w17605;
assign w17607 = w17602 & w17606;
assign w17608 = (~w17600 & ~w17602) | (~w17600 & w36012) | (~w17602 & w36012);
assign w17609 = ~w17022 & w17056;
assign w17610 = ~w17057 & ~w17609;
assign w17611 = w17608 & ~w17610;
assign w17612 = ~w17090 & w17611;
assign w17613 = w17058 & ~w17089;
assign w17614 = ~w17070 & ~w17073;
assign w17615 = ~w15814 & ~w15823;
assign w17616 = ~w15824 & ~w17615;
assign w17617 = w17614 & ~w17616;
assign w17618 = ~w17614 & w17616;
assign w17619 = ~w17617 & ~w17618;
assign w17620 = (~w13173 & w36015) | (~w13173 & w36016) | (w36015 & w36016);
assign w17621 = (~w13173 & w36017) | (~w13173 & w36018) | (w36017 & w36018);
assign w17622 = ~w17620 & w17621;
assign w17623 = ~w13946 & ~w17622;
assign w17624 = w17619 & w17623;
assign w17625 = ~w17619 & ~w17623;
assign w17626 = ~w17624 & ~w17625;
assign w17627 = (~w17075 & ~w17076) | (~w17075 & w36019) | (~w17076 & w36019);
assign w17628 = ~w17085 & ~w17627;
assign w17629 = w17626 & w17628;
assign w17630 = ~w17626 & ~w17628;
assign w17631 = ~w17629 & ~w17630;
assign w17632 = ~w17613 & w17631;
assign w17633 = ~w17612 & w17632;
assign w17634 = (~w17618 & ~w17619) | (~w17618 & w36020) | (~w17619 & w36020);
assign w17635 = ~w15828 & ~w15830;
assign w17636 = ~w15831 & ~w17635;
assign w17637 = w17634 & ~w17636;
assign w17638 = ~w12914 & w36021;
assign w17639 = w8298 & ~w12910;
assign w17640 = ~w12905 & w36022;
assign w17641 = (w8278 & w13518) | (w8278 & w36023) | (w13518 & w36023);
assign w17642 = ~w17639 & ~w17640;
assign w17643 = ~w17638 & w17642;
assign w17644 = ~w17641 & w36024;
assign w17645 = (a_8 & w17641) | (a_8 & w36025) | (w17641 & w36025);
assign w17646 = ~w17644 & ~w17645;
assign w17647 = w7511 & ~w12878;
assign w17648 = w7489 & w12874;
assign w17649 = w7192 & w12869;
assign w17650 = ~w17648 & ~w17649;
assign w17651 = ~w17647 & w17650;
assign w17652 = (w17651 & ~w13771) | (w17651 & w36026) | (~w13771 & w36026);
assign w17653 = a_11 & ~w17652;
assign w17654 = (~w13771 & w36027) | (~w13771 & w36028) | (w36027 & w36028);
assign w17655 = ~w17653 & ~w17654;
assign w17656 = ~w17422 & ~w17439;
assign w17657 = ~w17440 & ~w17656;
assign w17658 = w8391 & w14614;
assign w17659 = w6304 & w12651;
assign w17660 = w6059 & w12793;
assign w17661 = w6061 & ~w12830;
assign w17662 = ~w17659 & ~w17660;
assign w17663 = ~w17661 & w36029;
assign w17664 = (~a_17 & w17661) | (~a_17 & w36030) | (w17661 & w36030);
assign w17665 = ~w17663 & ~w17664;
assign w17666 = (w17665 & ~w14614) | (w17665 & w36031) | (~w14614 & w36031);
assign w17667 = ~w17658 & ~w17666;
assign w17668 = ~w17657 & ~w17667;
assign w17669 = w17397 & ~w17414;
assign w17670 = ~w17415 & ~w17669;
assign w17671 = w8391 & ~w15101;
assign w17672 = w6061 & w12789;
assign w17673 = ~w12770 & w36032;
assign w17674 = w6304 & w12793;
assign w17675 = ~w17672 & ~w17673;
assign w17676 = (~a_17 & ~w17675) | (~a_17 & w36033) | (~w17675 & w36033);
assign w17677 = w17675 & w36034;
assign w17678 = ~w17676 & ~w17677;
assign w17679 = (w17678 & w15101) | (w17678 & w36035) | (w15101 & w36035);
assign w17680 = ~w17671 & ~w17679;
assign w17681 = ~w17670 & ~w17680;
assign w17682 = ~w17376 & ~w17377;
assign w17683 = ~w17394 & w17682;
assign w17684 = w17394 & ~w17682;
assign w17685 = ~w17683 & ~w17684;
assign w17686 = ~w12770 & w31873;
assign w17687 = w6059 & w12732;
assign w17688 = w6061 & ~w12774;
assign w17689 = ~w17686 & ~w17687;
assign w17690 = (~a_17 & ~w17689) | (~a_17 & w36036) | (~w17689 & w36036);
assign w17691 = w17689 & w36037;
assign w17692 = ~w17690 & ~w17691;
assign w17693 = ~w15435 & w17692;
assign w17694 = ~a_17 & ~w6063;
assign w17695 = ~w8391 & ~w17694;
assign w17696 = w17689 & w36038;
assign w17697 = ~w17690 & ~w17696;
assign w17698 = w15435 & w17697;
assign w17699 = ~w17693 & ~w17698;
assign w17700 = w17685 & ~w17699;
assign w17701 = w12679 & w36039;
assign w17702 = w17352 & ~w17701;
assign w17703 = (a_20 & ~w17352) | (a_20 & w36040) | (~w17352 & w36040);
assign w17704 = ~w17346 & w17703;
assign w17705 = w17346 & ~w17703;
assign w17706 = ~w17704 & ~w17705;
assign w17707 = w6059 & w12701;
assign w17708 = w6304 & w12732;
assign w17709 = (~w17707 & ~w12739) | (~w17707 & w36041) | (~w12739 & w36041);
assign w17710 = ~w17708 & w17709;
assign w17711 = a_17 & w17710;
assign w17712 = w17706 & w17711;
assign w17713 = (w17712 & w15977) | (w17712 & w36042) | (w15977 & w36042);
assign w17714 = w8419 & w17706;
assign w17715 = ~a_17 & ~w17710;
assign w17716 = w17706 & w17715;
assign w17717 = (~w17716 & w15977) | (~w17716 & w36043) | (w15977 & w36043);
assign w17718 = ~w17713 & w17717;
assign w17719 = ~a_17 & w17710;
assign w17720 = ~w17706 & w17719;
assign w17721 = (w17720 & w15977) | (w17720 & w36044) | (w15977 & w36044);
assign w17722 = w8391 & ~w17706;
assign w17723 = a_17 & ~w17710;
assign w17724 = ~w17706 & w17723;
assign w17725 = (~w17724 & w15977) | (~w17724 & w36045) | (w15977 & w36045);
assign w17726 = ~w17721 & w17725;
assign w17727 = ~w17352 & w17701;
assign w17728 = ~w17702 & ~w17727;
assign w17729 = w12702 & w31874;
assign w17730 = w6063 & w15385;
assign w17731 = ~w12702 & w17730;
assign w17732 = w6059 & w12679;
assign w17733 = w6304 & w11683;
assign w17734 = w11678 & w17733;
assign w17735 = w6304 & ~w12675;
assign w17736 = ~w12674 & w17735;
assign w17737 = w6061 & ~w11501;
assign w17738 = w12684 & w17737;
assign w17739 = ~w17732 & ~w17734;
assign w17740 = ~w17736 & ~w17738;
assign w17741 = w17739 & w17740;
assign w17742 = ~w17731 & w17741;
assign w17743 = ~w17729 & w17742;
assign w17744 = w6054 & w12679;
assign w17745 = w12684 & w31875;
assign w17746 = w6061 & w12679;
assign w17747 = w6063 & ~w15324;
assign w17748 = ~w17745 & ~w17746;
assign w17749 = ~w17747 & w17748;
assign w17750 = (a_17 & ~w12679) | (a_17 & w36046) | (~w12679 & w36046);
assign w17751 = w17749 & w17750;
assign w17752 = (~w17347 & ~w17743) | (~w17347 & w31876) | (~w17743 & w31876);
assign w17753 = w6063 & w15283;
assign w17754 = w6063 & ~w12681;
assign w17755 = w12688 & w17754;
assign w17756 = ~w15282 & w17755;
assign w17757 = w6304 & ~w11825;
assign w17758 = ~w12699 & w17757;
assign w17759 = w11825 & w17733;
assign w17760 = ~w11678 & w17759;
assign w17761 = w15293 & w17737;
assign w17762 = ~w12674 & w31877;
assign w17763 = w12684 & w31878;
assign w17764 = ~w17760 & ~w17761;
assign w17765 = ~w17758 & w17764;
assign w17766 = ~w17762 & ~w17763;
assign w17767 = w17765 & w17766;
assign w17768 = ~w17756 & w17767;
assign w17769 = ~w17753 & w17768;
assign w17770 = a_17 & ~w17769;
assign w17771 = ~a_17 & w17769;
assign w17772 = ~w17770 & ~w17771;
assign w17773 = (~w17728 & ~w17772) | (~w17728 & w31879) | (~w17772 & w31879);
assign w17774 = w17772 & w31880;
assign w17775 = w6063 & w12715;
assign w17776 = w6304 & w12739;
assign w17777 = w6059 & w12702;
assign w17778 = w6061 & w12701;
assign w17779 = w6063 & ~w12700;
assign w17780 = w12711 & ~w17779;
assign w17781 = w6063 & w12700;
assign w17782 = ~w12711 & ~w17781;
assign w17783 = ~w17780 & ~w17782;
assign w17784 = ~w12704 & w17783;
assign w17785 = ~w17777 & ~w17778;
assign w17786 = ~w17776 & w17785;
assign w17787 = ~w17784 & w17786;
assign w17788 = ~w17775 & w17787;
assign w17789 = a_17 & ~w17788;
assign w17790 = ~a_17 & w17788;
assign w17791 = ~w17789 & ~w17790;
assign w17792 = (~w17773 & w17791) | (~w17773 & w31881) | (w17791 & w31881);
assign w17793 = w17726 & w17792;
assign w17794 = w17718 & ~w17793;
assign w17795 = w6061 & w12732;
assign w17796 = w6059 & w12739;
assign w17797 = w6304 & ~w12774;
assign w17798 = ~w17795 & ~w17796;
assign w17799 = ~w17797 & w17798;
assign w17800 = (w17799 & w15157) | (w17799 & w36047) | (w15157 & w36047);
assign w17801 = w17346 & w31882;
assign w17802 = ~w17355 & ~w17801;
assign w17803 = w17375 & w17802;
assign w17804 = ~w17375 & ~w17802;
assign w17805 = ~w17803 & ~w17804;
assign w17806 = ~a_17 & w17805;
assign w17807 = a_17 & ~w17805;
assign w17808 = ~w17806 & ~w17807;
assign w17809 = w17800 & w17808;
assign w17810 = ~w17800 & ~w17808;
assign w17811 = ~w17809 & ~w17810;
assign w17812 = ~w17794 & w17811;
assign w17813 = ~w17685 & w17699;
assign w17814 = ~w17800 & ~w17806;
assign w17815 = a_17 & w17805;
assign w17816 = w17800 & ~w17815;
assign w17817 = ~w17814 & ~w17816;
assign w17818 = ~w17813 & ~w17817;
assign w17819 = (~w17700 & w17812) | (~w17700 & w31883) | (w17812 & w31883);
assign w17820 = w6059 & ~w12774;
assign w17821 = w6304 & w12789;
assign w17822 = ~w12770 & w36048;
assign w17823 = ~w17821 & w36049;
assign w17824 = ~w6063 & w17823;
assign w17825 = ~w15127 & w17823;
assign w17826 = (~w17824 & ~w17825) | (~w17824 & w31884) | (~w17825 & w31884);
assign w17827 = ~a_17 & w17826;
assign w17828 = a_17 & ~w17826;
assign w17829 = ~w17827 & ~w17828;
assign w17830 = w17321 & w17329;
assign w17831 = ~w17395 & w17830;
assign w17832 = w17395 & ~w17830;
assign w17833 = ~w17831 & ~w17832;
assign w17834 = ~w17829 & ~w17833;
assign w17835 = w17829 & w17833;
assign w17836 = ~w17834 & ~w17835;
assign w17837 = w17819 & w17836;
assign w17838 = w17670 & w17680;
assign w17839 = (~w17834 & ~w17670) | (~w17834 & w36050) | (~w17670 & w36050);
assign w17840 = ~w17837 & w17839;
assign w17841 = ~w17681 & ~w17840;
assign w17842 = w8391 & w15071;
assign w17843 = w6061 & w12793;
assign w17844 = w6059 & w12789;
assign w17845 = w6304 & ~w12830;
assign w17846 = ~w17843 & ~w17844;
assign w17847 = (~a_17 & w17845) | (~a_17 & w36051) | (w17845 & w36051);
assign w17848 = ~w17845 & w36052;
assign w17849 = ~w17847 & ~w17848;
assign w17850 = (w17849 & ~w15071) | (w17849 & w36053) | (~w15071 & w36053);
assign w17851 = ~w17842 & ~w17850;
assign w17852 = ~w17303 & ~w17416;
assign w17853 = ~w17415 & w31885;
assign w17854 = (~w17852 & w17415) | (~w17852 & w31886) | (w17415 & w31886);
assign w17855 = ~w17853 & ~w17854;
assign w17856 = w17851 & ~w17855;
assign w17857 = ~w17851 & w17855;
assign w17858 = ~w17856 & ~w17857;
assign w17859 = w17841 & w17858;
assign w17860 = w17657 & w17667;
assign w17861 = (~w17856 & ~w17657) | (~w17856 & w31887) | (~w17657 & w31887);
assign w17862 = (~w17668 & w17859) | (~w17668 & w31888) | (w17859 & w31888);
assign w17863 = (~w17437 & ~w17439) | (~w17437 & w36054) | (~w17439 & w36054);
assign w17864 = ~w17285 & ~w17441;
assign w17865 = ~w15044 & w36055;
assign w17866 = ~w15044 & w36056;
assign w17867 = w6304 & w12646;
assign w17868 = w6061 & w12651;
assign w17869 = (~w17867 & w12830) | (~w17867 & w36057) | (w12830 & w36057);
assign w17870 = (~a_17 & ~w17869) | (~a_17 & w36058) | (~w17869 & w36058);
assign w17871 = w17869 & w36059;
assign w17872 = ~w17870 & ~w17871;
assign w17873 = ~w17866 & w17872;
assign w17874 = ~w17865 & ~w17873;
assign w17875 = w17864 & ~w17874;
assign w17876 = ~w17864 & w17874;
assign w17877 = ~w17875 & ~w17876;
assign w17878 = w17863 & w17877;
assign w17879 = ~w17863 & ~w17877;
assign w17880 = ~w17878 & ~w17879;
assign w17881 = w17862 & w17880;
assign w17882 = ~w17862 & ~w17880;
assign w17883 = ~w17881 & ~w17882;
assign w17884 = w8564 & w14393;
assign w17885 = w6998 & ~w12661;
assign w17886 = w6446 & ~w12637;
assign w17887 = w6996 & ~w12668;
assign w17888 = ~w17885 & ~w17886;
assign w17889 = w17888 & w36060;
assign w17890 = (~a_14 & ~w17888) | (~a_14 & w36061) | (~w17888 & w36061);
assign w17891 = ~w17889 & ~w17890;
assign w17892 = (w17891 & ~w14393) | (w17891 & w36062) | (~w14393 & w36062);
assign w17893 = ~w17884 & ~w17892;
assign w17894 = ~w17883 & ~w17893;
assign w17895 = ~w17819 & ~w17836;
assign w17896 = ~w17837 & ~w17895;
assign w17897 = w8564 & w14614;
assign w17898 = w6996 & w12651;
assign w17899 = w6446 & w12793;
assign w17900 = w6998 & ~w12830;
assign w17901 = ~w17898 & ~w17899;
assign w17902 = ~w17900 & w36063;
assign w17903 = (~a_14 & w17900) | (~a_14 & w36064) | (w17900 & w36064);
assign w17904 = ~w17902 & ~w17903;
assign w17905 = (w17904 & ~w14614) | (w17904 & w36065) | (~w14614 & w36065);
assign w17906 = ~w17897 & ~w17905;
assign w17907 = ~w17896 & ~w17906;
assign w17908 = w17794 & ~w17811;
assign w17909 = ~w17812 & ~w17908;
assign w17910 = w8564 & ~w15101;
assign w17911 = w6998 & w12789;
assign w17912 = ~w12770 & w36066;
assign w17913 = w6996 & w12793;
assign w17914 = ~w17911 & ~w17912;
assign w17915 = (~a_14 & ~w17914) | (~a_14 & w36067) | (~w17914 & w36067);
assign w17916 = w17914 & w36068;
assign w17917 = ~w17915 & ~w17916;
assign w17918 = (w17917 & w15101) | (w17917 & w36069) | (w15101 & w36069);
assign w17919 = ~w17910 & ~w17918;
assign w17920 = ~w17909 & ~w17919;
assign w17921 = ~w17773 & ~w17774;
assign w17922 = ~w17791 & w17921;
assign w17923 = w17791 & ~w17921;
assign w17924 = ~w17922 & ~w17923;
assign w17925 = ~w12770 & w31889;
assign w17926 = w6446 & w12732;
assign w17927 = w6998 & ~w12774;
assign w17928 = ~w17925 & ~w17926;
assign w17929 = (~a_14 & ~w17928) | (~a_14 & w36070) | (~w17928 & w36070);
assign w17930 = w17928 & w36071;
assign w17931 = ~w17929 & ~w17930;
assign w17932 = ~w15435 & w17931;
assign w17933 = (~a_14 & ~w6441) | (~a_14 & w36072) | (~w6441 & w36072);
assign w17934 = ~w8564 & ~w17933;
assign w17935 = w17928 & w36073;
assign w17936 = ~w17929 & ~w17935;
assign w17937 = w15435 & w17936;
assign w17938 = ~w17932 & ~w17937;
assign w17939 = w17924 & ~w17938;
assign w17940 = w12679 & w36074;
assign w17941 = w17749 & ~w17940;
assign w17942 = (a_17 & ~w17749) | (a_17 & w36075) | (~w17749 & w36075);
assign w17943 = ~w17743 & w17942;
assign w17944 = w17743 & ~w17942;
assign w17945 = ~w17943 & ~w17944;
assign w17946 = w6446 & w12701;
assign w17947 = w6996 & w12732;
assign w17948 = (~w17946 & ~w12739) | (~w17946 & w36076) | (~w12739 & w36076);
assign w17949 = ~w17947 & w17948;
assign w17950 = a_14 & w17949;
assign w17951 = w17945 & w17950;
assign w17952 = (w17951 & w15977) | (w17951 & w36077) | (w15977 & w36077);
assign w17953 = w8592 & w17945;
assign w17954 = ~a_14 & ~w17949;
assign w17955 = w17945 & w17954;
assign w17956 = (~w17955 & w15977) | (~w17955 & w36078) | (w15977 & w36078);
assign w17957 = ~w17952 & w17956;
assign w17958 = ~a_14 & w17949;
assign w17959 = ~w17945 & w17958;
assign w17960 = (w17959 & w15977) | (w17959 & w36079) | (w15977 & w36079);
assign w17961 = w8564 & ~w17945;
assign w17962 = a_14 & ~w17949;
assign w17963 = ~w17945 & w17962;
assign w17964 = (~w17963 & w15977) | (~w17963 & w36080) | (w15977 & w36080);
assign w17965 = ~w17960 & w17964;
assign w17966 = ~w17749 & w17940;
assign w17967 = ~w17941 & ~w17966;
assign w17968 = w12702 & w31890;
assign w17969 = w6447 & w15385;
assign w17970 = ~w12702 & w17969;
assign w17971 = w6996 & ~w12675;
assign w17972 = ~w12674 & w17971;
assign w17973 = w6446 & w12679;
assign w17974 = w6996 & w11683;
assign w17975 = w11678 & w17974;
assign w17976 = w6998 & ~w11501;
assign w17977 = w12684 & w17976;
assign w17978 = ~w17972 & ~w17973;
assign w17979 = ~w17975 & ~w17977;
assign w17980 = w17978 & w17979;
assign w17981 = ~w17970 & w17980;
assign w17982 = ~w17968 & w17981;
assign w17983 = w6441 & w12679;
assign w17984 = w12684 & w31891;
assign w17985 = w6998 & w12679;
assign w17986 = w6447 & ~w15324;
assign w17987 = ~w17984 & ~w17985;
assign w17988 = ~w17986 & w17987;
assign w17989 = (a_14 & ~w12679) | (a_14 & w36081) | (~w12679 & w36081);
assign w17990 = w17988 & w17989;
assign w17991 = (~w17744 & ~w17982) | (~w17744 & w31892) | (~w17982 & w31892);
assign w17992 = w6447 & w15283;
assign w17993 = w6447 & ~w12681;
assign w17994 = w12688 & w17993;
assign w17995 = ~w15282 & w17994;
assign w17996 = w6996 & ~w11825;
assign w17997 = ~w12699 & w17996;
assign w17998 = w11825 & w17974;
assign w17999 = ~w11678 & w17998;
assign w18000 = w15293 & w17976;
assign w18001 = ~w12674 & w31893;
assign w18002 = w12684 & w31894;
assign w18003 = ~w17999 & ~w18000;
assign w18004 = ~w17997 & w18003;
assign w18005 = ~w18001 & ~w18002;
assign w18006 = w18004 & w18005;
assign w18007 = ~w17995 & w18006;
assign w18008 = ~w17992 & w18007;
assign w18009 = a_14 & ~w18008;
assign w18010 = ~a_14 & w18008;
assign w18011 = ~w18009 & ~w18010;
assign w18012 = (~w17967 & ~w18011) | (~w17967 & w31895) | (~w18011 & w31895);
assign w18013 = w18011 & w31896;
assign w18014 = w6447 & w12715;
assign w18015 = w6996 & w12739;
assign w18016 = w6446 & w12702;
assign w18017 = w6998 & w12701;
assign w18018 = w6447 & ~w12700;
assign w18019 = w12711 & ~w18018;
assign w18020 = w6447 & w12700;
assign w18021 = ~w12711 & ~w18020;
assign w18022 = ~w18019 & ~w18021;
assign w18023 = ~w12704 & w18022;
assign w18024 = ~w18016 & ~w18017;
assign w18025 = ~w18015 & w18024;
assign w18026 = ~w18023 & w18025;
assign w18027 = ~w18014 & w18026;
assign w18028 = a_14 & ~w18027;
assign w18029 = ~a_14 & w18027;
assign w18030 = ~w18028 & ~w18029;
assign w18031 = (~w18012 & w18030) | (~w18012 & w31897) | (w18030 & w31897);
assign w18032 = w17965 & w18031;
assign w18033 = w17957 & ~w18032;
assign w18034 = w6998 & w12732;
assign w18035 = w6446 & w12739;
assign w18036 = w6996 & ~w12774;
assign w18037 = ~w18034 & ~w18035;
assign w18038 = ~w18036 & w18037;
assign w18039 = (w18038 & w15157) | (w18038 & w36082) | (w15157 & w36082);
assign w18040 = w17743 & w31898;
assign w18041 = ~w17752 & ~w18040;
assign w18042 = w17772 & w18041;
assign w18043 = ~w17772 & ~w18041;
assign w18044 = ~w18042 & ~w18043;
assign w18045 = ~a_14 & w18044;
assign w18046 = a_14 & ~w18044;
assign w18047 = ~w18045 & ~w18046;
assign w18048 = w18039 & w18047;
assign w18049 = ~w18039 & ~w18047;
assign w18050 = ~w18048 & ~w18049;
assign w18051 = ~w18033 & w18050;
assign w18052 = ~w17924 & w17938;
assign w18053 = ~w18039 & ~w18045;
assign w18054 = a_14 & w18044;
assign w18055 = w18039 & ~w18054;
assign w18056 = ~w18053 & ~w18055;
assign w18057 = ~w18052 & ~w18056;
assign w18058 = (~w17939 & w18051) | (~w17939 & w31899) | (w18051 & w31899);
assign w18059 = w6446 & ~w12774;
assign w18060 = w6996 & w12789;
assign w18061 = ~w12770 & w36083;
assign w18062 = ~w18060 & w36084;
assign w18063 = ~w6447 & w18062;
assign w18064 = ~w15127 & w18062;
assign w18065 = (~w18063 & ~w18064) | (~w18063 & w31900) | (~w18064 & w31900);
assign w18066 = ~a_14 & w18065;
assign w18067 = a_14 & ~w18065;
assign w18068 = ~w18066 & ~w18067;
assign w18069 = w17718 & w17726;
assign w18070 = ~w17792 & w18069;
assign w18071 = w17792 & ~w18069;
assign w18072 = ~w18070 & ~w18071;
assign w18073 = ~w18068 & ~w18072;
assign w18074 = w18068 & w18072;
assign w18075 = ~w18073 & ~w18074;
assign w18076 = w18058 & w18075;
assign w18077 = w17909 & w17919;
assign w18078 = (~w18073 & ~w17909) | (~w18073 & w36085) | (~w17909 & w36085);
assign w18079 = ~w18076 & w18078;
assign w18080 = ~w17920 & ~w18079;
assign w18081 = w8564 & w15071;
assign w18082 = w6998 & w12793;
assign w18083 = w6446 & w12789;
assign w18084 = w6996 & ~w12830;
assign w18085 = ~w18082 & ~w18083;
assign w18086 = (~a_14 & w18084) | (~a_14 & w36086) | (w18084 & w36086);
assign w18087 = ~w18084 & w36087;
assign w18088 = ~w18086 & ~w18087;
assign w18089 = (w18088 & ~w15071) | (w18088 & w36088) | (~w15071 & w36088);
assign w18090 = ~w18081 & ~w18089;
assign w18091 = ~w17700 & ~w17813;
assign w18092 = ~w17812 & w31901;
assign w18093 = (~w18091 & w17812) | (~w18091 & w31902) | (w17812 & w31902);
assign w18094 = ~w18092 & ~w18093;
assign w18095 = w18090 & ~w18094;
assign w18096 = ~w18090 & w18094;
assign w18097 = ~w18095 & ~w18096;
assign w18098 = w18080 & w18097;
assign w18099 = w17896 & w17906;
assign w18100 = (~w18095 & ~w17896) | (~w18095 & w31903) | (~w17896 & w31903);
assign w18101 = (~w17907 & w18098) | (~w17907 & w31904) | (w18098 & w31904);
assign w18102 = ~w17834 & ~w17837;
assign w18103 = ~w17681 & ~w17838;
assign w18104 = ~w15044 & w36089;
assign w18105 = ~w15044 & w36090;
assign w18106 = w6996 & w12646;
assign w18107 = w6998 & w12651;
assign w18108 = (~w18106 & w12830) | (~w18106 & w36091) | (w12830 & w36091);
assign w18109 = (~a_14 & ~w18108) | (~a_14 & w36092) | (~w18108 & w36092);
assign w18110 = w18108 & w36093;
assign w18111 = ~w18109 & ~w18110;
assign w18112 = ~w18105 & w18111;
assign w18113 = ~w18104 & ~w18112;
assign w18114 = w18103 & ~w18113;
assign w18115 = ~w18103 & w18113;
assign w18116 = ~w18114 & ~w18115;
assign w18117 = w18102 & w18116;
assign w18118 = ~w18102 & ~w18116;
assign w18119 = ~w18117 & ~w18118;
assign w18120 = w18101 & w18119;
assign w18121 = w18113 & ~w18119;
assign w18122 = ~w17841 & ~w17858;
assign w18123 = ~w17859 & ~w18122;
assign w18124 = w8564 & ~w15027;
assign w18125 = w6996 & ~w12637;
assign w18126 = w6446 & w12651;
assign w18127 = w6998 & w12646;
assign w18128 = ~w18125 & w36094;
assign w18129 = a_14 & w18128;
assign w18130 = ~a_14 & ~w18128;
assign w18131 = ~w18129 & ~w18130;
assign w18132 = (w18131 & w15027) | (w18131 & w36095) | (w15027 & w36095);
assign w18133 = ~w18124 & ~w18132;
assign w18134 = w18123 & w18133;
assign w18135 = ~w18121 & ~w18134;
assign w18136 = ~w18120 & w18135;
assign w18137 = ~w18123 & ~w18133;
assign w18138 = (~w17856 & ~w17841) | (~w17856 & w31905) | (~w17841 & w31905);
assign w18139 = ~w17668 & ~w17860;
assign w18140 = w6996 & ~w12661;
assign w18141 = w6998 & ~w12637;
assign w18142 = w6446 & w12646;
assign w18143 = ~w18141 & ~w18142;
assign w18144 = ~w18140 & w18143;
assign w18145 = (w18144 & w14641) | (w18144 & w36096) | (w14641 & w36096);
assign w18146 = ~a_14 & w18145;
assign w18147 = (~w14641 & w36097) | (~w14641 & w36098) | (w36097 & w36098);
assign w18148 = ~w18146 & ~w18147;
assign w18149 = ~w18139 & ~w18148;
assign w18150 = w18138 & w18149;
assign w18151 = w18139 & ~w18148;
assign w18152 = ~w18138 & w18151;
assign w18153 = ~w18150 & ~w18152;
assign w18154 = ~w18137 & w18153;
assign w18155 = ~w18136 & w18154;
assign w18156 = w18139 & w18148;
assign w18157 = w18138 & w18156;
assign w18158 = ~w18139 & w18148;
assign w18159 = ~w18138 & w18158;
assign w18160 = ~w18157 & ~w18159;
assign w18161 = ~w17880 & w17893;
assign w18162 = w17862 & w18161;
assign w18163 = w17880 & w17893;
assign w18164 = ~w17862 & w18163;
assign w18165 = ~w18162 & ~w18164;
assign w18166 = w18160 & w18165;
assign w18167 = ~w18155 & w18166;
assign w18168 = ~w17894 & ~w18167;
assign w18169 = w17874 & ~w17880;
assign w18170 = ~w17881 & ~w18169;
assign w18171 = ~w17444 & ~w17461;
assign w18172 = ~w17462 & ~w18171;
assign w18173 = w8391 & ~w15027;
assign w18174 = w6304 & ~w12637;
assign w18175 = w6059 & w12651;
assign w18176 = w6061 & w12646;
assign w18177 = ~w18174 & w36099;
assign w18178 = a_17 & w18177;
assign w18179 = ~a_17 & ~w18177;
assign w18180 = ~w18178 & ~w18179;
assign w18181 = (w18180 & w15027) | (w18180 & w36100) | (w15027 & w36100);
assign w18182 = ~w18173 & ~w18181;
assign w18183 = w18172 & w18182;
assign w18184 = ~w18172 & ~w18182;
assign w18185 = ~w18183 & ~w18184;
assign w18186 = w8564 & ~w14535;
assign w18187 = w6998 & ~w12668;
assign w18188 = w6446 & ~w12661;
assign w18189 = w6996 & ~w12630;
assign w18190 = ~w18187 & ~w18188;
assign w18191 = (~a_14 & ~w18190) | (~a_14 & w36101) | (~w18190 & w36101);
assign w18192 = w18190 & w36102;
assign w18193 = ~w18191 & ~w18192;
assign w18194 = (w18193 & w14535) | (w18193 & w36103) | (w14535 & w36103);
assign w18195 = ~w18186 & ~w18194;
assign w18196 = w18185 & ~w18195;
assign w18197 = ~w18185 & w18195;
assign w18198 = ~w18196 & ~w18197;
assign w18199 = w18170 & ~w18198;
assign w18200 = ~w18170 & w18198;
assign w18201 = ~w18199 & ~w18200;
assign w18202 = w18168 & ~w18201;
assign w18203 = w18170 & ~w18185;
assign w18204 = w18195 & ~w18203;
assign w18205 = ~w18200 & w18204;
assign w18206 = ~w18169 & ~w18183;
assign w18207 = ~w17881 & w18206;
assign w18208 = (~w18184 & ~w18206) | (~w18184 & w31906) | (~w18206 & w31906);
assign w18209 = (~w17459 & ~w17444) | (~w17459 & w31907) | (~w17444 & w31907);
assign w18210 = ~w17272 & ~w17463;
assign w18211 = w6304 & ~w12661;
assign w18212 = w6061 & ~w12637;
assign w18213 = w6059 & w12646;
assign w18214 = ~w18212 & ~w18213;
assign w18215 = ~w18211 & w18214;
assign w18216 = (w18215 & w14641) | (w18215 & w36104) | (w14641 & w36104);
assign w18217 = ~a_17 & w18216;
assign w18218 = (~w14641 & w36105) | (~w14641 & w36106) | (w36105 & w36106);
assign w18219 = ~w18217 & ~w18218;
assign w18220 = w18210 & ~w18219;
assign w18221 = ~w18210 & w18219;
assign w18222 = ~w18220 & ~w18221;
assign w18223 = ~w18209 & w18222;
assign w18224 = w18209 & ~w18222;
assign w18225 = ~w18223 & ~w18224;
assign w18226 = w8564 & ~w14412;
assign w18227 = w6998 & ~w12630;
assign w18228 = w6446 & ~w12668;
assign w18229 = w6996 & w12622;
assign w18230 = ~w18227 & ~w18228;
assign w18231 = w18230 & w36107;
assign w18232 = (~a_14 & ~w18230) | (~a_14 & w36108) | (~w18230 & w36108);
assign w18233 = ~w18231 & ~w18232;
assign w18234 = (w18233 & w14412) | (w18233 & w36109) | (w14412 & w36109);
assign w18235 = ~w18226 & ~w18234;
assign w18236 = w18225 & w18235;
assign w18237 = w18208 & w18236;
assign w18238 = ~w18225 & w18235;
assign w18239 = ~w18208 & w18238;
assign w18240 = ~w18237 & ~w18239;
assign w18241 = ~w18205 & w18240;
assign w18242 = ~w18202 & w18241;
assign w18243 = w18208 & ~w18225;
assign w18244 = ~w18208 & w18225;
assign w18245 = ~w18243 & ~w18244;
assign w18246 = ~w18235 & ~w18245;
assign w18247 = w18209 & ~w18210;
assign w18248 = w18219 & ~w18247;
assign w18249 = ~w18223 & w18248;
assign w18250 = ~w18219 & w18247;
assign w18251 = ~w18209 & w18220;
assign w18252 = ~w18184 & ~w18251;
assign w18253 = ~w18250 & w18252;
assign w18254 = ~w18207 & w18253;
assign w18255 = ~w18249 & ~w18254;
assign w18256 = w6996 & w12856;
assign w18257 = w6998 & w12622;
assign w18258 = w6446 & ~w12630;
assign w18259 = ~w18257 & ~w18258;
assign w18260 = ~w18256 & w18259;
assign w18261 = (w18260 & ~w14091) | (w18260 & w36110) | (~w14091 & w36110);
assign w18262 = a_14 & ~w18261;
assign w18263 = (~w14091 & w36111) | (~w14091 & w36112) | (w36111 & w36112);
assign w18264 = ~w18262 & ~w18263;
assign w18265 = w8391 & w14393;
assign w18266 = w6061 & ~w12661;
assign w18267 = w6059 & ~w12637;
assign w18268 = w6304 & ~w12668;
assign w18269 = ~w18266 & ~w18267;
assign w18270 = w18269 & w36113;
assign w18271 = (~a_17 & ~w18269) | (~a_17 & w36114) | (~w18269 & w36114);
assign w18272 = ~w18270 & ~w18271;
assign w18273 = (w18272 & ~w14393) | (w18272 & w36115) | (~w14393 & w36115);
assign w18274 = ~w18265 & ~w18273;
assign w18275 = w17484 & w18274;
assign w18276 = w17466 & w18275;
assign w18277 = ~w17484 & w18274;
assign w18278 = ~w17466 & w18277;
assign w18279 = ~w18276 & ~w18278;
assign w18280 = ~w17484 & ~w18274;
assign w18281 = w17466 & w18280;
assign w18282 = w17484 & ~w18274;
assign w18283 = ~w17466 & w18282;
assign w18284 = ~w18281 & ~w18283;
assign w18285 = w18279 & w18284;
assign w18286 = ~w18264 & ~w18285;
assign w18287 = w18255 & ~w18286;
assign w18288 = ~w18264 & w18285;
assign w18289 = ~w18255 & ~w18288;
assign w18290 = ~w18287 & ~w18289;
assign w18291 = ~w18246 & ~w18290;
assign w18292 = ~w18242 & w18291;
assign w18293 = w18264 & ~w18285;
assign w18294 = ~w18288 & ~w18293;
assign w18295 = w18255 & ~w18294;
assign w18296 = ~w18287 & ~w18293;
assign w18297 = ~w18295 & ~w18296;
assign w18298 = ~w18292 & ~w18297;
assign w18299 = ~w18249 & w18279;
assign w18300 = ~w18254 & w18299;
assign w18301 = w18284 & ~w18300;
assign w18302 = w8564 & w14442;
assign w18303 = w6998 & w12856;
assign w18304 = w6446 & w12622;
assign w18305 = w6996 & ~w12860;
assign w18306 = ~w18303 & ~w18304;
assign w18307 = ~w18305 & w36116;
assign w18308 = (~a_14 & w18305) | (~a_14 & w36117) | (w18305 & w36117);
assign w18309 = ~w18307 & ~w18308;
assign w18310 = (w18309 & ~w14442) | (w18309 & w36118) | (~w14442 & w36118);
assign w18311 = ~w18302 & ~w18310;
assign w18312 = w17467 & w17479;
assign w18313 = w17468 & ~w17478;
assign w18314 = ~w17467 & w18313;
assign w18315 = ~w17272 & ~w18312;
assign w18316 = ~w18314 & w18315;
assign w18317 = ~w17465 & w18316;
assign w18318 = ~w17486 & ~w18317;
assign w18319 = w8391 & ~w14535;
assign w18320 = ~w14391 & w36119;
assign w18321 = w8419 & ~w14532;
assign w18322 = w6061 & ~w12668;
assign w18323 = w6059 & ~w12661;
assign w18324 = w6304 & ~w12630;
assign w18325 = ~w18322 & ~w18323;
assign w18326 = (a_17 & ~w18325) | (a_17 & w36121) | (~w18325 & w36121);
assign w18327 = w18325 & w36122;
assign w18328 = ~w18326 & ~w18327;
assign w18329 = (~w14391 & w36123) | (~w14391 & w36124) | (w36123 & w36124);
assign w18330 = ~w18320 & w18329;
assign w18331 = ~w18319 & ~w18330;
assign w18332 = w17498 & ~w18331;
assign w18333 = ~w17498 & w18331;
assign w18334 = ~w18332 & ~w18333;
assign w18335 = w17488 & ~w18334;
assign w18336 = ~w17488 & w18334;
assign w18337 = ~w18335 & ~w18336;
assign w18338 = w18318 & w18337;
assign w18339 = ~w18318 & ~w18337;
assign w18340 = ~w18338 & ~w18339;
assign w18341 = ~w18311 & w18340;
assign w18342 = w18301 & w18341;
assign w18343 = ~w18311 & ~w18340;
assign w18344 = ~w18301 & w18343;
assign w18345 = ~w18342 & ~w18344;
assign w18346 = w18311 & ~w18340;
assign w18347 = w18301 & w18346;
assign w18348 = w18311 & w18340;
assign w18349 = ~w18301 & w18348;
assign w18350 = ~w18347 & ~w18349;
assign w18351 = w18345 & w18350;
assign w18352 = ~w17655 & ~w18351;
assign w18353 = w17655 & w18351;
assign w18354 = ~w18352 & ~w18353;
assign w18355 = w18298 & w18354;
assign w18356 = ~w18298 & ~w18354;
assign w18357 = ~w18355 & ~w18356;
assign w18358 = w17655 & w18357;
assign w18359 = ~w18058 & ~w18075;
assign w18360 = ~w18076 & ~w18359;
assign w18361 = w9061 & w14614;
assign w18362 = w7511 & w12651;
assign w18363 = w7192 & w12793;
assign w18364 = w7489 & ~w12830;
assign w18365 = ~w18362 & ~w18363;
assign w18366 = ~w18364 & w36125;
assign w18367 = (~a_11 & w18364) | (~a_11 & w36126) | (w18364 & w36126);
assign w18368 = ~w18366 & ~w18367;
assign w18369 = (w18368 & ~w14614) | (w18368 & w36127) | (~w14614 & w36127);
assign w18370 = ~w18361 & ~w18369;
assign w18371 = ~w18360 & ~w18370;
assign w18372 = w18033 & ~w18050;
assign w18373 = ~w18051 & ~w18372;
assign w18374 = w9061 & ~w15101;
assign w18375 = w7489 & w12789;
assign w18376 = ~w12770 & w36128;
assign w18377 = w7511 & w12793;
assign w18378 = ~w18375 & ~w18376;
assign w18379 = (~a_11 & ~w18378) | (~a_11 & w36129) | (~w18378 & w36129);
assign w18380 = w18378 & w36130;
assign w18381 = ~w18379 & ~w18380;
assign w18382 = (w18381 & w15101) | (w18381 & w36131) | (w15101 & w36131);
assign w18383 = ~w18374 & ~w18382;
assign w18384 = ~w18373 & ~w18383;
assign w18385 = ~w18012 & ~w18013;
assign w18386 = ~w18030 & w18385;
assign w18387 = w18030 & ~w18385;
assign w18388 = ~w18386 & ~w18387;
assign w18389 = ~w12770 & w31908;
assign w18390 = w7192 & w12732;
assign w18391 = w7489 & ~w12774;
assign w18392 = ~w18389 & ~w18390;
assign w18393 = (~a_11 & ~w18392) | (~a_11 & w36132) | (~w18392 & w36132);
assign w18394 = w18392 & w36133;
assign w18395 = ~w18393 & ~w18394;
assign w18396 = ~w15435 & w18395;
assign w18397 = (~a_11 & ~w7187) | (~a_11 & w36134) | (~w7187 & w36134);
assign w18398 = ~w9061 & ~w18397;
assign w18399 = w18392 & w36135;
assign w18400 = ~w18393 & ~w18399;
assign w18401 = w15435 & w18400;
assign w18402 = ~w18396 & ~w18401;
assign w18403 = w18388 & ~w18402;
assign w18404 = w12679 & w36136;
assign w18405 = w17988 & ~w18404;
assign w18406 = (a_14 & ~w17988) | (a_14 & w36137) | (~w17988 & w36137);
assign w18407 = ~w17982 & w18406;
assign w18408 = w17982 & ~w18406;
assign w18409 = ~w18407 & ~w18408;
assign w18410 = w7192 & w12701;
assign w18411 = w7511 & w12732;
assign w18412 = (~w18410 & ~w12739) | (~w18410 & w36138) | (~w12739 & w36138);
assign w18413 = ~w18411 & w18412;
assign w18414 = a_11 & w18413;
assign w18415 = w18409 & w18414;
assign w18416 = (w18415 & w15977) | (w18415 & w36139) | (w15977 & w36139);
assign w18417 = w9089 & w18409;
assign w18418 = ~a_11 & ~w18413;
assign w18419 = w18409 & w18418;
assign w18420 = (~w18419 & w15977) | (~w18419 & w36140) | (w15977 & w36140);
assign w18421 = ~w18416 & w18420;
assign w18422 = ~a_11 & w18413;
assign w18423 = ~w18409 & w18422;
assign w18424 = (w18423 & w15977) | (w18423 & w36141) | (w15977 & w36141);
assign w18425 = w9061 & ~w18409;
assign w18426 = a_11 & ~w18413;
assign w18427 = ~w18409 & w18426;
assign w18428 = (~w18427 & w15977) | (~w18427 & w36142) | (w15977 & w36142);
assign w18429 = ~w18424 & w18428;
assign w18430 = ~w17988 & w18404;
assign w18431 = ~w18405 & ~w18430;
assign w18432 = w12702 & w31909;
assign w18433 = w7193 & w15385;
assign w18434 = ~w12702 & w18433;
assign w18435 = w7511 & ~w12675;
assign w18436 = ~w12674 & w18435;
assign w18437 = w7192 & w12679;
assign w18438 = w7511 & w11683;
assign w18439 = w11678 & w18438;
assign w18440 = w7489 & ~w11501;
assign w18441 = w12684 & w18440;
assign w18442 = ~w18436 & ~w18437;
assign w18443 = ~w18439 & ~w18441;
assign w18444 = w18442 & w18443;
assign w18445 = ~w18434 & w18444;
assign w18446 = ~w18432 & w18445;
assign w18447 = w7187 & w12679;
assign w18448 = w12684 & w31910;
assign w18449 = w7489 & w12679;
assign w18450 = w7193 & ~w15324;
assign w18451 = ~w18448 & ~w18449;
assign w18452 = ~w18450 & w18451;
assign w18453 = (a_11 & ~w12679) | (a_11 & w36143) | (~w12679 & w36143);
assign w18454 = w18452 & w18453;
assign w18455 = (~w17983 & ~w18446) | (~w17983 & w31911) | (~w18446 & w31911);
assign w18456 = w7193 & w15283;
assign w18457 = w7193 & ~w12681;
assign w18458 = w12688 & w18457;
assign w18459 = ~w15282 & w18458;
assign w18460 = w7511 & ~w11825;
assign w18461 = ~w12699 & w18460;
assign w18462 = w11825 & w18438;
assign w18463 = ~w11678 & w18462;
assign w18464 = w15293 & w18440;
assign w18465 = ~w12674 & w31912;
assign w18466 = w12684 & w36144;
assign w18467 = ~w18463 & ~w18464;
assign w18468 = ~w18461 & w18467;
assign w18469 = ~w18465 & ~w18466;
assign w18470 = w18468 & w18469;
assign w18471 = ~w18459 & w18470;
assign w18472 = ~w18456 & w18471;
assign w18473 = a_11 & ~w18472;
assign w18474 = ~a_11 & w18472;
assign w18475 = ~w18473 & ~w18474;
assign w18476 = w18475 & w31913;
assign w18477 = (~w18431 & ~w18475) | (~w18431 & w31914) | (~w18475 & w31914);
assign w18478 = w7193 & w12715;
assign w18479 = w7511 & w12739;
assign w18480 = w7192 & w12702;
assign w18481 = w7489 & w12701;
assign w18482 = w7193 & ~w12700;
assign w18483 = w12711 & ~w18482;
assign w18484 = w7193 & w12700;
assign w18485 = ~w12711 & ~w18484;
assign w18486 = ~w18483 & ~w18485;
assign w18487 = ~w12704 & w18486;
assign w18488 = ~w18480 & ~w18481;
assign w18489 = ~w18479 & w18488;
assign w18490 = ~w18487 & w18489;
assign w18491 = ~w18478 & w18490;
assign w18492 = a_11 & ~w18491;
assign w18493 = ~a_11 & w18491;
assign w18494 = ~w18492 & ~w18493;
assign w18495 = (~w18476 & ~w18494) | (~w18476 & w31915) | (~w18494 & w31915);
assign w18496 = w18429 & ~w18495;
assign w18497 = w18421 & ~w18496;
assign w18498 = w7489 & w12732;
assign w18499 = w7192 & w12739;
assign w18500 = w7511 & ~w12774;
assign w18501 = ~w18498 & ~w18499;
assign w18502 = ~w18500 & w18501;
assign w18503 = (w18502 & w15157) | (w18502 & w36145) | (w15157 & w36145);
assign w18504 = w17982 & w31916;
assign w18505 = ~w17991 & ~w18504;
assign w18506 = w18011 & w18505;
assign w18507 = ~w18011 & ~w18505;
assign w18508 = ~w18506 & ~w18507;
assign w18509 = ~a_11 & w18508;
assign w18510 = a_11 & ~w18508;
assign w18511 = ~w18509 & ~w18510;
assign w18512 = w18503 & w18511;
assign w18513 = ~w18503 & ~w18511;
assign w18514 = ~w18512 & ~w18513;
assign w18515 = ~w18497 & w18514;
assign w18516 = ~w18388 & w18402;
assign w18517 = ~w18503 & ~w18509;
assign w18518 = a_11 & w18508;
assign w18519 = w18503 & ~w18518;
assign w18520 = ~w18517 & ~w18519;
assign w18521 = ~w18516 & ~w18520;
assign w18522 = (~w18403 & w18515) | (~w18403 & w31917) | (w18515 & w31917);
assign w18523 = w7192 & ~w12774;
assign w18524 = w7511 & w12789;
assign w18525 = ~w12770 & w36146;
assign w18526 = ~w18524 & w36147;
assign w18527 = ~w7193 & w18526;
assign w18528 = ~w15127 & w18526;
assign w18529 = (~w18527 & ~w18528) | (~w18527 & w31918) | (~w18528 & w31918);
assign w18530 = ~a_11 & w18529;
assign w18531 = a_11 & ~w18529;
assign w18532 = ~w18530 & ~w18531;
assign w18533 = w17957 & w17965;
assign w18534 = ~w18031 & w18533;
assign w18535 = w18031 & ~w18533;
assign w18536 = ~w18534 & ~w18535;
assign w18537 = ~w18532 & ~w18536;
assign w18538 = w18532 & w18536;
assign w18539 = ~w18537 & ~w18538;
assign w18540 = w18522 & w18539;
assign w18541 = w18373 & w18383;
assign w18542 = (~w18537 & ~w18373) | (~w18537 & w36148) | (~w18373 & w36148);
assign w18543 = ~w18540 & w18542;
assign w18544 = ~w18384 & ~w18543;
assign w18545 = w9061 & w15071;
assign w18546 = w7489 & w12793;
assign w18547 = w7192 & w12789;
assign w18548 = w7511 & ~w12830;
assign w18549 = ~w18546 & ~w18547;
assign w18550 = (~a_11 & w18548) | (~a_11 & w36149) | (w18548 & w36149);
assign w18551 = ~w18548 & w36150;
assign w18552 = ~w18550 & ~w18551;
assign w18553 = (w18552 & ~w15071) | (w18552 & w36151) | (~w15071 & w36151);
assign w18554 = ~w18545 & ~w18553;
assign w18555 = ~w17939 & ~w18052;
assign w18556 = ~w18051 & w31919;
assign w18557 = (~w18555 & w18051) | (~w18555 & w31920) | (w18051 & w31920);
assign w18558 = ~w18556 & ~w18557;
assign w18559 = w18554 & ~w18558;
assign w18560 = ~w18554 & w18558;
assign w18561 = ~w18559 & ~w18560;
assign w18562 = w18544 & w18561;
assign w18563 = w18360 & w18370;
assign w18564 = (~w18559 & ~w18360) | (~w18559 & w31921) | (~w18360 & w31921);
assign w18565 = (~w18371 & w18562) | (~w18371 & w31922) | (w18562 & w31922);
assign w18566 = ~w18073 & ~w18076;
assign w18567 = ~w17920 & ~w18077;
assign w18568 = ~w15044 & w36152;
assign w18569 = ~w15044 & w36153;
assign w18570 = w7511 & w12646;
assign w18571 = w7489 & w12651;
assign w18572 = (~w18570 & w12830) | (~w18570 & w36154) | (w12830 & w36154);
assign w18573 = (~a_11 & ~w18572) | (~a_11 & w36155) | (~w18572 & w36155);
assign w18574 = w18572 & w36156;
assign w18575 = ~w18573 & ~w18574;
assign w18576 = ~w18569 & w18575;
assign w18577 = ~w18568 & ~w18576;
assign w18578 = w18567 & ~w18577;
assign w18579 = ~w18567 & w18577;
assign w18580 = ~w18578 & ~w18579;
assign w18581 = w18566 & w18580;
assign w18582 = ~w18566 & ~w18580;
assign w18583 = ~w18581 & ~w18582;
assign w18584 = w18565 & w18583;
assign w18585 = w18577 & ~w18583;
assign w18586 = ~w18080 & ~w18097;
assign w18587 = ~w18098 & ~w18586;
assign w18588 = w9061 & ~w15027;
assign w18589 = w7511 & ~w12637;
assign w18590 = w7192 & w12651;
assign w18591 = w7489 & w12646;
assign w18592 = ~w18589 & w36157;
assign w18593 = a_11 & w18592;
assign w18594 = ~a_11 & ~w18592;
assign w18595 = ~w18593 & ~w18594;
assign w18596 = (w18595 & w15027) | (w18595 & w36158) | (w15027 & w36158);
assign w18597 = ~w18588 & ~w18596;
assign w18598 = w18587 & w18597;
assign w18599 = ~w18585 & ~w18598;
assign w18600 = ~w18584 & w18599;
assign w18601 = ~w18587 & ~w18597;
assign w18602 = (~w18095 & ~w18080) | (~w18095 & w31923) | (~w18080 & w31923);
assign w18603 = ~w17907 & ~w18099;
assign w18604 = w7511 & ~w12661;
assign w18605 = w7489 & ~w12637;
assign w18606 = w7192 & w12646;
assign w18607 = ~w18605 & ~w18606;
assign w18608 = ~w18604 & w18607;
assign w18609 = (w18608 & w14641) | (w18608 & w36159) | (w14641 & w36159);
assign w18610 = ~a_11 & w18609;
assign w18611 = (~w14641 & w36160) | (~w14641 & w36161) | (w36160 & w36161);
assign w18612 = ~w18610 & ~w18611;
assign w18613 = ~w18603 & ~w18612;
assign w18614 = w18602 & w18613;
assign w18615 = w18603 & ~w18612;
assign w18616 = ~w18602 & w18615;
assign w18617 = ~w18614 & ~w18616;
assign w18618 = ~w18601 & w18617;
assign w18619 = ~w18600 & w18618;
assign w18620 = w18603 & w18612;
assign w18621 = w18602 & w18620;
assign w18622 = ~w18603 & w18612;
assign w18623 = ~w18602 & w18622;
assign w18624 = ~w18621 & ~w18623;
assign w18625 = w9061 & w14393;
assign w18626 = w7489 & ~w12661;
assign w18627 = w7192 & ~w12637;
assign w18628 = w7511 & ~w12668;
assign w18629 = ~w18626 & ~w18627;
assign w18630 = w18629 & w36162;
assign w18631 = (~a_11 & ~w18629) | (~a_11 & w36163) | (~w18629 & w36163);
assign w18632 = ~w18630 & ~w18631;
assign w18633 = (w18632 & ~w14393) | (w18632 & w36164) | (~w14393 & w36164);
assign w18634 = ~w18625 & ~w18633;
assign w18635 = ~w18119 & w18634;
assign w18636 = w18101 & w18635;
assign w18637 = w18119 & w18634;
assign w18638 = ~w18101 & w18637;
assign w18639 = ~w18636 & ~w18638;
assign w18640 = w18624 & w18639;
assign w18641 = ~w18619 & w18640;
assign w18642 = w18119 & ~w18634;
assign w18643 = w18101 & w18642;
assign w18644 = ~w18119 & ~w18634;
assign w18645 = ~w18101 & w18644;
assign w18646 = ~w18643 & ~w18645;
assign w18647 = ~w18641 & w18646;
assign w18648 = ~w18120 & ~w18121;
assign w18649 = ~w18134 & ~w18137;
assign w18650 = w9061 & ~w14535;
assign w18651 = w7489 & ~w12668;
assign w18652 = w7192 & ~w12661;
assign w18653 = w7511 & ~w12630;
assign w18654 = ~w18651 & ~w18652;
assign w18655 = (~a_11 & ~w18654) | (~a_11 & w36165) | (~w18654 & w36165);
assign w18656 = w18654 & w36166;
assign w18657 = ~w18655 & ~w18656;
assign w18658 = (w18657 & w14535) | (w18657 & w36167) | (w14535 & w36167);
assign w18659 = ~w18650 & ~w18658;
assign w18660 = w18649 & ~w18659;
assign w18661 = ~w18649 & w18659;
assign w18662 = ~w18660 & ~w18661;
assign w18663 = w18648 & ~w18662;
assign w18664 = ~w18648 & w18662;
assign w18665 = ~w18663 & ~w18664;
assign w18666 = w18647 & ~w18665;
assign w18667 = (w18659 & ~w18648) | (w18659 & w36168) | (~w18648 & w36168);
assign w18668 = ~w18664 & w18667;
assign w18669 = (~w18137 & ~w18135) | (~w18137 & w31924) | (~w18135 & w31924);
assign w18670 = w18153 & w18160;
assign w18671 = w9061 & ~w14412;
assign w18672 = w7489 & ~w12630;
assign w18673 = w7192 & ~w12668;
assign w18674 = w7511 & w12622;
assign w18675 = ~w18672 & ~w18673;
assign w18676 = w18675 & w36169;
assign w18677 = (~a_11 & ~w18675) | (~a_11 & w36170) | (~w18675 & w36170);
assign w18678 = ~w18676 & ~w18677;
assign w18679 = (w18678 & w14412) | (w18678 & w36171) | (w14412 & w36171);
assign w18680 = ~w18671 & ~w18679;
assign w18681 = ~w18670 & w18680;
assign w18682 = w18669 & w18681;
assign w18683 = w18670 & w18680;
assign w18684 = ~w18669 & w18683;
assign w18685 = ~w18682 & ~w18684;
assign w18686 = ~w18668 & w18685;
assign w18687 = ~w18666 & w18686;
assign w18688 = ~w18669 & w18670;
assign w18689 = w18669 & ~w18670;
assign w18690 = ~w18688 & ~w18689;
assign w18691 = ~w18680 & w18690;
assign w18692 = (w18160 & w18136) | (w18160 & w37570) | (w18136 & w37570);
assign w18693 = w7489 & w12622;
assign w18694 = w7192 & ~w12630;
assign w18695 = w7511 & w12856;
assign w18696 = ~w18693 & ~w18694;
assign w18697 = (a_11 & ~w18696) | (a_11 & w36172) | (~w18696 & w36172);
assign w18698 = w7193 & w14091;
assign w18699 = w18696 & w36173;
assign w18700 = ~w18698 & w18699;
assign w18701 = (~w18697 & ~w14091) | (~w18697 & w36174) | (~w14091 & w36174);
assign w18702 = ~w18700 & w18701;
assign w18703 = (w17893 & w18700) | (w17893 & w36175) | (w18700 & w36175);
assign w18704 = ~w18700 & w36176;
assign w18705 = ~w18703 & ~w18704;
assign w18706 = w17883 & ~w18705;
assign w18707 = ~w17883 & w18705;
assign w18708 = ~w18706 & ~w18707;
assign w18709 = w18692 & w18708;
assign w18710 = ~w18692 & ~w18708;
assign w18711 = ~w18709 & ~w18710;
assign w18712 = ~w18691 & ~w18711;
assign w18713 = ~w18687 & w18712;
assign w18714 = w9061 & w14442;
assign w18715 = w7489 & w12856;
assign w18716 = w7192 & w12622;
assign w18717 = w7511 & ~w12860;
assign w18718 = ~w18715 & ~w18716;
assign w18719 = ~w18717 & w36177;
assign w18720 = (~a_11 & w18717) | (~a_11 & w36178) | (w18717 & w36178);
assign w18721 = ~w18719 & ~w18720;
assign w18722 = (w18721 & ~w14442) | (w18721 & w36179) | (~w14442 & w36179);
assign w18723 = ~w18714 & ~w18722;
assign w18724 = w18170 & w18723;
assign w18725 = w18198 & ~w18724;
assign w18726 = ~w18170 & w18723;
assign w18727 = ~w18198 & ~w18726;
assign w18728 = ~w18725 & ~w18727;
assign w18729 = w18168 & ~w18728;
assign w18730 = w18198 & ~w18726;
assign w18731 = ~w18198 & ~w18724;
assign w18732 = ~w18730 & ~w18731;
assign w18733 = ~w18168 & ~w18732;
assign w18734 = ~w18729 & ~w18733;
assign w18735 = ~w17894 & w18165;
assign w18736 = ~w18692 & ~w18735;
assign w18737 = w18692 & w18735;
assign w18738 = ~w18736 & ~w18737;
assign w18739 = w18702 & ~w18738;
assign w18740 = ~w18734 & ~w18739;
assign w18741 = ~w18713 & w18740;
assign w18742 = w18170 & ~w18723;
assign w18743 = w18198 & ~w18742;
assign w18744 = ~w18170 & ~w18723;
assign w18745 = ~w18198 & ~w18744;
assign w18746 = ~w18743 & ~w18745;
assign w18747 = ~w18168 & w18746;
assign w18748 = w18198 & ~w18744;
assign w18749 = ~w18198 & ~w18742;
assign w18750 = ~w18748 & ~w18749;
assign w18751 = w18168 & w18750;
assign w18752 = ~w18747 & ~w18751;
assign w18753 = ~w18741 & w18752;
assign w18754 = (~w18205 & ~w18168) | (~w18205 & w37571) | (~w18168 & w37571);
assign w18755 = w9061 & w13979;
assign w18756 = w7511 & w12869;
assign w18757 = w7192 & w12856;
assign w18758 = w7489 & ~w12860;
assign w18759 = ~w18756 & ~w18757;
assign w18760 = ~w18758 & w18759;
assign w18761 = a_11 & ~w18760;
assign w18762 = ~a_11 & w18760;
assign w18763 = (w18762 & ~w13979) | (w18762 & w36180) | (~w13979 & w36180);
assign w18764 = ~w18755 & ~w18761;
assign w18765 = ~w18763 & w18764;
assign w18766 = (w18235 & ~w18764) | (w18235 & w36181) | (~w18764 & w36181);
assign w18767 = w18764 & w36182;
assign w18768 = ~w18766 & ~w18767;
assign w18769 = w18245 & ~w18768;
assign w18770 = ~w18245 & w18768;
assign w18771 = ~w18769 & ~w18770;
assign w18772 = w18754 & w18771;
assign w18773 = ~w18754 & ~w18771;
assign w18774 = ~w18772 & ~w18773;
assign w18775 = ~w18741 & w37572;
assign w18776 = w18765 & w18774;
assign w18777 = ~w18242 & ~w18246;
assign w18778 = w7511 & w12874;
assign w18779 = w7192 & ~w12860;
assign w18780 = w7489 & w12869;
assign w18781 = w7193 & w13965;
assign w18782 = ~w18779 & w36183;
assign w18783 = (a_11 & w18781) | (a_11 & w36184) | (w18781 & w36184);
assign w18784 = ~w18781 & w36185;
assign w18785 = ~w18783 & ~w18784;
assign w18786 = ~w18255 & w18294;
assign w18787 = ~w18295 & ~w18786;
assign w18788 = w18785 & w18787;
assign w18789 = w18777 & w18788;
assign w18790 = w18785 & ~w18787;
assign w18791 = ~w18777 & w18790;
assign w18792 = ~w18789 & ~w18791;
assign w18793 = ~w18776 & w18792;
assign w18794 = ~w18775 & w18793;
assign w18795 = w18298 & w18352;
assign w18796 = ~w17655 & w18351;
assign w18797 = ~w18298 & w18796;
assign w18798 = ~w18785 & ~w18787;
assign w18799 = w18777 & w18798;
assign w18800 = ~w18785 & w18787;
assign w18801 = ~w18777 & w18800;
assign w18802 = ~w18799 & ~w18801;
assign w18803 = ~w18795 & ~w18797;
assign w18804 = w18802 & w18803;
assign w18805 = ~w18794 & w18804;
assign w18806 = ~w18358 & ~w18805;
assign w18807 = ~w18297 & w18350;
assign w18808 = w18345 & ~w18807;
assign w18809 = w18345 & ~w18787;
assign w18810 = w18777 & w18809;
assign w18811 = ~w18808 & ~w18810;
assign w18812 = w6061 & ~w12630;
assign w18813 = w6059 & ~w12668;
assign w18814 = w6304 & w12622;
assign w18815 = ~w18812 & ~w18813;
assign w18816 = ~w18814 & w18815;
assign w18817 = (w18816 & w14412) | (w18816 & w36186) | (w14412 & w36186);
assign w18818 = a_17 & ~w18817;
assign w18819 = (w14412 & w36187) | (w14412 & w36188) | (w36187 & w36188);
assign w18820 = ~w18818 & ~w18819;
assign w18821 = w17503 & ~w17505;
assign w18822 = ~w17503 & w17505;
assign w18823 = ~w18821 & ~w18822;
assign w18824 = w18820 & w18823;
assign w18825 = ~w18820 & ~w18823;
assign w18826 = ~w18824 & ~w18825;
assign w18827 = w18331 & ~w18340;
assign w18828 = ~w17498 & ~w18331;
assign w18829 = w17488 & ~w18828;
assign w18830 = ~w17488 & ~w18332;
assign w18831 = ~w18829 & ~w18830;
assign w18832 = w18318 & w18831;
assign w18833 = (~w18331 & w17488) | (~w18331 & w18828) | (w17488 & w18828);
assign w18834 = ~w17502 & w18833;
assign w18835 = ~w18318 & w18834;
assign w18836 = w18284 & ~w18832;
assign w18837 = ~w18835 & w18836;
assign w18838 = ~w18300 & w18837;
assign w18839 = ~w18827 & ~w18838;
assign w18840 = w6446 & w12856;
assign w18841 = w6996 & w12869;
assign w18842 = (~w18840 & w12860) | (~w18840 & w36189) | (w12860 & w36189);
assign w18843 = ~w18841 & w18842;
assign w18844 = (w18843 & ~w13979) | (w18843 & w36190) | (~w13979 & w36190);
assign w18845 = a_14 & w18844;
assign w18846 = (w13979 & w36191) | (w13979 & w36192) | (w36191 & w36192);
assign w18847 = ~w18845 & ~w18846;
assign w18848 = ~w18838 & w31925;
assign w18849 = (w18847 & w18838) | (w18847 & w31926) | (w18838 & w31926);
assign w18850 = ~w18848 & ~w18849;
assign w18851 = w18826 & w18850;
assign w18852 = ~w18826 & ~w18850;
assign w18853 = ~w18851 & ~w18852;
assign w18854 = ~w18811 & ~w18853;
assign w18855 = w18811 & w18853;
assign w18856 = ~w18854 & ~w18855;
assign w18857 = ~w12892 & w36193;
assign w18858 = w7489 & ~w12878;
assign w18859 = w7192 & w12874;
assign w18860 = ~w18858 & ~w18859;
assign w18861 = ~w18857 & w18860;
assign w18862 = (w18861 & ~w13787) | (w18861 & w36194) | (~w13787 & w36194);
assign w18863 = a_11 & ~w18862;
assign w18864 = (~w13787 & w36195) | (~w13787 & w36196) | (w36195 & w36196);
assign w18865 = ~w18863 & ~w18864;
assign w18866 = w18856 & w18865;
assign w18867 = ~w18856 & ~w18865;
assign w18868 = ~w18866 & ~w18867;
assign w18869 = ~w18806 & w18868;
assign w18870 = w18806 & ~w18868;
assign w18871 = ~w18869 & ~w18870;
assign w18872 = w17646 & w18871;
assign w18873 = ~w17646 & ~w18871;
assign w18874 = ~w18872 & ~w18873;
assign w18875 = (w18802 & ~w18793) | (w18802 & w37573) | (~w18793 & w37573);
assign w18876 = ~w18357 & ~w18875;
assign w18877 = w18357 & w18875;
assign w18878 = ~w18876 & ~w18877;
assign w18879 = ~w12905 & w36197;
assign w18880 = ~w12892 & w36198;
assign w18881 = w8295 & ~w12910;
assign w18882 = w8278 & w13815;
assign w18883 = ~w18881 & w36199;
assign w18884 = ~w18882 & w36200;
assign w18885 = (a_8 & w18882) | (a_8 & w36201) | (w18882 & w36201);
assign w18886 = ~w18884 & ~w18885;
assign w18887 = w18878 & ~w18886;
assign w18888 = (~w18739 & w18687) | (~w18739 & w37574) | (w18687 & w37574);
assign w18889 = w8295 & ~w12878;
assign w18890 = w8298 & w12874;
assign w18891 = w8277 & w12869;
assign w18892 = ~w18890 & ~w18891;
assign w18893 = ~w18889 & w18892;
assign w18894 = (w18893 & ~w13771) | (w18893 & w36202) | (~w13771 & w36202);
assign w18895 = a_8 & ~w18894;
assign w18896 = (~w13771 & w36203) | (~w13771 & w36204) | (w36203 & w36204);
assign w18897 = ~w18895 & ~w18896;
assign w18898 = ~w18734 & w18752;
assign w18899 = w18897 & ~w18898;
assign w18900 = ~w18897 & w18898;
assign w18901 = ~w18899 & ~w18900;
assign w18902 = ~w18888 & w18901;
assign w18903 = (w18897 & ~w18888) | (w18897 & w31927) | (~w18888 & w31927);
assign w18904 = ~w18902 & w18903;
assign w18905 = ~w12892 & w36205;
assign w18906 = w8298 & ~w12878;
assign w18907 = w8277 & w12874;
assign w18908 = ~w18906 & ~w18907;
assign w18909 = ~w18905 & w18908;
assign w18910 = (w18909 & ~w13787) | (w18909 & w36206) | (~w13787 & w36206);
assign w18911 = a_8 & ~w18910;
assign w18912 = (~w13787 & w36207) | (~w13787 & w36208) | (w36207 & w36208);
assign w18913 = ~w18911 & ~w18912;
assign w18914 = w18774 & w18913;
assign w18915 = w18753 & w18914;
assign w18916 = ~w18774 & w18913;
assign w18917 = ~w18753 & w18916;
assign w18918 = ~w18915 & ~w18917;
assign w18919 = ~w18904 & w18918;
assign w18920 = ~w18774 & ~w18913;
assign w18921 = w18753 & w18920;
assign w18922 = w18774 & ~w18913;
assign w18923 = ~w18753 & w18922;
assign w18924 = ~w18921 & ~w18923;
assign w18925 = ~w18919 & w18924;
assign w18926 = w8295 & w12874;
assign w18927 = w8277 & ~w12860;
assign w18928 = w8298 & w12869;
assign w18929 = w8278 & w13965;
assign w18930 = ~w18927 & w36209;
assign w18931 = ~w18929 & w36210;
assign w18932 = (a_8 & w18929) | (a_8 & w36211) | (w18929 & w36211);
assign w18933 = ~w18931 & ~w18932;
assign w18934 = ~w18687 & w37575;
assign w18935 = (~w18691 & w18666) | (~w18691 & w37576) | (w18666 & w37576);
assign w18936 = w18711 & ~w18933;
assign w18937 = ~w18935 & w18936;
assign w18938 = ~w18934 & ~w18937;
assign w18939 = w9456 & w14442;
assign w18940 = w8298 & w12856;
assign w18941 = w8277 & w12622;
assign w18942 = w8295 & ~w12860;
assign w18943 = ~w18940 & ~w18941;
assign w18944 = ~w18942 & w36212;
assign w18945 = (~a_8 & w18942) | (~a_8 & w36213) | (w18942 & w36213);
assign w18946 = ~w18944 & ~w18945;
assign w18947 = (w18946 & ~w14442) | (w18946 & w36214) | (~w14442 & w36214);
assign w18948 = ~w18939 & ~w18947;
assign w18949 = w18648 & w18948;
assign w18950 = w18662 & ~w18949;
assign w18951 = ~w18648 & w18948;
assign w18952 = ~w18662 & ~w18951;
assign w18953 = ~w18950 & ~w18952;
assign w18954 = w18647 & w18953;
assign w18955 = w18662 & ~w18951;
assign w18956 = ~w18662 & ~w18949;
assign w18957 = ~w18955 & ~w18956;
assign w18958 = ~w18647 & w18957;
assign w18959 = ~w18954 & ~w18958;
assign w18960 = w8295 & w12856;
assign w18961 = w8298 & w12622;
assign w18962 = w8277 & ~w12630;
assign w18963 = ~w18961 & ~w18962;
assign w18964 = ~w18960 & w18963;
assign w18965 = (w18964 & ~w14091) | (w18964 & w36215) | (~w14091 & w36215);
assign w18966 = a_8 & ~w18965;
assign w18967 = (~w14091 & w36216) | (~w14091 & w36217) | (w36216 & w36217);
assign w18968 = ~w18966 & ~w18967;
assign w18969 = (w18624 & w18600) | (w18624 & w36218) | (w18600 & w36218);
assign w18970 = w18639 & w18646;
assign w18971 = ~w18969 & ~w18970;
assign w18972 = w18969 & w18970;
assign w18973 = ~w18971 & ~w18972;
assign w18974 = w18968 & ~w18973;
assign w18975 = w18959 & ~w18974;
assign w18976 = w18648 & ~w18948;
assign w18977 = w18662 & ~w18976;
assign w18978 = ~w18648 & ~w18948;
assign w18979 = ~w18662 & ~w18978;
assign w18980 = ~w18977 & ~w18979;
assign w18981 = ~w18647 & w18980;
assign w18982 = w18662 & ~w18978;
assign w18983 = ~w18662 & ~w18976;
assign w18984 = ~w18982 & ~w18983;
assign w18985 = w18647 & w18984;
assign w18986 = ~w18981 & ~w18985;
assign w18987 = ~w18975 & w18986;
assign w18988 = (~w18601 & ~w18599) | (~w18601 & w31928) | (~w18599 & w31928);
assign w18989 = w18617 & w18624;
assign w18990 = w18988 & ~w18989;
assign w18991 = ~w18988 & w18989;
assign w18992 = ~w18990 & ~w18991;
assign w18993 = w9456 & ~w14412;
assign w18994 = w8295 & w12622;
assign w18995 = w8277 & ~w12668;
assign w18996 = w8298 & ~w12630;
assign w18997 = ~w18994 & ~w18995;
assign w18998 = w18997 & w36219;
assign w18999 = (~a_8 & ~w18997) | (~a_8 & w36220) | (~w18997 & w36220);
assign w19000 = ~w18998 & ~w18999;
assign w19001 = (w19000 & w14412) | (w19000 & w36221) | (w14412 & w36221);
assign w19002 = ~w18993 & ~w19001;
assign w19003 = w18992 & ~w19002;
assign w19004 = w9456 & w14393;
assign w19005 = w8298 & ~w12661;
assign w19006 = w8277 & ~w12637;
assign w19007 = w8295 & ~w12668;
assign w19008 = ~w19005 & ~w19006;
assign w19009 = w19008 & w36222;
assign w19010 = (~a_8 & ~w19008) | (~a_8 & w36223) | (~w19008 & w36223);
assign w19011 = ~w19009 & ~w19010;
assign w19012 = (w19011 & ~w14393) | (w19011 & w36224) | (~w14393 & w36224);
assign w19013 = ~w19004 & ~w19012;
assign w19014 = w18583 & w19013;
assign w19015 = ~w18565 & w19014;
assign w19016 = ~w18583 & w19013;
assign w19017 = w18565 & w19016;
assign w19018 = ~w19015 & ~w19017;
assign w19019 = w18583 & ~w19013;
assign w19020 = ~w19016 & ~w19019;
assign w19021 = w18565 & w19020;
assign w19022 = ~w18565 & ~w19020;
assign w19023 = ~w19021 & ~w19022;
assign w19024 = w19018 & w19023;
assign w19025 = ~w18522 & ~w18539;
assign w19026 = ~w18540 & ~w19025;
assign w19027 = w9456 & w14614;
assign w19028 = w8295 & w12651;
assign w19029 = w8277 & w12793;
assign w19030 = w8298 & ~w12830;
assign w19031 = ~w19028 & ~w19029;
assign w19032 = ~w19030 & w36225;
assign w19033 = (~a_8 & w19030) | (~a_8 & w36226) | (w19030 & w36226);
assign w19034 = ~w19032 & ~w19033;
assign w19035 = (w19034 & ~w14614) | (w19034 & w36227) | (~w14614 & w36227);
assign w19036 = ~w19027 & ~w19035;
assign w19037 = ~w19026 & ~w19036;
assign w19038 = w18497 & ~w18514;
assign w19039 = ~w18515 & ~w19038;
assign w19040 = w9456 & ~w15101;
assign w19041 = w8298 & w12789;
assign w19042 = ~w12770 & w36228;
assign w19043 = w8295 & w12793;
assign w19044 = ~w19041 & ~w19042;
assign w19045 = (~a_8 & ~w19044) | (~a_8 & w36229) | (~w19044 & w36229);
assign w19046 = w19044 & w36230;
assign w19047 = ~w19045 & ~w19046;
assign w19048 = (w19047 & w15101) | (w19047 & w36231) | (w15101 & w36231);
assign w19049 = ~w19040 & ~w19048;
assign w19050 = ~w19039 & ~w19049;
assign w19051 = ~w18476 & ~w18477;
assign w19052 = w18494 & w19051;
assign w19053 = ~w18494 & ~w19051;
assign w19054 = ~w19052 & ~w19053;
assign w19055 = ~w12770 & w31929;
assign w19056 = w8277 & w12732;
assign w19057 = w8298 & ~w12774;
assign w19058 = ~w19055 & ~w19056;
assign w19059 = (~a_8 & ~w19058) | (~a_8 & w36232) | (~w19058 & w36232);
assign w19060 = w19058 & w36233;
assign w19061 = ~w19059 & ~w19060;
assign w19062 = ~w15435 & w19061;
assign w19063 = (~a_8 & w8272) | (~a_8 & w36234) | (w8272 & w36234);
assign w19064 = ~w9456 & ~w19063;
assign w19065 = w19058 & w36235;
assign w19066 = ~w19059 & ~w19065;
assign w19067 = w15435 & w19066;
assign w19068 = ~w19062 & ~w19067;
assign w19069 = ~w19054 & ~w19068;
assign w19070 = w12679 & w36236;
assign w19071 = w18452 & ~w19070;
assign w19072 = (a_11 & ~w18452) | (a_11 & w36237) | (~w18452 & w36237);
assign w19073 = ~w18446 & w19072;
assign w19074 = w18446 & ~w19072;
assign w19075 = ~w19073 & ~w19074;
assign w19076 = w8277 & w12701;
assign w19077 = w8295 & w12732;
assign w19078 = (~w19076 & ~w12739) | (~w19076 & w36238) | (~w12739 & w36238);
assign w19079 = ~w19077 & w19078;
assign w19080 = a_8 & w19079;
assign w19081 = w19075 & w19080;
assign w19082 = (w19081 & w15977) | (w19081 & w36239) | (w15977 & w36239);
assign w19083 = w9484 & w19075;
assign w19084 = ~a_8 & ~w19079;
assign w19085 = w19075 & w19084;
assign w19086 = (~w19085 & w15977) | (~w19085 & w36240) | (w15977 & w36240);
assign w19087 = ~w19082 & w19086;
assign w19088 = w12702 & w31930;
assign w19089 = w8278 & w15385;
assign w19090 = ~w12702 & w19089;
assign w19091 = w8277 & w12679;
assign w19092 = w8295 & w12675;
assign w19093 = w12674 & w19092;
assign w19094 = w8295 & ~w12675;
assign w19095 = ~w12674 & w19094;
assign w19096 = w8298 & ~w11501;
assign w19097 = w12684 & w19096;
assign w19098 = ~w19091 & ~w19093;
assign w19099 = ~w19095 & ~w19097;
assign w19100 = w19098 & w19099;
assign w19101 = ~w19090 & w19100;
assign w19102 = ~w19088 & w19101;
assign w19103 = w8298 & w12679;
assign w19104 = (~w19103 & w15324) | (~w19103 & w31931) | (w15324 & w31931);
assign w19105 = a_8 & ~w8272;
assign w19106 = w12679 & w19105;
assign w19107 = w12684 & w31932;
assign w19108 = ~w19106 & ~w19107;
assign w19109 = w19104 & w19108;
assign w19110 = a_8 & w19109;
assign w19111 = w19102 & w31933;
assign w19112 = (~w18447 & ~w19102) | (~w18447 & w31934) | (~w19102 & w31934);
assign w19113 = ~w19111 & ~w19112;
assign w19114 = w8278 & w15283;
assign w19115 = w8278 & ~w12681;
assign w19116 = w12688 & w19115;
assign w19117 = ~w15282 & w19116;
assign w19118 = w8295 & ~w11825;
assign w19119 = ~w12699 & w19118;
assign w19120 = w8298 & ~w12675;
assign w19121 = ~w12674 & w19120;
assign w19122 = w15293 & w19096;
assign w19123 = w8295 & w11825;
assign w19124 = w12699 & w19123;
assign w19125 = w12684 & w31935;
assign w19126 = ~w19121 & ~w19122;
assign w19127 = ~w19119 & w19126;
assign w19128 = ~w19124 & ~w19125;
assign w19129 = w19127 & w19128;
assign w19130 = ~w19117 & w19129;
assign w19131 = ~w19114 & w19130;
assign w19132 = a_8 & ~w19131;
assign w19133 = ~a_8 & w19131;
assign w19134 = ~w19132 & ~w19133;
assign w19135 = w19113 & w19134;
assign w19136 = (~w19111 & ~w19134) | (~w19111 & w31936) | (~w19134 & w31936);
assign w19137 = w8278 & w12715;
assign w19138 = w8295 & w12739;
assign w19139 = w8277 & w12702;
assign w19140 = w8298 & w12701;
assign w19141 = w8278 & ~w12700;
assign w19142 = w12711 & ~w19141;
assign w19143 = w8278 & w12700;
assign w19144 = ~w12711 & ~w19143;
assign w19145 = ~w19142 & ~w19144;
assign w19146 = ~w12704 & w19145;
assign w19147 = ~w19139 & ~w19140;
assign w19148 = ~w19138 & w19147;
assign w19149 = ~w19146 & w19148;
assign w19150 = ~w19137 & w19149;
assign w19151 = ~w18452 & w19070;
assign w19152 = ~w19071 & ~w19151;
assign w19153 = ~a_8 & ~w19152;
assign w19154 = w19150 & w19153;
assign w19155 = a_8 & ~w19152;
assign w19156 = ~w19150 & w19155;
assign w19157 = ~w19154 & ~w19156;
assign w19158 = ~w19136 & w19157;
assign w19159 = a_8 & w19152;
assign w19160 = w19150 & w19159;
assign w19161 = ~a_8 & w19152;
assign w19162 = ~w19150 & w19161;
assign w19163 = ~w19160 & ~w19162;
assign w19164 = ~w19158 & w19163;
assign w19165 = ~a_8 & w19079;
assign w19166 = ~w19075 & w19165;
assign w19167 = (w19166 & w15977) | (w19166 & w36241) | (w15977 & w36241);
assign w19168 = w9456 & ~w19075;
assign w19169 = a_8 & ~w19079;
assign w19170 = ~w19075 & w19169;
assign w19171 = (~w19170 & w15977) | (~w19170 & w36242) | (w15977 & w36242);
assign w19172 = ~w19167 & w19171;
assign w19173 = (w19087 & w19164) | (w19087 & w36243) | (w19164 & w36243);
assign w19174 = w8298 & w12732;
assign w19175 = w8277 & w12739;
assign w19176 = w8295 & ~w12774;
assign w19177 = ~w19174 & ~w19175;
assign w19178 = ~w19176 & w19177;
assign w19179 = (w19178 & w15157) | (w19178 & w36244) | (w15157 & w36244);
assign w19180 = w18446 & w31937;
assign w19181 = ~w18455 & ~w19180;
assign w19182 = w18475 & w19181;
assign w19183 = ~w18475 & ~w19181;
assign w19184 = ~w19182 & ~w19183;
assign w19185 = ~a_8 & w19184;
assign w19186 = a_8 & ~w19184;
assign w19187 = ~w19185 & ~w19186;
assign w19188 = w19179 & w19187;
assign w19189 = ~w19179 & ~w19187;
assign w19190 = ~w19188 & ~w19189;
assign w19191 = ~w19173 & w19190;
assign w19192 = w19054 & w19068;
assign w19193 = ~w19179 & ~w19185;
assign w19194 = a_8 & w19184;
assign w19195 = w19179 & ~w19194;
assign w19196 = ~w19193 & ~w19195;
assign w19197 = ~w19192 & ~w19196;
assign w19198 = (~w19069 & w19191) | (~w19069 & w31938) | (w19191 & w31938);
assign w19199 = w8277 & ~w12774;
assign w19200 = ~w12770 & w36245;
assign w19201 = w8295 & w12789;
assign w19202 = ~w19199 & ~w19200;
assign w19203 = ~w19201 & w19202;
assign w19204 = ~w8278 & w19203;
assign w19205 = ~w15127 & w19203;
assign w19206 = (~w19204 & ~w19205) | (~w19204 & w31939) | (~w19205 & w31939);
assign w19207 = ~a_8 & w19206;
assign w19208 = a_8 & ~w19206;
assign w19209 = ~w19207 & ~w19208;
assign w19210 = w18421 & w18429;
assign w19211 = ~w18495 & w19210;
assign w19212 = w18495 & ~w19210;
assign w19213 = ~w19211 & ~w19212;
assign w19214 = ~w19209 & w19213;
assign w19215 = w19209 & ~w19213;
assign w19216 = ~w19214 & ~w19215;
assign w19217 = w19198 & w19216;
assign w19218 = w19039 & w19049;
assign w19219 = (~w19214 & ~w19039) | (~w19214 & w36246) | (~w19039 & w36246);
assign w19220 = ~w19217 & w19219;
assign w19221 = ~w19050 & ~w19220;
assign w19222 = w9456 & w15071;
assign w19223 = w8298 & w12793;
assign w19224 = w8277 & w12789;
assign w19225 = w8295 & ~w12830;
assign w19226 = ~w19223 & ~w19224;
assign w19227 = (~a_8 & w19225) | (~a_8 & w36247) | (w19225 & w36247);
assign w19228 = ~w19225 & w36248;
assign w19229 = ~w19227 & ~w19228;
assign w19230 = (w19229 & ~w15071) | (w19229 & w36249) | (~w15071 & w36249);
assign w19231 = ~w19222 & ~w19230;
assign w19232 = ~w18403 & ~w18516;
assign w19233 = ~w18515 & w31940;
assign w19234 = (~w19232 & w18515) | (~w19232 & w31941) | (w18515 & w31941);
assign w19235 = ~w19233 & ~w19234;
assign w19236 = w19231 & ~w19235;
assign w19237 = ~w19231 & w19235;
assign w19238 = ~w19236 & ~w19237;
assign w19239 = w19221 & w19238;
assign w19240 = w19026 & w19036;
assign w19241 = (~w19236 & ~w19026) | (~w19236 & w31942) | (~w19026 & w31942);
assign w19242 = (~w19037 & w19239) | (~w19037 & w31943) | (w19239 & w31943);
assign w19243 = ~w18537 & ~w18540;
assign w19244 = ~w18384 & ~w18541;
assign w19245 = ~w15044 & w36250;
assign w19246 = ~w15044 & w36251;
assign w19247 = w8295 & w12646;
assign w19248 = w8298 & w12651;
assign w19249 = (~w19247 & w12830) | (~w19247 & w36252) | (w12830 & w36252);
assign w19250 = (~a_8 & ~w19249) | (~a_8 & w36253) | (~w19249 & w36253);
assign w19251 = w19249 & w36254;
assign w19252 = ~w19250 & ~w19251;
assign w19253 = ~w19246 & w19252;
assign w19254 = ~w19245 & ~w19253;
assign w19255 = w19244 & ~w19254;
assign w19256 = ~w19244 & w19254;
assign w19257 = ~w19255 & ~w19256;
assign w19258 = w19243 & w19257;
assign w19259 = ~w19243 & ~w19257;
assign w19260 = ~w19258 & ~w19259;
assign w19261 = w19242 & w19260;
assign w19262 = w19254 & ~w19260;
assign w19263 = ~w18544 & ~w18561;
assign w19264 = ~w18562 & ~w19263;
assign w19265 = w9456 & ~w15027;
assign w19266 = w8295 & ~w12637;
assign w19267 = w8277 & w12651;
assign w19268 = w8298 & w12646;
assign w19269 = ~w19266 & w36255;
assign w19270 = a_8 & w19269;
assign w19271 = ~a_8 & ~w19269;
assign w19272 = ~w19270 & ~w19271;
assign w19273 = (w19272 & w15027) | (w19272 & w36256) | (w15027 & w36256);
assign w19274 = ~w19265 & ~w19273;
assign w19275 = w19264 & w19274;
assign w19276 = ~w19262 & ~w19275;
assign w19277 = ~w19261 & w19276;
assign w19278 = ~w19264 & ~w19274;
assign w19279 = (~w18559 & ~w18544) | (~w18559 & w31944) | (~w18544 & w31944);
assign w19280 = ~w18371 & ~w18563;
assign w19281 = w8295 & ~w12661;
assign w19282 = w8298 & ~w12637;
assign w19283 = w8277 & w12646;
assign w19284 = ~w19282 & ~w19283;
assign w19285 = ~w19281 & w19284;
assign w19286 = (w19285 & w14641) | (w19285 & w36257) | (w14641 & w36257);
assign w19287 = a_8 & ~w19286;
assign w19288 = (w14641 & w36258) | (w14641 & w36259) | (w36258 & w36259);
assign w19289 = ~w19287 & ~w19288;
assign w19290 = ~w19280 & ~w19289;
assign w19291 = w19279 & w19290;
assign w19292 = w19280 & ~w19289;
assign w19293 = ~w19279 & w19292;
assign w19294 = ~w19291 & ~w19293;
assign w19295 = ~w19278 & w19294;
assign w19296 = ~w19277 & w19295;
assign w19297 = w19280 & w19289;
assign w19298 = w19279 & w19297;
assign w19299 = ~w19280 & w19289;
assign w19300 = ~w19279 & w19299;
assign w19301 = ~w19298 & ~w19300;
assign w19302 = w19018 & w19301;
assign w19303 = ~w19296 & w19302;
assign w19304 = ~w19024 & ~w19303;
assign w19305 = ~w18584 & ~w18585;
assign w19306 = ~w18598 & ~w18601;
assign w19307 = w9456 & ~w14535;
assign w19308 = w8298 & ~w12668;
assign w19309 = w8277 & ~w12661;
assign w19310 = w8295 & ~w12630;
assign w19311 = ~w19308 & ~w19309;
assign w19312 = (~a_8 & ~w19311) | (~a_8 & w36260) | (~w19311 & w36260);
assign w19313 = w19311 & w36261;
assign w19314 = ~w19312 & ~w19313;
assign w19315 = (w19314 & w14535) | (w19314 & w36262) | (w14535 & w36262);
assign w19316 = ~w19307 & ~w19315;
assign w19317 = ~w19306 & w19316;
assign w19318 = w19306 & ~w19316;
assign w19319 = ~w19317 & ~w19318;
assign w19320 = w19305 & ~w19319;
assign w19321 = ~w19305 & w19319;
assign w19322 = ~w19320 & ~w19321;
assign w19323 = w19304 & ~w19322;
assign w19324 = w18988 & w36263;
assign w19325 = w18989 & w19002;
assign w19326 = ~w18988 & w19325;
assign w19327 = (w19316 & w18587) | (w19316 & w36264) | (w18587 & w36264);
assign w19328 = w18599 & w36265;
assign w19329 = ~w19305 & w19317;
assign w19330 = ~w19328 & ~w19329;
assign w19331 = ~w19326 & w19330;
assign w19332 = ~w19324 & w19331;
assign w19333 = (~w19003 & w19323) | (~w19003 & w36266) | (w19323 & w36266);
assign w19334 = w18968 & w18970;
assign w19335 = ~w18968 & ~w18970;
assign w19336 = ~w19334 & ~w19335;
assign w19337 = w18969 & w19336;
assign w19338 = ~w18969 & ~w19336;
assign w19339 = ~w19337 & ~w19338;
assign w19340 = w18986 & ~w19339;
assign w19341 = w19333 & w19340;
assign w19342 = ~w18987 & ~w19341;
assign w19343 = (~w18668 & ~w18647) | (~w18668 & w36267) | (~w18647 & w36267);
assign w19344 = w9456 & w13979;
assign w19345 = w8295 & w12869;
assign w19346 = w8277 & w12856;
assign w19347 = w8298 & ~w12860;
assign w19348 = ~w19345 & ~w19346;
assign w19349 = ~w19347 & w19348;
assign w19350 = a_8 & ~w19349;
assign w19351 = ~a_8 & w19349;
assign w19352 = (w19351 & ~w13979) | (w19351 & w36268) | (~w13979 & w36268);
assign w19353 = ~w19344 & ~w19350;
assign w19354 = ~w19352 & w19353;
assign w19355 = (w18680 & ~w19353) | (w18680 & w36269) | (~w19353 & w36269);
assign w19356 = w19353 & w36270;
assign w19357 = ~w19355 & ~w19356;
assign w19358 = w18690 & ~w19357;
assign w19359 = ~w18690 & w19357;
assign w19360 = ~w19358 & ~w19359;
assign w19361 = w19343 & w19360;
assign w19362 = ~w19343 & ~w19360;
assign w19363 = ~w19361 & ~w19362;
assign w19364 = ~w19342 & w19363;
assign w19365 = w19354 & ~w19363;
assign w19366 = w18711 & w18933;
assign w19367 = w18935 & w19366;
assign w19368 = ~w18711 & w18933;
assign w19369 = ~w18935 & w19368;
assign w19370 = ~w19367 & ~w19369;
assign w19371 = ~w19365 & w19370;
assign w19372 = ~w19364 & w19371;
assign w19373 = (w18938 & w19364) | (w18938 & w37577) | (w19364 & w37577);
assign w19374 = w18888 & ~w18901;
assign w19375 = ~w18902 & ~w19374;
assign w19376 = w18924 & ~w19375;
assign w19377 = w19373 & w19376;
assign w19378 = ~w18925 & ~w19377;
assign w19379 = w18240 & ~w18246;
assign w19380 = w18242 & ~w18246;
assign w19381 = (~w18765 & w18754) | (~w18765 & w31945) | (w18754 & w31945);
assign w19382 = ~w19380 & w19381;
assign w19383 = (~w18776 & ~w18753) | (~w18776 & w37578) | (~w18753 & w37578);
assign w19384 = w18792 & w18802;
assign w19385 = ~w12905 & w36271;
assign w19386 = ~w12892 & w36272;
assign w19387 = w8277 & ~w12878;
assign w19388 = ~w13598 & w36273;
assign w19389 = ~w19386 & ~w19387;
assign w19390 = ~w19385 & w19389;
assign w19391 = (a_8 & w19388) | (a_8 & w36274) | (w19388 & w36274);
assign w19392 = ~w19388 & w36275;
assign w19393 = ~w19391 & ~w19392;
assign w19394 = ~w19384 & ~w19393;
assign w19395 = w19383 & w19394;
assign w19396 = w19384 & ~w19393;
assign w19397 = ~w19383 & w19396;
assign w19398 = ~w19395 & ~w19397;
assign w19399 = ~w19378 & w19398;
assign w19400 = w18875 & w31946;
assign w19401 = ~w18357 & w18886;
assign w19402 = ~w18875 & w19401;
assign w19403 = w19384 & w19393;
assign w19404 = w19383 & w19403;
assign w19405 = ~w19384 & w19393;
assign w19406 = ~w19383 & w19405;
assign w19407 = ~w19404 & ~w19406;
assign w19408 = ~w19402 & w19407;
assign w19409 = ~w19400 & w19408;
assign w19410 = ~w19399 & w19409;
assign w19411 = ~w18887 & ~w19410;
assign w19412 = w18874 & w19411;
assign w19413 = ~w18874 & ~w19411;
assign w19414 = ~w19412 & ~w19413;
assign w19415 = (w9788 & w12616) | (w9788 & w36276) | (w12616 & w36276);
assign w19416 = (w9780 & w12612) | (w9780 & w36277) | (w12612 & w36277);
assign w19417 = ~w12930 & w36278;
assign w19418 = ~w19416 & ~w19417;
assign w19419 = ~w19415 & w19418;
assign w19420 = (w19419 & ~w13389) | (w19419 & w36279) | (~w13389 & w36279);
assign w19421 = a_5 & ~w19420;
assign w19422 = (~w13389 & w36280) | (~w13389 & w36281) | (w36280 & w36281);
assign w19423 = ~w19421 & ~w19422;
assign w19424 = w19414 & w19423;
assign w19425 = (w9788 & w12612) | (w9788 & w36282) | (w12612 & w36282);
assign w19426 = ~w12914 & w36283;
assign w19427 = ~w12930 & w36284;
assign w19428 = ~w19426 & ~w19427;
assign w19429 = ~w19425 & w19428;
assign w19430 = (w19429 & ~w13375) | (w19429 & w36285) | (~w13375 & w36285);
assign w19431 = a_5 & w19430;
assign w19432 = (w13375 & w36286) | (w13375 & w36287) | (w36286 & w36287);
assign w19433 = ~w19431 & ~w19432;
assign w19434 = (w19407 & w19378) | (w19407 & w31947) | (w19378 & w31947);
assign w19435 = ~w18886 & w19433;
assign w19436 = w18886 & ~w19433;
assign w19437 = ~w19435 & ~w19436;
assign w19438 = w18878 & w19437;
assign w19439 = ~w18878 & ~w19437;
assign w19440 = ~w19438 & ~w19439;
assign w19441 = w19434 & w19440;
assign w19442 = ~w19434 & ~w19440;
assign w19443 = ~w19441 & ~w19442;
assign w19444 = ~w19433 & ~w19443;
assign w19445 = ~w12892 & w36288;
assign w19446 = w9786 & w12874;
assign w19447 = w9780 & ~w12878;
assign w19448 = ~w19446 & ~w19447;
assign w19449 = ~w19445 & w19448;
assign w19450 = (w19449 & ~w13787) | (w19449 & w36289) | (~w13787 & w36289);
assign w19451 = a_5 & ~w19450;
assign w19452 = (~w13787 & w36290) | (~w13787 & w36291) | (w36290 & w36291);
assign w19453 = ~w19451 & ~w19452;
assign w19454 = w19363 & w19453;
assign w19455 = w19342 & w19454;
assign w19456 = ~w19363 & w19453;
assign w19457 = ~w19342 & w19456;
assign w19458 = ~w19455 & ~w19457;
assign w19459 = w19333 & ~w19339;
assign w19460 = (~w18974 & ~w19333) | (~w18974 & w31948) | (~w19333 & w31948);
assign w19461 = w18959 & w18986;
assign w19462 = w9788 & ~w12878;
assign w19463 = w9786 & w12869;
assign w19464 = w9780 & w12874;
assign w19465 = ~w19463 & ~w19464;
assign w19466 = ~w19462 & w19465;
assign w19467 = (w19466 & ~w13771) | (w19466 & w36292) | (~w13771 & w36292);
assign w19468 = a_5 & w19467;
assign w19469 = (w13771 & w36293) | (w13771 & w36294) | (w36293 & w36294);
assign w19470 = ~w19468 & ~w19469;
assign w19471 = ~w19461 & ~w19470;
assign w19472 = ~w19460 & w19471;
assign w19473 = w19461 & ~w19470;
assign w19474 = w19460 & w19473;
assign w19475 = ~w19472 & ~w19474;
assign w19476 = w19458 & w19475;
assign w19477 = ~w19363 & ~w19453;
assign w19478 = w19342 & w19477;
assign w19479 = w19363 & ~w19453;
assign w19480 = ~w19342 & w19479;
assign w19481 = ~w19478 & ~w19480;
assign w19482 = ~w19476 & w19481;
assign w19483 = ~w19333 & w19339;
assign w19484 = ~w19459 & ~w19483;
assign w19485 = w9788 & w12874;
assign w19486 = w9786 & ~w12860;
assign w19487 = w9780 & w12869;
assign w19488 = w9790 & w13965;
assign w19489 = ~w19486 & w36295;
assign w19490 = ~w19488 & w36296;
assign w19491 = (a_5 & w19488) | (a_5 & w36297) | (w19488 & w36297);
assign w19492 = ~w19490 & ~w19491;
assign w19493 = ~w19484 & ~w19492;
assign w19494 = w9788 & w12856;
assign w19495 = w9786 & ~w12630;
assign w19496 = w9780 & w12622;
assign w19497 = ~w19495 & ~w19496;
assign w19498 = ~w19494 & w19497;
assign w19499 = (w19498 & ~w14091) | (w19498 & w36298) | (~w14091 & w36298);
assign w19500 = a_5 & ~w19499;
assign w19501 = (~w14091 & w36299) | (~w14091 & w36300) | (w36299 & w36300);
assign w19502 = ~w19500 & ~w19501;
assign w19503 = (w19301 & w19277) | (w19301 & w36301) | (w19277 & w36301);
assign w19504 = w19023 & ~w19503;
assign w19505 = ~w19023 & w19503;
assign w19506 = ~w19504 & ~w19505;
assign w19507 = w19502 & ~w19506;
assign w19508 = ~w19502 & w19506;
assign w19509 = ~w19507 & ~w19508;
assign w19510 = ~w19221 & ~w19238;
assign w19511 = ~w19239 & ~w19510;
assign w19512 = w10033 & ~w15027;
assign w19513 = w9788 & ~w12637;
assign w19514 = w9786 & w12651;
assign w19515 = w9780 & w12646;
assign w19516 = ~w19513 & w36302;
assign w19517 = a_5 & w19516;
assign w19518 = ~a_5 & ~w19516;
assign w19519 = ~w19517 & ~w19518;
assign w19520 = (w19519 & w15027) | (w19519 & w36303) | (w15027 & w36303);
assign w19521 = ~w19512 & ~w19520;
assign w19522 = ~w19511 & ~w19521;
assign w19523 = ~w19198 & ~w19216;
assign w19524 = ~w19217 & ~w19523;
assign w19525 = w10033 & w14614;
assign w19526 = w9788 & w12651;
assign w19527 = w9786 & w12793;
assign w19528 = w9780 & ~w12830;
assign w19529 = ~w19526 & ~w19527;
assign w19530 = ~w19528 & w36304;
assign w19531 = (~a_5 & w19528) | (~a_5 & w36305) | (w19528 & w36305);
assign w19532 = ~w19530 & ~w19531;
assign w19533 = (w19532 & ~w14614) | (w19532 & w36306) | (~w14614 & w36306);
assign w19534 = ~w19525 & ~w19533;
assign w19535 = ~w19524 & ~w19534;
assign w19536 = w19173 & ~w19190;
assign w19537 = ~w19191 & ~w19536;
assign w19538 = w10033 & ~w15101;
assign w19539 = ~w12770 & w36307;
assign w19540 = w9780 & w12789;
assign w19541 = w9788 & w12793;
assign w19542 = ~w19539 & ~w19540;
assign w19543 = (~a_5 & ~w19542) | (~a_5 & w36308) | (~w19542 & w36308);
assign w19544 = w19542 & w36309;
assign w19545 = ~w19543 & ~w19544;
assign w19546 = (w19545 & w15101) | (w19545 & w36310) | (w15101 & w36310);
assign w19547 = ~w19538 & ~w19546;
assign w19548 = ~w19537 & ~w19547;
assign w19549 = w19157 & w19163;
assign w19550 = w19136 & ~w19549;
assign w19551 = ~w19136 & w19549;
assign w19552 = ~w19550 & ~w19551;
assign w19553 = w9780 & ~w12774;
assign w19554 = w9786 & w12732;
assign w19555 = ~w12770 & w36311;
assign w19556 = ~w19553 & ~w19554;
assign w19557 = (~a_5 & ~w19556) | (~a_5 & w36312) | (~w19556 & w36312);
assign w19558 = w19556 & w36313;
assign w19559 = ~w19557 & ~w19558;
assign w19560 = ~w15435 & w19559;
assign w19561 = (~a_5 & ~w9776) | (~a_5 & w36314) | (~w9776 & w36314);
assign w19562 = ~w10033 & ~w19561;
assign w19563 = w19556 & w36315;
assign w19564 = ~w19557 & ~w19563;
assign w19565 = w15435 & w19564;
assign w19566 = ~w19560 & ~w19565;
assign w19567 = ~w19552 & ~w19566;
assign w19568 = w9786 & w12701;
assign w19569 = w9788 & w12732;
assign w19570 = (~w19568 & ~w12739) | (~w19568 & w36316) | (~w12739 & w36316);
assign w19571 = ~w19569 & w19570;
assign w19572 = (~w15977 & w19583) | (~w15977 & w36317) | (w19583 & w36317);
assign w19573 = ~a_5 & w19571;
assign w19574 = a_8 & ~w19109;
assign w19575 = ~w19102 & w19574;
assign w19576 = w19102 & ~w19574;
assign w19577 = ~w19575 & ~w19576;
assign w19578 = (~w15977 & w36318) | (~w15977 & w36319) | (w36318 & w36319);
assign w19579 = ~w19572 & w19578;
assign w19580 = w19573 & ~w19577;
assign w19581 = (w19580 & w15977) | (w19580 & w36320) | (w15977 & w36320);
assign w19582 = w10033 & ~w19577;
assign w19583 = a_5 & ~w19571;
assign w19584 = ~w19577 & w19583;
assign w19585 = (~w19584 & w15977) | (~w19584 & w36321) | (w15977 & w36321);
assign w19586 = ~w19581 & w19585;
assign w19587 = (w19106 & ~w19104) | (w19106 & w36322) | (~w19104 & w36322);
assign w19588 = ~w19109 & ~w19587;
assign w19589 = w12689 & ~w15282;
assign w19590 = ~w15283 & ~w19589;
assign w19591 = w12684 & w36323;
assign w19592 = w9788 & w12701;
assign w19593 = (~w19591 & ~w12702) | (~w19591 & w36324) | (~w12702 & w36324);
assign w19594 = ~w19592 & w19593;
assign w19595 = (w19594 & w19590) | (w19594 & w36325) | (w19590 & w36325);
assign w19596 = w8270 & w12679;
assign w19597 = w9788 & w12702;
assign w19598 = w9780 & ~w11501;
assign w19599 = w12684 & w19598;
assign w19600 = w9786 & w12679;
assign w19601 = ~w19599 & ~w19600;
assign w19602 = w9776 & w12679;
assign w19603 = w9780 & w12679;
assign w19604 = w12684 & w36326;
assign w19605 = (~w19603 & w15324) | (~w19603 & w31951) | (w15324 & w31951);
assign w19606 = ~w19604 & w19605;
assign w19607 = (a_5 & ~w12679) | (a_5 & w36327) | (~w12679 & w36327);
assign w19608 = ~w19599 & w36328;
assign w19609 = ~w19597 & w19608;
assign w19610 = w19606 & w19609;
assign w19611 = ~w12702 & w15385;
assign w19612 = ~w15386 & ~w19611;
assign w19613 = w9790 & ~w19612;
assign w19614 = w19610 & ~w19613;
assign w19615 = ~w19596 & ~w19614;
assign w19616 = w19595 & ~w19615;
assign w19617 = w8271 & w12679;
assign w19618 = w19609 & w31952;
assign w19619 = ~w19617 & ~w19618;
assign w19620 = ~w19595 & ~w19619;
assign w19621 = ~w19616 & w36329;
assign w19622 = (w19588 & w19616) | (w19588 & w36330) | (w19616 & w36330);
assign w19623 = w9790 & w12715;
assign w19624 = w9788 & w12739;
assign w19625 = w9780 & w12701;
assign w19626 = w9786 & w12702;
assign w19627 = w9790 & ~w12700;
assign w19628 = w12711 & ~w19627;
assign w19629 = w9790 & w12700;
assign w19630 = ~w12711 & ~w19629;
assign w19631 = ~w19628 & ~w19630;
assign w19632 = ~w12704 & w19631;
assign w19633 = ~w19625 & ~w19626;
assign w19634 = ~w19624 & w19633;
assign w19635 = ~w19632 & w19634;
assign w19636 = ~w19623 & w19635;
assign w19637 = a_5 & ~w19636;
assign w19638 = ~a_5 & w19636;
assign w19639 = ~w19637 & ~w19638;
assign w19640 = (~w19621 & w19639) | (~w19621 & w36331) | (w19639 & w36331);
assign w19641 = w19586 & w19640;
assign w19642 = ~w19579 & ~w19641;
assign w19643 = w9780 & w12732;
assign w19644 = w9786 & w12739;
assign w19645 = w9788 & ~w12774;
assign w19646 = ~w19643 & ~w19644;
assign w19647 = ~w19645 & w19646;
assign w19648 = (w19647 & w15157) | (w19647 & w36332) | (w15157 & w36332);
assign w19649 = ~w19113 & ~w19134;
assign w19650 = ~w19135 & ~w19649;
assign w19651 = ~a_5 & w19650;
assign w19652 = a_5 & ~w19650;
assign w19653 = ~w19651 & ~w19652;
assign w19654 = w19648 & w19653;
assign w19655 = ~w19648 & ~w19653;
assign w19656 = ~w19654 & ~w19655;
assign w19657 = ~w19642 & w19656;
assign w19658 = w19552 & w19566;
assign w19659 = a_5 & w19650;
assign w19660 = w19648 & ~w19659;
assign w19661 = ~w19648 & ~w19651;
assign w19662 = ~w19660 & ~w19661;
assign w19663 = ~w19658 & ~w19662;
assign w19664 = ~w19657 & w19663;
assign w19665 = ~w19567 & ~w19664;
assign w19666 = w9786 & ~w12774;
assign w19667 = w9788 & w12789;
assign w19668 = ~w12770 & w36333;
assign w19669 = ~w19667 & w36334;
assign w19670 = ~w9790 & w19669;
assign w19671 = ~w15127 & w19669;
assign w19672 = (~w19670 & ~w19671) | (~w19670 & w31953) | (~w19671 & w31953);
assign w19673 = ~a_5 & w19672;
assign w19674 = a_5 & ~w19672;
assign w19675 = ~w19673 & ~w19674;
assign w19676 = w19087 & w19172;
assign w19677 = w19164 & ~w19676;
assign w19678 = ~w19164 & w19676;
assign w19679 = ~w19677 & ~w19678;
assign w19680 = ~w19675 & w19679;
assign w19681 = w19675 & ~w19679;
assign w19682 = ~w19680 & ~w19681;
assign w19683 = w19665 & w19682;
assign w19684 = w19537 & w19547;
assign w19685 = (~w19680 & ~w19537) | (~w19680 & w36335) | (~w19537 & w36335);
assign w19686 = (~w19548 & w19683) | (~w19548 & w36336) | (w19683 & w36336);
assign w19687 = w10033 & w15071;
assign w19688 = w9780 & w12793;
assign w19689 = w9786 & w12789;
assign w19690 = w9788 & ~w12830;
assign w19691 = ~w19688 & ~w19689;
assign w19692 = (~a_5 & w19690) | (~a_5 & w36337) | (w19690 & w36337);
assign w19693 = ~w19690 & w36338;
assign w19694 = ~w19692 & ~w19693;
assign w19695 = (w19694 & ~w15071) | (w19694 & w36339) | (~w15071 & w36339);
assign w19696 = ~w19687 & ~w19695;
assign w19697 = ~w19069 & ~w19192;
assign w19698 = (w19697 & w19191) | (w19697 & w31954) | (w19191 & w31954);
assign w19699 = ~w19191 & w31955;
assign w19700 = ~w19698 & ~w19699;
assign w19701 = w19696 & w19700;
assign w19702 = ~w19696 & ~w19700;
assign w19703 = ~w19701 & ~w19702;
assign w19704 = w19686 & w19703;
assign w19705 = w19524 & w19534;
assign w19706 = (~w19701 & ~w19524) | (~w19701 & w31956) | (~w19524 & w31956);
assign w19707 = (~w19535 & w19704) | (~w19535 & w31957) | (w19704 & w31957);
assign w19708 = ~w15044 & w36340;
assign w19709 = ~w15044 & w36341;
assign w19710 = w9788 & w12646;
assign w19711 = w9780 & w12651;
assign w19712 = (~w19710 & w12830) | (~w19710 & w36342) | (w12830 & w36342);
assign w19713 = w19712 & w36343;
assign w19714 = (~a_5 & ~w19712) | (~a_5 & w36344) | (~w19712 & w36344);
assign w19715 = ~w19713 & ~w19714;
assign w19716 = ~w19709 & w19715;
assign w19717 = ~w19708 & ~w19716;
assign w19718 = ~w19050 & ~w19218;
assign w19719 = (~w19214 & ~w19216) | (~w19214 & w31958) | (~w19216 & w31958);
assign w19720 = w19718 & w19719;
assign w19721 = ~w19718 & ~w19719;
assign w19722 = ~w19720 & ~w19721;
assign w19723 = w19717 & ~w19722;
assign w19724 = ~w19717 & w19722;
assign w19725 = ~w19723 & ~w19724;
assign w19726 = w19707 & w19725;
assign w19727 = w19511 & w19521;
assign w19728 = (~w19723 & ~w19511) | (~w19723 & w31959) | (~w19511 & w31959);
assign w19729 = ~w19726 & w19728;
assign w19730 = ~w19522 & ~w19729;
assign w19731 = w10033 & w14393;
assign w19732 = w9780 & ~w12661;
assign w19733 = w9786 & ~w12637;
assign w19734 = w9788 & ~w12668;
assign w19735 = ~w19732 & ~w19733;
assign w19736 = w19735 & w36345;
assign w19737 = (~a_5 & ~w19735) | (~a_5 & w36346) | (~w19735 & w36346);
assign w19738 = ~w19736 & ~w19737;
assign w19739 = (w19738 & ~w14393) | (w19738 & w36347) | (~w14393 & w36347);
assign w19740 = ~w19731 & ~w19739;
assign w19741 = w19260 & ~w19740;
assign w19742 = w19242 & w19741;
assign w19743 = ~w19260 & ~w19740;
assign w19744 = ~w19242 & w19743;
assign w19745 = ~w19742 & ~w19744;
assign w19746 = (~w19236 & ~w19221) | (~w19236 & w31960) | (~w19221 & w31960);
assign w19747 = ~w19037 & ~w19240;
assign w19748 = w9788 & ~w12661;
assign w19749 = w9780 & ~w12637;
assign w19750 = w9786 & w12646;
assign w19751 = ~w19749 & ~w19750;
assign w19752 = ~w19748 & w19751;
assign w19753 = (w19752 & w14641) | (w19752 & w36348) | (w14641 & w36348);
assign w19754 = a_5 & ~w19753;
assign w19755 = (w14641 & w36349) | (w14641 & w36350) | (w36349 & w36350);
assign w19756 = ~w19754 & ~w19755;
assign w19757 = w19747 & w19756;
assign w19758 = ~w19747 & ~w19756;
assign w19759 = ~w19757 & ~w19758;
assign w19760 = w19746 & w19759;
assign w19761 = ~w19746 & ~w19759;
assign w19762 = ~w19760 & ~w19761;
assign w19763 = w19745 & ~w19762;
assign w19764 = w19730 & w19763;
assign w19765 = ~w19260 & w19740;
assign w19766 = w19242 & w19765;
assign w19767 = w19260 & w19740;
assign w19768 = ~w19242 & w19767;
assign w19769 = ~w19766 & ~w19768;
assign w19770 = ~w19746 & ~w19747;
assign w19771 = w19746 & w19747;
assign w19772 = ~w19770 & ~w19771;
assign w19773 = w19756 & ~w19772;
assign w19774 = w19769 & ~w19773;
assign w19775 = w19745 & ~w19774;
assign w19776 = ~w19764 & ~w19775;
assign w19777 = ~w19261 & ~w19262;
assign w19778 = ~w19275 & ~w19278;
assign w19779 = w10033 & ~w14535;
assign w19780 = w9780 & ~w12668;
assign w19781 = w9786 & ~w12661;
assign w19782 = w9788 & ~w12630;
assign w19783 = ~w19780 & ~w19781;
assign w19784 = (~a_5 & ~w19783) | (~a_5 & w36351) | (~w19783 & w36351);
assign w19785 = w19783 & w36352;
assign w19786 = ~w19784 & ~w19785;
assign w19787 = (w19786 & w14535) | (w19786 & w36353) | (w14535 & w36353);
assign w19788 = ~w19779 & ~w19787;
assign w19789 = ~w19778 & w19788;
assign w19790 = w19778 & ~w19788;
assign w19791 = ~w19789 & ~w19790;
assign w19792 = w19777 & ~w19791;
assign w19793 = ~w19777 & w19791;
assign w19794 = ~w19792 & ~w19793;
assign w19795 = ~w19776 & ~w19794;
assign w19796 = (~w19278 & ~w19276) | (~w19278 & w31961) | (~w19276 & w31961);
assign w19797 = w19294 & w19301;
assign w19798 = w10033 & ~w14412;
assign w19799 = w9780 & ~w12630;
assign w19800 = w9786 & ~w12668;
assign w19801 = w9788 & w12622;
assign w19802 = ~w19799 & ~w19800;
assign w19803 = (~a_5 & ~w19802) | (~a_5 & w36354) | (~w19802 & w36354);
assign w19804 = w19802 & w36355;
assign w19805 = ~w19803 & ~w19804;
assign w19806 = (w19805 & w14412) | (w19805 & w36356) | (w14412 & w36356);
assign w19807 = ~w19798 & ~w19806;
assign w19808 = ~w19797 & w19807;
assign w19809 = w19796 & w19808;
assign w19810 = w19797 & w19807;
assign w19811 = ~w19796 & w19810;
assign w19812 = ~w19809 & ~w19811;
assign w19813 = ~w19777 & w19789;
assign w19814 = (w19788 & w19264) | (w19788 & w36357) | (w19264 & w36357);
assign w19815 = w19276 & w36358;
assign w19816 = ~w19813 & ~w19815;
assign w19817 = w19812 & w19816;
assign w19818 = ~w19796 & ~w19797;
assign w19819 = w19796 & w19797;
assign w19820 = ~w19818 & ~w19819;
assign w19821 = ~w19807 & ~w19820;
assign w19822 = (~w19821 & w19795) | (~w19821 & w36359) | (w19795 & w36359);
assign w19823 = w19509 & w19822;
assign w19824 = ~w19304 & w19322;
assign w19825 = ~w19323 & ~w19824;
assign w19826 = w10033 & w14442;
assign w19827 = w9780 & w12856;
assign w19828 = w9786 & w12622;
assign w19829 = w9788 & ~w12860;
assign w19830 = ~w19827 & ~w19828;
assign w19831 = ~w19829 & w36360;
assign w19832 = (~a_5 & w19829) | (~a_5 & w36361) | (w19829 & w36361);
assign w19833 = ~w19831 & ~w19832;
assign w19834 = (w19833 & ~w14442) | (w19833 & w36362) | (~w14442 & w36362);
assign w19835 = ~w19826 & ~w19834;
assign w19836 = w19825 & w19835;
assign w19837 = (~w19507 & ~w19825) | (~w19507 & w36363) | (~w19825 & w36363);
assign w19838 = ~w19823 & w19837;
assign w19839 = ~w19825 & ~w19835;
assign w19840 = (w19330 & ~w19304) | (w19330 & w36364) | (~w19304 & w36364);
assign w19841 = w10033 & w13979;
assign w19842 = w9788 & w12869;
assign w19843 = w9786 & w12856;
assign w19844 = w9780 & ~w12860;
assign w19845 = ~w19842 & ~w19843;
assign w19846 = ~w19844 & w19845;
assign w19847 = a_5 & ~w19846;
assign w19848 = ~a_5 & w19846;
assign w19849 = (w19848 & ~w13979) | (w19848 & w36365) | (~w13979 & w36365);
assign w19850 = ~w19841 & ~w19847;
assign w19851 = ~w19849 & w19850;
assign w19852 = (w19002 & ~w19850) | (w19002 & w36366) | (~w19850 & w36366);
assign w19853 = w19850 & w36367;
assign w19854 = ~w19852 & ~w19853;
assign w19855 = w18992 & ~w19854;
assign w19856 = ~w18992 & w19854;
assign w19857 = ~w19855 & ~w19856;
assign w19858 = w19840 & w19857;
assign w19859 = ~w19840 & ~w19857;
assign w19860 = ~w19858 & ~w19859;
assign w19861 = ~w19839 & w19860;
assign w19862 = ~w19838 & w19861;
assign w19863 = w19851 & ~w19860;
assign w19864 = w19339 & w19492;
assign w19865 = w19333 & w19864;
assign w19866 = ~w19339 & w19492;
assign w19867 = ~w19333 & w19866;
assign w19868 = ~w19865 & ~w19867;
assign w19869 = ~w19863 & w19868;
assign w19870 = (~w19493 & ~w19869) | (~w19493 & w36368) | (~w19869 & w36368);
assign w19871 = ~w19461 & w19470;
assign w19872 = ~w19473 & ~w19871;
assign w19873 = w19460 & w19872;
assign w19874 = ~w19460 & ~w19872;
assign w19875 = ~w19873 & ~w19874;
assign w19876 = w19481 & ~w19875;
assign w19877 = w19870 & w19876;
assign w19878 = ~w19482 & ~w19877;
assign w19879 = w18685 & ~w18691;
assign w19880 = ~w19343 & ~w19879;
assign w19881 = w18687 & ~w18691;
assign w19882 = ~w19354 & ~w19880;
assign w19883 = ~w19881 & w19882;
assign w19884 = (~w19883 & ~w19342) | (~w19883 & w36369) | (~w19342 & w36369);
assign w19885 = w18938 & w19370;
assign w19886 = ~w12905 & w36370;
assign w19887 = w9786 & ~w12878;
assign w19888 = ~w12892 & w36371;
assign w19889 = ~w13598 & w36372;
assign w19890 = ~w19887 & ~w19888;
assign w19891 = ~w19886 & w19890;
assign w19892 = ~w19889 & w36373;
assign w19893 = (~a_5 & w19889) | (~a_5 & w36374) | (w19889 & w36374);
assign w19894 = ~w19892 & ~w19893;
assign w19895 = w19885 & ~w19894;
assign w19896 = ~w19885 & w19894;
assign w19897 = ~w19895 & ~w19896;
assign w19898 = w19884 & w19897;
assign w19899 = ~w19884 & ~w19897;
assign w19900 = ~w19898 & ~w19899;
assign w19901 = ~w19878 & w19900;
assign w19902 = ~w12905 & w36375;
assign w19903 = ~w12892 & w36376;
assign w19904 = w9788 & ~w12910;
assign w19905 = w9790 & w13815;
assign w19906 = ~w19904 & w36377;
assign w19907 = ~w19905 & w36378;
assign w19908 = (a_5 & w19905) | (a_5 & w36379) | (w19905 & w36379);
assign w19909 = ~w19907 & ~w19908;
assign w19910 = w19375 & w19909;
assign w19911 = w19373 & w19910;
assign w19912 = ~w19375 & w19909;
assign w19913 = ~w19373 & w19912;
assign w19914 = ~w19911 & ~w19913;
assign w19915 = w19884 & w19885;
assign w19916 = (~w19894 & w19884) | (~w19894 & w19895) | (w19884 & w19895);
assign w19917 = ~w19915 & w19916;
assign w19918 = w19914 & ~w19917;
assign w19919 = ~w19901 & w19918;
assign w19920 = ~w19375 & ~w19909;
assign w19921 = w19373 & w19920;
assign w19922 = w19375 & ~w19909;
assign w19923 = ~w19373 & w19922;
assign w19924 = ~w19921 & ~w19923;
assign w19925 = ~w19919 & w19924;
assign w19926 = w18888 & w31962;
assign w19927 = ~w18888 & w18900;
assign w19928 = w18938 & ~w19927;
assign w19929 = ~w19926 & w19928;
assign w19930 = ~w19372 & w19929;
assign w19931 = ~w18904 & ~w19930;
assign w19932 = w18918 & w18924;
assign w19933 = ~w12914 & w36380;
assign w19934 = w9780 & ~w12910;
assign w19935 = ~w12905 & w36381;
assign w19936 = (w9790 & w13518) | (w9790 & w36382) | (w13518 & w36382);
assign w19937 = ~w19934 & ~w19935;
assign w19938 = ~w19933 & w19937;
assign w19939 = ~w19936 & w36383;
assign w19940 = (a_5 & w19936) | (a_5 & w36384) | (w19936 & w36384);
assign w19941 = ~w19939 & ~w19940;
assign w19942 = ~w19932 & ~w19941;
assign w19943 = w19932 & w19941;
assign w19944 = ~w19942 & ~w19943;
assign w19945 = w19931 & w19944;
assign w19946 = ~w19931 & ~w19944;
assign w19947 = ~w19945 & ~w19946;
assign w19948 = w19925 & ~w19947;
assign w19949 = w19941 & w19947;
assign w19950 = ~w12930 & w36385;
assign w19951 = w9786 & ~w12910;
assign w19952 = ~w12914 & w36386;
assign w19953 = ~w13501 & w36387;
assign w19954 = ~w19951 & ~w19952;
assign w19955 = ~w19950 & w19954;
assign w19956 = ~w19953 & w36388;
assign w19957 = (a_5 & w19953) | (a_5 & w36389) | (w19953 & w36389);
assign w19958 = ~w19956 & ~w19957;
assign w19959 = w19398 & w19407;
assign w19960 = w19378 & ~w19959;
assign w19961 = ~w19378 & w19959;
assign w19962 = ~w19960 & ~w19961;
assign w19963 = w19958 & w19962;
assign w19964 = ~w19949 & ~w19963;
assign w19965 = ~w19948 & w19964;
assign w19966 = w19440 & w31963;
assign w19967 = ~w19958 & ~w19962;
assign w19968 = w18886 & w19433;
assign w19969 = w18878 & w19968;
assign w19970 = ~w18878 & w19435;
assign w19971 = ~w19969 & ~w19970;
assign w19972 = ~w19434 & ~w19971;
assign w19973 = ~w19967 & ~w19972;
assign w19974 = ~w19966 & w19973;
assign w19975 = ~w19965 & w19974;
assign w19976 = ~w19444 & ~w19975;
assign w19977 = ~w19414 & ~w19423;
assign w19978 = ~w19976 & ~w19977;
assign w19979 = (~w19424 & w19976) | (~w19424 & w31964) | (w19976 & w31964);
assign w19980 = w18806 & ~w18866;
assign w19981 = (~w18867 & ~w18806) | (~w18867 & w31965) | (~w18806 & w31965);
assign w19982 = ~w18826 & ~w18839;
assign w19983 = w18826 & w18839;
assign w19984 = ~w19982 & ~w19983;
assign w19985 = ~w18847 & ~w19984;
assign w19986 = (~w19985 & w18811) | (~w19985 & w31966) | (w18811 & w31966);
assign w19987 = ~w18825 & ~w18839;
assign w19988 = (~w18824 & w18839) | (~w18824 & w31967) | (w18839 & w31967);
assign w19989 = w6996 & w12874;
assign w19990 = w6446 & ~w12860;
assign w19991 = w6998 & w12869;
assign w19992 = w6447 & w13965;
assign w19993 = ~w19990 & w36390;
assign w19994 = (a_14 & w19992) | (a_14 & w36391) | (w19992 & w36391);
assign w19995 = ~w19992 & w36392;
assign w19996 = ~w19994 & ~w19995;
assign w19997 = ~w16798 & w31968;
assign w19998 = w16798 & w17247;
assign w19999 = ~w17502 & ~w19998;
assign w20000 = ~w19997 & w19999;
assign w20001 = ~w17501 & w20000;
assign w20002 = ~w17252 & ~w20001;
assign w20003 = w17236 & w17257;
assign w20004 = w6304 & w12856;
assign w20005 = w6061 & w12622;
assign w20006 = w6059 & ~w12630;
assign w20007 = ~w20005 & ~w20006;
assign w20008 = ~w20004 & w20007;
assign w20009 = (w20008 & ~w14091) | (w20008 & w36393) | (~w14091 & w36393);
assign w20010 = a_17 & ~w20009;
assign w20011 = (~w14091 & w36394) | (~w14091 & w36395) | (w36394 & w36395);
assign w20012 = ~w20010 & ~w20011;
assign w20013 = w20003 & w20012;
assign w20014 = ~w20003 & ~w20012;
assign w20015 = ~w20013 & ~w20014;
assign w20016 = w20002 & w20015;
assign w20017 = ~w20002 & ~w20015;
assign w20018 = ~w20016 & ~w20017;
assign w20019 = w19996 & ~w20018;
assign w20020 = w19988 & w20019;
assign w20021 = w19996 & w20018;
assign w20022 = ~w19988 & w20021;
assign w20023 = ~w20020 & ~w20022;
assign w20024 = ~w19996 & w20018;
assign w20025 = w19988 & w20024;
assign w20026 = ~w19996 & ~w20018;
assign w20027 = ~w19988 & w20026;
assign w20028 = ~w20025 & ~w20027;
assign w20029 = w20023 & w20028;
assign w20030 = ~w12905 & w36396;
assign w20031 = ~w12892 & w36397;
assign w20032 = w7192 & ~w12878;
assign w20033 = ~w13598 & w36398;
assign w20034 = ~w20031 & ~w20032;
assign w20035 = ~w20030 & w20034;
assign w20036 = (a_11 & w20033) | (a_11 & w36399) | (w20033 & w36399);
assign w20037 = ~w20033 & w36400;
assign w20038 = ~w20036 & ~w20037;
assign w20039 = ~w20029 & ~w20038;
assign w20040 = w20029 & w20038;
assign w20041 = ~w20039 & ~w20040;
assign w20042 = w19986 & w20041;
assign w20043 = ~w19986 & ~w20041;
assign w20044 = ~w20042 & ~w20043;
assign w20045 = ~w12930 & w36401;
assign w20046 = w8277 & ~w12910;
assign w20047 = ~w12914 & w36402;
assign w20048 = ~w13501 & w36403;
assign w20049 = ~w20046 & ~w20047;
assign w20050 = ~w20045 & w20049;
assign w20051 = ~w20048 & w36404;
assign w20052 = (~a_8 & w20048) | (~a_8 & w36405) | (w20048 & w36405);
assign w20053 = ~w20051 & ~w20052;
assign w20054 = ~w20044 & w20053;
assign w20055 = w19981 & w20054;
assign w20056 = w20044 & w20053;
assign w20057 = ~w19981 & w20056;
assign w20058 = ~w20055 & ~w20057;
assign w20059 = w20044 & ~w20053;
assign w20060 = w19981 & w20059;
assign w20061 = ~w20044 & ~w20053;
assign w20062 = ~w19981 & w20061;
assign w20063 = ~w20060 & ~w20062;
assign w20064 = ~w18872 & w20063;
assign w20065 = ~w19412 & w20064;
assign w20066 = w20058 & ~w20065;
assign w20067 = ~w19986 & w20029;
assign w20068 = w20038 & ~w20067;
assign w20069 = ~w20042 & w20068;
assign w20070 = ~w20038 & w20067;
assign w20071 = w19986 & w20039;
assign w20072 = ~w18867 & ~w20071;
assign w20073 = ~w20070 & w20072;
assign w20074 = ~w19980 & w20073;
assign w20075 = ~w20069 & ~w20074;
assign w20076 = (w8295 & w12612) | (w8295 & w36406) | (w12612 & w36406);
assign w20077 = ~w12914 & w36407;
assign w20078 = ~w12930 & w36408;
assign w20079 = ~w20077 & ~w20078;
assign w20080 = ~w20076 & w20079;
assign w20081 = (w20080 & ~w13375) | (w20080 & w36409) | (~w13375 & w36409);
assign w20082 = a_8 & ~w20081;
assign w20083 = (~w13375 & w36410) | (~w13375 & w36411) | (w36410 & w36411);
assign w20084 = ~w20082 & ~w20083;
assign w20085 = ~w19985 & w20023;
assign w20086 = ~w18854 & w20085;
assign w20087 = w20028 & ~w20086;
assign w20088 = ~w12905 & w36412;
assign w20089 = w7511 & ~w12910;
assign w20090 = ~w12892 & w36413;
assign w20091 = w7193 & w13815;
assign w20092 = ~w20089 & w36414;
assign w20093 = (a_11 & w20091) | (a_11 & w36415) | (w20091 & w36415);
assign w20094 = ~w20091 & w36416;
assign w20095 = ~w20093 & ~w20094;
assign w20096 = ~w20003 & w20012;
assign w20097 = ~w20002 & w20096;
assign w20098 = w20002 & w20013;
assign w20099 = ~w20097 & ~w20098;
assign w20100 = w20018 & w20099;
assign w20101 = ~w18824 & w20099;
assign w20102 = ~w19987 & w20101;
assign w20103 = ~w20100 & ~w20102;
assign w20104 = w17508 & ~w17530;
assign w20105 = ~w17531 & ~w20104;
assign w20106 = w6998 & w12874;
assign w20107 = w6446 & w12869;
assign w20108 = w6996 & ~w12878;
assign w20109 = ~w20106 & ~w20107;
assign w20110 = w20109 & w36417;
assign w20111 = (w20110 & ~w13771) | (w20110 & w36418) | (~w13771 & w36418);
assign w20112 = w8564 & w13771;
assign w20113 = (a_14 & ~w20109) | (a_14 & w36419) | (~w20109 & w36419);
assign w20114 = ~w20112 & ~w20113;
assign w20115 = ~w20111 & w20114;
assign w20116 = w8391 & w14442;
assign w20117 = w6061 & w12856;
assign w20118 = w6059 & w12622;
assign w20119 = w6304 & ~w12860;
assign w20120 = ~w20117 & ~w20118;
assign w20121 = ~w20119 & w36420;
assign w20122 = (~a_17 & w20119) | (~a_17 & w36421) | (w20119 & w36421);
assign w20123 = ~w20121 & ~w20122;
assign w20124 = (w20123 & ~w14442) | (w20123 & w36422) | (~w14442 & w36422);
assign w20125 = ~w20116 & ~w20124;
assign w20126 = w20114 & w36423;
assign w20127 = (w20125 & ~w20114) | (w20125 & w36424) | (~w20114 & w36424);
assign w20128 = ~w20126 & ~w20127;
assign w20129 = w20105 & ~w20128;
assign w20130 = ~w20105 & w20128;
assign w20131 = ~w20129 & ~w20130;
assign w20132 = w20103 & w20131;
assign w20133 = ~w20103 & ~w20131;
assign w20134 = ~w20132 & ~w20133;
assign w20135 = w20095 & ~w20134;
assign w20136 = ~w20095 & w20134;
assign w20137 = ~w20135 & ~w20136;
assign w20138 = w20087 & w20137;
assign w20139 = ~w20087 & ~w20137;
assign w20140 = ~w20138 & ~w20139;
assign w20141 = w20084 & w20140;
assign w20142 = ~w20084 & ~w20140;
assign w20143 = ~w20141 & ~w20142;
assign w20144 = ~w20075 & w20143;
assign w20145 = w20075 & ~w20143;
assign w20146 = ~w20144 & ~w20145;
assign w20147 = w9788 & w12604;
assign w20148 = (w9786 & w12616) | (w9786 & w36425) | (w12616 & w36425);
assign w20149 = ~w12589 & w36426;
assign w20150 = ~w20148 & ~w20149;
assign w20151 = ~w20147 & w20150;
assign w20152 = (w20151 & w13288) | (w20151 & w36427) | (w13288 & w36427);
assign w20153 = a_5 & w20152;
assign w20154 = (~w13288 & w36428) | (~w13288 & w36429) | (w36428 & w36429);
assign w20155 = ~w20153 & ~w20154;
assign w20156 = w20146 & w20155;
assign w20157 = ~w20066 & w20156;
assign w20158 = ~w20146 & w20155;
assign w20159 = w20066 & w20158;
assign w20160 = ~w20157 & ~w20159;
assign w20161 = ~w18872 & ~w19412;
assign w20162 = w20058 & w20063;
assign w20163 = (w9780 & w12616) | (w9780 & w36430) | (w12616 & w36430);
assign w20164 = (w9786 & w12612) | (w9786 & w36431) | (w12612 & w36431);
assign w20165 = ~w12589 & w36432;
assign w20166 = ~w20163 & ~w20164;
assign w20167 = ~w20165 & w20166;
assign w20168 = (w20167 & ~w13123) | (w20167 & w36433) | (~w13123 & w36433);
assign w20169 = a_5 & w20168;
assign w20170 = (w13123 & w36434) | (w13123 & w36435) | (w36434 & w36435);
assign w20171 = ~w20169 & ~w20170;
assign w20172 = w20162 & ~w20171;
assign w20173 = ~w20162 & w20171;
assign w20174 = ~w20172 & ~w20173;
assign w20175 = ~w20161 & ~w20174;
assign w20176 = w20161 & w20174;
assign w20177 = ~w20175 & ~w20176;
assign w20178 = w20160 & ~w20177;
assign w20179 = ~w19979 & w20178;
assign w20180 = ~w20162 & ~w20171;
assign w20181 = ~w20161 & w20180;
assign w20182 = w20161 & w20172;
assign w20183 = ~w20181 & ~w20182;
assign w20184 = w20146 & ~w20155;
assign w20185 = ~w20158 & ~w20184;
assign w20186 = w20066 & w20185;
assign w20187 = ~w20066 & ~w20185;
assign w20188 = ~w20186 & ~w20187;
assign w20189 = w20183 & ~w20188;
assign w20190 = w20160 & ~w20189;
assign w20191 = ~w20179 & ~w20190;
assign w20192 = ~w20069 & ~w20140;
assign w20193 = ~w20074 & w20192;
assign w20194 = ~w20084 & ~w20193;
assign w20195 = ~w20144 & w20194;
assign w20196 = w20058 & ~w20195;
assign w20197 = ~w20065 & w20196;
assign w20198 = w20084 & w20146;
assign w20199 = ~w20095 & w20140;
assign w20200 = ~w20193 & ~w20199;
assign w20201 = (w8295 & w12616) | (w8295 & w36436) | (w12616 & w36436);
assign w20202 = (w8298 & w12612) | (w8298 & w36437) | (w12612 & w36437);
assign w20203 = ~w12930 & w36438;
assign w20204 = ~w20202 & ~w20203;
assign w20205 = ~w20201 & w20204;
assign w20206 = (w20205 & ~w13389) | (w20205 & w36439) | (~w13389 & w36439);
assign w20207 = a_8 & w20206;
assign w20208 = (w13389 & w36440) | (w13389 & w36441) | (w36440 & w36441);
assign w20209 = ~w20207 & ~w20208;
assign w20210 = w20115 & ~w20134;
assign w20211 = w20028 & w20134;
assign w20212 = ~w20086 & w20211;
assign w20213 = ~w20210 & ~w20212;
assign w20214 = ~w17530 & ~w20125;
assign w20215 = w17508 & w20214;
assign w20216 = w17530 & ~w20125;
assign w20217 = ~w17508 & w20216;
assign w20218 = ~w20215 & ~w20217;
assign w20219 = ~w20018 & w20218;
assign w20220 = ~w19988 & w20219;
assign w20221 = w20099 & ~w20125;
assign w20222 = ~w20099 & w20125;
assign w20223 = ~w20105 & ~w20222;
assign w20224 = ~w20221 & ~w20223;
assign w20225 = ~w20220 & ~w20224;
assign w20226 = (~w17532 & w17508) | (~w17532 & w31969) | (w17508 & w31969);
assign w20227 = w6059 & w12856;
assign w20228 = w6304 & w12869;
assign w20229 = (~w20227 & w12860) | (~w20227 & w36442) | (w12860 & w36442);
assign w20230 = ~w20228 & w20229;
assign w20231 = (w20230 & ~w13979) | (w20230 & w36443) | (~w13979 & w36443);
assign w20232 = a_17 & ~w20231;
assign w20233 = (~w13979 & w36444) | (~w13979 & w36445) | (w36444 & w36445);
assign w20234 = ~w20232 & ~w20233;
assign w20235 = w17218 & w31970;
assign w20236 = (w20234 & ~w17218) | (w20234 & w31971) | (~w17218 & w31971);
assign w20237 = ~w20235 & ~w20236;
assign w20238 = w20226 & ~w20237;
assign w20239 = ~w20226 & w20237;
assign w20240 = ~w20238 & ~w20239;
assign w20241 = ~w20225 & ~w20240;
assign w20242 = w20225 & w20240;
assign w20243 = ~w20241 & ~w20242;
assign w20244 = ~w12892 & w36446;
assign w20245 = w6998 & ~w12878;
assign w20246 = w6446 & w12874;
assign w20247 = ~w20245 & ~w20246;
assign w20248 = ~w20244 & w20247;
assign w20249 = (w20248 & ~w13787) | (w20248 & w36447) | (~w13787 & w36447);
assign w20250 = a_14 & ~w20249;
assign w20251 = (~w13787 & w36448) | (~w13787 & w36449) | (w36448 & w36449);
assign w20252 = ~w20250 & ~w20251;
assign w20253 = (w9061 & w13518) | (w9061 & w36450) | (w13518 & w36450);
assign w20254 = ~w12905 & w36451;
assign w20255 = w7489 & ~w12910;
assign w20256 = ~w12914 & w36452;
assign w20257 = ~w20254 & ~w20255;
assign w20258 = (a_11 & ~w20257) | (a_11 & w36453) | (~w20257 & w36453);
assign w20259 = (w7193 & w13518) | (w7193 & w36454) | (w13518 & w36454);
assign w20260 = w20257 & w36455;
assign w20261 = ~w20259 & w20260;
assign w20262 = ~w20253 & ~w20258;
assign w20263 = ~w20261 & w20262;
assign w20264 = w20252 & ~w20263;
assign w20265 = ~w20252 & w20263;
assign w20266 = ~w20264 & ~w20265;
assign w20267 = w20243 & ~w20266;
assign w20268 = ~w20243 & w20266;
assign w20269 = ~w20267 & ~w20268;
assign w20270 = w20213 & w20269;
assign w20271 = ~w20213 & ~w20269;
assign w20272 = ~w20270 & ~w20271;
assign w20273 = ~w20209 & ~w20272;
assign w20274 = w20209 & w20272;
assign w20275 = ~w20273 & ~w20274;
assign w20276 = ~w20200 & w20275;
assign w20277 = ~w20199 & ~w20272;
assign w20278 = ~w20193 & w20277;
assign w20279 = ~w20209 & ~w20278;
assign w20280 = ~w20276 & w20279;
assign w20281 = ~w20198 & ~w20280;
assign w20282 = ~w20197 & w20281;
assign w20283 = w20200 & ~w20275;
assign w20284 = ~w20276 & ~w20283;
assign w20285 = ~w20279 & w20284;
assign w20286 = w20263 & w20272;
assign w20287 = w20243 & w20252;
assign w20288 = w20213 & ~w20287;
assign w20289 = ~w20243 & ~w20252;
assign w20290 = (~w20289 & ~w20213) | (~w20289 & w31972) | (~w20213 & w31972);
assign w20291 = w17218 & w20234;
assign w20292 = ~w17531 & w36456;
assign w20293 = ~w20226 & w20236;
assign w20294 = ~w20292 & ~w20293;
assign w20295 = (w20294 & w20225) | (w20294 & w31973) | (w20225 & w31973);
assign w20296 = w6304 & w12874;
assign w20297 = w6059 & ~w12860;
assign w20298 = w6061 & w12869;
assign w20299 = w6063 & w13965;
assign w20300 = ~w20297 & w36457;
assign w20301 = ~w20299 & w36458;
assign w20302 = (a_17 & w20299) | (a_17 & w36459) | (w20299 & w36459);
assign w20303 = ~w20301 & ~w20302;
assign w20304 = ~w17541 & w20303;
assign w20305 = w17541 & ~w20303;
assign w20306 = ~w20304 & ~w20305;
assign w20307 = w17539 & w20306;
assign w20308 = ~w17539 & ~w20306;
assign w20309 = ~w20307 & ~w20308;
assign w20310 = ~w13598 & w36460;
assign w20311 = ~w12892 & w36461;
assign w20312 = w6446 & ~w12878;
assign w20313 = ~w12905 & w36462;
assign w20314 = ~w20311 & ~w20312;
assign w20315 = (a_14 & ~w20314) | (a_14 & w36463) | (~w20314 & w36463);
assign w20316 = ~w13598 & w36464;
assign w20317 = w20314 & w36465;
assign w20318 = ~w20316 & w20317;
assign w20319 = ~w20310 & ~w20315;
assign w20320 = ~w20318 & w20319;
assign w20321 = w20309 & ~w20320;
assign w20322 = ~w20309 & w20320;
assign w20323 = ~w20321 & ~w20322;
assign w20324 = w20295 & w20323;
assign w20325 = ~w20295 & ~w20323;
assign w20326 = ~w20324 & ~w20325;
assign w20327 = ~w12589 & w36466;
assign w20328 = (w8277 & w12612) | (w8277 & w36467) | (w12612 & w36467);
assign w20329 = (w8298 & w12616) | (w8298 & w36468) | (w12616 & w36468);
assign w20330 = ~w20327 & ~w20328;
assign w20331 = w20330 & w36469;
assign w20332 = (w20331 & ~w13123) | (w20331 & w36470) | (~w13123 & w36470);
assign w20333 = w9456 & w13123;
assign w20334 = (a_8 & ~w20330) | (a_8 & w36471) | (~w20330 & w36471);
assign w20335 = ~w20333 & ~w20334;
assign w20336 = ~w20332 & w20335;
assign w20337 = ~w12930 & w36472;
assign w20338 = w7192 & ~w12910;
assign w20339 = ~w12914 & w36473;
assign w20340 = ~w13501 & w36474;
assign w20341 = ~w20338 & ~w20339;
assign w20342 = ~w20337 & w20341;
assign w20343 = ~w20340 & w36475;
assign w20344 = (a_11 & w20340) | (a_11 & w36476) | (w20340 & w36476);
assign w20345 = ~w20343 & ~w20344;
assign w20346 = w20336 & ~w20345;
assign w20347 = ~w20336 & w20345;
assign w20348 = ~w20346 & ~w20347;
assign w20349 = w20326 & ~w20348;
assign w20350 = ~w20326 & w20348;
assign w20351 = ~w20349 & ~w20350;
assign w20352 = w20290 & ~w20351;
assign w20353 = ~w20290 & w20351;
assign w20354 = ~w20352 & ~w20353;
assign w20355 = ~w20278 & w36477;
assign w20356 = (~w20354 & w20278) | (~w20354 & w36478) | (w20278 & w36478);
assign w20357 = ~w20355 & ~w20356;
assign w20358 = ~w20285 & w20357;
assign w20359 = ~w20282 & w20358;
assign w20360 = w9788 & w12598;
assign w20361 = w9786 & w12604;
assign w20362 = w9780 & w12601;
assign w20363 = ~w20361 & ~w20362;
assign w20364 = ~w20360 & w20363;
assign w20365 = (w20364 & ~w12961) | (w20364 & w36479) | (~w12961 & w36479);
assign w20366 = ~a_5 & w20365;
assign w20367 = (w12961 & w36480) | (w12961 & w36481) | (w36480 & w36481);
assign w20368 = ~w20366 & ~w20367;
assign w20369 = w20359 & ~w20368;
assign w20370 = ~w20357 & ~w20368;
assign w20371 = (w20370 & w20282) | (w20370 & w36482) | (w20282 & w36482);
assign w20372 = ~w20369 & ~w20371;
assign w20373 = ~w20197 & ~w20198;
assign w20374 = w9788 & w12601;
assign w20375 = ~w12589 & w36483;
assign w20376 = w9780 & w12604;
assign w20377 = ~w20375 & ~w20376;
assign w20378 = ~w20374 & w20377;
assign w20379 = (w20378 & w13140) | (w20378 & w36484) | (w13140 & w36484);
assign w20380 = ~a_5 & w20379;
assign w20381 = (~w13140 & w36485) | (~w13140 & w36486) | (w36485 & w36486);
assign w20382 = ~w20380 & ~w20381;
assign w20383 = w20284 & w20382;
assign w20384 = ~w20284 & ~w20382;
assign w20385 = ~w20383 & ~w20384;
assign w20386 = w20373 & w20385;
assign w20387 = ~w20373 & ~w20385;
assign w20388 = ~w20386 & ~w20387;
assign w20389 = w20372 & w20388;
assign w20390 = ~w20191 & w20389;
assign w20391 = w20382 & ~w20388;
assign w20392 = ~w20357 & w20368;
assign w20393 = ~w20282 & w36487;
assign w20394 = w20357 & w20368;
assign w20395 = (w20394 & w20282) | (w20394 & w36488) | (w20282 & w36488);
assign w20396 = ~w20393 & ~w20395;
assign w20397 = ~w20391 & w20396;
assign w20398 = w20372 & ~w20397;
assign w20399 = ~w20390 & ~w20398;
assign w20400 = w20336 & ~w20357;
assign w20401 = ~w20359 & ~w20400;
assign w20402 = ~w20289 & w20326;
assign w20403 = ~w20288 & w20402;
assign w20404 = ~w20288 & w36489;
assign w20405 = ~w20326 & ~w20345;
assign w20406 = ~w20290 & w20405;
assign w20407 = ~w20404 & ~w20406;
assign w20408 = w20278 & w20407;
assign w20409 = (~w20345 & ~w20272) | (~w20345 & w36490) | (~w20272 & w36490);
assign w20410 = w20272 & w31974;
assign w20411 = ~w20290 & ~w20326;
assign w20412 = ~w20403 & ~w20411;
assign w20413 = ~w20410 & ~w20412;
assign w20414 = ~w20409 & ~w20413;
assign w20415 = ~w20408 & ~w20414;
assign w20416 = w20320 & ~w20326;
assign w20417 = (~w20416 & w20288) | (~w20416 & w36491) | (w20288 & w36491);
assign w20418 = ~w20303 & ~w20309;
assign w20419 = w20306 & w31975;
assign w20420 = ~w17539 & w20304;
assign w20421 = w20294 & ~w20420;
assign w20422 = ~w20419 & w20421;
assign w20423 = (~w20418 & w20241) | (~w20418 & w36492) | (w20241 & w36492);
assign w20424 = w6998 & w12906;
assign w20425 = w6996 & ~w12910;
assign w20426 = ~w12892 & w36493;
assign w20427 = ~w20425 & ~w20426;
assign w20428 = ~w20424 & w20427;
assign w20429 = (w20428 & ~w13815) | (w20428 & w36494) | (~w13815 & w36494);
assign w20430 = ~a_14 & w20429;
assign w20431 = (w13815 & w36495) | (w13815 & w36496) | (w36495 & w36496);
assign w20432 = ~w20430 & ~w20431;
assign w20433 = ~w17181 & w17199;
assign w20434 = ~w17200 & ~w20433;
assign w20435 = ~w17191 & ~w20434;
assign w20436 = (~w17202 & ~w17539) | (~w17202 & w36497) | (~w17539 & w36497);
assign w20437 = w17175 & w17180;
assign w20438 = w6304 & ~w12878;
assign w20439 = w6061 & w12874;
assign w20440 = w6059 & w12869;
assign w20441 = ~w20439 & ~w20440;
assign w20442 = ~w20438 & w20441;
assign w20443 = (w20442 & ~w13771) | (w20442 & w36498) | (~w13771 & w36498);
assign w20444 = a_17 & ~w20443;
assign w20445 = (~w13771 & w36499) | (~w13771 & w36500) | (w36499 & w36500);
assign w20446 = ~w20444 & ~w20445;
assign w20447 = w20437 & w20446;
assign w20448 = ~w20437 & ~w20446;
assign w20449 = ~w20447 & ~w20448;
assign w20450 = w20436 & w20449;
assign w20451 = ~w20436 & ~w20449;
assign w20452 = ~w20450 & ~w20451;
assign w20453 = ~w20432 & ~w20452;
assign w20454 = w20423 & w20453;
assign w20455 = ~w20432 & w20452;
assign w20456 = ~w20423 & w20455;
assign w20457 = ~w20454 & ~w20456;
assign w20458 = w20432 & w20452;
assign w20459 = w20423 & w20458;
assign w20460 = w20432 & ~w20452;
assign w20461 = ~w20423 & w20460;
assign w20462 = ~w20459 & ~w20461;
assign w20463 = w20457 & w20462;
assign w20464 = (w7511 & w12612) | (w7511 & w36501) | (w12612 & w36501);
assign w20465 = ~w12914 & w36502;
assign w20466 = ~w12930 & w36503;
assign w20467 = ~w20465 & ~w20466;
assign w20468 = ~w20464 & w20467;
assign w20469 = (w20468 & ~w13375) | (w20468 & w36504) | (~w13375 & w36504);
assign w20470 = ~a_11 & w20469;
assign w20471 = (w13375 & w36505) | (w13375 & w36506) | (w36505 & w36506);
assign w20472 = ~w20470 & ~w20471;
assign w20473 = w20463 & w20472;
assign w20474 = ~w20463 & ~w20472;
assign w20475 = ~w20473 & ~w20474;
assign w20476 = w20417 & w20475;
assign w20477 = ~w20417 & ~w20475;
assign w20478 = ~w20476 & ~w20477;
assign w20479 = w9780 & w12598;
assign w20480 = w9786 & w12601;
assign w20481 = ~w13011 & w36507;
assign w20482 = ~w20479 & ~w20480;
assign w20483 = ~w20481 & w20482;
assign w20484 = (w20483 & w13021) | (w20483 & w36508) | (w13021 & w36508);
assign w20485 = ~w12589 & w36509;
assign w20486 = (w8277 & w12616) | (w8277 & w36510) | (w12616 & w36510);
assign w20487 = w8295 & w12604;
assign w20488 = ~w20485 & ~w20486;
assign w20489 = ~w20487 & w20488;
assign w20490 = (w20489 & w13288) | (w20489 & w36511) | (w13288 & w36511);
assign w20491 = a_8 & ~w20490;
assign w20492 = (w13288 & w36512) | (w13288 & w36513) | (w36512 & w36513);
assign w20493 = ~w20491 & ~w20492;
assign w20494 = (a_5 & w20491) | (a_5 & w36514) | (w20491 & w36514);
assign w20495 = ~w20491 & w36515;
assign w20496 = ~w20494 & ~w20495;
assign w20497 = w20484 & ~w20496;
assign w20498 = ~w20484 & w20496;
assign w20499 = ~w20497 & ~w20498;
assign w20500 = w20478 & ~w20499;
assign w20501 = ~w20478 & w20499;
assign w20502 = ~w20500 & ~w20501;
assign w20503 = w20415 & ~w20502;
assign w20504 = ~w20415 & w20502;
assign w20505 = ~w20503 & ~w20504;
assign w20506 = w20401 & w20505;
assign w20507 = ~w20401 & ~w20505;
assign w20508 = ~w20506 & ~w20507;
assign w20509 = ~w20399 & w20508;
assign w20510 = (~w13021 & w36516) | (~w13021 & w36517) | (w36516 & w36517);
assign w20511 = (w13021 & w36518) | (w13021 & w36519) | (w36518 & w36519);
assign w20512 = ~w20510 & ~w20511;
assign w20513 = ~w20508 & w20512;
assign w20514 = (~w20513 & w20399) | (~w20513 & w31976) | (w20399 & w31976);
assign w20515 = w20415 & ~w20478;
assign w20516 = ~w20415 & w20478;
assign w20517 = ~w20515 & ~w20516;
assign w20518 = w20493 & ~w20517;
assign w20519 = w20401 & ~w20518;
assign w20520 = ~w20493 & w20517;
assign w20521 = (~w20520 & ~w20401) | (~w20520 & w31977) | (~w20401 & w31977);
assign w20522 = ~w13174 & w36520;
assign w20523 = w9786 & w12598;
assign w20524 = ~w13011 & w36521;
assign w20525 = ~w13205 & w36522;
assign w20526 = ~w20524 & w36523;
assign w20527 = ~w20525 & w36524;
assign w20528 = (~a_5 & w20525) | (~a_5 & w36525) | (w20525 & w36525);
assign w20529 = ~w20527 & ~w20528;
assign w20530 = ~w20463 & w20472;
assign w20531 = ~w20417 & w20530;
assign w20532 = w20417 & w20473;
assign w20533 = ~w20531 & ~w20532;
assign w20534 = w20478 & w20533;
assign w20535 = ~w20408 & w20533;
assign w20536 = ~w20414 & w20535;
assign w20537 = ~w20534 & ~w20536;
assign w20538 = ~w20416 & w20462;
assign w20539 = ~w20403 & w20538;
assign w20540 = (w20457 & w20403) | (w20457 & w36526) | (w20403 & w36526);
assign w20541 = ~w20437 & w20446;
assign w20542 = ~w20436 & w20541;
assign w20543 = w20436 & w20447;
assign w20544 = ~w20542 & ~w20543;
assign w20545 = (w20544 & ~w20423) | (w20544 & w31978) | (~w20423 & w31978);
assign w20546 = ~w12892 & w36527;
assign w20547 = w6061 & ~w12878;
assign w20548 = w6059 & w12874;
assign w20549 = ~w20547 & ~w20548;
assign w20550 = ~w20546 & w20549;
assign w20551 = (w20550 & ~w13787) | (w20550 & w36528) | (~w13787 & w36528);
assign w20552 = a_17 & w20551;
assign w20553 = (w13787 & w36529) | (w13787 & w36530) | (w36529 & w36530);
assign w20554 = ~w20552 & ~w20553;
assign w20555 = w17153 & w20554;
assign w20556 = ~w17153 & ~w20554;
assign w20557 = ~w20555 & ~w20556;
assign w20558 = ~w12914 & w36531;
assign w20559 = w6998 & ~w12910;
assign w20560 = ~w12905 & w36532;
assign w20561 = (w6447 & w13518) | (w6447 & w36533) | (w13518 & w36533);
assign w20562 = ~w20559 & ~w20560;
assign w20563 = ~w20558 & w20562;
assign w20564 = ~w20561 & w36534;
assign w20565 = (a_14 & w20561) | (a_14 & w36535) | (w20561 & w36535);
assign w20566 = ~w20564 & ~w20565;
assign w20567 = w17544 & ~w20566;
assign w20568 = ~w17544 & w20566;
assign w20569 = ~w20567 & ~w20568;
assign w20570 = w20557 & w20569;
assign w20571 = ~w20557 & ~w20569;
assign w20572 = ~w20570 & ~w20571;
assign w20573 = w20545 & w20572;
assign w20574 = ~w20545 & ~w20572;
assign w20575 = ~w20573 & ~w20574;
assign w20576 = ~w20539 & w31979;
assign w20577 = (~w20575 & w20539) | (~w20575 & w31980) | (w20539 & w31980);
assign w20578 = ~w20576 & ~w20577;
assign w20579 = w8295 & w12601;
assign w20580 = w8298 & w12604;
assign w20581 = ~w12589 & w36536;
assign w20582 = ~w20580 & ~w20581;
assign w20583 = ~w20579 & w20582;
assign w20584 = (w20583 & w13140) | (w20583 & w36537) | (w13140 & w36537);
assign w20585 = ~a_8 & w20584;
assign w20586 = (~w13140 & w36538) | (~w13140 & w36539) | (w36538 & w36539);
assign w20587 = ~w20585 & ~w20586;
assign w20588 = (w7511 & w12616) | (w7511 & w36540) | (w12616 & w36540);
assign w20589 = (w7489 & w12612) | (w7489 & w36541) | (w12612 & w36541);
assign w20590 = ~w12930 & w36542;
assign w20591 = ~w20589 & ~w20590;
assign w20592 = ~w20588 & w20591;
assign w20593 = (w20592 & ~w13389) | (w20592 & w36543) | (~w13389 & w36543);
assign w20594 = ~a_11 & w20593;
assign w20595 = (w13389 & w36544) | (w13389 & w36545) | (w36544 & w36545);
assign w20596 = ~w20594 & ~w20595;
assign w20597 = ~w20587 & w20596;
assign w20598 = w20587 & ~w20596;
assign w20599 = ~w20597 & ~w20598;
assign w20600 = w20578 & ~w20599;
assign w20601 = ~w20578 & w20599;
assign w20602 = ~w20600 & ~w20601;
assign w20603 = w20537 & w20602;
assign w20604 = ~w20537 & ~w20602;
assign w20605 = ~w20603 & ~w20604;
assign w20606 = w20529 & w20605;
assign w20607 = ~w20529 & ~w20605;
assign w20608 = ~w20606 & ~w20607;
assign w20609 = w20521 & w20608;
assign w20610 = ~w20521 & ~w20608;
assign w20611 = ~w20609 & ~w20610;
assign w20612 = (w13201 & w36548) | (w13201 & w36549) | (w36548 & w36549);
assign w20613 = (~w13173 & w36550) | (~w13173 & w36551) | (w36550 & w36551);
assign w20614 = ~w20612 & w20613;
assign w20615 = (a_2 & ~w13177) | (a_2 & w34211) | (~w13177 & w34211);
assign w20616 = w20614 & ~w20615;
assign w20617 = (a_2 & w20612) | (a_2 & w36552) | (w20612 & w36552);
assign w20618 = ~w20616 & ~w20617;
assign w20619 = w20611 & w20618;
assign w20620 = ~w20514 & w20619;
assign w20621 = (w20618 & w20508) | (w20618 & w31981) | (w20508 & w31981);
assign w20622 = ~w20611 & w20621;
assign w20623 = ~w20509 & w20622;
assign w20624 = (w13173 & w36553) | (w13173 & w36554) | (w36553 & w36554);
assign w20625 = w10837 & ~w13264;
assign w20626 = (~w20624 & ~w13177) | (~w20624 & w36555) | (~w13177 & w36555);
assign w20627 = ~w13174 & w36556;
assign w20628 = a_2 & ~w20627;
assign w20629 = ~w20625 & w36557;
assign w20630 = (a_2 & w20625) | (a_2 & w36558) | (w20625 & w36558);
assign w20631 = ~w20629 & ~w20630;
assign w20632 = w20508 & w20631;
assign w20633 = w20399 & w20632;
assign w20634 = ~w20508 & w20631;
assign w20635 = ~w20399 & w20634;
assign w20636 = ~w20633 & ~w20635;
assign w20637 = ~w20623 & w20636;
assign w20638 = ~w20620 & w20637;
assign w20639 = w20611 & ~w20618;
assign w20640 = w20514 & w20639;
assign w20641 = ~w20611 & ~w20618;
assign w20642 = ~w20514 & w20641;
assign w20643 = ~w20640 & ~w20642;
assign w20644 = ~w20638 & w20643;
assign w20645 = ~w19665 & ~w19682;
assign w20646 = ~w19683 & ~w20645;
assign w20647 = w3 & w12651;
assign w20648 = w10837 & w14614;
assign w20649 = (~w20647 & w12830) | (~w20647 & w36559) | (w12830 & w36559);
assign w20650 = ~w20648 & w20649;
assign w20651 = (a_2 & ~w12793) | (a_2 & w34211) | (~w12793 & w34211);
assign w20652 = w20650 & ~w20651;
assign w20653 = (a_2 & w20648) | (a_2 & w36560) | (w20648 & w36560);
assign w20654 = ~w20652 & ~w20653;
assign w20655 = ~w20646 & ~w20654;
assign w20656 = w10835 & w12651;
assign w20657 = w3 & w12646;
assign w20658 = ~w15044 & w36561;
assign w20659 = ~w20656 & ~w20657;
assign w20660 = ~w20658 & w20659;
assign w20661 = (a_2 & w12830) | (a_2 & w34211) | (w12830 & w34211);
assign w20662 = w20660 & ~w20661;
assign w20663 = (a_2 & w20658) | (a_2 & w36562) | (w20658 & w36562);
assign w20664 = ~w20662 & ~w20663;
assign w20665 = ~w19548 & ~w19684;
assign w20666 = (~w19680 & ~w19665) | (~w19680 & w36563) | (~w19665 & w36563);
assign w20667 = ~w20665 & w20666;
assign w20668 = w20665 & ~w20666;
assign w20669 = ~w20667 & ~w20668;
assign w20670 = ~w20664 & ~w20669;
assign w20671 = w10909 & w12789;
assign w20672 = w10835 & w12793;
assign w20673 = w10837 & w15071;
assign w20674 = (~w20672 & w12830) | (~w20672 & w36564) | (w12830 & w36564);
assign w20675 = (~a_2 & w20673) | (~a_2 & w36565) | (w20673 & w36565);
assign w20676 = ~w20673 & w36566;
assign w20677 = ~w20675 & ~w20676;
assign w20678 = ~w20671 & ~w20677;
assign w20679 = ~w19567 & ~w19658;
assign w20680 = (~w19662 & ~w19656) | (~w19662 & w36567) | (~w19656 & w36567);
assign w20681 = w20679 & w20680;
assign w20682 = ~w20679 & ~w20680;
assign w20683 = ~w20681 & ~w20682;
assign w20684 = w20678 & ~w20683;
assign w20685 = ~w20678 & w20683;
assign w20686 = w19642 & ~w19656;
assign w20687 = ~w19657 & ~w20686;
assign w20688 = ~w12770 & w36568;
assign w20689 = w3 & w12793;
assign w20690 = w10835 & w12789;
assign w20691 = ~w20689 & ~w20690;
assign w20692 = (w20691 & w15101) | (w20691 & w36569) | (w15101 & w36569);
assign w20693 = ~a_2 & ~w20692;
assign w20694 = (w15101 & w36570) | (w15101 & w36571) | (w36570 & w36571);
assign w20695 = (~w20688 & w20693) | (~w20688 & w36572) | (w20693 & w36572);
assign w20696 = ~w20687 & ~w20695;
assign w20697 = ~w12770 & w36573;
assign w20698 = w3 & w12789;
assign w20699 = ~w20697 & ~w20698;
assign w20700 = (w20699 & w15128) | (w20699 & w36574) | (w15128 & w36574);
assign w20701 = (a_2 & w12774) | (a_2 & w34211) | (w12774 & w34211);
assign w20702 = w20700 & ~w20701;
assign w20703 = (~w15128 & w36575) | (~w15128 & w36576) | (w36575 & w36576);
assign w20704 = ~w19579 & w19586;
assign w20705 = w19640 & ~w20704;
assign w20706 = ~w19640 & w20704;
assign w20707 = ~w20705 & ~w20706;
assign w20708 = w10909 & w12732;
assign w20709 = ~w12770 & w36577;
assign w20710 = w10835 & ~w12774;
assign w20711 = ~w20709 & ~w20710;
assign w20712 = (w20711 & ~w15435) | (w20711 & w36578) | (~w15435 & w36578);
assign w20713 = ~a_2 & ~w20712;
assign w20714 = (~w15435 & w36579) | (~w15435 & w36580) | (w36579 & w36580);
assign w20715 = (~w20708 & w20713) | (~w20708 & w36581) | (w20713 & w36581);
assign w20716 = ~w19621 & ~w19622;
assign w20717 = ~w19639 & w20716;
assign w20718 = w19639 & ~w20716;
assign w20719 = ~w20717 & ~w20718;
assign w20720 = ~w20715 & w20719;
assign w20721 = w20715 & ~w20719;
assign w20722 = ~w19614 & w36582;
assign w20723 = (w19595 & w20722) | (w19595 & w36583) | (w20722 & w36583);
assign w20724 = ~w20722 & w36584;
assign w20725 = ~w20723 & ~w20724;
assign w20726 = w10909 & w12739;
assign w20727 = w3 & ~w12774;
assign w20728 = w10835 & w12732;
assign w20729 = ~w20727 & ~w20728;
assign w20730 = (w20729 & w15157) | (w20729 & w36585) | (w15157 & w36585);
assign w20731 = ~a_2 & ~w20730;
assign w20732 = (w15157 & w36586) | (w15157 & w36587) | (w36586 & w36587);
assign w20733 = (~w20726 & w20731) | (~w20726 & w36588) | (w20731 & w36588);
assign w20734 = ~w20725 & w20733;
assign w20735 = w20725 & ~w20733;
assign w20736 = w12679 & w36589;
assign w20737 = w19605 & w36590;
assign w20738 = a_5 & ~w20737;
assign w20739 = ~w19597 & w19601;
assign w20740 = ~w19613 & w36591;
assign w20741 = (w20738 & w19613) | (w20738 & w36592) | (w19613 & w36592);
assign w20742 = ~w20740 & ~w20741;
assign w20743 = (a_2 & ~w12701) | (a_2 & w34211) | (~w12701 & w34211);
assign w20744 = w3 & w12732;
assign w20745 = w10835 & w12739;
assign w20746 = ~w20744 & ~w20745;
assign w20747 = (w20746 & w15977) | (w20746 & w36593) | (w15977 & w36593);
assign w20748 = ~w20743 & w20747;
assign w20749 = (~w15977 & w36594) | (~w15977 & w36595) | (w36594 & w36595);
assign w20750 = ~w20748 & w36596;
assign w20751 = (w20736 & ~w19605) | (w20736 & w36597) | (~w19605 & w36597);
assign w20752 = ~w20737 & ~w20751;
assign w20753 = w12684 & w36598;
assign w20754 = w10835 & w12702;
assign w20755 = w3 & w12701;
assign w20756 = ~w20754 & ~w20755;
assign w20757 = (w20756 & w19590) | (w20756 & w36599) | (w19590 & w36599);
assign w20758 = ~a_2 & w20757;
assign w20759 = w12679 & w36600;
assign w20760 = ~w20757 & ~w20759;
assign w20761 = ~a_1 & ~w15324;
assign w20762 = ~w12702 & ~w20761;
assign w20763 = w12684 & w36601;
assign w20764 = ~w12679 & ~w20763;
assign w20765 = (w20764 & w20762) | (w20764 & w36602) | (w20762 & w36602);
assign w20766 = (~w20753 & w20765) | (~w20753 & w36603) | (w20765 & w36603);
assign w20767 = ~w20758 & w20766;
assign w20768 = (~w20752 & ~w20767) | (~w20752 & w36604) | (~w20767 & w36604);
assign w20769 = w20767 & w36605;
assign w20770 = w10909 & w12702;
assign w20771 = w10835 & w12701;
assign w20772 = w10837 & ~w15278;
assign w20773 = (~w20771 & ~w12739) | (~w20771 & w36606) | (~w12739 & w36606);
assign w20774 = (a_2 & w20772) | (a_2 & w36607) | (w20772 & w36607);
assign w20775 = ~w20772 & w36608;
assign w20776 = ~w20770 & ~w20774;
assign w20777 = (~w20769 & ~w20776) | (~w20769 & w36609) | (~w20776 & w36609);
assign w20778 = ~w20768 & ~w20777;
assign w20779 = ~w20750 & ~w20778;
assign w20780 = (~w20742 & w20748) | (~w20742 & w36610) | (w20748 & w36610);
assign w20781 = ~w20779 & ~w20780;
assign w20782 = ~w20735 & w20781;
assign w20783 = ~w20721 & ~w20734;
assign w20784 = ~w20782 & w20783;
assign w20785 = ~w20702 & ~w20703;
assign w20786 = (~w20784 & w36612) | (~w20784 & w36613) | (w36612 & w36613);
assign w20787 = w20687 & w20695;
assign w20788 = ~w20784 & w36614;
assign w20789 = ~w20787 & ~w20788;
assign w20790 = ~w20786 & w20789;
assign w20791 = ~w20685 & ~w20696;
assign w20792 = ~w20790 & w20791;
assign w20793 = (~w20684 & ~w20646) | (~w20684 & w36615) | (~w20646 & w36615);
assign w20794 = ~w20792 & w20793;
assign w20795 = ~w20655 & ~w20670;
assign w20796 = ~w20794 & w20795;
assign w20797 = w20664 & w20669;
assign w20798 = ~w19686 & ~w19703;
assign w20799 = ~w19704 & ~w20798;
assign w20800 = w10909 & w12651;
assign w20801 = w3 & ~w12637;
assign w20802 = w10835 & w12646;
assign w20803 = ~w20801 & ~w20802;
assign w20804 = (w20803 & w15027) | (w20803 & w36616) | (w15027 & w36616);
assign w20805 = ~a_2 & ~w20804;
assign w20806 = (w15027 & w36617) | (w15027 & w36618) | (w36617 & w36618);
assign w20807 = (~w20800 & w20805) | (~w20800 & w36619) | (w20805 & w36619);
assign w20808 = w20799 & w20807;
assign w20809 = ~w20797 & ~w20808;
assign w20810 = ~w20796 & w20809;
assign w20811 = ~w20799 & ~w20807;
assign w20812 = ~w19535 & ~w19705;
assign w20813 = ~w19701 & ~w19704;
assign w20814 = ~w20812 & w20813;
assign w20815 = w20812 & ~w20813;
assign w20816 = ~w20814 & ~w20815;
assign w20817 = w3 & ~w12661;
assign w20818 = w10835 & ~w12637;
assign w20819 = ~w20817 & ~w20818;
assign w20820 = (w20819 & w14641) | (w20819 & w36620) | (w14641 & w36620);
assign w20821 = (a_2 & ~w12646) | (a_2 & w34211) | (~w12646 & w34211);
assign w20822 = w20820 & ~w20821;
assign w20823 = (~w14641 & w36621) | (~w14641 & w36622) | (w36621 & w36622);
assign w20824 = ~w20822 & ~w20823;
assign w20825 = (~w20811 & w20816) | (~w20811 & w36623) | (w20816 & w36623);
assign w20826 = ~w20810 & w20825;
assign w20827 = w20816 & w20824;
assign w20828 = ~w19707 & ~w19725;
assign w20829 = ~w19726 & ~w20828;
assign w20830 = w3 & ~w12668;
assign w20831 = w10835 & ~w12661;
assign w20832 = ~w20830 & ~w20831;
assign w20833 = (w20832 & ~w14393) | (w20832 & w36624) | (~w14393 & w36624);
assign w20834 = (a_2 & w12637) | (a_2 & w34211) | (w12637 & w34211);
assign w20835 = w20833 & ~w20834;
assign w20836 = (w14393 & w36625) | (w14393 & w36626) | (w36625 & w36626);
assign w20837 = ~w20835 & ~w20836;
assign w20838 = w20829 & w20837;
assign w20839 = ~w20827 & ~w20838;
assign w20840 = ~w20826 & w20839;
assign w20841 = ~w20829 & ~w20837;
assign w20842 = ~w19522 & ~w19727;
assign w20843 = ~w19723 & ~w19726;
assign w20844 = ~w20842 & w20843;
assign w20845 = w20842 & ~w20843;
assign w20846 = ~w20844 & ~w20845;
assign w20847 = w3 & ~w12630;
assign w20848 = w10835 & ~w12668;
assign w20849 = ~w20847 & ~w20848;
assign w20850 = (w20849 & w14535) | (w20849 & w36627) | (w14535 & w36627);
assign w20851 = (a_2 & w12661) | (a_2 & w34211) | (w12661 & w34211);
assign w20852 = w20850 & ~w20851;
assign w20853 = (~w14535 & w36628) | (~w14535 & w36629) | (w36628 & w36629);
assign w20854 = ~w20852 & ~w20853;
assign w20855 = (~w20841 & w20846) | (~w20841 & w36630) | (w20846 & w36630);
assign w20856 = ~w20840 & w20855;
assign w20857 = w20846 & w20854;
assign w20858 = w19730 & ~w19762;
assign w20859 = ~w19730 & w19762;
assign w20860 = ~w20858 & ~w20859;
assign w20861 = w10835 & ~w12630;
assign w20862 = w3 & w12622;
assign w20863 = ~w20861 & ~w20862;
assign w20864 = (w20863 & w14412) | (w20863 & w36631) | (w14412 & w36631);
assign w20865 = (a_2 & w12668) | (a_2 & w34211) | (w12668 & w34211);
assign w20866 = w20864 & ~w20865;
assign w20867 = (~w14412 & w36632) | (~w14412 & w36633) | (w36632 & w36633);
assign w20868 = ~w20866 & ~w20867;
assign w20869 = w20860 & w20868;
assign w20870 = ~w20857 & ~w20869;
assign w20871 = ~w20860 & ~w20868;
assign w20872 = w19745 & w19769;
assign w20873 = (~w19773 & ~w19730) | (~w19773 & w36634) | (~w19730 & w36634);
assign w20874 = ~w20872 & w20873;
assign w20875 = w20872 & ~w20873;
assign w20876 = ~w20874 & ~w20875;
assign w20877 = w3 & w12856;
assign w20878 = w10835 & w12622;
assign w20879 = ~w20877 & ~w20878;
assign w20880 = (w20879 & ~w14091) | (w20879 & w36635) | (~w14091 & w36635);
assign w20881 = (a_2 & w12630) | (a_2 & w34211) | (w12630 & w34211);
assign w20882 = w20880 & ~w20881;
assign w20883 = (w14091 & w36636) | (w14091 & w36637) | (w36636 & w36637);
assign w20884 = ~w20882 & ~w20883;
assign w20885 = ~w20876 & ~w20884;
assign w20886 = (~w20871 & ~w20870) | (~w20871 & w36638) | (~w20870 & w36638);
assign w20887 = ~w20885 & w20886;
assign w20888 = w20876 & w20884;
assign w20889 = w19776 & w19794;
assign w20890 = ~w19795 & ~w20889;
assign w20891 = w10835 & w12856;
assign w20892 = w10837 & w14442;
assign w20893 = (~w20891 & w12860) | (~w20891 & w36639) | (w12860 & w36639);
assign w20894 = ~w20892 & w20893;
assign w20895 = (a_2 & ~w12622) | (a_2 & w34211) | (~w12622 & w34211);
assign w20896 = w20894 & ~w20895;
assign w20897 = (a_2 & w20892) | (a_2 & w36640) | (w20892 & w36640);
assign w20898 = ~w20896 & ~w20897;
assign w20899 = (~w20888 & ~w20890) | (~w20888 & w36641) | (~w20890 & w36641);
assign w20900 = ~w20887 & w20899;
assign w20901 = ~w20890 & ~w20898;
assign w20902 = w19812 & ~w19821;
assign w20903 = (w19816 & w19776) | (w19816 & w36642) | (w19776 & w36642);
assign w20904 = ~w20902 & w20903;
assign w20905 = w20902 & ~w20903;
assign w20906 = ~w20904 & ~w20905;
assign w20907 = w10835 & ~w12860;
assign w20908 = w3 & w12869;
assign w20909 = ~w20907 & ~w20908;
assign w20910 = (w20909 & ~w13979) | (w20909 & w36643) | (~w13979 & w36643);
assign w20911 = (a_2 & ~w12856) | (a_2 & w34211) | (~w12856 & w34211);
assign w20912 = w20910 & ~w20911;
assign w20913 = (w13979 & w36644) | (w13979 & w36645) | (w36644 & w36645);
assign w20914 = ~w20912 & ~w20913;
assign w20915 = (~w20901 & w20906) | (~w20901 & w31982) | (w20906 & w31982);
assign w20916 = ~w20900 & w20915;
assign w20917 = w20906 & w20914;
assign w20918 = ~w19509 & ~w19822;
assign w20919 = ~w19823 & ~w20918;
assign w20920 = w3 & w12874;
assign w20921 = w10835 & w12869;
assign w20922 = ~w20920 & ~w20921;
assign w20923 = (w20922 & ~w13965) | (w20922 & w36646) | (~w13965 & w36646);
assign w20924 = (a_2 & w12860) | (a_2 & w34211) | (w12860 & w34211);
assign w20925 = w20923 & ~w20924;
assign w20926 = (w13965 & w36647) | (w13965 & w36648) | (w36647 & w36648);
assign w20927 = ~w20925 & ~w20926;
assign w20928 = w20919 & w20927;
assign w20929 = ~w20917 & ~w20928;
assign w20930 = ~w20919 & ~w20927;
assign w20931 = ~w19836 & ~w19839;
assign w20932 = ~w19507 & ~w19823;
assign w20933 = w20931 & w20932;
assign w20934 = ~w20931 & ~w20932;
assign w20935 = ~w20933 & ~w20934;
assign w20936 = w3 & ~w12878;
assign w20937 = w10835 & w12874;
assign w20938 = ~w20936 & ~w20937;
assign w20939 = (w20938 & ~w13771) | (w20938 & w36649) | (~w13771 & w36649);
assign w20940 = (a_2 & ~w12869) | (a_2 & w34211) | (~w12869 & w34211);
assign w20941 = w20939 & ~w20940;
assign w20942 = (w13771 & w36650) | (w13771 & w36651) | (w36650 & w36651);
assign w20943 = ~w20941 & ~w20942;
assign w20944 = w20935 & ~w20943;
assign w20945 = (~w20930 & ~w20929) | (~w20930 & w31983) | (~w20929 & w31983);
assign w20946 = ~w20944 & w20945;
assign w20947 = ~w20935 & w20943;
assign w20948 = (~w19860 & w19838) | (~w19860 & w31984) | (w19838 & w31984);
assign w20949 = ~w19862 & ~w20948;
assign w20950 = ~w12892 & w36652;
assign w20951 = w10835 & ~w12878;
assign w20952 = ~w20950 & ~w20951;
assign w20953 = (w20952 & ~w13787) | (w20952 & w36653) | (~w13787 & w36653);
assign w20954 = (a_2 & ~w12874) | (a_2 & w34211) | (~w12874 & w34211);
assign w20955 = w20953 & ~w20954;
assign w20956 = (w13787 & w36654) | (w13787 & w36655) | (w36654 & w36655);
assign w20957 = ~w20955 & ~w20956;
assign w20958 = w20949 & w20957;
assign w20959 = ~w20947 & ~w20958;
assign w20960 = ~w20946 & w20959;
assign w20961 = ~w20949 & ~w20957;
assign w20962 = ~w19493 & w19868;
assign w20963 = ~w19862 & ~w19863;
assign w20964 = ~w20962 & w20963;
assign w20965 = w20962 & ~w20963;
assign w20966 = ~w20964 & ~w20965;
assign w20967 = ~w12905 & w36656;
assign w20968 = ~w12892 & w36657;
assign w20969 = ~w13598 & w36658;
assign w20970 = ~w20967 & ~w20968;
assign w20971 = ~w20969 & w20970;
assign w20972 = (a_2 & w12878) | (a_2 & w34211) | (w12878 & w34211);
assign w20973 = w20971 & ~w20972;
assign w20974 = (a_2 & w20969) | (a_2 & w36659) | (w20969 & w36659);
assign w20975 = ~w20973 & ~w20974;
assign w20976 = (~w20961 & w20966) | (~w20961 & w31985) | (w20966 & w31985);
assign w20977 = ~w20960 & w20976;
assign w20978 = w20966 & w20975;
assign w20979 = w19870 & ~w19875;
assign w20980 = ~w19870 & w19875;
assign w20981 = ~w20979 & ~w20980;
assign w20982 = ~w12905 & w36660;
assign w20983 = w3 & ~w12910;
assign w20984 = ~w20982 & ~w20983;
assign w20985 = (w20984 & ~w13815) | (w20984 & w36661) | (~w13815 & w36661);
assign w20986 = (a_2 & ~w12894) | (a_2 & w34211) | (~w12894 & w34211);
assign w20987 = w20985 & ~w20986;
assign w20988 = (w13815 & w36662) | (w13815 & w36663) | (w36662 & w36663);
assign w20989 = ~w20987 & ~w20988;
assign w20990 = w20981 & w20989;
assign w20991 = ~w20978 & ~w20990;
assign w20992 = ~w20977 & w20991;
assign w20993 = (w19475 & ~w19870) | (w19475 & w31986) | (~w19870 & w31986);
assign w20994 = w19458 & w19481;
assign w20995 = ~w12914 & w36664;
assign w20996 = w10835 & ~w12910;
assign w20997 = (w10837 & w13518) | (w10837 & w36665) | (w13518 & w36665);
assign w20998 = ~w20995 & ~w20996;
assign w20999 = ~w12905 & w36666;
assign w21000 = a_2 & ~w20999;
assign w21001 = ~w20997 & w36667;
assign w21002 = (a_2 & w20997) | (a_2 & w36668) | (w20997 & w36668);
assign w21003 = ~w21001 & ~w21002;
assign w21004 = w20993 & w36669;
assign w21005 = w20994 & ~w21003;
assign w21006 = ~w20993 & w21005;
assign w21007 = ~w20981 & ~w20989;
assign w21008 = ~w21006 & ~w21007;
assign w21009 = ~w21004 & w21008;
assign w21010 = ~w20992 & w21009;
assign w21011 = w19878 & ~w19900;
assign w21012 = ~w19901 & ~w21011;
assign w21013 = ~w12930 & w36670;
assign w21014 = ~w12914 & w36671;
assign w21015 = ~w13501 & w36672;
assign w21016 = ~w21013 & ~w21014;
assign w21017 = ~w21015 & w21016;
assign w21018 = (a_2 & w12910) | (a_2 & w34211) | (w12910 & w34211);
assign w21019 = w21017 & ~w21018;
assign w21020 = (a_2 & w21015) | (a_2 & w36673) | (w21015 & w36673);
assign w21021 = ~w21019 & ~w21020;
assign w21022 = ~w20993 & w20994;
assign w21023 = (w21003 & ~w20993) | (w21003 & w36674) | (~w20993 & w36674);
assign w21024 = ~w21022 & w21023;
assign w21025 = (~w21024 & ~w21012) | (~w21024 & w36675) | (~w21012 & w36675);
assign w21026 = ~w21010 & w21025;
assign w21027 = (~w19917 & w19878) | (~w19917 & w37579) | (w19878 & w37579);
assign w21028 = w19914 & w19924;
assign w21029 = (w3 & w12612) | (w3 & w36676) | (w12612 & w36676);
assign w21030 = ~w12930 & w36677;
assign w21031 = ~w21029 & ~w21030;
assign w21032 = (w21031 & ~w13375) | (w21031 & w36678) | (~w13375 & w36678);
assign w21033 = (a_2 & ~w12916) | (a_2 & w34211) | (~w12916 & w34211);
assign w21034 = w21032 & ~w21033;
assign w21035 = (w13375 & w36679) | (w13375 & w36680) | (w36679 & w36680);
assign w21036 = ~w21034 & ~w21035;
assign w21037 = w21027 & w31987;
assign w21038 = w21028 & ~w21036;
assign w21039 = ~w21027 & w21038;
assign w21040 = ~w21012 & ~w21021;
assign w21041 = ~w21039 & ~w21040;
assign w21042 = ~w21037 & w21041;
assign w21043 = ~w21026 & w21042;
assign w21044 = (w3 & w12616) | (w3 & w36681) | (w12616 & w36681);
assign w21045 = (w10835 & w12612) | (w10835 & w36682) | (w12612 & w36682);
assign w21046 = ~w21044 & ~w21045;
assign w21047 = (w21046 & ~w13389) | (w21046 & w36683) | (~w13389 & w36683);
assign w21048 = (a_2 & ~w12931) | (a_2 & w34211) | (~w12931 & w34211);
assign w21049 = w21047 & ~w21048;
assign w21050 = (w13389 & w36684) | (w13389 & w36685) | (w36684 & w36685);
assign w21051 = ~w21049 & ~w21050;
assign w21052 = w19947 & w21051;
assign w21053 = w19925 & w21052;
assign w21054 = ~w19947 & w21051;
assign w21055 = ~w19925 & w21054;
assign w21056 = ~w21027 & w21028;
assign w21057 = (w21036 & ~w21027) | (w21036 & w31988) | (~w21027 & w31988);
assign w21058 = ~w21056 & w21057;
assign w21059 = ~w21053 & ~w21055;
assign w21060 = ~w21058 & w21059;
assign w21061 = ~w21043 & w21060;
assign w21062 = w19931 & w19942;
assign w21063 = w19932 & ~w19941;
assign w21064 = ~w19931 & w21063;
assign w21065 = w19924 & ~w21062;
assign w21066 = ~w21064 & w21065;
assign w21067 = ~w19919 & w21066;
assign w21068 = ~w19949 & ~w21067;
assign w21069 = ~w19963 & ~w19967;
assign w21070 = ~w21068 & w21069;
assign w21071 = (w10835 & w12616) | (w10835 & w36686) | (w12616 & w36686);
assign w21072 = ~w12589 & w36687;
assign w21073 = ~w21071 & ~w21072;
assign w21074 = (w21073 & ~w13123) | (w21073 & w36688) | (~w13123 & w36688);
assign w21075 = (a_2 & w12613) | (a_2 & w34211) | (w12613 & w34211);
assign w21076 = w21074 & ~w21075;
assign w21077 = (w13123 & w36689) | (w13123 & w36690) | (w36689 & w36690);
assign w21078 = ~w21076 & ~w21077;
assign w21079 = w21070 & ~w21078;
assign w21080 = w19947 & ~w21051;
assign w21081 = ~w19925 & w21080;
assign w21082 = ~w19947 & ~w21051;
assign w21083 = w19925 & w21082;
assign w21084 = w19958 & ~w21078;
assign w21085 = w19962 & ~w21084;
assign w21086 = ~w19958 & ~w21078;
assign w21087 = ~w19962 & ~w21086;
assign w21088 = ~w21085 & ~w21087;
assign w21089 = w21068 & w21088;
assign w21090 = ~w21081 & ~w21083;
assign w21091 = ~w21089 & w21090;
assign w21092 = ~w21079 & w21091;
assign w21093 = ~w21061 & w21092;
assign w21094 = w21068 & ~w21069;
assign w21095 = ~w21070 & w21078;
assign w21096 = ~w21094 & w21095;
assign w21097 = ~w21093 & ~w21096;
assign w21098 = ~w19965 & ~w19967;
assign w21099 = w3 & w12604;
assign w21100 = ~w12589 & w36691;
assign w21101 = ~w21099 & ~w21100;
assign w21102 = (w21101 & w13288) | (w21101 & w36692) | (w13288 & w36692);
assign w21103 = (a_2 & w12617) | (a_2 & w34211) | (w12617 & w34211);
assign w21104 = w21102 & ~w21103;
assign w21105 = (~w13288 & w36693) | (~w13288 & w36694) | (w36693 & w36694);
assign w21106 = ~w21104 & ~w21105;
assign w21107 = w19443 & ~w21106;
assign w21108 = ~w19443 & w21106;
assign w21109 = ~w21107 & ~w21108;
assign w21110 = w21098 & ~w21109;
assign w21111 = ~w21098 & w21109;
assign w21112 = ~w21110 & ~w21111;
assign w21113 = ~w21097 & w21112;
assign w21114 = w21106 & ~w21112;
assign w21115 = w3 & w12601;
assign w21116 = w10835 & w12604;
assign w21117 = ~w21115 & ~w21116;
assign w21118 = (w21117 & w13140) | (w21117 & w36695) | (w13140 & w36695);
assign w21119 = (a_2 & ~w12607) | (a_2 & w34211) | (~w12607 & w34211);
assign w21120 = w21118 & ~w21119;
assign w21121 = (~w13140 & w36696) | (~w13140 & w36697) | (w36696 & w36697);
assign w21122 = ~w21120 & ~w21121;
assign w21123 = w19423 & w21122;
assign w21124 = w19414 & ~w21123;
assign w21125 = ~w19423 & w21122;
assign w21126 = ~w19414 & ~w21125;
assign w21127 = ~w21124 & ~w21126;
assign w21128 = ~w19976 & ~w21127;
assign w21129 = w19414 & ~w21125;
assign w21130 = ~w19414 & ~w21123;
assign w21131 = ~w21129 & ~w21130;
assign w21132 = w19976 & ~w21131;
assign w21133 = ~w21128 & ~w21132;
assign w21134 = ~w21114 & ~w21133;
assign w21135 = ~w21113 & w21134;
assign w21136 = ~w19424 & ~w19977;
assign w21137 = w19976 & ~w21136;
assign w21138 = ~w19976 & w21136;
assign w21139 = ~w21137 & ~w21138;
assign w21140 = ~w21122 & ~w21139;
assign w21141 = ~w21135 & ~w21140;
assign w21142 = w3 & w12598;
assign w21143 = w10835 & w12601;
assign w21144 = ~w21142 & ~w21143;
assign w21145 = (w21144 & ~w12961) | (w21144 & w36698) | (~w12961 & w36698);
assign w21146 = (a_2 & ~w12604) | (a_2 & w34211) | (~w12604 & w34211);
assign w21147 = w21145 & ~w21146;
assign w21148 = (w12961 & w36699) | (w12961 & w36700) | (w36699 & w36700);
assign w21149 = ~w21147 & ~w21148;
assign w21150 = w20177 & ~w21149;
assign w21151 = ~w20177 & w21149;
assign w21152 = ~w21150 & ~w21151;
assign w21153 = w19979 & ~w21152;
assign w21154 = ~w19979 & w21152;
assign w21155 = ~w21153 & ~w21154;
assign w21156 = w21141 & w21155;
assign w21157 = w20177 & w20183;
assign w21158 = ~w19424 & w20183;
assign w21159 = ~w19978 & w21158;
assign w21160 = ~w21157 & ~w21159;
assign w21161 = ~w13011 & w36701;
assign w21162 = w10835 & w12598;
assign w21163 = ~w21161 & ~w21162;
assign w21164 = (w21163 & w13021) | (w21163 & w36702) | (w13021 & w36702);
assign w21165 = (a_2 & ~w12601) | (a_2 & w34211) | (~w12601 & w34211);
assign w21166 = w21164 & ~w21165;
assign w21167 = (~w13021 & w36703) | (~w13021 & w36704) | (w36703 & w36704);
assign w21168 = ~w21166 & ~w21167;
assign w21169 = ~w20188 & w21168;
assign w21170 = ~w21160 & ~w21169;
assign w21171 = w20188 & w21168;
assign w21172 = w21160 & ~w21171;
assign w21173 = ~w21170 & ~w21172;
assign w21174 = w19979 & ~w20177;
assign w21175 = ~w19979 & w20177;
assign w21176 = ~w21174 & ~w21175;
assign w21177 = w21149 & ~w21176;
assign w21178 = ~w21173 & ~w21177;
assign w21179 = ~w21156 & w21178;
assign w21180 = w20188 & ~w21168;
assign w21181 = ~w21169 & ~w21180;
assign w21182 = w21160 & w21181;
assign w21183 = ~w21160 & ~w21181;
assign w21184 = ~w21182 & ~w21183;
assign w21185 = ~w21173 & ~w21184;
assign w21186 = ~w13174 & w36705;
assign w21187 = ~w13011 & w36706;
assign w21188 = ~w13205 & w36707;
assign w21189 = ~w21186 & ~w21187;
assign w21190 = ~w21188 & w21189;
assign w21191 = (a_2 & ~w12598) | (a_2 & w34211) | (~w12598 & w34211);
assign w21192 = w21190 & ~w21191;
assign w21193 = (a_2 & w21188) | (a_2 & w36708) | (w21188 & w36708);
assign w21194 = ~w21192 & ~w21193;
assign w21195 = ~w20388 & ~w21194;
assign w21196 = w20191 & w21195;
assign w21197 = w20388 & ~w21194;
assign w21198 = ~w20191 & w21197;
assign w21199 = ~w21196 & ~w21198;
assign w21200 = ~w21185 & w21199;
assign w21201 = ~w21179 & w21200;
assign w21202 = w20388 & w21194;
assign w21203 = w20191 & w21202;
assign w21204 = ~w20388 & w21194;
assign w21205 = ~w20191 & w21204;
assign w21206 = ~w21203 & ~w21205;
assign w21207 = ~w21201 & w21206;
assign w21208 = ~w20191 & w20388;
assign w21209 = (~w20391 & w20191) | (~w20391 & w31989) | (w20191 & w31989);
assign w21210 = w20372 & w20396;
assign w21211 = w3 & w13177;
assign w21212 = ~w13174 & w36709;
assign w21213 = ~w21211 & ~w21212;
assign w21214 = (w21213 & ~w13207) | (w21213 & w36710) | (~w13207 & w36710);
assign w21215 = (a_2 & ~w13013) | (a_2 & w34211) | (~w13013 & w34211);
assign w21216 = w21214 & ~w21215;
assign w21217 = (w13207 & w36711) | (w13207 & w36712) | (w36711 & w36712);
assign w21218 = ~w21216 & ~w21217;
assign w21219 = w20372 & w36713;
assign w21220 = (w21218 & ~w20372) | (w21218 & w36714) | (~w20372 & w36714);
assign w21221 = ~w21219 & ~w21220;
assign w21222 = w21209 & ~w21221;
assign w21223 = ~w21209 & w21221;
assign w21224 = ~w21222 & ~w21223;
assign w21225 = (~w21224 & w21201) | (~w21224 & w36715) | (w21201 & w36715);
assign w21226 = ~w21209 & w21220;
assign w21227 = (w21218 & w20388) | (w21218 & w31990) | (w20388 & w31990);
assign w21228 = w21210 & w21227;
assign w21229 = ~w21208 & w21228;
assign w21230 = ~w21226 & ~w21229;
assign w21231 = (w21230 & w21207) | (w21230 & w31991) | (w21207 & w31991);
assign w21232 = ~w20508 & ~w20631;
assign w21233 = w20399 & w21232;
assign w21234 = w20508 & ~w20631;
assign w21235 = ~w20399 & w21234;
assign w21236 = ~w21233 & ~w21235;
assign w21237 = w20636 & w21236;
assign w21238 = w20643 & w21237;
assign w21239 = ~w21231 & w21238;
assign w21240 = ~w20644 & ~w21239;
assign w21241 = ~w20520 & w20605;
assign w21242 = ~w20519 & w21241;
assign w21243 = ~w20529 & ~w21242;
assign w21244 = ~w20610 & w21243;
assign w21245 = ~w20513 & ~w21244;
assign w21246 = ~w20509 & w21245;
assign w21247 = w20611 & ~w21243;
assign w21248 = ~w21246 & ~w21247;
assign w21249 = (w13173 & w36718) | (w13173 & w36719) | (w36718 & w36719);
assign w21250 = w20587 & ~w20605;
assign w21251 = ~w21242 & ~w21250;
assign w21252 = w20575 & ~w20596;
assign w21253 = w20540 & ~w21252;
assign w21254 = ~w20575 & ~w20596;
assign w21255 = ~w20540 & ~w21254;
assign w21256 = ~w21253 & ~w21255;
assign w21257 = ~w20478 & ~w21256;
assign w21258 = ~w20415 & w21257;
assign w21259 = w20533 & ~w20596;
assign w21260 = ~w20533 & w20596;
assign w21261 = ~w20578 & ~w21260;
assign w21262 = ~w21259 & ~w21261;
assign w21263 = ~w21258 & ~w21262;
assign w21264 = w20566 & w20572;
assign w21265 = w20545 & w21264;
assign w21266 = w20566 & ~w20572;
assign w21267 = ~w20545 & w21266;
assign w21268 = ~w21265 & ~w21267;
assign w21269 = (w21268 & w20539) | (w21268 & w36720) | (w20539 & w36720);
assign w21270 = ~w17544 & ~w20555;
assign w21271 = ~w17153 & w20554;
assign w21272 = w17544 & ~w21271;
assign w21273 = ~w21270 & ~w21272;
assign w21274 = ~w20452 & ~w21273;
assign w21275 = w20423 & w21274;
assign w21276 = w17153 & ~w20554;
assign w21277 = w17544 & ~w21276;
assign w21278 = ~w17544 & ~w20556;
assign w21279 = ~w21277 & ~w21278;
assign w21280 = w20544 & ~w21279;
assign w21281 = ~w21273 & ~w21280;
assign w21282 = ~w21275 & ~w21281;
assign w21283 = ~w12930 & w36721;
assign w21284 = w6446 & ~w12910;
assign w21285 = ~w12914 & w36722;
assign w21286 = ~w13501 & w36723;
assign w21287 = ~w21284 & ~w21285;
assign w21288 = ~w21283 & w21287;
assign w21289 = ~w21286 & w36724;
assign w21290 = (a_14 & w21286) | (a_14 & w36725) | (w21286 & w36725);
assign w21291 = ~w21289 & ~w21290;
assign w21292 = w17133 & w17138;
assign w21293 = ~w12905 & w36726;
assign w21294 = ~w12892 & w36727;
assign w21295 = w6059 & ~w12878;
assign w21296 = ~w13598 & w36728;
assign w21297 = ~w21294 & ~w21295;
assign w21298 = ~w21293 & w21297;
assign w21299 = ~w21296 & w36729;
assign w21300 = (a_17 & w21296) | (a_17 & w36730) | (w21296 & w36730);
assign w21301 = ~w21299 & ~w21300;
assign w21302 = w21292 & ~w21301;
assign w21303 = ~w21292 & w21301;
assign w21304 = ~w21302 & ~w21303;
assign w21305 = w17545 & w21304;
assign w21306 = ~w17545 & ~w21304;
assign w21307 = ~w21305 & ~w21306;
assign w21308 = ~w21291 & w21307;
assign w21309 = w21282 & w21308;
assign w21310 = ~w21291 & ~w21307;
assign w21311 = ~w21282 & w21310;
assign w21312 = ~w21309 & ~w21311;
assign w21313 = w21291 & ~w21307;
assign w21314 = w21282 & w21313;
assign w21315 = w21291 & w21307;
assign w21316 = ~w21282 & w21315;
assign w21317 = ~w21314 & ~w21316;
assign w21318 = w21312 & w21317;
assign w21319 = (w7489 & w12616) | (w7489 & w36731) | (w12616 & w36731);
assign w21320 = (w7192 & w12612) | (w7192 & w36732) | (w12612 & w36732);
assign w21321 = ~w12589 & w36733;
assign w21322 = ~w21319 & ~w21320;
assign w21323 = ~w21321 & w21322;
assign w21324 = (w21323 & ~w13123) | (w21323 & w36734) | (~w13123 & w36734);
assign w21325 = ~a_11 & w21324;
assign w21326 = (w13123 & w36735) | (w13123 & w36736) | (w36735 & w36736);
assign w21327 = ~w21325 & ~w21326;
assign w21328 = w21318 & ~w21327;
assign w21329 = ~w21318 & w21327;
assign w21330 = ~w21328 & ~w21329;
assign w21331 = w21269 & w21330;
assign w21332 = ~w21269 & ~w21330;
assign w21333 = ~w21331 & ~w21332;
assign w21334 = w21263 & ~w21333;
assign w21335 = ~w21263 & w21333;
assign w21336 = ~w21334 & ~w21335;
assign w21337 = w8295 & w12598;
assign w21338 = w8298 & w12601;
assign w21339 = w8277 & w12604;
assign w21340 = ~w21338 & ~w21339;
assign w21341 = ~w21337 & w21340;
assign w21342 = (w21341 & ~w12961) | (w21341 & w36737) | (~w12961 & w36737);
assign w21343 = ~a_8 & w21342;
assign w21344 = (w12961 & w36738) | (w12961 & w36739) | (w36738 & w36739);
assign w21345 = ~w21343 & ~w21344;
assign w21346 = ~w13174 & w36740;
assign w21347 = ~w13011 & w36741;
assign w21348 = w9788 & w13177;
assign w21349 = ~w21346 & ~w21347;
assign w21350 = (a_5 & ~w21349) | (a_5 & w36742) | (~w21349 & w36742);
assign w21351 = w10061 & w13207;
assign w21352 = w21349 & w36743;
assign w21353 = ~w21351 & w21352;
assign w21354 = (~w21350 & ~w13207) | (~w21350 & w36744) | (~w13207 & w36744);
assign w21355 = ~w21353 & w21354;
assign w21356 = (w21345 & w21353) | (w21345 & w36745) | (w21353 & w36745);
assign w21357 = ~w21353 & w36746;
assign w21358 = ~w21356 & ~w21357;
assign w21359 = w21336 & ~w21358;
assign w21360 = ~w21336 & w21358;
assign w21361 = ~w21359 & ~w21360;
assign w21362 = w21251 & w21361;
assign w21363 = ~w21251 & ~w21361;
assign w21364 = ~w21362 & ~w21363;
assign w21365 = w21249 & w21364;
assign w21366 = ~w21249 & ~w21364;
assign w21367 = ~w21365 & ~w21366;
assign w21368 = w21248 & ~w21367;
assign w21369 = ~w21248 & w21367;
assign w21370 = ~w21368 & ~w21369;
assign w21371 = ~w21247 & ~w21364;
assign w21372 = ~w21246 & w21371;
assign w21373 = w21355 & w21364;
assign w21374 = ~w21372 & ~w21373;
assign w21375 = ~w21336 & ~w21345;
assign w21376 = w21333 & w21345;
assign w21377 = w21263 & ~w21376;
assign w21378 = ~w21333 & w21345;
assign w21379 = ~w21263 & ~w21378;
assign w21380 = ~w21377 & ~w21379;
assign w21381 = ~w21250 & ~w21380;
assign w21382 = ~w21242 & w21381;
assign w21383 = ~w21375 & ~w21382;
assign w21384 = w21327 & ~w21333;
assign w21385 = ~w21335 & ~w21384;
assign w21386 = w10033 & ~w13264;
assign w21387 = (w13173 & w36747) | (w13173 & w36748) | (w36747 & w36748);
assign w21388 = ~w13174 & w36749;
assign w21389 = w9780 & w13177;
assign w21390 = ~w21387 & ~w21388;
assign w21391 = ~w21389 & w21390;
assign w21392 = a_5 & w21391;
assign w21393 = ~a_5 & ~w21391;
assign w21394 = ~w21392 & ~w21393;
assign w21395 = (w21394 & w13264) | (w21394 & w36750) | (w13264 & w36750);
assign w21396 = ~w21386 & ~w21395;
assign w21397 = w21268 & w21317;
assign w21398 = w21312 & ~w21397;
assign w21399 = w20575 & w21312;
assign w21400 = w20540 & w21399;
assign w21401 = ~w21398 & ~w21400;
assign w21402 = ~w21282 & ~w21307;
assign w21403 = w21301 & w21307;
assign w21404 = ~w21402 & ~w21403;
assign w21405 = (w6996 & w12612) | (w6996 & w36751) | (w12612 & w36751);
assign w21406 = ~w12914 & w36752;
assign w21407 = ~w12930 & w36753;
assign w21408 = ~w21406 & ~w21407;
assign w21409 = ~w21405 & w21408;
assign w21410 = (w21409 & ~w13375) | (w21409 & w36754) | (~w13375 & w36754);
assign w21411 = ~a_14 & w21410;
assign w21412 = (w13375 & w36755) | (w13375 & w36756) | (w36755 & w36756);
assign w21413 = ~w21411 & ~w21412;
assign w21414 = ~w12905 & w36757;
assign w21415 = w6304 & ~w12910;
assign w21416 = ~w12892 & w36758;
assign w21417 = w6063 & w13815;
assign w21418 = ~w21415 & w36759;
assign w21419 = ~w21417 & w36760;
assign w21420 = (a_17 & w21417) | (a_17 & w36761) | (w21417 & w36761);
assign w21421 = ~w21419 & ~w21420;
assign w21422 = ~w17561 & w21421;
assign w21423 = w17561 & ~w21421;
assign w21424 = ~w21422 & ~w21423;
assign w21425 = w17546 & w21424;
assign w21426 = ~w17546 & ~w21424;
assign w21427 = ~w21425 & ~w21426;
assign w21428 = w21413 & ~w21427;
assign w21429 = ~w21413 & w21427;
assign w21430 = ~w21428 & ~w21429;
assign w21431 = w21404 & w21430;
assign w21432 = ~w21404 & ~w21430;
assign w21433 = ~w21431 & ~w21432;
assign w21434 = w21401 & ~w21433;
assign w21435 = ~w21401 & w21433;
assign w21436 = ~w21434 & ~w21435;
assign w21437 = w7511 & w12604;
assign w21438 = ~w12589 & w36762;
assign w21439 = (w7192 & w12616) | (w7192 & w36763) | (w12616 & w36763);
assign w21440 = ~w21438 & ~w21439;
assign w21441 = ~w21437 & w21440;
assign w21442 = (w21441 & w13288) | (w21441 & w36764) | (w13288 & w36764);
assign w21443 = a_11 & ~w21442;
assign w21444 = (w13288 & w36765) | (w13288 & w36766) | (w36765 & w36766);
assign w21445 = ~w21443 & ~w21444;
assign w21446 = w8298 & w12598;
assign w21447 = w8277 & w12601;
assign w21448 = ~w13011 & w36767;
assign w21449 = ~w21446 & ~w21447;
assign w21450 = ~w21448 & w21449;
assign w21451 = (w21450 & w13021) | (w21450 & w36768) | (w13021 & w36768);
assign w21452 = a_8 & ~w21451;
assign w21453 = (w13021 & w36769) | (w13021 & w36770) | (w36769 & w36770);
assign w21454 = ~w21452 & ~w21453;
assign w21455 = w21445 & w21454;
assign w21456 = ~w21445 & ~w21454;
assign w21457 = ~w21455 & ~w21456;
assign w21458 = w21436 & w21457;
assign w21459 = ~w21436 & ~w21457;
assign w21460 = ~w21458 & ~w21459;
assign w21461 = w21396 & ~w21460;
assign w21462 = ~w21396 & w21460;
assign w21463 = ~w21461 & ~w21462;
assign w21464 = w21385 & ~w21463;
assign w21465 = ~w21385 & w21463;
assign w21466 = ~w21464 & ~w21465;
assign w21467 = w21383 & w21466;
assign w21468 = ~w21383 & ~w21466;
assign w21469 = ~w21467 & ~w21468;
assign w21470 = w14339 & ~w21469;
assign w21471 = ~w14339 & w21469;
assign w21472 = ~w21470 & ~w21471;
assign w21473 = w21374 & ~w21472;
assign w21474 = ~w21370 & ~w21473;
assign w21475 = ~w21240 & w21474;
assign w21476 = ~w21374 & w21472;
assign w21477 = ~w21249 & ~w21372;
assign w21478 = ~w21369 & w21477;
assign w21479 = ~w21476 & ~w21478;
assign w21480 = ~w21473 & ~w21479;
assign w21481 = w21396 & w21469;
assign w21482 = ~w21470 & ~w21481;
assign w21483 = w21436 & w21445;
assign w21484 = ~w21384 & ~w21483;
assign w21485 = ~w21335 & w21484;
assign w21486 = ~w21436 & ~w21445;
assign w21487 = ~w21485 & ~w21486;
assign w21488 = w21413 & ~w21433;
assign w21489 = ~w17120 & ~w17564;
assign w21490 = ~w17565 & ~w21489;
assign w21491 = w8564 & w13389;
assign w21492 = (w6998 & w12612) | (w6998 & w36771) | (w12612 & w36771);
assign w21493 = ~w12930 & w36772;
assign w21494 = (w6996 & w12616) | (w6996 & w36773) | (w12616 & w36773);
assign w21495 = ~w21492 & ~w21493;
assign w21496 = ~w21494 & w21495;
assign w21497 = a_14 & ~w21496;
assign w21498 = ~a_14 & w21496;
assign w21499 = (w21498 & ~w13389) | (w21498 & w36774) | (~w13389 & w36774);
assign w21500 = ~w21491 & ~w21497;
assign w21501 = ~w21499 & w21500;
assign w21502 = ~w21490 & ~w21501;
assign w21503 = w21490 & w21501;
assign w21504 = ~w21502 & ~w21503;
assign w21505 = ~w21421 & ~w21427;
assign w21506 = ~w21402 & w36775;
assign w21507 = ~w21505 & ~w21506;
assign w21508 = w21504 & ~w21507;
assign w21509 = ~w21504 & w21507;
assign w21510 = ~w21508 & ~w21509;
assign w21511 = (~w21510 & w21435) | (~w21510 & w36776) | (w21435 & w36776);
assign w21512 = ~w21435 & w36777;
assign w21513 = ~w21511 & ~w21512;
assign w21514 = ~w13174 & w36778;
assign w21515 = ~w13011 & w36779;
assign w21516 = w8277 & w12598;
assign w21517 = ~w13205 & w36780;
assign w21518 = ~w21515 & w36781;
assign w21519 = (a_8 & w21517) | (a_8 & w36782) | (w21517 & w36782);
assign w21520 = ~w21517 & w36783;
assign w21521 = ~w21519 & ~w21520;
assign w21522 = w7511 & w12601;
assign w21523 = w7489 & w12604;
assign w21524 = ~w12589 & w36784;
assign w21525 = ~w21523 & ~w21524;
assign w21526 = ~w21522 & w21525;
assign w21527 = (w21526 & w13140) | (w21526 & w36785) | (w13140 & w36785);
assign w21528 = a_11 & ~w21527;
assign w21529 = (w13140 & w36786) | (w13140 & w36787) | (w36786 & w36787);
assign w21530 = ~w21528 & ~w21529;
assign w21531 = w21521 & ~w21530;
assign w21532 = ~w21521 & w21530;
assign w21533 = ~w21531 & ~w21532;
assign w21534 = w21513 & w21533;
assign w21535 = ~w21513 & ~w21533;
assign w21536 = ~w21534 & ~w21535;
assign w21537 = w21487 & ~w21536;
assign w21538 = ~w21487 & w21536;
assign w21539 = ~w21537 & ~w21538;
assign w21540 = w9786 & w13177;
assign w21541 = (w13201 & w36790) | (w13201 & w36791) | (w36790 & w36791);
assign w21542 = (~w13173 & w36792) | (~w13173 & w36793) | (w36792 & w36793);
assign w21543 = ~w21540 & w21542;
assign w21544 = (a_5 & w21541) | (a_5 & w36794) | (w21541 & w36794);
assign w21545 = ~w21541 & w36795;
assign w21546 = ~w21544 & ~w21545;
assign w21547 = w21539 & w21546;
assign w21548 = ~w21539 & ~w21546;
assign w21549 = ~w21547 & ~w21548;
assign w21550 = w21385 & ~w21460;
assign w21551 = ~w21385 & w21460;
assign w21552 = ~w21550 & ~w21551;
assign w21553 = w21454 & ~w21552;
assign w21554 = ~w21382 & w36796;
assign w21555 = ~w21553 & ~w21554;
assign w21556 = w21549 & ~w21555;
assign w21557 = ~w21549 & w21555;
assign w21558 = ~w21556 & ~w21557;
assign w21559 = ~w21482 & w21558;
assign w21560 = w21521 & w21536;
assign w21561 = (~w21502 & w21507) | (~w21502 & w36797) | (w21507 & w36797);
assign w21562 = ~w17571 & ~w17580;
assign w21563 = ~w17581 & ~w21562;
assign w21564 = w21561 & ~w21563;
assign w21565 = ~w21561 & w21563;
assign w21566 = ~w21564 & ~w21565;
assign w21567 = w7511 & w12598;
assign w21568 = w7489 & w12601;
assign w21569 = w7192 & w12604;
assign w21570 = ~w21568 & ~w21569;
assign w21571 = ~w21567 & w21570;
assign w21572 = (w21571 & ~w12961) | (w21571 & w36798) | (~w12961 & w36798);
assign w21573 = a_11 & ~w21572;
assign w21574 = (~w12961 & w36799) | (~w12961 & w36800) | (w36799 & w36800);
assign w21575 = ~w21573 & ~w21574;
assign w21576 = ~w13174 & w36801;
assign w21577 = ~w13011 & w36802;
assign w21578 = w8295 & w13177;
assign w21579 = ~w21576 & ~w21577;
assign w21580 = ~w21578 & w21579;
assign w21581 = (w21580 & ~w13207) | (w21580 & w36803) | (~w13207 & w36803);
assign w21582 = a_8 & ~w21581;
assign w21583 = (~w13207 & w36804) | (~w13207 & w36805) | (w36804 & w36805);
assign w21584 = ~w21582 & ~w21583;
assign w21585 = (w21575 & w21582) | (w21575 & w36806) | (w21582 & w36806);
assign w21586 = ~w21582 & w36807;
assign w21587 = ~w21585 & ~w21586;
assign w21588 = w21566 & w21587;
assign w21589 = ~w21566 & ~w21587;
assign w21590 = ~w21588 & ~w21589;
assign w21591 = ~w21511 & ~w21530;
assign w21592 = ~w21512 & ~w21591;
assign w21593 = ~w21590 & w21592;
assign w21594 = w21590 & ~w21592;
assign w21595 = ~w21593 & ~w21594;
assign w21596 = ~w21537 & w36808;
assign w21597 = (w21595 & w21537) | (w21595 & w36809) | (w21537 & w36809);
assign w21598 = ~w21596 & ~w21597;
assign w21599 = (~w13173 & w36812) | (~w13173 & w36813) | (w36812 & w36813);
assign w21600 = (~w13173 & w36814) | (~w13173 & w36815) | (w36814 & w36815);
assign w21601 = ~w21599 & w21600;
assign w21602 = ~w14377 & ~w21601;
assign w21603 = w21598 & ~w21602;
assign w21604 = ~w21598 & w21602;
assign w21605 = ~w21603 & ~w21604;
assign w21606 = ~w21547 & ~w21556;
assign w21607 = ~w21605 & ~w21606;
assign w21608 = ~w17587 & w17596;
assign w21609 = ~w17597 & ~w21608;
assign w21610 = ~w21564 & ~w21575;
assign w21611 = ~w21565 & ~w21610;
assign w21612 = w21609 & ~w21611;
assign w21613 = ~w21609 & w21611;
assign w21614 = ~w21612 & ~w21613;
assign w21615 = w8298 & w13177;
assign w21616 = ~w13174 & w36816;
assign w21617 = (w13173 & w36817) | (w13173 & w36818) | (w36817 & w36818);
assign w21618 = ~w21616 & ~w21617;
assign w21619 = ~w21615 & w21618;
assign w21620 = (w21619 & w13264) | (w21619 & w36819) | (w13264 & w36819);
assign w21621 = a_8 & ~w21620;
assign w21622 = (w13264 & w36820) | (w13264 & w36821) | (w36820 & w36821);
assign w21623 = ~w21621 & ~w21622;
assign w21624 = w21614 & w21623;
assign w21625 = ~w21614 & ~w21623;
assign w21626 = ~w21624 & ~w21625;
assign w21627 = w21584 & w21590;
assign w21628 = (w14379 & w21593) | (w14379 & w36822) | (w21593 & w36822);
assign w21629 = ~w21593 & w36823;
assign w21630 = ~w21628 & ~w21629;
assign w21631 = w21626 & w21630;
assign w21632 = ~w21626 & ~w21630;
assign w21633 = ~w21631 & ~w21632;
assign w21634 = (~w21596 & ~w21598) | (~w21596 & w31992) | (~w21598 & w31992);
assign w21635 = w21633 & w21634;
assign w21636 = (~w21635 & w21606) | (~w21635 & w36824) | (w21606 & w36824);
assign w21637 = ~w21559 & w21636;
assign w21638 = ~w21480 & w21637;
assign w21639 = ~w21475 & w21638;
assign w21640 = w21482 & ~w21558;
assign w21641 = w21605 & w21606;
assign w21642 = ~w21607 & ~w21641;
assign w21643 = ~w21640 & w21642;
assign w21644 = (~w21628 & ~w21630) | (~w21628 & w36825) | (~w21630 & w36825);
assign w21645 = (~w21613 & ~w21614) | (~w21613 & w36826) | (~w21614 & w36826);
assign w21646 = w8277 & w13177;
assign w21647 = (w13201 & w36829) | (w13201 & w36830) | (w36829 & w36830);
assign w21648 = (~w13173 & w36831) | (~w13173 & w36832) | (w36831 & w36832);
assign w21649 = ~w21646 & w21648;
assign w21650 = (a_8 & w21647) | (a_8 & w36833) | (w21647 & w36833);
assign w21651 = ~w21647 & w36834;
assign w21652 = ~w21650 & ~w21651;
assign w21653 = ~w17105 & ~w17106;
assign w21654 = w17598 & ~w21653;
assign w21655 = ~w17598 & w21653;
assign w21656 = ~w21654 & ~w21655;
assign w21657 = ~w21652 & w21656;
assign w21658 = w21652 & ~w21656;
assign w21659 = ~w21657 & ~w21658;
assign w21660 = w21645 & ~w21659;
assign w21661 = ~w21645 & w21659;
assign w21662 = ~w21660 & ~w21661;
assign w21663 = w21644 & ~w21662;
assign w21664 = ~w17602 & ~w17606;
assign w21665 = ~w17607 & ~w21664;
assign w21666 = (~w21658 & w21645) | (~w21658 & w36835) | (w21645 & w36835);
assign w21667 = w21665 & ~w21666;
assign w21668 = ~w21665 & w21666;
assign w21669 = ~w21667 & ~w21668;
assign w21670 = ~w21633 & ~w21634;
assign w21671 = (~w21663 & w21634) | (~w21663 & w36836) | (w21634 & w36836);
assign w21672 = w21669 & w21671;
assign w21673 = (w21672 & w21643) | (w21672 & w32455) | (w21643 & w32455);
assign w21674 = (w21673 & ~w21638) | (w21673 & w36837) | (~w21638 & w36837);
assign w21675 = ~w21644 & w21662;
assign w21676 = w21669 & w21675;
assign w21677 = (~w21667 & ~w21675) | (~w21667 & w36838) | (~w21675 & w36838);
assign w21678 = ~w17608 & w17610;
assign w21679 = ~w17090 & ~w21678;
assign w21680 = w21677 & w21679;
assign w21681 = w17633 & ~w17637;
assign w21682 = ~w15832 & w15834;
assign w21683 = ~w17634 & w17636;
assign w21684 = ~w17637 & ~w21683;
assign w21685 = ~w17629 & w21684;
assign w21686 = ~w17637 & ~w21685;
assign w21687 = (~w21682 & w21685) | (~w21682 & w36839) | (w21685 & w36839);
assign w21688 = (w21639 & w36840) | (w21639 & w36841) | (w36840 & w36841);
assign w21689 = ~w15839 & w36842;
assign w21690 = ~w14872 & ~w14884;
assign w21691 = w15844 & w21690;
assign w21692 = w14890 & ~w21691;
assign w21693 = w14880 & ~w14882;
assign w21694 = w14885 & ~w14887;
assign w21695 = ~w14883 & ~w21693;
assign w21696 = w21694 & w21695;
assign w21697 = ~w21693 & ~w21696;
assign w21698 = w14315 & ~w14317;
assign w21699 = ~w14318 & ~w21698;
assign w21700 = ~w14229 & w21699;
assign w21701 = ~w21696 & w36846;
assign w21702 = ~w14205 & ~w14226;
assign w21703 = w13707 & ~w13709;
assign w21704 = ~w13710 & ~w21703;
assign w21705 = (~w14212 & ~w14213) | (~w14212 & w36851) | (~w14213 & w36851);
assign w21706 = w5016 & w13177;
assign w21707 = (w13173 & w36852) | (w13173 & w36853) | (w36852 & w36853);
assign w21708 = (w13201 & w36854) | (w13201 & w36855) | (w36854 & w36855);
assign w21709 = ~w5286 & ~w21707;
assign w21710 = ~w21706 & w21709;
assign w21711 = (a_23 & w21708) | (a_23 & w36856) | (w21708 & w36856);
assign w21712 = ~w21708 & w36857;
assign w21713 = ~w21711 & ~w21712;
assign w21714 = w21705 & ~w21713;
assign w21715 = ~w21705 & w21713;
assign w21716 = ~w21714 & ~w21715;
assign w21717 = w21704 & w21716;
assign w21718 = ~w21704 & ~w21716;
assign w21719 = ~w21717 & ~w21718;
assign w21720 = ~w21702 & w21719;
assign w21721 = w21702 & ~w21719;
assign w21722 = ~w13714 & w13718;
assign w21723 = ~w13719 & ~w21722;
assign w21724 = (~w21715 & ~w21716) | (~w21715 & w36860) | (~w21716 & w36860);
assign w21725 = ~w21723 & ~w21724;
assign w21726 = w21723 & w21724;
assign w21727 = ~w21725 & ~w21726;
assign w21728 = ~w21721 & w21727;
assign w21729 = (~w21688 & w36861) | (~w21688 & w36862) | (w36861 & w36862);
assign w21730 = ~w13721 & ~w13722;
assign w21731 = ~w21725 & w21730;
assign w21732 = w21725 & ~w21730;
assign w21733 = ~w21731 & ~w21732;
assign w21734 = (w21688 & w36863) | (w21688 & w36864) | (w36863 & w36864);
assign w21735 = (w21688 & w36867) | (w21688 & w36868) | (w36867 & w36868);
assign w21736 = w13667 & ~w21735;
assign w21737 = (~w21735 & w36870) | (~w21735 & w36871) | (w36870 & w36871);
assign w21738 = w13330 & ~w13332;
assign w21739 = ~w13333 & ~w21738;
assign w21740 = (~w21735 & w36874) | (~w21735 & w36875) | (w36874 & w36875);
assign w21741 = (~w21735 & w36878) | (~w21735 & w36879) | (w36878 & w36879);
assign w21742 = (w21735 & w36880) | (w21735 & w36881) | (w36880 & w36881);
assign w21743 = ~w21741 & ~w21742;
assign w21744 = w3 & ~w21743;
assign w21745 = (w21735 & w36882) | (w21735 & w36883) | (w36882 & w36883);
assign w21746 = ~w21740 & ~w21745;
assign w21747 = w10835 & w21746;
assign w21748 = ~w21743 & w21746;
assign w21749 = w21743 & ~w21746;
assign w21750 = ~w21748 & ~w21749;
assign w21751 = (w21735 & w36884) | (w21735 & w36885) | (w36884 & w36885);
assign w21752 = ~w21737 & ~w21751;
assign w21753 = ~w21746 & ~w21752;
assign w21754 = (w21688 & w36886) | (w21688 & w36887) | (w36886 & w36887);
assign w21755 = ~w21736 & ~w21754;
assign w21756 = (~w21688 & w36888) | (~w21688 & w36889) | (w36888 & w36889);
assign w21757 = ~w21734 & ~w21756;
assign w21758 = ~w21755 & w21757;
assign w21759 = (~w21688 & w36890) | (~w21688 & w36891) | (w36890 & w36891);
assign w21760 = ~w21699 & ~w21759;
assign w21761 = (~w21688 & w36892) | (~w21688 & w36893) | (w36892 & w36893);
assign w21762 = ~w21760 & ~w21761;
assign w21763 = ~w14888 & ~w21694;
assign w21764 = (w15848 & ~w21688) | (w15848 & w36894) | (~w21688 & w36894);
assign w21765 = (w21690 & w21764) | (w21690 & w21691) | (w21764 & w21691);
assign w21766 = (~w21764 & w36897) | (~w21764 & w36898) | (w36897 & w36898);
assign w21767 = (~w21764 & w36899) | (~w21764 & w36900) | (w36899 & w36900);
assign w21768 = ~w21694 & ~w21695;
assign w21769 = ~w21696 & ~w21768;
assign w21770 = (w21764 & w36901) | (w21764 & w36902) | (w36901 & w36902);
assign w21771 = ~w21767 & ~w21770;
assign w21772 = ~w21762 & ~w21771;
assign w21773 = (w21764 & w36903) | (w21764 & w36904) | (w36903 & w36904);
assign w21774 = w21770 & ~w21773;
assign w21775 = ~w21772 & ~w21774;
assign w21776 = w14318 & ~w14320;
assign w21777 = ~w14321 & ~w21776;
assign w21778 = ~w21759 & w36905;
assign w21779 = (~w21777 & w21759) | (~w21777 & w36906) | (w21759 & w36906);
assign w21780 = ~w21778 & ~w21779;
assign w21781 = ~w21772 & w36907;
assign w21782 = ~w21760 & w22034;
assign w21783 = ~w21781 & ~w21782;
assign w21784 = ~w21240 & ~w21370;
assign w21785 = ~w20644 & w21370;
assign w21786 = ~w21239 & w21785;
assign w21787 = ~w21784 & ~w21786;
assign w21788 = ~w21473 & ~w21476;
assign w21789 = ~w21478 & w21788;
assign w21790 = w21478 & ~w21788;
assign w21791 = ~w21789 & ~w21790;
assign w21792 = w21787 & ~w21791;
assign w21793 = w21177 & w21184;
assign w21794 = ~w21177 & ~w21184;
assign w21795 = ~w21793 & ~w21794;
assign w21796 = ~w21156 & ~w21795;
assign w21797 = w21156 & w21184;
assign w21798 = ~w21796 & ~w21797;
assign w21799 = ~w21179 & ~w21185;
assign w21800 = w21199 & w21206;
assign w21801 = ~w21799 & w21800;
assign w21802 = w21799 & ~w21800;
assign w21803 = ~w21801 & ~w21802;
assign w21804 = ~w21798 & w21803;
assign w21805 = w21798 & ~w21803;
assign w21806 = ~w21141 & ~w21155;
assign w21807 = ~w21156 & ~w21806;
assign w21808 = w21795 & w21807;
assign w21809 = ~w21113 & ~w21114;
assign w21810 = ~w21133 & ~w21140;
assign w21811 = w21809 & ~w21810;
assign w21812 = ~w21809 & w21810;
assign w21813 = ~w21811 & ~w21812;
assign w21814 = w21097 & ~w21112;
assign w21815 = ~w21113 & ~w21814;
assign w21816 = w21813 & ~w21815;
assign w21817 = ~w21807 & w21816;
assign w21818 = w21813 & ~w21817;
assign w21819 = ~w21808 & ~w21818;
assign w21820 = ~w21795 & w21806;
assign w21821 = ~w21797 & ~w21820;
assign w21822 = ~w21819 & w21821;
assign w21823 = ~w21805 & ~w21822;
assign w21824 = ~w21804 & ~w21823;
assign w21825 = ~w21179 & w31994;
assign w21826 = (~w21199 & w21179) | (~w21199 & w31995) | (w21179 & w31995);
assign w21827 = ~w21825 & ~w21826;
assign w21828 = w21224 & w21827;
assign w21829 = ~w21224 & ~w21827;
assign w21830 = ~w21828 & ~w21829;
assign w21831 = ~w21823 & w31996;
assign w21832 = ~w21201 & w36908;
assign w21833 = ~w21225 & ~w21832;
assign w21834 = ~w21803 & w21833;
assign w21835 = ~w21831 & ~w21834;
assign w21836 = w21230 & w21237;
assign w21837 = ~w21225 & w21836;
assign w21838 = ~w21231 & ~w21237;
assign w21839 = ~w21837 & ~w21838;
assign w21840 = w21206 & ~w21229;
assign w21841 = ~w21226 & w21840;
assign w21842 = ~w21201 & w21841;
assign w21843 = ~w21209 & w21219;
assign w21844 = (~w21218 & ~w20372) | (~w21218 & w36909) | (~w20372 & w36909);
assign w21845 = w21209 & w21844;
assign w21846 = ~w21843 & ~w21845;
assign w21847 = w21236 & w21846;
assign w21848 = ~w21842 & w21847;
assign w21849 = w20636 & ~w21848;
assign w21850 = ~w20620 & ~w20623;
assign w21851 = w20643 & w21850;
assign w21852 = w21849 & ~w21851;
assign w21853 = ~w21849 & w21851;
assign w21854 = ~w21852 & ~w21853;
assign w21855 = w21839 & ~w21854;
assign w21856 = ~w21230 & ~w21237;
assign w21857 = w21833 & w21856;
assign w21858 = (~w21230 & ~w21207) | (~w21230 & w31997) | (~w21207 & w31997);
assign w21859 = ~w21201 & w31998;
assign w21860 = w21237 & ~w21859;
assign w21861 = ~w21858 & w21860;
assign w21862 = ~w21225 & w21237;
assign w21863 = ~w21237 & ~w21859;
assign w21864 = ~w21862 & ~w21863;
assign w21865 = ~w21861 & ~w21864;
assign w21866 = ~w21857 & w21865;
assign w21867 = ~w21855 & w21866;
assign w21868 = ~w21835 & w21867;
assign w21869 = ~w21839 & w21854;
assign w21870 = ~w21836 & ~w21856;
assign w21871 = w21833 & ~w21870;
assign w21872 = (~w21871 & ~w21854) | (~w21871 & w31999) | (~w21854 & w31999);
assign w21873 = ~w21786 & w21854;
assign w21874 = ~w21784 & w21873;
assign w21875 = w21872 & ~w21874;
assign w21876 = ~w21868 & w21875;
assign w21877 = ~w21792 & w21876;
assign w21878 = ~w21787 & ~w21854;
assign w21879 = w21240 & ~w21791;
assign w21880 = ~w21370 & w21788;
assign w21881 = ~w21786 & ~w21880;
assign w21882 = ~w21879 & ~w21881;
assign w21883 = ~w21878 & ~w21882;
assign w21884 = ~w21877 & w21883;
assign w21885 = ~w21559 & ~w21607;
assign w21886 = ~w21480 & w21885;
assign w21887 = (w21643 & ~w21886) | (w21643 & w32000) | (~w21886 & w32000);
assign w21888 = ~w21559 & ~w21642;
assign w21889 = ~w21480 & w21888;
assign w21890 = w21640 & ~w21642;
assign w21891 = (~w21890 & ~w21889) | (~w21890 & w32001) | (~w21889 & w32001);
assign w21892 = ~w21887 & w21891;
assign w21893 = ~w21784 & w21791;
assign w21894 = ~w21882 & ~w21893;
assign w21895 = ~w21892 & w21894;
assign w21896 = ~w21884 & ~w21895;
assign w21897 = ~w21559 & ~w21640;
assign w21898 = ~w21475 & ~w21480;
assign w21899 = ~w21897 & w21898;
assign w21900 = w21897 & ~w21898;
assign w21901 = ~w21899 & ~w21900;
assign w21902 = ~w21892 & ~w21901;
assign w21903 = w21894 & ~w21901;
assign w21904 = (w21892 & ~w21894) | (w21892 & w21914) | (~w21894 & w21914);
assign w21905 = ~w21902 & ~w21904;
assign w21906 = ~w21896 & w21905;
assign w21907 = ~w21635 & ~w21670;
assign w21908 = (w32002 & ~w21886) | (w32002 & w36910) | (~w21886 & w36910);
assign w21909 = (w21886 & w36911) | (w21886 & w36912) | (w36911 & w36912);
assign w21910 = ~w21908 & ~w21909;
assign w21911 = ~w21892 & w21910;
assign w21912 = ~w21896 & w32004;
assign w21913 = w21892 & ~w21910;
assign w21914 = w21892 & w21901;
assign w21915 = ~w21913 & ~w21914;
assign w21916 = ~w21663 & ~w21675;
assign w21917 = ~w21670 & w21916;
assign w21918 = (w21917 & w21643) | (w21917 & w32457) | (w21643 & w32457);
assign w21919 = (w21918 & ~w21638) | (w21918 & w36913) | (~w21638 & w36913);
assign w21920 = (w21638 & w36914) | (w21638 & w36915) | (w36914 & w36915);
assign w21921 = ~w21919 & ~w21920;
assign w21922 = ~w21910 & w21921;
assign w21923 = w21915 & ~w21922;
assign w21924 = ~w21912 & w21923;
assign w21925 = (w17633 & w21674) | (w17633 & w32007) | (w21674 & w32007);
assign w21926 = ~w17090 & ~w17631;
assign w21927 = ~w17090 & ~w17613;
assign w21928 = ~w17611 & w21927;
assign w21929 = w21926 & ~w21928;
assign w21930 = ~w17611 & ~w21678;
assign w21931 = w21677 & w21930;
assign w21932 = w21677 & w36916;
assign w21933 = (~w21929 & w21674) | (~w21929 & w32458) | (w21674 & w32458);
assign w21934 = ~w21925 & w21933;
assign w21935 = w17611 & ~w21927;
assign w21936 = ~w21928 & ~w21935;
assign w21937 = (w21931 & w21639) | (w21931 & w32459) | (w21639 & w32459);
assign w21938 = (~w21639 & w36917) | (~w21639 & w36918) | (w36917 & w36918);
assign w21939 = (w21639 & w36919) | (w21639 & w36920) | (w36919 & w36920);
assign w21940 = ~w21938 & ~w21939;
assign w21941 = w21934 & ~w21940;
assign w21942 = ~w21934 & w21940;
assign w21943 = ~w21941 & ~w21942;
assign w21944 = (~w21639 & w32460) | (~w21639 & w32461) | (w32460 & w32461);
assign w21945 = ~w21937 & ~w21944;
assign w21946 = ~w21936 & w21945;
assign w21947 = w21943 & ~w21946;
assign w21948 = ~w21669 & ~w21675;
assign w21949 = (w21948 & w21639) | (w21948 & w32462) | (w21639 & w32462);
assign w21950 = (~w21676 & w21639) | (~w21676 & w32463) | (w21639 & w32463);
assign w21951 = ~w21949 & w21950;
assign w21952 = w21921 & w21951;
assign w21953 = w21910 & ~w21921;
assign w21954 = ~w21921 & ~w21951;
assign w21955 = ~w21953 & ~w21954;
assign w21956 = w21945 & ~w21951;
assign w21957 = w21955 & w32009;
assign w21958 = w21947 & w21957;
assign w21959 = ~w21924 & w21958;
assign w21960 = ~w21940 & ~w21945;
assign w21961 = ~w21945 & w21951;
assign w21962 = ~w21960 & w32010;
assign w21963 = w21947 & ~w21962;
assign w21964 = w17629 & ~w21684;
assign w21965 = ~w21685 & ~w21964;
assign w21966 = (w21674 & w36921) | (w21674 & w36922) | (w36921 & w36922);
assign w21967 = (~w21674 & w36923) | (~w21674 & w36924) | (w36923 & w36924);
assign w21968 = ~w21966 & ~w21967;
assign w21969 = ~w15835 & ~w21682;
assign w21970 = (w21639 & w36925) | (w21639 & w36926) | (w36925 & w36926);
assign w21971 = w21969 & w21970;
assign w21972 = ~w21969 & ~w21970;
assign w21973 = ~w21971 & ~w21972;
assign w21974 = ~w21968 & ~w21973;
assign w21975 = w21934 & ~w21965;
assign w21976 = ~w21941 & ~w21975;
assign w21977 = ~w21974 & w21976;
assign w21978 = ~w21963 & w21977;
assign w21979 = ~w21959 & w21978;
assign w21980 = w15838 & ~w21688;
assign w21981 = w15835 & ~w15837;
assign w21982 = (w21685 & w36927) | (w21685 & w36928) | (w36927 & w36928);
assign w21983 = (w21639 & w36929) | (w21639 & w36930) | (w36929 & w36930);
assign w21984 = ~w21981 & ~w21983;
assign w21985 = ~w21980 & w21984;
assign w21986 = ~w15566 & ~w15840;
assign w21987 = (w21685 & w36931) | (w21685 & w36932) | (w36931 & w36932);
assign w21988 = (w21639 & w36933) | (w21639 & w36934) | (w36933 & w36934);
assign w21989 = ~w15702 & ~w15838;
assign w21990 = (w21986 & w21988) | (w21986 & w36935) | (w21988 & w36935);
assign w21991 = ~w21988 & w36936;
assign w21992 = ~w21990 & ~w21991;
assign w21993 = w21985 & ~w21992;
assign w21994 = ~w21985 & w21992;
assign w21995 = ~w21993 & ~w21994;
assign w21996 = ~w21973 & w21985;
assign w21997 = w21973 & ~w21985;
assign w21998 = ~w21996 & ~w21997;
assign w21999 = (w21968 & w21973) | (w21968 & w22926) | (w21973 & w22926);
assign w22000 = w21998 & ~w21999;
assign w22001 = w21995 & w22000;
assign w22002 = (w22001 & w21959) | (w22001 & w36937) | (w21959 & w36937);
assign w22003 = w15840 & ~w15846;
assign w22004 = w15703 & ~w15846;
assign w22005 = (w22004 & w21688) | (w22004 & w36938) | (w21688 & w36938);
assign w22006 = (w21688 & w36939) | (w21688 & w36940) | (w36939 & w36940);
assign w22007 = ~w22005 & w22006;
assign w22008 = w21992 & ~w22007;
assign w22009 = ~w21992 & w22007;
assign w22010 = ~w22008 & ~w22009;
assign w22011 = ~w21993 & ~w21996;
assign w22012 = w22010 & w22011;
assign w22013 = ~w21764 & w36941;
assign w22014 = ~w21765 & ~w22013;
assign w22015 = w22007 & w22014;
assign w22016 = ~w22007 & ~w22014;
assign w22017 = ~w22015 & ~w22016;
assign w22018 = ~w22008 & w22017;
assign w22019 = (w22018 & w22002) | (w22018 & w36942) | (w22002 & w36942);
assign w22020 = ~w21766 & ~w21773;
assign w22021 = ~w22014 & w22020;
assign w22022 = (w32014 & w22002) | (w32014 & w36943) | (w22002 & w36943);
assign w22023 = w22014 & ~w22020;
assign w22024 = ~w22015 & ~w22023;
assign w22025 = w21771 & ~w22020;
assign w22026 = w21762 & w21771;
assign w22027 = ~w22025 & ~w22026;
assign w22028 = ~w21782 & w22027;
assign w22029 = ~w21720 & ~w21721;
assign w22030 = (~w21688 & w36946) | (~w21688 & w36947) | (w36946 & w36947);
assign w22031 = (w21688 & w36948) | (w21688 & w36949) | (w36948 & w36949);
assign w22032 = ~w22030 & ~w22031;
assign w22033 = (~w21688 & w36950) | (~w21688 & w36951) | (w36950 & w36951);
assign w22034 = (w21688 & w36952) | (w21688 & w36953) | (w36952 & w36953);
assign w22035 = ~w22033 & ~w22034;
assign w22036 = w22032 & ~w22035;
assign w22037 = ~w21720 & ~w21727;
assign w22038 = (w21688 & w36954) | (w21688 & w36955) | (w36954 & w36955);
assign w22039 = ~w21729 & ~w22038;
assign w22040 = w22032 & w22039;
assign w22041 = ~w22036 & ~w22040;
assign w22042 = (~w22022 & w36956) | (~w22022 & w36957) | (w36956 & w36957);
assign w22043 = ~w22032 & w22035;
assign w22044 = ~w22032 & ~w22039;
assign w22045 = ~w22043 & ~w22044;
assign w22046 = w21757 & ~w22039;
assign w22047 = w21734 & ~w22038;
assign w22048 = ~w22046 & ~w22047;
assign w22049 = w21755 & ~w21757;
assign w22050 = ~w21758 & ~w22049;
assign w22051 = w22048 & w22050;
assign w22052 = w21755 & w22046;
assign w22053 = (~w22042 & w36959) | (~w22042 & w36960) | (w36959 & w36960);
assign w22054 = w21752 & w21755;
assign w22055 = ~w21752 & ~w21755;
assign w22056 = ~w22054 & ~w22055;
assign w22057 = w22053 & w36961;
assign w22058 = w21746 & w21752;
assign w22059 = ~w21753 & ~w22058;
assign w22060 = ~w22054 & w22059;
assign w22061 = (w22060 & ~w22053) | (w22060 & w36962) | (~w22053 & w36962);
assign w22062 = (w22053 & w36963) | (w22053 & w36964) | (w36963 & w36964);
assign w22063 = (w22053 & w36965) | (w22053 & w36966) | (w36965 & w36966);
assign w22064 = (~w22053 & w36967) | (~w22053 & w36968) | (w36967 & w36968);
assign w22065 = ~w22063 & ~w22064;
assign w22066 = ~w21744 & ~w21747;
assign w22067 = (w22066 & ~w22065) | (w22066 & w36969) | (~w22065 & w36969);
assign w22068 = (a_2 & ~w21752) | (a_2 & w34211) | (~w21752 & w34211);
assign w22069 = w22067 & ~w22068;
assign w22070 = (w22065 & w36970) | (w22065 & w36971) | (w36970 & w36971);
assign w22071 = ~w22069 & ~w22070;
assign w22072 = w7511 & ~w21945;
assign w22073 = w7489 & w21951;
assign w22074 = w7192 & w21921;
assign w22075 = ~w21922 & ~w21952;
assign w22076 = w21915 & w22075;
assign w22077 = w21955 & ~w22076;
assign w22078 = ~w21954 & w32015;
assign w22079 = ~w21896 & w36972;
assign w22080 = ~w21956 & ~w21961;
assign w22081 = (w22080 & w22079) | (w22080 & w32464) | (w22079 & w32464);
assign w22082 = ~w22079 & w32465;
assign w22083 = ~w22081 & ~w22082;
assign w22084 = ~w22073 & ~w22074;
assign w22085 = ~w22072 & w22084;
assign w22086 = (w22085 & ~w22083) | (w22085 & w36973) | (~w22083 & w36973);
assign w22087 = a_11 & ~w22086;
assign w22088 = (~w22083 & w36974) | (~w22083 & w36975) | (w36974 & w36975);
assign w22089 = ~w22087 & ~w22088;
assign w22090 = ~w21894 & w21901;
assign w22091 = ~w21903 & ~w22090;
assign w22092 = w21884 & ~w22091;
assign w22093 = ~w21894 & w21914;
assign w22094 = ~w21902 & ~w22093;
assign w22095 = ~w22092 & ~w22094;
assign w22096 = ~w21906 & ~w22095;
assign w22097 = w6998 & w21901;
assign w22098 = w6996 & w21892;
assign w22099 = ~w21882 & w36976;
assign w22100 = ~w22097 & ~w22098;
assign w22101 = ~w22099 & w22100;
assign w22102 = (w22096 & w32466) | (w22096 & w32467) | (w32466 & w32467);
assign w22103 = (~w22096 & w32468) | (~w22096 & w32469) | (w32468 & w32469);
assign w22104 = ~w22102 & ~w22103;
assign w22105 = (w21872 & ~w21867) | (w21872 & w32017) | (~w21867 & w32017);
assign w22106 = ~w21874 & ~w21878;
assign w22107 = w22105 & w22106;
assign w22108 = w6063 & w22107;
assign w22109 = w21873 & w32018;
assign w22110 = w6063 & ~w21854;
assign w22111 = ~w21787 & w22110;
assign w22112 = ~w22109 & ~w22111;
assign w22113 = ~w22105 & ~w22112;
assign w22114 = w6059 & ~w21839;
assign w22115 = w6061 & w21854;
assign w22116 = w6304 & w21787;
assign w22117 = ~w22114 & ~w22115;
assign w22118 = ~w22116 & w22117;
assign w22119 = ~w22113 & w22118;
assign w22120 = ~w22108 & w22119;
assign w22121 = a_17 & ~w22120;
assign w22122 = ~a_17 & w22120;
assign w22123 = ~w22121 & ~w22122;
assign w22124 = ~w21813 & w21815;
assign w22125 = ~w21813 & w32019;
assign w22126 = w5286 & w21813;
assign w22127 = ~w22125 & ~w22126;
assign w22128 = w21813 & w32020;
assign w22129 = w504 & w21815;
assign w22130 = w21815 & w35960;
assign w22131 = w5080 & w21815;
assign w22132 = ~w22130 & ~w22131;
assign w22133 = ~w22128 & w22132;
assign w22134 = w22127 & w22133;
assign w22135 = ~w22127 & w22130;
assign w22136 = ~w22134 & ~w22135;
assign w22137 = ~w21808 & w21821;
assign w22138 = w21818 & ~w22137;
assign w22139 = ~w22137 & w32021;
assign w22140 = ~w21796 & w32022;
assign w22141 = w5308 & w21813;
assign w22142 = w5818 & w21807;
assign w22143 = (w5309 & w21817) | (w5309 & w32023) | (w21817 & w32023);
assign w22144 = w22137 & w22143;
assign w22145 = ~w22141 & ~w22142;
assign w22146 = ~w22140 & w22145;
assign w22147 = ~w22144 & w22146;
assign w22148 = ~w22139 & w22147;
assign w22149 = ~w21813 & w32024;
assign w22150 = w5816 & w21813;
assign w22151 = ~w22149 & ~w22150;
assign w22152 = w21813 & w32025;
assign w22153 = w5300 & w21815;
assign w22154 = w21815 & w36039;
assign w22155 = w5818 & w21815;
assign w22156 = ~w22154 & ~w22155;
assign w22157 = ~w22152 & w22156;
assign w22158 = w22151 & w22157;
assign w22159 = a_20 & ~w22158;
assign w22160 = w21807 & ~w21816;
assign w22161 = ~w21817 & ~w22160;
assign w22162 = w5309 & ~w22161;
assign w22163 = w5308 & w21815;
assign w22164 = w5816 & w21807;
assign w22165 = (~w22163 & ~w21813) | (~w22163 & w36977) | (~w21813 & w36977);
assign w22166 = ~w22164 & w22165;
assign w22167 = ~w22162 & w22166;
assign w22168 = ~w22159 & w22167;
assign w22169 = (w22167 & w32470) | (w22167 & w32471) | (w32470 & w32471);
assign w22170 = ~w22148 & ~w22169;
assign w22171 = w22147 & w32027;
assign w22172 = (~w22129 & ~w22167) | (~w22129 & w32472) | (~w22167 & w32472);
assign w22173 = ~w22171 & ~w22172;
assign w22174 = ~w22170 & w22173;
assign w22175 = ~w22136 & ~w22174;
assign w22176 = w22136 & w22174;
assign w22177 = ~w21804 & ~w21805;
assign w22178 = w21822 & ~w22177;
assign w22179 = (w5309 & ~w21803) | (w5309 & w32029) | (~w21803 & w32029);
assign w22180 = w21823 & w22179;
assign w22181 = ~w21796 & w36978;
assign w22182 = w5308 & w21807;
assign w22183 = w5816 & ~w21803;
assign w22184 = ~w22181 & ~w22182;
assign w22185 = ~w22183 & w22184;
assign w22186 = ~w22180 & w22185;
assign w22187 = (a_20 & ~w22186) | (a_20 & w32030) | (~w22186 & w32030);
assign w22188 = w22186 & w32031;
assign w22189 = ~w22187 & ~w22188;
assign w22190 = ~w22176 & ~w22189;
assign w22191 = ~w22175 & ~w22190;
assign w22192 = a_23 & ~w22134;
assign w22193 = w5017 & ~w22161;
assign w22194 = w5016 & w21815;
assign w22195 = w5286 & w21807;
assign w22196 = (~w22194 & ~w21813) | (~w22194 & w36979) | (~w21813 & w36979);
assign w22197 = ~w22195 & w22196;
assign w22198 = ~w22193 & w22197;
assign w22199 = w22192 & ~w22198;
assign w22200 = ~w22192 & w22198;
assign w22201 = ~w22199 & ~w22200;
assign w22202 = w8311 & w21830;
assign w22203 = w21824 & w22202;
assign w22204 = w8311 & ~w21830;
assign w22205 = ~w21824 & w22204;
assign w22206 = ~w22203 & ~w22205;
assign w22207 = ~w22201 & ~w22206;
assign w22208 = w8339 & w21830;
assign w22209 = w21824 & w22208;
assign w22210 = w8339 & ~w21830;
assign w22211 = ~w21824 & w22210;
assign w22212 = ~w22209 & ~w22211;
assign w22213 = w5816 & ~w21224;
assign w22214 = w21207 & w22213;
assign w22215 = w5818 & ~w21800;
assign w22216 = w21799 & w22215;
assign w22217 = w5818 & w21800;
assign w22218 = ~w21799 & w22217;
assign w22219 = w5816 & w21224;
assign w22220 = ~w21207 & w22219;
assign w22221 = ~w21796 & w32032;
assign w22222 = ~w22216 & ~w22218;
assign w22223 = ~w22214 & w22222;
assign w22224 = ~w22220 & ~w22221;
assign w22225 = w22223 & w22224;
assign w22226 = a_20 & ~w22225;
assign w22227 = ~a_20 & w22225;
assign w22228 = ~w22226 & ~w22227;
assign w22229 = ~w22201 & ~w22228;
assign w22230 = w22212 & w22229;
assign w22231 = ~w22207 & ~w22230;
assign w22232 = w22212 & ~w22228;
assign w22233 = w22201 & w22206;
assign w22234 = ~w22232 & w22233;
assign w22235 = w22231 & ~w22234;
assign w22236 = w22191 & ~w22235;
assign w22237 = ~w22191 & w22235;
assign w22238 = ~w22236 & ~w22237;
assign w22239 = w22123 & ~w22238;
assign w22240 = ~w22123 & w22238;
assign w22241 = ~w22239 & ~w22240;
assign w22242 = ~w21865 & ~w21871;
assign w22243 = ~w21834 & ~w21871;
assign w22244 = ~w21831 & w22243;
assign w22245 = ~w22242 & ~w22244;
assign w22246 = ~w21855 & ~w21869;
assign w22247 = ~w22245 & w22246;
assign w22248 = w6063 & w22247;
assign w22249 = w6063 & ~w22246;
assign w22250 = w6059 & w21833;
assign w22251 = w6304 & w21854;
assign w22252 = (~w22250 & w21839) | (~w22250 & w36980) | (w21839 & w36980);
assign w22253 = ~w22251 & w22252;
assign w22254 = (w22253 & ~w22249) | (w22253 & w32033) | (~w22249 & w32033);
assign w22255 = ~w22248 & w22254;
assign w22256 = ~a_17 & w22255;
assign w22257 = a_17 & ~w22255;
assign w22258 = ~w22256 & ~w22257;
assign w22259 = ~w22175 & ~w22176;
assign w22260 = ~w22189 & w22259;
assign w22261 = w22189 & ~w22259;
assign w22262 = ~w22260 & ~w22261;
assign w22263 = w22258 & ~w22262;
assign w22264 = ~w22258 & w22262;
assign w22265 = (~w22167 & w36981) | (~w22167 & w36982) | (w36981 & w36982);
assign w22266 = ~w22169 & ~w22265;
assign w22267 = w22148 & w22266;
assign w22268 = ~w22148 & ~w22266;
assign w22269 = ~w22267 & ~w22268;
assign w22270 = w6304 & ~w21839;
assign w22271 = w6061 & w21833;
assign w22272 = w6059 & ~w21803;
assign w22273 = ~w22271 & ~w22272;
assign w22274 = (a_17 & w22270) | (a_17 & w36983) | (w22270 & w36983);
assign w22275 = ~w22270 & w36984;
assign w22276 = w21835 & ~w21866;
assign w22277 = ~w21835 & w21866;
assign w22278 = ~w22276 & ~w22277;
assign w22279 = ~w22274 & ~w22275;
assign w22280 = ~w22278 & w22279;
assign w22281 = ~w22270 & w36985;
assign w22282 = ~w22274 & ~w22281;
assign w22283 = w22278 & w22282;
assign w22284 = ~w22280 & ~w22283;
assign w22285 = w22269 & ~w22284;
assign w22286 = ~w22269 & w22284;
assign w22287 = w22159 & ~w22167;
assign w22288 = ~w22168 & ~w22287;
assign w22289 = (~w21830 & w21823) | (~w21830 & w32034) | (w21823 & w32034);
assign w22290 = w8391 & w22289;
assign w22291 = w8391 & w21830;
assign w22292 = w21824 & w22291;
assign w22293 = w6304 & ~w21224;
assign w22294 = w21207 & w22293;
assign w22295 = w6304 & w21224;
assign w22296 = ~w21207 & w22295;
assign w22297 = ~w22294 & ~w22296;
assign w22298 = (w6059 & ~w21156) | (w6059 & w32035) | (~w21156 & w32035);
assign w22299 = ~w21796 & w22298;
assign w22300 = w6061 & ~w21800;
assign w22301 = w21799 & w22300;
assign w22302 = w6061 & w21800;
assign w22303 = ~w21799 & w22302;
assign w22304 = ~w22301 & ~w22303;
assign w22305 = ~w22299 & w22304;
assign w22306 = w22297 & w22305;
assign w22307 = w17694 & w22306;
assign w22308 = a_17 & ~w22306;
assign w22309 = ~w22307 & ~w22308;
assign w22310 = ~w22292 & w22309;
assign w22311 = ~w22290 & w22310;
assign w22312 = (~a_17 & w21796) | (~a_17 & w32036) | (w21796 & w32036);
assign w22313 = w22304 & w22312;
assign w22314 = w22297 & w22313;
assign w22315 = ~w21830 & w22314;
assign w22316 = w21824 & w22315;
assign w22317 = w21830 & w22314;
assign w22318 = ~w21824 & w22317;
assign w22319 = ~w22316 & ~w22318;
assign w22320 = (~w22288 & ~w22311) | (~w22288 & w32473) | (~w22311 & w32473);
assign w22321 = ~w22137 & w32037;
assign w22322 = ~w21796 & w32038;
assign w22323 = w6059 & w21813;
assign w22324 = w6061 & w21807;
assign w22325 = (w6063 & w21817) | (w6063 & w32039) | (w21817 & w32039);
assign w22326 = w22137 & w22325;
assign w22327 = ~w22323 & ~w22324;
assign w22328 = ~w22322 & w22327;
assign w22329 = ~w22326 & w22328;
assign w22330 = ~w22321 & w22329;
assign w22331 = ~w21816 & ~w22124;
assign w22332 = w6063 & ~w22331;
assign w22333 = w6054 & w21815;
assign w22334 = w21815 & w36074;
assign w22335 = w6061 & w21815;
assign w22336 = (~w22335 & ~w21813) | (~w22335 & w32040) | (~w21813 & w32040);
assign w22337 = (~w21813 & w36986) | (~w21813 & w36987) | (w36986 & w36987);
assign w22338 = (w22337 & w22331) | (w22337 & w36988) | (w22331 & w36988);
assign w22339 = (a_17 & w22332) | (a_17 & w32041) | (w22332 & w32041);
assign w22340 = w6063 & ~w22161;
assign w22341 = w6059 & w21815;
assign w22342 = w6304 & w21807;
assign w22343 = (~w22341 & ~w21813) | (~w22341 & w36989) | (~w21813 & w36989);
assign w22344 = ~w22342 & w22343;
assign w22345 = ~w22340 & w22344;
assign w22346 = ~w22339 & w22345;
assign w22347 = (w22345 & w32474) | (w22345 & w32475) | (w32474 & w32475);
assign w22348 = ~w22330 & ~w22347;
assign w22349 = w22329 & w32043;
assign w22350 = (~w22153 & ~w22345) | (~w22153 & w36990) | (~w22345 & w36990);
assign w22351 = ~w22349 & ~w22350;
assign w22352 = ~w22348 & w22351;
assign w22353 = ~w22151 & w22154;
assign w22354 = ~w22158 & ~w22353;
assign w22355 = ~w22352 & ~w22354;
assign w22356 = ~w22177 & w32044;
assign w22357 = (w6063 & w21819) | (w6063 & w32045) | (w21819 & w32045);
assign w22358 = w22177 & w22357;
assign w22359 = ~w21796 & w36991;
assign w22360 = w6304 & ~w21803;
assign w22361 = w6059 & w21807;
assign w22362 = ~w22359 & ~w22361;
assign w22363 = ~w22360 & w22362;
assign w22364 = ~w22358 & w22363;
assign w22365 = (a_17 & ~w22364) | (a_17 & w32046) | (~w22364 & w32046);
assign w22366 = w22364 & w32047;
assign w22367 = ~w22365 & ~w22366;
assign w22368 = ~w22355 & w22367;
assign w22369 = w22352 & w22354;
assign w22370 = w22288 & w22319;
assign w22371 = w22311 & w22370;
assign w22372 = ~w22369 & ~w22371;
assign w22373 = (~w22320 & ~w22372) | (~w22320 & w32476) | (~w22372 & w32476);
assign w22374 = (~w22285 & ~w22373) | (~w22285 & w32048) | (~w22373 & w32048);
assign w22375 = ~w22264 & ~w22374;
assign w22376 = ~w22263 & ~w22375;
assign w22377 = w22241 & ~w22376;
assign w22378 = ~w22241 & w22376;
assign w22379 = ~w22377 & ~w22378;
assign w22380 = w22104 & w22379;
assign w22381 = ~w21876 & ~w21878;
assign w22382 = ~w21792 & ~w21882;
assign w22383 = w22381 & ~w22382;
assign w22384 = ~w21882 & w32050;
assign w22385 = ~w22381 & w22384;
assign w22386 = ~w21882 & w32051;
assign w22387 = w6446 & w21854;
assign w22388 = w6998 & w21787;
assign w22389 = ~w22387 & ~w22388;
assign w22390 = ~w22386 & w22389;
assign w22391 = ~w22385 & w22390;
assign w22392 = (a_14 & ~w22391) | (a_14 & w32052) | (~w22391 & w32052);
assign w22393 = w22391 & w32053;
assign w22394 = ~w22392 & ~w22393;
assign w22395 = ~w22285 & ~w22286;
assign w22396 = w22373 & w22395;
assign w22397 = ~w22373 & ~w22395;
assign w22398 = ~w22396 & ~w22397;
assign w22399 = ~w22394 & ~w22398;
assign w22400 = w6447 & w22107;
assign w22401 = w21873 & w32054;
assign w22402 = w6447 & ~w21854;
assign w22403 = ~w21787 & w22402;
assign w22404 = ~w22401 & ~w22403;
assign w22405 = ~w22105 & ~w22404;
assign w22406 = w6446 & ~w21839;
assign w22407 = w6998 & w21854;
assign w22408 = w6996 & w21787;
assign w22409 = ~w22406 & ~w22407;
assign w22410 = ~w22408 & w22409;
assign w22411 = ~w22405 & w22410;
assign w22412 = ~w22400 & w22411;
assign w22413 = a_14 & ~w22412;
assign w22414 = ~a_14 & w22412;
assign w22415 = ~w22413 & ~w22414;
assign w22416 = ~w22368 & ~w22369;
assign w22417 = ~w22320 & ~w22371;
assign w22418 = w22416 & ~w22417;
assign w22419 = ~w22416 & w22417;
assign w22420 = ~w22418 & ~w22419;
assign w22421 = ~w22415 & ~w22420;
assign w22422 = w6447 & w22247;
assign w22423 = w6447 & ~w22246;
assign w22424 = w6446 & w21833;
assign w22425 = w6996 & w21854;
assign w22426 = (~w22424 & w21839) | (~w22424 & w36992) | (w21839 & w36992);
assign w22427 = ~w22425 & w22426;
assign w22428 = (w22427 & ~w22423) | (w22427 & w32055) | (~w22423 & w32055);
assign w22429 = ~w22422 & w22428;
assign w22430 = a_14 & ~w22429;
assign w22431 = ~a_14 & w22429;
assign w22432 = ~w22430 & ~w22431;
assign w22433 = ~w22355 & ~w22369;
assign w22434 = w22367 & w22433;
assign w22435 = ~w22367 & ~w22433;
assign w22436 = ~w22434 & ~w22435;
assign w22437 = ~w22432 & ~w22436;
assign w22438 = w22432 & w22436;
assign w22439 = (~w22345 & w32477) | (~w22345 & w32478) | (w32477 & w32478);
assign w22440 = ~w22347 & ~w22439;
assign w22441 = w22330 & w22440;
assign w22442 = ~w22330 & ~w22440;
assign w22443 = ~w22441 & ~w22442;
assign w22444 = w22278 & w32479;
assign w22445 = w8592 & w22278;
assign w22446 = w6996 & ~w21839;
assign w22447 = w6998 & w21833;
assign w22448 = w6446 & ~w21803;
assign w22449 = ~w22447 & ~w22448;
assign w22450 = ~w22446 & w36993;
assign w22451 = (a_14 & w22446) | (a_14 & w36994) | (w22446 & w36994);
assign w22452 = ~w22450 & ~w22451;
assign w22453 = ~w22443 & ~w22452;
assign w22454 = ~w22445 & w22453;
assign w22455 = ~w22444 & ~w22454;
assign w22456 = ~w22137 & w32056;
assign w22457 = ~w21796 & w32057;
assign w22458 = w6446 & w21813;
assign w22459 = w6998 & w21807;
assign w22460 = (w6447 & w21817) | (w6447 & w32058) | (w21817 & w32058);
assign w22461 = w22137 & w22460;
assign w22462 = ~w22458 & ~w22459;
assign w22463 = ~w22457 & w22462;
assign w22464 = ~w22461 & w22463;
assign w22465 = ~w22456 & w22464;
assign w22466 = w6447 & ~w22331;
assign w22467 = w6441 & w21815;
assign w22468 = w21815 & w36136;
assign w22469 = w6998 & w21815;
assign w22470 = (~w22469 & ~w21813) | (~w22469 & w32059) | (~w21813 & w32059);
assign w22471 = (~w21813 & w36995) | (~w21813 & w36996) | (w36995 & w36996);
assign w22472 = (w22471 & w22331) | (w22471 & w36997) | (w22331 & w36997);
assign w22473 = (a_14 & w22466) | (a_14 & w32060) | (w22466 & w32060);
assign w22474 = w6447 & ~w22161;
assign w22475 = w6446 & w21815;
assign w22476 = w6996 & w21807;
assign w22477 = (~w22475 & ~w21813) | (~w22475 & w36998) | (~w21813 & w36998);
assign w22478 = ~w22476 & w22477;
assign w22479 = ~w22474 & w22478;
assign w22480 = ~w22473 & w22479;
assign w22481 = (w22479 & w32480) | (w22479 & w32481) | (w32480 & w32481);
assign w22482 = ~w22465 & ~w22481;
assign w22483 = w22464 & w32062;
assign w22484 = (~w22333 & ~w22479) | (~w22333 & w32482) | (~w22479 & w32482);
assign w22485 = ~w22483 & ~w22484;
assign w22486 = ~w22482 & w22485;
assign w22487 = (w22336 & w22331) | (w22336 & w36999) | (w22331 & w36999);
assign w22488 = w22334 & ~w22487;
assign w22489 = ~w22338 & ~w22488;
assign w22490 = w22486 & w22489;
assign w22491 = (w6447 & w21819) | (w6447 & w32064) | (w21819 & w32064);
assign w22492 = w22177 & w22491;
assign w22493 = ~w21796 & w37000;
assign w22494 = w6996 & ~w21803;
assign w22495 = w6446 & w21807;
assign w22496 = ~w22493 & ~w22495;
assign w22497 = ~w22494 & w22496;
assign w22498 = ~w22492 & w22497;
assign w22499 = (a_14 & ~w22498) | (a_14 & w32065) | (~w22498 & w32065);
assign w22500 = w22498 & w32066;
assign w22501 = ~w22499 & ~w22500;
assign w22502 = ~w22490 & ~w22501;
assign w22503 = w22339 & ~w22345;
assign w22504 = ~w22346 & ~w22503;
assign w22505 = w8564 & w21830;
assign w22506 = w21824 & w22505;
assign w22507 = w8564 & ~w21830;
assign w22508 = ~w21824 & w22507;
assign w22509 = ~w22506 & ~w22508;
assign w22510 = ~w22504 & ~w22509;
assign w22511 = w8592 & w21830;
assign w22512 = w21824 & w22511;
assign w22513 = w8592 & ~w21830;
assign w22514 = ~w21824 & w22513;
assign w22515 = ~w22512 & ~w22514;
assign w22516 = w6996 & ~w21224;
assign w22517 = w21207 & w22516;
assign w22518 = w6998 & ~w21800;
assign w22519 = w21799 & w22518;
assign w22520 = w6998 & w21800;
assign w22521 = ~w21799 & w22520;
assign w22522 = w6996 & w21224;
assign w22523 = ~w21207 & w22522;
assign w22524 = ~w21796 & w32067;
assign w22525 = ~w22519 & ~w22521;
assign w22526 = ~w22517 & w22525;
assign w22527 = ~w22523 & ~w22524;
assign w22528 = w22526 & w22527;
assign w22529 = a_14 & ~w22528;
assign w22530 = ~a_14 & w22528;
assign w22531 = ~w22529 & ~w22530;
assign w22532 = ~w22504 & ~w22531;
assign w22533 = w22515 & w22532;
assign w22534 = ~w22510 & ~w22533;
assign w22535 = ~w22486 & ~w22489;
assign w22536 = w22534 & ~w22535;
assign w22537 = w22515 & ~w22531;
assign w22538 = w22504 & w22509;
assign w22539 = ~w22537 & w22538;
assign w22540 = (~w22539 & ~w22536) | (~w22539 & w32068) | (~w22536 & w32068);
assign w22541 = (~w22452 & ~w22278) | (~w22452 & w37001) | (~w22278 & w37001);
assign w22542 = (w22443 & ~w22278) | (w22443 & w32483) | (~w22278 & w32483);
assign w22543 = ~w22541 & w22542;
assign w22544 = w22540 & ~w22543;
assign w22545 = w22455 & ~w22544;
assign w22546 = ~w22438 & ~w22545;
assign w22547 = ~w22437 & ~w22546;
assign w22548 = ~w22421 & w22547;
assign w22549 = w22415 & w22420;
assign w22550 = w22394 & w22398;
assign w22551 = ~w22549 & ~w22550;
assign w22552 = ~w22548 & w22551;
assign w22553 = ~w22399 & ~w22552;
assign w22554 = ~w21884 & w22091;
assign w22555 = ~w22092 & ~w22554;
assign w22556 = w8564 & w22555;
assign w22557 = w6446 & w21787;
assign w22558 = ~w21882 & w37002;
assign w22559 = (~w22557 & ~w21901) | (~w22557 & w37003) | (~w21901 & w37003);
assign w22560 = ~w22558 & w22559;
assign w22561 = a_14 & w22560;
assign w22562 = ~a_14 & ~w22560;
assign w22563 = ~w22561 & ~w22562;
assign w22564 = (w22563 & ~w22555) | (w22563 & w37004) | (~w22555 & w37004);
assign w22565 = ~w22556 & ~w22564;
assign w22566 = ~w22263 & ~w22264;
assign w22567 = ~w22374 & w22566;
assign w22568 = w22374 & ~w22566;
assign w22569 = ~w22567 & ~w22568;
assign w22570 = w22565 & w22569;
assign w22571 = ~w22553 & ~w22570;
assign w22572 = ~w22565 & ~w22569;
assign w22573 = ~w22104 & ~w22379;
assign w22574 = ~w22572 & ~w22573;
assign w22575 = ~w22571 & w22574;
assign w22576 = ~w22380 & ~w22575;
assign w22577 = ~w21911 & ~w21913;
assign w22578 = (w21896 & w32484) | (w21896 & w32485) | (w32484 & w32485);
assign w22579 = (~w21896 & w32486) | (~w21896 & w32487) | (w32486 & w32487);
assign w22580 = ~w22578 & ~w22579;
assign w22581 = w8564 & ~w22580;
assign w22582 = w6998 & w21892;
assign w22583 = w6446 & w21901;
assign w22584 = w6996 & ~w21910;
assign w22585 = ~w22582 & ~w22583;
assign w22586 = w22585 & w37005;
assign w22587 = (~a_14 & ~w22585) | (~a_14 & w37006) | (~w22585 & w37006);
assign w22588 = ~w22586 & ~w22587;
assign w22589 = (w22588 & w22580) | (w22588 & w37007) | (w22580 & w37007);
assign w22590 = ~w22581 & ~w22589;
assign w22591 = ~w21882 & w32071;
assign w22592 = ~w22381 & w22591;
assign w22593 = ~w21882 & w32072;
assign w22594 = w6059 & w21854;
assign w22595 = w6061 & w21787;
assign w22596 = ~w22594 & ~w22595;
assign w22597 = ~w22593 & w22596;
assign w22598 = ~w22592 & w22597;
assign w22599 = (a_17 & ~w22598) | (a_17 & w32073) | (~w22598 & w32073);
assign w22600 = w22598 & w32074;
assign w22601 = ~w22599 & ~w22600;
assign w22602 = ~w22175 & w22231;
assign w22603 = (~w22234 & ~w22602) | (~w22234 & w32075) | (~w22602 & w32075);
assign w22604 = ~w22137 & w37008;
assign w22605 = ~w21796 & w32076;
assign w22606 = w5080 & w21807;
assign w22607 = w5016 & w21813;
assign w22608 = (w5017 & w21817) | (w5017 & w32077) | (w21817 & w32077);
assign w22609 = w22137 & w22608;
assign w22610 = ~w22606 & ~w22607;
assign w22611 = ~w22605 & w22610;
assign w22612 = ~w22609 & w22611;
assign w22613 = ~w22604 & w22612;
assign w22614 = ~w1222 & w21815;
assign w22615 = (a_23 & ~w22198) | (a_23 & w32078) | (~w22198 & w32078);
assign w22616 = w22614 & ~w22615;
assign w22617 = ~w22614 & w22615;
assign w22618 = ~w22616 & ~w22617;
assign w22619 = w22613 & w22618;
assign w22620 = ~w22613 & ~w22618;
assign w22621 = ~w22619 & ~w22620;
assign w22622 = w5816 & ~w21839;
assign w22623 = w5818 & w21833;
assign w22624 = w5308 & ~w21803;
assign w22625 = ~w22623 & ~w22624;
assign w22626 = (a_20 & w22622) | (a_20 & w37009) | (w22622 & w37009);
assign w22627 = ~w22622 & w37010;
assign w22628 = ~w22626 & ~w22627;
assign w22629 = ~w22278 & w22628;
assign w22630 = ~w22622 & w37011;
assign w22631 = ~w22626 & ~w22630;
assign w22632 = w22278 & w22631;
assign w22633 = ~w22629 & ~w22632;
assign w22634 = w22621 & ~w22633;
assign w22635 = ~w22621 & w22633;
assign w22636 = ~w22634 & ~w22635;
assign w22637 = w22603 & w22636;
assign w22638 = ~w22603 & ~w22636;
assign w22639 = ~w22637 & ~w22638;
assign w22640 = ~w22601 & w22639;
assign w22641 = w22601 & ~w22639;
assign w22642 = ~w22640 & ~w22641;
assign w22643 = ~w22240 & ~w22376;
assign w22644 = (~w22239 & w22376) | (~w22239 & w32488) | (w22376 & w32488);
assign w22645 = w22642 & w22644;
assign w22646 = ~w22642 & ~w22644;
assign w22647 = ~w22645 & ~w22646;
assign w22648 = ~w22590 & w22647;
assign w22649 = w22590 & ~w22647;
assign w22650 = ~w22648 & ~w22649;
assign w22651 = w22576 & ~w22650;
assign w22652 = ~w22576 & w22650;
assign w22653 = ~w22651 & ~w22652;
assign w22654 = w22089 & w22653;
assign w22655 = w7511 & w21921;
assign w22656 = w7192 & w21892;
assign w22657 = w7489 & ~w21910;
assign w22658 = ~w21922 & ~w21953;
assign w22659 = w21915 & ~w22658;
assign w22660 = ~w21912 & w22659;
assign w22661 = ~w21915 & w22658;
assign w22662 = ~w21911 & w22658;
assign w22663 = (~w22661 & ~w21906) | (~w22661 & w32079) | (~w21906 & w32079);
assign w22664 = ~w22660 & w22663;
assign w22665 = ~w22655 & ~w22656;
assign w22666 = ~w22657 & w22665;
assign w22667 = (w22666 & ~w22664) | (w22666 & w37012) | (~w22664 & w37012);
assign w22668 = a_11 & w22667;
assign w22669 = (w22664 & w37013) | (w22664 & w37014) | (w37013 & w37014);
assign w22670 = ~w22668 & ~w22669;
assign w22671 = ~w22570 & ~w22572;
assign w22672 = w22553 & ~w22671;
assign w22673 = ~w22553 & w22671;
assign w22674 = ~w22672 & ~w22673;
assign w22675 = ~w22670 & ~w22674;
assign w22676 = w7489 & w21901;
assign w22677 = ~w21882 & w37015;
assign w22678 = w7511 & w21892;
assign w22679 = ~w22676 & ~w22677;
assign w22680 = ~w22678 & w22679;
assign w22681 = (w22096 & w32489) | (w22096 & w32490) | (w32489 & w32490);
assign w22682 = (~w22096 & w32491) | (~w22096 & w32492) | (w32491 & w32492);
assign w22683 = ~w22681 & ~w22682;
assign w22684 = ~w22421 & ~w22549;
assign w22685 = w22547 & ~w22684;
assign w22686 = ~w22547 & w22684;
assign w22687 = ~w22685 & ~w22686;
assign w22688 = w22683 & ~w22687;
assign w22689 = w9061 & w22555;
assign w22690 = w7192 & w21787;
assign w22691 = ~w21882 & w37016;
assign w22692 = (~w22690 & ~w21901) | (~w22690 & w37017) | (~w21901 & w37017);
assign w22693 = ~w22691 & w22692;
assign w22694 = a_11 & w22693;
assign w22695 = ~a_11 & ~w22693;
assign w22696 = ~w22694 & ~w22695;
assign w22697 = (w22696 & ~w22555) | (w22696 & w37018) | (~w22555 & w37018);
assign w22698 = ~w22689 & ~w22697;
assign w22699 = ~w22437 & ~w22438;
assign w22700 = w22545 & w22699;
assign w22701 = ~w22545 & ~w22699;
assign w22702 = ~w22700 & ~w22701;
assign w22703 = w22698 & w22702;
assign w22704 = ~w21882 & w32082;
assign w22705 = ~w22381 & w22704;
assign w22706 = ~w21882 & w32083;
assign w22707 = w7192 & w21854;
assign w22708 = w7489 & w21787;
assign w22709 = ~w22707 & ~w22708;
assign w22710 = ~w22706 & w22709;
assign w22711 = ~w22705 & w22710;
assign w22712 = w22711 & w32084;
assign w22713 = (a_11 & ~w22711) | (a_11 & w32085) | (~w22711 & w32085);
assign w22714 = ~w22712 & ~w22713;
assign w22715 = w22455 & ~w22543;
assign w22716 = w22540 & ~w22715;
assign w22717 = ~w22540 & w22715;
assign w22718 = ~w22716 & ~w22717;
assign w22719 = ~w22714 & ~w22718;
assign w22720 = ~w22502 & ~w22535;
assign w22721 = w22534 & ~w22539;
assign w22722 = w22720 & ~w22721;
assign w22723 = ~w22720 & w22721;
assign w22724 = ~w22722 & ~w22723;
assign w22725 = ~w22105 & ~w22106;
assign w22726 = ~w22107 & ~w22725;
assign w22727 = w9061 & ~w22726;
assign w22728 = w9089 & ~w22726;
assign w22729 = w7192 & ~w21839;
assign w22730 = w7489 & w21854;
assign w22731 = w7511 & w21787;
assign w22732 = ~w22729 & ~w22730;
assign w22733 = ~w22731 & w22732;
assign w22734 = ~a_11 & ~w22733;
assign w22735 = a_11 & w22733;
assign w22736 = ~w22734 & ~w22735;
assign w22737 = ~w22728 & w22736;
assign w22738 = ~w22727 & ~w22737;
assign w22739 = ~w22724 & w22738;
assign w22740 = w22724 & ~w22738;
assign w22741 = ~w22739 & ~w22740;
assign w22742 = w7193 & w22247;
assign w22743 = w7193 & ~w22246;
assign w22744 = w7192 & w21833;
assign w22745 = w7511 & w21854;
assign w22746 = (~w22744 & w21839) | (~w22744 & w37019) | (w21839 & w37019);
assign w22747 = ~w22745 & w22746;
assign w22748 = (w22747 & ~w22743) | (w22747 & w32086) | (~w22743 & w32086);
assign w22749 = ~w22742 & w22748;
assign w22750 = ~a_11 & w22749;
assign w22751 = a_11 & ~w22749;
assign w22752 = ~w22750 & ~w22751;
assign w22753 = ~w22490 & ~w22535;
assign w22754 = w22501 & ~w22753;
assign w22755 = ~w22501 & w22753;
assign w22756 = ~w22754 & ~w22755;
assign w22757 = w22752 & ~w22756;
assign w22758 = ~w22752 & w22756;
assign w22759 = w7489 & w21833;
assign w22760 = w7192 & ~w21803;
assign w22761 = w7511 & ~w21839;
assign w22762 = ~w22759 & ~w22760;
assign w22763 = ~w22761 & w37020;
assign w22764 = (a_11 & w22761) | (a_11 & w37021) | (w22761 & w37021);
assign w22765 = ~w22763 & ~w22764;
assign w22766 = (~w22765 & ~w22278) | (~w22765 & w37022) | (~w22278 & w37022);
assign w22767 = w9061 & w22278;
assign w22768 = (~w22479 & w37023) | (~w22479 & w37024) | (w37023 & w37024);
assign w22769 = ~w22481 & ~w22768;
assign w22770 = w22465 & w22769;
assign w22771 = ~w22465 & ~w22769;
assign w22772 = ~w22770 & ~w22771;
assign w22773 = (w22772 & ~w22278) | (w22772 & w37025) | (~w22278 & w37025);
assign w22774 = ~w22766 & w22773;
assign w22775 = ~w22137 & w32087;
assign w22776 = ~w21796 & w32088;
assign w22777 = w7192 & w21813;
assign w22778 = w7489 & w21807;
assign w22779 = (w7193 & w21817) | (w7193 & w32089) | (w21817 & w32089);
assign w22780 = w22137 & w22779;
assign w22781 = ~w22777 & ~w22778;
assign w22782 = ~w22776 & w22781;
assign w22783 = ~w22780 & w22782;
assign w22784 = ~w22775 & w22783;
assign w22785 = w7193 & ~w22331;
assign w22786 = w7187 & w21815;
assign w22787 = w21815 & w36236;
assign w22788 = w7489 & w21815;
assign w22789 = (~w22788 & ~w21813) | (~w22788 & w32090) | (~w21813 & w32090);
assign w22790 = (~w21813 & w37026) | (~w21813 & w37027) | (w37026 & w37027);
assign w22791 = (w22790 & w22331) | (w22790 & w37028) | (w22331 & w37028);
assign w22792 = (a_11 & w22785) | (a_11 & w32091) | (w22785 & w32091);
assign w22793 = w7193 & ~w22161;
assign w22794 = w7192 & w21815;
assign w22795 = w7511 & w21807;
assign w22796 = (~w22794 & ~w21813) | (~w22794 & w37029) | (~w21813 & w37029);
assign w22797 = ~w22795 & w22796;
assign w22798 = ~w22793 & w22797;
assign w22799 = ~w22792 & w22798;
assign w22800 = (w22798 & w32493) | (w22798 & w32494) | (w32493 & w32494);
assign w22801 = ~w22784 & ~w22800;
assign w22802 = w22783 & w32093;
assign w22803 = (~w22467 & ~w22798) | (~w22467 & w32495) | (~w22798 & w32495);
assign w22804 = ~w22802 & ~w22803;
assign w22805 = ~w22801 & w22804;
assign w22806 = (w22470 & w22331) | (w22470 & w37030) | (w22331 & w37030);
assign w22807 = w22468 & ~w22806;
assign w22808 = ~w22472 & ~w22807;
assign w22809 = w22805 & w22808;
assign w22810 = (w7193 & w21819) | (w7193 & w32095) | (w21819 & w32095);
assign w22811 = w22177 & w22810;
assign w22812 = ~w21796 & w37031;
assign w22813 = w7511 & ~w21803;
assign w22814 = w7192 & w21807;
assign w22815 = ~w22812 & ~w22814;
assign w22816 = ~w22813 & w22815;
assign w22817 = ~w22811 & w22816;
assign w22818 = (a_11 & ~w22817) | (a_11 & w32096) | (~w22817 & w32096);
assign w22819 = w22817 & w32097;
assign w22820 = ~w22818 & ~w22819;
assign w22821 = ~w22809 & ~w22820;
assign w22822 = w22473 & ~w22479;
assign w22823 = ~w22480 & ~w22822;
assign w22824 = w9061 & w21830;
assign w22825 = w21824 & w22824;
assign w22826 = w9061 & ~w21830;
assign w22827 = ~w21824 & w22826;
assign w22828 = ~w22825 & ~w22827;
assign w22829 = ~w22823 & ~w22828;
assign w22830 = w9089 & w21830;
assign w22831 = w21824 & w22830;
assign w22832 = w9089 & ~w21830;
assign w22833 = ~w21824 & w22832;
assign w22834 = ~w22831 & ~w22833;
assign w22835 = w7511 & ~w21224;
assign w22836 = w21207 & w22835;
assign w22837 = w7489 & ~w21800;
assign w22838 = w21799 & w22837;
assign w22839 = w7489 & w21800;
assign w22840 = ~w21799 & w22839;
assign w22841 = w7511 & w21224;
assign w22842 = ~w21207 & w22841;
assign w22843 = ~w21796 & w32098;
assign w22844 = ~w22838 & ~w22840;
assign w22845 = ~w22836 & w22844;
assign w22846 = ~w22842 & ~w22843;
assign w22847 = w22845 & w22846;
assign w22848 = a_11 & ~w22847;
assign w22849 = ~a_11 & w22847;
assign w22850 = ~w22848 & ~w22849;
assign w22851 = ~w22823 & ~w22850;
assign w22852 = w22834 & w22851;
assign w22853 = ~w22829 & ~w22852;
assign w22854 = ~w22805 & ~w22808;
assign w22855 = w22853 & ~w22854;
assign w22856 = w22834 & ~w22850;
assign w22857 = w22823 & w22828;
assign w22858 = ~w22856 & w22857;
assign w22859 = (~w22858 & ~w22855) | (~w22858 & w32099) | (~w22855 & w32099);
assign w22860 = ~w22774 & w22859;
assign w22861 = (~w22772 & w22766) | (~w22772 & w32496) | (w22766 & w32496);
assign w22862 = ~w22860 & ~w22861;
assign w22863 = ~w22758 & w22862;
assign w22864 = ~w22757 & ~w22863;
assign w22865 = w22741 & ~w22864;
assign w22866 = w22714 & w22718;
assign w22867 = ~w22739 & ~w22866;
assign w22868 = ~w22865 & w22867;
assign w22869 = ~w22719 & ~w22868;
assign w22870 = ~w22703 & ~w22869;
assign w22871 = ~w22698 & ~w22702;
assign w22872 = ~w22683 & w22687;
assign w22873 = ~w22871 & ~w22872;
assign w22874 = ~w22870 & w22873;
assign w22875 = ~w22688 & ~w22874;
assign w22876 = w9061 & ~w22580;
assign w22877 = w7489 & w21892;
assign w22878 = w7192 & w21901;
assign w22879 = w7511 & ~w21910;
assign w22880 = ~w22877 & ~w22878;
assign w22881 = (~a_11 & ~w22880) | (~a_11 & w37032) | (~w22880 & w37032);
assign w22882 = w22880 & w37033;
assign w22883 = ~w22881 & ~w22882;
assign w22884 = (w22883 & w22580) | (w22883 & w37034) | (w22580 & w37034);
assign w22885 = ~w22876 & ~w22884;
assign w22886 = ~w22399 & ~w22550;
assign w22887 = (~w22549 & ~w22547) | (~w22549 & w32497) | (~w22547 & w32497);
assign w22888 = w22886 & w22887;
assign w22889 = ~w22886 & ~w22887;
assign w22890 = ~w22888 & ~w22889;
assign w22891 = w22885 & ~w22890;
assign w22892 = ~w22874 & w32498;
assign w22893 = ~w22885 & w22890;
assign w22894 = w22670 & w22674;
assign w22895 = (~w22893 & ~w22674) | (~w22893 & w32499) | (~w22674 & w32499);
assign w22896 = ~w22892 & w22895;
assign w22897 = ~w22675 & ~w22896;
assign w22898 = w7511 & w21951;
assign w22899 = w7489 & w21921;
assign w22900 = w7192 & ~w21910;
assign w22901 = (~w21952 & w22079) | (~w21952 & w32500) | (w22079 & w32500);
assign w22902 = w21951 & w37035;
assign w22903 = ~w21954 & ~w22902;
assign w22904 = (~w21906 & w37036) | (~w21906 & w37037) | (w37036 & w37037);
assign w22905 = ~w22901 & ~w22904;
assign w22906 = ~w22901 & w37038;
assign w22907 = ~w22898 & w37039;
assign w22908 = ~w22906 & w37040;
assign w22909 = (~a_11 & w22906) | (~a_11 & w37041) | (w22906 & w37041);
assign w22910 = ~w22908 & ~w22909;
assign w22911 = (~w22572 & w22553) | (~w22572 & w32501) | (w22553 & w32501);
assign w22912 = ~w22380 & ~w22573;
assign w22913 = w22911 & ~w22912;
assign w22914 = ~w22911 & w22912;
assign w22915 = ~w22913 & ~w22914;
assign w22916 = ~w22910 & ~w22915;
assign w22917 = w22897 & ~w22916;
assign w22918 = w22910 & w22915;
assign w22919 = (~w22918 & w22653) | (~w22918 & w32502) | (w22653 & w32502);
assign w22920 = ~w22917 & w22919;
assign w22921 = ~w22654 & ~w22920;
assign w22922 = ~w21934 & w21973;
assign w22923 = w21999 & ~w22922;
assign w22924 = ~w21974 & ~w22923;
assign w22925 = (~w21963 & w21924) | (~w21963 & w37042) | (w21924 & w37042);
assign w22926 = ~w21934 & w21968;
assign w22927 = w21976 & ~w22926;
assign w22928 = (~w22924 & w21959) | (~w22924 & w37043) | (w21959 & w37043);
assign w22929 = ~w21959 & w37044;
assign w22930 = ~w22928 & ~w22929;
assign w22931 = w9456 & ~w22930;
assign w22932 = w8298 & ~w21968;
assign w22933 = w8277 & w21934;
assign w22934 = w8295 & ~w21973;
assign w22935 = ~w22932 & ~w22933;
assign w22936 = ~w22934 & w22935;
assign w22937 = a_8 & w22936;
assign w22938 = ~a_8 & ~w22936;
assign w22939 = ~w22937 & ~w22938;
assign w22940 = (w22939 & w22930) | (w22939 & w37045) | (w22930 & w37045);
assign w22941 = ~w22931 & ~w22940;
assign w22942 = ~w22575 & w32503;
assign w22943 = ~w22648 & ~w22942;
assign w22944 = w6998 & ~w21910;
assign w22945 = w6446 & w21892;
assign w22946 = w6996 & w21921;
assign w22947 = ~w22944 & ~w22945;
assign w22948 = ~w22946 & w22947;
assign w22949 = (w22948 & ~w22664) | (w22948 & w37046) | (~w22664 & w37046);
assign w22950 = a_14 & ~w22949;
assign w22951 = (~w22664 & w37047) | (~w22664 & w37048) | (w37047 & w37048);
assign w22952 = ~w22950 & ~w22951;
assign w22953 = ~w22239 & ~w22641;
assign w22954 = ~w22643 & w22953;
assign w22955 = ~w22640 & ~w22954;
assign w22956 = w8391 & w22555;
assign w22957 = w6059 & w21787;
assign w22958 = ~w21882 & w37049;
assign w22959 = (~w22957 & ~w21901) | (~w22957 & w37050) | (~w21901 & w37050);
assign w22960 = ~w22958 & w22959;
assign w22961 = a_17 & w22960;
assign w22962 = ~a_17 & ~w22960;
assign w22963 = ~w22961 & ~w22962;
assign w22964 = (w22963 & ~w22555) | (w22963 & w37051) | (~w22555 & w37051);
assign w22965 = ~w22956 & ~w22964;
assign w22966 = w5309 & w22247;
assign w22967 = w5309 & ~w22246;
assign w22968 = w5308 & w21833;
assign w22969 = w5816 & w21854;
assign w22970 = (~w22968 & w21839) | (~w22968 & w37052) | (w21839 & w37052);
assign w22971 = ~w22969 & w22970;
assign w22972 = (w22971 & ~w22967) | (w22971 & w32101) | (~w22967 & w32101);
assign w22973 = ~w22966 & w22972;
assign w22974 = a_20 & ~w22973;
assign w22975 = ~a_20 & w22973;
assign w22976 = ~w22974 & ~w22975;
assign w22977 = w21815 & w35766;
assign w22978 = w1226 & ~w22331;
assign w22979 = w4638 & w21815;
assign w22980 = (~w22979 & ~w21813) | (~w22979 & w37053) | (~w21813 & w37053);
assign w22981 = (w22977 & w22978) | (w22977 & w37054) | (w22978 & w37054);
assign w22982 = ~w22978 & w32102;
assign w22983 = ~w22981 & ~w22982;
assign w22984 = ~w22613 & ~w22616;
assign w22985 = w22612 & w37055;
assign w22986 = ~w22617 & ~w22985;
assign w22987 = (~w22983 & ~w22986) | (~w22983 & w32103) | (~w22986 & w32103);
assign w22988 = w22986 & w32104;
assign w22989 = ~w22987 & ~w22988;
assign w22990 = ~w22177 & w32105;
assign w22991 = (w5017 & w21819) | (w5017 & w32106) | (w21819 & w32106);
assign w22992 = w22177 & w22991;
assign w22993 = w5016 & w21807;
assign w22994 = w5286 & ~w21803;
assign w22995 = ~w21796 & w37056;
assign w22996 = ~w22993 & ~w22995;
assign w22997 = ~w22994 & w22996;
assign w22998 = ~w22992 & w22997;
assign w22999 = w22998 & w32107;
assign w23000 = (a_23 & ~w22998) | (a_23 & w32108) | (~w22998 & w32108);
assign w23001 = ~w22999 & ~w23000;
assign w23002 = w22989 & w23001;
assign w23003 = ~w22989 & ~w23001;
assign w23004 = ~w23002 & ~w23003;
assign w23005 = w22976 & w23004;
assign w23006 = ~w22976 & ~w23004;
assign w23007 = ~w23005 & ~w23006;
assign w23008 = ~w22603 & ~w22635;
assign w23009 = ~w22634 & ~w23008;
assign w23010 = w23007 & ~w23009;
assign w23011 = ~w23007 & w23009;
assign w23012 = ~w23010 & ~w23011;
assign w23013 = w22965 & w23012;
assign w23014 = ~w22965 & ~w23012;
assign w23015 = ~w23013 & ~w23014;
assign w23016 = w22955 & ~w23015;
assign w23017 = ~w22955 & w23015;
assign w23018 = ~w23016 & ~w23017;
assign w23019 = w22952 & ~w23018;
assign w23020 = ~w22952 & w23018;
assign w23021 = ~w23019 & ~w23020;
assign w23022 = w7489 & ~w21945;
assign w23023 = w7192 & w21951;
assign w23024 = w7511 & ~w21940;
assign w23025 = w22075 & w32109;
assign w23026 = ~w21912 & w23025;
assign w23027 = ~w21946 & ~w21960;
assign w23028 = (~w21961 & ~w21955) | (~w21961 & w32110) | (~w21955 & w32110);
assign w23029 = w23027 & ~w23028;
assign w23030 = ~w23026 & w23029;
assign w23031 = (~w23027 & w23026) | (~w23027 & w32504) | (w23026 & w32504);
assign w23032 = ~w23030 & ~w23031;
assign w23033 = ~w23022 & ~w23023;
assign w23034 = ~w23024 & w23033;
assign w23035 = (w23034 & ~w23032) | (w23034 & w37057) | (~w23032 & w37057);
assign w23036 = a_11 & ~w23035;
assign w23037 = (~w23032 & w37058) | (~w23032 & w37059) | (w37058 & w37059);
assign w23038 = ~w23036 & ~w23037;
assign w23039 = w23021 & w23038;
assign w23040 = ~w23021 & ~w23038;
assign w23041 = ~w23039 & ~w23040;
assign w23042 = w22943 & w23041;
assign w23043 = ~w22943 & ~w23041;
assign w23044 = ~w23042 & ~w23043;
assign w23045 = ~w22941 & ~w23044;
assign w23046 = w22921 & w23045;
assign w23047 = ~w22941 & w23044;
assign w23048 = ~w22921 & w23047;
assign w23049 = ~w23046 & ~w23048;
assign w23050 = w8295 & ~w21945;
assign w23051 = w8298 & w21951;
assign w23052 = w8277 & w21921;
assign w23053 = ~w23051 & ~w23052;
assign w23054 = ~w23050 & w23053;
assign w23055 = (w23054 & ~w22083) | (w23054 & w37060) | (~w22083 & w37060);
assign w23056 = a_8 & ~w23055;
assign w23057 = (~w22083 & w37061) | (~w22083 & w37062) | (w37061 & w37062);
assign w23058 = ~w23056 & ~w23057;
assign w23059 = ~w22891 & ~w22893;
assign w23060 = w22875 & ~w23059;
assign w23061 = ~w22875 & w23059;
assign w23062 = ~w23060 & ~w23061;
assign w23063 = ~w23058 & ~w23062;
assign w23064 = ~w22741 & w22864;
assign w23065 = ~w22865 & ~w23064;
assign w23066 = w8295 & w21892;
assign w23067 = w8298 & w21901;
assign w23068 = ~w21882 & w37063;
assign w23069 = ~w23066 & ~w23067;
assign w23070 = ~w23068 & w23069;
assign w23071 = (w22096 & w32505) | (w22096 & w32506) | (w32505 & w32506);
assign w23072 = (~w22096 & w32507) | (~w22096 & w32508) | (w32507 & w32508);
assign w23073 = ~w23071 & ~w23072;
assign w23074 = w23065 & w23073;
assign w23075 = ~w21882 & w37064;
assign w23076 = w8298 & w21787;
assign w23077 = w8277 & w21854;
assign w23078 = ~w22381 & w22382;
assign w23079 = ~w22383 & ~w23078;
assign w23080 = ~w23076 & ~w23077;
assign w23081 = ~w23075 & w23080;
assign w23082 = (~w23079 & w37065) | (~w23079 & w37066) | (w37065 & w37066);
assign w23083 = (w23079 & w37067) | (w23079 & w37068) | (w37067 & w37068);
assign w23084 = ~w23082 & ~w23083;
assign w23085 = ~w22774 & ~w22861;
assign w23086 = ~w22859 & w23085;
assign w23087 = w22859 & ~w23085;
assign w23088 = ~w23086 & ~w23087;
assign w23089 = ~w23084 & ~w23088;
assign w23090 = w8278 & w22107;
assign w23091 = w21873 & w32112;
assign w23092 = w8278 & ~w21854;
assign w23093 = ~w21787 & w23092;
assign w23094 = ~w23091 & ~w23093;
assign w23095 = ~w22105 & ~w23094;
assign w23096 = w8277 & ~w21839;
assign w23097 = w8298 & w21854;
assign w23098 = w8295 & w21787;
assign w23099 = ~w23096 & ~w23097;
assign w23100 = ~w23098 & w23099;
assign w23101 = ~w23095 & w23100;
assign w23102 = ~w23090 & w23101;
assign w23103 = a_8 & ~w23102;
assign w23104 = ~a_8 & w23102;
assign w23105 = ~w23103 & ~w23104;
assign w23106 = ~w22821 & ~w22854;
assign w23107 = w22853 & ~w22858;
assign w23108 = w23106 & ~w23107;
assign w23109 = ~w23106 & w23107;
assign w23110 = ~w23108 & ~w23109;
assign w23111 = w23105 & ~w23110;
assign w23112 = w8278 & w22247;
assign w23113 = w8278 & ~w22246;
assign w23114 = w8277 & w21833;
assign w23115 = w8295 & w21854;
assign w23116 = (~w23114 & w21839) | (~w23114 & w37069) | (w21839 & w37069);
assign w23117 = ~w23115 & w23116;
assign w23118 = (w23117 & ~w23113) | (w23117 & w32113) | (~w23113 & w32113);
assign w23119 = ~w23112 & w23118;
assign w23120 = a_8 & ~w23119;
assign w23121 = ~a_8 & w23119;
assign w23122 = ~w23120 & ~w23121;
assign w23123 = ~w22809 & ~w22854;
assign w23124 = w22820 & ~w23123;
assign w23125 = ~w22820 & w23123;
assign w23126 = ~w23124 & ~w23125;
assign w23127 = ~w23122 & w23126;
assign w23128 = w23122 & ~w23126;
assign w23129 = ~w23127 & ~w23128;
assign w23130 = (~w22798 & w37070) | (~w22798 & w37071) | (w37070 & w37071);
assign w23131 = ~w22800 & ~w23130;
assign w23132 = w22784 & w23131;
assign w23133 = ~w22784 & ~w23131;
assign w23134 = ~w23132 & ~w23133;
assign w23135 = w9456 & w22278;
assign w23136 = w8298 & w21833;
assign w23137 = w8277 & ~w21803;
assign w23138 = w8295 & ~w21839;
assign w23139 = ~w23136 & ~w23137;
assign w23140 = (~a_8 & w23138) | (~a_8 & w37072) | (w23138 & w37072);
assign w23141 = ~w23138 & w37073;
assign w23142 = ~w23140 & ~w23141;
assign w23143 = (w23142 & ~w22278) | (w23142 & w37074) | (~w22278 & w37074);
assign w23144 = ~w23135 & ~w23143;
assign w23145 = w23134 & w23144;
assign w23146 = (~w23134 & w23143) | (~w23134 & w32510) | (w23143 & w32510);
assign w23147 = w22792 & ~w22798;
assign w23148 = ~w22799 & ~w23147;
assign w23149 = ~w21823 & w32114;
assign w23150 = ~w22289 & ~w23149;
assign w23151 = w9456 & ~w23150;
assign w23152 = w9484 & ~w23150;
assign w23153 = ~w21796 & w37075;
assign w23154 = w8295 & w21833;
assign w23155 = (~w23153 & w21803) | (~w23153 & w37076) | (w21803 & w37076);
assign w23156 = ~w23154 & w23155;
assign w23157 = ~a_8 & ~w23156;
assign w23158 = a_8 & w23156;
assign w23159 = ~w23157 & ~w23158;
assign w23160 = ~w23152 & w23159;
assign w23161 = ~w23160 & w37077;
assign w23162 = (~w23148 & w23160) | (~w23148 & w32511) | (w23160 & w32511);
assign w23163 = ~w22137 & w32115;
assign w23164 = ~w21796 & w32116;
assign w23165 = w8277 & w21813;
assign w23166 = w8298 & w21807;
assign w23167 = (w8278 & w21817) | (w8278 & w32117) | (w21817 & w32117);
assign w23168 = w22137 & w23167;
assign w23169 = ~w23165 & ~w23166;
assign w23170 = ~w23164 & w23169;
assign w23171 = ~w23168 & w23170;
assign w23172 = ~w23163 & w23171;
assign w23173 = w8278 & ~w22331;
assign w23174 = w8298 & w21815;
assign w23175 = (~w23174 & ~w21813) | (~w23174 & w32118) | (~w21813 & w32118);
assign w23176 = ~w8272 & w21815;
assign w23177 = w21815 & w19105;
assign w23178 = (~w21813 & w37078) | (~w21813 & w37079) | (w37078 & w37079);
assign w23179 = (w23178 & w22331) | (w23178 & w37080) | (w22331 & w37080);
assign w23180 = (a_8 & w23173) | (a_8 & w32119) | (w23173 & w32119);
assign w23181 = w8278 & ~w22161;
assign w23182 = w8277 & w21815;
assign w23183 = w8295 & w21807;
assign w23184 = (~w23182 & ~w21813) | (~w23182 & w37081) | (~w21813 & w37081);
assign w23185 = ~w23183 & w23184;
assign w23186 = ~w23181 & w23185;
assign w23187 = ~w23180 & w23186;
assign w23188 = (w23186 & w32512) | (w23186 & w32513) | (w32512 & w32513);
assign w23189 = ~w23172 & ~w23188;
assign w23190 = w23171 & w32121;
assign w23191 = (~w22786 & ~w23186) | (~w22786 & w32514) | (~w23186 & w32514);
assign w23192 = ~w23190 & ~w23191;
assign w23193 = ~w23189 & w23192;
assign w23194 = (w22789 & w22331) | (w22789 & w37082) | (w22331 & w37082);
assign w23195 = w22787 & ~w23194;
assign w23196 = ~w22791 & ~w23195;
assign w23197 = w23193 & w23196;
assign w23198 = ~w23193 & ~w23196;
assign w23199 = (w8278 & w21819) | (w8278 & w32123) | (w21819 & w32123);
assign w23200 = w22177 & w23199;
assign w23201 = ~w21796 & w37083;
assign w23202 = w8295 & ~w21803;
assign w23203 = w8277 & w21807;
assign w23204 = ~w23201 & ~w23203;
assign w23205 = ~w23202 & w23204;
assign w23206 = ~w23200 & w23205;
assign w23207 = (a_8 & ~w23206) | (a_8 & w32124) | (~w23206 & w32124);
assign w23208 = w23206 & w32125;
assign w23209 = ~w23207 & ~w23208;
assign w23210 = ~w23198 & w23209;
assign w23211 = ~w23197 & ~w23210;
assign w23212 = (~w23161 & w23211) | (~w23161 & w37084) | (w23211 & w37084);
assign w23213 = ~w23146 & ~w23212;
assign w23214 = ~w23145 & ~w23213;
assign w23215 = w23129 & w23214;
assign w23216 = ~w23105 & w23110;
assign w23217 = ~w23127 & ~w23216;
assign w23218 = ~w23215 & w23217;
assign w23219 = ~w23111 & ~w23218;
assign w23220 = (~w23089 & w23218) | (~w23089 & w37085) | (w23218 & w37085);
assign w23221 = w23084 & w23088;
assign w23222 = w9456 & w22555;
assign w23223 = w8277 & w21787;
assign w23224 = ~w21882 & w37086;
assign w23225 = (~w23223 & ~w21901) | (~w23223 & w37087) | (~w21901 & w37087);
assign w23226 = ~w23224 & w23225;
assign w23227 = a_8 & w23226;
assign w23228 = ~a_8 & ~w23226;
assign w23229 = ~w23227 & ~w23228;
assign w23230 = (w23229 & ~w22555) | (w23229 & w37088) | (~w22555 & w37088);
assign w23231 = ~w23222 & ~w23230;
assign w23232 = ~w22757 & ~w22758;
assign w23233 = w22862 & w23232;
assign w23234 = ~w22862 & ~w23232;
assign w23235 = ~w23233 & ~w23234;
assign w23236 = w23231 & w23235;
assign w23237 = (~w23221 & ~w23235) | (~w23221 & w37089) | (~w23235 & w37089);
assign w23238 = ~w23220 & w23237;
assign w23239 = ~w23065 & ~w23073;
assign w23240 = ~w23231 & ~w23235;
assign w23241 = ~w23239 & ~w23240;
assign w23242 = (~w23074 & ~w23241) | (~w23074 & w37090) | (~w23241 & w37090);
assign w23243 = w9456 & ~w22580;
assign w23244 = w8298 & w21892;
assign w23245 = w8277 & w21901;
assign w23246 = w8295 & ~w21910;
assign w23247 = ~w23244 & ~w23245;
assign w23248 = w23247 & w37091;
assign w23249 = (~a_8 & ~w23247) | (~a_8 & w37092) | (~w23247 & w37092);
assign w23250 = ~w23248 & ~w23249;
assign w23251 = (w23250 & w22580) | (w23250 & w37093) | (w22580 & w37093);
assign w23252 = ~w23243 & ~w23251;
assign w23253 = ~w22739 & ~w22865;
assign w23254 = ~w22719 & ~w22866;
assign w23255 = w23253 & ~w23254;
assign w23256 = ~w23253 & w23254;
assign w23257 = ~w23255 & ~w23256;
assign w23258 = ~w23252 & ~w23257;
assign w23259 = w23252 & w23257;
assign w23260 = ~w23258 & ~w23259;
assign w23261 = w23242 & w23260;
assign w23262 = w8298 & ~w21910;
assign w23263 = w8277 & w21892;
assign w23264 = w8295 & w21921;
assign w23265 = ~w23262 & ~w23263;
assign w23266 = ~w23264 & w23265;
assign w23267 = (w23266 & ~w22664) | (w23266 & w37094) | (~w22664 & w37094);
assign w23268 = a_8 & ~w23267;
assign w23269 = (~w22664 & w37095) | (~w22664 & w37096) | (w37095 & w37096);
assign w23270 = ~w23268 & ~w23269;
assign w23271 = ~w22703 & ~w22871;
assign w23272 = w22869 & ~w23271;
assign w23273 = ~w22869 & w23271;
assign w23274 = ~w23272 & ~w23273;
assign w23275 = ~w23270 & w23274;
assign w23276 = ~w23258 & ~w23275;
assign w23277 = ~w23261 & w23276;
assign w23278 = w23270 & ~w23274;
assign w23279 = (~w22871 & w22869) | (~w22871 & w32515) | (w22869 & w32515);
assign w23280 = w8277 & ~w21910;
assign w23281 = w8298 & w21921;
assign w23282 = w8295 & w21951;
assign w23283 = ~w23280 & ~w23281;
assign w23284 = ~w23282 & w23283;
assign w23285 = ~a_8 & w23284;
assign w23286 = (w23285 & ~w32126) | (w23285 & w32516) | (~w32126 & w32516);
assign w23287 = ~w22901 & w32127;
assign w23288 = a_8 & ~w23284;
assign w23289 = ~w23287 & ~w23288;
assign w23290 = ~w23286 & w23289;
assign w23291 = ~w22688 & ~w22872;
assign w23292 = w23290 & ~w23291;
assign w23293 = w23279 & w23292;
assign w23294 = w23290 & w23291;
assign w23295 = ~w23279 & w23294;
assign w23296 = ~w23293 & ~w23295;
assign w23297 = ~w23278 & w23296;
assign w23298 = ~w23277 & w23297;
assign w23299 = ~w23279 & ~w23291;
assign w23300 = w23279 & w23291;
assign w23301 = ~w23299 & ~w23300;
assign w23302 = ~w23290 & ~w23301;
assign w23303 = ~w23298 & ~w23302;
assign w23304 = w23058 & w23062;
assign w23305 = ~w23063 & ~w23304;
assign w23306 = ~w23303 & w23305;
assign w23307 = ~w23063 & ~w23306;
assign w23308 = ~w21943 & ~w21960;
assign w23309 = (w23308 & w23026) | (w23308 & w32517) | (w23026 & w32517);
assign w23310 = w22925 & ~w23309;
assign w23311 = w8277 & ~w21945;
assign w23312 = w8295 & w21934;
assign w23313 = w8298 & ~w21940;
assign w23314 = ~w23311 & ~w23312;
assign w23315 = (a_8 & ~w23314) | (a_8 & w37097) | (~w23314 & w37097);
assign w23316 = w8278 & w23310;
assign w23317 = w23314 & w37098;
assign w23318 = ~w23316 & w23317;
assign w23319 = (~w23315 & ~w23310) | (~w23315 & w37099) | (~w23310 & w37099);
assign w23320 = ~w23318 & w23319;
assign w23321 = w22910 & ~w23320;
assign w23322 = w22915 & ~w23321;
assign w23323 = ~w22910 & ~w23320;
assign w23324 = ~w22915 & ~w23323;
assign w23325 = ~w23322 & ~w23324;
assign w23326 = w22897 & ~w23325;
assign w23327 = w22915 & ~w23323;
assign w23328 = ~w22915 & ~w23321;
assign w23329 = ~w23327 & ~w23328;
assign w23330 = ~w22897 & ~w23329;
assign w23331 = ~w23326 & ~w23330;
assign w23332 = ~w22892 & ~w22893;
assign w23333 = ~w22675 & ~w22894;
assign w23334 = w8298 & ~w21945;
assign w23335 = w8277 & w21951;
assign w23336 = w8295 & ~w21940;
assign w23337 = ~w23334 & ~w23335;
assign w23338 = ~w23336 & w23337;
assign w23339 = (w23338 & ~w23032) | (w23338 & w37100) | (~w23032 & w37100);
assign w23340 = ~a_8 & w23339;
assign w23341 = (w23032 & w37101) | (w23032 & w37102) | (w37101 & w37102);
assign w23342 = ~w23340 & ~w23341;
assign w23343 = w23333 & w23342;
assign w23344 = ~w23333 & ~w23342;
assign w23345 = ~w23343 & ~w23344;
assign w23346 = w23332 & w23345;
assign w23347 = ~w23332 & ~w23345;
assign w23348 = ~w23346 & ~w23347;
assign w23349 = ~w23331 & w23348;
assign w23350 = w23307 & w23349;
assign w23351 = w23332 & ~w23333;
assign w23352 = ~w23332 & w23333;
assign w23353 = ~w23351 & ~w23352;
assign w23354 = w23342 & ~w23353;
assign w23355 = ~w23331 & w23354;
assign w23356 = ~w22916 & ~w22918;
assign w23357 = ~w22897 & ~w23356;
assign w23358 = w22897 & w23356;
assign w23359 = ~w23357 & ~w23358;
assign w23360 = w23320 & ~w23359;
assign w23361 = ~w23355 & ~w23360;
assign w23362 = (~w22918 & ~w22897) | (~w22918 & w37103) | (~w22897 & w37103);
assign w23363 = ~w21940 & w21975;
assign w23364 = ~w22925 & ~w22927;
assign w23365 = (~w23363 & w21959) | (~w23363 & w37104) | (w21959 & w37104);
assign w23366 = ~w23364 & w23365;
assign w23367 = w9456 & ~w23366;
assign w23368 = w8298 & w21934;
assign w23369 = w8277 & ~w21940;
assign w23370 = w8295 & ~w21968;
assign w23371 = ~w23368 & ~w23369;
assign w23372 = (~a_8 & ~w23371) | (~a_8 & w37105) | (~w23371 & w37105);
assign w23373 = w23371 & w37106;
assign w23374 = ~w23372 & ~w23373;
assign w23375 = (w23374 & w23366) | (w23374 & w37107) | (w23366 & w37107);
assign w23376 = ~w23367 & ~w23375;
assign w23377 = ~w22089 & ~w23376;
assign w23378 = w22089 & w23376;
assign w23379 = ~w23377 & ~w23378;
assign w23380 = ~w22653 & w23379;
assign w23381 = w22653 & ~w23379;
assign w23382 = ~w23380 & ~w23381;
assign w23383 = w23362 & w23382;
assign w23384 = ~w23362 & ~w23382;
assign w23385 = ~w23383 & ~w23384;
assign w23386 = (~w23385 & w23350) | (~w23385 & w32518) | (w23350 & w32518);
assign w23387 = w23376 & w23385;
assign w23388 = w22941 & w23044;
assign w23389 = w22921 & w23388;
assign w23390 = w22941 & ~w23044;
assign w23391 = ~w22921 & w23390;
assign w23392 = ~w23389 & ~w23391;
assign w23393 = ~w23387 & w23392;
assign w23394 = (w23049 & ~w23393) | (w23049 & w32519) | (~w23393 & w32519);
assign w23395 = (~w21979 & w37108) | (~w21979 & w37109) | (w37108 & w37109);
assign w23396 = ~w22009 & ~w22017;
assign w23397 = ~w23395 & w23396;
assign w23398 = ~w22019 & ~w23397;
assign w23399 = ~w23397 & w37110;
assign w23400 = ~w23397 & w37111;
assign w23401 = w9780 & w22007;
assign w23402 = w9786 & ~w21992;
assign w23403 = w9788 & w22014;
assign w23404 = ~w23401 & ~w23402;
assign w23405 = ~w23403 & w23404;
assign w23406 = a_5 & w23405;
assign w23407 = ~a_5 & ~w23405;
assign w23408 = ~w23406 & ~w23407;
assign w23409 = ~w23400 & w23408;
assign w23410 = ~w23399 & ~w23409;
assign w23411 = ~w22921 & w23044;
assign w23412 = w22943 & ~w23021;
assign w23413 = ~w22943 & w23021;
assign w23414 = ~w23412 & ~w23413;
assign w23415 = w23038 & ~w23414;
assign w23416 = ~w23411 & ~w23415;
assign w23417 = (~w22648 & ~w23018) | (~w22648 & w32520) | (~w23018 & w32520);
assign w23418 = ~w22942 & w23417;
assign w23419 = ~w23019 & ~w23418;
assign w23420 = w6998 & w21921;
assign w23421 = w6996 & w21951;
assign w23422 = w6446 & ~w21910;
assign w23423 = ~w22901 & w37112;
assign w23424 = ~w23421 & w37113;
assign w23425 = ~w23423 & w37114;
assign w23426 = (a_14 & w23423) | (a_14 & w37115) | (w23423 & w37115);
assign w23427 = ~w23425 & ~w23426;
assign w23428 = w7192 & ~w21945;
assign w23429 = w7511 & w21934;
assign w23430 = w7489 & ~w21940;
assign w23431 = ~w23428 & ~w23429;
assign w23432 = (a_11 & ~w23431) | (a_11 & w37116) | (~w23431 & w37116);
assign w23433 = w7193 & w23310;
assign w23434 = w23431 & w37117;
assign w23435 = ~w23433 & w23434;
assign w23436 = (~w23432 & ~w23310) | (~w23432 & w37118) | (~w23310 & w37118);
assign w23437 = ~w23435 & w23436;
assign w23438 = w23427 & ~w23437;
assign w23439 = ~w22955 & ~w23013;
assign w23440 = (~w23014 & w22955) | (~w23014 & w32521) | (w22955 & w32521);
assign w23441 = w5309 & w22107;
assign w23442 = w21873 & w32129;
assign w23443 = w5309 & ~w21854;
assign w23444 = ~w21787 & w23443;
assign w23445 = ~w23442 & ~w23444;
assign w23446 = ~w22105 & ~w23445;
assign w23447 = w5308 & ~w21839;
assign w23448 = w5818 & w21854;
assign w23449 = w5816 & w21787;
assign w23450 = ~w23447 & ~w23448;
assign w23451 = ~w23449 & w23450;
assign w23452 = ~w23446 & w23451;
assign w23453 = ~w23441 & w23452;
assign w23454 = a_20 & ~w23453;
assign w23455 = ~a_20 & w23453;
assign w23456 = ~w23454 & ~w23455;
assign w23457 = ~w22987 & w23001;
assign w23458 = ~w22988 & ~w23457;
assign w23459 = (a_26 & w22978) | (a_26 & w37119) | (w22978 & w37119);
assign w23460 = w4666 & w21807;
assign w23461 = ~w518 & w21815;
assign w23462 = w1226 & ~w22161;
assign w23463 = (~w23461 & ~w21813) | (~w23461 & w37120) | (~w21813 & w37120);
assign w23464 = ~w23460 & w23463;
assign w23465 = ~w23462 & w23464;
assign w23466 = ~w23459 & w23465;
assign w23467 = w23459 & ~w23465;
assign w23468 = ~w23466 & ~w23467;
assign w23469 = w7961 & w22289;
assign w23470 = w7961 & w21830;
assign w23471 = w21824 & w23470;
assign w23472 = w5286 & ~w21224;
assign w23473 = w21207 & w23472;
assign w23474 = w5286 & w21224;
assign w23475 = ~w21207 & w23474;
assign w23476 = ~w23473 & ~w23475;
assign w23477 = (w5016 & ~w21156) | (w5016 & w32130) | (~w21156 & w32130);
assign w23478 = ~w21796 & w23477;
assign w23479 = w5080 & ~w21800;
assign w23480 = w21799 & w23479;
assign w23481 = w5080 & w21800;
assign w23482 = ~w21799 & w23481;
assign w23483 = ~w23480 & ~w23482;
assign w23484 = ~w23478 & w23483;
assign w23485 = w23476 & w23484;
assign w23486 = w7962 & w23485;
assign w23487 = a_23 & ~w23485;
assign w23488 = ~w23486 & ~w23487;
assign w23489 = ~w23471 & w23488;
assign w23490 = ~w23469 & w23489;
assign w23491 = (~a_23 & w21796) | (~a_23 & w32131) | (w21796 & w32131);
assign w23492 = w23483 & w23491;
assign w23493 = w23476 & w23492;
assign w23494 = ~w21830 & w23493;
assign w23495 = w21824 & w23494;
assign w23496 = w21830 & w23493;
assign w23497 = ~w21824 & w23496;
assign w23498 = ~w23495 & ~w23497;
assign w23499 = (~w23468 & ~w23490) | (~w23468 & w32522) | (~w23490 & w32522);
assign w23500 = w23468 & w23498;
assign w23501 = w23490 & w23500;
assign w23502 = ~w23499 & ~w23501;
assign w23503 = w23458 & ~w23502;
assign w23504 = ~w23458 & w23502;
assign w23505 = ~w23503 & ~w23504;
assign w23506 = ~w23456 & ~w23505;
assign w23507 = w23456 & w23505;
assign w23508 = ~w23506 & ~w23507;
assign w23509 = ~w23006 & ~w23009;
assign w23510 = ~w23005 & ~w23509;
assign w23511 = w23508 & w23510;
assign w23512 = ~w23508 & ~w23510;
assign w23513 = ~w23511 & ~w23512;
assign w23514 = w6061 & w21901;
assign w23515 = w6304 & w21892;
assign w23516 = ~w21882 & w37121;
assign w23517 = ~w23514 & ~w23515;
assign w23518 = ~w23516 & w23517;
assign w23519 = (w22096 & w32523) | (w22096 & w32524) | (w32523 & w32524);
assign w23520 = (~w22096 & w32525) | (~w22096 & w32526) | (w32525 & w32526);
assign w23521 = ~w23519 & ~w23520;
assign w23522 = ~w23513 & w23521;
assign w23523 = w23513 & ~w23521;
assign w23524 = ~w23522 & ~w23523;
assign w23525 = w23440 & w23524;
assign w23526 = ~w23440 & ~w23524;
assign w23527 = ~w23525 & ~w23526;
assign w23528 = ~w23438 & w23527;
assign w23529 = ~w23427 & ~w23437;
assign w23530 = ~w23527 & ~w23529;
assign w23531 = ~w23528 & ~w23530;
assign w23532 = w23419 & ~w23531;
assign w23533 = w23527 & ~w23529;
assign w23534 = ~w23438 & ~w23527;
assign w23535 = ~w23533 & ~w23534;
assign w23536 = ~w23419 & ~w23535;
assign w23537 = ~w23532 & ~w23536;
assign w23538 = ~w23427 & w23437;
assign w23539 = w23527 & ~w23538;
assign w23540 = w23427 & w23437;
assign w23541 = ~w23527 & ~w23540;
assign w23542 = ~w23539 & ~w23541;
assign w23543 = w23419 & w23542;
assign w23544 = w23527 & ~w23540;
assign w23545 = ~w23527 & ~w23538;
assign w23546 = ~w23544 & ~w23545;
assign w23547 = ~w23419 & w23546;
assign w23548 = ~w23543 & ~w23547;
assign w23549 = ~w23537 & w23548;
assign w23550 = (~w21999 & w21959) | (~w21999 & w37122) | (w21959 & w37122);
assign w23551 = ~w21998 & ~w23550;
assign w23552 = (w22000 & w21959) | (w22000 & w37123) | (w21959 & w37123);
assign w23553 = ~w23551 & ~w23552;
assign w23554 = ~w23551 & w37124;
assign w23555 = ~w23551 & w37125;
assign w23556 = w8295 & w21985;
assign w23557 = w8277 & ~w21968;
assign w23558 = w8298 & ~w21973;
assign w23559 = ~w23556 & ~w23557;
assign w23560 = w23559 & w37126;
assign w23561 = (~a_8 & ~w23559) | (~a_8 & w37127) | (~w23559 & w37127);
assign w23562 = ~w23560 & ~w23561;
assign w23563 = ~w23555 & w23562;
assign w23564 = ~w23554 & ~w23563;
assign w23565 = ~w23549 & w23564;
assign w23566 = w23549 & ~w23564;
assign w23567 = ~w23565 & ~w23566;
assign w23568 = w23416 & ~w23567;
assign w23569 = ~w23416 & w23567;
assign w23570 = ~w23568 & ~w23569;
assign w23571 = w23410 & w23570;
assign w23572 = w23394 & w23571;
assign w23573 = w23410 & ~w23570;
assign w23574 = ~w23394 & w23573;
assign w23575 = ~w23572 & ~w23574;
assign w23576 = w9788 & w22007;
assign w23577 = w9780 & ~w21992;
assign w23578 = w9786 & w21985;
assign w23579 = (w21979 & w37128) | (w21979 & w37129) | (w37128 & w37129);
assign w23580 = ~w23395 & ~w23579;
assign w23581 = ~w23577 & ~w23578;
assign w23582 = ~w23576 & w23581;
assign w23583 = (w23582 & ~w23580) | (w23582 & w37130) | (~w23580 & w37130);
assign w23584 = a_5 & ~w23583;
assign w23585 = (~w23580 & w37131) | (~w23580 & w37132) | (w37131 & w37132);
assign w23586 = ~w23584 & ~w23585;
assign w23587 = ~w23386 & ~w23387;
assign w23588 = w23049 & w23392;
assign w23589 = ~w23587 & ~w23588;
assign w23590 = w23587 & w23588;
assign w23591 = ~w23589 & ~w23590;
assign w23592 = w23586 & ~w23591;
assign w23593 = w23575 & ~w23592;
assign w23594 = ~w23410 & ~w23570;
assign w23595 = w23394 & w23594;
assign w23596 = ~w23410 & w23570;
assign w23597 = ~w23394 & w23596;
assign w23598 = ~w23595 & ~w23597;
assign w23599 = ~w23593 & w23598;
assign w23600 = w23586 & w23588;
assign w23601 = ~w23586 & ~w23588;
assign w23602 = ~w23600 & ~w23601;
assign w23603 = w23587 & w23602;
assign w23604 = ~w23587 & ~w23602;
assign w23605 = ~w23603 & ~w23604;
assign w23606 = w23307 & w23348;
assign w23607 = ~w23307 & ~w23348;
assign w23608 = ~w23606 & ~w23607;
assign w23609 = w10033 & ~w22930;
assign w23610 = w9780 & ~w21968;
assign w23611 = w9786 & w21934;
assign w23612 = w9788 & ~w21973;
assign w23613 = ~w23610 & ~w23611;
assign w23614 = ~w23612 & w23613;
assign w23615 = a_5 & w23614;
assign w23616 = ~a_5 & ~w23614;
assign w23617 = ~w23615 & ~w23616;
assign w23618 = (w23617 & w22930) | (w23617 & w37133) | (w22930 & w37133);
assign w23619 = ~w23609 & ~w23618;
assign w23620 = ~w23608 & ~w23619;
assign w23621 = w9786 & ~w21945;
assign w23622 = w9788 & w21934;
assign w23623 = w9780 & ~w21940;
assign w23624 = ~w23621 & ~w23622;
assign w23625 = ~w23623 & w23624;
assign w23626 = (w23625 & ~w23310) | (w23625 & w37134) | (~w23310 & w37134);
assign w23627 = a_5 & ~w23626;
assign w23628 = (~w23310 & w37135) | (~w23310 & w37136) | (w37135 & w37136);
assign w23629 = ~w23627 & ~w23628;
assign w23630 = ~w23277 & ~w23278;
assign w23631 = w23296 & ~w23302;
assign w23632 = w23630 & ~w23631;
assign w23633 = ~w23630 & w23631;
assign w23634 = ~w23632 & ~w23633;
assign w23635 = w23629 & w23634;
assign w23636 = w10033 & ~w22580;
assign w23637 = w9786 & w21901;
assign w23638 = w9780 & w21892;
assign w23639 = w9788 & ~w21910;
assign w23640 = ~w23637 & ~w23638;
assign w23641 = w23640 & w37137;
assign w23642 = (~a_5 & ~w23640) | (~a_5 & w37138) | (~w23640 & w37138);
assign w23643 = ~w23641 & ~w23642;
assign w23644 = (w23643 & w22580) | (w23643 & w37139) | (w22580 & w37139);
assign w23645 = ~w23636 & ~w23644;
assign w23646 = ~w23089 & ~w23221;
assign w23647 = w23219 & ~w23646;
assign w23648 = ~w23219 & w23646;
assign w23649 = ~w23647 & ~w23648;
assign w23650 = ~w23645 & ~w23649;
assign w23651 = ~w23129 & ~w23214;
assign w23652 = ~w23215 & ~w23651;
assign w23653 = w10033 & w22555;
assign w23654 = w9786 & w21787;
assign w23655 = ~w21882 & w37140;
assign w23656 = (~w23654 & ~w21901) | (~w23654 & w37141) | (~w21901 & w37141);
assign w23657 = ~w23655 & w23656;
assign w23658 = a_5 & w23657;
assign w23659 = ~a_5 & ~w23657;
assign w23660 = ~w23658 & ~w23659;
assign w23661 = (w23660 & ~w22555) | (w23660 & w37142) | (~w22555 & w37142);
assign w23662 = ~w23653 & ~w23661;
assign w23663 = w23652 & ~w23662;
assign w23664 = ~w21882 & w37143;
assign w23665 = w9786 & w21854;
assign w23666 = w9780 & w21787;
assign w23667 = ~w23665 & ~w23666;
assign w23668 = ~w23664 & w23667;
assign w23669 = (~w23079 & w37144) | (~w23079 & w37145) | (w37144 & w37145);
assign w23670 = (w23079 & w37146) | (w23079 & w37147) | (w37146 & w37147);
assign w23671 = ~w23669 & ~w23670;
assign w23672 = ~w23145 & ~w23146;
assign w23673 = ~w23212 & w23672;
assign w23674 = w23212 & ~w23672;
assign w23675 = ~w23673 & ~w23674;
assign w23676 = w23671 & w23675;
assign w23677 = ~w23671 & ~w23675;
assign w23678 = ~w23676 & ~w23677;
assign w23679 = w10033 & ~w22726;
assign w23680 = w9786 & ~w21839;
assign w23681 = w9780 & w21854;
assign w23682 = w9788 & w21787;
assign w23683 = ~w23680 & ~w23681;
assign w23684 = ~w23682 & w23683;
assign w23685 = a_5 & ~w23684;
assign w23686 = ~a_5 & w23684;
assign w23687 = (w23686 & w22726) | (w23686 & w37148) | (w22726 & w37148);
assign w23688 = ~w23679 & ~w23685;
assign w23689 = ~w23687 & w23688;
assign w23690 = ~w23161 & ~w23162;
assign w23691 = ~w23211 & w23690;
assign w23692 = w23211 & ~w23690;
assign w23693 = ~w23691 & ~w23692;
assign w23694 = ~w23689 & ~w23693;
assign w23695 = w23689 & w23693;
assign w23696 = ~w23694 & ~w23695;
assign w23697 = w22245 & ~w22246;
assign w23698 = ~w22247 & ~w23697;
assign w23699 = w9786 & w21833;
assign w23700 = w9780 & ~w21839;
assign w23701 = (~w23699 & ~w21854) | (~w23699 & w37149) | (~w21854 & w37149);
assign w23702 = ~w23700 & w23701;
assign w23703 = (~w23698 & w37150) | (~w23698 & w37151) | (w37150 & w37151);
assign w23704 = (w23698 & w37152) | (w23698 & w37153) | (w37152 & w37153);
assign w23705 = ~w23703 & ~w23704;
assign w23706 = ~w23197 & ~w23198;
assign w23707 = w23209 & w23706;
assign w23708 = ~w23209 & ~w23706;
assign w23709 = ~w23707 & ~w23708;
assign w23710 = ~w23705 & ~w23709;
assign w23711 = w23705 & w23709;
assign w23712 = (~w23186 & w37154) | (~w23186 & w37155) | (w37154 & w37155);
assign w23713 = ~w23188 & ~w23712;
assign w23714 = w23172 & w23713;
assign w23715 = ~w23172 & ~w23713;
assign w23716 = ~w23714 & ~w23715;
assign w23717 = w10033 & w22278;
assign w23718 = w9780 & w21833;
assign w23719 = w9786 & ~w21803;
assign w23720 = w9788 & ~w21839;
assign w23721 = ~w23718 & ~w23719;
assign w23722 = (~a_5 & w23720) | (~a_5 & w37156) | (w23720 & w37156);
assign w23723 = ~w23720 & w37157;
assign w23724 = ~w23722 & ~w23723;
assign w23725 = (w23724 & ~w22278) | (w23724 & w37158) | (~w22278 & w37158);
assign w23726 = ~w23717 & ~w23725;
assign w23727 = ~w23716 & ~w23726;
assign w23728 = ~w23725 & w32529;
assign w23729 = ~w21818 & w22137;
assign w23730 = ~w22138 & ~w23729;
assign w23731 = w9780 & w21807;
assign w23732 = w9786 & w21813;
assign w23733 = ~w21796 & w37159;
assign w23734 = ~w23731 & ~w23732;
assign w23735 = ~w23733 & w23734;
assign w23736 = (w23735 & w23730) | (w23735 & w32133) | (w23730 & w32133);
assign w23737 = w9776 & w21815;
assign w23738 = w21815 & w36589;
assign w23739 = w9790 & ~w22331;
assign w23740 = w9788 & w21813;
assign w23741 = w9780 & w21815;
assign w23742 = (~w23741 & ~w21813) | (~w23741 & w37160) | (~w21813 & w37160);
assign w23743 = (w23742 & w22331) | (w23742 & w37161) | (w22331 & w37161);
assign w23744 = ~w23739 & w32134;
assign w23745 = (a_5 & w23739) | (a_5 & w32530) | (w23739 & w32530);
assign w23746 = w9788 & w21807;
assign w23747 = w9786 & w21815;
assign w23748 = w9790 & ~w22161;
assign w23749 = (~w23747 & ~w21813) | (~w23747 & w37162) | (~w21813 & w37162);
assign w23750 = ~w23746 & w23749;
assign w23751 = ~w23748 & w23750;
assign w23752 = ~w23745 & w23751;
assign w23753 = (a_5 & ~w23751) | (a_5 & w32531) | (~w23751 & w32531);
assign w23754 = w23176 & ~w23753;
assign w23755 = ~w23736 & ~w23754;
assign w23756 = (~w23176 & ~w23751) | (~w23176 & w37163) | (~w23751 & w37163);
assign w23757 = (w23730 & w32532) | (w23730 & w32533) | (w32532 & w32533);
assign w23758 = ~w23756 & ~w23757;
assign w23759 = ~w23755 & w23758;
assign w23760 = (w23175 & w22331) | (w23175 & w37164) | (w22331 & w37164);
assign w23761 = w23177 & ~w23760;
assign w23762 = ~w23179 & ~w23761;
assign w23763 = w23759 & w23762;
assign w23764 = ~w21822 & w22177;
assign w23765 = ~w22178 & ~w23764;
assign w23766 = w9786 & w21807;
assign w23767 = w9788 & ~w21803;
assign w23768 = ~w21796 & w37165;
assign w23769 = ~w23766 & ~w23768;
assign w23770 = ~w23767 & w23769;
assign w23771 = (w23765 & w32534) | (w23765 & w32535) | (w32534 & w32535);
assign w23772 = (~w23765 & w32536) | (~w23765 & w32537) | (w32536 & w32537);
assign w23773 = ~w23771 & ~w23772;
assign w23774 = ~w23763 & ~w23773;
assign w23775 = w10061 & ~w23150;
assign w23776 = w23180 & ~w23186;
assign w23777 = ~w23187 & ~w23776;
assign w23778 = w9788 & w21833;
assign w23779 = ~w21796 & w37166;
assign w23780 = (~w23779 & w21803) | (~w23779 & w37167) | (w21803 & w37167);
assign w23781 = ~w23778 & w23780;
assign w23782 = ~a_5 & w23781;
assign w23783 = a_5 & ~w23781;
assign w23784 = ~w23782 & ~w23783;
assign w23785 = ~w23777 & ~w23784;
assign w23786 = ~w23775 & w23785;
assign w23787 = ~w23150 & w37168;
assign w23788 = ~w23786 & ~w23787;
assign w23789 = ~w23759 & ~w23762;
assign w23790 = ~w23786 & w32538;
assign w23791 = ~w23775 & ~w23784;
assign w23792 = (w23777 & w23150) | (w23777 & w37169) | (w23150 & w37169);
assign w23793 = ~w23791 & w23792;
assign w23794 = (~w23793 & ~w23790) | (~w23793 & w32136) | (~w23790 & w32136);
assign w23795 = ~w23728 & w23794;
assign w23796 = ~w23727 & ~w23795;
assign w23797 = (~w23710 & w23796) | (~w23710 & w37170) | (w23796 & w37170);
assign w23798 = w23696 & ~w23797;
assign w23799 = (~w23694 & ~w23696) | (~w23694 & w37171) | (~w23696 & w37171);
assign w23800 = w23678 & w23799;
assign w23801 = ~w23652 & w23662;
assign w23802 = (~w23676 & w23652) | (~w23676 & w37172) | (w23652 & w37172);
assign w23803 = ~w23800 & w23802;
assign w23804 = ~w23663 & ~w23803;
assign w23805 = ~w21882 & w37173;
assign w23806 = w9780 & w21901;
assign w23807 = w9788 & w21892;
assign w23808 = ~w23805 & ~w23806;
assign w23809 = ~w23807 & w23808;
assign w23810 = (w23809 & ~w22096) | (w23809 & w37174) | (~w22096 & w37174);
assign w23811 = a_5 & w23810;
assign w23812 = (w22096 & w37175) | (w22096 & w37176) | (w37175 & w37176);
assign w23813 = ~w23811 & ~w23812;
assign w23814 = ~w23111 & ~w23216;
assign w23815 = (~w23127 & ~w23129) | (~w23127 & w37177) | (~w23129 & w37177);
assign w23816 = ~w23814 & w23815;
assign w23817 = w23814 & ~w23815;
assign w23818 = ~w23816 & ~w23817;
assign w23819 = ~w23813 & ~w23818;
assign w23820 = w23813 & w23818;
assign w23821 = ~w23819 & ~w23820;
assign w23822 = w23804 & w23821;
assign w23823 = w23645 & w23649;
assign w23824 = (~w23819 & ~w23649) | (~w23819 & w37178) | (~w23649 & w37178);
assign w23825 = ~w23822 & w23824;
assign w23826 = ~w23650 & ~w23825;
assign w23827 = w9780 & ~w21910;
assign w23828 = w9786 & w21892;
assign w23829 = w9788 & w21921;
assign w23830 = ~w23827 & ~w23828;
assign w23831 = ~w23829 & w23830;
assign w23832 = (w23831 & ~w22664) | (w23831 & w37179) | (~w22664 & w37179);
assign w23833 = a_5 & w23832;
assign w23834 = (w22664 & w37180) | (w22664 & w37181) | (w37180 & w37181);
assign w23835 = ~w23833 & ~w23834;
assign w23836 = ~w23236 & ~w23240;
assign w23837 = (~w23221 & w23219) | (~w23221 & w32539) | (w23219 & w32539);
assign w23838 = ~w23836 & w23837;
assign w23839 = w23836 & ~w23837;
assign w23840 = ~w23838 & ~w23839;
assign w23841 = ~w23835 & w23840;
assign w23842 = w23835 & ~w23840;
assign w23843 = ~w23841 & ~w23842;
assign w23844 = ~w22901 & w37182;
assign w23845 = w9786 & ~w21910;
assign w23846 = w9788 & w21951;
assign w23847 = w9780 & w21921;
assign w23848 = ~w23846 & w37183;
assign w23849 = a_5 & ~w23848;
assign w23850 = ~w22901 & w37184;
assign w23851 = ~a_5 & w23848;
assign w23852 = ~w23850 & w23851;
assign w23853 = ~w23844 & ~w23849;
assign w23854 = ~w23852 & w23853;
assign w23855 = ~w23238 & ~w23240;
assign w23856 = ~w23074 & ~w23239;
assign w23857 = w23855 & w23856;
assign w23858 = ~w23855 & ~w23856;
assign w23859 = ~w23857 & ~w23858;
assign w23860 = ~w23854 & ~w23859;
assign w23861 = w23843 & ~w23860;
assign w23862 = w23826 & w23861;
assign w23863 = w23854 & w23859;
assign w23864 = (~w23841 & ~w23859) | (~w23841 & w32540) | (~w23859 & w32540);
assign w23865 = ~w23860 & ~w23864;
assign w23866 = ~w23862 & ~w23865;
assign w23867 = ~w23242 & ~w23260;
assign w23868 = ~w23261 & ~w23867;
assign w23869 = w9788 & ~w21945;
assign w23870 = w9786 & w21921;
assign w23871 = w9780 & w21951;
assign w23872 = ~w23870 & ~w23871;
assign w23873 = ~w23869 & w23872;
assign w23874 = (w23873 & ~w22083) | (w23873 & w37185) | (~w22083 & w37185);
assign w23875 = a_5 & ~w23874;
assign w23876 = (~w22083 & w37186) | (~w22083 & w37187) | (w37186 & w37187);
assign w23877 = ~w23875 & ~w23876;
assign w23878 = ~w23868 & w23877;
assign w23879 = w23868 & ~w23877;
assign w23880 = ~w23878 & ~w23879;
assign w23881 = ~w23866 & w23880;
assign w23882 = w9780 & ~w21945;
assign w23883 = w9786 & w21951;
assign w23884 = w9788 & ~w21940;
assign w23885 = ~w23882 & ~w23883;
assign w23886 = ~w23884 & w23885;
assign w23887 = (w23886 & ~w23032) | (w23886 & w37188) | (~w23032 & w37188);
assign w23888 = a_5 & ~w23887;
assign w23889 = (~w23032 & w37189) | (~w23032 & w37190) | (w37189 & w37190);
assign w23890 = ~w23888 & ~w23889;
assign w23891 = (~w23258 & ~w23260) | (~w23258 & w37191) | (~w23260 & w37191);
assign w23892 = ~w23275 & ~w23278;
assign w23893 = w23891 & w23892;
assign w23894 = ~w23891 & ~w23892;
assign w23895 = ~w23893 & ~w23894;
assign w23896 = w23890 & w23895;
assign w23897 = (~w23878 & ~w23895) | (~w23878 & w32541) | (~w23895 & w32541);
assign w23898 = ~w23881 & w23897;
assign w23899 = ~w23890 & ~w23895;
assign w23900 = ~w23629 & ~w23634;
assign w23901 = (~w23899 & w23634) | (~w23899 & w37192) | (w23634 & w37192);
assign w23902 = ~w23898 & w23901;
assign w23903 = ~w23635 & ~w23902;
assign w23904 = w23303 & ~w23305;
assign w23905 = ~w23306 & ~w23904;
assign w23906 = w9780 & w21934;
assign w23907 = w9786 & ~w21940;
assign w23908 = w9788 & ~w21968;
assign w23909 = ~w23906 & ~w23907;
assign w23910 = (a_5 & ~w23909) | (a_5 & w37193) | (~w23909 & w37193);
assign w23911 = w9790 & ~w23366;
assign w23912 = w23909 & w37194;
assign w23913 = ~w23911 & w23912;
assign w23914 = (~w23910 & w23366) | (~w23910 & w37195) | (w23366 & w37195);
assign w23915 = ~w23913 & w23914;
assign w23916 = ~w23905 & w23915;
assign w23917 = w23905 & ~w23915;
assign w23918 = ~w23916 & ~w23917;
assign w23919 = ~w23903 & w23918;
assign w23920 = w23608 & w23619;
assign w23921 = (~w23916 & ~w23608) | (~w23916 & w32542) | (~w23608 & w32542);
assign w23922 = (~w23620 & w23919) | (~w23620 & w32543) | (w23919 & w32543);
assign w23923 = ~w23350 & w37196;
assign w23924 = ~w23386 & ~w23923;
assign w23925 = w9788 & ~w21992;
assign w23926 = w9786 & ~w21973;
assign w23927 = w9780 & w21985;
assign w23928 = ~w23552 & w37197;
assign w23929 = (~w21995 & w23552) | (~w21995 & w37198) | (w23552 & w37198);
assign w23930 = ~w23928 & ~w23929;
assign w23931 = ~w23926 & ~w23927;
assign w23932 = ~w23925 & w23931;
assign w23933 = (w23932 & w23930) | (w23932 & w37199) | (w23930 & w37199);
assign w23934 = a_5 & w23933;
assign w23935 = (~w23930 & w37200) | (~w23930 & w37201) | (w37200 & w37201);
assign w23936 = ~w23934 & ~w23935;
assign w23937 = (w23936 & w23923) | (w23936 & w32544) | (w23923 & w32544);
assign w23938 = (~w23354 & ~w23307) | (~w23354 & w32545) | (~w23307 & w32545);
assign w23939 = ~w23331 & ~w23360;
assign w23940 = w9788 & w21985;
assign w23941 = w9786 & ~w21968;
assign w23942 = w9780 & ~w21973;
assign w23943 = ~w23551 & w37202;
assign w23944 = ~w23940 & ~w23941;
assign w23945 = ~w23942 & w23944;
assign w23946 = ~w23943 & w37203;
assign w23947 = (a_5 & w23943) | (a_5 & w37204) | (w23943 & w37204);
assign w23948 = ~w23946 & ~w23947;
assign w23949 = ~w23360 & w37205;
assign w23950 = (~w23948 & w23360) | (~w23948 & w37206) | (w23360 & w37206);
assign w23951 = ~w23949 & ~w23950;
assign w23952 = w23938 & w23951;
assign w23953 = ~w23938 & ~w23951;
assign w23954 = ~w23952 & ~w23953;
assign w23955 = ~w23937 & ~w23954;
assign w23956 = w23922 & w23955;
assign w23957 = w23924 & ~w23936;
assign w23958 = ~w23938 & ~w23939;
assign w23959 = w23938 & w23939;
assign w23960 = ~w23958 & ~w23959;
assign w23961 = w23948 & ~w23960;
assign w23962 = ~w23937 & w23961;
assign w23963 = ~w23957 & ~w23962;
assign w23964 = ~w23956 & w23963;
assign w23965 = w23598 & ~w23605;
assign w23966 = ~w23964 & w23965;
assign w23967 = ~w23599 & ~w23966;
assign w23968 = ~w23416 & w23565;
assign w23969 = w23549 & w23564;
assign w23970 = w23416 & w23969;
assign w23971 = ~w23968 & ~w23970;
assign w23972 = (w23971 & ~w23394) | (w23971 & w37207) | (~w23394 & w37207);
assign w23973 = w23044 & ~w23537;
assign w23974 = ~w22921 & w23973;
assign w23975 = ~w23415 & w23548;
assign w23976 = ~w23537 & ~w23975;
assign w23977 = ~w23974 & ~w23976;
assign w23978 = w23427 & w23527;
assign w23979 = w23419 & ~w23978;
assign w23980 = ~w23427 & ~w23527;
assign w23981 = (~w23980 & ~w23419) | (~w23980 & w37208) | (~w23419 & w37208);
assign w23982 = w9456 & ~w23930;
assign w23983 = w8298 & w21985;
assign w23984 = w8277 & ~w21973;
assign w23985 = w8295 & ~w21992;
assign w23986 = ~w23983 & ~w23984;
assign w23987 = w23986 & w37209;
assign w23988 = (~a_8 & ~w23986) | (~a_8 & w37210) | (~w23986 & w37210);
assign w23989 = ~w23987 & ~w23988;
assign w23990 = (w23989 & w23930) | (w23989 & w37211) | (w23930 & w37211);
assign w23991 = ~w23982 & ~w23990;
assign w23992 = w23981 & ~w23991;
assign w23993 = ~w23014 & ~w23523;
assign w23994 = ~w23439 & w23993;
assign w23995 = ~w23522 & ~w23994;
assign w23996 = w8391 & ~w22580;
assign w23997 = w6061 & w21892;
assign w23998 = w6059 & w21901;
assign w23999 = w6304 & ~w21910;
assign w24000 = ~w23997 & ~w23998;
assign w24001 = w24000 & w37212;
assign w24002 = (~a_17 & ~w24000) | (~a_17 & w37213) | (~w24000 & w37213);
assign w24003 = ~w24001 & ~w24002;
assign w24004 = (w24003 & w22580) | (w24003 & w37214) | (w22580 & w37214);
assign w24005 = ~w23996 & ~w24004;
assign w24006 = ~w21882 & w32138;
assign w24007 = ~w22381 & w24006;
assign w24008 = ~w21882 & w32139;
assign w24009 = w5308 & w21854;
assign w24010 = w5818 & w21787;
assign w24011 = ~w24009 & ~w24010;
assign w24012 = ~w24008 & w24011;
assign w24013 = ~w24007 & w24012;
assign w24014 = (a_20 & ~w24013) | (a_20 & w32140) | (~w24013 & w32140);
assign w24015 = w24013 & w32141;
assign w24016 = ~w24014 & ~w24015;
assign w24017 = ~w22988 & ~w23501;
assign w24018 = (~w23499 & ~w24017) | (~w23499 & w32546) | (~w24017 & w32546);
assign w24019 = (a_26 & ~w23465) | (a_26 & w37215) | (~w23465 & w37215);
assign w24020 = w3954 & w21815;
assign w24021 = ~w22137 & w32142;
assign w24022 = ~w21796 & w32143;
assign w24023 = w4638 & w21807;
assign w24024 = ~w518 & w21813;
assign w24025 = (w1226 & w21817) | (w1226 & w32144) | (w21817 & w32144);
assign w24026 = w22137 & w24025;
assign w24027 = ~w24023 & ~w24024;
assign w24028 = ~w24022 & w24027;
assign w24029 = ~w24026 & w24028;
assign w24030 = w24029 & w32145;
assign w24031 = (~w24020 & ~w24029) | (~w24020 & w32146) | (~w24029 & w32146);
assign w24032 = ~w24030 & ~w24031;
assign w24033 = ~w24019 & w24032;
assign w24034 = w24019 & ~w24032;
assign w24035 = ~w24033 & ~w24034;
assign w24036 = w5286 & ~w21839;
assign w24037 = w5080 & w21833;
assign w24038 = w5016 & ~w21803;
assign w24039 = ~w24037 & ~w24038;
assign w24040 = (a_23 & w24036) | (a_23 & w37216) | (w24036 & w37216);
assign w24041 = ~w24036 & w37217;
assign w24042 = ~w24040 & ~w24041;
assign w24043 = ~w22278 & w24042;
assign w24044 = ~w7961 & ~w7962;
assign w24045 = ~w24036 & w37218;
assign w24046 = ~w24040 & ~w24045;
assign w24047 = w22278 & w24046;
assign w24048 = ~w24043 & ~w24047;
assign w24049 = w24035 & ~w24048;
assign w24050 = ~w24035 & w24048;
assign w24051 = ~w24049 & ~w24050;
assign w24052 = w24018 & ~w24051;
assign w24053 = ~w24018 & w24051;
assign w24054 = ~w24052 & ~w24053;
assign w24055 = w24016 & ~w24054;
assign w24056 = ~w24016 & w24054;
assign w24057 = ~w24055 & ~w24056;
assign w24058 = ~w23506 & ~w23511;
assign w24059 = w24057 & w24058;
assign w24060 = ~w24057 & ~w24058;
assign w24061 = ~w24059 & ~w24060;
assign w24062 = ~w24005 & ~w24061;
assign w24063 = w24005 & w24061;
assign w24064 = ~w24062 & ~w24063;
assign w24065 = w23995 & w24064;
assign w24066 = ~w23995 & ~w24064;
assign w24067 = ~w24065 & ~w24066;
assign w24068 = w6996 & ~w21945;
assign w24069 = w6998 & w21951;
assign w24070 = w6446 & w21921;
assign w24071 = ~w24069 & ~w24070;
assign w24072 = ~w24068 & w24071;
assign w24073 = (w24072 & ~w22083) | (w24072 & w37219) | (~w22083 & w37219);
assign w24074 = a_14 & ~w24073;
assign w24075 = (~w22083 & w37220) | (~w22083 & w37221) | (w37220 & w37221);
assign w24076 = ~w24074 & ~w24075;
assign w24077 = ~w24067 & w24076;
assign w24078 = w24067 & ~w24076;
assign w24079 = ~w24077 & ~w24078;
assign w24080 = w9061 & ~w23366;
assign w24081 = w7489 & w21934;
assign w24082 = w7192 & ~w21940;
assign w24083 = w7511 & ~w21968;
assign w24084 = ~w24081 & ~w24082;
assign w24085 = w24084 & w37222;
assign w24086 = (~a_11 & ~w24084) | (~a_11 & w37223) | (~w24084 & w37223);
assign w24087 = ~w24085 & ~w24086;
assign w24088 = (w24087 & w23366) | (w24087 & w37224) | (w23366 & w37224);
assign w24089 = ~w24080 & ~w24088;
assign w24090 = w24079 & w24089;
assign w24091 = ~w24079 & ~w24089;
assign w24092 = ~w24090 & ~w24091;
assign w24093 = ~w23992 & w24092;
assign w24094 = ~w23981 & ~w23991;
assign w24095 = ~w24092 & ~w24094;
assign w24096 = ~w24093 & ~w24095;
assign w24097 = w23977 & ~w24096;
assign w24098 = w24092 & ~w24094;
assign w24099 = ~w23992 & ~w24092;
assign w24100 = ~w24098 & ~w24099;
assign w24101 = ~w23977 & ~w24100;
assign w24102 = ~w24097 & ~w24101;
assign w24103 = w23981 & w23991;
assign w24104 = w24092 & ~w24103;
assign w24105 = ~w23981 & w23991;
assign w24106 = ~w24092 & ~w24105;
assign w24107 = ~w24104 & ~w24106;
assign w24108 = ~w23977 & w24107;
assign w24109 = w24092 & ~w24105;
assign w24110 = ~w24092 & ~w24103;
assign w24111 = ~w24109 & ~w24110;
assign w24112 = w23977 & w24111;
assign w24113 = ~w24108 & ~w24112;
assign w24114 = ~w24102 & w24113;
assign w24115 = w9788 & ~w22020;
assign w24116 = w9786 & w22007;
assign w24117 = w9780 & w22014;
assign w24118 = (~w22002 & w37225) | (~w22002 & w37226) | (w37225 & w37226);
assign w24119 = ~w22021 & ~w22023;
assign w24120 = w24118 & ~w24119;
assign w24121 = ~w24118 & w24119;
assign w24122 = ~w24120 & ~w24121;
assign w24123 = ~w24116 & ~w24117;
assign w24124 = ~w24115 & w24123;
assign w24125 = (w24124 & ~w24122) | (w24124 & w37227) | (~w24122 & w37227);
assign w24126 = ~a_5 & w24125;
assign w24127 = (w24122 & w37228) | (w24122 & w37229) | (w37228 & w37229);
assign w24128 = ~w24126 & ~w24127;
assign w24129 = w24114 & ~w24128;
assign w24130 = ~w24114 & w24128;
assign w24131 = ~w24129 & ~w24130;
assign w24132 = w23972 & w24131;
assign w24133 = ~w23972 & ~w24131;
assign w24134 = ~w24132 & ~w24133;
assign w24135 = ~w23967 & w24134;
assign w24136 = w24128 & ~w24134;
assign w24137 = w23971 & w24113;
assign w24138 = ~w24102 & ~w24137;
assign w24139 = ~w23570 & ~w24102;
assign w24140 = w23394 & w24139;
assign w24141 = ~w24138 & ~w24140;
assign w24142 = ~w23981 & w24092;
assign w24143 = w23981 & ~w24092;
assign w24144 = ~w24142 & ~w24143;
assign w24145 = ~w23977 & ~w24144;
assign w24146 = (w24089 & ~w24079) | (w24089 & w37230) | (~w24079 & w37230);
assign w24147 = ~w24142 & w24146;
assign w24148 = ~w24145 & ~w24147;
assign w24149 = (~w23980 & ~w24067) | (~w23980 & w32547) | (~w24067 & w32547);
assign w24150 = ~w23979 & w24149;
assign w24151 = ~w24077 & ~w24150;
assign w24152 = w9061 & ~w22930;
assign w24153 = w7489 & ~w21968;
assign w24154 = w7192 & w21934;
assign w24155 = w7511 & ~w21973;
assign w24156 = ~w24153 & ~w24154;
assign w24157 = ~w24155 & w24156;
assign w24158 = ~a_11 & ~w24157;
assign w24159 = a_11 & w24157;
assign w24160 = ~w24158 & ~w24159;
assign w24161 = (w24160 & w22930) | (w24160 & w37231) | (w22930 & w37231);
assign w24162 = ~w24152 & ~w24161;
assign w24163 = ~w24062 & ~w24065;
assign w24164 = w6304 & w21921;
assign w24165 = w6059 & w21892;
assign w24166 = w6061 & ~w21910;
assign w24167 = ~w24164 & ~w24165;
assign w24168 = ~w24166 & w24167;
assign w24169 = (w24168 & ~w22664) | (w24168 & w37232) | (~w22664 & w37232);
assign w24170 = ~a_17 & w24169;
assign w24171 = (w22664 & w37233) | (w22664 & w37234) | (w37233 & w37234);
assign w24172 = ~w24170 & ~w24171;
assign w24173 = ~w23506 & ~w24056;
assign w24174 = ~w23511 & w24173;
assign w24175 = ~w24055 & ~w24174;
assign w24176 = w8311 & w22555;
assign w24177 = w5308 & w21787;
assign w24178 = ~w21882 & w37235;
assign w24179 = (~w24177 & ~w21901) | (~w24177 & w37236) | (~w21901 & w37236);
assign w24180 = ~w24178 & w24179;
assign w24181 = a_20 & w24180;
assign w24182 = ~a_20 & ~w24180;
assign w24183 = ~w24181 & ~w24182;
assign w24184 = (w24183 & ~w22555) | (w24183 & w37237) | (~w22555 & w37237);
assign w24185 = ~w24176 & ~w24184;
assign w24186 = w5017 & w22247;
assign w24187 = w5017 & ~w22246;
assign w24188 = w5016 & w21833;
assign w24189 = w5286 & w21854;
assign w24190 = (~w24188 & w21839) | (~w24188 & w37238) | (w21839 & w37238);
assign w24191 = ~w24189 & w24190;
assign w24192 = (w24191 & ~w24187) | (w24191 & w32147) | (~w24187 & w32147);
assign w24193 = ~w24186 & w24192;
assign w24194 = ~a_23 & w24193;
assign w24195 = a_23 & ~w24193;
assign w24196 = ~w24194 & ~w24195;
assign w24197 = w24019 & ~w24030;
assign w24198 = w24029 & w32148;
assign w24199 = ~w24031 & ~w24198;
assign w24200 = ~w24197 & w24199;
assign w24201 = w21815 & w35763;
assign w24202 = w4446 & w21813;
assign w24203 = w4070 & ~w21815;
assign w24204 = w21813 & w24203;
assign w24205 = w4070 & w21815;
assign w24206 = ~w21813 & w24205;
assign w24207 = ~w24204 & ~w24206;
assign w24208 = w4068 & w21815;
assign w24209 = (~w24208 & ~w21813) | (~w24208 & w37239) | (~w21813 & w37239);
assign w24210 = (w24201 & ~w24207) | (w24201 & w37240) | (~w24207 & w37240);
assign w24211 = w24207 & w37241;
assign w24212 = ~w24210 & ~w24211;
assign w24213 = w24200 & w24212;
assign w24214 = ~w24200 & ~w24212;
assign w24215 = ~w24213 & ~w24214;
assign w24216 = ~w22177 & w32149;
assign w24217 = (w1226 & w21819) | (w1226 & w32150) | (w21819 & w32150);
assign w24218 = w22177 & w24217;
assign w24219 = ~w518 & w21807;
assign w24220 = w4666 & ~w21803;
assign w24221 = ~w21796 & w37242;
assign w24222 = ~w24219 & ~w24221;
assign w24223 = ~w24220 & w24222;
assign w24224 = ~w24218 & w24223;
assign w24225 = (a_26 & ~w24224) | (a_26 & w32151) | (~w24224 & w32151);
assign w24226 = w24224 & w32152;
assign w24227 = ~w24225 & ~w24226;
assign w24228 = w24215 & w24227;
assign w24229 = ~w24215 & ~w24227;
assign w24230 = ~w24228 & ~w24229;
assign w24231 = w24196 & w24230;
assign w24232 = ~w24196 & ~w24230;
assign w24233 = ~w24231 & ~w24232;
assign w24234 = (~w24049 & ~w24018) | (~w24049 & w32153) | (~w24018 & w32153);
assign w24235 = w24233 & ~w24234;
assign w24236 = ~w24233 & w24234;
assign w24237 = ~w24235 & ~w24236;
assign w24238 = ~w24185 & ~w24237;
assign w24239 = w24185 & w24237;
assign w24240 = ~w24238 & ~w24239;
assign w24241 = w24175 & ~w24240;
assign w24242 = ~w24175 & w24240;
assign w24243 = ~w24241 & ~w24242;
assign w24244 = w24172 & w24243;
assign w24245 = ~w24172 & ~w24243;
assign w24246 = ~w24244 & ~w24245;
assign w24247 = w6998 & ~w21945;
assign w24248 = w6446 & w21951;
assign w24249 = w6996 & ~w21940;
assign w24250 = ~w24247 & ~w24248;
assign w24251 = ~w24249 & w24250;
assign w24252 = (w24251 & ~w23032) | (w24251 & w37243) | (~w23032 & w37243);
assign w24253 = a_14 & w24252;
assign w24254 = (w23032 & w37244) | (w23032 & w37245) | (w37244 & w37245);
assign w24255 = ~w24253 & ~w24254;
assign w24256 = w24246 & ~w24255;
assign w24257 = ~w24246 & w24255;
assign w24258 = ~w24256 & ~w24257;
assign w24259 = w24163 & ~w24258;
assign w24260 = ~w24163 & w24258;
assign w24261 = ~w24259 & ~w24260;
assign w24262 = w24162 & ~w24261;
assign w24263 = w24151 & w24262;
assign w24264 = w24162 & w24261;
assign w24265 = ~w24151 & w24264;
assign w24266 = ~w24263 & ~w24265;
assign w24267 = ~w24162 & w24261;
assign w24268 = w24151 & w24267;
assign w24269 = ~w24162 & ~w24261;
assign w24270 = ~w24151 & w24269;
assign w24271 = ~w24268 & ~w24270;
assign w24272 = w24266 & w24271;
assign w24273 = w9456 & w23580;
assign w24274 = w8298 & ~w21992;
assign w24275 = w8277 & w21985;
assign w24276 = w8295 & w22007;
assign w24277 = ~w24274 & ~w24275;
assign w24278 = w24277 & w37246;
assign w24279 = (~a_8 & ~w24277) | (~a_8 & w37247) | (~w24277 & w37247);
assign w24280 = ~w24278 & ~w24279;
assign w24281 = (w24280 & ~w23580) | (w24280 & w37248) | (~w23580 & w37248);
assign w24282 = ~w24273 & ~w24281;
assign w24283 = w24272 & ~w24282;
assign w24284 = ~w24272 & w24282;
assign w24285 = ~w24283 & ~w24284;
assign w24286 = w24148 & w24285;
assign w24287 = ~w24148 & ~w24285;
assign w24288 = ~w24286 & ~w24287;
assign w24289 = ~w24141 & w24288;
assign w24290 = w24141 & ~w24288;
assign w24291 = ~w24289 & ~w24290;
assign w24292 = ~w21774 & ~w22025;
assign w24293 = ~w22022 & w37249;
assign w24294 = (w24292 & w22022) | (w24292 & w37250) | (w22022 & w37250);
assign w24295 = ~w24293 & ~w24294;
assign w24296 = w10033 & w24295;
assign w24297 = w9780 & ~w22020;
assign w24298 = w9786 & w22014;
assign w24299 = w9788 & w21771;
assign w24300 = ~w24297 & ~w24298;
assign w24301 = w24300 & w37251;
assign w24302 = (~a_5 & ~w24300) | (~a_5 & w37252) | (~w24300 & w37252);
assign w24303 = ~w24301 & ~w24302;
assign w24304 = (w24303 & ~w24295) | (w24303 & w37253) | (~w24295 & w37253);
assign w24305 = ~w24296 & ~w24304;
assign w24306 = w24291 & w24305;
assign w24307 = ~w24136 & ~w24306;
assign w24308 = ~w24135 & w24307;
assign w24309 = ~w24291 & ~w24305;
assign w24310 = ~w24148 & ~w24272;
assign w24311 = w24148 & w24272;
assign w24312 = ~w24310 & ~w24311;
assign w24313 = w24282 & ~w24312;
assign w24314 = ~w24289 & ~w24313;
assign w24315 = ~w24147 & w24266;
assign w24316 = ~w24145 & w24315;
assign w24317 = ~w24163 & w24256;
assign w24318 = ~w24246 & ~w24255;
assign w24319 = w24163 & w24318;
assign w24320 = ~w24317 & ~w24319;
assign w24321 = w24261 & w24320;
assign w24322 = ~w24077 & w24320;
assign w24323 = ~w24150 & w24322;
assign w24324 = ~w24321 & ~w24323;
assign w24325 = ~w24062 & ~w24245;
assign w24326 = ~w24065 & w24325;
assign w24327 = ~w24244 & ~w24326;
assign w24328 = ~w23551 & w37254;
assign w24329 = ~w23551 & w37255;
assign w24330 = w7511 & w21985;
assign w24331 = w7192 & ~w21968;
assign w24332 = w7489 & ~w21973;
assign w24333 = ~w24330 & ~w24331;
assign w24334 = w24333 & w37256;
assign w24335 = (~a_11 & ~w24333) | (~a_11 & w37257) | (~w24333 & w37257);
assign w24336 = ~w24334 & ~w24335;
assign w24337 = ~w24329 & w24336;
assign w24338 = ~w24328 & ~w24337;
assign w24339 = (~w24338 & w24326) | (~w24338 & w32548) | (w24326 & w32548);
assign w24340 = ~w24326 & w32549;
assign w24341 = ~w24339 & ~w24340;
assign w24342 = w24175 & ~w24239;
assign w24343 = (~w24238 & ~w24175) | (~w24238 & w32550) | (~w24175 & w32550);
assign w24344 = w5017 & w22107;
assign w24345 = w21873 & w32154;
assign w24346 = w5017 & ~w21854;
assign w24347 = ~w21787 & w24346;
assign w24348 = ~w24345 & ~w24347;
assign w24349 = ~w22105 & ~w24348;
assign w24350 = w5016 & ~w21839;
assign w24351 = w5080 & w21854;
assign w24352 = w5286 & w21787;
assign w24353 = ~w24350 & ~w24351;
assign w24354 = ~w24352 & w24353;
assign w24355 = ~w24349 & w24354;
assign w24356 = ~w24344 & w24355;
assign w24357 = a_23 & ~w24356;
assign w24358 = ~a_23 & w24356;
assign w24359 = ~w24357 & ~w24358;
assign w24360 = w4403 & w22289;
assign w24361 = w4403 & w21830;
assign w24362 = w21824 & w24361;
assign w24363 = w4666 & ~w21224;
assign w24364 = w21207 & w24363;
assign w24365 = w4666 & w21224;
assign w24366 = ~w21207 & w24365;
assign w24367 = ~w24364 & ~w24366;
assign w24368 = (~w518 & ~w21156) | (~w518 & w32155) | (~w21156 & w32155);
assign w24369 = ~w21796 & w24368;
assign w24370 = w4638 & ~w21800;
assign w24371 = w21799 & w24370;
assign w24372 = w4638 & w21800;
assign w24373 = ~w21799 & w24372;
assign w24374 = ~w24371 & ~w24373;
assign w24375 = ~w24369 & w24374;
assign w24376 = w24367 & w24375;
assign w24377 = w7680 & w24376;
assign w24378 = a_26 & ~w24376;
assign w24379 = ~w24377 & ~w24378;
assign w24380 = ~w24362 & w24379;
assign w24381 = ~w24360 & w24380;
assign w24382 = (~a_26 & w21796) | (~a_26 & w32156) | (w21796 & w32156);
assign w24383 = w24374 & w24382;
assign w24384 = w24367 & w24383;
assign w24385 = ~w21830 & w24384;
assign w24386 = w21824 & w24385;
assign w24387 = w21830 & w24384;
assign w24388 = ~w21824 & w24387;
assign w24389 = ~w24386 & ~w24388;
assign w24390 = (a_29 & ~w21815) | (a_29 & w37258) | (~w21815 & w37258);
assign w24391 = ~w24202 & w24390;
assign w24392 = w24207 & w24391;
assign w24393 = a_29 & ~w24392;
assign w24394 = w4070 & ~w22161;
assign w24395 = w4446 & w21807;
assign w24396 = w3957 & w21815;
assign w24397 = (~w24396 & ~w21813) | (~w24396 & w32157) | (~w21813 & w32157);
assign w24398 = ~w24395 & w24397;
assign w24399 = ~w24394 & w24398;
assign w24400 = ~w24393 & w24399;
assign w24401 = w24393 & ~w24399;
assign w24402 = ~w24400 & ~w24401;
assign w24403 = (~w24402 & ~w24381) | (~w24402 & w32551) | (~w24381 & w32551);
assign w24404 = w24389 & w24402;
assign w24405 = w24381 & w24404;
assign w24406 = ~w24403 & ~w24405;
assign w24407 = ~w24214 & w24227;
assign w24408 = ~w24213 & ~w24407;
assign w24409 = ~w24406 & w24408;
assign w24410 = w24406 & ~w24408;
assign w24411 = ~w24409 & ~w24410;
assign w24412 = w24359 & w24411;
assign w24413 = ~w24359 & ~w24411;
assign w24414 = ~w24412 & ~w24413;
assign w24415 = ~w24232 & ~w24234;
assign w24416 = ~w24231 & ~w24415;
assign w24417 = w24414 & w24416;
assign w24418 = ~w24414 & ~w24416;
assign w24419 = ~w24417 & ~w24418;
assign w24420 = w5816 & w21892;
assign w24421 = w5818 & w21901;
assign w24422 = ~w21882 & w37259;
assign w24423 = ~w24420 & ~w24421;
assign w24424 = ~w24422 & w24423;
assign w24425 = (w22096 & w32552) | (w22096 & w32553) | (w32552 & w32553);
assign w24426 = (~w22096 & w32554) | (~w22096 & w32555) | (w32554 & w32555);
assign w24427 = ~w24425 & ~w24426;
assign w24428 = ~w24419 & w24427;
assign w24429 = w24419 & ~w24427;
assign w24430 = ~w24428 & ~w24429;
assign w24431 = ~w22901 & w37260;
assign w24432 = ~w22901 & w32159;
assign w24433 = w6059 & ~w21910;
assign w24434 = w6304 & w21951;
assign w24435 = w6061 & w21921;
assign w24436 = ~w24434 & w37261;
assign w24437 = ~a_17 & ~w24436;
assign w24438 = a_17 & w24436;
assign w24439 = ~w24437 & ~w24438;
assign w24440 = ~w24432 & w24439;
assign w24441 = ~w24431 & ~w24440;
assign w24442 = w24430 & ~w24441;
assign w24443 = w24343 & w24442;
assign w24444 = ~w24430 & ~w24441;
assign w24445 = ~w24343 & w24444;
assign w24446 = ~w24443 & ~w24445;
assign w24447 = ~w24430 & w24441;
assign w24448 = w24343 & w24447;
assign w24449 = w24430 & w24441;
assign w24450 = ~w24343 & w24449;
assign w24451 = ~w24448 & ~w24450;
assign w24452 = w24446 & w24451;
assign w24453 = w6446 & ~w21945;
assign w24454 = w6996 & w21934;
assign w24455 = w6998 & ~w21940;
assign w24456 = ~w24453 & ~w24454;
assign w24457 = (a_14 & ~w24456) | (a_14 & w37262) | (~w24456 & w37262);
assign w24458 = w6447 & w23310;
assign w24459 = w24456 & w37263;
assign w24460 = ~w24458 & w24459;
assign w24461 = (~w24457 & ~w23310) | (~w24457 & w37264) | (~w23310 & w37264);
assign w24462 = ~w24460 & w24461;
assign w24463 = w24452 & ~w24462;
assign w24464 = ~w24452 & w24462;
assign w24465 = ~w24463 & ~w24464;
assign w24466 = w24341 & ~w24465;
assign w24467 = ~w24341 & w24465;
assign w24468 = ~w24466 & ~w24467;
assign w24469 = w24324 & w24468;
assign w24470 = ~w24324 & ~w24468;
assign w24471 = ~w24469 & ~w24470;
assign w24472 = w24271 & ~w24471;
assign w24473 = ~w24316 & w24472;
assign w24474 = ~w23397 & w37265;
assign w24475 = ~w23397 & w37266;
assign w24476 = w8298 & w22007;
assign w24477 = w8277 & ~w21992;
assign w24478 = w8295 & w22014;
assign w24479 = ~w24476 & ~w24477;
assign w24480 = ~w24478 & w24479;
assign w24481 = ~a_8 & ~w24480;
assign w24482 = a_8 & w24480;
assign w24483 = ~w24481 & ~w24482;
assign w24484 = ~w24475 & w24483;
assign w24485 = ~w24474 & ~w24484;
assign w24486 = w24473 & ~w24485;
assign w24487 = w24271 & ~w24316;
assign w24488 = w24471 & ~w24485;
assign w24489 = ~w24487 & w24488;
assign w24490 = ~w24486 & ~w24489;
assign w24491 = w24471 & w24485;
assign w24492 = w24487 & w24491;
assign w24493 = ~w24471 & w24485;
assign w24494 = ~w24487 & w24493;
assign w24495 = ~w24492 & ~w24494;
assign w24496 = w24490 & w24495;
assign w24497 = ~w22022 & w37267;
assign w24498 = ~w24497 & w37268;
assign w24499 = ~w21772 & ~w22026;
assign w24500 = ~w22025 & ~w24499;
assign w24501 = (~w22022 & w37269) | (~w22022 & w37270) | (w37269 & w37270);
assign w24502 = ~w24498 & ~w24501;
assign w24503 = ~w24498 & w37271;
assign w24504 = ~w24498 & w37272;
assign w24505 = w9786 & ~w22020;
assign w24506 = ~w21760 & w37273;
assign w24507 = w9780 & w21771;
assign w24508 = ~w24505 & ~w24506;
assign w24509 = w24508 & w37274;
assign w24510 = (~a_5 & ~w24508) | (~a_5 & w37275) | (~w24508 & w37275);
assign w24511 = ~w24509 & ~w24510;
assign w24512 = ~w24504 & w24511;
assign w24513 = ~w24503 & ~w24512;
assign w24514 = ~w24496 & ~w24513;
assign w24515 = w24314 & w24514;
assign w24516 = w24496 & ~w24513;
assign w24517 = ~w24314 & w24516;
assign w24518 = ~w24515 & ~w24517;
assign w24519 = ~w24309 & w24518;
assign w24520 = ~w24308 & w24519;
assign w24521 = ~w24313 & w24495;
assign w24522 = ~w24289 & w24521;
assign w24523 = w24490 & ~w24522;
assign w24524 = w9786 & w21771;
assign w24525 = w9788 & ~w22035;
assign w24526 = ~w21760 & w37276;
assign w24527 = ~w24497 & w37277;
assign w24528 = (~w21780 & w24497) | (~w21780 & w37278) | (w24497 & w37278);
assign w24529 = ~w24527 & ~w24528;
assign w24530 = ~w24525 & ~w24526;
assign w24531 = ~w24524 & w24530;
assign w24532 = (w24531 & ~w24529) | (w24531 & w37279) | (~w24529 & w37279);
assign w24533 = a_5 & ~w24532;
assign w24534 = (~w24529 & w37280) | (~w24529 & w37281) | (w37280 & w37281);
assign w24535 = ~w24533 & ~w24534;
assign w24536 = ~w24327 & w24463;
assign w24537 = ~w24452 & ~w24462;
assign w24538 = w24327 & w24537;
assign w24539 = ~w24536 & ~w24538;
assign w24540 = ~w24327 & w24464;
assign w24541 = w24452 & w24462;
assign w24542 = w24327 & w24541;
assign w24543 = ~w24540 & ~w24542;
assign w24544 = w24539 & w24543;
assign w24545 = w24324 & ~w24544;
assign w24546 = ~w24324 & w24544;
assign w24547 = ~w24545 & ~w24546;
assign w24548 = w24338 & ~w24547;
assign w24549 = ~w24473 & ~w24548;
assign w24550 = ~w24261 & w24539;
assign w24551 = ~w24151 & w24550;
assign w24552 = w24320 & w24543;
assign w24553 = w24539 & ~w24552;
assign w24554 = ~w24551 & ~w24553;
assign w24555 = w9061 & ~w23930;
assign w24556 = w7489 & w21985;
assign w24557 = w7192 & ~w21973;
assign w24558 = w7511 & ~w21992;
assign w24559 = ~w24556 & ~w24557;
assign w24560 = w24559 & w37282;
assign w24561 = (~a_11 & ~w24559) | (~a_11 & w37283) | (~w24559 & w37283);
assign w24562 = ~w24560 & ~w24561;
assign w24563 = (w24562 & w23930) | (w24562 & w37284) | (w23930 & w37284);
assign w24564 = ~w24555 & ~w24563;
assign w24565 = ~w24326 & w37285;
assign w24566 = w24446 & ~w24565;
assign w24567 = w8564 & ~w23366;
assign w24568 = w6446 & ~w21940;
assign w24569 = w6998 & w21934;
assign w24570 = w6996 & ~w21968;
assign w24571 = ~w24568 & ~w24569;
assign w24572 = w24571 & w37286;
assign w24573 = (~a_14 & ~w24571) | (~a_14 & w37287) | (~w24571 & w37287);
assign w24574 = ~w24572 & ~w24573;
assign w24575 = (w24574 & w23366) | (w24574 & w37288) | (w23366 & w37288);
assign w24576 = ~w24567 & ~w24575;
assign w24577 = ~w24238 & ~w24429;
assign w24578 = ~w24342 & w24577;
assign w24579 = ~w24428 & ~w24578;
assign w24580 = ~w24413 & ~w24417;
assign w24581 = ~w21882 & w32161;
assign w24582 = ~w22381 & w24581;
assign w24583 = ~w21882 & w32162;
assign w24584 = w5080 & w21787;
assign w24585 = w5016 & w21854;
assign w24586 = ~w24584 & ~w24585;
assign w24587 = ~w24583 & w24586;
assign w24588 = ~w24582 & w24587;
assign w24589 = w24588 & w32163;
assign w24590 = (a_23 & ~w24588) | (a_23 & w32164) | (~w24588 & w32164);
assign w24591 = ~w24589 & ~w24590;
assign w24592 = ~w24213 & ~w24405;
assign w24593 = (~w24403 & ~w24592) | (~w24403 & w32556) | (~w24592 & w32556);
assign w24594 = ~w21796 & w32165;
assign w24595 = w3957 & w21813;
assign w24596 = w4068 & w21807;
assign w24597 = ~w24595 & ~w24596;
assign w24598 = ~w24594 & w24597;
assign w24599 = ~w21817 & w32166;
assign w24600 = ~w22137 & w24599;
assign w24601 = ~w21820 & w32167;
assign w24602 = w21819 & w24601;
assign w24603 = ~w24600 & ~w24602;
assign w24604 = (a_29 & ~w24603) | (a_29 & w32168) | (~w24603 & w32168);
assign w24605 = ~a_29 & w24598;
assign w24606 = w24603 & w24605;
assign w24607 = ~w1477 & w21815;
assign w24608 = w24392 & w24398;
assign w24609 = ~w24394 & w24608;
assign w24610 = w24607 & w24609;
assign w24611 = ~w24607 & ~w24609;
assign w24612 = ~w24610 & ~w24611;
assign w24613 = ~w24606 & w24612;
assign w24614 = ~w24604 & w24613;
assign w24615 = ~w24604 & ~w24606;
assign w24616 = ~w24612 & ~w24615;
assign w24617 = ~w24614 & ~w24616;
assign w24618 = w4666 & ~w21237;
assign w24619 = ~w21231 & w24618;
assign w24620 = ~w518 & ~w21803;
assign w24621 = w4638 & w21833;
assign w24622 = w21836 & w37289;
assign w24623 = ~w24619 & ~w24620;
assign w24624 = ~w24621 & ~w24622;
assign w24625 = (a_26 & ~w24624) | (a_26 & w32169) | (~w24624 & w32169);
assign w24626 = w24624 & w32557;
assign w24627 = ~w24625 & ~w24626;
assign w24628 = ~w22278 & ~w24627;
assign w24629 = w24624 & w32558;
assign w24630 = (~w32169 & w32424) | (~w32169 & w37290) | (w32424 & w37290);
assign w24631 = ~w24629 & w24630;
assign w24632 = w22278 & ~w24631;
assign w24633 = ~w24628 & ~w24632;
assign w24634 = w24617 & w24633;
assign w24635 = ~w24617 & ~w24633;
assign w24636 = ~w24634 & ~w24635;
assign w24637 = w24593 & ~w24636;
assign w24638 = ~w24593 & w24636;
assign w24639 = ~w24637 & ~w24638;
assign w24640 = w24591 & ~w24639;
assign w24641 = ~w24591 & w24639;
assign w24642 = ~w24640 & ~w24641;
assign w24643 = w8339 & ~w22577;
assign w24644 = (~w21896 & w37291) | (~w21896 & w37292) | (w37291 & w37292);
assign w24645 = w8339 & ~w21914;
assign w24646 = w22577 & w24645;
assign w24647 = (w24646 & w21896) | (w24646 & w37293) | (w21896 & w37293);
assign w24648 = w5816 & ~w21910;
assign w24649 = w5308 & w21901;
assign w24650 = w5818 & w21892;
assign w24651 = ~w24649 & ~w24650;
assign w24652 = w24651 & w37294;
assign w24653 = (a_20 & ~w24651) | (a_20 & w37295) | (~w24651 & w37295);
assign w24654 = ~w24652 & ~w24653;
assign w24655 = ~w24647 & ~w24654;
assign w24656 = ~w24644 & w24655;
assign w24657 = w8311 & w22577;
assign w24658 = (w21896 & w37296) | (w21896 & w37297) | (w37296 & w37297);
assign w24659 = w8311 & ~w22577;
assign w24660 = (~w21896 & w37298) | (~w21896 & w37299) | (w37298 & w37299);
assign w24661 = ~w24658 & ~w24660;
assign w24662 = ~w24656 & w24661;
assign w24663 = w24642 & ~w24662;
assign w24664 = w24580 & w24663;
assign w24665 = ~w24642 & ~w24662;
assign w24666 = ~w24580 & w24665;
assign w24667 = ~w24664 & ~w24666;
assign w24668 = ~w24642 & w24662;
assign w24669 = w24580 & w24668;
assign w24670 = w24642 & w24662;
assign w24671 = ~w24580 & w24670;
assign w24672 = ~w24669 & ~w24671;
assign w24673 = w24667 & w24672;
assign w24674 = w6061 & w21951;
assign w24675 = w6059 & w21921;
assign w24676 = w6304 & ~w21945;
assign w24677 = ~w24674 & ~w24675;
assign w24678 = ~w24676 & w24677;
assign w24679 = (~w22083 & w37300) | (~w22083 & w37301) | (w37300 & w37301);
assign w24680 = (w22083 & w37302) | (w22083 & w37303) | (w37302 & w37303);
assign w24681 = ~w24679 & ~w24680;
assign w24682 = w24673 & ~w24681;
assign w24683 = ~w24673 & w24681;
assign w24684 = ~w24682 & ~w24683;
assign w24685 = w24579 & w24684;
assign w24686 = ~w24579 & ~w24684;
assign w24687 = ~w24685 & ~w24686;
assign w24688 = w24576 & ~w24687;
assign w24689 = ~w24576 & w24687;
assign w24690 = ~w24688 & ~w24689;
assign w24691 = w24566 & w24690;
assign w24692 = ~w24566 & ~w24690;
assign w24693 = ~w24691 & ~w24692;
assign w24694 = w24564 & ~w24693;
assign w24695 = w24554 & w24694;
assign w24696 = w24564 & w24693;
assign w24697 = ~w24554 & w24696;
assign w24698 = ~w24695 & ~w24697;
assign w24699 = ~w24564 & w24693;
assign w24700 = w24554 & w24699;
assign w24701 = ~w24564 & ~w24693;
assign w24702 = ~w24554 & w24701;
assign w24703 = ~w24700 & ~w24702;
assign w24704 = w24698 & w24703;
assign w24705 = w9456 & w24122;
assign w24706 = w8298 & w22014;
assign w24707 = w8277 & w22007;
assign w24708 = w8295 & ~w22020;
assign w24709 = ~w24706 & ~w24707;
assign w24710 = w24709 & w37304;
assign w24711 = (~a_8 & ~w24709) | (~a_8 & w37305) | (~w24709 & w37305);
assign w24712 = ~w24710 & ~w24711;
assign w24713 = (w24712 & ~w24122) | (w24712 & w37306) | (~w24122 & w37306);
assign w24714 = ~w24705 & ~w24713;
assign w24715 = ~w24704 & w24714;
assign w24716 = w24704 & ~w24714;
assign w24717 = ~w24715 & ~w24716;
assign w24718 = w24549 & w24717;
assign w24719 = ~w24549 & ~w24717;
assign w24720 = ~w24718 & ~w24719;
assign w24721 = w24535 & ~w24720;
assign w24722 = w24523 & w24721;
assign w24723 = w24535 & w24720;
assign w24724 = ~w24523 & w24723;
assign w24725 = ~w24722 & ~w24724;
assign w24726 = ~w24314 & ~w24496;
assign w24727 = w24314 & w24496;
assign w24728 = ~w24726 & ~w24727;
assign w24729 = w24513 & ~w24728;
assign w24730 = w24725 & ~w24729;
assign w24731 = ~w24520 & w24730;
assign w24732 = w24523 & w24720;
assign w24733 = ~w24549 & w24715;
assign w24734 = w24704 & w24714;
assign w24735 = w24549 & w24734;
assign w24736 = ~w24733 & ~w24735;
assign w24737 = ~w24548 & w24698;
assign w24738 = ~w24473 & w24737;
assign w24739 = (w24703 & ~w24737) | (w24703 & w32171) | (~w24737 & w32171);
assign w24740 = ~w24554 & ~w24693;
assign w24741 = w24576 & w24693;
assign w24742 = ~w24740 & ~w24741;
assign w24743 = w9456 & w24295;
assign w24744 = w8298 & ~w22020;
assign w24745 = w8277 & w22014;
assign w24746 = w8295 & w21771;
assign w24747 = ~w24744 & ~w24745;
assign w24748 = w24747 & w37307;
assign w24749 = (~a_8 & ~w24747) | (~a_8 & w37308) | (~w24747 & w37308);
assign w24750 = ~w24748 & ~w24749;
assign w24751 = (w24750 & ~w24295) | (w24750 & w37309) | (~w24295 & w37309);
assign w24752 = ~w24743 & ~w24751;
assign w24753 = ~w22036 & ~w22043;
assign w24754 = (w22022 & w37310) | (w22022 & w37311) | (w37310 & w37311);
assign w24755 = (~w22022 & w37312) | (~w22022 & w37313) | (w37312 & w37313);
assign w24756 = ~w24754 & ~w24755;
assign w24757 = w10033 & w24756;
assign w24758 = ~w21760 & w37314;
assign w24759 = w9780 & ~w22035;
assign w24760 = w9788 & w22032;
assign w24761 = ~w24758 & ~w24759;
assign w24762 = (~a_5 & ~w24761) | (~a_5 & w37315) | (~w24761 & w37315);
assign w24763 = w24761 & w37316;
assign w24764 = ~w24762 & ~w24763;
assign w24765 = (w24764 & ~w24756) | (w24764 & w37317) | (~w24756 & w37317);
assign w24766 = ~w24757 & ~w24765;
assign w24767 = w24752 & ~w24766;
assign w24768 = ~w24752 & w24766;
assign w24769 = ~w24767 & ~w24768;
assign w24770 = w24681 & ~w24687;
assign w24771 = w24446 & w24687;
assign w24772 = ~w24565 & w24771;
assign w24773 = ~w24770 & ~w24772;
assign w24774 = ~w24428 & w24672;
assign w24775 = (w24667 & ~w24774) | (w24667 & w32172) | (~w24774 & w32172);
assign w24776 = ~w24413 & ~w24641;
assign w24777 = ~w24417 & w24776;
assign w24778 = ~w24640 & ~w24777;
assign w24779 = w5016 & w21787;
assign w24780 = ~w21882 & w37318;
assign w24781 = (~w24779 & ~w21901) | (~w24779 & w37319) | (~w21901 & w37319);
assign w24782 = ~w24780 & w24781;
assign w24783 = a_23 & ~w24782;
assign w24784 = ~a_23 & w24782;
assign w24785 = (w24784 & ~w22555) | (w24784 & w32559) | (~w22555 & w32559);
assign w24786 = (~w24783 & ~w22555) | (~w24783 & w32635) | (~w22555 & w32635);
assign w24787 = ~w24785 & w24786;
assign w24788 = w1226 & w22247;
assign w24789 = w1226 & ~w22246;
assign w24790 = ~w518 & w21833;
assign w24791 = w4666 & w21854;
assign w24792 = (~w24790 & w21839) | (~w24790 & w37320) | (w21839 & w37320);
assign w24793 = ~w24791 & w24792;
assign w24794 = (w24793 & ~w24789) | (w24793 & w32173) | (~w24789 & w32173);
assign w24795 = ~w24788 & w24794;
assign w24796 = ~a_26 & w24795;
assign w24797 = a_26 & ~w24795;
assign w24798 = ~w24796 & ~w24797;
assign w24799 = (~w24610 & ~w24613) | (~w24610 & w32174) | (~w24613 & w32174);
assign w24800 = ~w21813 & w32175;
assign w24801 = w1327 & w21815;
assign w24802 = (~w1477 & ~w21815) | (~w1477 & w32176) | (~w21815 & w32176);
assign w24803 = (~w24801 & ~w21813) | (~w24801 & w32177) | (~w21813 & w32177);
assign w24804 = ~w24800 & w24803;
assign w24805 = w87 & w37321;
assign w24806 = w1125 & w1152;
assign w24807 = w1287 & w1949;
assign w24808 = w2418 & w3560;
assign w24809 = w3892 & w4152;
assign w24810 = w4539 & ~w24805;
assign w24811 = w24809 & w24810;
assign w24812 = w24807 & w24808;
assign w24813 = w2556 & w24806;
assign w24814 = w4711 & w24813;
assign w24815 = w24811 & w24812;
assign w24816 = w13728 & w24815;
assign w24817 = w24814 & w24816;
assign w24818 = ~w191 & ~w319;
assign w24819 = w648 & w24818;
assign w24820 = w1686 & w1777;
assign w24821 = w1821 & w2379;
assign w24822 = w5188 & w24821;
assign w24823 = w24819 & w24820;
assign w24824 = w729 & w24823;
assign w24825 = w24822 & w24824;
assign w24826 = ~w75 & ~w349;
assign w24827 = ~w355 & w24826;
assign w24828 = w51 & w2609;
assign w24829 = w3568 & w5387;
assign w24830 = w24828 & w24829;
assign w24831 = w2311 & w24827;
assign w24832 = w3064 & w6606;
assign w24833 = w24831 & w24832;
assign w24834 = w2181 & w24830;
assign w24835 = w15244 & w24834;
assign w24836 = w24833 & w24835;
assign w24837 = w24825 & w24836;
assign w24838 = w15174 & w24817;
assign w24839 = w24837 & w24838;
assign w24840 = ~w24804 & ~w24839;
assign w24841 = w24804 & w24839;
assign w24842 = ~w24840 & ~w24841;
assign w24843 = w24799 & ~w24842;
assign w24844 = ~w24799 & w24842;
assign w24845 = ~w24843 & ~w24844;
assign w24846 = (w4070 & w21819) | (w4070 & w32179) | (w21819 & w32179);
assign w24847 = w22177 & w24846;
assign w24848 = ~w21796 & w37322;
assign w24849 = w4446 & ~w21803;
assign w24850 = w3957 & w21807;
assign w24851 = ~w24848 & ~w24850;
assign w24852 = ~w24849 & w24851;
assign w24853 = ~w24847 & w24852;
assign w24854 = w24853 & w32180;
assign w24855 = (a_29 & ~w24853) | (a_29 & w32181) | (~w24853 & w32181);
assign w24856 = ~w24854 & ~w24855;
assign w24857 = w24845 & ~w24856;
assign w24858 = ~w24845 & w24856;
assign w24859 = ~w24857 & ~w24858;
assign w24860 = w24798 & ~w24859;
assign w24861 = ~w24798 & w24859;
assign w24862 = ~w24860 & ~w24861;
assign w24863 = (~w24635 & w24593) | (~w24635 & w32182) | (w24593 & w32182);
assign w24864 = w24862 & w24863;
assign w24865 = ~w24862 & ~w24863;
assign w24866 = ~w24864 & ~w24865;
assign w24867 = ~w24787 & ~w24866;
assign w24868 = w24787 & w24866;
assign w24869 = ~w24867 & ~w24868;
assign w24870 = w24778 & ~w24869;
assign w24871 = ~w24778 & w24869;
assign w24872 = ~w24870 & ~w24871;
assign w24873 = w5816 & w21921;
assign w24874 = w5308 & w21892;
assign w24875 = w5818 & ~w21910;
assign w24876 = ~w24873 & ~w24874;
assign w24877 = ~w24875 & w24876;
assign w24878 = (w24877 & ~w22664) | (w24877 & w37323) | (~w22664 & w37323);
assign w24879 = a_20 & w24878;
assign w24880 = (w22664 & w37324) | (w22664 & w37325) | (w37324 & w37325);
assign w24881 = ~w24879 & ~w24880;
assign w24882 = w24872 & ~w24881;
assign w24883 = ~w24872 & w24881;
assign w24884 = ~w24882 & ~w24883;
assign w24885 = w24775 & w24884;
assign w24886 = ~w24775 & ~w24884;
assign w24887 = ~w24885 & ~w24886;
assign w24888 = w9061 & w23580;
assign w24889 = w7489 & ~w21992;
assign w24890 = w7192 & w21985;
assign w24891 = w7511 & w22007;
assign w24892 = ~w24889 & ~w24890;
assign w24893 = (~a_11 & ~w24892) | (~a_11 & w37326) | (~w24892 & w37326);
assign w24894 = w24892 & w37327;
assign w24895 = ~w24893 & ~w24894;
assign w24896 = (w24895 & ~w23580) | (w24895 & w37328) | (~w23580 & w37328);
assign w24897 = ~w24888 & ~w24896;
assign w24898 = w8564 & ~w22930;
assign w24899 = w8592 & w22928;
assign w24900 = ~w22923 & w37329;
assign w24901 = ~w21959 & w37330;
assign w24902 = w6998 & ~w21968;
assign w24903 = w6446 & w21934;
assign w24904 = w6996 & ~w21973;
assign w24905 = ~w24902 & ~w24903;
assign w24906 = ~w24904 & w24905;
assign w24907 = a_14 & ~w24906;
assign w24908 = ~a_14 & w24906;
assign w24909 = ~w24907 & ~w24908;
assign w24910 = ~w24901 & ~w24909;
assign w24911 = ~w24899 & w24910;
assign w24912 = ~w24898 & ~w24911;
assign w24913 = w6061 & ~w21945;
assign w24914 = w6059 & w21951;
assign w24915 = w6304 & ~w21940;
assign w24916 = ~w24913 & ~w24914;
assign w24917 = ~w24915 & w24916;
assign w24918 = (w24917 & ~w23032) | (w24917 & w37331) | (~w23032 & w37331);
assign w24919 = ~a_17 & w24918;
assign w24920 = (w23032 & w37332) | (w23032 & w37333) | (w37332 & w37333);
assign w24921 = ~w24919 & ~w24920;
assign w24922 = w24912 & ~w24921;
assign w24923 = ~w24912 & w24921;
assign w24924 = ~w24922 & ~w24923;
assign w24925 = w24897 & ~w24924;
assign w24926 = ~w24897 & w24924;
assign w24927 = ~w24925 & ~w24926;
assign w24928 = w24887 & ~w24927;
assign w24929 = ~w24887 & w24927;
assign w24930 = ~w24928 & ~w24929;
assign w24931 = ~w24772 & w32560;
assign w24932 = (~w24930 & w24772) | (~w24930 & w32561) | (w24772 & w32561);
assign w24933 = ~w24931 & ~w24932;
assign w24934 = w24769 & ~w24933;
assign w24935 = ~w24769 & w24933;
assign w24936 = ~w24934 & ~w24935;
assign w24937 = w24742 & ~w24936;
assign w24938 = ~w24742 & w24936;
assign w24939 = ~w24937 & ~w24938;
assign w24940 = w24739 & w24939;
assign w24941 = ~w24739 & ~w24939;
assign w24942 = ~w24940 & ~w24941;
assign w24943 = w24736 & ~w24942;
assign w24944 = ~w24732 & w24943;
assign w24945 = w24720 & w24942;
assign w24946 = ~w24736 & w24942;
assign w24947 = (~w24946 & ~w24945) | (~w24946 & w32183) | (~w24945 & w32183);
assign w24948 = ~w24944 & w24947;
assign w24949 = ~w24523 & ~w24720;
assign w24950 = ~w24732 & ~w24949;
assign w24951 = ~w24535 & ~w24950;
assign w24952 = w24948 & ~w24951;
assign w24953 = ~w24731 & w24952;
assign w24954 = w24766 & ~w24948;
assign w24955 = w9788 & w22039;
assign w24956 = w9786 & ~w22035;
assign w24957 = w9780 & w22032;
assign w24958 = ~w22042 & w37334;
assign w24959 = ~w22040 & ~w22044;
assign w24960 = ~w22036 & ~w24959;
assign w24961 = ~w24754 & w24960;
assign w24962 = ~w24958 & ~w24961;
assign w24963 = ~w24956 & ~w24957;
assign w24964 = ~w24955 & w24963;
assign w24965 = (w24964 & ~w24962) | (w24964 & w37335) | (~w24962 & w37335);
assign w24966 = ~a_5 & w24965;
assign w24967 = (w24962 & w37336) | (w24962 & w37337) | (w37336 & w37337);
assign w24968 = ~w24966 & ~w24967;
assign w24969 = (w24933 & w24740) | (w24933 & w37338) | (w24740 & w37338);
assign w24970 = ~w24741 & ~w24933;
assign w24971 = ~w24740 & w24970;
assign w24972 = w24703 & ~w24971;
assign w24973 = ~w24969 & w24972;
assign w24974 = ~w24738 & w24973;
assign w24975 = ~w24969 & ~w24971;
assign w24976 = w24897 & ~w24975;
assign w24977 = ~w24974 & ~w24976;
assign w24978 = w8298 & w21771;
assign w24979 = ~w21760 & w37339;
assign w24980 = w8277 & ~w22020;
assign w24981 = ~w24498 & w37340;
assign w24982 = ~w24979 & ~w24980;
assign w24983 = ~w24978 & w24982;
assign w24984 = ~w24981 & w37341;
assign w24985 = (a_8 & w24981) | (a_8 & w37342) | (w24981 & w37342);
assign w24986 = ~w24984 & ~w24985;
assign w24987 = ~w24887 & ~w24921;
assign w24988 = w24887 & w24921;
assign w24989 = ~w24987 & ~w24988;
assign w24990 = w24912 & w24989;
assign w24991 = w24773 & w24990;
assign w24992 = w24912 & ~w24989;
assign w24993 = ~w24773 & w24992;
assign w24994 = ~w24991 & ~w24993;
assign w24995 = ~w24741 & w24994;
assign w24996 = ~w24740 & w24995;
assign w24997 = ~w24772 & w32184;
assign w24998 = (w24989 & w24772) | (w24989 & w32185) | (w24772 & w32185);
assign w24999 = ~w24997 & ~w24998;
assign w25000 = ~w24912 & ~w24999;
assign w25001 = (~w25000 & ~w24995) | (~w25000 & w32186) | (~w24995 & w32186);
assign w25002 = ~w24770 & ~w24988;
assign w25003 = ~w24772 & w25002;
assign w25004 = ~w24882 & ~w24885;
assign w25005 = w5080 & w21901;
assign w25006 = ~w21882 & w37343;
assign w25007 = w5286 & w21892;
assign w25008 = ~w25005 & ~w25006;
assign w25009 = ~w25007 & w25008;
assign w25010 = (w22096 & w32562) | (w22096 & w32563) | (w32562 & w32563);
assign w25011 = (~w22096 & w32564) | (~w22096 & w32565) | (w32564 & w32565);
assign w25012 = ~w25010 & ~w25011;
assign w25013 = w1226 & w22107;
assign w25014 = w21873 & w32188;
assign w25015 = w1226 & ~w21854;
assign w25016 = ~w21787 & w25015;
assign w25017 = ~w25014 & ~w25016;
assign w25018 = ~w22105 & ~w25017;
assign w25019 = ~w518 & ~w21839;
assign w25020 = w4638 & w21854;
assign w25021 = w4666 & w21787;
assign w25022 = ~w25019 & ~w25020;
assign w25023 = ~w25021 & w25022;
assign w25024 = ~w25018 & w25023;
assign w25025 = ~w25013 & w25024;
assign w25026 = a_26 & ~w25025;
assign w25027 = ~a_26 & w25025;
assign w25028 = ~w25026 & ~w25027;
assign w25029 = ~w21796 & w37344;
assign w25030 = w4446 & w21833;
assign w25031 = (~w25029 & w21803) | (~w25029 & w37345) | (w21803 & w37345);
assign w25032 = ~w25030 & w25031;
assign w25033 = (w25032 & w23150) | (w25032 & w32566) | (w23150 & w32566);
assign w25034 = ~w62 & w13336;
assign w25035 = w387 & w935;
assign w25036 = w1344 & w1360;
assign w25037 = w2151 & w3274;
assign w25038 = w3518 & w3979;
assign w25039 = w4912 & w25038;
assign w25040 = w25036 & w25037;
assign w25041 = w25034 & w25035;
assign w25042 = w25040 & w25041;
assign w25043 = w2188 & w25039;
assign w25044 = w4145 & w4524;
assign w25045 = w25043 & w25044;
assign w25046 = w5530 & w25042;
assign w25047 = w25045 & w25046;
assign w25048 = w6707 & w25047;
assign w25049 = w15174 & w25048;
assign w25050 = ~w24804 & w37346;
assign w25051 = (w25049 & w24804) | (w25049 & w37347) | (w24804 & w37347);
assign w25052 = ~w25050 & ~w25051;
assign w25053 = w1478 & ~w22161;
assign w25054 = w21815 & w1399;
assign w25055 = w668 & w21807;
assign w25056 = (~w25054 & ~w21813) | (~w25054 & w37348) | (~w21813 & w37348);
assign w25057 = ~w25055 & w25056;
assign w25058 = ~w25053 & w25057;
assign w25059 = w25052 & ~w25058;
assign w25060 = ~w25052 & w25058;
assign w25061 = ~w25059 & ~w25060;
assign w25062 = a_29 & w25061;
assign w25063 = w25033 & w25062;
assign w25064 = ~a_29 & w25061;
assign w25065 = ~w25033 & w25064;
assign w25066 = ~w25063 & ~w25065;
assign w25067 = ~a_29 & ~w25061;
assign w25068 = w25033 & w25067;
assign w25069 = a_29 & ~w25061;
assign w25070 = ~w25033 & w25069;
assign w25071 = ~w25068 & ~w25070;
assign w25072 = w25066 & w25071;
assign w25073 = ~w24844 & ~w24856;
assign w25074 = ~w24843 & ~w25073;
assign w25075 = w25072 & ~w25074;
assign w25076 = ~w25072 & w25074;
assign w25077 = ~w25075 & ~w25076;
assign w25078 = w25028 & ~w25077;
assign w25079 = ~w25028 & w25077;
assign w25080 = ~w25078 & ~w25079;
assign w25081 = ~w24861 & w24863;
assign w25082 = ~w24860 & ~w25081;
assign w25083 = w25080 & w25082;
assign w25084 = ~w25080 & ~w25082;
assign w25085 = ~w25083 & ~w25084;
assign w25086 = w25012 & ~w25085;
assign w25087 = ~w25012 & w25085;
assign w25088 = ~w25086 & ~w25087;
assign w25089 = ~w24868 & ~w24871;
assign w25090 = w25088 & w25089;
assign w25091 = ~w25088 & ~w25089;
assign w25092 = ~w25090 & ~w25091;
assign w25093 = ~w22901 & w32189;
assign w25094 = w5818 & w21921;
assign w25095 = w5308 & ~w21910;
assign w25096 = w5816 & w21951;
assign w25097 = ~w25094 & ~w25095;
assign w25098 = ~w25096 & w25097;
assign w25099 = (a_20 & w25093) | (a_20 & w37349) | (w25093 & w37349);
assign w25100 = ~w25093 & w37350;
assign w25101 = ~w25099 & ~w25100;
assign w25102 = w8391 & w23310;
assign w25103 = w6059 & ~w21945;
assign w25104 = w6061 & ~w21940;
assign w25105 = w6304 & w21934;
assign w25106 = ~w25103 & ~w25104;
assign w25107 = (~a_17 & ~w25106) | (~a_17 & w37351) | (~w25106 & w37351);
assign w25108 = w25106 & w37352;
assign w25109 = ~w25107 & ~w25108;
assign w25110 = (w25109 & ~w32190) | (w25109 & w37353) | (~w32190 & w37353);
assign w25111 = ~w25102 & ~w25110;
assign w25112 = w25101 & ~w25111;
assign w25113 = ~w25101 & w25111;
assign w25114 = ~w25112 & ~w25113;
assign w25115 = w25092 & w25114;
assign w25116 = ~w25092 & ~w25114;
assign w25117 = ~w25115 & ~w25116;
assign w25118 = w25004 & ~w25117;
assign w25119 = ~w25004 & w25117;
assign w25120 = ~w25118 & ~w25119;
assign w25121 = (~w25120 & w25003) | (~w25120 & w32191) | (w25003 & w32191);
assign w25122 = ~w25003 & w32192;
assign w25123 = ~w25121 & ~w25122;
assign w25124 = w7511 & w22014;
assign w25125 = w7192 & ~w21992;
assign w25126 = w7489 & w22007;
assign w25127 = ~w23397 & w37354;
assign w25128 = ~w25125 & ~w25126;
assign w25129 = ~w25124 & w25128;
assign w25130 = ~w25127 & w37355;
assign w25131 = (~a_11 & w25127) | (~a_11 & w37356) | (w25127 & w37356);
assign w25132 = ~w25130 & ~w25131;
assign w25133 = w6996 & w21985;
assign w25134 = w6446 & ~w21968;
assign w25135 = w6998 & ~w21973;
assign w25136 = ~w23551 & w37357;
assign w25137 = ~w25133 & ~w25134;
assign w25138 = ~w25135 & w25137;
assign w25139 = (a_14 & w25136) | (a_14 & w37358) | (w25136 & w37358);
assign w25140 = ~w25136 & w37359;
assign w25141 = ~w25139 & ~w25140;
assign w25142 = w25132 & ~w25141;
assign w25143 = ~w25132 & w25141;
assign w25144 = ~w25142 & ~w25143;
assign w25145 = w25123 & ~w25144;
assign w25146 = ~w25123 & w25144;
assign w25147 = ~w25145 & ~w25146;
assign w25148 = w25001 & w25147;
assign w25149 = ~w25001 & ~w25147;
assign w25150 = ~w25148 & ~w25149;
assign w25151 = w24986 & ~w25150;
assign w25152 = ~w24986 & w25150;
assign w25153 = ~w25151 & ~w25152;
assign w25154 = w24977 & w25153;
assign w25155 = ~w24977 & ~w25153;
assign w25156 = ~w25154 & ~w25155;
assign w25157 = ~w24752 & w24975;
assign w25158 = w24739 & ~w25157;
assign w25159 = ~w24752 & ~w24975;
assign w25160 = ~w24739 & ~w25159;
assign w25161 = ~w25158 & ~w25160;
assign w25162 = w24720 & ~w25161;
assign w25163 = w24523 & w25162;
assign w25164 = ~w24736 & w24752;
assign w25165 = w24736 & ~w24752;
assign w25166 = (~w32171 & w37360) | (~w32171 & w37361) | (w37360 & w37361);
assign w25167 = ~w24974 & ~w25166;
assign w25168 = ~w25165 & w25167;
assign w25169 = ~w25164 & ~w25168;
assign w25170 = ~w25163 & w25169;
assign w25171 = w24968 & ~w25156;
assign w25172 = w25170 & w25171;
assign w25173 = w24968 & w25156;
assign w25174 = ~w25170 & w25173;
assign w25175 = ~w25172 & ~w25174;
assign w25176 = ~w24954 & w25175;
assign w25177 = ~w24953 & w25176;
assign w25178 = ~w25156 & ~w25170;
assign w25179 = w24986 & w25156;
assign w25180 = ~w25132 & w25150;
assign w25181 = (~w25150 & w24974) | (~w25150 & w32193) | (w24974 & w32193);
assign w25182 = ~w25180 & ~w25181;
assign w25183 = w25123 & w25141;
assign w25184 = ~w25003 & w32194;
assign w25185 = ~w25120 & ~w25141;
assign w25186 = (~w25185 & w25003) | (~w25185 & w32195) | (w25003 & w32195);
assign w25187 = ~w25184 & ~w25186;
assign w25188 = ~w25000 & ~w25187;
assign w25189 = ~w24996 & w25188;
assign w25190 = (~w25183 & w24996) | (~w25183 & w32196) | (w24996 & w32196);
assign w25191 = w8277 & w21771;
assign w25192 = ~w21760 & w37362;
assign w25193 = w8295 & ~w22035;
assign w25194 = ~w25192 & ~w25193;
assign w25195 = ~w25191 & w25194;
assign w25196 = (w25195 & ~w24529) | (w25195 & w37363) | (~w24529 & w37363);
assign w25197 = ~a_8 & w25196;
assign w25198 = (w24529 & w37364) | (w24529 & w37365) | (w37364 & w37365);
assign w25199 = ~w25197 & ~w25198;
assign w25200 = w9788 & ~w21757;
assign w25201 = w9780 & w22039;
assign w25202 = w9786 & w22032;
assign w25203 = (w22048 & w22042) | (w22048 & w37366) | (w22042 & w37366);
assign w25204 = ~w22042 & w37367;
assign w25205 = ~w25203 & ~w25204;
assign w25206 = ~w25201 & ~w25202;
assign w25207 = ~w25200 & w25206;
assign w25208 = (w25207 & w25205) | (w25207 & w37368) | (w25205 & w37368);
assign w25209 = a_5 & ~w25208;
assign w25210 = (w25205 & w37369) | (w25205 & w37370) | (w37369 & w37370);
assign w25211 = ~w25209 & ~w25210;
assign w25212 = ~w25199 & ~w25211;
assign w25213 = (~w32196 & w37371) | (~w32196 & w37372) | (w37371 & w37372);
assign w25214 = w25199 & ~w25211;
assign w25215 = (w32196 & w37373) | (w32196 & w37374) | (w37373 & w37374);
assign w25216 = ~w25213 & ~w25215;
assign w25217 = w25111 & ~w25120;
assign w25218 = ~w25111 & w25118;
assign w25219 = w25092 & w25112;
assign w25220 = ~w25101 & ~w25111;
assign w25221 = ~w25092 & w25220;
assign w25222 = ~w25219 & ~w25221;
assign w25223 = ~w25004 & ~w25222;
assign w25224 = ~w24987 & ~w25223;
assign w25225 = ~w25218 & w25224;
assign w25226 = (~w25217 & w25003) | (~w25217 & w32197) | (w25003 & w32197);
assign w25227 = w25092 & ~w25101;
assign w25228 = ~w25092 & w25101;
assign w25229 = w25004 & ~w25228;
assign w25230 = (~w25227 & ~w25004) | (~w25227 & w32567) | (~w25004 & w32567);
assign w25231 = w5816 & ~w21945;
assign w25232 = w5818 & w21951;
assign w25233 = w5308 & w21921;
assign w25234 = ~w25232 & ~w25233;
assign w25235 = ~w25231 & w25234;
assign w25236 = (w25235 & ~w22083) | (w25235 & w37375) | (~w22083 & w37375);
assign w25237 = a_20 & ~w25236;
assign w25238 = (~w22083 & w37376) | (~w22083 & w37377) | (w37376 & w37377);
assign w25239 = ~w25237 & ~w25238;
assign w25240 = w5016 & w21901;
assign w25241 = w5080 & w21892;
assign w25242 = w5286 & ~w21910;
assign w25243 = ~w25240 & ~w25241;
assign w25244 = (a_23 & ~w25243) | (a_23 & w37378) | (~w25243 & w37378);
assign w25245 = w5017 & ~w22580;
assign w25246 = w25243 & w37379;
assign w25247 = ~w25245 & w25246;
assign w25248 = (~w25244 & w22580) | (~w25244 & w37380) | (w22580 & w37380);
assign w25249 = ~w25247 & w25248;
assign w25250 = ~w25079 & ~w25082;
assign w25251 = (~w25078 & w25082) | (~w25078 & w32568) | (w25082 & w32568);
assign w25252 = w4446 & ~w21839;
assign w25253 = w4068 & w21833;
assign w25254 = w3957 & ~w21803;
assign w25255 = ~w25253 & ~w25254;
assign w25256 = (a_29 & w25252) | (a_29 & w37381) | (w25252 & w37381);
assign w25257 = ~w25252 & w37382;
assign w25258 = ~w25256 & ~w25257;
assign w25259 = ~w22278 & w25258;
assign w25260 = ~w7268 & ~w7269;
assign w25261 = ~w25252 & w37383;
assign w25262 = ~w25256 & ~w25261;
assign w25263 = w22278 & w25262;
assign w25264 = ~w25259 & ~w25263;
assign w25265 = ~w21817 & w32198;
assign w25266 = ~w22137 & w25265;
assign w25267 = (w1478 & w21817) | (w1478 & w32199) | (w21817 & w32199);
assign w25268 = w22137 & w25267;
assign w25269 = ~w25266 & ~w25268;
assign w25270 = ~w21796 & w32200;
assign w25271 = w1399 & w21813;
assign w25272 = w1327 & w21807;
assign w25273 = ~w25271 & ~w25272;
assign w25274 = ~w25270 & w25273;
assign w25275 = w340 & w1153;
assign w25276 = ~w67 & ~w83;
assign w25277 = w2621 & w25276;
assign w25278 = w753 & w1663;
assign w25279 = w1686 & w1960;
assign w25280 = w3209 & w5390;
assign w25281 = w6635 & w25280;
assign w25282 = w25278 & w25279;
assign w25283 = w91 & w25275;
assign w25284 = w25277 & w25283;
assign w25285 = w25281 & w25282;
assign w25286 = w3492 & w4547;
assign w25287 = w25285 & w25286;
assign w25288 = w5585 & w25284;
assign w25289 = w25287 & w25288;
assign w25290 = w3699 & w25289;
assign w25291 = w3206 & w25290;
assign w25292 = w25274 & w25291;
assign w25293 = w25269 & w25292;
assign w25294 = (~w25291 & ~w25269) | (~w25291 & w32201) | (~w25269 & w32201);
assign w25295 = ~w25293 & ~w25294;
assign w25296 = (~w25050 & w25058) | (~w25050 & w32202) | (w25058 & w32202);
assign w25297 = w25295 & ~w25296;
assign w25298 = ~w25295 & w25296;
assign w25299 = ~w25297 & ~w25298;
assign w25300 = ~w25264 & w25299;
assign w25301 = w25264 & ~w25299;
assign w25302 = ~w25300 & ~w25301;
assign w25303 = (w25071 & w25074) | (w25071 & w32569) | (w25074 & w32569);
assign w25304 = ~w25302 & ~w25303;
assign w25305 = w25302 & w25303;
assign w25306 = ~w25304 & ~w25305;
assign w25307 = ~w21882 & w32204;
assign w25308 = ~w22381 & w25307;
assign w25309 = ~w21882 & w32205;
assign w25310 = w4638 & w21787;
assign w25311 = ~w518 & w21854;
assign w25312 = ~w25310 & ~w25311;
assign w25313 = ~w25309 & w25312;
assign w25314 = ~w25308 & w25313;
assign w25315 = (a_26 & ~w25314) | (a_26 & w32206) | (~w25314 & w32206);
assign w25316 = w25314 & w32207;
assign w25317 = ~w25315 & ~w25316;
assign w25318 = w25306 & w25317;
assign w25319 = ~w25306 & ~w25317;
assign w25320 = ~w25318 & ~w25319;
assign w25321 = w25251 & ~w25320;
assign w25322 = ~w25251 & w25320;
assign w25323 = ~w25321 & ~w25322;
assign w25324 = w25249 & w25323;
assign w25325 = ~w25249 & ~w25323;
assign w25326 = ~w25324 & ~w25325;
assign w25327 = ~w24868 & ~w25086;
assign w25328 = ~w24871 & w25327;
assign w25329 = ~w25087 & ~w25328;
assign w25330 = w25326 & ~w25329;
assign w25331 = ~w25326 & w25329;
assign w25332 = ~w25330 & ~w25331;
assign w25333 = w25239 & ~w25332;
assign w25334 = ~w25239 & w25332;
assign w25335 = ~w25333 & ~w25334;
assign w25336 = w6304 & ~w21968;
assign w25337 = w6061 & w21934;
assign w25338 = w6059 & ~w21940;
assign w25339 = ~w25337 & ~w25338;
assign w25340 = ~w25336 & w25339;
assign w25341 = (w25340 & w23366) | (w25340 & w37384) | (w23366 & w37384);
assign w25342 = a_17 & ~w25341;
assign w25343 = (w23366 & w37385) | (w23366 & w37386) | (w37385 & w37386);
assign w25344 = ~w25342 & ~w25343;
assign w25345 = w6998 & w21985;
assign w25346 = w6446 & ~w21973;
assign w25347 = w6996 & ~w21992;
assign w25348 = ~w25345 & ~w25346;
assign w25349 = (a_14 & ~w25348) | (a_14 & w37387) | (~w25348 & w37387);
assign w25350 = w8592 & ~w23930;
assign w25351 = w25348 & w37388;
assign w25352 = ~w25350 & w25351;
assign w25353 = (~w25349 & w23930) | (~w25349 & w37389) | (w23930 & w37389);
assign w25354 = ~w25352 & w25353;
assign w25355 = w25344 & w25354;
assign w25356 = ~w25335 & w25355;
assign w25357 = ~w25344 & w25354;
assign w25358 = w25335 & w25357;
assign w25359 = ~w25356 & ~w25358;
assign w25360 = w25230 & w25359;
assign w25361 = w25335 & w25355;
assign w25362 = ~w25335 & w25357;
assign w25363 = ~w25361 & ~w25362;
assign w25364 = ~w25230 & w25363;
assign w25365 = ~w25360 & ~w25364;
assign w25366 = ~w25226 & w25365;
assign w25367 = w25230 & ~w25363;
assign w25368 = ~w25230 & ~w25359;
assign w25369 = ~w25367 & ~w25368;
assign w25370 = w25226 & ~w25369;
assign w25371 = ~w25366 & ~w25370;
assign w25372 = ~w25344 & ~w25354;
assign w25373 = ~w25335 & w25372;
assign w25374 = w25344 & ~w25354;
assign w25375 = w25335 & w25374;
assign w25376 = ~w25373 & ~w25375;
assign w25377 = w25230 & w25376;
assign w25378 = w25335 & w25372;
assign w25379 = ~w25335 & w25374;
assign w25380 = ~w25378 & ~w25379;
assign w25381 = ~w25230 & w25380;
assign w25382 = ~w25377 & ~w25381;
assign w25383 = ~w25226 & w25382;
assign w25384 = w25230 & ~w25380;
assign w25385 = ~w25230 & ~w25376;
assign w25386 = ~w25384 & ~w25385;
assign w25387 = w25226 & ~w25386;
assign w25388 = ~w25383 & ~w25387;
assign w25389 = w25371 & w25388;
assign w25390 = w9061 & w24122;
assign w25391 = w7489 & w22014;
assign w25392 = w7192 & w22007;
assign w25393 = w7511 & ~w22020;
assign w25394 = ~w25391 & ~w25392;
assign w25395 = w25394 & w37390;
assign w25396 = (~a_11 & ~w25394) | (~a_11 & w37391) | (~w25394 & w37391);
assign w25397 = ~w25395 & ~w25396;
assign w25398 = (w25397 & ~w24122) | (w25397 & w37392) | (~w24122 & w37392);
assign w25399 = ~w25390 & ~w25398;
assign w25400 = w25389 & ~w25399;
assign w25401 = ~w25389 & w25399;
assign w25402 = ~w25400 & ~w25401;
assign w25403 = ~w25216 & ~w25402;
assign w25404 = (~w32196 & w37393) | (~w32196 & w37394) | (w37393 & w37394);
assign w25405 = (w32196 & w37395) | (w32196 & w37396) | (w37395 & w37396);
assign w25406 = ~w25404 & ~w25405;
assign w25407 = w25402 & w25406;
assign w25408 = ~w25403 & ~w25407;
assign w25409 = w25182 & ~w25408;
assign w25410 = ~w25402 & w25406;
assign w25411 = ~w25216 & w25402;
assign w25412 = ~w25410 & ~w25411;
assign w25413 = ~w25182 & ~w25412;
assign w25414 = ~w25409 & ~w25413;
assign w25415 = ~w25179 & ~w25414;
assign w25416 = ~w25178 & w25415;
assign w25417 = ~w24968 & w25156;
assign w25418 = w25170 & w25417;
assign w25419 = ~w24968 & ~w25156;
assign w25420 = ~w25170 & w25419;
assign w25421 = ~w25418 & ~w25420;
assign w25422 = (~w25179 & w25170) | (~w25179 & w32208) | (w25170 & w32208);
assign w25423 = w25182 & w25412;
assign w25424 = ~w25182 & w25408;
assign w25425 = ~w25423 & ~w25424;
assign w25426 = (~w32208 & w37397) | (~w32208 & w37398) | (w37397 & w37398);
assign w25427 = ~w25416 & w25421;
assign w25428 = ~w25426 & w25427;
assign w25429 = ~w25177 & w25428;
assign w25430 = ~w25190 & w25400;
assign w25431 = ~w25389 & ~w25399;
assign w25432 = w25190 & w25431;
assign w25433 = ~w25430 & ~w25432;
assign w25434 = ~w25190 & w25401;
assign w25435 = w25389 & w25399;
assign w25436 = w25190 & w25435;
assign w25437 = ~w25434 & ~w25436;
assign w25438 = w25433 & w25437;
assign w25439 = w25199 & w25438;
assign w25440 = w25182 & w25439;
assign w25441 = w25199 & ~w25438;
assign w25442 = ~w25182 & w25441;
assign w25443 = ~w25440 & ~w25442;
assign w25444 = ~w25199 & ~w25438;
assign w25445 = w25182 & w25444;
assign w25446 = ~w25199 & w25438;
assign w25447 = ~w25182 & w25446;
assign w25448 = ~w25445 & ~w25447;
assign w25449 = w25443 & w25448;
assign w25450 = w25211 & w25449;
assign w25451 = w25422 & w25450;
assign w25452 = w25211 & ~w25449;
assign w25453 = ~w25422 & w25452;
assign w25454 = ~w25451 & ~w25453;
assign w25455 = ~w25429 & w25454;
assign w25456 = ~w25179 & w25443;
assign w25457 = ~w25178 & w25456;
assign w25458 = ~w25180 & w25437;
assign w25459 = ~w25181 & w25458;
assign w25460 = w25433 & ~w25459;
assign w25461 = ~w25335 & w25344;
assign w25462 = w25230 & w25461;
assign w25463 = w25335 & w25344;
assign w25464 = ~w25230 & w25463;
assign w25465 = ~w25462 & ~w25464;
assign w25466 = ~w25217 & w25465;
assign w25467 = ~w25230 & ~w25335;
assign w25468 = w25230 & w25335;
assign w25469 = ~w25467 & ~w25468;
assign w25470 = ~w25344 & ~w25469;
assign w25471 = (~w25470 & ~w25466) | (~w25470 & w37399) | (~w25466 & w37399);
assign w25472 = ~w25227 & ~w25334;
assign w25473 = ~w25229 & w25472;
assign w25474 = ~w25333 & ~w25473;
assign w25475 = (~w25324 & w25328) | (~w25324 & w32570) | (w25328 & w32570);
assign w25476 = ~w25325 & ~w25475;
assign w25477 = w5080 & ~w21910;
assign w25478 = w5016 & w21892;
assign w25479 = w5286 & w21921;
assign w25480 = ~w25477 & ~w25478;
assign w25481 = ~w25479 & w25480;
assign w25482 = (w25481 & ~w22664) | (w25481 & w37400) | (~w22664 & w37400);
assign w25483 = a_23 & w25482;
assign w25484 = (w22664 & w37401) | (w22664 & w37402) | (w37401 & w37402);
assign w25485 = ~w25483 & ~w25484;
assign w25486 = ~w25300 & ~w25303;
assign w25487 = w4070 & w22247;
assign w25488 = w4070 & ~w22246;
assign w25489 = w3957 & w21833;
assign w25490 = w4068 & ~w21839;
assign w25491 = (~w25489 & ~w21854) | (~w25489 & w37403) | (~w21854 & w37403);
assign w25492 = ~w25490 & w25491;
assign w25493 = (w25492 & ~w25488) | (w25492 & w37404) | (~w25488 & w37404);
assign w25494 = ~w25487 & w25493;
assign w25495 = ~w21819 & w32210;
assign w25496 = ~w22177 & w25495;
assign w25497 = (w1478 & w21819) | (w1478 & w32211) | (w21819 & w32211);
assign w25498 = w22177 & w25497;
assign w25499 = ~w21796 & w37405;
assign w25500 = w668 & ~w21803;
assign w25501 = w1399 & w21807;
assign w25502 = ~w25499 & ~w25501;
assign w25503 = ~w25500 & w25502;
assign w25504 = ~w25498 & w25503;
assign w25505 = ~w164 & ~w239;
assign w25506 = ~w316 & ~w355;
assign w25507 = w25505 & w25506;
assign w25508 = w945 & w2527;
assign w25509 = w3080 & w25508;
assign w25510 = w5857 & w25507;
assign w25511 = w13059 & w25510;
assign w25512 = w2575 & w25509;
assign w25513 = w13055 & w25512;
assign w25514 = w25511 & w25513;
assign w25515 = w111 & w25514;
assign w25516 = w15221 & w25515;
assign w25517 = (~w25516 & ~w25504) | (~w25516 & w32212) | (~w25504 & w32212);
assign w25518 = (w25516 & w22177) | (w25516 & w32571) | (w22177 & w32571);
assign w25519 = w25504 & w25518;
assign w25520 = ~w25517 & ~w25519;
assign w25521 = ~w25293 & ~w25296;
assign w25522 = ~w25294 & ~w25521;
assign w25523 = (a_29 & w25521) | (a_29 & w32213) | (w25521 & w32213);
assign w25524 = ~w25521 & w32214;
assign w25525 = ~w25523 & ~w25524;
assign w25526 = w25520 & ~w25525;
assign w25527 = ~w25520 & w25525;
assign w25528 = ~w25526 & ~w25527;
assign w25529 = w25494 & w25528;
assign w25530 = ~w25494 & ~w25528;
assign w25531 = ~w25529 & ~w25530;
assign w25532 = ~w25301 & w25531;
assign w25533 = w25531 & w32572;
assign w25534 = ~w25300 & ~w25531;
assign w25535 = ~w25305 & w25534;
assign w25536 = ~w25533 & ~w25535;
assign w25537 = ~w518 & w21787;
assign w25538 = ~w21882 & w37406;
assign w25539 = (~w25537 & ~w21901) | (~w25537 & w37407) | (~w21901 & w37407);
assign w25540 = ~w25538 & w25539;
assign w25541 = ~a_26 & w25540;
assign w25542 = (w25541 & ~w22555) | (w25541 & w32215) | (~w22555 & w32215);
assign w25543 = a_26 & ~w25540;
assign w25544 = (~w25543 & ~w22555) | (~w25543 & w32216) | (~w22555 & w32216);
assign w25545 = ~w25542 & w25544;
assign w25546 = w25536 & w25545;
assign w25547 = ~w25536 & ~w25545;
assign w25548 = ~w25546 & ~w25547;
assign w25549 = ~w25078 & ~w25318;
assign w25550 = ~w25250 & w25549;
assign w25551 = ~w25319 & ~w25550;
assign w25552 = w25548 & ~w25551;
assign w25553 = ~w25548 & w25551;
assign w25554 = ~w25552 & ~w25553;
assign w25555 = ~w25485 & ~w25554;
assign w25556 = w25485 & w25554;
assign w25557 = ~w25555 & ~w25556;
assign w25558 = w25476 & ~w25557;
assign w25559 = ~w25476 & w25557;
assign w25560 = ~w25558 & ~w25559;
assign w25561 = w5818 & ~w21945;
assign w25562 = w5308 & w21951;
assign w25563 = w5816 & ~w21940;
assign w25564 = ~w25561 & ~w25562;
assign w25565 = ~w25563 & w25564;
assign w25566 = (w25565 & ~w23032) | (w25565 & w37408) | (~w23032 & w37408);
assign w25567 = a_20 & ~w25566;
assign w25568 = (~w23032 & w37409) | (~w23032 & w37410) | (w37409 & w37410);
assign w25569 = ~w25567 & ~w25568;
assign w25570 = w8391 & ~w22930;
assign w25571 = w6061 & ~w21968;
assign w25572 = w6059 & w21934;
assign w25573 = w6304 & ~w21973;
assign w25574 = ~w25571 & ~w25572;
assign w25575 = ~w25573 & w25574;
assign w25576 = ~a_17 & ~w25575;
assign w25577 = a_17 & w25575;
assign w25578 = ~w25576 & ~w25577;
assign w25579 = (w25578 & w22930) | (w25578 & w37411) | (w22930 & w37411);
assign w25580 = ~w25570 & ~w25579;
assign w25581 = ~w25569 & ~w25580;
assign w25582 = w25560 & ~w25581;
assign w25583 = w25569 & ~w25580;
assign w25584 = ~w25560 & ~w25583;
assign w25585 = ~w25582 & ~w25584;
assign w25586 = w25474 & ~w25585;
assign w25587 = w25560 & ~w25583;
assign w25588 = ~w25560 & ~w25581;
assign w25589 = ~w25587 & ~w25588;
assign w25590 = ~w25474 & ~w25589;
assign w25591 = ~w25586 & ~w25590;
assign w25592 = w25569 & w25580;
assign w25593 = w25560 & ~w25592;
assign w25594 = ~w25569 & w25580;
assign w25595 = ~w25560 & ~w25594;
assign w25596 = ~w25593 & ~w25595;
assign w25597 = w25474 & w25596;
assign w25598 = w25560 & ~w25594;
assign w25599 = ~w25560 & ~w25592;
assign w25600 = ~w25598 & ~w25599;
assign w25601 = ~w25474 & w25600;
assign w25602 = ~w25597 & ~w25601;
assign w25603 = ~w25591 & w25602;
assign w25604 = w6996 & w22007;
assign w25605 = w6998 & ~w21992;
assign w25606 = w6446 & w21985;
assign w25607 = ~w25605 & ~w25606;
assign w25608 = ~w25604 & w25607;
assign w25609 = (w25608 & ~w23580) | (w25608 & w37412) | (~w23580 & w37412);
assign w25610 = a_14 & ~w25609;
assign w25611 = (~w23580 & w37413) | (~w23580 & w37414) | (w37413 & w37414);
assign w25612 = ~w25610 & ~w25611;
assign w25613 = w9061 & w24295;
assign w25614 = w7489 & ~w22020;
assign w25615 = w7192 & w22014;
assign w25616 = w7511 & w21771;
assign w25617 = ~w25614 & ~w25615;
assign w25618 = w25617 & w37415;
assign w25619 = (~a_11 & ~w25617) | (~a_11 & w37416) | (~w25617 & w37416);
assign w25620 = ~w25618 & ~w25619;
assign w25621 = (w25620 & ~w24295) | (w25620 & w37417) | (~w24295 & w37417);
assign w25622 = ~w25613 & ~w25621;
assign w25623 = w25612 & ~w25622;
assign w25624 = ~w25603 & w25623;
assign w25625 = ~w25612 & ~w25622;
assign w25626 = w25603 & w25625;
assign w25627 = ~w25624 & ~w25626;
assign w25628 = ~w25471 & w25627;
assign w25629 = ~w25603 & w25625;
assign w25630 = w25603 & w25623;
assign w25631 = ~w25629 & ~w25630;
assign w25632 = w25471 & w25631;
assign w25633 = ~w25628 & ~w25632;
assign w25634 = ~w25612 & w25622;
assign w25635 = ~w25603 & w25634;
assign w25636 = w25612 & w25622;
assign w25637 = w25603 & w25636;
assign w25638 = ~w25635 & ~w25637;
assign w25639 = ~w25471 & w25638;
assign w25640 = ~w25603 & w25636;
assign w25641 = w25603 & w25634;
assign w25642 = ~w25640 & ~w25641;
assign w25643 = w25471 & w25642;
assign w25644 = ~w25639 & ~w25643;
assign w25645 = ~w25633 & ~w25644;
assign w25646 = ~w25183 & w25371;
assign w25647 = (w25388 & w25189) | (w25388 & w32217) | (w25189 & w32217);
assign w25648 = w8295 & w22032;
assign w25649 = ~w21760 & w37418;
assign w25650 = w8298 & ~w22035;
assign w25651 = ~w25648 & ~w25649;
assign w25652 = ~w25650 & w25651;
assign w25653 = (w25652 & ~w24756) | (w25652 & w37419) | (~w24756 & w37419);
assign w25654 = a_8 & ~w25653;
assign w25655 = (~w24756 & w37420) | (~w24756 & w37421) | (w37420 & w37421);
assign w25656 = ~w25654 & ~w25655;
assign w25657 = (w32217 & w37422) | (w32217 & w37423) | (w37422 & w37423);
assign w25658 = (~w32217 & w37424) | (~w32217 & w37425) | (w37424 & w37425);
assign w25659 = ~w25657 & ~w25658;
assign w25660 = w25645 & ~w25659;
assign w25661 = ~w25645 & w25659;
assign w25662 = ~w25660 & ~w25661;
assign w25663 = w25460 & w25662;
assign w25664 = ~w25460 & ~w25662;
assign w25665 = ~w25663 & ~w25664;
assign w25666 = (~w32209 & w37426) | (~w32209 & w37427) | (w37426 & w37427);
assign w25667 = w25448 & ~w25665;
assign w25668 = ~w25457 & w25667;
assign w25669 = ~w25666 & ~w25668;
assign w25670 = ~w21736 & w37428;
assign w25671 = w9780 & ~w21757;
assign w25672 = w9786 & w22039;
assign w25673 = ~w22046 & ~w22050;
assign w25674 = (~w22042 & w37429) | (~w22042 & w37430) | (w37429 & w37430);
assign w25675 = w22053 & ~w25674;
assign w25676 = ~w25671 & ~w25672;
assign w25677 = ~w25670 & w25676;
assign w25678 = (w25677 & w25675) | (w25677 & w37431) | (w25675 & w37431);
assign w25679 = ~a_5 & w25678;
assign w25680 = (~w25675 & w37432) | (~w25675 & w37433) | (w37432 & w37433);
assign w25681 = ~w25679 & ~w25680;
assign w25682 = ~w25669 & ~w25681;
assign w25683 = w25669 & w25681;
assign w25684 = ~w25682 & ~w25683;
assign w25685 = w25455 & w25684;
assign w25686 = ~w25455 & ~w25684;
assign w25687 = ~w25685 & ~w25686;
assign w25688 = w22071 & ~w25687;
assign w25689 = ~w22071 & w25687;
assign w25690 = ~w25688 & ~w25689;
assign w25691 = ~w25177 & w25421;
assign w25692 = ~w25416 & ~w25426;
assign w25693 = w25454 & w25692;
assign w25694 = w25691 & ~w25693;
assign w25695 = ~w25691 & w25693;
assign w25696 = ~w25694 & ~w25695;
assign w25697 = w3 & w21746;
assign w25698 = w10835 & w21752;
assign w25699 = (w22053 & w37435) | (w22053 & w37436) | (w37435 & w37436);
assign w25700 = ~w22061 & ~w25699;
assign w25701 = ~w25697 & ~w25698;
assign w25702 = (w25701 & w25700) | (w25701 & w37437) | (w25700 & w37437);
assign w25703 = (a_2 & ~w21755) | (a_2 & w34211) | (~w21755 & w34211);
assign w25704 = w25702 & ~w25703;
assign w25705 = (~w25700 & w37438) | (~w25700 & w37439) | (w37438 & w37439);
assign w25706 = ~w25704 & ~w25705;
assign w25707 = w25696 & ~w25706;
assign w25708 = ~w24306 & ~w24309;
assign w25709 = ~w24135 & ~w24136;
assign w25710 = w25708 & w25709;
assign w25711 = ~w25708 & ~w25709;
assign w25712 = ~w25710 & ~w25711;
assign w25713 = w3 & w22032;
assign w25714 = w10835 & ~w22035;
assign w25715 = ~w25713 & ~w25714;
assign w25716 = (w25715 & ~w24756) | (w25715 & w37440) | (~w24756 & w37440);
assign w25717 = (a_2 & ~w21762) | (a_2 & w34211) | (~w21762 & w34211);
assign w25718 = w25716 & ~w25717;
assign w25719 = (w24756 & w37441) | (w24756 & w37442) | (w37441 & w37442);
assign w25720 = ~w25718 & ~w25719;
assign w25721 = w25712 & ~w25720;
assign w25722 = ~w23605 & ~w23964;
assign w25723 = w23605 & w23964;
assign w25724 = ~w25722 & ~w25723;
assign w25725 = w3 & w21771;
assign w25726 = w10835 & ~w22020;
assign w25727 = ~w25725 & ~w25726;
assign w25728 = (w25727 & ~w24295) | (w25727 & w37443) | (~w24295 & w37443);
assign w25729 = (a_2 & ~w22014) | (a_2 & w34211) | (~w22014 & w34211);
assign w25730 = w25728 & ~w25729;
assign w25731 = (w24295 & w37444) | (w24295 & w37445) | (w37444 & w37445);
assign w25732 = ~w25730 & ~w25731;
assign w25733 = w25724 & w25732;
assign w25734 = w3 & ~w22020;
assign w25735 = w10835 & w22014;
assign w25736 = ~w25734 & ~w25735;
assign w25737 = (w25736 & ~w24122) | (w25736 & w37446) | (~w24122 & w37446);
assign w25738 = (a_2 & ~w22007) | (a_2 & w34211) | (~w22007 & w34211);
assign w25739 = w25737 & ~w25738;
assign w25740 = (w24122 & w37447) | (w24122 & w37448) | (w37447 & w37448);
assign w25741 = ~w25739 & ~w25740;
assign w25742 = ~w23937 & ~w23957;
assign w25743 = (w32543 & w37449) | (w32543 & w37450) | (w37449 & w37450);
assign w25744 = ~w23961 & ~w25743;
assign w25745 = w25742 & ~w25744;
assign w25746 = ~w25742 & w25744;
assign w25747 = ~w25745 & ~w25746;
assign w25748 = w25741 & w25747;
assign w25749 = w23903 & ~w23918;
assign w25750 = ~w23919 & ~w25749;
assign w25751 = w3 & ~w21992;
assign w25752 = w10835 & w21985;
assign w25753 = ~w25751 & ~w25752;
assign w25754 = (w25753 & w23930) | (w25753 & w37451) | (w23930 & w37451);
assign w25755 = (a_2 & w21973) | (a_2 & w34211) | (w21973 & w34211);
assign w25756 = w25754 & ~w25755;
assign w25757 = (~w23930 & w37452) | (~w23930 & w37453) | (w37452 & w37453);
assign w25758 = ~w25756 & ~w25757;
assign w25759 = ~w25750 & ~w25758;
assign w25760 = ~w23804 & ~w23821;
assign w25761 = ~w23822 & ~w25760;
assign w25762 = w10835 & w21921;
assign w25763 = w3 & w21951;
assign w25764 = ~w22901 & w37454;
assign w25765 = ~w25762 & ~w25763;
assign w25766 = ~w25764 & w25765;
assign w25767 = (a_2 & w21910) | (a_2 & w34211) | (w21910 & w34211);
assign w25768 = w25766 & ~w25767;
assign w25769 = (a_2 & w25764) | (a_2 & w37455) | (w25764 & w37455);
assign w25770 = ~w25768 & ~w25769;
assign w25771 = w25761 & w25770;
assign w25772 = w3 & ~w21945;
assign w25773 = w10835 & w21951;
assign w25774 = ~w25772 & ~w25773;
assign w25775 = (w25774 & ~w22083) | (w25774 & w37456) | (~w22083 & w37456);
assign w25776 = (a_2 & ~w21921) | (a_2 & w34211) | (~w21921 & w34211);
assign w25777 = w25775 & ~w25776;
assign w25778 = (w22083 & w37457) | (w22083 & w37458) | (w37457 & w37458);
assign w25779 = ~w25777 & ~w25778;
assign w25780 = ~w23650 & ~w23823;
assign w25781 = ~w23819 & ~w23822;
assign w25782 = ~w25780 & w25781;
assign w25783 = w25780 & ~w25781;
assign w25784 = ~w25782 & ~w25783;
assign w25785 = w25779 & w25784;
assign w25786 = ~w25761 & ~w25770;
assign w25787 = ~w23678 & ~w23799;
assign w25788 = ~w23800 & ~w25787;
assign w25789 = w3 & ~w21910;
assign w25790 = w10835 & w21892;
assign w25791 = ~w25789 & ~w25790;
assign w25792 = (w25791 & w22580) | (w25791 & w37459) | (w22580 & w37459);
assign w25793 = (a_2 & ~w21901) | (a_2 & w34211) | (~w21901 & w34211);
assign w25794 = w25792 & ~w25793;
assign w25795 = (~w22580 & w37460) | (~w22580 & w37461) | (w37460 & w37461);
assign w25796 = ~w25794 & ~w25795;
assign w25797 = ~w25788 & ~w25796;
assign w25798 = w25788 & w25796;
assign w25799 = ~w23696 & w23797;
assign w25800 = ~w23798 & ~w25799;
assign w25801 = ~w21882 & w37462;
assign w25802 = w10835 & w21901;
assign w25803 = w3 & w21892;
assign w25804 = ~w25802 & ~w25803;
assign w25805 = (w22096 & w32573) | (w22096 & w32574) | (w32573 & w32574);
assign w25806 = (~w22096 & w32575) | (~w22096 & w32576) | (w32575 & w32576);
assign w25807 = ~w25805 & ~w25806;
assign w25808 = ~w25801 & ~w25807;
assign w25809 = w25800 & ~w25808;
assign w25810 = ~w21882 & w37463;
assign w25811 = w3 & w21901;
assign w25812 = ~w25810 & ~w25811;
assign w25813 = (w25812 & ~w22555) | (w25812 & w32577) | (~w22555 & w32577);
assign w25814 = (a_2 & ~w21787) | (a_2 & w34211) | (~w21787 & w34211);
assign w25815 = w25813 & ~w25814;
assign w25816 = (w22555 & w37464) | (w22555 & w37465) | (w37464 & w37465);
assign w25817 = ~w25815 & ~w25816;
assign w25818 = ~w23710 & ~w23711;
assign w25819 = ~w23796 & w25818;
assign w25820 = w23796 & ~w25818;
assign w25821 = ~w25819 & ~w25820;
assign w25822 = w25817 & ~w25821;
assign w25823 = ~w25800 & w25808;
assign w25824 = ~w25817 & w25821;
assign w25825 = ~w23727 & ~w23728;
assign w25826 = ~w23794 & w25825;
assign w25827 = w23794 & ~w25825;
assign w25828 = ~w25826 & ~w25827;
assign w25829 = w10909 & w21854;
assign w25830 = ~w21882 & w37466;
assign w25831 = w10835 & w21787;
assign w25832 = ~w25830 & ~w25831;
assign w25833 = (~w23079 & w32578) | (~w23079 & w32579) | (w32578 & w32579);
assign w25834 = (w23079 & w32580) | (w23079 & w32581) | (w32580 & w32581);
assign w25835 = ~w25833 & ~w25834;
assign w25836 = ~w25829 & ~w25835;
assign w25837 = ~w25828 & ~w25836;
assign w25838 = w3 & w21787;
assign w25839 = w10835 & w21854;
assign w25840 = ~w25838 & ~w25839;
assign w25841 = (w25840 & w22726) | (w25840 & w37467) | (w22726 & w37467);
assign w25842 = a_2 & ~w25841;
assign w25843 = (a_2 & w21839) | (a_2 & w34211) | (w21839 & w34211);
assign w25844 = w25841 & ~w25843;
assign w25845 = ~w25842 & ~w25844;
assign w25846 = ~w23774 & ~w23789;
assign w25847 = w23788 & ~w23793;
assign w25848 = w25846 & ~w25847;
assign w25849 = ~w25846 & w25847;
assign w25850 = ~w25848 & ~w25849;
assign w25851 = w25845 & ~w25850;
assign w25852 = w10909 & w21833;
assign w25853 = w3 & w21854;
assign w25854 = w10835 & ~w21839;
assign w25855 = ~w25853 & ~w25854;
assign w25856 = (w25855 & w23698) | (w25855 & w37468) | (w23698 & w37468);
assign w25857 = ~a_2 & ~w25856;
assign w25858 = (w23698 & w37469) | (w23698 & w37470) | (w37469 & w37470);
assign w25859 = (~w25852 & w25857) | (~w25852 & w37471) | (w25857 & w37471);
assign w25860 = ~w23763 & ~w23789;
assign w25861 = w23773 & ~w25860;
assign w25862 = ~w23773 & w25860;
assign w25863 = ~w25861 & ~w25862;
assign w25864 = w25859 & ~w25863;
assign w25865 = ~w23176 & w23753;
assign w25866 = ~w23754 & ~w25865;
assign w25867 = w23736 & w25866;
assign w25868 = ~w23736 & ~w25866;
assign w25869 = ~w25867 & ~w25868;
assign w25870 = w10835 & w21833;
assign w25871 = w10837 & w22278;
assign w25872 = (~w25870 & w21839) | (~w25870 & w37472) | (w21839 & w37472);
assign w25873 = ~w25871 & w25872;
assign w25874 = (a_2 & w25871) | (a_2 & w37473) | (w25871 & w37473);
assign w25875 = (a_2 & w21803) | (a_2 & w34211) | (w21803 & w34211);
assign w25876 = w25873 & ~w25875;
assign w25877 = (~w25869 & w25876) | (~w25869 & w37474) | (w25876 & w37474);
assign w25878 = ~w25876 & w37475;
assign w25879 = w23745 & ~w23751;
assign w25880 = ~w23752 & ~w25879;
assign w25881 = ~w21796 & w37476;
assign w25882 = a_2 & ~w25881;
assign w25883 = w3 & w21833;
assign w25884 = w10835 & ~w21803;
assign w25885 = ~w25883 & ~w25884;
assign w25886 = (w25885 & w23150) | (w25885 & w37477) | (w23150 & w37477);
assign w25887 = ~w25882 & w25886;
assign w25888 = (~w23150 & w37478) | (~w23150 & w37479) | (w37478 & w37479);
assign w25889 = (~w25880 & w25887) | (~w25880 & w37480) | (w25887 & w37480);
assign w25890 = ~w25887 & w37481;
assign w25891 = w23738 & ~w23743;
assign w25892 = ~w23744 & ~w25891;
assign w25893 = w10835 & w21807;
assign w25894 = ~w21796 & w37482;
assign w25895 = ~w25893 & ~w25894;
assign w25896 = (w25895 & w23730) | (w25895 & w32582) | (w23730 & w32582);
assign w25897 = (~w23730 & w37483) | (~w23730 & w37484) | (w37483 & w37484);
assign w25898 = (a_2 & ~w21813) | (a_2 & w34211) | (~w21813 & w34211);
assign w25899 = w25896 & ~w25898;
assign w25900 = a_0 & w21807;
assign w25901 = a_2 & ~w21815;
assign w25902 = (w25901 & ~w21813) | (w25901 & w37485) | (~w21813 & w37485);
assign w25903 = (~w23737 & w25900) | (~w23737 & w37486) | (w25900 & w37486);
assign w25904 = ~w25897 & ~w25903;
assign w25905 = ~w25899 & w25904;
assign w25906 = w25892 & w25905;
assign w25907 = ~w25892 & ~w25905;
assign w25908 = ~w21796 & w37487;
assign w25909 = (~w25908 & w21803) | (~w25908 & w37488) | (w21803 & w37488);
assign w25910 = (w25909 & w23765) | (w25909 & w32583) | (w23765 & w32583);
assign w25911 = (a_2 & ~w21807) | (a_2 & w34211) | (~w21807 & w34211);
assign w25912 = w25910 & w25911;
assign w25913 = (~w23765 & w37489) | (~w23765 & w37490) | (w37489 & w37490);
assign w25914 = ~w25912 & ~w25913;
assign w25915 = (~w25906 & w25914) | (~w25906 & w37491) | (w25914 & w37491);
assign w25916 = (~w25889 & ~w25915) | (~w25889 & w37492) | (~w25915 & w37492);
assign w25917 = ~w25878 & ~w25916;
assign w25918 = ~w25877 & ~w25917;
assign w25919 = ~w25864 & ~w25918;
assign w25920 = ~w25859 & w25863;
assign w25921 = ~w25845 & w25850;
assign w25922 = ~w25920 & ~w25921;
assign w25923 = ~w25919 & w25922;
assign w25924 = (~w25851 & ~w25836) | (~w25851 & w37493) | (~w25836 & w37493);
assign w25925 = ~w25923 & w25924;
assign w25926 = ~w25824 & ~w25837;
assign w25927 = ~w25925 & w25926;
assign w25928 = ~w25822 & ~w25823;
assign w25929 = ~w25927 & w25928;
assign w25930 = (~w25798 & w25929) | (~w25798 & w37494) | (w25929 & w37494);
assign w25931 = ~w25797 & ~w25930;
assign w25932 = w10909 & w21892;
assign w25933 = w10835 & ~w21910;
assign w25934 = w3 & w21921;
assign w25935 = ~w25933 & ~w25934;
assign w25936 = (w25935 & ~w22664) | (w25935 & w37495) | (~w22664 & w37495);
assign w25937 = ~a_2 & ~w25936;
assign w25938 = (~w22664 & w37496) | (~w22664 & w37497) | (w37496 & w37497);
assign w25939 = (~w25932 & w25937) | (~w25932 & w37498) | (w25937 & w37498);
assign w25940 = ~w25931 & ~w25939;
assign w25941 = ~w23663 & ~w23801;
assign w25942 = ~w23676 & ~w23800;
assign w25943 = ~w25941 & ~w25942;
assign w25944 = w25941 & w25942;
assign w25945 = ~w25943 & ~w25944;
assign w25946 = (w25945 & w25930) | (w25945 & w37500) | (w25930 & w37500);
assign w25947 = ~w25940 & w37501;
assign w25948 = ~w25771 & ~w25785;
assign w25949 = ~w25947 & w25948;
assign w25950 = ~w25779 & ~w25784;
assign w25951 = w23826 & w23843;
assign w25952 = ~w23826 & ~w23843;
assign w25953 = ~w25951 & ~w25952;
assign w25954 = w10835 & ~w21945;
assign w25955 = w3 & ~w21940;
assign w25956 = ~w25954 & ~w25955;
assign w25957 = (w25956 & ~w23032) | (w25956 & w37502) | (~w23032 & w37502);
assign w25958 = (a_2 & ~w21951) | (a_2 & w34211) | (~w21951 & w34211);
assign w25959 = w25957 & ~w25958;
assign w25960 = (w23032 & w37503) | (w23032 & w37504) | (w37503 & w37504);
assign w25961 = ~w25959 & ~w25960;
assign w25962 = ~w25953 & ~w25961;
assign w25963 = ~w25950 & ~w25962;
assign w25964 = ~w25949 & w25963;
assign w25965 = w25953 & w25961;
assign w25966 = ~w23860 & ~w23863;
assign w25967 = ~w23841 & ~w25951;
assign w25968 = w25966 & ~w25967;
assign w25969 = ~w25966 & w25967;
assign w25970 = ~w25968 & ~w25969;
assign w25971 = w10835 & ~w21940;
assign w25972 = w3 & w21934;
assign w25973 = ~w25971 & ~w25972;
assign w25974 = (w25973 & ~w23310) | (w25973 & w37505) | (~w23310 & w37505);
assign w25975 = (a_2 & w21945) | (a_2 & w34211) | (w21945 & w34211);
assign w25976 = w25974 & ~w25975;
assign w25977 = (w23310 & w37506) | (w23310 & w37507) | (w37506 & w37507);
assign w25978 = ~w25976 & ~w25977;
assign w25979 = w25970 & w25978;
assign w25980 = ~w25964 & ~w25965;
assign w25981 = ~w25979 & w25980;
assign w25982 = ~w25970 & ~w25978;
assign w25983 = w23866 & ~w23880;
assign w25984 = ~w23881 & ~w25983;
assign w25985 = w3 & ~w21968;
assign w25986 = w10835 & w21934;
assign w25987 = ~w25985 & ~w25986;
assign w25988 = (w25987 & w23366) | (w25987 & w37508) | (w23366 & w37508);
assign w25989 = (a_2 & w21940) | (a_2 & w34211) | (w21940 & w34211);
assign w25990 = w25988 & ~w25989;
assign w25991 = (~w23366 & w37509) | (~w23366 & w37510) | (w37509 & w37510);
assign w25992 = ~w25990 & ~w25991;
assign w25993 = ~w25984 & ~w25992;
assign w25994 = ~w25982 & ~w25993;
assign w25995 = ~w25981 & w25994;
assign w25996 = w25984 & w25992;
assign w25997 = w3 & ~w21973;
assign w25998 = w10835 & ~w21968;
assign w25999 = ~w25997 & ~w25998;
assign w26000 = (w25999 & w22930) | (w25999 & w37511) | (w22930 & w37511);
assign w26001 = (a_2 & ~w21934) | (a_2 & w34211) | (~w21934 & w34211);
assign w26002 = w26000 & ~w26001;
assign w26003 = (~w22930 & w37512) | (~w22930 & w37513) | (w37512 & w37513);
assign w26004 = ~w26002 & ~w26003;
assign w26005 = ~w23896 & ~w23899;
assign w26006 = (~w23878 & w23866) | (~w23878 & w32584) | (w23866 & w32584);
assign w26007 = w26005 & w26006;
assign w26008 = ~w26005 & ~w26006;
assign w26009 = ~w26007 & ~w26008;
assign w26010 = (~w25996 & w26009) | (~w25996 & w37514) | (w26009 & w37514);
assign w26011 = ~w25995 & w26010;
assign w26012 = ~w26004 & w26009;
assign w26013 = w10835 & ~w21973;
assign w26014 = w3 & w21985;
assign w26015 = ~w23551 & w37515;
assign w26016 = ~w26013 & ~w26014;
assign w26017 = ~w26015 & w26016;
assign w26018 = (a_2 & w21968) | (a_2 & w34211) | (w21968 & w34211);
assign w26019 = w26017 & ~w26018;
assign w26020 = (a_2 & w26015) | (a_2 & w37516) | (w26015 & w37516);
assign w26021 = ~w26019 & ~w26020;
assign w26022 = (~w23899 & w23881) | (~w23899 & w32585) | (w23881 & w32585);
assign w26023 = ~w23635 & ~w23900;
assign w26024 = w26022 & w26023;
assign w26025 = ~w26022 & ~w26023;
assign w26026 = ~w26024 & ~w26025;
assign w26027 = ~w26021 & ~w26026;
assign w26028 = ~w26012 & ~w26027;
assign w26029 = ~w26011 & w26028;
assign w26030 = w26021 & w26026;
assign w26031 = (~w26030 & ~w25750) | (~w26030 & w32586) | (~w25750 & w32586);
assign w26032 = ~w26029 & w26031;
assign w26033 = w3 & w22014;
assign w26034 = w10835 & w22007;
assign w26035 = ~w23397 & w37517;
assign w26036 = ~w26033 & ~w26034;
assign w26037 = ~w26035 & w26036;
assign w26038 = (a_2 & w21992) | (a_2 & w34211) | (w21992 & w34211);
assign w26039 = w26037 & ~w26038;
assign w26040 = (a_2 & w26035) | (a_2 & w37518) | (w26035 & w37518);
assign w26041 = ~w26039 & ~w26040;
assign w26042 = ~w23954 & ~w26041;
assign w26043 = w23922 & w26042;
assign w26044 = w23954 & ~w26041;
assign w26045 = ~w23922 & w26044;
assign w26046 = ~w26043 & ~w26045;
assign w26047 = w3 & w22007;
assign w26048 = w10835 & ~w21992;
assign w26049 = ~w26047 & ~w26048;
assign w26050 = (w26049 & ~w23580) | (w26049 & w37519) | (~w23580 & w37519);
assign w26051 = (a_2 & ~w21985) | (a_2 & w34211) | (~w21985 & w34211);
assign w26052 = w26050 & ~w26051;
assign w26053 = (w23580 & w37520) | (w23580 & w37521) | (w37520 & w37521);
assign w26054 = ~w26052 & ~w26053;
assign w26055 = (~w23916 & w23903) | (~w23916 & w32587) | (w23903 & w32587);
assign w26056 = ~w23620 & ~w23920;
assign w26057 = w26055 & ~w26056;
assign w26058 = ~w26055 & w26056;
assign w26059 = ~w26057 & ~w26058;
assign w26060 = ~w26054 & ~w26059;
assign w26061 = ~w25759 & ~w26032;
assign w26062 = w26046 & ~w26060;
assign w26063 = w26061 & w26062;
assign w26064 = w26054 & w26059;
assign w26065 = w26046 & w26064;
assign w26066 = (~w32543 & w37522) | (~w32543 & w37523) | (w37522 & w37523);
assign w26067 = ~w25743 & w26041;
assign w26068 = ~w26066 & w26067;
assign w26069 = ~w26065 & ~w26068;
assign w26070 = ~w26063 & w26069;
assign w26071 = ~w25748 & w26070;
assign w26072 = ~w25724 & ~w25732;
assign w26073 = ~w25741 & ~w25747;
assign w26074 = ~w26072 & ~w26073;
assign w26075 = ~w26071 & w26074;
assign w26076 = ~w25733 & ~w26075;
assign w26077 = w23967 & ~w24134;
assign w26078 = ~w24135 & ~w26077;
assign w26079 = w3 & ~w22035;
assign w26080 = ~w21760 & w37524;
assign w26081 = ~w26079 & ~w26080;
assign w26082 = (w26081 & ~w24529) | (w26081 & w37525) | (~w24529 & w37525);
assign w26083 = (a_2 & ~w21771) | (a_2 & w34211) | (~w21771 & w34211);
assign w26084 = w26082 & ~w26083;
assign w26085 = (w24529 & w37526) | (w24529 & w37527) | (w37526 & w37527);
assign w26086 = ~w26084 & ~w26085;
assign w26087 = w23575 & w23598;
assign w26088 = ~w25722 & w37528;
assign w26089 = (w26087 & w25722) | (w26087 & w37529) | (w25722 & w37529);
assign w26090 = ~w26088 & ~w26089;
assign w26091 = w10835 & w21771;
assign w26092 = ~w21760 & w37530;
assign w26093 = ~w24498 & w37531;
assign w26094 = ~w26091 & ~w26092;
assign w26095 = ~w26093 & w26094;
assign w26096 = (a_2 & w22020) | (a_2 & w34211) | (w22020 & w34211);
assign w26097 = w26095 & ~w26096;
assign w26098 = (a_2 & w26093) | (a_2 & w37532) | (w26093 & w37532);
assign w26099 = ~w26097 & ~w26098;
assign w26100 = ~w26090 & ~w26099;
assign w26101 = (~w26100 & w26078) | (~w26100 & w37533) | (w26078 & w37533);
assign w26102 = ~w26076 & w26101;
assign w26103 = w26078 & w26086;
assign w26104 = w26090 & w26099;
assign w26105 = (w26104 & w26078) | (w26104 & w37534) | (w26078 & w37534);
assign w26106 = ~w26103 & ~w26105;
assign w26107 = ~w26102 & w26106;
assign w26108 = ~w25721 & ~w26107;
assign w26109 = ~w25712 & w25720;
assign w26110 = ~w24308 & ~w24309;
assign w26111 = w24518 & ~w24729;
assign w26112 = w26110 & ~w26111;
assign w26113 = ~w26110 & w26111;
assign w26114 = ~w26112 & ~w26113;
assign w26115 = w3 & w22039;
assign w26116 = w10835 & w22032;
assign w26117 = ~w26115 & ~w26116;
assign w26118 = (w26117 & ~w24962) | (w26117 & w37535) | (~w24962 & w37535);
assign w26119 = (a_2 & w22035) | (a_2 & w34211) | (w22035 & w34211);
assign w26120 = w26118 & ~w26119;
assign w26121 = (w24962 & w37536) | (w24962 & w37537) | (w37536 & w37537);
assign w26122 = ~w26120 & ~w26121;
assign w26123 = ~w26114 & w26122;
assign w26124 = ~w26109 & ~w26123;
assign w26125 = ~w26108 & w26124;
assign w26126 = w26114 & ~w26122;
assign w26127 = ~w24520 & ~w24729;
assign w26128 = w24725 & ~w24951;
assign w26129 = w26127 & ~w26128;
assign w26130 = ~w26127 & w26128;
assign w26131 = ~w26129 & ~w26130;
assign w26132 = w3 & ~w21757;
assign w26133 = w10835 & w22039;
assign w26134 = ~w26132 & ~w26133;
assign w26135 = (w26134 & w25205) | (w26134 & w37538) | (w25205 & w37538);
assign w26136 = (a_2 & ~w22032) | (a_2 & w34211) | (~w22032 & w34211);
assign w26137 = w26135 & ~w26136;
assign w26138 = (~w25205 & w37539) | (~w25205 & w37540) | (w37539 & w37540);
assign w26139 = ~w26137 & ~w26138;
assign w26140 = ~w26131 & ~w26139;
assign w26141 = ~w26126 & ~w26140;
assign w26142 = ~w26125 & w26141;
assign w26143 = w26131 & w26139;
assign w26144 = (~w32220 & w37541) | (~w32220 & w37542) | (w37541 & w37542);
assign w26145 = ~w24953 & ~w26144;
assign w26146 = ~w21736 & w37543;
assign w26147 = w10835 & ~w21757;
assign w26148 = ~w26146 & ~w26147;
assign w26149 = (w26148 & w25675) | (w26148 & w37544) | (w25675 & w37544);
assign w26150 = (a_2 & ~w22039) | (a_2 & w34211) | (~w22039 & w34211);
assign w26151 = w26149 & ~w26150;
assign w26152 = (~w25675 & w37545) | (~w25675 & w37546) | (w37545 & w37546);
assign w26153 = ~w26151 & ~w26152;
assign w26154 = w26145 & w26153;
assign w26155 = ~w26143 & ~w26154;
assign w26156 = ~w26142 & w26155;
assign w26157 = ~w26145 & ~w26153;
assign w26158 = w25175 & w25421;
assign w26159 = (~w24954 & w24731) | (~w24954 & w32221) | (w24731 & w32221);
assign w26160 = w26158 & ~w26159;
assign w26161 = ~w26158 & w26159;
assign w26162 = ~w26160 & ~w26161;
assign w26163 = w3 & w21752;
assign w26164 = ~w21736 & w37547;
assign w26165 = (~w22056 & ~w22053) | (~w22056 & w37548) | (~w22053 & w37548);
assign w26166 = ~w22057 & ~w26165;
assign w26167 = ~w26163 & ~w26164;
assign w26168 = (w26167 & ~w26166) | (w26167 & w37549) | (~w26166 & w37549);
assign w26169 = (a_2 & w21757) | (a_2 & w34211) | (w21757 & w34211);
assign w26170 = w26168 & ~w26169;
assign w26171 = (w26166 & w37550) | (w26166 & w37551) | (w37550 & w37551);
assign w26172 = ~w26170 & ~w26171;
assign w26173 = (~w26157 & w26162) | (~w26157 & w37552) | (w26162 & w37552);
assign w26174 = ~w26156 & w26173;
assign w26175 = w26162 & w26172;
assign w26176 = (~w26175 & w25696) | (~w26175 & w32222) | (w25696 & w32222);
assign w26177 = (~w25707 & w26174) | (~w25707 & w37553) | (w26174 & w37553);
assign w26178 = w25690 & w26177;
assign w26179 = ~w25690 & ~w26177;
assign w26180 = ~w26178 & ~w26179;
assign w26181 = ~w25688 & ~w26178;
assign w26182 = w25455 & ~w25683;
assign w26183 = w25471 & w25627;
assign w26184 = ~w25471 & w25631;
assign w26185 = ~w26183 & ~w26184;
assign w26186 = ~w25647 & ~w26185;
assign w26187 = ~w25633 & w25647;
assign w26188 = ~w26186 & ~w26187;
assign w26189 = w25471 & w25638;
assign w26190 = ~w25471 & w25642;
assign w26191 = ~w26189 & ~w26190;
assign w26192 = ~w25647 & ~w26191;
assign w26193 = ~w25644 & w25647;
assign w26194 = ~w26192 & ~w26193;
assign w26195 = ~w26188 & ~w26194;
assign w26196 = w25460 & w26195;
assign w26197 = (w25656 & w25460) | (w25656 & w32588) | (w25460 & w32588);
assign w26198 = ~w26196 & w26197;
assign w26199 = (~w26198 & w25457) | (~w26198 & w32223) | (w25457 & w32223);
assign w26200 = w25437 & ~w26194;
assign w26201 = ~w26188 & ~w26200;
assign w26202 = w25438 & ~w26188;
assign w26203 = ~w25182 & w26202;
assign w26204 = ~w26201 & ~w26203;
assign w26205 = w10033 & w26166;
assign w26206 = ~w21736 & w37554;
assign w26207 = w9786 & ~w21757;
assign w26208 = w9788 & w21752;
assign w26209 = ~w26206 & ~w26207;
assign w26210 = ~w26208 & w26209;
assign w26211 = a_5 & ~w26210;
assign w26212 = ~a_5 & w26210;
assign w26213 = (w26212 & ~w26166) | (w26212 & w37555) | (~w26166 & w37555);
assign w26214 = ~w26205 & ~w26211;
assign w26215 = ~w26213 & w26214;
assign w26216 = ~w26204 & w26215;
assign w26217 = w26204 & ~w26215;
assign w26218 = ~w26216 & ~w26217;
assign w26219 = w8295 & w22039;
assign w26220 = w8277 & ~w22035;
assign w26221 = w8298 & w22032;
assign w26222 = ~w26220 & ~w26221;
assign w26223 = ~w26219 & w26222;
assign w26224 = (w26223 & ~w24962) | (w26223 & w37556) | (~w24962 & w37556);
assign w26225 = ~a_8 & w26224;
assign w26226 = (w24962 & w37557) | (w24962 & w37558) | (w37557 & w37558);
assign w26227 = ~w26225 & ~w26226;
assign w26228 = w25471 & ~w25603;
assign w26229 = ~w25471 & w25603;
assign w26230 = ~w26228 & ~w26229;
assign w26231 = w25612 & ~w26230;
assign w26232 = ~w25612 & w26230;
assign w26233 = w25647 & ~w26232;
assign w26234 = (~w26231 & ~w25647) | (~w26231 & w37559) | (~w25647 & w37559);
assign w26235 = w7489 & w21771;
assign w26236 = ~w21760 & w37560;
assign w26237 = w7192 & ~w22020;
assign w26238 = ~w24498 & w37561;
assign w26239 = ~w26236 & ~w26237;
assign w26240 = ~w26235 & w26239;
assign w26241 = ~w26238 & w26240;
assign w26242 = ~w26238 & w37562;
assign w26243 = a_11 & ~w26241;
assign w26244 = ~w26242 & ~w26243;
assign w26245 = ~w25226 & ~w25470;
assign w26246 = w25465 & w25602;
assign w26247 = ~w26245 & w26246;
assign w26248 = ~w25591 & ~w26247;
assign w26249 = w6996 & w22014;
assign w26250 = w6446 & ~w21992;
assign w26251 = w6998 & w22007;
assign w26252 = w6447 & w23398;
assign w26253 = ~w26250 & ~w26251;
assign w26254 = ~w26249 & w26253;
assign w26255 = ~w26252 & w26254;
assign w26256 = a_14 & ~w26255;
assign w26257 = ~a_14 & w26255;
assign w26258 = ~w26256 & ~w26257;
assign w26259 = w25560 & ~w25569;
assign w26260 = w25558 & w25569;
assign w26261 = w25557 & w25569;
assign w26262 = ~w25476 & w26261;
assign w26263 = ~w25333 & ~w26262;
assign w26264 = ~w26260 & w26263;
assign w26265 = ~w25473 & w26264;
assign w26266 = ~w26259 & ~w26265;
assign w26267 = (~w25319 & w25536) | (~w25319 & w32224) | (w25536 & w32224);
assign w26268 = ~w25550 & w26267;
assign w26269 = ~w25546 & ~w26268;
assign w26270 = w4666 & w21892;
assign w26271 = ~w518 & w21894;
assign w26272 = w4638 & w21901;
assign w26273 = ~w26270 & ~w26271;
assign w26274 = ~w26272 & w26273;
assign w26275 = (w22096 & w32589) | (w22096 & w32590) | (w32589 & w32590);
assign w26276 = (~w22096 & w32591) | (~w22096 & w32592) | (w32591 & w32592);
assign w26277 = ~w26275 & ~w26276;
assign w26278 = w25493 & w32226;
assign w26279 = (~a_29 & ~w25493) | (~a_29 & w32227) | (~w25493 & w32227);
assign w26280 = ~w26278 & ~w26279;
assign w26281 = ~w25520 & ~w25522;
assign w26282 = w25520 & w25522;
assign w26283 = ~w26281 & ~w26282;
assign w26284 = ~w26280 & ~w26283;
assign w26285 = (~w26284 & ~w25532) | (~w26284 & w32228) | (~w25532 & w32228);
assign w26286 = w4070 & w22107;
assign w26287 = w21873 & w32229;
assign w26288 = w4070 & ~w21854;
assign w26289 = ~w21787 & w26288;
assign w26290 = ~w26287 & ~w26289;
assign w26291 = ~w22105 & ~w26290;
assign w26292 = w3957 & ~w21839;
assign w26293 = w4068 & w21854;
assign w26294 = w4446 & w21787;
assign w26295 = ~w26292 & ~w26293;
assign w26296 = ~w26294 & w26295;
assign w26297 = ~w26291 & w26296;
assign w26298 = ~w26286 & w26297;
assign w26299 = ~w25519 & ~w25522;
assign w26300 = ~w25517 & ~w26299;
assign w26301 = w668 & ~w21224;
assign w26302 = w21207 & w26301;
assign w26303 = w1327 & ~w21800;
assign w26304 = w21799 & w26303;
assign w26305 = w1327 & w21800;
assign w26306 = ~w21799 & w26305;
assign w26307 = w668 & w21224;
assign w26308 = ~w21207 & w26307;
assign w26309 = ~w21796 & w32230;
assign w26310 = ~w26304 & ~w26306;
assign w26311 = ~w26302 & w26310;
assign w26312 = ~w26308 & ~w26309;
assign w26313 = w26311 & w26312;
assign w26314 = w1478 & ~w21224;
assign w26315 = w21827 & ~w26314;
assign w26316 = w1478 & w21224;
assign w26317 = ~w21827 & ~w26316;
assign w26318 = ~w26315 & ~w26317;
assign w26319 = w26313 & ~w26318;
assign w26320 = w21824 & ~w26319;
assign w26321 = w21827 & ~w26316;
assign w26322 = ~w21827 & ~w26314;
assign w26323 = ~w26321 & ~w26322;
assign w26324 = w26313 & ~w26323;
assign w26325 = ~w21824 & ~w26324;
assign w26326 = ~w26320 & ~w26325;
assign w26327 = ~w216 & ~w741;
assign w26328 = w628 & w26327;
assign w26329 = w819 & w2404;
assign w26330 = w26328 & w26329;
assign w26331 = w1716 & w2037;
assign w26332 = w3026 & w3602;
assign w26333 = w5171 & w26332;
assign w26334 = w26330 & w26331;
assign w26335 = w13451 & w26334;
assign w26336 = w4392 & w26333;
assign w26337 = w26335 & w26336;
assign w26338 = w4863 & w26337;
assign w26339 = w13534 & w26338;
assign w26340 = ~w26326 & ~w26339;
assign w26341 = w26326 & w26339;
assign w26342 = ~w26340 & ~w26341;
assign w26343 = w26300 & w26342;
assign w26344 = ~w26300 & ~w26342;
assign w26345 = ~w26343 & ~w26344;
assign w26346 = a_29 & ~w26345;
assign w26347 = w26298 & w26346;
assign w26348 = ~a_29 & ~w26345;
assign w26349 = ~w26298 & w26348;
assign w26350 = ~w26347 & ~w26349;
assign w26351 = ~a_29 & ~w26298;
assign w26352 = a_29 & w26298;
assign w26353 = w26345 & ~w26351;
assign w26354 = ~w26352 & w26353;
assign w26355 = w26350 & ~w26354;
assign w26356 = w26285 & ~w26355;
assign w26357 = ~w26285 & w26355;
assign w26358 = ~w26356 & ~w26357;
assign w26359 = w26277 & w26358;
assign w26360 = ~w26277 & ~w26358;
assign w26361 = ~w26359 & ~w26360;
assign w26362 = ~w26269 & w26361;
assign w26363 = w26269 & ~w26361;
assign w26364 = ~w26362 & ~w26363;
assign w26365 = w7961 & w22905;
assign w26366 = w5016 & ~w21910;
assign w26367 = w5080 & w21921;
assign w26368 = w5286 & w21951;
assign w26369 = ~w26366 & ~w26367;
assign w26370 = ~w26368 & w26369;
assign w26371 = a_23 & ~w26370;
assign w26372 = w5017 & w22905;
assign w26373 = ~a_23 & w26370;
assign w26374 = ~w26372 & w26373;
assign w26375 = ~w26365 & ~w26371;
assign w26376 = ~w26374 & w26375;
assign w26377 = w26364 & w26376;
assign w26378 = ~w26364 & ~w26376;
assign w26379 = ~w26377 & ~w26378;
assign w26380 = (~w25325 & ~w25554) | (~w25325 & w32593) | (~w25554 & w32593);
assign w26381 = ~w25475 & w26380;
assign w26382 = ~w25555 & ~w26381;
assign w26383 = w26379 & w26382;
assign w26384 = ~w26379 & ~w26382;
assign w26385 = ~w26383 & ~w26384;
assign w26386 = w5308 & ~w21945;
assign w26387 = w5816 & w21934;
assign w26388 = w5818 & ~w21940;
assign w26389 = w5309 & w23310;
assign w26390 = ~w26386 & ~w26387;
assign w26391 = ~w26388 & w26390;
assign w26392 = ~w26389 & w26391;
assign w26393 = a_20 & ~w26392;
assign w26394 = ~a_20 & w26392;
assign w26395 = ~w26393 & ~w26394;
assign w26396 = w6304 & w21985;
assign w26397 = w6059 & ~w21968;
assign w26398 = w6061 & ~w21973;
assign w26399 = w6063 & w23553;
assign w26400 = ~w26396 & ~w26397;
assign w26401 = ~w26398 & w26400;
assign w26402 = ~w26399 & w26401;
assign w26403 = a_17 & ~w26402;
assign w26404 = ~a_17 & w26402;
assign w26405 = ~w26403 & ~w26404;
assign w26406 = ~w26395 & w26405;
assign w26407 = w26395 & ~w26405;
assign w26408 = ~w26406 & ~w26407;
assign w26409 = w26385 & ~w26408;
assign w26410 = ~w26385 & w26408;
assign w26411 = ~w26409 & ~w26410;
assign w26412 = w26266 & w26411;
assign w26413 = ~w26266 & ~w26411;
assign w26414 = ~w26412 & ~w26413;
assign w26415 = w26258 & ~w26414;
assign w26416 = ~w26258 & w26414;
assign w26417 = ~w26415 & ~w26416;
assign w26418 = w26248 & w26417;
assign w26419 = ~w26248 & ~w26417;
assign w26420 = ~w26418 & ~w26419;
assign w26421 = w26244 & ~w26420;
assign w26422 = ~w26244 & w26420;
assign w26423 = ~w26421 & ~w26422;
assign w26424 = w26234 & w26423;
assign w26425 = ~w26234 & ~w26423;
assign w26426 = ~w26424 & ~w26425;
assign w26427 = w26227 & w26426;
assign w26428 = ~w26227 & ~w26426;
assign w26429 = ~w26427 & ~w26428;
assign w26430 = w26218 & ~w26429;
assign w26431 = ~w26218 & w26429;
assign w26432 = ~w26430 & ~w26431;
assign w26433 = w26199 & w26432;
assign w26434 = ~w26199 & ~w26432;
assign w26435 = ~w26433 & ~w26434;
assign w26436 = ~w25682 & w26435;
assign w26437 = ~w26182 & w26436;
assign w26438 = (~w25682 & ~w25455) | (~w25682 & w32231) | (~w25455 & w32231);
assign w26439 = ~w26435 & ~w26438;
assign w26440 = ~w26437 & ~w26439;
assign w26441 = ~w13251 & ~w13255;
assign w26442 = ~w13232 & ~w13241;
assign w26443 = ~w13225 & ~w13228;
assign w26444 = w1258 & w1694;
assign w26445 = w3932 & w26444;
assign w26446 = w13219 & w26445;
assign w26447 = w26443 & ~w26446;
assign w26448 = ~w26443 & w26446;
assign w26449 = ~w26447 & ~w26448;
assign w26450 = w668 & w13177;
assign w26451 = w1327 & w13180;
assign w26452 = w1478 & w13207;
assign w26453 = ~w13236 & ~w26451;
assign w26454 = ~w26450 & w26453;
assign w26455 = ~w26452 & w26454;
assign w26456 = w26449 & ~w26455;
assign w26457 = ~w26449 & w26455;
assign w26458 = ~w26456 & ~w26457;
assign w26459 = w26442 & ~w26458;
assign w26460 = ~w26442 & w26458;
assign w26461 = ~w26459 & ~w26460;
assign w26462 = a_29 & ~w3956;
assign w26463 = ~a_26 & w7;
assign w26464 = ~w26462 & ~w26463;
assign w26465 = w26461 & w26464;
assign w26466 = ~w26461 & ~w26464;
assign w26467 = ~w26465 & ~w26466;
assign w26468 = w26441 & ~w26467;
assign w26469 = ~w26441 & w26467;
assign w26470 = ~w26468 & ~w26469;
assign w26471 = ~w13278 & w26470;
assign w26472 = ~w21742 & w26471;
assign w26473 = w13278 & ~w26470;
assign w26474 = ~w26472 & ~w26473;
assign w26475 = w21742 & ~w26470;
assign w26476 = w26474 & ~w26475;
assign w26477 = w3 & w26476;
assign w26478 = w10835 & ~w21743;
assign w26479 = ~w21743 & w26476;
assign w26480 = ~w21741 & ~w26474;
assign w26481 = ~w21749 & ~w26480;
assign w26482 = w22062 & w26481;
assign w26483 = ~w21748 & ~w26479;
assign w26484 = ~w26482 & w26483;
assign w26485 = ~w26479 & ~w26484;
assign w26486 = ~w21746 & w26479;
assign w26487 = ~w26480 & ~w26486;
assign w26488 = ~w22063 & ~w26487;
assign w26489 = ~w26485 & ~w26488;
assign w26490 = w10837 & w26489;
assign w26491 = ~w26477 & ~w26478;
assign w26492 = ~w26490 & w26491;
assign w26493 = w10839 & w21746;
assign w26494 = a_2 & ~w26493;
assign w26495 = w26492 & ~w26494;
assign w26496 = a_2 & ~w26492;
assign w26497 = ~w26495 & ~w26496;
assign w26498 = ~w26440 & ~w26497;
assign w26499 = w26440 & w26497;
assign w26500 = ~w26498 & ~w26499;
assign w26501 = w26181 & ~w26500;
assign w26502 = ~w26181 & w26500;
assign w26503 = ~w26501 & ~w26502;
assign w26504 = w26180 & w26503;
assign w26505 = ~w26180 & ~w26503;
assign w26506 = ~w26504 & ~w26505;
assign w26507 = ~w25688 & ~w26499;
assign w26508 = ~w26178 & w26507;
assign w26509 = w26216 & ~w26429;
assign w26510 = w26204 & ~w26428;
assign w26511 = (w26215 & ~w26426) | (w26215 & w32594) | (~w26426 & w32594);
assign w26512 = w26510 & w26511;
assign w26513 = ~w26509 & ~w26512;
assign w26514 = w26215 & w26513;
assign w26515 = ~w26199 & w26514;
assign w26516 = w26199 & ~w26513;
assign w26517 = ~w26515 & ~w26516;
assign w26518 = (w26517 & w26182) | (w26517 & w32595) | (w26182 & w32595);
assign w26519 = w26204 & w26427;
assign w26520 = w26227 & ~w26426;
assign w26521 = ~w26204 & w26520;
assign w26522 = ~w26519 & ~w26521;
assign w26523 = ~w26198 & w26522;
assign w26524 = ~w25668 & w26523;
assign w26525 = ~w26227 & w26426;
assign w26526 = ~w26204 & ~w26525;
assign w26527 = ~w26510 & ~w26526;
assign w26528 = (~w26527 & w25668) | (~w26527 & w32232) | (w25668 & w32232);
assign w26529 = ~w26204 & w26426;
assign w26530 = w26244 & ~w26426;
assign w26531 = ~w26529 & ~w26530;
assign w26532 = w9788 & w21746;
assign w26533 = w9786 & w21755;
assign w26534 = w9780 & w21752;
assign w26535 = w9790 & ~w25700;
assign w26536 = ~w26533 & ~w26534;
assign w26537 = ~w26532 & w26536;
assign w26538 = ~w26535 & w26537;
assign w26539 = ~a_5 & w26538;
assign w26540 = a_5 & ~w26538;
assign w26541 = ~w26539 & ~w26540;
assign w26542 = w26258 & w26414;
assign w26543 = w26248 & w26542;
assign w26544 = ~w26248 & w26415;
assign w26545 = ~w26543 & ~w26544;
assign w26546 = ~w26231 & w26545;
assign w26547 = ~w26233 & w26546;
assign w26548 = ~w26258 & ~w26420;
assign w26549 = ~w26547 & ~w26548;
assign w26550 = ~w25591 & ~w26414;
assign w26551 = ~w26247 & w26550;
assign w26552 = w26405 & w26414;
assign w26553 = ~w26551 & ~w26552;
assign w26554 = ~w25555 & ~w26377;
assign w26555 = (~w26378 & ~w26554) | (~w26378 & w32596) | (~w26554 & w32596);
assign w26556 = w5816 & ~w21968;
assign w26557 = w5308 & ~w21940;
assign w26558 = w5818 & w21934;
assign w26559 = w5309 & ~w23366;
assign w26560 = ~w26557 & ~w26558;
assign w26561 = ~w26556 & w26560;
assign w26562 = ~w26559 & w26561;
assign w26563 = a_20 & w26562;
assign w26564 = ~a_20 & ~w26562;
assign w26565 = ~w26563 & ~w26564;
assign w26566 = ~w26359 & ~w26362;
assign w26567 = ~w26284 & w26350;
assign w26568 = (~w26354 & ~w26567) | (~w26354 & w32597) | (~w26567 & w32597);
assign w26569 = w4068 & w21787;
assign w26570 = w3957 & w21854;
assign w26571 = w4446 & w21894;
assign w26572 = ~w26569 & ~w26570;
assign w26573 = ~w26571 & w26572;
assign w26574 = (w26573 & w23079) | (w26573 & w32233) | (w23079 & w32233);
assign w26575 = w1478 & w22278;
assign w26576 = w1327 & w21833;
assign w26577 = w1399 & ~w21803;
assign w26578 = w668 & ~w21839;
assign w26579 = ~w26576 & ~w26577;
assign w26580 = ~w26578 & w26579;
assign w26581 = (w26580 & ~w22278) | (w26580 & w32598) | (~w22278 & w32598);
assign w26582 = w63 & w3517;
assign w26583 = ~w195 & ~w475;
assign w26584 = ~w568 & ~w590;
assign w26585 = ~w834 & w26584;
assign w26586 = w158 & w934;
assign w26587 = w2454 & w5187;
assign w26588 = w13985 & w26583;
assign w26589 = w26587 & w26588;
assign w26590 = w26585 & w26586;
assign w26591 = w2808 & w3767;
assign w26592 = w26582 & w26591;
assign w26593 = w26589 & w26590;
assign w26594 = w6709 & w26593;
assign w26595 = w6610 & w26592;
assign w26596 = w26594 & w26595;
assign w26597 = w2795 & w14029;
assign w26598 = w26596 & w26597;
assign w26599 = w1794 & w26598;
assign w26600 = ~w26581 & ~w26599;
assign w26601 = w26580 & w26599;
assign w26602 = ~w26575 & w26601;
assign w26603 = ~w26600 & ~w26602;
assign w26604 = ~w26341 & ~w26343;
assign w26605 = (a_29 & w26343) | (a_29 & w32234) | (w26343 & w32234);
assign w26606 = ~w26343 & w32235;
assign w26607 = ~w26605 & ~w26606;
assign w26608 = w26603 & ~w26607;
assign w26609 = ~w26603 & w26607;
assign w26610 = ~w26608 & ~w26609;
assign w26611 = w26574 & w26610;
assign w26612 = ~w26574 & ~w26610;
assign w26613 = ~w26611 & ~w26612;
assign w26614 = ~w26568 & w26613;
assign w26615 = w26568 & ~w26613;
assign w26616 = ~w26614 & ~w26615;
assign w26617 = w1226 & ~w22580;
assign w26618 = ~w518 & w21901;
assign w26619 = w4638 & w21892;
assign w26620 = w4666 & ~w21910;
assign w26621 = ~w26618 & ~w26619;
assign w26622 = ~w26620 & w26621;
assign w26623 = ~a_26 & w26622;
assign w26624 = ~w26617 & w26623;
assign w26625 = w4403 & ~w22580;
assign w26626 = a_26 & ~w26622;
assign w26627 = ~w26625 & ~w26626;
assign w26628 = ~w26624 & w26627;
assign w26629 = w26616 & w26628;
assign w26630 = ~w26616 & ~w26628;
assign w26631 = ~w26629 & ~w26630;
assign w26632 = w5016 & w21921;
assign w26633 = w5080 & w21951;
assign w26634 = w5286 & ~w21945;
assign w26635 = ~w26632 & ~w26633;
assign w26636 = ~w26634 & w26635;
assign w26637 = (w26636 & ~w22083) | (w26636 & w32236) | (~w22083 & w32236);
assign w26638 = ~a_23 & w26637;
assign w26639 = a_23 & ~w26637;
assign w26640 = ~w26638 & ~w26639;
assign w26641 = w26631 & ~w26640;
assign w26642 = ~w26631 & w26640;
assign w26643 = ~w26641 & ~w26642;
assign w26644 = w26566 & w26643;
assign w26645 = ~w26566 & ~w26643;
assign w26646 = ~w26644 & ~w26645;
assign w26647 = w26565 & w26646;
assign w26648 = w26555 & w26647;
assign w26649 = w26565 & ~w26646;
assign w26650 = ~w26555 & w26649;
assign w26651 = ~w26648 & ~w26650;
assign w26652 = ~w26565 & ~w26646;
assign w26653 = w26555 & w26652;
assign w26654 = ~w26565 & w26646;
assign w26655 = ~w26555 & w26654;
assign w26656 = ~w26653 & ~w26655;
assign w26657 = w26651 & w26656;
assign w26658 = w6304 & ~w21992;
assign w26659 = w6061 & w21985;
assign w26660 = w6059 & ~w21973;
assign w26661 = w6063 & ~w23930;
assign w26662 = ~w26659 & ~w26660;
assign w26663 = ~w26658 & w26662;
assign w26664 = ~w26661 & w26663;
assign w26665 = a_17 & ~w26664;
assign w26666 = ~a_17 & w26664;
assign w26667 = ~w26665 & ~w26666;
assign w26668 = ~w26657 & ~w26667;
assign w26669 = w26657 & w26667;
assign w26670 = ~w26668 & ~w26669;
assign w26671 = ~w26379 & ~w26395;
assign w26672 = w26382 & w26671;
assign w26673 = w26379 & ~w26395;
assign w26674 = ~w26382 & w26673;
assign w26675 = ~w26672 & ~w26674;
assign w26676 = ~w26259 & w26675;
assign w26677 = ~w26265 & w26676;
assign w26678 = ~w26385 & w26395;
assign w26679 = ~w26677 & ~w26678;
assign w26680 = w8564 & w24122;
assign w26681 = w8592 & w24122;
assign w26682 = w6998 & w22014;
assign w26683 = w6446 & w22007;
assign w26684 = w6996 & ~w22020;
assign w26685 = ~w26682 & ~w26683;
assign w26686 = ~w26684 & w26685;
assign w26687 = a_14 & w26686;
assign w26688 = ~a_14 & ~w26686;
assign w26689 = ~w26687 & ~w26688;
assign w26690 = ~w26681 & w26689;
assign w26691 = ~w26680 & ~w26690;
assign w26692 = ~w26677 & w32599;
assign w26693 = (w26691 & w26677) | (w26691 & w32600) | (w26677 & w32600);
assign w26694 = ~w26692 & ~w26693;
assign w26695 = w26670 & ~w26694;
assign w26696 = ~w26670 & w26694;
assign w26697 = ~w26695 & ~w26696;
assign w26698 = ~w26553 & w26697;
assign w26699 = w26553 & ~w26697;
assign w26700 = ~w26698 & ~w26699;
assign w26701 = w7192 & w21771;
assign w26702 = w7489 & w21762;
assign w26703 = w7511 & ~w22035;
assign w26704 = w7193 & w24529;
assign w26705 = ~w26702 & ~w26703;
assign w26706 = ~w26701 & w26705;
assign w26707 = ~w26704 & w26706;
assign w26708 = a_11 & ~w26707;
assign w26709 = ~a_11 & w26707;
assign w26710 = ~w26708 & ~w26709;
assign w26711 = w9456 & ~w25205;
assign w26712 = w8298 & w22039;
assign w26713 = w8277 & w22032;
assign w26714 = w8295 & ~w21757;
assign w26715 = ~w26712 & ~w26713;
assign w26716 = ~w26714 & w26715;
assign w26717 = a_8 & ~w26716;
assign w26718 = w8278 & ~w25205;
assign w26719 = ~a_8 & w26716;
assign w26720 = ~w26718 & w26719;
assign w26721 = ~w26711 & ~w26717;
assign w26722 = ~w26720 & w26721;
assign w26723 = w26710 & ~w26722;
assign w26724 = ~w26710 & w26722;
assign w26725 = ~w26723 & ~w26724;
assign w26726 = w26700 & ~w26725;
assign w26727 = ~w26700 & w26725;
assign w26728 = ~w26726 & ~w26727;
assign w26729 = w26549 & w26728;
assign w26730 = ~w26549 & ~w26728;
assign w26731 = ~w26729 & ~w26730;
assign w26732 = w26541 & ~w26731;
assign w26733 = ~w26541 & w26731;
assign w26734 = ~w26732 & ~w26733;
assign w26735 = w26531 & w26734;
assign w26736 = ~w26531 & ~w26734;
assign w26737 = ~w26735 & ~w26736;
assign w26738 = w26528 & ~w26737;
assign w26739 = ~w26528 & w26737;
assign w26740 = ~w26738 & ~w26739;
assign w26741 = ~w26469 & ~w26472;
assign w26742 = ~w26460 & ~w26465;
assign w26743 = ~w26448 & ~w26456;
assign w26744 = w3887 & w3934;
assign w26745 = w26446 & ~w26744;
assign w26746 = ~w26446 & w26744;
assign w26747 = ~w26745 & ~w26746;
assign w26748 = ~w26743 & w26747;
assign w26749 = w26743 & ~w26747;
assign w26750 = ~w26748 & ~w26749;
assign w26751 = w1399 & w13180;
assign w26752 = w1478 & ~w13264;
assign w26753 = ~w667 & ~w26751;
assign w26754 = ~w26752 & w26753;
assign w26755 = w26464 & w26754;
assign w26756 = ~w26464 & ~w26754;
assign w26757 = ~w26755 & ~w26756;
assign w26758 = w26750 & ~w26757;
assign w26759 = ~w26750 & w26757;
assign w26760 = ~w26758 & ~w26759;
assign w26761 = ~w26742 & w26760;
assign w26762 = w26742 & ~w26760;
assign w26763 = ~w26761 & ~w26762;
assign w26764 = w26741 & ~w26763;
assign w26765 = ~w26741 & w26763;
assign w26766 = ~w26764 & ~w26765;
assign w26767 = w3 & w26766;
assign w26768 = w10835 & w26476;
assign w26769 = ~w26476 & ~w26766;
assign w26770 = w26476 & w26766;
assign w26771 = ~w26769 & ~w26770;
assign w26772 = ~w26484 & ~w26771;
assign w26773 = w26484 & w26771;
assign w26774 = ~w26772 & ~w26773;
assign w26775 = w10837 & ~w26774;
assign w26776 = ~w26767 & ~w26768;
assign w26777 = ~w26775 & w26776;
assign w26778 = w10839 & ~w21743;
assign w26779 = a_2 & ~w26778;
assign w26780 = w26777 & ~w26779;
assign w26781 = a_2 & ~w26777;
assign w26782 = ~w26780 & ~w26781;
assign w26783 = w26740 & w26782;
assign w26784 = ~w26740 & ~w26782;
assign w26785 = ~w26783 & ~w26784;
assign w26786 = w26518 & w26785;
assign w26787 = ~w26518 & ~w26785;
assign w26788 = ~w26786 & ~w26787;
assign w26789 = ~w26498 & ~w26788;
assign w26790 = ~w26508 & w26789;
assign w26791 = (w26788 & w26508) | (w26788 & w32601) | (w26508 & w32601);
assign w26792 = ~w26790 & ~w26791;
assign w26793 = w26504 & w26792;
assign w26794 = ~w26504 & ~w26792;
assign w26795 = ~w26793 & ~w26794;
assign w26796 = w26782 & w26788;
assign w26797 = (~w26796 & w26508) | (~w26796 & w32602) | (w26508 & w32602);
assign w26798 = ~w26541 & ~w26740;
assign w26799 = w26528 & w32603;
assign w26800 = w26541 & w26737;
assign w26801 = ~w26528 & w26800;
assign w26802 = w26517 & ~w26801;
assign w26803 = ~w26799 & w26802;
assign w26804 = (~w26798 & w26437) | (~w26798 & w32237) | (w26437 & w32237);
assign w26805 = ~w26531 & ~w26731;
assign w26806 = ~w26530 & w26731;
assign w26807 = ~w26529 & w26806;
assign w26808 = ~w26527 & ~w26807;
assign w26809 = ~w26805 & w26808;
assign w26810 = ~w26524 & w26809;
assign w26811 = ~w26805 & ~w26807;
assign w26812 = w26722 & ~w26811;
assign w26813 = ~w26810 & ~w26812;
assign w26814 = w26700 & w26710;
assign w26815 = w26549 & w26814;
assign w26816 = ~w26700 & w26710;
assign w26817 = ~w26549 & w26816;
assign w26818 = ~w26815 & ~w26817;
assign w26819 = ~w26530 & w26818;
assign w26820 = ~w26529 & w26819;
assign w26821 = ~w26549 & ~w26700;
assign w26822 = w26549 & w26700;
assign w26823 = ~w26710 & ~w26821;
assign w26824 = ~w26822 & w26823;
assign w26825 = ~w26820 & ~w26824;
assign w26826 = w26657 & ~w26667;
assign w26827 = ~w26679 & w26826;
assign w26828 = w26668 & w26679;
assign w26829 = ~w26827 & ~w26828;
assign w26830 = ~w26657 & w26667;
assign w26831 = ~w26679 & w26830;
assign w26832 = w26669 & w26679;
assign w26833 = ~w26831 & ~w26832;
assign w26834 = w26829 & w26833;
assign w26835 = w26553 & ~w26834;
assign w26836 = ~w26553 & w26834;
assign w26837 = ~w26835 & ~w26836;
assign w26838 = ~w26691 & ~w26837;
assign w26839 = (w26691 & w26553) | (w26691 & w32604) | (w26553 & w32604);
assign w26840 = ~w26835 & w26839;
assign w26841 = (~w26840 & ~w26549) | (~w26840 & w32605) | (~w26549 & w32605);
assign w26842 = ~w26552 & w26833;
assign w26843 = ~w26551 & w26842;
assign w26844 = (w26829 & ~w26842) | (w26829 & w32238) | (~w26842 & w32238);
assign w26845 = w8564 & w24295;
assign w26846 = w8592 & w24295;
assign w26847 = w6998 & ~w22020;
assign w26848 = w6446 & w22014;
assign w26849 = w6996 & w21771;
assign w26850 = ~w26847 & ~w26848;
assign w26851 = ~w26849 & w26850;
assign w26852 = a_14 & w26851;
assign w26853 = ~a_14 & ~w26851;
assign w26854 = ~w26852 & ~w26853;
assign w26855 = ~w26846 & w26854;
assign w26856 = ~w26845 & ~w26855;
assign w26857 = w26656 & ~w26678;
assign w26858 = (w26651 & ~w26857) | (w26651 & w32239) | (~w26857 & w32239);
assign w26859 = w6304 & w22007;
assign w26860 = w6061 & ~w21992;
assign w26861 = w6059 & w21985;
assign w26862 = w6063 & w23580;
assign w26863 = ~w26860 & ~w26861;
assign w26864 = ~w26859 & w26863;
assign w26865 = ~w26862 & w26864;
assign w26866 = a_17 & ~w26865;
assign w26867 = ~a_17 & w26865;
assign w26868 = ~w26866 & ~w26867;
assign w26869 = w26640 & ~w26646;
assign w26870 = w26555 & w26646;
assign w26871 = ~w26869 & ~w26870;
assign w26872 = w4666 & w21921;
assign w26873 = ~w518 & w21892;
assign w26874 = w4638 & ~w21910;
assign w26875 = w1226 & w22664;
assign w26876 = ~w26872 & ~w26873;
assign w26877 = ~w26874 & w26876;
assign w26878 = ~w26875 & w26877;
assign w26879 = a_26 & w26878;
assign w26880 = ~a_26 & ~w26878;
assign w26881 = ~w26879 & ~w26880;
assign w26882 = (~w23079 & w32606) | (~w23079 & w32607) | (w32606 & w32607);
assign w26883 = (w23079 & w32608) | (w23079 & w32609) | (w32608 & w32609);
assign w26884 = ~w26882 & ~w26883;
assign w26885 = ~w26603 & ~w26604;
assign w26886 = w26603 & w26604;
assign w26887 = ~w26885 & ~w26886;
assign w26888 = ~w26884 & w26887;
assign w26889 = (~w26888 & ~w26568) | (~w26888 & w32240) | (~w26568 & w32240);
assign w26890 = w4446 & w21901;
assign w26891 = w3957 & w21787;
assign w26892 = w4068 & w21894;
assign w26893 = ~w26890 & ~w26891;
assign w26894 = ~w26892 & w26893;
assign w26895 = ~a_29 & w26894;
assign w26896 = (w26895 & ~w22555) | (w26895 & w32241) | (~w22555 & w32241);
assign w26897 = a_29 & ~w26894;
assign w26898 = (~w26897 & ~w22555) | (~w26897 & w32242) | (~w22555 & w32242);
assign w26899 = ~w26896 & w26898;
assign w26900 = (~w26600 & ~w26604) | (~w26600 & w32610) | (~w26604 & w32610);
assign w26901 = w668 & w21854;
assign w26902 = w1399 & w21833;
assign w26903 = w1327 & ~w21839;
assign w26904 = ~w26901 & ~w26902;
assign w26905 = ~w26903 & w26904;
assign w26906 = (w26905 & w23698) | (w26905 & w32611) | (w23698 & w32611);
assign w26907 = w320 & w1343;
assign w26908 = w1454 & w1588;
assign w26909 = w1954 & w14055;
assign w26910 = w26908 & w26909;
assign w26911 = w344 & w26907;
assign w26912 = w1986 & w3867;
assign w26913 = w6643 & w13562;
assign w26914 = w26912 & w26913;
assign w26915 = w26910 & w26911;
assign w26916 = w3432 & w26915;
assign w26917 = w4352 & w26914;
assign w26918 = w26916 & w26917;
assign w26919 = w3180 & w26918;
assign w26920 = w4384 & w26919;
assign w26921 = ~w26906 & ~w26920;
assign w26922 = w26906 & w26920;
assign w26923 = ~w26921 & ~w26922;
assign w26924 = w26900 & ~w26923;
assign w26925 = ~w26900 & w26923;
assign w26926 = ~w26924 & ~w26925;
assign w26927 = w26899 & w26926;
assign w26928 = ~w26899 & ~w26926;
assign w26929 = ~w26927 & ~w26928;
assign w26930 = w26889 & w26929;
assign w26931 = ~w26889 & ~w26929;
assign w26932 = ~w26930 & ~w26931;
assign w26933 = ~w26881 & ~w26932;
assign w26934 = w26881 & w26932;
assign w26935 = ~w26933 & ~w26934;
assign w26936 = (~w26359 & ~w26616) | (~w26359 & w32243) | (~w26616 & w32243);
assign w26937 = ~w26362 & w26936;
assign w26938 = ~w26630 & ~w26937;
assign w26939 = w26935 & w26938;
assign w26940 = ~w26935 & ~w26938;
assign w26941 = ~w26939 & ~w26940;
assign w26942 = w5080 & ~w21945;
assign w26943 = w5016 & w21951;
assign w26944 = w5286 & ~w21940;
assign w26945 = w5017 & w23032;
assign w26946 = ~w26942 & ~w26943;
assign w26947 = ~w26944 & w26946;
assign w26948 = ~w26945 & w26947;
assign w26949 = a_23 & ~w26948;
assign w26950 = ~a_23 & w26948;
assign w26951 = ~w26949 & ~w26950;
assign w26952 = w8311 & ~w22930;
assign w26953 = w8339 & ~w22930;
assign w26954 = w5818 & ~w21968;
assign w26955 = w5308 & w21934;
assign w26956 = w5816 & ~w21973;
assign w26957 = ~w26954 & ~w26955;
assign w26958 = ~w26956 & w26957;
assign w26959 = a_20 & w26958;
assign w26960 = ~a_20 & ~w26958;
assign w26961 = ~w26959 & ~w26960;
assign w26962 = ~w26953 & w26961;
assign w26963 = ~w26952 & ~w26962;
assign w26964 = w26951 & ~w26963;
assign w26965 = ~w26951 & w26963;
assign w26966 = ~w26964 & ~w26965;
assign w26967 = w26941 & ~w26966;
assign w26968 = ~w26941 & w26966;
assign w26969 = ~w26967 & ~w26968;
assign w26970 = w26871 & w26969;
assign w26971 = ~w26871 & ~w26969;
assign w26972 = ~w26970 & ~w26971;
assign w26973 = w26868 & ~w26972;
assign w26974 = ~w26868 & w26972;
assign w26975 = ~w26973 & ~w26974;
assign w26976 = w26858 & w26975;
assign w26977 = ~w26858 & ~w26975;
assign w26978 = ~w26976 & ~w26977;
assign w26979 = ~w26856 & w26978;
assign w26980 = w26844 & w26979;
assign w26981 = ~w26856 & ~w26978;
assign w26982 = ~w26844 & w26981;
assign w26983 = ~w26980 & ~w26982;
assign w26984 = w26856 & ~w26978;
assign w26985 = w26844 & w26984;
assign w26986 = w26856 & w26978;
assign w26987 = ~w26844 & w26986;
assign w26988 = ~w26985 & ~w26987;
assign w26989 = w26983 & w26988;
assign w26990 = w9061 & w24756;
assign w26991 = w9089 & w24756;
assign w26992 = w7192 & w21762;
assign w26993 = w7489 & ~w22035;
assign w26994 = w7511 & w22032;
assign w26995 = ~w26992 & ~w26993;
assign w26996 = ~w26994 & w26995;
assign w26997 = a_11 & w26996;
assign w26998 = ~a_11 & ~w26996;
assign w26999 = ~w26997 & ~w26998;
assign w27000 = ~w26991 & w26999;
assign w27001 = ~w26990 & ~w27000;
assign w27002 = ~w26989 & w27001;
assign w27003 = w26989 & ~w27001;
assign w27004 = ~w27002 & ~w27003;
assign w27005 = w26841 & w27004;
assign w27006 = ~w26841 & ~w27004;
assign w27007 = ~w27005 & ~w27006;
assign w27008 = ~w26825 & ~w27007;
assign w27009 = w26825 & w27007;
assign w27010 = ~w27008 & ~w27009;
assign w27011 = w8295 & w21755;
assign w27012 = w8298 & ~w21757;
assign w27013 = w8277 & w22039;
assign w27014 = w8278 & ~w25675;
assign w27015 = ~w27012 & ~w27013;
assign w27016 = ~w27011 & w27015;
assign w27017 = ~w27014 & w27016;
assign w27018 = a_8 & w27017;
assign w27019 = ~a_8 & ~w27017;
assign w27020 = ~w27018 & ~w27019;
assign w27021 = w9788 & ~w21743;
assign w27022 = w9786 & w21752;
assign w27023 = w9780 & w21746;
assign w27024 = w9790 & w22065;
assign w27025 = ~w27022 & ~w27023;
assign w27026 = ~w27021 & w27025;
assign w27027 = ~w27024 & w27026;
assign w27028 = a_5 & w27027;
assign w27029 = ~a_5 & ~w27027;
assign w27030 = ~w27028 & ~w27029;
assign w27031 = w27020 & ~w27030;
assign w27032 = ~w27020 & w27030;
assign w27033 = ~w27031 & ~w27032;
assign w27034 = w27010 & ~w27033;
assign w27035 = ~w27010 & w27033;
assign w27036 = ~w27034 & ~w27035;
assign w27037 = w26813 & w27036;
assign w27038 = ~w26813 & ~w27036;
assign w27039 = ~w27037 & ~w27038;
assign w27040 = ~w26804 & w27039;
assign w27041 = w26804 & ~w27039;
assign w27042 = ~w27040 & ~w27041;
assign w27043 = ~w26761 & ~w26765;
assign w27044 = ~w26746 & ~w26748;
assign w27045 = ~a_31 & w35;
assign w27046 = w3887 & w3958;
assign w27047 = ~w27045 & ~w27046;
assign w27048 = w27044 & ~w27047;
assign w27049 = ~w27044 & w27047;
assign w27050 = ~w27048 & ~w27049;
assign w27051 = ~w26750 & w26755;
assign w27052 = w26750 & w26756;
assign w27053 = ~w27051 & ~w27052;
assign w27054 = w27050 & ~w27053;
assign w27055 = ~w27050 & w27053;
assign w27056 = ~w27054 & ~w27055;
assign w27057 = w27043 & w27056;
assign w27058 = ~w27043 & ~w27056;
assign w27059 = ~w27057 & ~w27058;
assign w27060 = w3 & w27059;
assign w27061 = w10835 & w26766;
assign w27062 = ~w26769 & ~w26773;
assign w27063 = ~w26766 & ~w27059;
assign w27064 = w26766 & w27059;
assign w27065 = ~w27063 & ~w27064;
assign w27066 = w27062 & w27065;
assign w27067 = ~w27062 & ~w27065;
assign w27068 = ~w27066 & ~w27067;
assign w27069 = w10837 & w27068;
assign w27070 = ~w27060 & ~w27061;
assign w27071 = ~w27069 & w27070;
assign w27072 = w10839 & w26476;
assign w27073 = a_2 & ~w27072;
assign w27074 = w27071 & ~w27073;
assign w27075 = a_2 & ~w27071;
assign w27076 = ~w27074 & ~w27075;
assign w27077 = w27042 & w27076;
assign w27078 = ~w27042 & ~w27076;
assign w27079 = ~w27077 & ~w27078;
assign w27080 = w26797 & ~w27079;
assign w27081 = ~w26797 & w27079;
assign w27082 = ~w27080 & ~w27081;
assign w27083 = w26793 & w27082;
assign w27084 = ~w26793 & ~w27082;
assign w27085 = ~w27083 & ~w27084;
assign w27086 = ~w26796 & ~w27077;
assign w27087 = ~w26790 & w27086;
assign w27088 = ~w27030 & w27039;
assign w27089 = ~w27041 & ~w27088;
assign w27090 = w3 & w27063;
assign w27091 = w10835 & w27059;
assign w27092 = w27059 & w27062;
assign w27093 = ~w26476 & w26773;
assign w27094 = ~w27092 & ~w27093;
assign w27095 = w10837 & w27094;
assign w27096 = ~w27090 & ~w27091;
assign w27097 = ~w27095 & w27096;
assign w27098 = w10839 & w26766;
assign w27099 = a_2 & ~w27098;
assign w27100 = w27097 & ~w27099;
assign w27101 = a_2 & ~w27097;
assign w27102 = ~w27100 & ~w27101;
assign w27103 = w27010 & ~w27020;
assign w27104 = ~w27010 & w27020;
assign w27105 = (~w27103 & w26813) | (~w27103 & w32244) | (w26813 & w32244);
assign w27106 = (w32244 & w37580) | (w32244 & w37581) | (w37580 & w37581);
assign w27107 = (~w32244 & w37582) | (~w32244 & w37583) | (w37582 & w37583);
assign w27108 = ~w27106 & ~w27107;
assign w27109 = w9788 & w26476;
assign w27110 = w9780 & ~w21743;
assign w27111 = w9786 & w21746;
assign w27112 = w9790 & w26489;
assign w27113 = ~w27110 & ~w27111;
assign w27114 = ~w27109 & w27113;
assign w27115 = ~w27112 & w27114;
assign w27116 = a_5 & ~w27115;
assign w27117 = ~a_5 & w27115;
assign w27118 = ~w27116 & ~w27117;
assign w27119 = ~w26841 & w27002;
assign w27120 = w26989 & w27001;
assign w27121 = w26841 & w27120;
assign w27122 = ~w27119 & ~w27121;
assign w27123 = (w27122 & ~w26825) | (w27122 & w32612) | (~w26825 & w32612);
assign w27124 = ~w26840 & w26988;
assign w27125 = w26983 & ~w27124;
assign w27126 = ~w26700 & w26983;
assign w27127 = w26549 & w27126;
assign w27128 = ~w27125 & ~w27127;
assign w27129 = w7511 & w22039;
assign w27130 = w7192 & ~w22035;
assign w27131 = w7489 & w22032;
assign w27132 = w7193 & w24962;
assign w27133 = ~w27130 & ~w27131;
assign w27134 = ~w27129 & w27133;
assign w27135 = ~w27132 & w27134;
assign w27136 = a_11 & ~w27135;
assign w27137 = ~a_11 & w27135;
assign w27138 = ~w27136 & ~w27137;
assign w27139 = (w32239 & w32613) | (w32239 & w32614) | (w32613 & w32614);
assign w27140 = ~w26858 & w26972;
assign w27141 = ~w27139 & ~w27140;
assign w27142 = w26868 & w27141;
assign w27143 = w26843 & ~w27142;
assign w27144 = ~w26829 & ~w26868;
assign w27145 = w26829 & w26868;
assign w27146 = ~w27141 & ~w27145;
assign w27147 = ~w27144 & ~w27146;
assign w27148 = ~w27143 & w27147;
assign w27149 = w6998 & w21771;
assign w27150 = w6996 & w21762;
assign w27151 = w6446 & ~w22020;
assign w27152 = w6447 & w24502;
assign w27153 = ~w27150 & ~w27151;
assign w27154 = ~w27149 & w27153;
assign w27155 = ~w27152 & w27154;
assign w27156 = ~a_14 & w27155;
assign w27157 = a_14 & ~w27155;
assign w27158 = ~w27156 & ~w27157;
assign w27159 = w26963 & w26972;
assign w27160 = ~w27139 & ~w27159;
assign w27161 = w26941 & w26951;
assign w27162 = ~w26869 & ~w27161;
assign w27163 = ~w26870 & w27162;
assign w27164 = ~w26941 & ~w26951;
assign w27165 = ~w26933 & ~w26939;
assign w27166 = ~w26888 & ~w26927;
assign w27167 = ~w26615 & w27166;
assign w27168 = (~w26928 & w26615) | (~w26928 & w32245) | (w26615 & w32245);
assign w27169 = w1102 & w1261;
assign w27170 = w1772 & w27169;
assign w27171 = w1454 & w4009;
assign w27172 = w4847 & w27171;
assign w27173 = w3372 & w3385;
assign w27174 = w3443 & w5173;
assign w27175 = w27173 & w27174;
assign w27176 = w15082 & w27172;
assign w27177 = w27170 & w27176;
assign w27178 = w27175 & w27177;
assign w27179 = w2950 & w27178;
assign w27180 = w4176 & w6656;
assign w27181 = w27179 & w27180;
assign w27182 = w1399 & ~w21839;
assign w27183 = w1327 & w21854;
assign w27184 = w668 & w21787;
assign w27185 = ~w27182 & ~w27183;
assign w27186 = ~w27184 & w27185;
assign w27187 = ~w27181 & ~w27186;
assign w27188 = w1478 & ~w27181;
assign w27189 = (~w27187 & w22726) | (~w27187 & w32615) | (w22726 & w32615);
assign w27190 = w1478 & ~w22726;
assign w27191 = w27181 & w27186;
assign w27192 = ~w27190 & w27191;
assign w27193 = w27189 & ~w27192;
assign w27194 = ~w26900 & ~w26922;
assign w27195 = (~w26921 & w26900) | (~w26921 & w32246) | (w26900 & w32246);
assign w27196 = ~w27193 & w27195;
assign w27197 = w27193 & ~w27195;
assign w27198 = ~w27196 & ~w27197;
assign w27199 = w7268 & w22096;
assign w27200 = w3957 & w21894;
assign w27201 = w4446 & w21892;
assign w27202 = w4068 & w21901;
assign w27203 = ~w27200 & ~w27201;
assign w27204 = ~w27202 & w27203;
assign w27205 = w7269 & w27204;
assign w27206 = a_29 & ~w27204;
assign w27207 = ~a_29 & w27204;
assign w27208 = ~w22096 & w27207;
assign w27209 = ~w27205 & ~w27206;
assign w27210 = ~w27199 & w27209;
assign w27211 = ~w27208 & w27210;
assign w27212 = w27210 & w32616;
assign w27213 = (~w27198 & ~w27210) | (~w27198 & w32617) | (~w27210 & w32617);
assign w27214 = ~w27212 & ~w27213;
assign w27215 = w27168 & w27214;
assign w27216 = ~w27168 & ~w27214;
assign w27217 = ~w27215 & ~w27216;
assign w27218 = ~w22901 & w32247;
assign w27219 = w4666 & w21951;
assign w27220 = w4638 & w21921;
assign w27221 = ~w518 & ~w21910;
assign w27222 = ~w27219 & ~w27220;
assign w27223 = ~w27221 & w27222;
assign w27224 = ~w27218 & w27223;
assign w27225 = ~a_26 & w27224;
assign w27226 = a_26 & ~w27224;
assign w27227 = ~w27225 & ~w27226;
assign w27228 = w5016 & ~w21945;
assign w27229 = w5080 & ~w21940;
assign w27230 = w5286 & w21934;
assign w27231 = ~w27228 & ~w27229;
assign w27232 = ~w27230 & w27231;
assign w27233 = ~a_23 & w27232;
assign w27234 = (w27233 & ~w22925) | (w27233 & w32248) | (~w22925 & w32248);
assign w27235 = w7961 & w23310;
assign w27236 = w7962 & w27232;
assign w27237 = a_23 & ~w27232;
assign w27238 = ~w27236 & ~w27237;
assign w27239 = ~w27234 & w27238;
assign w27240 = ~w27235 & w27239;
assign w27241 = w27227 & ~w27240;
assign w27242 = ~w27227 & w27240;
assign w27243 = ~w27241 & ~w27242;
assign w27244 = w27217 & ~w27243;
assign w27245 = ~w27217 & w27243;
assign w27246 = ~w27244 & ~w27245;
assign w27247 = w27165 & w27246;
assign w27248 = ~w27165 & ~w27246;
assign w27249 = ~w27247 & ~w27248;
assign w27250 = ~w27164 & ~w27249;
assign w27251 = ~w27163 & w27250;
assign w27252 = (~w27164 & ~w27162) | (~w27164 & w32249) | (~w27162 & w32249);
assign w27253 = w27249 & ~w27252;
assign w27254 = ~w27251 & ~w27253;
assign w27255 = w6304 & w22014;
assign w27256 = w6059 & ~w21992;
assign w27257 = w6061 & w22007;
assign w27258 = w6063 & w23398;
assign w27259 = ~w27256 & ~w27257;
assign w27260 = ~w27255 & w27259;
assign w27261 = ~w27258 & w27260;
assign w27262 = a_17 & w27261;
assign w27263 = ~a_17 & ~w27261;
assign w27264 = ~w27262 & ~w27263;
assign w27265 = w5816 & w21985;
assign w27266 = w5308 & ~w21968;
assign w27267 = w5818 & ~w21973;
assign w27268 = w5309 & w23553;
assign w27269 = ~w27265 & ~w27266;
assign w27270 = ~w27267 & w27269;
assign w27271 = ~w27268 & w27270;
assign w27272 = a_20 & ~w27271;
assign w27273 = ~a_20 & w27271;
assign w27274 = ~w27272 & ~w27273;
assign w27275 = w27264 & ~w27274;
assign w27276 = ~w27264 & w27274;
assign w27277 = ~w27275 & ~w27276;
assign w27278 = w27254 & ~w27277;
assign w27279 = ~w27254 & w27277;
assign w27280 = ~w27278 & ~w27279;
assign w27281 = w27160 & w27280;
assign w27282 = ~w27160 & ~w27280;
assign w27283 = ~w27281 & ~w27282;
assign w27284 = w27158 & ~w27283;
assign w27285 = ~w27158 & w27283;
assign w27286 = ~w27284 & ~w27285;
assign w27287 = w27148 & w27286;
assign w27288 = ~w27148 & ~w27286;
assign w27289 = ~w27287 & ~w27288;
assign w27290 = ~w27138 & w27289;
assign w27291 = w27128 & w27290;
assign w27292 = ~w27138 & ~w27289;
assign w27293 = ~w27128 & w27292;
assign w27294 = ~w27291 & ~w27293;
assign w27295 = w27138 & ~w27289;
assign w27296 = w27128 & w27295;
assign w27297 = w27138 & w27289;
assign w27298 = ~w27128 & w27297;
assign w27299 = ~w27296 & ~w27298;
assign w27300 = w27294 & w27299;
assign w27301 = w9456 & w26166;
assign w27302 = w8298 & w21755;
assign w27303 = w8277 & ~w21757;
assign w27304 = w8295 & w21752;
assign w27305 = ~w27302 & ~w27303;
assign w27306 = ~w27304 & w27305;
assign w27307 = a_8 & ~w27306;
assign w27308 = w8278 & w26166;
assign w27309 = ~a_8 & w27306;
assign w27310 = ~w27308 & w27309;
assign w27311 = ~w27301 & ~w27307;
assign w27312 = ~w27310 & w27311;
assign w27313 = ~w27300 & w27312;
assign w27314 = w27300 & ~w27312;
assign w27315 = ~w27313 & ~w27314;
assign w27316 = w27123 & w27315;
assign w27317 = ~w27123 & ~w27315;
assign w27318 = ~w27316 & ~w27317;
assign w27319 = w27118 & ~w27318;
assign w27320 = ~w27118 & w27318;
assign w27321 = ~w27319 & ~w27320;
assign w27322 = w27108 & ~w27321;
assign w27323 = ~w27108 & w27321;
assign w27324 = ~w27322 & ~w27323;
assign w27325 = w27089 & w27324;
assign w27326 = ~w27089 & ~w27324;
assign w27327 = ~w27325 & ~w27326;
assign w27328 = ~w27078 & ~w27327;
assign w27329 = ~w27087 & w27328;
assign w27330 = ~w27077 & w27327;
assign w27331 = ~w27081 & w27330;
assign w27332 = ~w27329 & ~w27331;
assign w27333 = w27083 & w27332;
assign w27334 = ~w27083 & ~w27332;
assign w27335 = ~w27333 & ~w27334;
assign w27336 = w27102 & w27327;
assign w27337 = ~w27329 & ~w27336;
assign w27338 = w27118 & w27318;
assign w27339 = w27105 & ~w27338;
assign w27340 = ~w27105 & ~w27319;
assign w27341 = ~w27339 & ~w27340;
assign w27342 = ~w27088 & ~w27341;
assign w27343 = ~w27041 & w27342;
assign w27344 = ~w27118 & ~w27318;
assign w27345 = w27105 & ~w27344;
assign w27346 = ~w27105 & ~w27320;
assign w27347 = ~w27345 & ~w27346;
assign w27348 = ~w27343 & ~w27347;
assign w27349 = w10835 & w27063;
assign w27350 = w27065 & ~w27092;
assign w27351 = w10837 & ~w27350;
assign w27352 = ~w27349 & ~w27351;
assign w27353 = w10839 & w27059;
assign w27354 = a_2 & ~w27353;
assign w27355 = w27352 & ~w27354;
assign w27356 = a_2 & ~w27352;
assign w27357 = ~w27355 & ~w27356;
assign w27358 = w27122 & w27299;
assign w27359 = w27294 & ~w27358;
assign w27360 = w27007 & w27294;
assign w27361 = w26825 & w27360;
assign w27362 = ~w27359 & ~w27361;
assign w27363 = w8295 & w21746;
assign w27364 = w8298 & w21752;
assign w27365 = w8277 & w21755;
assign w27366 = w8278 & ~w25700;
assign w27367 = ~w27364 & ~w27365;
assign w27368 = ~w27363 & w27367;
assign w27369 = ~w27366 & w27368;
assign w27370 = ~a_8 & w27369;
assign w27371 = a_8 & ~w27369;
assign w27372 = ~w27370 & ~w27371;
assign w27373 = ~w27128 & ~w27289;
assign w27374 = w27158 & w27289;
assign w27375 = (~w27374 & w27128) | (~w27374 & w32618) | (w27128 & w32618);
assign w27376 = w7511 & ~w21757;
assign w27377 = w7192 & w22032;
assign w27378 = w7489 & w22039;
assign w27379 = w7193 & ~w25205;
assign w27380 = ~w27377 & ~w27378;
assign w27381 = ~w27376 & w27380;
assign w27382 = ~w27379 & w27381;
assign w27383 = a_11 & w27382;
assign w27384 = ~a_11 & ~w27382;
assign w27385 = ~w27383 & ~w27384;
assign w27386 = w27148 & w27283;
assign w27387 = ~w27264 & ~w27283;
assign w27388 = (~w27387 & ~w27148) | (~w27387 & w32250) | (~w27148 & w32250);
assign w27389 = w6446 & w21771;
assign w27390 = w6998 & w21762;
assign w27391 = w6996 & ~w22035;
assign w27392 = w6447 & w24529;
assign w27393 = ~w27390 & ~w27391;
assign w27394 = ~w27389 & w27393;
assign w27395 = ~w27392 & w27394;
assign w27396 = a_14 & ~w27395;
assign w27397 = ~a_14 & w27395;
assign w27398 = ~w27396 & ~w27397;
assign w27399 = ~w27254 & ~w27274;
assign w27400 = (w27274 & w27163) | (w27274 & w32251) | (w27163 & w32251);
assign w27401 = ~w27253 & w27400;
assign w27402 = ~w27159 & ~w27401;
assign w27403 = ~w27139 & w27402;
assign w27404 = ~w27399 & ~w27403;
assign w27405 = w8391 & w24122;
assign w27406 = w8419 & w24122;
assign w27407 = w6061 & w22014;
assign w27408 = w6059 & w22007;
assign w27409 = w6304 & ~w22020;
assign w27410 = ~w27407 & ~w27408;
assign w27411 = ~w27409 & w27410;
assign w27412 = a_17 & w27411;
assign w27413 = ~a_17 & ~w27411;
assign w27414 = ~w27412 & ~w27413;
assign w27415 = ~w27406 & w27414;
assign w27416 = ~w27405 & ~w27415;
assign w27417 = w27240 & w27249;
assign w27418 = (~w27417 & w27163) | (~w27417 & w32252) | (w27163 & w32252);
assign w27419 = w27217 & w27227;
assign w27420 = ~w26933 & ~w27419;
assign w27421 = ~w26939 & w27420;
assign w27422 = ~w27217 & ~w27227;
assign w27423 = ~w27421 & ~w27422;
assign w27424 = ~w26921 & w27189;
assign w27425 = (~w27192 & w27194) | (~w27192 & w32253) | (w27194 & w32253);
assign w27426 = w1327 & w21787;
assign w27427 = w1399 & w21854;
assign w27428 = w668 & w21894;
assign w27429 = ~w27426 & ~w27427;
assign w27430 = ~w27428 & w27429;
assign w27431 = ~w83 & ~w237;
assign w27432 = w1362 & w27431;
assign w27433 = w1769 & w2942;
assign w27434 = w3631 & w13930;
assign w27435 = w27433 & w27434;
assign w27436 = w26582 & w27432;
assign w27437 = w27435 & w27436;
assign w27438 = w263 & w317;
assign w27439 = w808 & w1400;
assign w27440 = w1585 & w1605;
assign w27441 = w1689 & w2552;
assign w27442 = w3630 & w3678;
assign w27443 = w14598 & w27442;
assign w27444 = w27440 & w27441;
assign w27445 = w27438 & w27439;
assign w27446 = w2009 & w3563;
assign w27447 = w27445 & w27446;
assign w27448 = w27443 & w27444;
assign w27449 = w3153 & w27448;
assign w27450 = w27437 & w27447;
assign w27451 = w27449 & w27450;
assign w27452 = w4326 & w27451;
assign w27453 = w4923 & w27452;
assign w27454 = (~w23079 & w32619) | (~w23079 & w32620) | (w32619 & w32620);
assign w27455 = (w23079 & w32621) | (w23079 & w32622) | (w32621 & w32622);
assign w27456 = ~w27454 & ~w27455;
assign w27457 = w27425 & w27456;
assign w27458 = ~w27425 & ~w27456;
assign w27459 = ~w27457 & ~w27458;
assign w27460 = w4070 & ~w22580;
assign w27461 = w4068 & w21892;
assign w27462 = w3957 & w21901;
assign w27463 = w4446 & ~w21910;
assign w27464 = ~w27461 & ~w27462;
assign w27465 = ~w27463 & w27464;
assign w27466 = ~w27460 & w27465;
assign w27467 = ~a_29 & w27466;
assign w27468 = a_29 & ~w27466;
assign w27469 = ~w27467 & ~w27468;
assign w27470 = ~w27459 & ~w27469;
assign w27471 = w27459 & w27469;
assign w27472 = ~w27470 & ~w27471;
assign w27473 = (~w26928 & w27211) | (~w26928 & w32255) | (w27211 & w32255);
assign w27474 = (~w27212 & w27167) | (~w27212 & w32256) | (w27167 & w32256);
assign w27475 = ~w518 & w21921;
assign w27476 = w4638 & w21951;
assign w27477 = w4666 & ~w21945;
assign w27478 = ~w27475 & ~w27476;
assign w27479 = ~w27477 & w27478;
assign w27480 = (w27479 & ~w22083) | (w27479 & w32257) | (~w22083 & w32257);
assign w27481 = a_26 & ~w27480;
assign w27482 = ~a_26 & w27480;
assign w27483 = ~w27481 & ~w27482;
assign w27484 = w27474 & ~w27483;
assign w27485 = ~w27474 & w27483;
assign w27486 = ~w27484 & ~w27485;
assign w27487 = w27472 & w27486;
assign w27488 = ~w27472 & ~w27486;
assign w27489 = ~w27487 & ~w27488;
assign w27490 = w27423 & w27489;
assign w27491 = ~w27423 & ~w27489;
assign w27492 = ~w27490 & ~w27491;
assign w27493 = w5286 & ~w21968;
assign w27494 = w5016 & ~w21940;
assign w27495 = w5080 & w21934;
assign w27496 = w5017 & ~w23366;
assign w27497 = ~w27494 & ~w27495;
assign w27498 = ~w27493 & w27497;
assign w27499 = ~w27496 & w27498;
assign w27500 = a_23 & w27499;
assign w27501 = ~a_23 & ~w27499;
assign w27502 = ~w27500 & ~w27501;
assign w27503 = w5818 & w21985;
assign w27504 = w5308 & ~w21973;
assign w27505 = w5816 & ~w21992;
assign w27506 = ~w27503 & ~w27504;
assign w27507 = ~w27505 & w27506;
assign w27508 = a_20 & ~w27507;
assign w27509 = w8311 & ~w23930;
assign w27510 = w8339 & ~w23930;
assign w27511 = ~a_20 & w27507;
assign w27512 = ~w27510 & w27511;
assign w27513 = ~w27508 & ~w27509;
assign w27514 = ~w27512 & w27513;
assign w27515 = w27502 & ~w27514;
assign w27516 = ~w27502 & w27514;
assign w27517 = ~w27515 & ~w27516;
assign w27518 = w27492 & ~w27517;
assign w27519 = ~w27492 & w27517;
assign w27520 = ~w27518 & ~w27519;
assign w27521 = w27418 & w27520;
assign w27522 = ~w27418 & ~w27520;
assign w27523 = ~w27521 & ~w27522;
assign w27524 = w27416 & ~w27523;
assign w27525 = ~w27416 & w27523;
assign w27526 = ~w27524 & ~w27525;
assign w27527 = w27404 & w27526;
assign w27528 = ~w27404 & ~w27526;
assign w27529 = ~w27527 & ~w27528;
assign w27530 = w27398 & ~w27529;
assign w27531 = ~w27398 & w27529;
assign w27532 = ~w27530 & ~w27531;
assign w27533 = w27388 & w27532;
assign w27534 = ~w27388 & ~w27532;
assign w27535 = ~w27533 & ~w27534;
assign w27536 = w27385 & ~w27535;
assign w27537 = ~w27385 & w27535;
assign w27538 = ~w27536 & ~w27537;
assign w27539 = w27375 & w27538;
assign w27540 = ~w27375 & ~w27538;
assign w27541 = ~w27539 & ~w27540;
assign w27542 = w27372 & w27541;
assign w27543 = w27362 & w27542;
assign w27544 = w27372 & ~w27541;
assign w27545 = ~w27362 & w27544;
assign w27546 = ~w27543 & ~w27545;
assign w27547 = ~w27372 & ~w27541;
assign w27548 = w27362 & w27547;
assign w27549 = ~w27372 & w27541;
assign w27550 = ~w27362 & w27549;
assign w27551 = ~w27548 & ~w27550;
assign w27552 = w27546 & w27551;
assign w27553 = w10033 & ~w26774;
assign w27554 = w9780 & w26476;
assign w27555 = w9786 & ~w21743;
assign w27556 = w9788 & w26766;
assign w27557 = ~w27554 & ~w27555;
assign w27558 = ~w27556 & w27557;
assign w27559 = a_5 & ~w27558;
assign w27560 = w9790 & ~w26774;
assign w27561 = ~a_5 & w27558;
assign w27562 = ~w27560 & w27561;
assign w27563 = ~w27553 & ~w27559;
assign w27564 = ~w27562 & w27563;
assign w27565 = w27552 & ~w27564;
assign w27566 = ~w27552 & w27564;
assign w27567 = ~w27565 & ~w27566;
assign w27568 = ~w27105 & w27318;
assign w27569 = ~w27123 & w27313;
assign w27570 = w27300 & w27312;
assign w27571 = w27123 & w27570;
assign w27572 = ~w27569 & ~w27571;
assign w27573 = (w27572 & w27105) | (w27572 & w32623) | (w27105 & w32623);
assign w27574 = w27567 & ~w27573;
assign w27575 = ~w27567 & w27573;
assign w27576 = ~w27574 & ~w27575;
assign w27577 = w27357 & w27576;
assign w27578 = w27348 & w27577;
assign w27579 = w27357 & ~w27576;
assign w27580 = ~w27348 & w27579;
assign w27581 = ~w27578 & ~w27580;
assign w27582 = w27348 & ~w27576;
assign w27583 = ~w27348 & w27576;
assign w27584 = ~w27582 & ~w27583;
assign w27585 = ~w27357 & ~w27584;
assign w27586 = w27581 & ~w27585;
assign w27587 = w27337 & ~w27586;
assign w27588 = ~w27337 & w27586;
assign w27589 = ~w27587 & ~w27588;
assign w27590 = w27333 & w27589;
assign w27591 = ~w27333 & ~w27589;
assign w27592 = ~w27590 & ~w27591;
assign w27593 = ~w27336 & w27581;
assign w27594 = ~w27329 & w27593;
assign w27595 = ~w27585 & ~w27594;
assign w27596 = w27565 & ~w27573;
assign w27597 = ~w27564 & w27572;
assign w27598 = ~w27552 & w27597;
assign w27599 = ~w27568 & w27598;
assign w27600 = ~w27347 & ~w27599;
assign w27601 = ~w27596 & w27600;
assign w27602 = ~w27343 & w27601;
assign w27603 = w27566 & ~w27573;
assign w27604 = w27552 & w27564;
assign w27605 = w27573 & w27604;
assign w27606 = ~w27603 & ~w27605;
assign w27607 = ~w27602 & w27606;
assign w27608 = w27546 & w27572;
assign w27609 = w27551 & ~w27608;
assign w27610 = w27318 & w27551;
assign w27611 = ~w27105 & w27610;
assign w27612 = ~w27609 & ~w27611;
assign w27613 = w10839 & w27063;
assign w27614 = a_2 & ~w27613;
assign w27615 = w9788 & w27059;
assign w27616 = w9786 & w26476;
assign w27617 = w9780 & w26766;
assign w27618 = w9790 & w27068;
assign w27619 = ~w27616 & ~w27617;
assign w27620 = ~w27615 & w27619;
assign w27621 = ~w27618 & w27620;
assign w27622 = a_5 & w27621;
assign w27623 = ~a_5 & ~w27621;
assign w27624 = ~w27622 & ~w27623;
assign w27625 = w27614 & ~w27624;
assign w27626 = ~w27614 & w27624;
assign w27627 = ~w27625 & ~w27626;
assign w27628 = ~w27385 & ~w27541;
assign w27629 = w27385 & ~w27541;
assign w27630 = ~w27362 & ~w27629;
assign w27631 = ~w27628 & ~w27630;
assign w27632 = w8295 & ~w21743;
assign w27633 = w8298 & w21746;
assign w27634 = w8277 & w21752;
assign w27635 = w8278 & w22065;
assign w27636 = ~w27633 & ~w27634;
assign w27637 = ~w27632 & w27636;
assign w27638 = ~w27635 & w27637;
assign w27639 = ~a_8 & w27638;
assign w27640 = a_8 & ~w27638;
assign w27641 = ~w27639 & ~w27640;
assign w27642 = w27398 & w27529;
assign w27643 = ~w27388 & w27642;
assign w27644 = w27388 & w27530;
assign w27645 = ~w27643 & ~w27644;
assign w27646 = w27535 & w27645;
assign w27647 = ~w27374 & w27645;
assign w27648 = ~w27373 & w27647;
assign w27649 = ~w27646 & ~w27648;
assign w27650 = w27404 & ~w27524;
assign w27651 = w27416 & w27523;
assign w27652 = ~w27404 & ~w27651;
assign w27653 = ~w27650 & ~w27652;
assign w27654 = ~w27387 & ~w27653;
assign w27655 = ~w27386 & w27654;
assign w27656 = ~w27416 & w27529;
assign w27657 = (~w27656 & w27386) | (~w27656 & w32258) | (w27386 & w32258);
assign w27658 = w6996 & w22032;
assign w27659 = w6446 & w21762;
assign w27660 = w6998 & ~w22035;
assign w27661 = w6447 & w24756;
assign w27662 = ~w27658 & ~w27659;
assign w27663 = ~w27660 & w27662;
assign w27664 = ~w27661 & w27663;
assign w27665 = a_14 & ~w27664;
assign w27666 = ~a_14 & w27664;
assign w27667 = ~w27665 & ~w27666;
assign w27668 = ~w27399 & w27523;
assign w27669 = ~w27403 & w27668;
assign w27670 = w27514 & ~w27523;
assign w27671 = ~w27669 & ~w27670;
assign w27672 = ~w27492 & w27502;
assign w27673 = ~w27489 & ~w27502;
assign w27674 = w27423 & w27673;
assign w27675 = w27489 & ~w27502;
assign w27676 = ~w27423 & w27675;
assign w27677 = ~w27674 & ~w27676;
assign w27678 = ~w27417 & w27677;
assign w27679 = (~w27672 & w27251) | (~w27672 & w32259) | (w27251 & w32259);
assign w27680 = w27483 & ~w27489;
assign w27681 = ~w27490 & ~w27680;
assign w27682 = ~w27471 & w27474;
assign w27683 = (~w27470 & ~w27474) | (~w27470 & w32624) | (~w27474 & w32624);
assign w27684 = w4068 & ~w21910;
assign w27685 = w3957 & w21892;
assign w27686 = w4446 & w21921;
assign w27687 = ~w27684 & ~w27685;
assign w27688 = ~w27686 & w27687;
assign w27689 = (w27688 & ~w22664) | (w27688 & w32625) | (~w22664 & w32625);
assign w27690 = a_29 & ~w27689;
assign w27691 = ~a_29 & w27689;
assign w27692 = ~w27690 & ~w27691;
assign w27693 = ~w27454 & ~w27457;
assign w27694 = w668 & w21901;
assign w27695 = w1399 & w21787;
assign w27696 = w1327 & w21894;
assign w27697 = ~w27694 & ~w27695;
assign w27698 = ~w27696 & w27697;
assign w27699 = (w27698 & ~w22555) | (w27698 & w32260) | (~w22555 & w32260);
assign w27700 = w1534 & w2663;
assign w27701 = w3488 & w4159;
assign w27702 = w13348 & w27701;
assign w27703 = w1195 & w27700;
assign w27704 = w6138 & w27703;
assign w27705 = w1526 & w27702;
assign w27706 = w4155 & w27705;
assign w27707 = w4110 & w27704;
assign w27708 = w27706 & w27707;
assign w27709 = w5612 & w27708;
assign w27710 = w15258 & w27709;
assign w27711 = ~w27699 & ~w27710;
assign w27712 = w27699 & w27710;
assign w27713 = ~w27711 & ~w27712;
assign w27714 = w27693 & ~w27713;
assign w27715 = ~w27693 & w27713;
assign w27716 = ~w27714 & ~w27715;
assign w27717 = w27692 & w27716;
assign w27718 = ~w27692 & ~w27716;
assign w27719 = ~w27717 & ~w27718;
assign w27720 = w1226 & w23032;
assign w27721 = w4638 & ~w21945;
assign w27722 = ~w518 & w21951;
assign w27723 = w4666 & ~w21940;
assign w27724 = ~w27721 & ~w27722;
assign w27725 = ~w27723 & w27724;
assign w27726 = ~w27720 & w27725;
assign w27727 = ~a_26 & w27726;
assign w27728 = a_26 & ~w27726;
assign w27729 = ~w27727 & ~w27728;
assign w27730 = ~w27719 & w27729;
assign w27731 = w27683 & w27730;
assign w27732 = w27719 & w27729;
assign w27733 = ~w27683 & w27732;
assign w27734 = ~w27731 & ~w27733;
assign w27735 = w27719 & ~w27729;
assign w27736 = w27683 & w27735;
assign w27737 = ~w27719 & ~w27729;
assign w27738 = ~w27683 & w27737;
assign w27739 = ~w27736 & ~w27738;
assign w27740 = w27734 & w27739;
assign w27741 = w5286 & ~w21973;
assign w27742 = w5080 & ~w21968;
assign w27743 = w5016 & w21934;
assign w27744 = w5017 & ~w22930;
assign w27745 = ~w27742 & ~w27743;
assign w27746 = ~w27741 & w27745;
assign w27747 = ~w27744 & w27746;
assign w27748 = a_23 & ~w27747;
assign w27749 = ~a_23 & w27747;
assign w27750 = ~w27748 & ~w27749;
assign w27751 = w27740 & ~w27750;
assign w27752 = ~w27740 & w27750;
assign w27753 = ~w27751 & ~w27752;
assign w27754 = w27681 & w27753;
assign w27755 = ~w27681 & ~w27753;
assign w27756 = ~w27754 & ~w27755;
assign w27757 = w27679 & w27756;
assign w27758 = ~w27679 & ~w27756;
assign w27759 = ~w27757 & ~w27758;
assign w27760 = w6304 & w21771;
assign w27761 = w6059 & w22014;
assign w27762 = w6061 & ~w22020;
assign w27763 = w6063 & w24295;
assign w27764 = ~w27761 & ~w27762;
assign w27765 = ~w27760 & w27764;
assign w27766 = ~w27763 & w27765;
assign w27767 = a_17 & w27766;
assign w27768 = ~a_17 & ~w27766;
assign w27769 = ~w27767 & ~w27768;
assign w27770 = w5816 & w22007;
assign w27771 = w5818 & ~w21992;
assign w27772 = w5308 & w21985;
assign w27773 = w5309 & w23580;
assign w27774 = ~w27771 & ~w27772;
assign w27775 = ~w27770 & w27774;
assign w27776 = ~w27773 & w27775;
assign w27777 = ~a_20 & w27776;
assign w27778 = a_20 & ~w27776;
assign w27779 = ~w27777 & ~w27778;
assign w27780 = w27769 & ~w27779;
assign w27781 = ~w27769 & w27779;
assign w27782 = ~w27780 & ~w27781;
assign w27783 = w27759 & ~w27782;
assign w27784 = ~w27759 & w27782;
assign w27785 = ~w27783 & ~w27784;
assign w27786 = w27671 & w27785;
assign w27787 = ~w27671 & ~w27785;
assign w27788 = ~w27786 & ~w27787;
assign w27789 = ~w27667 & ~w27788;
assign w27790 = w27667 & w27788;
assign w27791 = ~w27789 & ~w27790;
assign w27792 = w27657 & ~w27791;
assign w27793 = ~w27657 & w27791;
assign w27794 = ~w27792 & ~w27793;
assign w27795 = w7511 & w21755;
assign w27796 = w7489 & ~w21757;
assign w27797 = w7192 & w22039;
assign w27798 = w7193 & ~w25675;
assign w27799 = ~w27796 & ~w27797;
assign w27800 = ~w27795 & w27799;
assign w27801 = ~w27798 & w27800;
assign w27802 = ~a_11 & w27801;
assign w27803 = a_11 & ~w27801;
assign w27804 = ~w27802 & ~w27803;
assign w27805 = w27794 & w27804;
assign w27806 = ~w27794 & ~w27804;
assign w27807 = ~w27805 & ~w27806;
assign w27808 = w27649 & w27807;
assign w27809 = ~w27649 & ~w27807;
assign w27810 = ~w27808 & ~w27809;
assign w27811 = w27641 & ~w27810;
assign w27812 = ~w27641 & w27810;
assign w27813 = ~w27811 & ~w27812;
assign w27814 = w27631 & w27813;
assign w27815 = ~w27631 & ~w27813;
assign w27816 = ~w27814 & ~w27815;
assign w27817 = w27627 & ~w27816;
assign w27818 = ~w27627 & w27816;
assign w27819 = ~w27817 & ~w27818;
assign w27820 = w27612 & w27819;
assign w27821 = ~w27612 & ~w27819;
assign w27822 = ~w27820 & ~w27821;
assign w27823 = ~w27607 & w27822;
assign w27824 = w27607 & ~w27822;
assign w27825 = ~w27823 & ~w27824;
assign w27826 = (w27825 & w27594) | (w27825 & w32626) | (w27594 & w32626);
assign w27827 = ~w27594 & w32627;
assign w27828 = ~w27826 & ~w27827;
assign w27829 = w27590 & w27828;
assign w27830 = ~w27590 & ~w27828;
assign w27831 = ~w27829 & ~w27830;
assign w27832 = ~w27612 & ~w27816;
assign w27833 = w27612 & w27816;
assign w27834 = ~w27832 & ~w27833;
assign w27835 = w27624 & ~w27834;
assign w27836 = w27602 & ~w27835;
assign w27837 = w27606 & w27624;
assign w27838 = w27564 & ~w27624;
assign w27839 = w27552 & w27838;
assign w27840 = w27573 & ~w27839;
assign w27841 = ~w27552 & w27838;
assign w27842 = ~w27573 & ~w27841;
assign w27843 = ~w27840 & ~w27842;
assign w27844 = ~w27834 & ~w27843;
assign w27845 = ~w27837 & ~w27844;
assign w27846 = ~w27836 & ~w27845;
assign w27847 = w27641 & w27816;
assign w27848 = ~w27832 & ~w27847;
assign w27849 = ~w27804 & w27810;
assign w27850 = ~w27628 & ~w27810;
assign w27851 = ~w27630 & w27850;
assign w27852 = ~w27849 & ~w27851;
assign w27853 = w9788 & w27063;
assign w27854 = w9780 & w27059;
assign w27855 = w9786 & w26766;
assign w27856 = w9790 & w27094;
assign w27857 = ~w27854 & ~w27855;
assign w27858 = ~w27853 & w27857;
assign w27859 = ~w27856 & w27858;
assign w27860 = ~a_5 & w27859;
assign w27861 = a_5 & ~w27859;
assign w27862 = ~w27860 & ~w27861;
assign w27863 = a_2 & w27862;
assign w27864 = ~a_2 & ~w27862;
assign w27865 = ~w27863 & ~w27864;
assign w27866 = ~w27656 & w27788;
assign w27867 = ~w27655 & w27866;
assign w27868 = (~w27789 & w27655) | (~w27789 & w32261) | (w27655 & w32261);
assign w27869 = ~w27792 & ~w27868;
assign w27870 = ~w27646 & ~w27869;
assign w27871 = ~w27648 & w27870;
assign w27872 = w27667 & w27794;
assign w27873 = ~w27871 & ~w27872;
assign w27874 = ~w27769 & ~w27788;
assign w27875 = (~w27874 & w27655) | (~w27874 & w32262) | (w27655 & w32262);
assign w27876 = w6996 & w22039;
assign w27877 = w6446 & ~w22035;
assign w27878 = w6998 & w22032;
assign w27879 = w6447 & w24962;
assign w27880 = ~w27877 & ~w27878;
assign w27881 = ~w27876 & w27880;
assign w27882 = ~w27879 & w27881;
assign w27883 = a_14 & ~w27882;
assign w27884 = ~a_14 & w27882;
assign w27885 = ~w27883 & ~w27884;
assign w27886 = ~w27759 & ~w27779;
assign w27887 = ~w27756 & w27779;
assign w27888 = w27679 & w27887;
assign w27889 = w27756 & w27779;
assign w27890 = ~w27679 & w27889;
assign w27891 = ~w27888 & ~w27890;
assign w27892 = ~w27670 & w27891;
assign w27893 = ~w27669 & w27892;
assign w27894 = ~w27886 & ~w27893;
assign w27895 = w27750 & ~w27756;
assign w27896 = ~w27757 & ~w27895;
assign w27897 = w5816 & w22014;
assign w27898 = w5308 & ~w21992;
assign w27899 = w5818 & w22007;
assign w27900 = w5309 & w23398;
assign w27901 = ~w27898 & ~w27899;
assign w27902 = ~w27897 & w27901;
assign w27903 = ~w27900 & w27902;
assign w27904 = a_20 & w27903;
assign w27905 = ~a_20 & ~w27903;
assign w27906 = ~w27904 & ~w27905;
assign w27907 = w6063 & w24502;
assign w27908 = w6059 & ~w22020;
assign w27909 = w6304 & w21762;
assign w27910 = w6061 & w21771;
assign w27911 = ~w27908 & ~w27909;
assign w27912 = ~w27910 & w27911;
assign w27913 = ~w27907 & w27912;
assign w27914 = a_17 & ~w27913;
assign w27915 = ~a_17 & w27913;
assign w27916 = ~w27914 & ~w27915;
assign w27917 = ~w27906 & ~w27916;
assign w27918 = w27906 & w27916;
assign w27919 = ~w27917 & ~w27918;
assign w27920 = ~w27680 & w27734;
assign w27921 = ~w27490 & w27920;
assign w27922 = w27739 & ~w27921;
assign w27923 = ~w27470 & ~w27718;
assign w27924 = ~w27682 & w27923;
assign w27925 = ~w27717 & ~w27924;
assign w27926 = ~w22901 & w32263;
assign w27927 = w4446 & w21951;
assign w27928 = w3957 & ~w21910;
assign w27929 = w4068 & w21921;
assign w27930 = ~w27927 & ~w27928;
assign w27931 = ~w27929 & w27930;
assign w27932 = ~w27926 & w27931;
assign w27933 = a_29 & ~w27932;
assign w27934 = ~a_29 & w27932;
assign w27935 = ~w27933 & ~w27934;
assign w27936 = ~w27454 & ~w27711;
assign w27937 = ~w27457 & w27936;
assign w27938 = ~w27712 & ~w27937;
assign w27939 = w1327 & w21901;
assign w27940 = w1399 & w21894;
assign w27941 = w668 & w21892;
assign w27942 = ~w27939 & ~w27940;
assign w27943 = ~w27941 & w27942;
assign w27944 = (w27943 & ~w22096) | (w27943 & w32264) | (~w22096 & w32264);
assign w27945 = ~w50 & ~w451;
assign w27946 = w735 & w27945;
assign w27947 = w3344 & w3518;
assign w27948 = w5373 & w27947;
assign w27949 = w27946 & w27948;
assign w27950 = ~w447 & w1111;
assign w27951 = w1206 & w1400;
assign w27952 = w1661 & w1821;
assign w27953 = w2362 & w3021;
assign w27954 = w27952 & w27953;
assign w27955 = w27950 & w27951;
assign w27956 = w1688 & w2163;
assign w27957 = w27955 & w27956;
assign w27958 = w14058 & w27954;
assign w27959 = w27170 & w27958;
assign w27960 = w27949 & w27957;
assign w27961 = w27959 & w27960;
assign w27962 = w2795 & w5398;
assign w27963 = w14349 & w27962;
assign w27964 = w27961 & w27963;
assign w27965 = ~w27944 & ~w27964;
assign w27966 = w27944 & w27964;
assign w27967 = ~w27965 & ~w27966;
assign w27968 = w27938 & ~w27967;
assign w27969 = ~w27938 & w27967;
assign w27970 = ~w27968 & ~w27969;
assign w27971 = w27935 & ~w27970;
assign w27972 = ~w27935 & w27970;
assign w27973 = ~w27971 & ~w27972;
assign w27974 = w4666 & w21934;
assign w27975 = ~w518 & ~w21945;
assign w27976 = w4638 & ~w21940;
assign w27977 = w1226 & w23310;
assign w27978 = ~w27974 & ~w27975;
assign w27979 = ~w27976 & w27978;
assign w27980 = ~w27977 & w27979;
assign w27981 = a_26 & ~w27980;
assign w27982 = ~a_26 & w27980;
assign w27983 = ~w27981 & ~w27982;
assign w27984 = w27973 & w27983;
assign w27985 = w27925 & w27984;
assign w27986 = ~w27973 & w27983;
assign w27987 = ~w27925 & w27986;
assign w27988 = ~w27985 & ~w27987;
assign w27989 = ~w27973 & ~w27983;
assign w27990 = w27925 & w27989;
assign w27991 = w27973 & ~w27983;
assign w27992 = ~w27925 & w27991;
assign w27993 = ~w27990 & ~w27992;
assign w27994 = w27988 & w27993;
assign w27995 = w5286 & w21985;
assign w27996 = w5016 & ~w21968;
assign w27997 = w5080 & ~w21973;
assign w27998 = w5017 & w23553;
assign w27999 = ~w27995 & ~w27996;
assign w28000 = ~w27997 & w27999;
assign w28001 = ~w27998 & w28000;
assign w28002 = a_23 & w28001;
assign w28003 = ~a_23 & ~w28001;
assign w28004 = ~w28002 & ~w28003;
assign w28005 = w27994 & ~w28004;
assign w28006 = ~w27994 & w28004;
assign w28007 = ~w28005 & ~w28006;
assign w28008 = w27922 & w28007;
assign w28009 = ~w27922 & ~w28007;
assign w28010 = ~w28008 & ~w28009;
assign w28011 = w27919 & ~w28010;
assign w28012 = ~w27919 & w28010;
assign w28013 = ~w28011 & ~w28012;
assign w28014 = w27896 & ~w28013;
assign w28015 = ~w27896 & w28013;
assign w28016 = ~w28014 & ~w28015;
assign w28017 = w27894 & w28016;
assign w28018 = ~w27894 & ~w28016;
assign w28019 = ~w28017 & ~w28018;
assign w28020 = w27885 & ~w28019;
assign w28021 = ~w27885 & w28019;
assign w28022 = ~w28020 & ~w28021;
assign w28023 = w27875 & w28022;
assign w28024 = ~w27875 & ~w28022;
assign w28025 = ~w28023 & ~w28024;
assign w28026 = w7511 & w21752;
assign w28027 = w7192 & ~w21757;
assign w28028 = w7489 & w21755;
assign w28029 = w7193 & w26166;
assign w28030 = ~w28027 & ~w28028;
assign w28031 = ~w28026 & w28030;
assign w28032 = ~w28029 & w28031;
assign w28033 = a_11 & w28032;
assign w28034 = ~a_11 & ~w28032;
assign w28035 = ~w28033 & ~w28034;
assign w28036 = w8295 & w26476;
assign w28037 = w8298 & ~w21743;
assign w28038 = w8277 & w21746;
assign w28039 = w8278 & w26489;
assign w28040 = ~w28037 & ~w28038;
assign w28041 = ~w28036 & w28040;
assign w28042 = ~w28039 & w28041;
assign w28043 = a_8 & ~w28042;
assign w28044 = ~a_8 & w28042;
assign w28045 = ~w28043 & ~w28044;
assign w28046 = w28035 & ~w28045;
assign w28047 = ~w28035 & w28045;
assign w28048 = ~w28046 & ~w28047;
assign w28049 = w28025 & ~w28048;
assign w28050 = ~w28025 & w28048;
assign w28051 = ~w28049 & ~w28050;
assign w28052 = w27873 & w28051;
assign w28053 = ~w27873 & ~w28051;
assign w28054 = ~w28052 & ~w28053;
assign w28055 = w27865 & ~w28054;
assign w28056 = ~w27865 & w28054;
assign w28057 = ~w28055 & ~w28056;
assign w28058 = w27852 & w28057;
assign w28059 = ~w27852 & ~w28057;
assign w28060 = ~w28058 & ~w28059;
assign w28061 = w27848 & ~w28060;
assign w28062 = (w28060 & w27832) | (w28060 & w32628) | (w27832 & w32628);
assign w28063 = ~w28061 & ~w28062;
assign w28064 = ~w27846 & ~w28063;
assign w28065 = w27846 & w28063;
assign w28066 = ~w28064 & ~w28065;
assign w28067 = w27614 & w27822;
assign w28068 = w27607 & w28067;
assign w28069 = w27614 & ~w27822;
assign w28070 = ~w27607 & w28069;
assign w28071 = ~w28068 & ~w28070;
assign w28072 = ~w28066 & ~w28071;
assign w28073 = w28066 & w28071;
assign w28074 = ~w28072 & ~w28073;
assign w28075 = ~w27827 & ~w28074;
assign w28076 = w27827 & ~w28066;
assign w28077 = ~w28075 & ~w28076;
assign w28078 = w27829 & ~w28077;
assign w28079 = ~w27829 & w28077;
assign w28080 = ~w28078 & ~w28079;
assign w28081 = ~w27863 & w28062;
assign w28082 = ~w27863 & ~w28060;
assign w28083 = (~w27864 & ~w27848) | (~w27864 & w32629) | (~w27848 & w32629);
assign w28084 = ~w28081 & w28083;
assign w28085 = w27804 & w27810;
assign w28086 = ~w27872 & w28025;
assign w28087 = ~w27871 & w28086;
assign w28088 = ~w28035 & w28087;
assign w28089 = ~w28025 & ~w28035;
assign w28090 = ~w27873 & w28089;
assign w28091 = ~w28088 & ~w28090;
assign w28092 = ~w28085 & w28091;
assign w28093 = ~w28025 & w28035;
assign w28094 = w27873 & w28093;
assign w28095 = w28025 & w28035;
assign w28096 = ~w27873 & w28095;
assign w28097 = ~w28094 & ~w28096;
assign w28098 = ~w28092 & w28097;
assign w28099 = ~w27810 & w28097;
assign w28100 = ~w27631 & w28099;
assign w28101 = ~w28098 & ~w28100;
assign w28102 = ~w27885 & ~w28025;
assign w28103 = ~w28087 & ~w28102;
assign w28104 = w8295 & w26766;
assign w28105 = w8277 & ~w21743;
assign w28106 = w8298 & w26476;
assign w28107 = w8278 & ~w26774;
assign w28108 = ~w28105 & ~w28106;
assign w28109 = ~w28104 & w28108;
assign w28110 = ~w28107 & w28109;
assign w28111 = a_8 & w28110;
assign w28112 = ~a_8 & ~w28110;
assign w28113 = ~w28111 & ~w28112;
assign w28114 = ~w27916 & ~w28019;
assign w28115 = ~w27874 & w28019;
assign w28116 = (~w28114 & w27867) | (~w28114 & w32265) | (w27867 & w32265);
assign w28117 = w7511 & w21746;
assign w28118 = w7489 & w21752;
assign w28119 = w7192 & w21755;
assign w28120 = w7193 & ~w25700;
assign w28121 = ~w28118 & ~w28119;
assign w28122 = ~w28117 & w28121;
assign w28123 = ~w28120 & w28122;
assign w28124 = a_11 & ~w28123;
assign w28125 = ~a_11 & w28123;
assign w28126 = ~w28124 & ~w28125;
assign w28127 = ~w27895 & w28010;
assign w28128 = ~w27757 & w28127;
assign w28129 = (~w28010 & w27757) | (~w28010 & w32266) | (w27757 & w32266);
assign w28130 = ~w28128 & ~w28129;
assign w28131 = ~w27906 & ~w28130;
assign w28132 = w27906 & w28130;
assign w28133 = (~w28131 & ~w27894) | (~w28131 & w32267) | (~w27894 & w32267);
assign w28134 = w28004 & ~w28010;
assign w28135 = ~w28128 & ~w28134;
assign w28136 = w5816 & ~w22020;
assign w28137 = w5818 & w22014;
assign w28138 = w5308 & w22007;
assign w28139 = w5309 & w24122;
assign w28140 = ~w28137 & ~w28138;
assign w28141 = ~w28136 & w28140;
assign w28142 = ~w28139 & w28141;
assign w28143 = a_20 & ~w28142;
assign w28144 = ~a_20 & w28142;
assign w28145 = ~w28143 & ~w28144;
assign w28146 = w6059 & w21771;
assign w28147 = w6061 & w21762;
assign w28148 = w6304 & ~w22035;
assign w28149 = w6063 & w24529;
assign w28150 = ~w28147 & ~w28148;
assign w28151 = ~w28146 & w28150;
assign w28152 = ~w28149 & w28151;
assign w28153 = a_17 & w28152;
assign w28154 = ~a_17 & ~w28152;
assign w28155 = ~w28153 & ~w28154;
assign w28156 = w28145 & ~w28155;
assign w28157 = ~w28145 & w28155;
assign w28158 = ~w28156 & ~w28157;
assign w28159 = ~w28128 & w32268;
assign w28160 = (~w28158 & w28128) | (~w28158 & w32269) | (w28128 & w32269);
assign w28161 = ~w28159 & ~w28160;
assign w28162 = w27739 & w27993;
assign w28163 = (w27988 & w27921) | (w27988 & w32270) | (w27921 & w32270);
assign w28164 = ~w27712 & ~w27966;
assign w28165 = ~w27937 & w28164;
assign w28166 = ~w27965 & ~w28165;
assign w28167 = ~w97 & w1266;
assign w28168 = w1562 & w2715;
assign w28169 = w2798 & w3444;
assign w28170 = w13564 & w13926;
assign w28171 = w28169 & w28170;
assign w28172 = w28167 & w28168;
assign w28173 = w1197 & w3091;
assign w28174 = w13470 & w28173;
assign w28175 = w28171 & w28172;
assign w28176 = w6631 & w13058;
assign w28177 = w28175 & w28176;
assign w28178 = w525 & w28174;
assign w28179 = w3312 & w28178;
assign w28180 = w2699 & w28177;
assign w28181 = w28179 & w28180;
assign w28182 = w1451 & w28181;
assign w28183 = a_2 & ~w28182;
assign w28184 = ~a_2 & w28182;
assign w28185 = ~w28183 & ~w28184;
assign w28186 = w1327 & w21892;
assign w28187 = w1399 & w21901;
assign w28188 = w668 & ~w21910;
assign w28189 = ~w28186 & ~w28187;
assign w28190 = ~w28188 & w28189;
assign w28191 = (w28190 & w22580) | (w28190 & w32271) | (w22580 & w32271);
assign w28192 = w28185 & ~w28191;
assign w28193 = ~w28185 & w28191;
assign w28194 = ~w28192 & ~w28193;
assign w28195 = w28166 & ~w28194;
assign w28196 = ~w28166 & w28194;
assign w28197 = ~w28195 & ~w28196;
assign w28198 = w4446 & ~w21945;
assign w28199 = w4068 & w21951;
assign w28200 = w3957 & w21921;
assign w28201 = ~w28199 & ~w28200;
assign w28202 = ~w28198 & w28201;
assign w28203 = (w28202 & ~w22083) | (w28202 & w32272) | (~w22083 & w32272);
assign w28204 = a_29 & ~w28203;
assign w28205 = ~a_29 & w28203;
assign w28206 = ~w28204 & ~w28205;
assign w28207 = ~w28197 & w28206;
assign w28208 = w28197 & ~w28206;
assign w28209 = ~w28207 & ~w28208;
assign w28210 = ~w518 & ~w21940;
assign w28211 = w4638 & w21934;
assign w28212 = w4666 & ~w21968;
assign w28213 = ~w28210 & ~w28211;
assign w28214 = ~w28212 & w28213;
assign w28215 = (w28214 & w23366) | (w28214 & w32273) | (w23366 & w32273);
assign w28216 = a_26 & ~w28215;
assign w28217 = ~a_26 & w28215;
assign w28218 = ~w28216 & ~w28217;
assign w28219 = w28209 & ~w28218;
assign w28220 = ~w28209 & w28218;
assign w28221 = ~w28219 & ~w28220;
assign w28222 = ~w27924 & w32274;
assign w28223 = ~w27972 & ~w28222;
assign w28224 = ~w28221 & w28223;
assign w28225 = w28221 & ~w28223;
assign w28226 = ~w28224 & ~w28225;
assign w28227 = w5286 & ~w21992;
assign w28228 = w5016 & ~w21973;
assign w28229 = w5080 & w21985;
assign w28230 = w5017 & ~w23930;
assign w28231 = ~w28228 & ~w28229;
assign w28232 = ~w28227 & w28231;
assign w28233 = ~w28230 & w28232;
assign w28234 = a_23 & w28233;
assign w28235 = ~a_23 & ~w28233;
assign w28236 = ~w28234 & ~w28235;
assign w28237 = w28226 & w28236;
assign w28238 = ~w28226 & ~w28236;
assign w28239 = ~w28237 & ~w28238;
assign w28240 = ~w28163 & ~w28239;
assign w28241 = w28163 & w28239;
assign w28242 = ~w28240 & ~w28241;
assign w28243 = w8564 & ~w25205;
assign w28244 = w8592 & ~w25205;
assign w28245 = w6998 & w22039;
assign w28246 = w6446 & w22032;
assign w28247 = w6996 & ~w21757;
assign w28248 = ~w28245 & ~w28246;
assign w28249 = ~w28247 & w28248;
assign w28250 = a_14 & w28249;
assign w28251 = ~a_14 & ~w28249;
assign w28252 = ~w28250 & ~w28251;
assign w28253 = ~w28244 & w28252;
assign w28254 = ~w28243 & ~w28253;
assign w28255 = w28242 & ~w28254;
assign w28256 = ~w28242 & w28254;
assign w28257 = ~w28255 & ~w28256;
assign w28258 = w28161 & ~w28257;
assign w28259 = ~w28161 & w28257;
assign w28260 = ~w28258 & ~w28259;
assign w28261 = w28133 & w28260;
assign w28262 = ~w28133 & ~w28260;
assign w28263 = ~w28261 & ~w28262;
assign w28264 = w28126 & ~w28263;
assign w28265 = ~w28126 & w28263;
assign w28266 = ~w28264 & ~w28265;
assign w28267 = w28116 & w28266;
assign w28268 = ~w28116 & ~w28266;
assign w28269 = ~w28267 & ~w28268;
assign w28270 = w28113 & w28269;
assign w28271 = ~w28113 & ~w28269;
assign w28272 = ~w28270 & ~w28271;
assign w28273 = ~w28103 & w28272;
assign w28274 = w28103 & ~w28272;
assign w28275 = ~w28273 & ~w28274;
assign w28276 = w9780 & w27063;
assign w28277 = w9786 & w27059;
assign w28278 = w9790 & ~w27350;
assign w28279 = ~w28276 & ~w28277;
assign w28280 = ~w28278 & w28279;
assign w28281 = ~a_5 & w28280;
assign w28282 = a_5 & ~w28280;
assign w28283 = ~w28281 & ~w28282;
assign w28284 = w28275 & ~w28283;
assign w28285 = w28101 & w28284;
assign w28286 = ~w28275 & ~w28283;
assign w28287 = ~w28101 & w28286;
assign w28288 = ~w28285 & ~w28287;
assign w28289 = ~w28101 & ~w28275;
assign w28290 = (w28283 & ~w28101) | (w28283 & w32275) | (~w28101 & w32275);
assign w28291 = ~w28289 & w28290;
assign w28292 = w28288 & ~w28291;
assign w28293 = ~w27851 & w32276;
assign w28294 = (~w28054 & w27851) | (~w28054 & w32277) | (w27851 & w32277);
assign w28295 = ~w28293 & ~w28294;
assign w28296 = ~w27847 & w28295;
assign w28297 = ~w27832 & w28296;
assign w28298 = ~w28045 & ~w28295;
assign w28299 = ~w28297 & ~w28298;
assign w28300 = ~w28292 & w28299;
assign w28301 = w28292 & ~w28299;
assign w28302 = ~w28300 & ~w28301;
assign w28303 = ~w28084 & w28302;
assign w28304 = w28084 & ~w28302;
assign w28305 = ~w28303 & ~w28304;
assign w28306 = ~w27825 & ~w28065;
assign w28307 = w27595 & w28306;
assign w28308 = ~w28065 & ~w28071;
assign w28309 = ~w28064 & ~w28308;
assign w28310 = ~w28307 & w28309;
assign w28311 = (w28305 & w28307) | (w28305 & w32278) | (w28307 & w32278);
assign w28312 = ~w28307 & w32279;
assign w28313 = ~w28311 & ~w28312;
assign w28314 = w28078 & w28313;
assign w28315 = ~w28078 & ~w28313;
assign w28316 = ~w28314 & ~w28315;
assign w28317 = ~w28307 & w32280;
assign w28318 = w28288 & ~w28298;
assign w28319 = ~w28297 & w28318;
assign w28320 = ~w28291 & ~w28319;
assign w28321 = w9785 & w27063;
assign w28322 = ~a_5 & ~w28321;
assign w28323 = w14378 & w27063;
assign w28324 = ~w28322 & ~w28323;
assign w28325 = ~w28087 & w32281;
assign w28326 = ~w28113 & ~w28325;
assign w28327 = ~w28273 & w28326;
assign w28328 = ~w28324 & w28327;
assign w28329 = w28324 & ~w28327;
assign w28330 = ~w28328 & ~w28329;
assign w28331 = ~w28289 & ~w28330;
assign w28332 = w28289 & w28330;
assign w28333 = ~w28331 & ~w28332;
assign w28334 = w28126 & w28269;
assign w28335 = ~w28325 & ~w28334;
assign w28336 = w9456 & w27068;
assign w28337 = w8298 & w26766;
assign w28338 = w8277 & w26476;
assign w28339 = w8295 & w27059;
assign w28340 = ~w28337 & ~w28338;
assign w28341 = ~w28339 & w28340;
assign w28342 = a_8 & ~w28341;
assign w28343 = w8278 & w27068;
assign w28344 = ~a_8 & w28341;
assign w28345 = ~w28343 & w28344;
assign w28346 = ~w28336 & ~w28342;
assign w28347 = ~w28345 & w28346;
assign w28348 = w28335 & ~w28347;
assign w28349 = ~w28335 & w28347;
assign w28350 = ~w28348 & ~w28349;
assign w28351 = w6996 & w21755;
assign w28352 = w6998 & ~w21757;
assign w28353 = w6446 & w22039;
assign w28354 = w6447 & ~w25675;
assign w28355 = ~w28352 & ~w28353;
assign w28356 = ~w28351 & w28355;
assign w28357 = ~w28354 & w28356;
assign w28358 = a_14 & ~w28357;
assign w28359 = ~a_14 & w28357;
assign w28360 = ~w28358 & ~w28359;
assign w28361 = w5816 & w21771;
assign w28362 = w5308 & w22014;
assign w28363 = w5818 & ~w22020;
assign w28364 = w5309 & w24295;
assign w28365 = ~w28362 & ~w28363;
assign w28366 = ~w28361 & w28365;
assign w28367 = ~w28364 & w28366;
assign w28368 = a_20 & w28367;
assign w28369 = ~a_20 & ~w28367;
assign w28370 = ~w28368 & ~w28369;
assign w28371 = w28239 & w32282;
assign w28372 = ~w28237 & ~w28370;
assign w28373 = w28237 & w28370;
assign w28374 = ~w28372 & ~w28373;
assign w28375 = ~w28241 & w28374;
assign w28376 = ~w28371 & ~w28375;
assign w28377 = ~w147 & w250;
assign w28378 = w560 & w28377;
assign w28379 = w472 & w28378;
assign w28380 = ~w191 & w1101;
assign w28381 = w1291 & w1454;
assign w28382 = w2017 & w2336;
assign w28383 = w3674 & w4152;
assign w28384 = w5365 & w28383;
assign w28385 = w28381 & w28382;
assign w28386 = w78 & w28380;
assign w28387 = w2455 & w25034;
assign w28388 = w28386 & w28387;
assign w28389 = w28384 & w28385;
assign w28390 = w28388 & w28389;
assign w28391 = w3281 & w28379;
assign w28392 = w28390 & w28391;
assign w28393 = w3078 & w28392;
assign w28394 = w15364 & w28393;
assign w28395 = ~a_2 & w28394;
assign w28396 = a_2 & ~w28394;
assign w28397 = ~w28395 & ~w28396;
assign w28398 = ~w28183 & ~w28192;
assign w28399 = w28397 & w28398;
assign w28400 = ~w28397 & ~w28398;
assign w28401 = ~w28399 & ~w28400;
assign w28402 = w1327 & ~w21910;
assign w28403 = w1399 & w21892;
assign w28404 = w668 & w21921;
assign w28405 = w1478 & w22664;
assign w28406 = ~w28402 & ~w28403;
assign w28407 = ~w28404 & w28406;
assign w28408 = ~w28405 & w28407;
assign w28409 = ~w28401 & ~w28408;
assign w28410 = w28401 & w28408;
assign w28411 = ~w28409 & ~w28410;
assign w28412 = (~w28195 & ~w28197) | (~w28195 & w32283) | (~w28197 & w32283);
assign w28413 = w28411 & ~w28412;
assign w28414 = ~w28411 & w28412;
assign w28415 = ~w28413 & ~w28414;
assign w28416 = w4666 & ~w21973;
assign w28417 = w4638 & ~w21968;
assign w28418 = ~w518 & w21934;
assign w28419 = w1226 & ~w22930;
assign w28420 = ~w28417 & ~w28418;
assign w28421 = ~w28416 & w28420;
assign w28422 = ~w28419 & w28421;
assign w28423 = a_26 & ~w28422;
assign w28424 = ~a_26 & w28422;
assign w28425 = ~w28423 & ~w28424;
assign w28426 = w4068 & ~w21945;
assign w28427 = w3957 & w21951;
assign w28428 = w4446 & ~w21940;
assign w28429 = w4070 & w23032;
assign w28430 = ~w28426 & ~w28427;
assign w28431 = ~w28428 & w28430;
assign w28432 = ~w28429 & w28431;
assign w28433 = a_29 & ~w28432;
assign w28434 = ~a_29 & w28432;
assign w28435 = ~w28433 & ~w28434;
assign w28436 = w28425 & w28435;
assign w28437 = ~w28425 & ~w28435;
assign w28438 = ~w28436 & ~w28437;
assign w28439 = ~w28415 & w28438;
assign w28440 = w28415 & ~w28438;
assign w28441 = ~w28439 & ~w28440;
assign w28442 = (~w28219 & ~w28221) | (~w28219 & w32284) | (~w28221 & w32284);
assign w28443 = w5286 & w22007;
assign w28444 = w5080 & ~w21992;
assign w28445 = w5016 & w21985;
assign w28446 = w5017 & w23580;
assign w28447 = ~w28444 & ~w28445;
assign w28448 = ~w28443 & w28447;
assign w28449 = ~w28446 & w28448;
assign w28450 = a_23 & ~w28449;
assign w28451 = ~a_23 & w28449;
assign w28452 = ~w28450 & ~w28451;
assign w28453 = ~w28442 & ~w28452;
assign w28454 = w28442 & w28452;
assign w28455 = ~w28453 & ~w28454;
assign w28456 = w28441 & ~w28455;
assign w28457 = ~w28441 & w28455;
assign w28458 = ~w28456 & ~w28457;
assign w28459 = ~w28375 & w32285;
assign w28460 = (w28458 & w28375) | (w28458 & w32286) | (w28375 & w32286);
assign w28461 = ~w28459 & ~w28460;
assign w28462 = w6304 & w22032;
assign w28463 = w6059 & w21762;
assign w28464 = w6061 & ~w22035;
assign w28465 = w6063 & w24756;
assign w28466 = ~w28462 & ~w28463;
assign w28467 = ~w28464 & w28466;
assign w28468 = ~w28465 & w28467;
assign w28469 = a_17 & ~w28468;
assign w28470 = ~a_17 & w28468;
assign w28471 = ~w28469 & ~w28470;
assign w28472 = ~w28461 & w28471;
assign w28473 = w28458 & ~w28471;
assign w28474 = w28376 & w28473;
assign w28475 = ~w28458 & ~w28471;
assign w28476 = ~w28376 & w28475;
assign w28477 = ~w28474 & ~w28476;
assign w28478 = ~w28472 & w28477;
assign w28479 = w28145 & ~w28242;
assign w28480 = ~w28145 & w28242;
assign w28481 = (~w28479 & ~w28135) | (~w28479 & w32287) | (~w28135 & w32287);
assign w28482 = ~w28478 & w28481;
assign w28483 = w28478 & ~w28481;
assign w28484 = ~w28482 & ~w28483;
assign w28485 = w28360 & w28484;
assign w28486 = ~w28360 & ~w28484;
assign w28487 = ~w28485 & ~w28486;
assign w28488 = w28161 & w28242;
assign w28489 = ~w28161 & ~w28242;
assign w28490 = ~w28488 & ~w28489;
assign w28491 = w28133 & ~w28490;
assign w28492 = w28155 & w28490;
assign w28493 = ~w28491 & ~w28492;
assign w28494 = w28487 & w28493;
assign w28495 = ~w28487 & ~w28493;
assign w28496 = ~w28494 & ~w28495;
assign w28497 = ~w28254 & ~w28263;
assign w28498 = (~w28497 & w28116) | (~w28497 & w32288) | (w28116 & w32288);
assign w28499 = ~w28496 & ~w28498;
assign w28500 = w28496 & w28498;
assign w28501 = ~w28499 & ~w28500;
assign w28502 = w7511 & ~w21743;
assign w28503 = w7489 & w21746;
assign w28504 = w7192 & w21752;
assign w28505 = w7193 & w22065;
assign w28506 = ~w28503 & ~w28504;
assign w28507 = ~w28502 & w28506;
assign w28508 = ~w28505 & w28507;
assign w28509 = ~a_11 & w28508;
assign w28510 = a_11 & ~w28508;
assign w28511 = ~w28509 & ~w28510;
assign w28512 = w28501 & ~w28511;
assign w28513 = ~w28501 & w28511;
assign w28514 = ~w28512 & ~w28513;
assign w28515 = w28350 & w28514;
assign w28516 = ~w28350 & ~w28514;
assign w28517 = ~w28515 & ~w28516;
assign w28518 = ~w28333 & ~w28517;
assign w28519 = w28333 & w28517;
assign w28520 = ~w28518 & ~w28519;
assign w28521 = w28320 & ~w28520;
assign w28522 = ~w28320 & w28520;
assign w28523 = ~w28521 & ~w28522;
assign w28524 = w28303 & ~w28523;
assign w28525 = ~w28303 & w28523;
assign w28526 = ~w28524 & ~w28525;
assign w28527 = ~w28317 & w28526;
assign w28528 = ~w28304 & w28523;
assign w28529 = w28310 & w28528;
assign w28530 = ~w28527 & ~w28529;
assign w28531 = w28314 & ~w28530;
assign w28532 = ~w28314 & w28530;
assign w28533 = ~w28531 & ~w28532;
assign w28534 = ~w28311 & w28528;
assign w28535 = w28324 & ~w28331;
assign w28536 = ~w28518 & ~w28535;
assign w28537 = ~w28485 & ~w28494;
assign w28538 = w6998 & w21755;
assign w28539 = w6446 & ~w21757;
assign w28540 = w6996 & w21752;
assign w28541 = ~w28538 & ~w28539;
assign w28542 = ~w28540 & w28541;
assign w28543 = (w28542 & ~w26166) | (w28542 & w32289) | (~w26166 & w32289);
assign w28544 = a_14 & ~w28543;
assign w28545 = ~a_14 & w28543;
assign w28546 = ~w28544 & ~w28545;
assign w28547 = w28472 & w28546;
assign w28548 = w28477 & w28546;
assign w28549 = ~w28481 & w28548;
assign w28550 = ~w28547 & ~w28549;
assign w28551 = w28477 & ~w28481;
assign w28552 = ~w28472 & ~w28546;
assign w28553 = ~w28551 & w28552;
assign w28554 = w28550 & ~w28553;
assign w28555 = ~w169 & ~w265;
assign w28556 = ~w2716 & w28555;
assign w28557 = w584 & w624;
assign w28558 = w757 & w13094;
assign w28559 = w28557 & w28558;
assign w28560 = w1114 & w28556;
assign w28561 = w5579 & w28560;
assign w28562 = w4087 & w28559;
assign w28563 = w14561 & w28562;
assign w28564 = w1902 & w28561;
assign w28565 = w5525 & w28564;
assign w28566 = w28563 & w28565;
assign w28567 = w3037 & w28566;
assign w28568 = w3646 & w28567;
assign w28569 = a_2 & ~w28568;
assign w28570 = ~a_2 & w28568;
assign w28571 = ~w28569 & ~w28570;
assign w28572 = ~w28395 & ~w28398;
assign w28573 = ~w28396 & ~w28572;
assign w28574 = w28571 & ~w28573;
assign w28575 = ~w28571 & w28573;
assign w28576 = ~w28574 & ~w28575;
assign w28577 = w1327 & w21921;
assign w28578 = w1399 & ~w21910;
assign w28579 = w668 & w21951;
assign w28580 = w1478 & w22905;
assign w28581 = ~w28577 & ~w28578;
assign w28582 = ~w28579 & w28581;
assign w28583 = ~w28580 & w28582;
assign w28584 = w28576 & ~w28583;
assign w28585 = ~w28576 & w28583;
assign w28586 = ~w28584 & ~w28585;
assign w28587 = ~w28410 & ~w28413;
assign w28588 = w28586 & ~w28587;
assign w28589 = ~w28586 & w28587;
assign w28590 = ~w28588 & ~w28589;
assign w28591 = w3957 & ~w21945;
assign w28592 = w4446 & w21934;
assign w28593 = w4068 & ~w21940;
assign w28594 = w4070 & w23310;
assign w28595 = ~w28591 & ~w28592;
assign w28596 = ~w28593 & w28595;
assign w28597 = ~w28594 & w28596;
assign w28598 = a_29 & ~w28597;
assign w28599 = ~a_29 & w28597;
assign w28600 = ~w28598 & ~w28599;
assign w28601 = w4666 & w21985;
assign w28602 = ~w518 & ~w21968;
assign w28603 = w4638 & ~w21973;
assign w28604 = w1226 & w23553;
assign w28605 = ~w28601 & ~w28602;
assign w28606 = ~w28603 & w28605;
assign w28607 = ~w28604 & w28606;
assign w28608 = a_26 & ~w28607;
assign w28609 = ~a_26 & w28607;
assign w28610 = ~w28608 & ~w28609;
assign w28611 = ~w28600 & ~w28610;
assign w28612 = w28600 & w28610;
assign w28613 = ~w28611 & ~w28612;
assign w28614 = ~w28590 & ~w28613;
assign w28615 = w28590 & w28613;
assign w28616 = ~w28614 & ~w28615;
assign w28617 = ~w28436 & ~w28439;
assign w28618 = w5286 & w22014;
assign w28619 = w5016 & ~w21992;
assign w28620 = w5080 & w22007;
assign w28621 = w5017 & w23398;
assign w28622 = ~w28619 & ~w28620;
assign w28623 = ~w28618 & w28622;
assign w28624 = ~w28621 & w28623;
assign w28625 = a_23 & w28624;
assign w28626 = ~a_23 & ~w28624;
assign w28627 = ~w28625 & ~w28626;
assign w28628 = w28617 & w28627;
assign w28629 = ~w28617 & ~w28627;
assign w28630 = ~w28628 & ~w28629;
assign w28631 = ~w28616 & w28630;
assign w28632 = w28616 & ~w28630;
assign w28633 = ~w28631 & ~w28632;
assign w28634 = ~w28453 & ~w28457;
assign w28635 = w5818 & w21771;
assign w28636 = w5816 & w21762;
assign w28637 = w5308 & ~w22020;
assign w28638 = w5309 & w24502;
assign w28639 = ~w28636 & ~w28637;
assign w28640 = ~w28635 & w28639;
assign w28641 = ~w28638 & w28640;
assign w28642 = ~a_20 & w28641;
assign w28643 = a_20 & ~w28641;
assign w28644 = ~w28642 & ~w28643;
assign w28645 = w28634 & w28644;
assign w28646 = ~w28634 & ~w28644;
assign w28647 = ~w28645 & ~w28646;
assign w28648 = w28633 & w28647;
assign w28649 = ~w28633 & ~w28647;
assign w28650 = ~w28648 & ~w28649;
assign w28651 = w28370 & ~w28375;
assign w28652 = ~w28460 & ~w28651;
assign w28653 = w6304 & w22039;
assign w28654 = w6059 & ~w22035;
assign w28655 = w6061 & w22032;
assign w28656 = w6063 & w24962;
assign w28657 = ~w28654 & ~w28655;
assign w28658 = ~w28653 & w28657;
assign w28659 = ~w28656 & w28658;
assign w28660 = ~a_17 & w28659;
assign w28661 = a_17 & ~w28659;
assign w28662 = ~w28660 & ~w28661;
assign w28663 = ~w28652 & ~w28662;
assign w28664 = w28652 & w28662;
assign w28665 = ~w28663 & ~w28664;
assign w28666 = w28650 & ~w28665;
assign w28667 = ~w28650 & w28665;
assign w28668 = ~w28666 & ~w28667;
assign w28669 = ~w28554 & w28668;
assign w28670 = w28554 & ~w28668;
assign w28671 = ~w28669 & ~w28670;
assign w28672 = w7511 & w26476;
assign w28673 = w7489 & ~w21743;
assign w28674 = w7192 & w21746;
assign w28675 = w7193 & w26489;
assign w28676 = ~w28673 & ~w28674;
assign w28677 = ~w28672 & w28676;
assign w28678 = ~w28675 & w28677;
assign w28679 = a_11 & ~w28678;
assign w28680 = ~a_11 & w28678;
assign w28681 = ~w28679 & ~w28680;
assign w28682 = w28671 & w28681;
assign w28683 = ~w28671 & ~w28681;
assign w28684 = ~w28682 & ~w28683;
assign w28685 = w28537 & ~w28684;
assign w28686 = ~w28537 & w28684;
assign w28687 = ~w28685 & ~w28686;
assign w28688 = w8295 & w27063;
assign w28689 = w8298 & w27059;
assign w28690 = w8277 & w26766;
assign w28691 = w8278 & w27094;
assign w28692 = ~w28689 & ~w28690;
assign w28693 = ~w28688 & w28692;
assign w28694 = ~w28691 & w28693;
assign w28695 = a_8 & ~w28694;
assign w28696 = ~a_8 & w28694;
assign w28697 = ~w28695 & ~w28696;
assign w28698 = w28687 & w28697;
assign w28699 = ~w28687 & ~w28697;
assign w28700 = ~w28698 & ~w28699;
assign w28701 = ~w28499 & w28511;
assign w28702 = ~w28500 & ~w28701;
assign w28703 = w28700 & ~w28702;
assign w28704 = ~w28700 & w28702;
assign w28705 = ~w28703 & ~w28704;
assign w28706 = a_5 & w28705;
assign w28707 = ~a_5 & ~w28705;
assign w28708 = ~w28706 & ~w28707;
assign w28709 = ~w28348 & ~w28514;
assign w28710 = ~w28349 & ~w28709;
assign w28711 = w28708 & ~w28710;
assign w28712 = ~w28708 & w28710;
assign w28713 = ~w28711 & ~w28712;
assign w28714 = w28536 & ~w28713;
assign w28715 = ~w28536 & w28713;
assign w28716 = ~w28714 & ~w28715;
assign w28717 = w28521 & ~w28716;
assign w28718 = ~w28521 & w28716;
assign w28719 = ~w28717 & ~w28718;
assign w28720 = w28534 & w28719;
assign w28721 = ~w28534 & ~w28719;
assign w28722 = ~w28720 & ~w28721;
assign w28723 = w28531 & w28722;
assign w28724 = ~w28531 & ~w28722;
assign w28725 = ~w28723 & ~w28724;
assign w28726 = ~w28707 & ~w28710;
assign w28727 = ~w28706 & ~w28726;
assign w28728 = w8298 & w27063;
assign w28729 = w8277 & w27059;
assign w28730 = w8278 & ~w27350;
assign w28731 = ~w28728 & ~w28729;
assign w28732 = ~w28730 & w28731;
assign w28733 = ~a_8 & w28732;
assign w28734 = a_8 & ~w28732;
assign w28735 = ~w28733 & ~w28734;
assign w28736 = ~w28699 & ~w28702;
assign w28737 = ~w28736 & w32290;
assign w28738 = (w28735 & w28736) | (w28735 & w32291) | (w28736 & w32291);
assign w28739 = ~w28737 & ~w28738;
assign w28740 = (w28550 & ~w28554) | (w28550 & w32292) | (~w28554 & w32292);
assign w28741 = w6996 & w21746;
assign w28742 = w6998 & w21752;
assign w28743 = w6446 & w21755;
assign w28744 = w6447 & ~w25700;
assign w28745 = ~w28742 & ~w28743;
assign w28746 = ~w28741 & w28745;
assign w28747 = ~w28744 & w28746;
assign w28748 = a_14 & ~w28747;
assign w28749 = ~a_14 & w28747;
assign w28750 = ~w28748 & ~w28749;
assign w28751 = ~w28740 & w28750;
assign w28752 = w28740 & ~w28750;
assign w28753 = ~w28751 & ~w28752;
assign w28754 = ~w28663 & ~w28667;
assign w28755 = w6304 & ~w21757;
assign w28756 = w6061 & w22039;
assign w28757 = w6059 & w22032;
assign w28758 = w6063 & ~w25205;
assign w28759 = ~w28756 & ~w28757;
assign w28760 = ~w28755 & w28759;
assign w28761 = ~w28758 & w28760;
assign w28762 = a_17 & ~w28761;
assign w28763 = ~a_17 & w28761;
assign w28764 = ~w28762 & ~w28763;
assign w28765 = w28754 & w28764;
assign w28766 = ~w28754 & ~w28764;
assign w28767 = ~w28765 & ~w28766;
assign w28768 = ~w28645 & ~w28648;
assign w28769 = ~w28585 & ~w28588;
assign w28770 = ~w195 & ~w878;
assign w28771 = w1585 & w28770;
assign w28772 = w2102 & w2185;
assign w28773 = w3237 & w4850;
assign w28774 = w28772 & w28773;
assign w28775 = w5389 & w28771;
assign w28776 = w15208 & w28775;
assign w28777 = w13569 & w28774;
assign w28778 = w28776 & w28777;
assign w28779 = w24825 & w28778;
assign w28780 = w4270 & w28779;
assign w28781 = w3455 & w28780;
assign w28782 = ~a_2 & ~w28781;
assign w28783 = a_2 & w28781;
assign w28784 = ~w28782 & ~w28783;
assign w28785 = ~a_5 & w28784;
assign w28786 = a_5 & ~w28784;
assign w28787 = ~w28785 & ~w28786;
assign w28788 = w668 & ~w21945;
assign w28789 = w1327 & w21951;
assign w28790 = w1399 & w21921;
assign w28791 = w1478 & w22083;
assign w28792 = ~w28789 & ~w28790;
assign w28793 = ~w28788 & w28792;
assign w28794 = ~w28791 & w28793;
assign w28795 = w28787 & ~w28794;
assign w28796 = ~w28787 & w28794;
assign w28797 = ~w28795 & ~w28796;
assign w28798 = ~w28569 & ~w28574;
assign w28799 = w28797 & w28798;
assign w28800 = ~w28797 & ~w28798;
assign w28801 = ~w28799 & ~w28800;
assign w28802 = w4446 & ~w21968;
assign w28803 = w4068 & w21934;
assign w28804 = w3957 & ~w21940;
assign w28805 = w4070 & ~w23366;
assign w28806 = ~w28803 & ~w28804;
assign w28807 = ~w28802 & w28806;
assign w28808 = ~w28805 & w28807;
assign w28809 = a_29 & ~w28808;
assign w28810 = ~a_29 & w28808;
assign w28811 = ~w28809 & ~w28810;
assign w28812 = ~w28801 & w28811;
assign w28813 = w28801 & ~w28811;
assign w28814 = ~w28812 & ~w28813;
assign w28815 = w28769 & w28814;
assign w28816 = ~w28769 & ~w28814;
assign w28817 = ~w28815 & ~w28816;
assign w28818 = w4666 & ~w21992;
assign w28819 = ~w518 & ~w21973;
assign w28820 = w4638 & w21985;
assign w28821 = w1226 & ~w23930;
assign w28822 = ~w28819 & ~w28820;
assign w28823 = ~w28818 & w28822;
assign w28824 = ~w28821 & w28823;
assign w28825 = a_26 & w28824;
assign w28826 = ~a_26 & ~w28824;
assign w28827 = ~w28825 & ~w28826;
assign w28828 = w28817 & ~w28827;
assign w28829 = ~w28817 & w28827;
assign w28830 = ~w28828 & ~w28829;
assign w28831 = ~w28611 & ~w28615;
assign w28832 = w5286 & ~w22020;
assign w28833 = w5016 & w22007;
assign w28834 = w5080 & w22014;
assign w28835 = w5017 & w24122;
assign w28836 = ~w28833 & ~w28834;
assign w28837 = ~w28832 & w28836;
assign w28838 = ~w28835 & w28837;
assign w28839 = a_23 & w28838;
assign w28840 = ~a_23 & ~w28838;
assign w28841 = ~w28839 & ~w28840;
assign w28842 = ~w28831 & w28841;
assign w28843 = ~w28830 & w28842;
assign w28844 = w28831 & w28841;
assign w28845 = w28830 & w28844;
assign w28846 = ~w28843 & ~w28845;
assign w28847 = w28831 & ~w28841;
assign w28848 = ~w28830 & w28847;
assign w28849 = ~w28831 & ~w28841;
assign w28850 = w28830 & w28849;
assign w28851 = ~w28848 & ~w28850;
assign w28852 = w28846 & w28851;
assign w28853 = ~w28629 & ~w28631;
assign w28854 = w5308 & w21771;
assign w28855 = w5818 & w21762;
assign w28856 = w5816 & ~w22035;
assign w28857 = w5309 & w24529;
assign w28858 = ~w28855 & ~w28856;
assign w28859 = ~w28854 & w28858;
assign w28860 = ~w28857 & w28859;
assign w28861 = a_20 & ~w28860;
assign w28862 = ~a_20 & w28860;
assign w28863 = ~w28861 & ~w28862;
assign w28864 = ~w28853 & ~w28863;
assign w28865 = w28852 & w28864;
assign w28866 = w28853 & ~w28863;
assign w28867 = ~w28852 & w28866;
assign w28868 = ~w28865 & ~w28867;
assign w28869 = ~w28853 & w28863;
assign w28870 = ~w28852 & w28869;
assign w28871 = w28853 & w28863;
assign w28872 = w28852 & w28871;
assign w28873 = ~w28870 & ~w28872;
assign w28874 = w28868 & w28873;
assign w28875 = w28768 & ~w28874;
assign w28876 = ~w28768 & w28874;
assign w28877 = ~w28875 & ~w28876;
assign w28878 = ~w28767 & w28877;
assign w28879 = w28767 & ~w28877;
assign w28880 = ~w28878 & ~w28879;
assign w28881 = w28753 & ~w28880;
assign w28882 = ~w28753 & w28880;
assign w28883 = ~w28881 & ~w28882;
assign w28884 = (~w28682 & ~w28684) | (~w28682 & w32293) | (~w28684 & w32293);
assign w28885 = ~w28883 & w28884;
assign w28886 = w28883 & ~w28884;
assign w28887 = ~w28885 & ~w28886;
assign w28888 = w7511 & w26766;
assign w28889 = w7192 & ~w21743;
assign w28890 = w7489 & w26476;
assign w28891 = w7193 & ~w26774;
assign w28892 = ~w28889 & ~w28890;
assign w28893 = ~w28888 & w28892;
assign w28894 = ~w28891 & w28893;
assign w28895 = a_11 & w28894;
assign w28896 = ~a_11 & ~w28894;
assign w28897 = ~w28895 & ~w28896;
assign w28898 = w28887 & ~w28897;
assign w28899 = ~w28887 & w28897;
assign w28900 = ~w28898 & ~w28899;
assign w28901 = w28739 & ~w28900;
assign w28902 = ~w28739 & w28900;
assign w28903 = ~w28901 & ~w28902;
assign w28904 = ~w28727 & ~w28903;
assign w28905 = w28727 & w28903;
assign w28906 = ~w28904 & ~w28905;
assign w28907 = ~w28521 & ~w28714;
assign w28908 = ~w28303 & w28907;
assign w28909 = w28306 & w28908;
assign w28910 = w27595 & w28909;
assign w28911 = ~w28309 & w28908;
assign w28912 = ~w28910 & ~w28911;
assign w28913 = ~w28528 & w28907;
assign w28914 = (~w28715 & w28528) | (~w28715 & w32294) | (w28528 & w32294);
assign w28915 = w28912 & w28914;
assign w28916 = ~w28906 & w28915;
assign w28917 = w28906 & ~w28915;
assign w28918 = ~w28916 & ~w28917;
assign w28919 = ~w28723 & ~w28918;
assign w28920 = w28723 & w28918;
assign w28921 = ~w28919 & ~w28920;
assign w28922 = w8276 & w27063;
assign w28923 = ~a_8 & ~w28922;
assign w28924 = w14078 & w27063;
assign w28925 = ~w28923 & ~w28924;
assign w28926 = ~w28885 & w28925;
assign w28927 = ~w28886 & ~w28925;
assign w28928 = ~w28926 & ~w28927;
assign w28929 = w28897 & w28925;
assign w28930 = ~w28886 & w28929;
assign w28931 = ~w28897 & ~w28925;
assign w28932 = ~w28885 & w28931;
assign w28933 = ~w28930 & ~w28932;
assign w28934 = ~w28928 & w28933;
assign w28935 = ~w28751 & ~w28881;
assign w28936 = w7511 & w27059;
assign w28937 = w7489 & w26766;
assign w28938 = w7192 & w26476;
assign w28939 = w7193 & w27068;
assign w28940 = ~w28937 & ~w28938;
assign w28941 = ~w28936 & w28940;
assign w28942 = ~w28939 & w28941;
assign w28943 = ~a_11 & w28942;
assign w28944 = a_11 & ~w28942;
assign w28945 = ~w28943 & ~w28944;
assign w28946 = w28935 & ~w28945;
assign w28947 = ~w28935 & w28945;
assign w28948 = ~w28946 & ~w28947;
assign w28949 = w6996 & ~w21743;
assign w28950 = w6998 & w21746;
assign w28951 = w6446 & w21752;
assign w28952 = w6447 & w22065;
assign w28953 = ~w28950 & ~w28951;
assign w28954 = ~w28949 & w28953;
assign w28955 = ~w28952 & w28954;
assign w28956 = ~a_14 & w28955;
assign w28957 = a_14 & ~w28955;
assign w28958 = ~w28956 & ~w28957;
assign w28959 = ~w28766 & w28877;
assign w28960 = ~w28765 & ~w28959;
assign w28961 = w28958 & ~w28960;
assign w28962 = ~w28958 & w28960;
assign w28963 = ~w28961 & ~w28962;
assign w28964 = ~w28768 & w28868;
assign w28965 = w28873 & ~w28964;
assign w28966 = w6304 & w21755;
assign w28967 = w6061 & ~w21757;
assign w28968 = w6059 & w22039;
assign w28969 = w6063 & ~w25675;
assign w28970 = ~w28967 & ~w28968;
assign w28971 = ~w28966 & w28970;
assign w28972 = ~w28969 & w28971;
assign w28973 = ~a_17 & w28972;
assign w28974 = a_17 & ~w28972;
assign w28975 = ~w28973 & ~w28974;
assign w28976 = ~w28965 & w28975;
assign w28977 = w28873 & ~w28975;
assign w28978 = ~w28964 & w28977;
assign w28979 = ~w28976 & ~w28978;
assign w28980 = w5816 & w22032;
assign w28981 = w5308 & w21762;
assign w28982 = w5818 & ~w22035;
assign w28983 = w5309 & w24756;
assign w28984 = ~w28980 & ~w28981;
assign w28985 = ~w28982 & w28984;
assign w28986 = ~w28983 & w28985;
assign w28987 = a_20 & ~w28986;
assign w28988 = ~a_20 & w28986;
assign w28989 = ~w28987 & ~w28988;
assign w28990 = ~w28846 & ~w28989;
assign w28991 = w28853 & ~w28989;
assign w28992 = w28851 & w28991;
assign w28993 = ~w28990 & ~w28992;
assign w28994 = w28851 & w28853;
assign w28995 = w28846 & w28989;
assign w28996 = ~w28994 & w28995;
assign w28997 = w28993 & ~w28996;
assign w28998 = ~w28812 & ~w28815;
assign w28999 = ~w28796 & ~w28799;
assign w29000 = w4068 & ~w21968;
assign w29001 = w3957 & w21934;
assign w29002 = w4446 & ~w21973;
assign w29003 = ~w29000 & ~w29001;
assign w29004 = ~w29002 & w29003;
assign w29005 = (w29004 & w22930) | (w29004 & w32295) | (w22930 & w32295);
assign w29006 = ~a_29 & w29005;
assign w29007 = a_29 & ~w29005;
assign w29008 = ~w29006 & ~w29007;
assign w29009 = ~w28782 & ~w28785;
assign w29010 = ~w23031 & w32296;
assign w29011 = w668 & ~w21940;
assign w29012 = w1399 & w21951;
assign w29013 = w1327 & ~w21945;
assign w29014 = ~w29011 & ~w29012;
assign w29015 = ~w29013 & w29014;
assign w29016 = ~w29010 & w29015;
assign w29017 = w569 & w1419;
assign w29018 = w1633 & w2729;
assign w29019 = w3567 & w3674;
assign w29020 = w14006 & w29019;
assign w29021 = w29017 & w29018;
assign w29022 = w2058 & w29021;
assign w29023 = w6140 & w29020;
assign w29024 = w6634 & w29023;
assign w29025 = w3745 & w29022;
assign w29026 = w29024 & w29025;
assign w29027 = ~w172 & ~w789;
assign w29028 = w367 & w29027;
assign w29029 = w809 & w934;
assign w29030 = w2405 & w2570;
assign w29031 = w3155 & w4257;
assign w29032 = w15222 & w29031;
assign w29033 = w29029 & w29030;
assign w29034 = w1455 & w29028;
assign w29035 = w2434 & w6613;
assign w29036 = w29034 & w29035;
assign w29037 = w29032 & w29033;
assign w29038 = w1946 & w29037;
assign w29039 = w2369 & w29036;
assign w29040 = w29038 & w29039;
assign w29041 = w1847 & w29040;
assign w29042 = w29026 & w29041;
assign w29043 = w29016 & ~w29042;
assign w29044 = ~w29016 & w29042;
assign w29045 = ~w29043 & ~w29044;
assign w29046 = ~w29009 & ~w29045;
assign w29047 = w29009 & w29045;
assign w29048 = ~w29046 & ~w29047;
assign w29049 = w29008 & ~w29048;
assign w29050 = ~w29008 & w29048;
assign w29051 = ~w29049 & ~w29050;
assign w29052 = w28999 & ~w29051;
assign w29053 = ~w28999 & w29051;
assign w29054 = ~w29052 & ~w29053;
assign w29055 = w4666 & w22007;
assign w29056 = w4638 & ~w21992;
assign w29057 = ~w518 & w21985;
assign w29058 = w1226 & w23580;
assign w29059 = ~w29056 & ~w29057;
assign w29060 = ~w29055 & w29059;
assign w29061 = ~w29058 & w29060;
assign w29062 = a_26 & w29061;
assign w29063 = ~a_26 & ~w29061;
assign w29064 = ~w29062 & ~w29063;
assign w29065 = w29054 & w29064;
assign w29066 = ~w29054 & ~w29064;
assign w29067 = ~w29065 & ~w29066;
assign w29068 = w28998 & ~w29067;
assign w29069 = ~w28998 & w29067;
assign w29070 = ~w29068 & ~w29069;
assign w29071 = w5286 & w21771;
assign w29072 = w5016 & w22014;
assign w29073 = w5080 & ~w22020;
assign w29074 = w5017 & w24295;
assign w29075 = ~w29072 & ~w29073;
assign w29076 = ~w29071 & w29075;
assign w29077 = ~w29074 & w29076;
assign w29078 = ~a_23 & w29077;
assign w29079 = a_23 & ~w29077;
assign w29080 = ~w29078 & ~w29079;
assign w29081 = w29070 & w29080;
assign w29082 = ~w29070 & ~w29080;
assign w29083 = ~w29081 & ~w29082;
assign w29084 = ~w28828 & ~w28831;
assign w29085 = ~w28829 & ~w29084;
assign w29086 = ~w29083 & ~w29085;
assign w29087 = w29083 & w29085;
assign w29088 = ~w29086 & ~w29087;
assign w29089 = ~w28997 & w29088;
assign w29090 = w28997 & ~w29088;
assign w29091 = ~w29089 & ~w29090;
assign w29092 = ~w28979 & w29091;
assign w29093 = w28979 & ~w29091;
assign w29094 = ~w29092 & ~w29093;
assign w29095 = w28963 & w29094;
assign w29096 = ~w28963 & ~w29094;
assign w29097 = ~w29095 & ~w29096;
assign w29098 = w28948 & ~w29097;
assign w29099 = ~w28948 & w29097;
assign w29100 = ~w29098 & ~w29099;
assign w29101 = ~w28934 & ~w29100;
assign w29102 = w28934 & w29100;
assign w29103 = ~w29101 & ~w29102;
assign w29104 = ~w28738 & ~w28900;
assign w29105 = ~w28737 & ~w29104;
assign w29106 = ~w29103 & ~w29105;
assign w29107 = w29103 & w29105;
assign w29108 = ~w29106 & ~w29107;
assign w29109 = w28906 & w29108;
assign w29110 = w28914 & w29109;
assign w29111 = w28912 & w29110;
assign w29112 = ~w28904 & w29108;
assign w29113 = w28904 & ~w29108;
assign w29114 = ~w29112 & ~w29113;
assign w29115 = ~w28906 & ~w29114;
assign w29116 = (w29115 & ~w28912) | (w29115 & w32297) | (~w28912 & w32297);
assign w29117 = ~w29111 & ~w29116;
assign w29118 = w28723 & ~w29117;
assign w29119 = ~w28917 & ~w29114;
assign w29120 = w28917 & ~w29108;
assign w29121 = ~w29119 & ~w29120;
assign w29122 = ~w28920 & w29121;
assign w29123 = ~w29118 & ~w29122;
assign w29124 = (~w29106 & w28904) | (~w29106 & w32298) | (w28904 & w32298);
assign w29125 = ~w29109 & ~w29124;
assign w29126 = w28926 & ~w28930;
assign w29127 = ~w29101 & ~w29126;
assign w29128 = ~w28947 & ~w29097;
assign w29129 = ~w28946 & ~w29128;
assign w29130 = a_8 & w29129;
assign w29131 = ~a_8 & ~w29129;
assign w29132 = ~w29130 & ~w29131;
assign w29133 = w7511 & w27063;
assign w29134 = w7192 & w26766;
assign w29135 = w7489 & w27059;
assign w29136 = w7193 & w27094;
assign w29137 = ~w29134 & ~w29135;
assign w29138 = ~w29133 & w29137;
assign w29139 = ~w29136 & w29138;
assign w29140 = ~a_11 & w29139;
assign w29141 = a_11 & ~w29139;
assign w29142 = ~w29140 & ~w29141;
assign w29143 = ~w28961 & ~w29094;
assign w29144 = ~w28962 & ~w29143;
assign w29145 = w29142 & w29144;
assign w29146 = ~w29142 & ~w29144;
assign w29147 = ~w29145 & ~w29146;
assign w29148 = w28993 & w29088;
assign w29149 = ~w28996 & ~w29148;
assign w29150 = w6304 & w21752;
assign w29151 = w6059 & ~w21757;
assign w29152 = w6061 & w21755;
assign w29153 = w6063 & w26166;
assign w29154 = ~w29151 & ~w29152;
assign w29155 = ~w29150 & w29154;
assign w29156 = ~w29153 & w29155;
assign w29157 = ~a_17 & w29156;
assign w29158 = a_17 & ~w29156;
assign w29159 = ~w29157 & ~w29158;
assign w29160 = w29149 & ~w29159;
assign w29161 = ~w29149 & w29159;
assign w29162 = ~w29160 & ~w29161;
assign w29163 = ~w29081 & ~w29087;
assign w29164 = w5816 & w22039;
assign w29165 = w5308 & ~w22035;
assign w29166 = w5818 & w22032;
assign w29167 = w5309 & w24962;
assign w29168 = ~w29165 & ~w29166;
assign w29169 = ~w29164 & w29168;
assign w29170 = ~w29167 & w29169;
assign w29171 = ~a_20 & w29170;
assign w29172 = a_20 & ~w29170;
assign w29173 = ~w29171 & ~w29172;
assign w29174 = ~w29163 & w29173;
assign w29175 = w29163 & ~w29173;
assign w29176 = ~w29174 & ~w29175;
assign w29177 = ~w29066 & ~w29069;
assign w29178 = w4666 & w22014;
assign w29179 = w4638 & w22007;
assign w29180 = ~w518 & ~w21992;
assign w29181 = w1226 & w23398;
assign w29182 = ~w29179 & ~w29180;
assign w29183 = ~w29178 & w29182;
assign w29184 = ~w29181 & w29183;
assign w29185 = a_26 & ~w29184;
assign w29186 = ~a_26 & w29184;
assign w29187 = ~w29185 & ~w29186;
assign w29188 = w4446 & w21985;
assign w29189 = w3957 & ~w21968;
assign w29190 = w4068 & ~w21973;
assign w29191 = w4070 & w23553;
assign w29192 = ~w29188 & ~w29189;
assign w29193 = ~w29190 & w29192;
assign w29194 = ~w29191 & w29193;
assign w29195 = ~a_29 & w29194;
assign w29196 = a_29 & ~w29194;
assign w29197 = ~w29195 & ~w29196;
assign w29198 = ~w29187 & ~w29197;
assign w29199 = w29187 & w29197;
assign w29200 = ~w29198 & ~w29199;
assign w29201 = ~w29050 & ~w29053;
assign w29202 = ~w50 & w253;
assign w29203 = w728 & w1113;
assign w29204 = w2216 & w2845;
assign w29205 = w3329 & w29204;
assign w29206 = w29202 & w29203;
assign w29207 = w985 & w4851;
assign w29208 = w29206 & w29207;
assign w29209 = w3684 & w29205;
assign w29210 = w29208 & w29209;
assign w29211 = w2735 & w29210;
assign w29212 = ~w76 & ~w458;
assign w29213 = ~w1051 & w29212;
assign w29214 = w2569 & w5558;
assign w29215 = w6117 & w29214;
assign w29216 = w29213 & w29215;
assign w29217 = ~w292 & ~w363;
assign w29218 = ~w389 & ~w431;
assign w29219 = ~w589 & ~w694;
assign w29220 = w29218 & w29219;
assign w29221 = w3910 & w29217;
assign w29222 = w5844 & w6742;
assign w29223 = w29221 & w29222;
assign w29224 = w13061 & w29220;
assign w29225 = w29223 & w29224;
assign w29226 = w4252 & w29225;
assign w29227 = w29216 & w29226;
assign w29228 = w4150 & w29227;
assign w29229 = w29211 & w29228;
assign w29230 = w13548 & w29229;
assign w29231 = w29042 & ~w29230;
assign w29232 = ~w29042 & w29230;
assign w29233 = ~w29231 & ~w29232;
assign w29234 = w29009 & ~w29044;
assign w29235 = ~w29043 & ~w29234;
assign w29236 = w29233 & ~w29235;
assign w29237 = ~w29233 & w29235;
assign w29238 = ~w29236 & ~w29237;
assign w29239 = w668 & w21934;
assign w29240 = w1399 & ~w21945;
assign w29241 = w1327 & ~w21940;
assign w29242 = w1478 & w23310;
assign w29243 = ~w29239 & ~w29240;
assign w29244 = ~w29241 & w29243;
assign w29245 = ~w29242 & w29244;
assign w29246 = ~w29238 & ~w29245;
assign w29247 = w29238 & w29245;
assign w29248 = ~w29246 & ~w29247;
assign w29249 = w29201 & w29248;
assign w29250 = ~w29201 & ~w29248;
assign w29251 = ~w29249 & ~w29250;
assign w29252 = w29200 & ~w29251;
assign w29253 = ~w29200 & w29251;
assign w29254 = ~w29252 & ~w29253;
assign w29255 = w29177 & w29254;
assign w29256 = ~w29177 & ~w29254;
assign w29257 = ~w29255 & ~w29256;
assign w29258 = w5080 & w21771;
assign w29259 = w5286 & w21762;
assign w29260 = w5016 & ~w22020;
assign w29261 = w5017 & w24502;
assign w29262 = ~w29259 & ~w29260;
assign w29263 = ~w29258 & w29262;
assign w29264 = ~w29261 & w29263;
assign w29265 = ~a_23 & w29264;
assign w29266 = a_23 & ~w29264;
assign w29267 = ~w29265 & ~w29266;
assign w29268 = w29257 & ~w29267;
assign w29269 = ~w29257 & w29267;
assign w29270 = ~w29268 & ~w29269;
assign w29271 = w29176 & ~w29270;
assign w29272 = ~w29176 & w29270;
assign w29273 = ~w29271 & ~w29272;
assign w29274 = w29162 & w29273;
assign w29275 = ~w29162 & ~w29273;
assign w29276 = ~w29274 & ~w29275;
assign w29277 = ~w28978 & ~w29091;
assign w29278 = ~w28976 & ~w29277;
assign w29279 = w6996 & w26476;
assign w29280 = w6998 & ~w21743;
assign w29281 = w6446 & w21746;
assign w29282 = w6447 & w26489;
assign w29283 = ~w29280 & ~w29281;
assign w29284 = ~w29279 & w29283;
assign w29285 = ~w29282 & w29284;
assign w29286 = a_14 & ~w29285;
assign w29287 = ~a_14 & w29285;
assign w29288 = ~w29286 & ~w29287;
assign w29289 = w29278 & ~w29288;
assign w29290 = ~w29278 & w29288;
assign w29291 = ~w29289 & ~w29290;
assign w29292 = w29276 & w29291;
assign w29293 = ~w29276 & ~w29291;
assign w29294 = ~w29292 & ~w29293;
assign w29295 = w29147 & ~w29294;
assign w29296 = ~w29147 & w29294;
assign w29297 = ~w29295 & ~w29296;
assign w29298 = w29132 & ~w29297;
assign w29299 = ~w29132 & w29297;
assign w29300 = ~w29298 & ~w29299;
assign w29301 = w29127 & ~w29300;
assign w29302 = ~w29127 & w29300;
assign w29303 = ~w29301 & ~w29302;
assign w29304 = ~w29125 & w29303;
assign w29305 = w29125 & ~w29303;
assign w29306 = ~w29304 & ~w29305;
assign w29307 = w28912 & w32299;
assign w29308 = (w29306 & ~w28912) | (w29306 & w32300) | (~w28912 & w32300);
assign w29309 = ~w29307 & ~w29308;
assign w29310 = ~w29118 & w29309;
assign w29311 = ~w29117 & ~w29309;
assign w29312 = w28723 & w29311;
assign w29313 = ~w29310 & ~w29312;
assign w29314 = w7489 & w27063;
assign w29315 = w7192 & w27059;
assign w29316 = w7193 & ~w27350;
assign w29317 = ~w29314 & ~w29315;
assign w29318 = ~w29316 & w29317;
assign w29319 = a_11 & ~w29318;
assign w29320 = ~a_11 & w29318;
assign w29321 = ~w29319 & ~w29320;
assign w29322 = ~w29145 & ~w29294;
assign w29323 = ~w29146 & ~w29322;
assign w29324 = w29321 & w29323;
assign w29325 = ~w29321 & ~w29323;
assign w29326 = ~w29324 & ~w29325;
assign w29327 = w6996 & w26766;
assign w29328 = w6446 & ~w21743;
assign w29329 = w6998 & w26476;
assign w29330 = w6447 & ~w26774;
assign w29331 = ~w29328 & ~w29329;
assign w29332 = ~w29327 & w29331;
assign w29333 = ~w29330 & w29332;
assign w29334 = a_14 & w29333;
assign w29335 = ~a_14 & ~w29333;
assign w29336 = ~w29334 & ~w29335;
assign w29337 = ~w29276 & ~w29290;
assign w29338 = ~w29289 & ~w29337;
assign w29339 = ~w29336 & w29338;
assign w29340 = w29336 & ~w29338;
assign w29341 = ~w29339 & ~w29340;
assign w29342 = ~w29161 & ~w29273;
assign w29343 = w6304 & w21746;
assign w29344 = w6061 & w21752;
assign w29345 = w6059 & w21755;
assign w29346 = w6063 & ~w25700;
assign w29347 = ~w29344 & ~w29345;
assign w29348 = ~w29343 & w29347;
assign w29349 = ~w29346 & w29348;
assign w29350 = ~a_17 & w29349;
assign w29351 = a_17 & ~w29349;
assign w29352 = ~w29350 & ~w29351;
assign w29353 = ~w29160 & w29352;
assign w29354 = ~w29342 & w29353;
assign w29355 = ~w29161 & ~w29352;
assign w29356 = ~w29274 & w29355;
assign w29357 = ~w29354 & ~w29356;
assign w29358 = ~w29255 & ~w29268;
assign w29359 = ~w29198 & ~w29252;
assign w29360 = w4666 & ~w22020;
assign w29361 = ~w518 & w22007;
assign w29362 = w4638 & w22014;
assign w29363 = w1226 & w24122;
assign w29364 = ~w29361 & ~w29362;
assign w29365 = ~w29360 & w29364;
assign w29366 = ~w29363 & w29365;
assign w29367 = a_26 & ~w29366;
assign w29368 = ~a_26 & w29366;
assign w29369 = ~w29367 & ~w29368;
assign w29370 = w29359 & w29369;
assign w29371 = ~w29359 & ~w29369;
assign w29372 = ~w29370 & ~w29371;
assign w29373 = ~w29246 & ~w29249;
assign w29374 = ~w118 & w1658;
assign w29375 = ~w356 & ~w470;
assign w29376 = w1405 & w29375;
assign w29377 = w3014 & w4346;
assign w29378 = w29376 & w29377;
assign w29379 = w1642 & w2381;
assign w29380 = w13532 & w29374;
assign w29381 = w29379 & w29380;
assign w29382 = w384 & w29378;
assign w29383 = w3738 & w29382;
assign w29384 = w29381 & w29383;
assign w29385 = w3151 & w29384;
assign w29386 = w1753 & w2465;
assign w29387 = w29385 & w29386;
assign w29388 = ~w29042 & ~w29387;
assign w29389 = w29042 & w29387;
assign w29390 = ~w29388 & ~w29389;
assign w29391 = ~a_8 & w29390;
assign w29392 = a_8 & ~w29390;
assign w29393 = ~w29391 & ~w29392;
assign w29394 = ~w29043 & ~w29232;
assign w29395 = ~w29234 & w29394;
assign w29396 = ~w29231 & ~w29395;
assign w29397 = w668 & ~w21968;
assign w29398 = w1327 & w21934;
assign w29399 = w1399 & ~w21940;
assign w29400 = w1478 & ~w23366;
assign w29401 = ~w29398 & ~w29399;
assign w29402 = ~w29397 & w29401;
assign w29403 = ~w29400 & w29402;
assign w29404 = ~w29396 & ~w29403;
assign w29405 = w29396 & w29403;
assign w29406 = ~w29404 & ~w29405;
assign w29407 = w29393 & w29406;
assign w29408 = ~w29393 & ~w29406;
assign w29409 = ~w29407 & ~w29408;
assign w29410 = w4446 & ~w21992;
assign w29411 = w4068 & w21985;
assign w29412 = w3957 & ~w21973;
assign w29413 = w4070 & ~w23930;
assign w29414 = ~w29411 & ~w29412;
assign w29415 = ~w29410 & w29414;
assign w29416 = ~w29413 & w29415;
assign w29417 = a_29 & ~w29416;
assign w29418 = ~a_29 & w29416;
assign w29419 = ~w29417 & ~w29418;
assign w29420 = w29409 & w29419;
assign w29421 = ~w29409 & ~w29419;
assign w29422 = ~w29420 & ~w29421;
assign w29423 = w29373 & ~w29422;
assign w29424 = ~w29373 & w29422;
assign w29425 = ~w29423 & ~w29424;
assign w29426 = w5016 & w21771;
assign w29427 = w5080 & w21762;
assign w29428 = w5286 & ~w22035;
assign w29429 = w5017 & w24529;
assign w29430 = ~w29427 & ~w29428;
assign w29431 = ~w29426 & w29430;
assign w29432 = ~w29429 & w29431;
assign w29433 = ~a_23 & w29432;
assign w29434 = a_23 & ~w29432;
assign w29435 = ~w29433 & ~w29434;
assign w29436 = w29425 & ~w29435;
assign w29437 = ~w29425 & w29435;
assign w29438 = ~w29436 & ~w29437;
assign w29439 = w29372 & w29438;
assign w29440 = ~w29372 & ~w29438;
assign w29441 = ~w29439 & ~w29440;
assign w29442 = w29358 & ~w29441;
assign w29443 = ~w29358 & w29441;
assign w29444 = ~w29442 & ~w29443;
assign w29445 = w5816 & ~w21757;
assign w29446 = w5818 & w22039;
assign w29447 = w5308 & w22032;
assign w29448 = w5309 & ~w25205;
assign w29449 = ~w29446 & ~w29447;
assign w29450 = ~w29445 & w29449;
assign w29451 = ~w29448 & w29450;
assign w29452 = a_20 & ~w29451;
assign w29453 = ~a_20 & w29451;
assign w29454 = ~w29452 & ~w29453;
assign w29455 = w29444 & w29454;
assign w29456 = ~w29444 & ~w29454;
assign w29457 = ~w29455 & ~w29456;
assign w29458 = ~w29175 & ~w29270;
assign w29459 = ~w29174 & ~w29458;
assign w29460 = w29457 & ~w29459;
assign w29461 = ~w29457 & w29459;
assign w29462 = ~w29460 & ~w29461;
assign w29463 = ~w29357 & w29462;
assign w29464 = w29357 & ~w29462;
assign w29465 = ~w29463 & ~w29464;
assign w29466 = w29341 & ~w29465;
assign w29467 = ~w29341 & w29465;
assign w29468 = ~w29466 & ~w29467;
assign w29469 = w29326 & w29468;
assign w29470 = ~w29326 & ~w29468;
assign w29471 = ~w29469 & ~w29470;
assign w29472 = ~w29130 & ~w29298;
assign w29473 = w29471 & ~w29472;
assign w29474 = ~w29471 & w29472;
assign w29475 = ~w29473 & ~w29474;
assign w29476 = ~w29302 & ~w29475;
assign w29477 = ~w29304 & w29476;
assign w29478 = ~w28715 & ~w29124;
assign w29479 = (w29478 & w28528) | (w29478 & w32301) | (w28528 & w32301);
assign w29480 = w29476 & w29479;
assign w29481 = ~w29302 & ~w29473;
assign w29482 = w29478 & w29481;
assign w29483 = ~w28913 & w29482;
assign w29484 = w29125 & w29481;
assign w29485 = ~w29301 & ~w29474;
assign w29486 = ~w29473 & w29485;
assign w29487 = ~w29484 & w29486;
assign w29488 = (w29487 & ~w28912) | (w29487 & w32302) | (~w28912 & w32302);
assign w29489 = (~w29477 & ~w28912) | (~w29477 & w32630) | (~w28912 & w32630);
assign w29490 = ~w29488 & w29489;
assign w29491 = w29312 & w29490;
assign w29492 = ~w29312 & ~w29490;
assign w29493 = ~w29491 & ~w29492;
assign w29494 = ~w29324 & ~w29469;
assign w29495 = w7191 & w27063;
assign w29496 = ~a_11 & ~w29495;
assign w29497 = w13947 & w27063;
assign w29498 = ~w29496 & ~w29497;
assign w29499 = ~w29339 & w29465;
assign w29500 = ~w29340 & ~w29499;
assign w29501 = w29498 & w29500;
assign w29502 = ~w29498 & ~w29500;
assign w29503 = ~w29501 & ~w29502;
assign w29504 = ~w29354 & ~w29462;
assign w29505 = ~w29356 & ~w29504;
assign w29506 = w6996 & w27059;
assign w29507 = w6998 & w26766;
assign w29508 = w6446 & w26476;
assign w29509 = w6447 & w27068;
assign w29510 = ~w29507 & ~w29508;
assign w29511 = ~w29506 & w29510;
assign w29512 = ~w29509 & w29511;
assign w29513 = a_14 & ~w29512;
assign w29514 = ~a_14 & w29512;
assign w29515 = ~w29513 & ~w29514;
assign w29516 = ~w29505 & ~w29515;
assign w29517 = w29505 & w29515;
assign w29518 = ~w29516 & ~w29517;
assign w29519 = w6304 & ~w21743;
assign w29520 = w6061 & w21746;
assign w29521 = w6059 & w21752;
assign w29522 = w6063 & w22065;
assign w29523 = ~w29520 & ~w29521;
assign w29524 = ~w29519 & w29523;
assign w29525 = ~w29522 & w29524;
assign w29526 = ~a_17 & w29525;
assign w29527 = a_17 & ~w29525;
assign w29528 = ~w29526 & ~w29527;
assign w29529 = ~w29456 & ~w29459;
assign w29530 = ~w29455 & ~w29529;
assign w29531 = ~w29528 & w29530;
assign w29532 = w29528 & ~w29530;
assign w29533 = ~w29531 & ~w29532;
assign w29534 = w29435 & w29441;
assign w29535 = ~w29442 & ~w29534;
assign w29536 = w5816 & w21755;
assign w29537 = w5818 & ~w21757;
assign w29538 = w5308 & w22039;
assign w29539 = w5309 & ~w25675;
assign w29540 = ~w29537 & ~w29538;
assign w29541 = ~w29536 & w29540;
assign w29542 = ~w29539 & w29541;
assign w29543 = a_20 & ~w29542;
assign w29544 = ~a_20 & w29542;
assign w29545 = ~w29543 & ~w29544;
assign w29546 = ~w29535 & w29545;
assign w29547 = w29535 & ~w29545;
assign w29548 = ~w29546 & ~w29547;
assign w29549 = ~w29420 & ~w29424;
assign w29550 = ~w29404 & ~w29407;
assign w29551 = ~w29388 & ~w29391;
assign w29552 = ~w88 & ~w95;
assign w29553 = ~w626 & w29552;
assign w29554 = w990 & w1331;
assign w29555 = w2183 & w14576;
assign w29556 = w29554 & w29555;
assign w29557 = w906 & w29553;
assign w29558 = w2242 & w15165;
assign w29559 = w29557 & w29558;
assign w29560 = w13929 & w29556;
assign w29561 = w29559 & w29560;
assign w29562 = w5167 & w29561;
assign w29563 = w1582 & w29562;
assign w29564 = w3363 & w29563;
assign w29565 = w29551 & ~w29564;
assign w29566 = ~w29551 & w29564;
assign w29567 = ~w29565 & ~w29566;
assign w29568 = w1327 & ~w21968;
assign w29569 = w1399 & w21934;
assign w29570 = w668 & ~w21973;
assign w29571 = ~w29568 & ~w29569;
assign w29572 = ~w29570 & w29571;
assign w29573 = (w29572 & w22930) | (w29572 & w32303) | (w22930 & w32303);
assign w29574 = w29567 & w29573;
assign w29575 = ~w29567 & ~w29573;
assign w29576 = ~w29574 & ~w29575;
assign w29577 = w4446 & w22007;
assign w29578 = w4068 & ~w21992;
assign w29579 = w3957 & w21985;
assign w29580 = w4070 & w23580;
assign w29581 = ~w29578 & ~w29579;
assign w29582 = ~w29577 & w29581;
assign w29583 = ~w29580 & w29582;
assign w29584 = a_29 & ~w29583;
assign w29585 = ~a_29 & w29583;
assign w29586 = ~w29584 & ~w29585;
assign w29587 = w29576 & ~w29586;
assign w29588 = ~w29576 & w29586;
assign w29589 = ~w29587 & ~w29588;
assign w29590 = ~w29550 & w29589;
assign w29591 = w29550 & ~w29589;
assign w29592 = ~w29590 & ~w29591;
assign w29593 = w4666 & w21771;
assign w29594 = ~w518 & w22014;
assign w29595 = w4638 & ~w22020;
assign w29596 = w1226 & w24295;
assign w29597 = ~w29594 & ~w29595;
assign w29598 = ~w29593 & w29597;
assign w29599 = ~w29596 & w29598;
assign w29600 = a_26 & w29599;
assign w29601 = ~a_26 & ~w29599;
assign w29602 = ~w29600 & ~w29601;
assign w29603 = ~w29592 & w29602;
assign w29604 = w29592 & ~w29602;
assign w29605 = ~w29603 & ~w29604;
assign w29606 = w29549 & w29605;
assign w29607 = ~w29549 & ~w29605;
assign w29608 = ~w29606 & ~w29607;
assign w29609 = ~w29371 & w29425;
assign w29610 = w5286 & w22032;
assign w29611 = w5016 & w21762;
assign w29612 = w5080 & ~w22035;
assign w29613 = w5017 & w24756;
assign w29614 = ~w29610 & ~w29611;
assign w29615 = ~w29612 & w29614;
assign w29616 = ~w29613 & w29615;
assign w29617 = a_23 & ~w29616;
assign w29618 = ~a_23 & w29616;
assign w29619 = ~w29617 & ~w29618;
assign w29620 = ~w29370 & ~w29619;
assign w29621 = ~w29609 & w29620;
assign w29622 = ~w29370 & ~w29609;
assign w29623 = w29619 & ~w29622;
assign w29624 = ~w29621 & ~w29623;
assign w29625 = w29608 & ~w29624;
assign w29626 = ~w29608 & w29624;
assign w29627 = ~w29625 & ~w29626;
assign w29628 = w29548 & w29627;
assign w29629 = ~w29548 & ~w29627;
assign w29630 = ~w29628 & ~w29629;
assign w29631 = w29533 & ~w29630;
assign w29632 = ~w29533 & w29630;
assign w29633 = ~w29631 & ~w29632;
assign w29634 = ~w29518 & w29633;
assign w29635 = w29518 & ~w29633;
assign w29636 = ~w29634 & ~w29635;
assign w29637 = w29503 & w29636;
assign w29638 = ~w29503 & ~w29636;
assign w29639 = ~w29637 & ~w29638;
assign w29640 = ~w29494 & w29639;
assign w29641 = w29481 & ~w29640;
assign w29642 = ~w29109 & w32304;
assign w29643 = w29494 & ~w29639;
assign w29644 = ~w29473 & ~w29640;
assign w29645 = ~w29485 & w29644;
assign w29646 = ~w29643 & ~w29645;
assign w29647 = ~w29642 & w29646;
assign w29648 = ~w29640 & w29647;
assign w29649 = ~w29640 & ~w29643;
assign w29650 = ~w29473 & ~w29485;
assign w29651 = ~w29649 & w29650;
assign w29652 = ~w29648 & ~w29651;
assign w29653 = ~w29481 & w29649;
assign w29654 = ~w29650 & w29653;
assign w29655 = ~w29651 & ~w29654;
assign w29656 = w29479 & w29655;
assign w29657 = (~w29652 & ~w28912) | (~w29652 & w32305) | (~w28912 & w32305);
assign w29658 = w29484 & ~w29649;
assign w29659 = ~w28913 & w32306;
assign w29660 = (~w29658 & ~w28912) | (~w29658 & w32307) | (~w28912 & w32307);
assign w29661 = ~w29657 & w29660;
assign w29662 = w29490 & w29661;
assign w29663 = w29311 & w29662;
assign w29664 = w28723 & w29663;
assign w29665 = ~w29491 & ~w29661;
assign w29666 = ~w29664 & ~w29665;
assign w29667 = ~w28715 & w32304;
assign w29668 = (w29667 & w28528) | (w29667 & w32308) | (w28528 & w32308);
assign w29669 = w29647 & w29668;
assign w29670 = ~w29501 & ~w29637;
assign w29671 = ~w29517 & w29633;
assign w29672 = ~w29516 & ~w29671;
assign w29673 = a_11 & w29672;
assign w29674 = ~a_11 & ~w29672;
assign w29675 = ~w29673 & ~w29674;
assign w29676 = w6996 & w27063;
assign w29677 = w6998 & w27059;
assign w29678 = w6446 & w26766;
assign w29679 = w6447 & w27094;
assign w29680 = ~w29677 & ~w29678;
assign w29681 = ~w29676 & w29680;
assign w29682 = ~w29679 & w29681;
assign w29683 = a_14 & ~w29682;
assign w29684 = ~a_14 & w29682;
assign w29685 = ~w29683 & ~w29684;
assign w29686 = ~w29531 & w29630;
assign w29687 = ~w29532 & ~w29686;
assign w29688 = w29685 & ~w29687;
assign w29689 = ~w29685 & w29687;
assign w29690 = ~w29688 & ~w29689;
assign w29691 = w6061 & ~w21743;
assign w29692 = w6059 & w21746;
assign w29693 = w6304 & w26476;
assign w29694 = ~w29691 & ~w29692;
assign w29695 = ~w29693 & w29694;
assign w29696 = ~a_17 & w29695;
assign w29697 = (w29696 & ~w26489) | (w29696 & w32309) | (~w26489 & w32309);
assign w29698 = a_17 & ~w29695;
assign w29699 = (~w29698 & ~w26489) | (~w29698 & w32310) | (~w26489 & w32310);
assign w29700 = ~w29697 & w29699;
assign w29701 = ~w29547 & w29627;
assign w29702 = ~w29546 & ~w29701;
assign w29703 = w29700 & ~w29702;
assign w29704 = ~w29546 & ~w29700;
assign w29705 = ~w29701 & w29704;
assign w29706 = ~w29703 & ~w29705;
assign w29707 = ~w29608 & ~w29621;
assign w29708 = ~w29623 & ~w29707;
assign w29709 = w5816 & w21752;
assign w29710 = w5308 & ~w21757;
assign w29711 = w5818 & w21755;
assign w29712 = w5309 & w26166;
assign w29713 = ~w29710 & ~w29711;
assign w29714 = ~w29709 & w29713;
assign w29715 = ~w29712 & w29714;
assign w29716 = a_20 & w29715;
assign w29717 = ~a_20 & ~w29715;
assign w29718 = ~w29716 & ~w29717;
assign w29719 = ~w29708 & ~w29718;
assign w29720 = w29708 & w29718;
assign w29721 = ~w29719 & ~w29720;
assign w29722 = ~w29588 & ~w29590;
assign w29723 = w4068 & w22007;
assign w29724 = w3957 & ~w21992;
assign w29725 = w4446 & w22014;
assign w29726 = ~w29723 & ~w29724;
assign w29727 = ~w29725 & w29726;
assign w29728 = (w29727 & ~w23398) | (w29727 & w32311) | (~w23398 & w32311);
assign w29729 = a_29 & ~w29728;
assign w29730 = ~a_29 & w29728;
assign w29731 = ~w29729 & ~w29730;
assign w29732 = w668 & w21985;
assign w29733 = w1399 & ~w21968;
assign w29734 = w1327 & ~w21973;
assign w29735 = w1478 & w23553;
assign w29736 = ~w29732 & ~w29733;
assign w29737 = ~w29734 & w29736;
assign w29738 = ~w29735 & w29737;
assign w29739 = ~w29731 & w29738;
assign w29740 = w29731 & ~w29738;
assign w29741 = ~w29739 & ~w29740;
assign w29742 = w520 & ~w541;
assign w29743 = w950 & w1109;
assign w29744 = w2193 & w2419;
assign w29745 = w2717 & w3274;
assign w29746 = w4158 & w4713;
assign w29747 = w29745 & w29746;
assign w29748 = w29743 & w29744;
assign w29749 = w2551 & w29742;
assign w29750 = w3771 & w29749;
assign w29751 = w29747 & w29748;
assign w29752 = w29750 & w29751;
assign w29753 = w14582 & w29752;
assign w29754 = w13531 & w29753;
assign w29755 = w5612 & w29026;
assign w29756 = w29754 & w29755;
assign w29757 = w29564 & ~w29756;
assign w29758 = ~w29564 & w29756;
assign w29759 = ~w29757 & ~w29758;
assign w29760 = ~w29565 & ~w29574;
assign w29761 = w29759 & w29760;
assign w29762 = ~w29759 & ~w29760;
assign w29763 = ~w29761 & ~w29762;
assign w29764 = w29741 & ~w29763;
assign w29765 = ~w29741 & w29763;
assign w29766 = ~w29764 & ~w29765;
assign w29767 = w29722 & w29766;
assign w29768 = ~w29722 & ~w29766;
assign w29769 = ~w29767 & ~w29768;
assign w29770 = w4638 & w21771;
assign w29771 = w4666 & w21762;
assign w29772 = ~w518 & ~w22020;
assign w29773 = w1226 & w24502;
assign w29774 = ~w29771 & ~w29772;
assign w29775 = ~w29770 & w29774;
assign w29776 = ~w29773 & w29775;
assign w29777 = ~a_26 & w29776;
assign w29778 = a_26 & ~w29776;
assign w29779 = ~w29777 & ~w29778;
assign w29780 = w29769 & w29779;
assign w29781 = ~w29769 & ~w29779;
assign w29782 = ~w29780 & ~w29781;
assign w29783 = w5286 & w22039;
assign w29784 = w5016 & ~w22035;
assign w29785 = w5080 & w22032;
assign w29786 = w5017 & w24962;
assign w29787 = ~w29784 & ~w29785;
assign w29788 = ~w29783 & w29787;
assign w29789 = ~w29786 & w29788;
assign w29790 = ~a_23 & w29789;
assign w29791 = a_23 & ~w29789;
assign w29792 = ~w29790 & ~w29791;
assign w29793 = w29782 & w29792;
assign w29794 = ~w29782 & ~w29792;
assign w29795 = ~w29793 & ~w29794;
assign w29796 = ~w29603 & ~w29606;
assign w29797 = ~w29795 & w29796;
assign w29798 = w29795 & ~w29796;
assign w29799 = ~w29797 & ~w29798;
assign w29800 = ~w29721 & w29799;
assign w29801 = w29721 & ~w29799;
assign w29802 = ~w29800 & ~w29801;
assign w29803 = w29706 & ~w29802;
assign w29804 = ~w29706 & w29802;
assign w29805 = ~w29803 & ~w29804;
assign w29806 = w29690 & ~w29805;
assign w29807 = ~w29690 & w29805;
assign w29808 = ~w29806 & ~w29807;
assign w29809 = w29675 & w29808;
assign w29810 = ~w29675 & ~w29808;
assign w29811 = ~w29809 & ~w29810;
assign w29812 = w29670 & ~w29811;
assign w29813 = ~w29670 & w29811;
assign w29814 = ~w29812 & ~w29813;
assign w29815 = w29647 & w29814;
assign w29816 = ~w29647 & ~w29814;
assign w29817 = ~w29815 & ~w29816;
assign w29818 = (~w29817 & ~w28912) | (~w29817 & w32312) | (~w28912 & w32312);
assign w29819 = w28912 & w32313;
assign w29820 = ~w29818 & ~w29819;
assign w29821 = w29664 & w29820;
assign w29822 = ~w29664 & ~w29820;
assign w29823 = ~w29821 & ~w29822;
assign w29824 = ~w29689 & ~w29805;
assign w29825 = ~w29688 & ~w29824;
assign w29826 = w5816 & w21746;
assign w29827 = w5818 & w21752;
assign w29828 = w5308 & w21755;
assign w29829 = w5309 & ~w25700;
assign w29830 = ~w29827 & ~w29828;
assign w29831 = ~w29826 & w29830;
assign w29832 = ~w29829 & w29831;
assign w29833 = ~a_20 & w29832;
assign w29834 = a_20 & ~w29832;
assign w29835 = ~w29833 & ~w29834;
assign w29836 = ~w29719 & w29799;
assign w29837 = ~w29720 & ~w29836;
assign w29838 = ~w29835 & ~w29837;
assign w29839 = w29835 & w29837;
assign w29840 = ~w29838 & ~w29839;
assign w29841 = w6304 & w26766;
assign w29842 = w6059 & ~w21743;
assign w29843 = w6061 & w26476;
assign w29844 = w6063 & ~w26774;
assign w29845 = ~w29842 & ~w29843;
assign w29846 = ~w29841 & w29845;
assign w29847 = ~w29844 & w29846;
assign w29848 = a_17 & w29847;
assign w29849 = ~a_17 & ~w29847;
assign w29850 = ~w29848 & ~w29849;
assign w29851 = ~w29793 & ~w29796;
assign w29852 = ~w29794 & ~w29851;
assign w29853 = ~w518 & w21771;
assign w29854 = w4638 & w21762;
assign w29855 = w4666 & ~w22035;
assign w29856 = w1226 & w24529;
assign w29857 = ~w29854 & ~w29855;
assign w29858 = ~w29853 & w29857;
assign w29859 = ~w29856 & w29858;
assign w29860 = a_26 & ~w29859;
assign w29861 = ~a_26 & w29859;
assign w29862 = ~w29860 & ~w29861;
assign w29863 = ~w29757 & ~w29761;
assign w29864 = ~w183 & ~w191;
assign w29865 = ~w287 & ~w870;
assign w29866 = w29864 & w29865;
assign w29867 = w390 & w2655;
assign w29868 = w6168 & w29867;
assign w29869 = w133 & w29866;
assign w29870 = w5366 & w13083;
assign w29871 = w29869 & w29870;
assign w29872 = w5377 & w29868;
assign w29873 = w29871 & w29872;
assign w29874 = w3012 & w29873;
assign w29875 = w2345 & w29874;
assign w29876 = w2328 & w3788;
assign w29877 = w29875 & w29876;
assign w29878 = ~w29564 & ~w29877;
assign w29879 = w29564 & w29877;
assign w29880 = ~w29878 & ~w29879;
assign w29881 = ~a_11 & w29880;
assign w29882 = a_11 & ~w29880;
assign w29883 = ~w29881 & ~w29882;
assign w29884 = w1399 & ~w21973;
assign w29885 = w1327 & w21985;
assign w29886 = w668 & ~w21992;
assign w29887 = ~w29884 & ~w29885;
assign w29888 = ~w29886 & w29887;
assign w29889 = (w29888 & w23930) | (w29888 & w32314) | (w23930 & w32314);
assign w29890 = w29883 & ~w29889;
assign w29891 = ~w29883 & w29889;
assign w29892 = ~w29890 & ~w29891;
assign w29893 = w29863 & ~w29892;
assign w29894 = ~w29863 & w29892;
assign w29895 = ~w29893 & ~w29894;
assign w29896 = ~w29740 & ~w29763;
assign w29897 = ~w29739 & ~w29896;
assign w29898 = w29895 & w29897;
assign w29899 = ~w29895 & ~w29897;
assign w29900 = ~w29898 & ~w29899;
assign w29901 = w4446 & ~w22020;
assign w29902 = w4068 & w22014;
assign w29903 = w3957 & w22007;
assign w29904 = w4070 & w24122;
assign w29905 = ~w29902 & ~w29903;
assign w29906 = ~w29901 & w29905;
assign w29907 = ~w29904 & w29906;
assign w29908 = a_29 & ~w29907;
assign w29909 = ~a_29 & w29907;
assign w29910 = ~w29908 & ~w29909;
assign w29911 = w29900 & w29910;
assign w29912 = ~w29900 & ~w29910;
assign w29913 = ~w29911 & ~w29912;
assign w29914 = w29862 & w29913;
assign w29915 = ~w29862 & ~w29913;
assign w29916 = ~w29914 & ~w29915;
assign w29917 = w5286 & ~w21757;
assign w29918 = w5016 & w22032;
assign w29919 = w5080 & w22039;
assign w29920 = w5017 & ~w25205;
assign w29921 = ~w29918 & ~w29919;
assign w29922 = ~w29917 & w29921;
assign w29923 = ~w29920 & w29922;
assign w29924 = a_23 & w29923;
assign w29925 = ~a_23 & ~w29923;
assign w29926 = ~w29924 & ~w29925;
assign w29927 = ~w29768 & ~w29780;
assign w29928 = ~w29926 & ~w29927;
assign w29929 = ~w29916 & w29928;
assign w29930 = ~w29926 & w29927;
assign w29931 = w29916 & w29930;
assign w29932 = ~w29929 & ~w29931;
assign w29933 = ~w29916 & ~w29927;
assign w29934 = w29916 & w29927;
assign w29935 = w29926 & ~w29933;
assign w29936 = ~w29934 & w29935;
assign w29937 = w29932 & ~w29936;
assign w29938 = w29852 & ~w29937;
assign w29939 = ~w29852 & w29937;
assign w29940 = ~w29938 & ~w29939;
assign w29941 = w29850 & ~w29940;
assign w29942 = w29840 & w29941;
assign w29943 = w29850 & w29940;
assign w29944 = ~w29840 & w29943;
assign w29945 = ~w29942 & ~w29944;
assign w29946 = ~w29850 & ~w29940;
assign w29947 = ~w29840 & w29946;
assign w29948 = ~w29839 & w29940;
assign w29949 = ~w29838 & ~w29850;
assign w29950 = w29948 & w29949;
assign w29951 = ~w29947 & ~w29950;
assign w29952 = w29945 & w29951;
assign w29953 = ~w29705 & w29802;
assign w29954 = ~w29703 & ~w29953;
assign w29955 = w6998 & w27063;
assign w29956 = w6446 & w27059;
assign w29957 = w6447 & ~w27350;
assign w29958 = ~w29955 & ~w29956;
assign w29959 = ~w29957 & w29958;
assign w29960 = a_14 & ~w29959;
assign w29961 = ~a_14 & w29959;
assign w29962 = ~w29960 & ~w29961;
assign w29963 = w29954 & ~w29962;
assign w29964 = ~w29954 & w29962;
assign w29965 = ~w29963 & ~w29964;
assign w29966 = w29952 & w29965;
assign w29967 = ~w29952 & ~w29965;
assign w29968 = ~w29966 & ~w29967;
assign w29969 = w29825 & ~w29968;
assign w29970 = ~w29825 & w29968;
assign w29971 = ~w29969 & ~w29970;
assign w29972 = ~w29673 & ~w29808;
assign w29973 = ~w29674 & ~w29972;
assign w29974 = w29971 & w29973;
assign w29975 = ~w29971 & ~w29973;
assign w29976 = ~w29974 & ~w29975;
assign w29977 = w29813 & w29976;
assign w29978 = ~w29812 & w29976;
assign w29979 = w29646 & w29978;
assign w29980 = ~w29642 & w29979;
assign w29981 = ~w29977 & ~w29980;
assign w29982 = w29668 & ~w29977;
assign w29983 = (~w29981 & ~w28912) | (~w29981 & w32315) | (~w28912 & w32315);
assign w29984 = ~w29813 & ~w29976;
assign w29985 = ~w29815 & w29984;
assign w29986 = w29668 & w29984;
assign w29987 = (~w29985 & ~w28912) | (~w29985 & w32316) | (~w28912 & w32316);
assign w29988 = ~w29983 & w29987;
assign w29989 = w29820 & w29988;
assign w29990 = w29664 & w29989;
assign w29991 = ~w29821 & ~w29988;
assign w29992 = ~w29990 & ~w29991;
assign w29993 = ~w29974 & ~w29977;
assign w29994 = w29667 & w29993;
assign w29995 = ~w28913 & w32317;
assign w29996 = w28912 & w29995;
assign w29997 = ~w29980 & w29993;
assign w29998 = w29962 & ~w29968;
assign w29999 = ~w29970 & ~w29998;
assign w30000 = w6445 & w27063;
assign w30001 = ~a_14 & ~w30000;
assign w30002 = w13585 & w27063;
assign w30003 = ~w30001 & ~w30002;
assign w30004 = ~w29951 & w30003;
assign w30005 = ~w29954 & w30003;
assign w30006 = w29945 & w30005;
assign w30007 = ~w30004 & ~w30006;
assign w30008 = w29945 & ~w29954;
assign w30009 = w29951 & ~w30003;
assign w30010 = ~w30008 & w30009;
assign w30011 = w30007 & ~w30010;
assign w30012 = ~w29852 & w29932;
assign w30013 = ~w29936 & ~w30012;
assign w30014 = w5816 & ~w21743;
assign w30015 = w5818 & w21746;
assign w30016 = w5308 & w21752;
assign w30017 = w5309 & w22065;
assign w30018 = ~w30015 & ~w30016;
assign w30019 = ~w30014 & w30018;
assign w30020 = ~w30017 & w30019;
assign w30021 = ~a_20 & w30020;
assign w30022 = a_20 & ~w30020;
assign w30023 = ~w30021 & ~w30022;
assign w30024 = w30013 & w30023;
assign w30025 = ~w30013 & ~w30023;
assign w30026 = ~w30024 & ~w30025;
assign w30027 = w5286 & w21755;
assign w30028 = w5080 & ~w21757;
assign w30029 = w5016 & w22039;
assign w30030 = w5017 & ~w25675;
assign w30031 = ~w30028 & ~w30029;
assign w30032 = ~w30027 & w30031;
assign w30033 = ~w30030 & w30032;
assign w30034 = a_23 & ~w30033;
assign w30035 = ~a_23 & w30033;
assign w30036 = ~w30034 & ~w30035;
assign w30037 = ~w29914 & w29927;
assign w30038 = ~w29915 & ~w30037;
assign w30039 = ~w29898 & ~w29910;
assign w30040 = ~w29899 & ~w30039;
assign w30041 = ~w29878 & ~w29881;
assign w30042 = w1778 & w2250;
assign w30043 = w419 & w753;
assign w30044 = w2263 & w2710;
assign w30045 = w3239 & w3347;
assign w30046 = w30044 & w30045;
assign w30047 = w1239 & w30043;
assign w30048 = w30042 & w30047;
assign w30049 = w13351 & w30046;
assign w30050 = w30048 & w30049;
assign w30051 = w27437 & w27949;
assign w30052 = w30050 & w30051;
assign w30053 = w13093 & w30052;
assign w30054 = w14593 & w30053;
assign w30055 = w30041 & ~w30054;
assign w30056 = ~w30041 & w30054;
assign w30057 = ~w30055 & ~w30056;
assign w30058 = w668 & w22007;
assign w30059 = w1327 & ~w21992;
assign w30060 = w1399 & w21985;
assign w30061 = w1478 & w23580;
assign w30062 = ~w30059 & ~w30060;
assign w30063 = ~w30058 & w30062;
assign w30064 = ~w30061 & w30063;
assign w30065 = ~w30057 & ~w30064;
assign w30066 = w30057 & w30064;
assign w30067 = ~w30065 & ~w30066;
assign w30068 = ~w29890 & ~w29894;
assign w30069 = w30067 & w30068;
assign w30070 = ~w30067 & ~w30068;
assign w30071 = ~w30069 & ~w30070;
assign w30072 = w4446 & w21771;
assign w30073 = w3957 & w22014;
assign w30074 = w4068 & ~w22020;
assign w30075 = w4070 & w24295;
assign w30076 = ~w30073 & ~w30074;
assign w30077 = ~w30072 & w30076;
assign w30078 = ~w30075 & w30077;
assign w30079 = ~a_29 & w30078;
assign w30080 = a_29 & ~w30078;
assign w30081 = ~w30079 & ~w30080;
assign w30082 = w30071 & ~w30081;
assign w30083 = ~w30071 & w30081;
assign w30084 = ~w30082 & ~w30083;
assign w30085 = w30040 & ~w30084;
assign w30086 = ~w30040 & w30084;
assign w30087 = ~w30085 & ~w30086;
assign w30088 = w4666 & w22032;
assign w30089 = ~w518 & w21762;
assign w30090 = w4638 & ~w22035;
assign w30091 = w1226 & w24756;
assign w30092 = ~w30088 & ~w30089;
assign w30093 = ~w30090 & w30092;
assign w30094 = ~w30091 & w30093;
assign w30095 = a_26 & ~w30094;
assign w30096 = ~a_26 & w30094;
assign w30097 = ~w30095 & ~w30096;
assign w30098 = w30087 & w30097;
assign w30099 = ~w30087 & ~w30097;
assign w30100 = ~w30098 & ~w30099;
assign w30101 = w30038 & w30100;
assign w30102 = ~w30038 & ~w30100;
assign w30103 = ~w30101 & ~w30102;
assign w30104 = w30036 & ~w30103;
assign w30105 = ~w30036 & w30103;
assign w30106 = ~w30104 & ~w30105;
assign w30107 = ~w30026 & w30106;
assign w30108 = w30026 & ~w30106;
assign w30109 = ~w30107 & ~w30108;
assign w30110 = w6061 & w26766;
assign w30111 = w6059 & w26476;
assign w30112 = w6304 & w27059;
assign w30113 = ~w30110 & ~w30111;
assign w30114 = ~w30112 & w30113;
assign w30115 = ~a_17 & w30114;
assign w30116 = (w30115 & ~w27068) | (w30115 & w32318) | (~w27068 & w32318);
assign w30117 = a_17 & ~w30114;
assign w30118 = (~w30117 & ~w27068) | (~w30117 & w32319) | (~w27068 & w32319);
assign w30119 = ~w30116 & w30118;
assign w30120 = ~w29838 & ~w29948;
assign w30121 = ~w30119 & ~w30120;
assign w30122 = ~w29838 & w30119;
assign w30123 = ~w29948 & w30122;
assign w30124 = ~w30121 & ~w30123;
assign w30125 = w30109 & ~w30124;
assign w30126 = ~w30109 & w30124;
assign w30127 = ~w30125 & ~w30126;
assign w30128 = w30011 & ~w30127;
assign w30129 = ~w30011 & w30127;
assign w30130 = ~w30128 & ~w30129;
assign w30131 = ~w29999 & w30130;
assign w30132 = w29999 & ~w30130;
assign w30133 = ~w30131 & ~w30132;
assign w30134 = w29997 & ~w30133;
assign w30135 = ~w29997 & w30133;
assign w30136 = ~w30134 & ~w30135;
assign w30137 = w29996 & ~w30136;
assign w30138 = ~w29996 & w30136;
assign w30139 = ~w30137 & ~w30138;
assign w30140 = ~w29990 & w30139;
assign w30141 = w29664 & w32320;
assign w30142 = ~w30140 & ~w30141;
assign w30143 = ~w30109 & ~w30123;
assign w30144 = ~w30121 & ~w30143;
assign w30145 = a_14 & w30144;
assign w30146 = ~a_14 & ~w30144;
assign w30147 = ~w30145 & ~w30146;
assign w30148 = ~w217 & ~w239;
assign w30149 = ~w368 & w30148;
assign w30150 = w1075 & w1128;
assign w30151 = w1405 & w2654;
assign w30152 = w3210 & w3911;
assign w30153 = w30151 & w30152;
assign w30154 = w30149 & w30150;
assign w30155 = w30153 & w30154;
assign w30156 = w1050 & w3020;
assign w30157 = w30155 & w30156;
assign w30158 = w601 & w830;
assign w30159 = w5530 & w30158;
assign w30160 = w2753 & w30157;
assign w30161 = w30159 & w30160;
assign w30162 = w4309 & w30161;
assign w30163 = w30054 & ~w30162;
assign w30164 = ~w30054 & w30162;
assign w30165 = ~w30163 & ~w30164;
assign w30166 = w668 & w22014;
assign w30167 = w1399 & ~w21992;
assign w30168 = w1327 & w22007;
assign w30169 = w1478 & w23398;
assign w30170 = ~w30167 & ~w30168;
assign w30171 = ~w30166 & w30170;
assign w30172 = ~w30169 & w30171;
assign w30173 = w30165 & ~w30172;
assign w30174 = ~w30165 & w30172;
assign w30175 = ~w30173 & ~w30174;
assign w30176 = ~w30055 & ~w30066;
assign w30177 = w30175 & w30176;
assign w30178 = ~w30175 & ~w30176;
assign w30179 = ~w30177 & ~w30178;
assign w30180 = ~w30070 & ~w30081;
assign w30181 = ~w30069 & ~w30180;
assign w30182 = w30179 & w30181;
assign w30183 = ~w30179 & ~w30181;
assign w30184 = ~w30182 & ~w30183;
assign w30185 = w4068 & w21771;
assign w30186 = w4446 & w21762;
assign w30187 = w3957 & ~w22020;
assign w30188 = w4070 & w24502;
assign w30189 = ~w30186 & ~w30187;
assign w30190 = ~w30185 & w30189;
assign w30191 = ~w30188 & w30190;
assign w30192 = a_29 & ~w30191;
assign w30193 = ~a_29 & w30191;
assign w30194 = ~w30192 & ~w30193;
assign w30195 = w30184 & w30194;
assign w30196 = ~w30184 & ~w30194;
assign w30197 = ~w30195 & ~w30196;
assign w30198 = w4666 & w22039;
assign w30199 = ~w518 & ~w22035;
assign w30200 = w4638 & w22032;
assign w30201 = w1226 & w24962;
assign w30202 = ~w30199 & ~w30200;
assign w30203 = ~w30198 & w30202;
assign w30204 = ~w30201 & w30203;
assign w30205 = a_26 & ~w30204;
assign w30206 = ~a_26 & w30204;
assign w30207 = ~w30205 & ~w30206;
assign w30208 = w30197 & w30207;
assign w30209 = ~w30197 & ~w30207;
assign w30210 = ~w30208 & ~w30209;
assign w30211 = w5080 & w21755;
assign w30212 = w5016 & ~w21757;
assign w30213 = w5286 & w21752;
assign w30214 = ~w30211 & ~w30212;
assign w30215 = ~w30213 & w30214;
assign w30216 = (w30215 & ~w26166) | (w30215 & w32321) | (~w26166 & w32321);
assign w30217 = ~a_23 & w30216;
assign w30218 = a_23 & ~w30216;
assign w30219 = ~w30217 & ~w30218;
assign w30220 = ~w30085 & ~w30097;
assign w30221 = ~w30086 & ~w30220;
assign w30222 = w30219 & w30221;
assign w30223 = ~w30219 & ~w30221;
assign w30224 = ~w30222 & ~w30223;
assign w30225 = w30210 & w30224;
assign w30226 = ~w30210 & ~w30224;
assign w30227 = ~w30225 & ~w30226;
assign w30228 = ~w30036 & ~w30101;
assign w30229 = ~w30102 & ~w30228;
assign w30230 = w30227 & w30229;
assign w30231 = ~w30227 & ~w30229;
assign w30232 = ~w30230 & ~w30231;
assign w30233 = w5816 & w26476;
assign w30234 = w5818 & ~w21743;
assign w30235 = w5308 & w21746;
assign w30236 = w5309 & w26489;
assign w30237 = ~w30234 & ~w30235;
assign w30238 = ~w30233 & w30237;
assign w30239 = ~w30236 & w30238;
assign w30240 = ~a_20 & w30239;
assign w30241 = a_20 & ~w30239;
assign w30242 = ~w30240 & ~w30241;
assign w30243 = w30232 & w30242;
assign w30244 = ~w30232 & ~w30242;
assign w30245 = ~w30243 & ~w30244;
assign w30246 = ~w30024 & ~w30108;
assign w30247 = w30245 & ~w30246;
assign w30248 = ~w30245 & w30246;
assign w30249 = ~w30247 & ~w30248;
assign w30250 = w6304 & w27063;
assign w30251 = w6061 & w27059;
assign w30252 = w6059 & w26766;
assign w30253 = w6063 & w27094;
assign w30254 = ~w30251 & ~w30252;
assign w30255 = ~w30250 & w30254;
assign w30256 = ~w30253 & w30255;
assign w30257 = ~a_17 & w30256;
assign w30258 = a_17 & ~w30256;
assign w30259 = ~w30257 & ~w30258;
assign w30260 = ~w30249 & w30259;
assign w30261 = w30249 & ~w30259;
assign w30262 = ~w30260 & ~w30261;
assign w30263 = w30147 & ~w30262;
assign w30264 = ~w30147 & w30262;
assign w30265 = ~w30263 & ~w30264;
assign w30266 = w30007 & ~w30128;
assign w30267 = ~w30265 & w30266;
assign w30268 = w30265 & ~w30266;
assign w30269 = ~w30267 & ~w30268;
assign w30270 = ~w30131 & ~w30135;
assign w30271 = ~w28913 & w32322;
assign w30272 = w28912 & w30271;
assign w30273 = ~w30270 & ~w30272;
assign w30274 = (~w30269 & w30272) | (~w30269 & w32323) | (w30272 & w32323);
assign w30275 = w30269 & w30273;
assign w30276 = ~w30274 & ~w30275;
assign w30277 = ~w30141 & ~w30276;
assign w30278 = ~w30139 & ~w30274;
assign w30279 = w29988 & ~w30275;
assign w30280 = w30278 & w30279;
assign w30281 = w29664 & w32324;
assign w30282 = ~w30277 & ~w30281;
assign w30283 = ~w30145 & ~w30263;
assign w30284 = w6061 & w27063;
assign w30285 = w6059 & w27059;
assign w30286 = w6063 & ~w27350;
assign w30287 = ~w30284 & ~w30285;
assign w30288 = ~w30286 & w30287;
assign w30289 = ~a_17 & w30288;
assign w30290 = a_17 & ~w30288;
assign w30291 = ~w30289 & ~w30290;
assign w30292 = ~w30248 & w30259;
assign w30293 = ~w30247 & ~w30292;
assign w30294 = w30291 & ~w30293;
assign w30295 = ~w30291 & w30293;
assign w30296 = ~w30294 & ~w30295;
assign w30297 = ~w30230 & ~w30243;
assign w30298 = ~w30195 & ~w30208;
assign w30299 = ~w30177 & ~w30182;
assign w30300 = ~w30163 & ~w30173;
assign w30301 = ~w195 & w675;
assign w30302 = w1754 & w30301;
assign w30303 = w1740 & w2529;
assign w30304 = w4253 & w14323;
assign w30305 = w30303 & w30304;
assign w30306 = w13987 & w30302;
assign w30307 = w30305 & w30306;
assign w30308 = w2224 & w6641;
assign w30309 = w30307 & w30308;
assign w30310 = w13740 & w30309;
assign w30311 = w3601 & w30310;
assign w30312 = ~w30054 & ~w30311;
assign w30313 = w30054 & w30311;
assign w30314 = ~w30312 & ~w30313;
assign w30315 = ~a_14 & w30314;
assign w30316 = a_14 & ~w30314;
assign w30317 = ~w30315 & ~w30316;
assign w30318 = w30300 & ~w30317;
assign w30319 = ~w30300 & w30317;
assign w30320 = ~w30318 & ~w30319;
assign w30321 = w668 & ~w22020;
assign w30322 = w1327 & w22014;
assign w30323 = w1399 & w22007;
assign w30324 = w1478 & w24122;
assign w30325 = ~w30322 & ~w30323;
assign w30326 = ~w30321 & w30325;
assign w30327 = ~w30324 & w30326;
assign w30328 = w30320 & w30327;
assign w30329 = ~w30320 & ~w30327;
assign w30330 = ~w30328 & ~w30329;
assign w30331 = w3957 & w21771;
assign w30332 = w4068 & w21762;
assign w30333 = w4446 & ~w22035;
assign w30334 = w4070 & w24529;
assign w30335 = ~w30332 & ~w30333;
assign w30336 = ~w30331 & w30335;
assign w30337 = ~w30334 & w30336;
assign w30338 = a_29 & ~w30337;
assign w30339 = ~a_29 & w30337;
assign w30340 = ~w30338 & ~w30339;
assign w30341 = w30330 & ~w30340;
assign w30342 = ~w30330 & w30340;
assign w30343 = ~w30341 & ~w30342;
assign w30344 = w30299 & ~w30343;
assign w30345 = ~w30299 & w30343;
assign w30346 = ~w30344 & ~w30345;
assign w30347 = w4666 & ~w21757;
assign w30348 = ~w518 & w22032;
assign w30349 = w4638 & w22039;
assign w30350 = w1226 & ~w25205;
assign w30351 = ~w30348 & ~w30349;
assign w30352 = ~w30347 & w30351;
assign w30353 = ~w30350 & w30352;
assign w30354 = ~a_26 & w30353;
assign w30355 = a_26 & ~w30353;
assign w30356 = ~w30354 & ~w30355;
assign w30357 = w30346 & w30356;
assign w30358 = ~w30346 & ~w30356;
assign w30359 = ~w30357 & ~w30358;
assign w30360 = w30298 & ~w30359;
assign w30361 = ~w30298 & w30359;
assign w30362 = ~w30360 & ~w30361;
assign w30363 = ~w30222 & ~w30225;
assign w30364 = w5286 & w21746;
assign w30365 = w5016 & w21755;
assign w30366 = w5080 & w21752;
assign w30367 = w5017 & ~w25700;
assign w30368 = ~w30365 & ~w30366;
assign w30369 = ~w30364 & w30368;
assign w30370 = ~w30367 & w30369;
assign w30371 = ~a_23 & w30370;
assign w30372 = a_23 & ~w30370;
assign w30373 = ~w30371 & ~w30372;
assign w30374 = w30363 & ~w30373;
assign w30375 = ~w30363 & w30373;
assign w30376 = ~w30374 & ~w30375;
assign w30377 = ~w30362 & ~w30376;
assign w30378 = w30362 & w30376;
assign w30379 = ~w30377 & ~w30378;
assign w30380 = w5816 & w26766;
assign w30381 = w5308 & ~w21743;
assign w30382 = w5818 & w26476;
assign w30383 = w5309 & ~w26774;
assign w30384 = ~w30381 & ~w30382;
assign w30385 = ~w30380 & w30384;
assign w30386 = ~w30383 & w30385;
assign w30387 = a_20 & w30386;
assign w30388 = ~a_20 & ~w30386;
assign w30389 = ~w30387 & ~w30388;
assign w30390 = w30379 & ~w30389;
assign w30391 = ~w30379 & w30389;
assign w30392 = ~w30390 & ~w30391;
assign w30393 = w30297 & w30392;
assign w30394 = ~w30297 & ~w30392;
assign w30395 = ~w30393 & ~w30394;
assign w30396 = w30296 & ~w30395;
assign w30397 = ~w30296 & w30395;
assign w30398 = ~w30396 & ~w30397;
assign w30399 = ~w30283 & w30398;
assign w30400 = w30283 & ~w30398;
assign w30401 = ~w30399 & ~w30400;
assign w30402 = ~w30268 & ~w30401;
assign w30403 = w30132 & ~w30268;
assign w30404 = ~w30267 & ~w30403;
assign w30405 = w30401 & w30404;
assign w30406 = ~w30131 & ~w30268;
assign w30407 = ~w29974 & w30406;
assign w30408 = ~w29977 & w30407;
assign w30409 = w30405 & ~w30408;
assign w30410 = w29980 & w30405;
assign w30411 = (w30410 & ~w28912) | (w30410 & w32325) | (~w28912 & w32325);
assign w30412 = ~w30409 & ~w30411;
assign w30413 = ~w30402 & w30412;
assign w30414 = w29989 & w30413;
assign w30415 = w30278 & w30414;
assign w30416 = w29664 & w30415;
assign w30417 = ~w30275 & w30402;
assign w30418 = w30412 & ~w30417;
assign w30419 = ~w30281 & ~w30418;
assign w30420 = ~w30416 & ~w30419;
assign w30421 = ~w30294 & ~w30396;
assign w30422 = ~w30375 & ~w30378;
assign w30423 = ~w30342 & ~w30345;
assign w30424 = ~w30312 & ~w30315;
assign w30425 = w77 & ~w156;
assign w30426 = w182 & w1054;
assign w30427 = w1951 & w2361;
assign w30428 = w4732 & w15350;
assign w30429 = w30427 & w30428;
assign w30430 = w30425 & w30426;
assign w30431 = w588 & w2430;
assign w30432 = w25275 & w30431;
assign w30433 = w30429 & w30430;
assign w30434 = w30432 & w30433;
assign w30435 = w5874 & w30434;
assign w30436 = w5386 & w14033;
assign w30437 = w30435 & w30436;
assign w30438 = w2465 & w30437;
assign w30439 = w30424 & ~w30438;
assign w30440 = ~w30424 & w30438;
assign w30441 = ~w30439 & ~w30440;
assign w30442 = w668 & w21771;
assign w30443 = w1399 & w22014;
assign w30444 = w1327 & ~w22020;
assign w30445 = w1478 & w24295;
assign w30446 = ~w30443 & ~w30444;
assign w30447 = ~w30442 & w30446;
assign w30448 = ~w30445 & w30447;
assign w30449 = ~w30441 & ~w30448;
assign w30450 = w30441 & w30448;
assign w30451 = ~w30449 & ~w30450;
assign w30452 = ~w30318 & ~w30328;
assign w30453 = w30451 & ~w30452;
assign w30454 = ~w30451 & w30452;
assign w30455 = ~w30453 & ~w30454;
assign w30456 = w4446 & w22032;
assign w30457 = w3957 & w21762;
assign w30458 = w4068 & ~w22035;
assign w30459 = w4070 & w24756;
assign w30460 = ~w30456 & ~w30457;
assign w30461 = ~w30458 & w30460;
assign w30462 = ~w30459 & w30461;
assign w30463 = a_29 & ~w30462;
assign w30464 = ~a_29 & w30462;
assign w30465 = ~w30463 & ~w30464;
assign w30466 = w30455 & w30465;
assign w30467 = ~w30455 & ~w30465;
assign w30468 = ~w30466 & ~w30467;
assign w30469 = w30423 & ~w30468;
assign w30470 = ~w30423 & w30468;
assign w30471 = ~w30469 & ~w30470;
assign w30472 = w4666 & w21755;
assign w30473 = ~w518 & w22039;
assign w30474 = w4638 & ~w21757;
assign w30475 = w1226 & ~w25675;
assign w30476 = ~w30473 & ~w30474;
assign w30477 = ~w30472 & w30476;
assign w30478 = ~w30475 & w30477;
assign w30479 = a_26 & w30478;
assign w30480 = ~a_26 & ~w30478;
assign w30481 = ~w30479 & ~w30480;
assign w30482 = w30471 & ~w30481;
assign w30483 = ~w30471 & w30481;
assign w30484 = ~w30482 & ~w30483;
assign w30485 = ~w30357 & ~w30361;
assign w30486 = w30484 & ~w30485;
assign w30487 = ~w30484 & w30485;
assign w30488 = ~w30486 & ~w30487;
assign w30489 = w5286 & ~w21743;
assign w30490 = w5016 & w21752;
assign w30491 = w5080 & w21746;
assign w30492 = w5017 & w22065;
assign w30493 = ~w30490 & ~w30491;
assign w30494 = ~w30489 & w30493;
assign w30495 = ~w30492 & w30494;
assign w30496 = a_23 & w30495;
assign w30497 = ~a_23 & ~w30495;
assign w30498 = ~w30496 & ~w30497;
assign w30499 = w30488 & ~w30498;
assign w30500 = ~w30488 & w30498;
assign w30501 = ~w30499 & ~w30500;
assign w30502 = w30422 & ~w30501;
assign w30503 = ~w30422 & w30501;
assign w30504 = ~w30502 & ~w30503;
assign w30505 = w5816 & w27059;
assign w30506 = w5818 & w26766;
assign w30507 = w5308 & w26476;
assign w30508 = w5309 & w27068;
assign w30509 = ~w30506 & ~w30507;
assign w30510 = ~w30505 & w30509;
assign w30511 = ~w30508 & w30510;
assign w30512 = a_20 & ~w30511;
assign w30513 = ~a_20 & w30511;
assign w30514 = ~w30512 & ~w30513;
assign w30515 = w30504 & ~w30514;
assign w30516 = ~w30504 & w30514;
assign w30517 = ~w30515 & ~w30516;
assign w30518 = w6058 & w27063;
assign w30519 = ~a_17 & ~w30518;
assign w30520 = w13488 & w27063;
assign w30521 = ~w30519 & ~w30520;
assign w30522 = ~w30391 & ~w30393;
assign w30523 = w30521 & w30522;
assign w30524 = ~w30521 & ~w30522;
assign w30525 = ~w30523 & ~w30524;
assign w30526 = ~w30517 & w30525;
assign w30527 = w30517 & ~w30525;
assign w30528 = ~w30526 & ~w30527;
assign w30529 = ~w30421 & w30528;
assign w30530 = w30421 & ~w30528;
assign w30531 = ~w30529 & ~w30530;
assign w30532 = w30410 & w30531;
assign w30533 = (w30532 & ~w28912) | (w30532 & w32326) | (~w28912 & w32326);
assign w30534 = ~w30399 & ~w30409;
assign w30535 = w30531 & ~w30534;
assign w30536 = ~w30533 & ~w30535;
assign w30537 = ~w30531 & w30534;
assign w30538 = ~w30411 & w30537;
assign w30539 = w30536 & ~w30538;
assign w30540 = w30278 & w30539;
assign w30541 = w30414 & w30540;
assign w30542 = w29664 & w30541;
assign w30543 = ~w30416 & ~w30539;
assign w30544 = ~w30542 & ~w30543;
assign w30545 = w30405 & ~w30530;
assign w30546 = ~w30408 & w30545;
assign w30547 = ~w30399 & ~w30529;
assign w30548 = ~w30530 & ~w30547;
assign w30549 = ~w30546 & ~w30548;
assign w30550 = w29668 & w30549;
assign w30551 = w28912 & w30550;
assign w30552 = ~w30523 & ~w30526;
assign w30553 = ~w30486 & ~w30499;
assign w30554 = ~w30470 & ~w30482;
assign w30555 = ~w30454 & ~w30466;
assign w30556 = ~w95 & w15259;
assign w30557 = ~w136 & ~w188;
assign w30558 = ~w264 & w30557;
assign w30559 = w1687 & w1815;
assign w30560 = w2274 & w2557;
assign w30561 = w14020 & w30560;
assign w30562 = w30558 & w30559;
assign w30563 = w30042 & w30562;
assign w30564 = w1440 & w30561;
assign w30565 = w2704 & w30556;
assign w30566 = w30564 & w30565;
assign w30567 = w30563 & w30566;
assign w30568 = w1165 & w30567;
assign w30569 = w2118 & w5557;
assign w30570 = w30568 & w30569;
assign w30571 = w30438 & ~w30570;
assign w30572 = ~w30438 & w30570;
assign w30573 = ~w30571 & ~w30572;
assign w30574 = ~w30439 & ~w30450;
assign w30575 = w30573 & w30574;
assign w30576 = ~w30573 & ~w30574;
assign w30577 = ~w30575 & ~w30576;
assign w30578 = w1327 & w21771;
assign w30579 = w668 & w21762;
assign w30580 = w1399 & ~w22020;
assign w30581 = w1478 & w24502;
assign w30582 = ~w30579 & ~w30580;
assign w30583 = ~w30578 & w30582;
assign w30584 = ~w30581 & w30583;
assign w30585 = w30577 & ~w30584;
assign w30586 = ~w30577 & w30584;
assign w30587 = ~w30585 & ~w30586;
assign w30588 = w4446 & w22039;
assign w30589 = w3957 & ~w22035;
assign w30590 = w4068 & w22032;
assign w30591 = w4070 & w24962;
assign w30592 = ~w30589 & ~w30590;
assign w30593 = ~w30588 & w30592;
assign w30594 = ~w30591 & w30593;
assign w30595 = ~a_29 & w30594;
assign w30596 = a_29 & ~w30594;
assign w30597 = ~w30595 & ~w30596;
assign w30598 = w30587 & w30597;
assign w30599 = ~w30587 & ~w30597;
assign w30600 = ~w30598 & ~w30599;
assign w30601 = w30555 & ~w30600;
assign w30602 = ~w30555 & w30600;
assign w30603 = ~w30601 & ~w30602;
assign w30604 = w4666 & w21752;
assign w30605 = ~w518 & ~w21757;
assign w30606 = w4638 & w21755;
assign w30607 = w1226 & w26166;
assign w30608 = ~w30605 & ~w30606;
assign w30609 = ~w30604 & w30608;
assign w30610 = ~w30607 & w30609;
assign w30611 = ~a_26 & w30610;
assign w30612 = a_26 & ~w30610;
assign w30613 = ~w30611 & ~w30612;
assign w30614 = w30603 & w30613;
assign w30615 = ~w30603 & ~w30613;
assign w30616 = ~w30614 & ~w30615;
assign w30617 = w30554 & ~w30616;
assign w30618 = ~w30554 & w30616;
assign w30619 = ~w30617 & ~w30618;
assign w30620 = w5286 & w26476;
assign w30621 = w5080 & ~w21743;
assign w30622 = w5016 & w21746;
assign w30623 = w5017 & w26489;
assign w30624 = ~w30621 & ~w30622;
assign w30625 = ~w30620 & w30624;
assign w30626 = ~w30623 & w30625;
assign w30627 = ~a_23 & w30626;
assign w30628 = a_23 & ~w30626;
assign w30629 = ~w30627 & ~w30628;
assign w30630 = w30619 & w30629;
assign w30631 = ~w30619 & ~w30629;
assign w30632 = ~w30630 & ~w30631;
assign w30633 = w30553 & ~w30632;
assign w30634 = ~w30553 & w30632;
assign w30635 = ~w30633 & ~w30634;
assign w30636 = w5816 & w27063;
assign w30637 = w5818 & w27059;
assign w30638 = w5308 & w26766;
assign w30639 = w5309 & w27094;
assign w30640 = ~w30637 & ~w30638;
assign w30641 = ~w30636 & w30640;
assign w30642 = ~w30639 & w30641;
assign w30643 = a_20 & ~w30642;
assign w30644 = ~a_20 & w30642;
assign w30645 = ~w30643 & ~w30644;
assign w30646 = w30635 & w30645;
assign w30647 = ~w30635 & ~w30645;
assign w30648 = ~w30646 & ~w30647;
assign w30649 = ~w30502 & ~w30515;
assign w30650 = a_17 & w30649;
assign w30651 = ~a_17 & ~w30649;
assign w30652 = ~w30650 & ~w30651;
assign w30653 = w30648 & w30652;
assign w30654 = ~w30648 & ~w30652;
assign w30655 = ~w30653 & ~w30654;
assign w30656 = w30552 & ~w30655;
assign w30657 = ~w30552 & w30655;
assign w30658 = ~w30656 & ~w30657;
assign w30659 = w29978 & w30545;
assign w30660 = w29646 & w30659;
assign w30661 = ~w29642 & w30660;
assign w30662 = w30549 & ~w30661;
assign w30663 = ~w30658 & ~w30662;
assign w30664 = (w30663 & ~w28912) | (w30663 & w32327) | (~w28912 & w32327);
assign w30665 = w30549 & w30658;
assign w30666 = w29667 & w30665;
assign w30667 = ~w28913 & w30666;
assign w30668 = ~w30661 & w30665;
assign w30669 = (~w30668 & ~w28912) | (~w30668 & w32328) | (~w28912 & w32328);
assign w30670 = ~w30664 & w30669;
assign w30671 = w30542 & ~w30670;
assign w30672 = ~w30542 & w30670;
assign w30673 = ~w30671 & ~w30672;
assign w30674 = ~w30618 & ~w30630;
assign w30675 = ~w30585 & ~w30598;
assign w30676 = ~w30572 & ~w30575;
assign w30677 = w2251 & w4544;
assign w30678 = w4712 & w30677;
assign w30679 = w2013 & w2432;
assign w30680 = w6685 & w25277;
assign w30681 = w30679 & w30680;
assign w30682 = w272 & w30678;
assign w30683 = w3681 & w30682;
assign w30684 = w1832 & w30681;
assign w30685 = w30683 & w30684;
assign w30686 = w5184 & w30685;
assign w30687 = w4538 & w30686;
assign w30688 = ~w30570 & ~w30687;
assign w30689 = w30570 & w30687;
assign w30690 = ~w30688 & ~w30689;
assign w30691 = ~a_17 & w30690;
assign w30692 = a_17 & ~w30690;
assign w30693 = ~w30691 & ~w30692;
assign w30694 = w1399 & w21771;
assign w30695 = w1327 & w21762;
assign w30696 = w668 & ~w22035;
assign w30697 = w1478 & w24529;
assign w30698 = ~w30695 & ~w30696;
assign w30699 = ~w30694 & w30698;
assign w30700 = ~w30697 & w30699;
assign w30701 = w30693 & ~w30700;
assign w30702 = ~w30693 & w30700;
assign w30703 = ~w30701 & ~w30702;
assign w30704 = w30676 & ~w30703;
assign w30705 = ~w30676 & w30703;
assign w30706 = ~w30704 & ~w30705;
assign w30707 = w30675 & ~w30706;
assign w30708 = ~w30675 & w30706;
assign w30709 = ~w30707 & ~w30708;
assign w30710 = w4446 & ~w21757;
assign w30711 = w3957 & w22032;
assign w30712 = w4068 & w22039;
assign w30713 = w4070 & ~w25205;
assign w30714 = ~w30711 & ~w30712;
assign w30715 = ~w30710 & w30714;
assign w30716 = ~w30713 & w30715;
assign w30717 = a_29 & w30716;
assign w30718 = ~a_29 & ~w30716;
assign w30719 = ~w30717 & ~w30718;
assign w30720 = w30709 & ~w30719;
assign w30721 = ~w30709 & w30719;
assign w30722 = ~w30720 & ~w30721;
assign w30723 = ~w30602 & ~w30614;
assign w30724 = w4666 & w21746;
assign w30725 = ~w518 & w21755;
assign w30726 = w4638 & w21752;
assign w30727 = w1226 & ~w25700;
assign w30728 = ~w30725 & ~w30726;
assign w30729 = ~w30724 & w30728;
assign w30730 = ~w30727 & w30729;
assign w30731 = ~a_26 & w30730;
assign w30732 = a_26 & ~w30730;
assign w30733 = ~w30731 & ~w30732;
assign w30734 = w30723 & ~w30733;
assign w30735 = ~w30723 & w30733;
assign w30736 = ~w30734 & ~w30735;
assign w30737 = w30722 & w30736;
assign w30738 = ~w30722 & ~w30736;
assign w30739 = ~w30737 & ~w30738;
assign w30740 = w5286 & w26766;
assign w30741 = w5016 & ~w21743;
assign w30742 = w5080 & w26476;
assign w30743 = w5017 & ~w26774;
assign w30744 = ~w30741 & ~w30742;
assign w30745 = ~w30740 & w30744;
assign w30746 = ~w30743 & w30745;
assign w30747 = a_23 & w30746;
assign w30748 = ~a_23 & ~w30746;
assign w30749 = ~w30747 & ~w30748;
assign w30750 = w30739 & ~w30749;
assign w30751 = ~w30739 & w30749;
assign w30752 = ~w30750 & ~w30751;
assign w30753 = w30674 & ~w30752;
assign w30754 = ~w30674 & w30752;
assign w30755 = ~w30753 & ~w30754;
assign w30756 = ~w30634 & ~w30646;
assign w30757 = w5818 & w27063;
assign w30758 = w5308 & w27059;
assign w30759 = w5309 & ~w27350;
assign w30760 = ~w30757 & ~w30758;
assign w30761 = ~w30759 & w30760;
assign w30762 = ~a_20 & w30761;
assign w30763 = a_20 & ~w30761;
assign w30764 = ~w30762 & ~w30763;
assign w30765 = w30756 & ~w30764;
assign w30766 = ~w30756 & w30764;
assign w30767 = ~w30765 & ~w30766;
assign w30768 = ~w30755 & ~w30767;
assign w30769 = w30755 & w30767;
assign w30770 = ~w30768 & ~w30769;
assign w30771 = ~w30650 & ~w30653;
assign w30772 = w30770 & ~w30771;
assign w30773 = ~w30770 & w30771;
assign w30774 = ~w30772 & ~w30773;
assign w30775 = w30668 & w30774;
assign w30776 = ~w28913 & w32329;
assign w30777 = ~w30656 & w30774;
assign w30778 = w30656 & ~w30774;
assign w30779 = ~w30777 & ~w30778;
assign w30780 = ~w30668 & w30779;
assign w30781 = (w30780 & ~w28912) | (w30780 & w32330) | (~w28912 & w32330);
assign w30782 = (~w30775 & ~w28912) | (~w30775 & w32631) | (~w28912 & w32631);
assign w30783 = ~w30781 & w30782;
assign w30784 = (w30783 & ~w30542) | (w30783 & w32331) | (~w30542 & w32331);
assign w30785 = ~w30670 & ~w30783;
assign w30786 = w30542 & w30785;
assign w30787 = ~w30784 & ~w30786;
assign w30788 = ~w30766 & ~w30769;
assign w30789 = ~w30735 & ~w30737;
assign w30790 = ~w30708 & ~w30720;
assign w30791 = ~w30688 & ~w30691;
assign w30792 = ~w623 & ~w732;
assign w30793 = w594 & w30792;
assign w30794 = w1152 & w1929;
assign w30795 = w2440 & w4714;
assign w30796 = w26583 & w30795;
assign w30797 = w30793 & w30794;
assign w30798 = w2644 & w13030;
assign w30799 = w30797 & w30798;
assign w30800 = w30796 & w30799;
assign w30801 = w2534 & w3777;
assign w30802 = w30800 & w30801;
assign w30803 = w6524 & w30802;
assign w30804 = w29211 & w30803;
assign w30805 = w30791 & ~w30804;
assign w30806 = ~w30791 & w30804;
assign w30807 = ~w30805 & ~w30806;
assign w30808 = w668 & w22032;
assign w30809 = w1399 & w21762;
assign w30810 = w1327 & ~w22035;
assign w30811 = w1478 & w24756;
assign w30812 = ~w30808 & ~w30809;
assign w30813 = ~w30810 & w30812;
assign w30814 = ~w30811 & w30813;
assign w30815 = ~w30807 & ~w30814;
assign w30816 = w30807 & w30814;
assign w30817 = ~w30815 & ~w30816;
assign w30818 = ~w30701 & ~w30705;
assign w30819 = ~w30817 & ~w30818;
assign w30820 = w30817 & w30818;
assign w30821 = ~w30819 & ~w30820;
assign w30822 = w4446 & w21755;
assign w30823 = w4068 & ~w21757;
assign w30824 = w3957 & w22039;
assign w30825 = w4070 & ~w25675;
assign w30826 = ~w30823 & ~w30824;
assign w30827 = ~w30822 & w30826;
assign w30828 = ~w30825 & w30827;
assign w30829 = ~a_29 & w30828;
assign w30830 = a_29 & ~w30828;
assign w30831 = ~w30829 & ~w30830;
assign w30832 = w30821 & w30831;
assign w30833 = ~w30821 & ~w30831;
assign w30834 = ~w30832 & ~w30833;
assign w30835 = w30790 & ~w30834;
assign w30836 = ~w30790 & w30834;
assign w30837 = ~w30835 & ~w30836;
assign w30838 = w4666 & ~w21743;
assign w30839 = ~w518 & w21752;
assign w30840 = w4638 & w21746;
assign w30841 = w1226 & w22065;
assign w30842 = ~w30839 & ~w30840;
assign w30843 = ~w30838 & w30842;
assign w30844 = ~w30841 & w30843;
assign w30845 = a_26 & w30844;
assign w30846 = ~a_26 & ~w30844;
assign w30847 = ~w30845 & ~w30846;
assign w30848 = w30837 & ~w30847;
assign w30849 = ~w30837 & w30847;
assign w30850 = ~w30848 & ~w30849;
assign w30851 = w30789 & ~w30850;
assign w30852 = ~w30789 & w30850;
assign w30853 = ~w30851 & ~w30852;
assign w30854 = w5286 & w27059;
assign w30855 = w5016 & w26476;
assign w30856 = w5080 & w26766;
assign w30857 = w5017 & w27068;
assign w30858 = ~w30855 & ~w30856;
assign w30859 = ~w30854 & w30858;
assign w30860 = ~w30857 & w30859;
assign w30861 = a_23 & w30860;
assign w30862 = ~a_23 & ~w30860;
assign w30863 = ~w30861 & ~w30862;
assign w30864 = w30853 & ~w30863;
assign w30865 = ~w30853 & w30863;
assign w30866 = ~w30864 & ~w30865;
assign w30867 = ~w30750 & ~w30754;
assign w30868 = w30866 & ~w30867;
assign w30869 = ~w30866 & w30867;
assign w30870 = ~w30868 & ~w30869;
assign w30871 = w5304 & w27063;
assign w30872 = ~a_20 & ~w30871;
assign w30873 = w13110 & w27063;
assign w30874 = ~w30872 & ~w30873;
assign w30875 = w30870 & w30874;
assign w30876 = ~w30870 & ~w30874;
assign w30877 = ~w30875 & ~w30876;
assign w30878 = w30788 & ~w30877;
assign w30879 = ~w30788 & w30877;
assign w30880 = ~w30878 & ~w30879;
assign w30881 = w30772 & w30880;
assign w30882 = ~w30772 & ~w30880;
assign w30883 = ~w30881 & ~w30882;
assign w30884 = w30410 & w30883;
assign w30885 = (w30884 & ~w28912) | (w30884 & w32332) | (~w28912 & w32332);
assign w30886 = ~w30537 & w30883;
assign w30887 = ~w30885 & ~w30886;
assign w30888 = w30536 & ~w30887;
assign w30889 = w30785 & w30888;
assign w30890 = w29664 & w32333;
assign w30891 = ~w30551 & ~w30662;
assign w30892 = ~w30657 & ~w30891;
assign w30893 = w30777 & ~w30892;
assign w30894 = w30883 & ~w30893;
assign w30895 = ~w30880 & w30893;
assign w30896 = ~w30894 & ~w30895;
assign w30897 = (w30896 & ~w30542) | (w30896 & w32334) | (~w30542 & w32334);
assign w30898 = ~w30890 & ~w30897;
assign w30899 = ~w30772 & ~w30879;
assign w30900 = ~w30657 & w30899;
assign w30901 = w30549 & w30900;
assign w30902 = w29667 & w30901;
assign w30903 = ~w28913 & w30902;
assign w30904 = w28912 & w30903;
assign w30905 = ~w30661 & w30901;
assign w30906 = ~w30836 & ~w30848;
assign w30907 = ~w30819 & ~w30832;
assign w30908 = ~w313 & ~w540;
assign w30909 = ~w694 & w30908;
assign w30910 = w209 & w1641;
assign w30911 = w2873 & w3426;
assign w30912 = w3434 & w30911;
assign w30913 = w30909 & w30910;
assign w30914 = w30912 & w30913;
assign w30915 = w30556 & w30914;
assign w30916 = w4520 & w28379;
assign w30917 = w30915 & w30916;
assign w30918 = w4933 & w30917;
assign w30919 = w1847 & w6753;
assign w30920 = w30918 & w30919;
assign w30921 = w30804 & ~w30920;
assign w30922 = ~w30804 & w30920;
assign w30923 = ~w30921 & ~w30922;
assign w30924 = w668 & w22039;
assign w30925 = w1399 & ~w22035;
assign w30926 = w1327 & w22032;
assign w30927 = w1478 & w24962;
assign w30928 = ~w30925 & ~w30926;
assign w30929 = ~w30924 & w30928;
assign w30930 = ~w30927 & w30929;
assign w30931 = w30923 & ~w30930;
assign w30932 = ~w30923 & w30930;
assign w30933 = ~w30931 & ~w30932;
assign w30934 = ~w30805 & ~w30816;
assign w30935 = w30933 & w30934;
assign w30936 = ~w30933 & ~w30934;
assign w30937 = ~w30935 & ~w30936;
assign w30938 = w30907 & ~w30937;
assign w30939 = ~w30907 & w30937;
assign w30940 = ~w30938 & ~w30939;
assign w30941 = w4446 & w21752;
assign w30942 = w3957 & ~w21757;
assign w30943 = w4068 & w21755;
assign w30944 = w4070 & w26166;
assign w30945 = ~w30942 & ~w30943;
assign w30946 = ~w30941 & w30945;
assign w30947 = ~w30944 & w30946;
assign w30948 = ~a_29 & w30947;
assign w30949 = a_29 & ~w30947;
assign w30950 = ~w30948 & ~w30949;
assign w30951 = w30940 & w30950;
assign w30952 = ~w30940 & ~w30950;
assign w30953 = ~w30951 & ~w30952;
assign w30954 = w4666 & w26476;
assign w30955 = ~w518 & w21746;
assign w30956 = w4638 & ~w21743;
assign w30957 = w1226 & w26489;
assign w30958 = ~w30955 & ~w30956;
assign w30959 = ~w30954 & w30958;
assign w30960 = ~w30957 & w30959;
assign w30961 = a_26 & w30960;
assign w30962 = ~a_26 & ~w30960;
assign w30963 = ~w30961 & ~w30962;
assign w30964 = w30953 & ~w30963;
assign w30965 = ~w30953 & w30963;
assign w30966 = ~w30964 & ~w30965;
assign w30967 = w30906 & ~w30966;
assign w30968 = ~w30906 & w30966;
assign w30969 = ~w30967 & ~w30968;
assign w30970 = w5286 & w27063;
assign w30971 = w5080 & w27059;
assign w30972 = w5016 & w26766;
assign w30973 = w5017 & w27094;
assign w30974 = ~w30971 & ~w30972;
assign w30975 = ~w30970 & w30974;
assign w30976 = ~w30973 & w30975;
assign w30977 = a_23 & ~w30976;
assign w30978 = ~a_23 & w30976;
assign w30979 = ~w30977 & ~w30978;
assign w30980 = w30969 & w30979;
assign w30981 = ~w30969 & ~w30979;
assign w30982 = ~w30980 & ~w30981;
assign w30983 = ~w30852 & ~w30864;
assign w30984 = a_20 & ~w30983;
assign w30985 = ~a_20 & w30983;
assign w30986 = ~w30984 & ~w30985;
assign w30987 = w30982 & w30986;
assign w30988 = ~w30982 & ~w30986;
assign w30989 = ~w30987 & ~w30988;
assign w30990 = ~w30868 & ~w30875;
assign w30991 = ~w30989 & w30990;
assign w30992 = w30989 & ~w30990;
assign w30993 = ~w30991 & ~w30992;
assign w30994 = ~w30777 & w30899;
assign w30995 = ~w30878 & ~w30994;
assign w30996 = w30993 & w30995;
assign w30997 = ~w30905 & w30996;
assign w30998 = (w30997 & ~w28912) | (w30997 & w32335) | (~w28912 & w32335);
assign w30999 = ~w30905 & w30995;
assign w31000 = ~w30993 & ~w30999;
assign w31001 = ~w28913 & w32336;
assign w31002 = w28912 & w31001;
assign w31003 = ~w31000 & ~w31002;
assign w31004 = ~w30998 & w31003;
assign w31005 = w30890 & ~w31004;
assign w31006 = ~w30890 & w31004;
assign w31007 = ~w31005 & ~w31006;
assign w31008 = ~w30984 & ~w30987;
assign w31009 = ~w30951 & ~w30964;
assign w31010 = ~w30921 & ~w30931;
assign w31011 = ~w281 & ~w400;
assign w31012 = w839 & w31011;
assign w31013 = w1007 & w1562;
assign w31014 = w1948 & w2078;
assign w31015 = w5613 & w31014;
assign w31016 = w31012 & w31013;
assign w31017 = w1108 & w1497;
assign w31018 = w1865 & w31017;
assign w31019 = w31015 & w31016;
assign w31020 = w2704 & w14353;
assign w31021 = w31019 & w31020;
assign w31022 = w15247 & w31018;
assign w31023 = w31021 & w31022;
assign w31024 = w2176 & w31023;
assign w31025 = w236 & w31024;
assign w31026 = ~w30804 & ~w31025;
assign w31027 = w30804 & w31025;
assign w31028 = ~w31026 & ~w31027;
assign w31029 = ~a_20 & w31028;
assign w31030 = a_20 & ~w31028;
assign w31031 = ~w31029 & ~w31030;
assign w31032 = w31010 & ~w31031;
assign w31033 = ~w31010 & w31031;
assign w31034 = ~w31032 & ~w31033;
assign w31035 = w668 & ~w21757;
assign w31036 = w1327 & w22039;
assign w31037 = w1399 & w22032;
assign w31038 = w1478 & ~w25205;
assign w31039 = ~w31036 & ~w31037;
assign w31040 = ~w31035 & w31039;
assign w31041 = ~w31038 & w31040;
assign w31042 = w31034 & w31041;
assign w31043 = ~w31034 & ~w31041;
assign w31044 = ~w31042 & ~w31043;
assign w31045 = ~w30935 & ~w30939;
assign w31046 = ~w31044 & ~w31045;
assign w31047 = w31044 & w31045;
assign w31048 = ~w31046 & ~w31047;
assign w31049 = w4446 & w21746;
assign w31050 = w4068 & w21752;
assign w31051 = w3957 & w21755;
assign w31052 = w4070 & ~w25700;
assign w31053 = ~w31050 & ~w31051;
assign w31054 = ~w31049 & w31053;
assign w31055 = ~w31052 & w31054;
assign w31056 = ~a_29 & w31055;
assign w31057 = a_29 & ~w31055;
assign w31058 = ~w31056 & ~w31057;
assign w31059 = w31048 & w31058;
assign w31060 = ~w31048 & ~w31058;
assign w31061 = ~w31059 & ~w31060;
assign w31062 = w4666 & w26766;
assign w31063 = w4638 & w26476;
assign w31064 = ~w518 & ~w21743;
assign w31065 = w1226 & ~w26774;
assign w31066 = ~w31063 & ~w31064;
assign w31067 = ~w31062 & w31066;
assign w31068 = ~w31065 & w31067;
assign w31069 = a_26 & ~w31068;
assign w31070 = ~a_26 & w31068;
assign w31071 = ~w31069 & ~w31070;
assign w31072 = w31061 & w31071;
assign w31073 = ~w31061 & ~w31071;
assign w31074 = ~w31072 & ~w31073;
assign w31075 = w31009 & ~w31074;
assign w31076 = ~w31009 & w31074;
assign w31077 = ~w31075 & ~w31076;
assign w31078 = ~w30968 & ~w30980;
assign w31079 = w5080 & w27063;
assign w31080 = w5016 & w27059;
assign w31081 = w5017 & ~w27350;
assign w31082 = ~w31079 & ~w31080;
assign w31083 = ~w31081 & w31082;
assign w31084 = ~a_23 & w31083;
assign w31085 = a_23 & ~w31083;
assign w31086 = ~w31084 & ~w31085;
assign w31087 = w31078 & ~w31086;
assign w31088 = ~w31078 & w31086;
assign w31089 = ~w31087 & ~w31088;
assign w31090 = ~w31077 & ~w31089;
assign w31091 = w31077 & w31089;
assign w31092 = ~w31090 & ~w31091;
assign w31093 = w31008 & ~w31092;
assign w31094 = ~w31008 & w31092;
assign w31095 = ~w31093 & ~w31094;
assign w31096 = w30992 & w31095;
assign w31097 = ~w30991 & w31095;
assign w31098 = w30995 & w31097;
assign w31099 = ~w30905 & w31098;
assign w31100 = ~w31096 & ~w31099;
assign w31101 = ~w28913 & w32337;
assign w31102 = w28912 & w31101;
assign w31103 = ~w31100 & ~w31102;
assign w31104 = ~w30992 & ~w31095;
assign w31105 = ~w28913 & w32338;
assign w31106 = w28912 & w31105;
assign w31107 = ~w30997 & w31104;
assign w31108 = ~w31106 & ~w31107;
assign w31109 = ~w31103 & w31108;
assign w31110 = ~w30890 & w31109;
assign w31111 = w31004 & w31109;
assign w31112 = ~w31004 & ~w31109;
assign w31113 = ~w31111 & ~w31112;
assign w31114 = w30890 & w31113;
assign w31115 = ~w31110 & ~w31114;
assign w31116 = ~w31088 & ~w31091;
assign w31117 = w508 & w27063;
assign w31118 = ~a_23 & ~w31117;
assign w31119 = w510 & w27063;
assign w31120 = ~w31118 & ~w31119;
assign w31121 = ~w31046 & ~w31059;
assign w31122 = ~w31026 & ~w31029;
assign w31123 = ~w393 & ~w463;
assign w31124 = w911 & w31123;
assign w31125 = w3369 & w3495;
assign w31126 = w5185 & w15222;
assign w31127 = w31125 & w31126;
assign w31128 = w2190 & w31124;
assign w31129 = w4084 & w31128;
assign w31130 = w3523 & w31127;
assign w31131 = w31129 & w31130;
assign w31132 = w4261 & w15354;
assign w31133 = w31131 & w31132;
assign w31134 = w377 & w3341;
assign w31135 = w31133 & w31134;
assign w31136 = w4537 & w31135;
assign w31137 = w31122 & ~w31136;
assign w31138 = ~w31122 & w31136;
assign w31139 = ~w31137 & ~w31138;
assign w31140 = w668 & w21755;
assign w31141 = w1327 & ~w21757;
assign w31142 = w1399 & w22039;
assign w31143 = w1478 & ~w25675;
assign w31144 = ~w31141 & ~w31142;
assign w31145 = ~w31140 & w31144;
assign w31146 = ~w31143 & w31145;
assign w31147 = ~w31139 & ~w31146;
assign w31148 = w31139 & w31146;
assign w31149 = ~w31147 & ~w31148;
assign w31150 = ~w31032 & ~w31042;
assign w31151 = w31149 & ~w31150;
assign w31152 = ~w31149 & w31150;
assign w31153 = ~w31151 & ~w31152;
assign w31154 = w4446 & ~w21743;
assign w31155 = w4068 & w21746;
assign w31156 = w3957 & w21752;
assign w31157 = w4070 & w22065;
assign w31158 = ~w31155 & ~w31156;
assign w31159 = ~w31154 & w31158;
assign w31160 = ~w31157 & w31159;
assign w31161 = ~a_29 & w31160;
assign w31162 = a_29 & ~w31160;
assign w31163 = ~w31161 & ~w31162;
assign w31164 = w31153 & w31163;
assign w31165 = ~w31153 & ~w31163;
assign w31166 = ~w31164 & ~w31165;
assign w31167 = w31121 & ~w31166;
assign w31168 = ~w31121 & w31166;
assign w31169 = ~w31167 & ~w31168;
assign w31170 = w4666 & w27059;
assign w31171 = ~w518 & w26476;
assign w31172 = w4638 & w26766;
assign w31173 = w1226 & w27068;
assign w31174 = ~w31171 & ~w31172;
assign w31175 = ~w31170 & w31174;
assign w31176 = ~w31173 & w31175;
assign w31177 = a_26 & ~w31176;
assign w31178 = ~a_26 & w31176;
assign w31179 = ~w31177 & ~w31178;
assign w31180 = w31169 & ~w31179;
assign w31181 = ~w31169 & w31179;
assign w31182 = ~w31180 & ~w31181;
assign w31183 = ~w31072 & ~w31076;
assign w31184 = ~w31182 & ~w31183;
assign w31185 = w31182 & w31183;
assign w31186 = ~w31184 & ~w31185;
assign w31187 = w31120 & w31186;
assign w31188 = ~w31120 & ~w31186;
assign w31189 = ~w31187 & ~w31188;
assign w31190 = w31116 & ~w31189;
assign w31191 = ~w31116 & w31189;
assign w31192 = ~w31190 & ~w31191;
assign w31193 = ~w31094 & ~w31096;
assign w31194 = ~w31192 & ~w31193;
assign w31195 = w31192 & w31193;
assign w31196 = ~w28913 & w32339;
assign w31197 = w28912 & w31196;
assign w31198 = ~w31099 & w31195;
assign w31199 = w31099 & ~w31192;
assign w31200 = ~w30904 & w31199;
assign w31201 = ~w31197 & w32340;
assign w31202 = ~w31200 & w31201;
assign w31203 = w31111 & ~w31202;
assign w31204 = w30889 & w31203;
assign w31205 = w30416 & w31204;
assign w31206 = w30889 & w31111;
assign w31207 = (w31202 & ~w30416) | (w31202 & w32341) | (~w30416 & w32341);
assign w31208 = ~w31205 & ~w31207;
assign w31209 = ~w31184 & ~w31187;
assign w31210 = ~w31152 & ~w31164;
assign w31211 = ~w56 & ~w62;
assign w31212 = ~w907 & w31211;
assign w31213 = w911 & w1109;
assign w31214 = w1572 & w1665;
assign w31215 = w2100 & w31214;
assign w31216 = w31212 & w31213;
assign w31217 = w1386 & w13032;
assign w31218 = w15163 & w31217;
assign w31219 = w31215 & w31216;
assign w31220 = w31218 & w31219;
assign w31221 = w556 & w29216;
assign w31222 = w31220 & w31221;
assign w31223 = w24817 & w31222;
assign w31224 = w772 & w31223;
assign w31225 = w31136 & ~w31224;
assign w31226 = ~w31136 & w31224;
assign w31227 = ~w31225 & ~w31226;
assign w31228 = ~w31137 & ~w31148;
assign w31229 = w31227 & w31228;
assign w31230 = ~w31227 & ~w31228;
assign w31231 = ~w31229 & ~w31230;
assign w31232 = w668 & w21752;
assign w31233 = w1399 & ~w21757;
assign w31234 = w1327 & w21755;
assign w31235 = w1478 & w26166;
assign w31236 = ~w31233 & ~w31234;
assign w31237 = ~w31232 & w31236;
assign w31238 = ~w31235 & w31237;
assign w31239 = w31231 & ~w31238;
assign w31240 = ~w31231 & w31238;
assign w31241 = ~w31239 & ~w31240;
assign w31242 = w31210 & ~w31241;
assign w31243 = ~w31210 & w31241;
assign w31244 = ~w31242 & ~w31243;
assign w31245 = w4446 & w26476;
assign w31246 = w4068 & ~w21743;
assign w31247 = w3957 & w21746;
assign w31248 = w4070 & w26489;
assign w31249 = ~w31246 & ~w31247;
assign w31250 = ~w31245 & w31249;
assign w31251 = ~w31248 & w31250;
assign w31252 = a_29 & ~w31251;
assign w31253 = ~a_29 & w31251;
assign w31254 = ~w31252 & ~w31253;
assign w31255 = w31244 & w31254;
assign w31256 = ~w31244 & ~w31254;
assign w31257 = ~w31255 & ~w31256;
assign w31258 = w4666 & w27063;
assign w31259 = ~w518 & w26766;
assign w31260 = w4638 & w27059;
assign w31261 = w1226 & w27094;
assign w31262 = ~w31259 & ~w31260;
assign w31263 = ~w31258 & w31262;
assign w31264 = ~w31261 & w31263;
assign w31265 = ~a_26 & w31264;
assign w31266 = a_26 & ~w31264;
assign w31267 = ~w31265 & ~w31266;
assign w31268 = w31257 & w31267;
assign w31269 = ~w31257 & ~w31267;
assign w31270 = ~w31268 & ~w31269;
assign w31271 = ~w31167 & ~w31180;
assign w31272 = a_23 & w31271;
assign w31273 = ~a_23 & ~w31271;
assign w31274 = ~w31272 & ~w31273;
assign w31275 = w31270 & w31274;
assign w31276 = ~w31270 & ~w31274;
assign w31277 = ~w31275 & ~w31276;
assign w31278 = w31209 & ~w31277;
assign w31279 = ~w31209 & w31277;
assign w31280 = ~w31278 & ~w31279;
assign w31281 = ~w31190 & w31280;
assign w31282 = w31190 & ~w31280;
assign w31283 = ~w31281 & ~w31282;
assign w31284 = ~w31197 & w32342;
assign w31285 = (~w31280 & w31197) | (~w31280 & w32343) | (w31197 & w32343);
assign w31286 = ~w31284 & ~w31285;
assign w31287 = (w31286 & ~w30416) | (w31286 & w32344) | (~w30416 & w32344);
assign w31288 = w30416 & w32345;
assign w31289 = ~w31287 & ~w31288;
assign w31290 = ~w31272 & ~w31275;
assign w31291 = ~w31239 & ~w31243;
assign w31292 = ~w31226 & ~w31229;
assign w31293 = w1249 & w5371;
assign w31294 = w674 & w31293;
assign w31295 = w1465 & w2135;
assign w31296 = w3868 & w31295;
assign w31297 = w521 & w31294;
assign w31298 = w31296 & w31297;
assign w31299 = w1300 & w31298;
assign w31300 = w3899 & w31299;
assign w31301 = w3849 & w31300;
assign w31302 = ~w31224 & ~w31301;
assign w31303 = w31224 & w31301;
assign w31304 = ~w31302 & ~w31303;
assign w31305 = ~a_23 & w31304;
assign w31306 = a_23 & ~w31304;
assign w31307 = ~w31305 & ~w31306;
assign w31308 = w31292 & ~w31307;
assign w31309 = ~w31292 & w31307;
assign w31310 = ~w31308 & ~w31309;
assign w31311 = w668 & w21746;
assign w31312 = w1327 & w21752;
assign w31313 = w1399 & w21755;
assign w31314 = w1478 & ~w25700;
assign w31315 = ~w31312 & ~w31313;
assign w31316 = ~w31311 & w31315;
assign w31317 = ~w31314 & w31316;
assign w31318 = w31310 & ~w31317;
assign w31319 = ~w31310 & w31317;
assign w31320 = ~w31318 & ~w31319;
assign w31321 = w31291 & ~w31320;
assign w31322 = ~w31291 & w31320;
assign w31323 = ~w31321 & ~w31322;
assign w31324 = w4446 & w26766;
assign w31325 = w3957 & ~w21743;
assign w31326 = w4068 & w26476;
assign w31327 = w4070 & ~w26774;
assign w31328 = ~w31325 & ~w31326;
assign w31329 = ~w31324 & w31328;
assign w31330 = ~w31327 & w31329;
assign w31331 = a_29 & w31330;
assign w31332 = ~a_29 & ~w31330;
assign w31333 = ~w31331 & ~w31332;
assign w31334 = w31323 & ~w31333;
assign w31335 = ~w31323 & w31333;
assign w31336 = ~w31334 & ~w31335;
assign w31337 = ~w31255 & ~w31268;
assign w31338 = w4638 & w27063;
assign w31339 = ~w518 & w27059;
assign w31340 = w1226 & ~w27350;
assign w31341 = ~w31338 & ~w31339;
assign w31342 = ~w31340 & w31341;
assign w31343 = ~a_26 & w31342;
assign w31344 = a_26 & ~w31342;
assign w31345 = ~w31343 & ~w31344;
assign w31346 = w31337 & ~w31345;
assign w31347 = ~w31337 & w31345;
assign w31348 = ~w31346 & ~w31347;
assign w31349 = w31336 & w31348;
assign w31350 = ~w31336 & ~w31348;
assign w31351 = ~w31349 & ~w31350;
assign w31352 = ~w31290 & w31351;
assign w31353 = w31290 & ~w31351;
assign w31354 = ~w31352 & ~w31353;
assign w31355 = ~w31279 & ~w31281;
assign w31356 = w31354 & ~w31355;
assign w31357 = w31099 & w31356;
assign w31358 = ~w31195 & w31281;
assign w31359 = ~w31279 & ~w31358;
assign w31360 = w31354 & ~w31359;
assign w31361 = (~w31360 & w30904) | (~w31360 & w32346) | (w30904 & w32346);
assign w31362 = ~w31354 & w31355;
assign w31363 = w31099 & ~w31362;
assign w31364 = ~w31354 & w31359;
assign w31365 = (w31364 & w30904) | (w31364 & w32347) | (w30904 & w32347);
assign w31366 = w31361 & ~w31365;
assign w31367 = (w31366 & ~w30416) | (w31366 & w32348) | (~w30416 & w32348);
assign w31368 = w31286 & w31366;
assign w31369 = ~w31286 & ~w31366;
assign w31370 = ~w31368 & ~w31369;
assign w31371 = w30416 & w32349;
assign w31372 = ~w31367 & ~w31371;
assign w31373 = ~w31347 & ~w31349;
assign w31374 = ~w31322 & ~w31334;
assign w31375 = ~w31302 & ~w31305;
assign w31376 = ~w190 & ~w389;
assign w31377 = w386 & w31376;
assign w31378 = w1487 & w2400;
assign w31379 = w4385 & w15414;
assign w31380 = w31378 & w31379;
assign w31381 = w29374 & w31377;
assign w31382 = w31380 & w31381;
assign w31383 = w1264 & w6695;
assign w31384 = w14324 & w31383;
assign w31385 = w1286 & w31382;
assign w31386 = w1383 & w31385;
assign w31387 = w31384 & w31386;
assign w31388 = w15183 & w31387;
assign w31389 = w13219 & w31388;
assign w31390 = w31375 & ~w31389;
assign w31391 = ~w31375 & w31389;
assign w31392 = ~w31390 & ~w31391;
assign w31393 = w668 & ~w21743;
assign w31394 = w1327 & w21746;
assign w31395 = w1399 & w21752;
assign w31396 = w1478 & w22065;
assign w31397 = ~w31394 & ~w31395;
assign w31398 = ~w31393 & w31397;
assign w31399 = ~w31396 & w31398;
assign w31400 = ~w31392 & ~w31399;
assign w31401 = w31392 & w31399;
assign w31402 = ~w31400 & ~w31401;
assign w31403 = ~w31309 & ~w31318;
assign w31404 = ~w31402 & ~w31403;
assign w31405 = w31402 & w31403;
assign w31406 = ~w31404 & ~w31405;
assign w31407 = w4446 & w27059;
assign w31408 = w4068 & w26766;
assign w31409 = w3957 & w26476;
assign w31410 = w4070 & w27068;
assign w31411 = ~w31408 & ~w31409;
assign w31412 = ~w31407 & w31411;
assign w31413 = ~w31410 & w31412;
assign w31414 = a_29 & ~w31413;
assign w31415 = ~a_29 & w31413;
assign w31416 = ~w31414 & ~w31415;
assign w31417 = w31406 & w31416;
assign w31418 = ~w31406 & ~w31416;
assign w31419 = ~w31417 & ~w31418;
assign w31420 = w31374 & ~w31419;
assign w31421 = ~w31374 & w31419;
assign w31422 = ~w31420 & ~w31421;
assign w31423 = ~w518 & w27063;
assign w31424 = a_26 & ~w31423;
assign w31425 = ~a_26 & w31423;
assign w31426 = ~w31424 & ~w31425;
assign w31427 = w31422 & ~w31426;
assign w31428 = ~w31422 & w31426;
assign w31429 = ~w31427 & ~w31428;
assign w31430 = w31373 & ~w31429;
assign w31431 = ~w31373 & w31429;
assign w31432 = ~w31430 & ~w31431;
assign w31433 = w31352 & ~w31432;
assign w31434 = ~w31352 & ~w31431;
assign w31435 = ~w31430 & w31434;
assign w31436 = ~w31433 & ~w31435;
assign w31437 = w31368 & ~w31436;
assign w31438 = w31204 & w31437;
assign w31439 = w30416 & w31438;
assign w31440 = w31203 & w32632;
assign w31441 = w31361 & ~w31436;
assign w31442 = ~w31361 & w31436;
assign w31443 = ~w31441 & ~w31442;
assign w31444 = (w31443 & ~w30416) | (w31443 & w32633) | (~w30416 & w32633);
assign w31445 = ~w31439 & ~w31444;
assign w31446 = ~w31356 & w31435;
assign w31447 = w31099 & ~w31446;
assign w31448 = ~w31360 & w31435;
assign w31449 = (w31448 & w30904) | (w31448 & w32350) | (w30904 & w32350);
assign w31450 = ~w31421 & ~w31427;
assign w31451 = ~w31404 & ~w31417;
assign w31452 = ~w31390 & ~w31401;
assign w31453 = w1335 & w1591;
assign w31454 = w2984 & w31453;
assign w31455 = w1259 & w1278;
assign w31456 = w3876 & w12983;
assign w31457 = w31455 & w31456;
assign w31458 = w31454 & w31457;
assign w31459 = ~w31388 & w31458;
assign w31460 = w31389 & ~w31458;
assign w31461 = ~w31459 & ~w31460;
assign w31462 = ~w31452 & w31461;
assign w31463 = w31452 & ~w31461;
assign w31464 = ~w31462 & ~w31463;
assign w31465 = w668 & w26476;
assign w31466 = w1327 & ~w21743;
assign w31467 = w1399 & w21746;
assign w31468 = w1478 & w26489;
assign w31469 = ~w31466 & ~w31467;
assign w31470 = ~w31465 & w31469;
assign w31471 = ~w31468 & w31470;
assign w31472 = ~w31464 & ~w31471;
assign w31473 = w31464 & w31471;
assign w31474 = ~w31472 & ~w31473;
assign w31475 = w31451 & ~w31474;
assign w31476 = ~w31451 & w31474;
assign w31477 = ~w31475 & ~w31476;
assign w31478 = w4446 & w27063;
assign w31479 = w4068 & w27059;
assign w31480 = w3957 & w26766;
assign w31481 = w4070 & w27094;
assign w31482 = ~w31479 & ~w31480;
assign w31483 = ~w31478 & w31482;
assign w31484 = ~w31481 & w31483;
assign w31485 = a_29 & ~w31484;
assign w31486 = ~a_29 & w31484;
assign w31487 = ~w31485 & ~w31486;
assign w31488 = a_26 & w31487;
assign w31489 = ~a_26 & ~w31487;
assign w31490 = ~w31488 & ~w31489;
assign w31491 = ~w31477 & ~w31490;
assign w31492 = w31477 & w31490;
assign w31493 = ~w31491 & ~w31492;
assign w31494 = w31450 & ~w31493;
assign w31495 = ~w31450 & w31493;
assign w31496 = ~w31494 & ~w31495;
assign w31497 = ~w31436 & w31496;
assign w31498 = w31449 & w31497;
assign w31499 = ~w31430 & w31496;
assign w31500 = w31430 & ~w31496;
assign w31501 = ~w31499 & ~w31500;
assign w31502 = ~w31436 & w31501;
assign w31503 = ~w31449 & w31502;
assign w31504 = ~w31498 & ~w31503;
assign w31505 = w31368 & ~w31504;
assign w31506 = w31204 & w31505;
assign w31507 = w30416 & w31506;
assign w31508 = w31449 & ~w31496;
assign w31509 = ~w31449 & ~w31501;
assign w31510 = ~w31508 & ~w31509;
assign w31511 = ~w31439 & ~w31510;
assign w31512 = ~w31507 & ~w31511;
assign w31513 = w31361 & w31434;
assign w31514 = w31499 & ~w31513;
assign w31515 = ~w31495 & ~w31514;
assign w31516 = ~w31488 & ~w31492;
assign w31517 = w3957 & w27059;
assign w31518 = w4070 & ~w27350;
assign w31519 = ~w31517 & ~w31518;
assign w31520 = w668 & w26766;
assign w31521 = w1399 & ~w21743;
assign w31522 = w1327 & w26476;
assign w31523 = w1478 & ~w26774;
assign w31524 = ~w31521 & ~w31522;
assign w31525 = ~w31520 & w31524;
assign w31526 = ~w31523 & w31525;
assign w31527 = w31519 & ~w31526;
assign w31528 = ~w31519 & w31526;
assign w31529 = ~w31527 & ~w31528;
assign w31530 = w31516 & ~w31529;
assign w31531 = ~w31516 & w31529;
assign w31532 = ~w31530 & ~w31531;
assign w31533 = w3903 & w3933;
assign w31534 = a_26 & ~a_29;
assign w31535 = ~a_26 & a_29;
assign w31536 = ~w31534 & ~w31535;
assign w31537 = ~w31472 & ~w31476;
assign w31538 = w31389 & ~w31401;
assign w31539 = ~w31389 & ~w31452;
assign w31540 = w31461 & ~w31538;
assign w31541 = ~w31539 & w31540;
assign w31542 = w31537 & ~w31541;
assign w31543 = ~w31537 & w31541;
assign w31544 = ~w31542 & ~w31543;
assign w31545 = w31536 & w31544;
assign w31546 = ~w31536 & ~w31544;
assign w31547 = ~w31545 & ~w31546;
assign w31548 = w31533 & ~w31547;
assign w31549 = ~w31533 & w31547;
assign w31550 = ~w31548 & ~w31549;
assign w31551 = w31532 & ~w31550;
assign w31552 = ~w31532 & w31550;
assign w31553 = ~w31551 & ~w31552;
assign w31554 = w31515 & ~w31553;
assign w31555 = ~w31515 & w31553;
assign w31556 = ~w31554 & ~w31555;
assign w31557 = w31507 & w31556;
assign w31558 = ~w31507 & ~w31556;
assign w31559 = ~w31557 & ~w31558;
assign w31560 = ~w68 & ~w458;
assign w31561 = a_26 & w14;
assign w31562 = ~w732 & ~w450;
assign w31563 = ~w239 & ~w356;
assign w31564 = ~w65 & ~w205;
assign w31565 = w2732 & w2277;
assign w31566 = a_26 & w1221;
assign w31567 = w1585 & w2985;
assign w31568 = ~w207 & ~w125;
assign w31569 = w1549 & w1025;
assign w31570 = ~w3202 & w3272;
assign w31571 = ~w1478 & w6199;
assign w31572 = w6188 & w6488;
assign w31573 = ~w6485 & w6487;
assign w31574 = w6501 & w6502;
assign w31575 = ~w6501 & ~w6502;
assign w31576 = w2918 & ~w3053;
assign w31577 = ~w6543 & w6544;
assign w31578 = w6543 & ~w6544;
assign w31579 = w6552 & w1478;
assign w31580 = w6553 & ~w6591;
assign w31581 = ~w6553 & w6591;
assign w31582 = ~w2465 & w1327;
assign w31583 = (w1399 & ~w2587) | (w1399 & w32351) | (~w2587 & w32351);
assign w31584 = ~w6604 & ~w6629;
assign w31585 = w6679 & w32352;
assign w31586 = ~w6734 & ~w6725;
assign w31587 = ~w7268 & w7278;
assign w31588 = w6552 & w4070;
assign w31589 = ~w7291 & a_29;
assign w31590 = w7291 & ~a_29;
assign w31591 = ~w2465 & w4068;
assign w31592 = ~w2588 & w3957;
assign w31593 = ~w2465 & w4446;
assign w31594 = ~w2588 & w4068;
assign w31595 = ~w2588 & w3954;
assign w31596 = ~w2736 & w4068;
assign w31597 = w7348 & a_29;
assign w31598 = ~w7364 & ~w7285;
assign w31599 = w6543 & w7369;
assign w31600 = ~w4070 & w7389;
assign w31601 = w6543 & w7579;
assign w31602 = ~w2588 & ~w518;
assign w31603 = ~w2465 & w4666;
assign w31604 = ~w2588 & w4638;
assign w31605 = ~w2588 & ~w1222;
assign w31606 = ~w1226 & w7630;
assign w31607 = ~w7637 & a_26;
assign w31608 = w7637 & ~a_26;
assign w31609 = w6782 & w1226;
assign w31610 = w7650 & a_26;
assign w31611 = ~w7650 & ~a_26;
assign w31612 = ~w2736 & w4638;
assign w31613 = w7674 & a_26;
assign w31614 = ~w7574 & ~w7591;
assign w31615 = ~w7697 & ~w7575;
assign w31616 = ~w6501 & w7703;
assign w31617 = w3273 & w7749;
assign w31618 = ~w7593 & ~w7591;
assign w31619 = w6543 & w7933;
assign w31620 = w7955 & a_23;
assign w31621 = ~w2465 & w5286;
assign w31622 = ~w2588 & w5080;
assign w31623 = ~w2588 & w504;
assign w31624 = w7983 & a_23;
assign w31625 = ~w7985 & ~w7617;
assign w31626 = ~w5017 & w8002;
assign w31627 = w8006 & ~a_23;
assign w31628 = ~w8006 & a_23;
assign w31629 = w8013 & ~w7968;
assign w31630 = w7644 & ~w7686;
assign w31631 = ~w6501 & w8050;
assign w31632 = ~w8070 & w8074;
assign w31633 = w7718 & w7740;
assign w31634 = ~w8195 & ~w8197;
assign w31635 = ~w5309 & w8309;
assign w31636 = ~w8311 & ~w8312;
assign w31637 = ~w2465 & w5816;
assign w31638 = ~w2588 & w5818;
assign w31639 = ~w2588 & w5300;
assign w31640 = w8334 & a_20;
assign w31641 = ~w8336 & ~w7981;
assign w31642 = ~w5309 & w8355;
assign w31643 = ~w8359 & a_20;
assign w31644 = w8359 & ~a_20;
assign w31645 = ~w6063 & w8389;
assign w31646 = ~w8391 & ~w8392;
assign w31647 = ~w2465 & w6304;
assign w31648 = ~w2588 & w6061;
assign w31649 = ~w2588 & w6054;
assign w31650 = w8414 & a_17;
assign w31651 = ~w8416 & ~w8332;
assign w31652 = ~w6063 & w8435;
assign w31653 = ~w8439 & a_17;
assign w31654 = w8439 & ~a_17;
assign w31655 = ~w6063 & w8456;
assign w31656 = w8336 & w7981;
assign w31657 = w6543 & w8471;
assign w31658 = ~w5309 & w8506;
assign w31659 = w7985 & w7617;
assign w31660 = ~w6447 & w8562;
assign w31661 = ~w8564 & ~w8565;
assign w31662 = ~w2465 & w6996;
assign w31663 = ~w2588 & w6998;
assign w31664 = ~w2588 & w6441;
assign w31665 = w8587 & a_14;
assign w31666 = ~w8589 & ~w8412;
assign w31667 = ~w6447 & w8608;
assign w31668 = ~w8612 & a_14;
assign w31669 = w8612 & ~a_14;
assign w31670 = w6543 & w8628;
assign w31671 = ~w6447 & w8645;
assign w31672 = w8416 & w8332;
assign w31673 = w6489 & w8697;
assign w31674 = w6543 & w8737;
assign w31675 = w6489 & w8758;
assign w31676 = ~w8339 & w8797;
assign w31677 = w8785 & w8809;
assign w31678 = ~w6501 & w8882;
assign w31679 = ~w7193 & w9059;
assign w31680 = ~w9061 & ~w9062;
assign w31681 = ~w2465 & w7511;
assign w31682 = ~w2588 & w7489;
assign w31683 = ~w2588 & w7187;
assign w31684 = w9084 & a_11;
assign w31685 = ~w9086 & ~w8585;
assign w31686 = ~w7193 & w9105;
assign w31687 = ~w9109 & a_11;
assign w31688 = w9109 & ~a_11;
assign w31689 = w6543 & w9125;
assign w31690 = ~w7193 & w9142;
assign w31691 = w8589 & w8412;
assign w31692 = w6489 & w9194;
assign w31693 = w8939 & ~w9264;
assign w31694 = w6489 & w9280;
assign w31695 = ~w9325 & ~w9335;
assign w31696 = w9325 & w9335;
assign w31697 = ~w8278 & w9454;
assign w31698 = ~w9456 & ~w9457;
assign w31699 = ~w2465 & w8295;
assign w31700 = ~w2588 & w8298;
assign w31701 = ~w2588 & ~w8272;
assign w31702 = w9479 & a_8;
assign w31703 = ~w9481 & ~w9082;
assign w31704 = ~w8278 & w9500;
assign w31705 = ~w9504 & a_8;
assign w31706 = w9504 & ~a_8;
assign w31707 = w6543 & w9520;
assign w31708 = ~w8278 & w9537;
assign w31709 = w9086 & w8585;
assign w31710 = w6489 & w9589;
assign w31711 = ~w9263 & ~w8304;
assign w31712 = ~w9790 & w10031;
assign w31713 = ~w10033 & ~w10034;
assign w31714 = w10049 & ~w10045;
assign w31715 = ~w9790 & w10077;
assign w31716 = ~w10081 & a_5;
assign w31717 = w10081 & ~a_5;
assign w31718 = ~w9790 & w10110;
assign w31719 = w9481 & w9082;
assign w31720 = w6489 & w10157;
assign w31721 = w9710 & ~w9744;
assign w31722 = w9743 & ~w9766;
assign w31723 = w9293 & w9855;
assign w31724 = w10504 & w10565;
assign w31725 = w10560 & ~w10650;
assign w31726 = ~w10560 & w10650;
assign w31727 = w10673 & w10635;
assign w31728 = w10616 & w10729;
assign w31729 = w10682 & w10813;
assign w31730 = ~w10837 & w10898;
assign w31731 = ~w10837 & w10913;
assign w31732 = ~w10341 & ~w11237;
assign w31733 = w10341 & ~w10394;
assign w31734 = ~w11269 & ~w11277;
assign w31735 = w11269 & w11277;
assign w31736 = w10543 & ~w10548;
assign w31737 = ~w10804 & w11384;
assign w31738 = ~w11557 & w11568;
assign w31739 = w11557 & ~w11568;
assign w31740 = ~w8155 & ~w11581;
assign w31741 = w8155 & w11581;
assign w31742 = w11609 & w11731;
assign w31743 = ~w11721 & ~w11744;
assign w31744 = w11721 & w11744;
assign w31745 = ~w8158 & w8178;
assign w31746 = w8158 & ~w8178;
assign w31747 = w11819 & ~w11829;
assign w31748 = ~w11709 & ~w11842;
assign w31749 = ~w11790 & w11756;
assign w31750 = w11758 & ~w11877;
assign w31751 = ~w8175 & ~w8179;
assign w31752 = w11708 & w11836;
assign w31753 = w12027 & ~w12026;
assign w31754 = w11981 & w12099;
assign w31755 = w12012 & w12110;
assign w31756 = ~w12012 & ~w12110;
assign w31757 = w12001 & ~w12000;
assign w31758 = ~w12119 & ~w12204;
assign w31759 = w12119 & ~w12204;
assign w31760 = ~w8294 & w12442;
assign w31761 = ~w8294 & w12623;
assign w31762 = ~w12431 & w12438;
assign w31763 = ~w12640 & w12642;
assign w31764 = ~w12640 & ~w12433;
assign w31765 = w8294 & ~w12623;
assign w31766 = w12675 & ~w11825;
assign w31767 = ~w11683 & w11825;
assign w31768 = w11968 & ~w12720;
assign w31769 = ~w11968 & w11976;
assign w31770 = w12721 & ~w12725;
assign w31771 = w11976 & ~w12718;
assign w31772 = ~w11976 & w12718;
assign w31773 = ~w12728 & ~w12741;
assign w31774 = ~w12747 & ~w12100;
assign w31775 = ~w12764 & ~w12779;
assign w31776 = w12397 & ~w12776;
assign w31777 = w12776 & ~w12397;
assign w31778 = ~w12404 & w12790;
assign w31779 = ~w12791 & ~w12796;
assign w31780 = w11976 & w12762;
assign w31781 = w12791 & w12825;
assign w31782 = ~w12847 & ~w12631;
assign w31783 = w14390 & w12673;
assign w31784 = ~w1478 & w14619;
assign w31785 = ~w12833 & w12836;
assign w31786 = ~w12833 & w12835;
assign w31787 = w12822 & ~w12831;
assign w31788 = w14637 & w4070;
assign w31789 = w12780 & w12760;
assign w31790 = ~w15151 & ~w15153;
assign w31791 = ~w12728 & w15155;
assign w31792 = w12728 & w1478;
assign w31793 = w15204 & ~w15240;
assign w31794 = ~w15204 & w15240;
assign w31795 = ~w11501 & w1399;
assign w31796 = ~w1327 & ~w15375;
assign w31797 = ~w15385 & w1478;
assign w31798 = w15242 & ~w15241;
assign w31799 = ~w15433 & ~w15432;
assign w31800 = ~w12763 & w4068;
assign w31801 = w12735 & w3957;
assign w31802 = ~w12732 & w4070;
assign w31803 = ~w12728 & w15931;
assign w31804 = ~w15948 & w15954;
assign w31805 = ~w4068 & ~w15973;
assign w31806 = ~w15385 & w4070;
assign w31807 = ~w4070 & ~w16012;
assign w31808 = w16016 & w15995;
assign w31809 = ~w16016 & ~w15995;
assign w31810 = ~w12675 & w4068;
assign w31811 = ~w11501 & w3957;
assign w31812 = ~w16019 & ~w16017;
assign w31813 = ~w16019 & w16043;
assign w31814 = w16049 & w7269;
assign w31815 = ~w16049 & a_29;
assign w31816 = ~w16086 & ~w15920;
assign w31817 = w14637 & w1226;
assign w31818 = ~w1226 & w16271;
assign w31819 = ~w16296 & ~w16297;
assign w31820 = ~w4638 & ~w16316;
assign w31821 = ~w11501 & ~w518;
assign w31822 = ~w12675 & w4638;
assign w31823 = ~w15385 & w1226;
assign w31824 = ~w11501 & ~w4666;
assign w31825 = w16385 & ~w16339;
assign w31826 = ~w16385 & w16339;
assign w31827 = w16392 & w7680;
assign w31828 = ~w16392 & a_26;
assign w31829 = w16387 & ~w16386;
assign w31830 = ~w16432 & ~w16312;
assign w31831 = ~w16509 & w16265;
assign w31832 = ~w16646 & ~w16647;
assign w31833 = ~w12764 & w5286;
assign w31834 = ~a_23 & w5017;
assign w31835 = ~w15385 & w5017;
assign w31836 = ~w11501 & w5286;
assign w31837 = ~w16705 & ~w16379;
assign w31838 = ~w12675 & w5080;
assign w31839 = ~w11501 & w5016;
assign w31840 = w16706 & ~w16682;
assign w31841 = ~w16706 & w16682;
assign w31842 = w16745 & ~w16727;
assign w31843 = ~w16772 & ~w16660;
assign w31844 = ~w5017 & w16778;
assign w31845 = ~w16314 & ~w16312;
assign w31846 = ~w7961 & w16809;
assign w31847 = ~w16438 & ~w16440;
assign w31848 = ~w14637 & w16872;
assign w31849 = w14637 & w16876;
assign w31850 = ~w16479 & ~w16910;
assign w31851 = w16862 & ~w16864;
assign w31852 = w17237 & ~w17246;
assign w31853 = ~w12764 & w5816;
assign w31854 = ~w15385 & w5309;
assign w31855 = ~w11501 & w5816;
assign w31856 = ~w17354 & ~w16698;
assign w31857 = ~w12675 & w5818;
assign w31858 = ~w11501 & w5308;
assign w31859 = w17355 & ~w17331;
assign w31860 = ~w17355 & w17331;
assign w31861 = w17377 & ~w17376;
assign w31862 = w16705 & w16379;
assign w31863 = ~w17421 & ~w17303;
assign w31864 = w15122 & ~w17427;
assign w31865 = ~w16770 & w17455;
assign w31866 = w16770 & ~w17455;
assign w31867 = ~w17271 & ~w17459;
assign w31868 = ~w17464 & ~w17272;
assign w31869 = ~w16773 & ~w16787;
assign w31870 = w17485 & ~w17502;
assign w31871 = ~w17538 & w17218;
assign w31872 = ~w17153 & ~w17154;
assign w31873 = ~w12764 & w6304;
assign w31874 = ~w15385 & w6063;
assign w31875 = ~w11501 & w6304;
assign w31876 = ~w17751 & ~w17347;
assign w31877 = ~w12675 & w6061;
assign w31878 = ~w11501 & w6059;
assign w31879 = w17752 & ~w17728;
assign w31880 = ~w17752 & w17728;
assign w31881 = w17774 & ~w17773;
assign w31882 = w17354 & w16698;
assign w31883 = ~w17818 & ~w17700;
assign w31884 = w15122 & ~w17824;
assign w31885 = ~w17420 & w17852;
assign w31886 = w17420 & ~w17852;
assign w31887 = ~w17667 & ~w17856;
assign w31888 = ~w17861 & ~w17668;
assign w31889 = ~w12764 & w6996;
assign w31890 = ~w15385 & w6447;
assign w31891 = ~w11501 & w6996;
assign w31892 = ~w17990 & ~w17744;
assign w31893 = ~w12675 & w6998;
assign w31894 = ~w11501 & w6446;
assign w31895 = w17991 & ~w17967;
assign w31896 = ~w17991 & w17967;
assign w31897 = w18013 & ~w18012;
assign w31898 = w17751 & w17347;
assign w31899 = ~w18057 & ~w17939;
assign w31900 = w15122 & ~w18063;
assign w31901 = ~w17817 & w18091;
assign w31902 = w17817 & ~w18091;
assign w31903 = ~w17906 & ~w18095;
assign w31904 = ~w18100 & ~w17907;
assign w31905 = ~w17858 & ~w17856;
assign w31906 = w17881 & ~w18184;
assign w31907 = ~w17461 & ~w17459;
assign w31908 = ~w12764 & w7511;
assign w31909 = ~w15385 & w7193;
assign w31910 = ~w11501 & w7511;
assign w31911 = ~w18454 & ~w17983;
assign w31912 = ~w12675 & w7489;
assign w31913 = ~w18455 & w18431;
assign w31914 = w18455 & ~w18431;
assign w31915 = w18477 & ~w18476;
assign w31916 = w17990 & w17744;
assign w31917 = ~w18521 & ~w18403;
assign w31918 = w15122 & ~w18527;
assign w31919 = ~w18056 & w18555;
assign w31920 = w18056 & ~w18555;
assign w31921 = ~w18370 & ~w18559;
assign w31922 = ~w18564 & ~w18371;
assign w31923 = ~w18097 & ~w18095;
assign w31924 = w18120 & ~w18137;
assign w31925 = ~w18827 & ~w18847;
assign w31926 = w18827 & w18847;
assign w31927 = w18898 & w18897;
assign w31928 = w18584 & ~w18601;
assign w31929 = ~w12764 & w8295;
assign w31930 = ~w15385 & w8278;
assign w31931 = ~w8278 & ~w19103;
assign w31932 = ~w11501 & w8295;
assign w31933 = w19110 & w18447;
assign w31934 = ~w19110 & ~w18447;
assign w31935 = ~w11501 & w8277;
assign w31936 = ~w19113 & ~w19111;
assign w31937 = w18454 & w17983;
assign w31938 = ~w19197 & ~w19069;
assign w31939 = w15122 & ~w19204;
assign w31940 = ~w18520 & w19232;
assign w31941 = w18520 & ~w19232;
assign w31942 = ~w19036 & ~w19236;
assign w31943 = ~w19241 & ~w19037;
assign w31944 = ~w18561 & ~w18559;
assign w31945 = w19379 & ~w18765;
assign w31946 = w18357 & w18886;
assign w31947 = ~w19398 & w19407;
assign w31948 = w19339 & ~w18974;
assign w31949 = ~w9790 & w19571;
assign w31950 = ~w9790 & w19573;
assign w31951 = ~w9790 & ~w19603;
assign w31952 = w19606 & w19596;
assign w31953 = w15122 & ~w19670;
assign w31954 = w19196 & w19697;
assign w31955 = ~w19196 & ~w19697;
assign w31956 = ~w19534 & ~w19701;
assign w31957 = ~w19706 & ~w19535;
assign w31958 = ~w19198 & ~w19214;
assign w31959 = ~w19521 & ~w19723;
assign w31960 = ~w19238 & ~w19236;
assign w31961 = w19261 & ~w19278;
assign w31962 = ~w18898 & ~w18897;
assign w31963 = w19434 & w19433;
assign w31964 = w19977 & ~w19424;
assign w31965 = w18866 & ~w18867;
assign w31966 = w18853 & ~w19985;
assign w31967 = w18825 & ~w18824;
assign w31968 = ~w17237 & w17246;
assign w31969 = ~w17530 & ~w17532;
assign w31970 = w17537 & ~w20234;
assign w31971 = ~w17537 & w20234;
assign w31972 = w20287 & ~w20289;
assign w31973 = w20240 & w20294;
assign w31974 = w20263 & w20345;
assign w31975 = w17539 & w17541;
assign w31976 = ~w20508 & ~w20513;
assign w31977 = w20518 & ~w20520;
assign w31978 = w20452 & w20544;
assign w31979 = w20457 & w20575;
assign w31980 = ~w20457 & ~w20575;
assign w31981 = ~w20512 & w20618;
assign w31982 = w20914 & ~w20901;
assign w31983 = w20916 & ~w20930;
assign w31984 = w19839 & ~w19860;
assign w31985 = w20975 & ~w20961;
assign w31986 = w19875 & w19475;
assign w31987 = ~w21028 & ~w21036;
assign w31988 = w21028 & w21036;
assign w31989 = ~w20388 & ~w20391;
assign w31990 = ~w20382 & w21218;
assign w31991 = w21224 & w21230;
assign w31992 = w21602 & ~w21596;
assign w31993 = ~w21681 & w21687;
assign w31994 = ~w21185 & ~w21206;
assign w31995 = w21185 & ~w21199;
assign w31996 = ~w21804 & ~w21830;
assign w31997 = ~w21224 & ~w21230;
assign w31998 = w21206 & ~w21846;
assign w31999 = w21839 & ~w21871;
assign w32000 = w21475 & w21643;
assign w32001 = w21475 & ~w21890;
assign w32002 = (~w21907 & w21643) | (~w21907 & w32353) | (w21643 & w32353);
assign w32003 = ~w21643 & w32354;
assign w32004 = w21905 & ~w21911;
assign w32005 = (~w21670 & w21607) | (~w21670 & w32355) | (w21607 & w32355);
assign w32006 = (~w21643 & w32356) | (~w21643 & w32357) | (w32356 & w32357);
assign w32007 = ~w21680 & w17633;
assign w32008 = ~w21677 & ~w21930;
assign w32009 = ~w21956 & ~w21952;
assign w32010 = ~w21952 & ~w21961;
assign w32011 = ~w21681 & ~w21686;
assign w32012 = ~w21681 & w21982;
assign w32013 = ~w21681 & w21987;
assign w32014 = w22018 & ~w22021;
assign w32015 = ~w21953 & ~w21911;
assign w32016 = ~w6447 & w22101;
assign w32017 = w21835 & w21872;
assign w32018 = (w6063 & w21240) | (w6063 & w32358) | (w21240 & w32358);
assign w32019 = w21815 & w5017;
assign w32020 = ~w21815 & w5017;
assign w32021 = ~w21817 & w32359;
assign w32022 = ~w21797 & w5816;
assign w32023 = ~w21813 & w5309;
assign w32024 = w21815 & w5309;
assign w32025 = ~w21815 & w5309;
assign w32026 = ~w22158 & a_20;
assign w32027 = (~a_20 & w22137) | (~a_20 & w32360) | (w22137 & w32360);
assign w32028 = ~w21819 & w32361;
assign w32029 = w21798 & w5309;
assign w32030 = ~w22177 & w32362;
assign w32031 = (~a_20 & w22177) | (~a_20 & w32363) | (w22177 & w32363);
assign w32032 = ~w21797 & w5308;
assign w32033 = ~w22245 & w22253;
assign w32034 = w21804 & ~w21830;
assign w32035 = ~w21184 & w6059;
assign w32036 = ~w22298 & ~a_17;
assign w32037 = w21818 & w6063;
assign w32038 = ~w21797 & w6304;
assign w32039 = ~w21813 & w6063;
assign w32040 = (~w6304 & ~w21815) | (~w6304 & w32364) | (~w21815 & w32364);
assign w32041 = (a_17 & ~w22336) | (a_17 & w32365) | (~w22336 & w32365);
assign w32042 = (a_17 & w22332) | (a_17 & w32366) | (w22332 & w32366);
assign w32043 = ~w22321 & ~a_17;
assign w32044 = w21822 & w6063;
assign w32045 = ~w21821 & w6063;
assign w32046 = w22356 & a_17;
assign w32047 = ~w22356 & ~a_17;
assign w32048 = w22286 & ~w22285;
assign w32049 = (w6447 & w21882) | (w6447 & w32367) | (w21882 & w32367);
assign w32050 = ~w21792 & w6447;
assign w32051 = ~w21893 & w6996;
assign w32052 = w22381 & w32368;
assign w32053 = (~a_14 & ~w22381) | (~a_14 & w32369) | (~w22381 & w32369);
assign w32054 = ~w21784 & w6447;
assign w32055 = ~w22245 & w22427;
assign w32056 = ~w21817 & w32370;
assign w32057 = ~w21797 & w6996;
assign w32058 = ~w21813 & w6447;
assign w32059 = (~w6996 & ~w21815) | (~w6996 & w32371) | (~w21815 & w32371);
assign w32060 = (a_14 & ~w22470) | (a_14 & w32372) | (~w22470 & w32372);
assign w32061 = (a_14 & w22466) | (a_14 & w32373) | (w22466 & w32373);
assign w32062 = (~a_14 & w22137) | (~a_14 & w32374) | (w22137 & w32374);
assign w32063 = ~w21819 & w32375;
assign w32064 = ~w21821 & w6447;
assign w32065 = ~w22177 & w32376;
assign w32066 = (~a_14 & w22177) | (~a_14 & w32377) | (w22177 & w32377);
assign w32067 = ~w21797 & w6446;
assign w32068 = w22502 & ~w22539;
assign w32069 = (~w21914 & w21904) | (~w21914 & w32378) | (w21904 & w32378);
assign w32070 = (w6063 & w21882) | (w6063 & w32379) | (w21882 & w32379);
assign w32071 = ~w21792 & w6063;
assign w32072 = ~w21893 & w6304;
assign w32073 = w22381 & w32380;
assign w32074 = (~a_17 & ~w22381) | (~a_17 & w32381) | (~w22381 & w32381);
assign w32075 = w22190 & ~w22234;
assign w32076 = ~w21797 & w5286;
assign w32077 = ~w21813 & w5017;
assign w32078 = w22192 & a_23;
assign w32079 = ~w22662 & ~w22661;
assign w32080 = ~w7193 & w22680;
assign w32081 = (w7193 & w21882) | (w7193 & w32382) | (w21882 & w32382);
assign w32082 = ~w21792 & w7193;
assign w32083 = ~w21893 & w7511;
assign w32084 = (~a_11 & ~w22381) | (~a_11 & w32383) | (~w22381 & w32383);
assign w32085 = w22381 & w32384;
assign w32086 = ~w22245 & w22747;
assign w32087 = ~w21817 & w32385;
assign w32088 = ~w21797 & w7511;
assign w32089 = ~w21813 & w7193;
assign w32090 = (~w7511 & ~w21815) | (~w7511 & w32386) | (~w21815 & w32386);
assign w32091 = (a_11 & ~w22789) | (a_11 & w32387) | (~w22789 & w32387);
assign w32092 = (a_11 & w22785) | (a_11 & w32388) | (w22785 & w32388);
assign w32093 = (~a_11 & w22137) | (~a_11 & w32389) | (w22137 & w32389);
assign w32094 = ~w21819 & w32390;
assign w32095 = ~w21821 & w7193;
assign w32096 = ~w22177 & w32391;
assign w32097 = (~a_11 & w22177) | (~a_11 & w32392) | (w22177 & w32392);
assign w32098 = ~w21797 & w7192;
assign w32099 = w22821 & ~w22858;
assign w32100 = ~w21963 & w22927;
assign w32101 = ~w22245 & w22971;
assign w32102 = w22980 & ~w22977;
assign w32103 = w22984 & ~w22983;
assign w32104 = ~w22984 & w22983;
assign w32105 = w21822 & w5017;
assign w32106 = ~w21821 & w5017;
assign w32107 = ~w22990 & ~a_23;
assign w32108 = w22990 & a_23;
assign w32109 = w21915 & ~w21961;
assign w32110 = w21956 & ~w21961;
assign w32111 = ~w8278 & w23070;
assign w32112 = (w8278 & w21240) | (w8278 & w32393) | (w21240 & w32393);
assign w32113 = ~w22245 & w23117;
assign w32114 = ~w21804 & w21830;
assign w32115 = ~w21817 & w32394;
assign w32116 = ~w21797 & w8295;
assign w32117 = ~w21813 & w8278;
assign w32118 = (~w8295 & ~w21815) | (~w8295 & w32395) | (~w21815 & w32395);
assign w32119 = (a_8 & ~w23175) | (a_8 & w32396) | (~w23175 & w32396);
assign w32120 = (a_8 & w23173) | (a_8 & w32397) | (w23173 & w32397);
assign w32121 = (~a_8 & w22137) | (~a_8 & w32398) | (w22137 & w32398);
assign w32122 = ~w21819 & w32399;
assign w32123 = ~w21821 & w8278;
assign w32124 = ~w22177 & w32400;
assign w32125 = (~a_8 & w22177) | (~a_8 & w32401) | (w22177 & w32401);
assign w32126 = ~w22904 & w9484;
assign w32127 = (w9456 & ~w22663) | (w9456 & w32402) | (~w22663 & w32402);
assign w32128 = ~w22001 & w22011;
assign w32129 = (w5309 & w21240) | (w5309 & w32403) | (w21240 & w32403);
assign w32130 = ~w21184 & w5016;
assign w32131 = ~w23477 & ~a_23;
assign w32132 = ~w6063 & w23518;
assign w32133 = ~w23733 & w32404;
assign w32134 = ~w23740 & w32405;
assign w32135 = ~w9790 & w23770;
assign w32136 = w23774 & ~w23793;
assign w32137 = (w5309 & w21882) | (w5309 & w32406) | (w21882 & w32406);
assign w32138 = ~w21792 & w5309;
assign w32139 = ~w21893 & w5816;
assign w32140 = w22381 & w32407;
assign w32141 = (~a_20 & ~w22381) | (~a_20 & w32408) | (~w22381 & w32408);
assign w32142 = w21818 & w1226;
assign w32143 = ~w21797 & w4666;
assign w32144 = ~w21813 & w1226;
assign w32145 = ~w24021 & w24020;
assign w32146 = w24021 & ~w24020;
assign w32147 = ~w22245 & w24191;
assign w32148 = ~w24021 & ~a_26;
assign w32149 = w21822 & w1226;
assign w32150 = ~w21821 & w1226;
assign w32151 = w24216 & a_26;
assign w32152 = ~w24216 & ~a_26;
assign w32153 = w24050 & ~w24049;
assign w32154 = (w5017 & w21240) | (w5017 & w32409) | (w21240 & w32409);
assign w32155 = ~w21184 & ~w518;
assign w32156 = ~w24368 & ~a_26;
assign w32157 = ~w4068 & ~w24396;
assign w32158 = ~w5309 & w24424;
assign w32159 = (w8419 & ~w22663) | (w8419 & w32410) | (~w22663 & w32410);
assign w32160 = (w5017 & w21882) | (w5017 & w32411) | (w21882 & w32411);
assign w32161 = ~w21792 & w5017;
assign w32162 = ~w21893 & w5286;
assign w32163 = (~a_23 & ~w22381) | (~a_23 & w32412) | (~w22381 & w32412);
assign w32164 = w22381 & w32413;
assign w32165 = ~w21797 & w4446;
assign w32166 = w21813 & w4070;
assign w32167 = ~w21797 & w4070;
assign w32168 = ~w24598 & a_29;
assign w32169 = ~w24623 & a_26;
assign w32170 = ~w6063 & w24678;
assign w32171 = w24473 & w24703;
assign w32172 = w24578 & w24667;
assign w32173 = ~w22245 & w24793;
assign w32174 = w24604 & ~w24610;
assign w32175 = w21815 & w1478;
assign w32176 = ~a_31 & ~w1477;
assign w32177 = ~w24802 & ~w24801;
assign w32178 = ~w21819 & w32414;
assign w32179 = ~w21821 & w4070;
assign w32180 = (~a_29 & w22177) | (~a_29 & w32415) | (w22177 & w32415);
assign w32181 = ~w22177 & w32416;
assign w32182 = w24634 & ~w24635;
assign w32183 = ~w24523 & ~w24946;
assign w32184 = ~w24770 & ~w24989;
assign w32185 = w24770 & w24989;
assign w32186 = w24740 & ~w25000;
assign w32187 = ~w5017 & w25009;
assign w32188 = (w1226 & w21240) | (w1226 & w32417) | (w21240 & w32417);
assign w32189 = (w5309 & ~w22663) | (w5309 & w32418) | (~w22663 & w32418);
assign w32190 = (w8419 & w23030) | (w8419 & w32419) | (w23030 & w32419);
assign w32191 = w24987 & ~w25120;
assign w32192 = ~w24987 & w25120;
assign w32193 = w24976 & ~w25150;
assign w32194 = (~w24987 & ~w25120) | (~w24987 & w32420) | (~w25120 & w32420);
assign w32195 = (w24987 & w25120) | (w24987 & w32634) | (w25120 & w32634);
assign w32196 = ~w25188 & ~w25183;
assign w32197 = ~w25225 & ~w25217;
assign w32198 = w21813 & w1478;
assign w32199 = ~w21813 & w1478;
assign w32200 = ~w21797 & w668;
assign w32201 = ~w25274 & ~w25291;
assign w32202 = w25051 & ~w25050;
assign w32203 = (w1226 & w21882) | (w1226 & w32421) | (w21882 & w32421);
assign w32204 = ~w21792 & w1226;
assign w32205 = ~w21893 & w4666;
assign w32206 = w22381 & w32422;
assign w32207 = (~a_26 & ~w22381) | (~a_26 & w32423) | (~w22381 & w32423);
assign w32208 = w25156 & ~w25179;
assign w32209 = ~w25456 & w25448;
assign w32210 = w21821 & w1478;
assign w32211 = ~w21821 & w1478;
assign w32212 = w25496 & ~w25516;
assign w32213 = w25294 & a_29;
assign w32214 = ~w25294 & ~a_29;
assign w32215 = w25540 & w7680;
assign w32216 = (~w4403 & w25540) | (~w4403 & w32424) | (w25540 & w32424);
assign w32217 = ~w25646 & w25388;
assign w32218 = ~w10837 & w25804;
assign w32219 = ~w25830 & w32425;
assign w32220 = w24520 & ~w24951;
assign w32221 = ~w24952 & ~w24954;
assign w32222 = (~w25706 & ~w26162) | (~w25706 & w32426) | (~w26162 & w32426);
assign w32223 = ~w25667 & ~w26198;
assign w32224 = w25545 & ~w25319;
assign w32225 = ~w1226 & w26274;
assign w32226 = (a_29 & ~w22247) | (a_29 & w32427) | (~w22247 & w32427);
assign w32227 = w22247 & w32428;
assign w32228 = w25486 & ~w26284;
assign w32229 = (w4070 & w21240) | (w4070 & w32429) | (w21240 & w32429);
assign w32230 = ~w21797 & w1399;
assign w32231 = w25683 & ~w25682;
assign w32232 = ~w26523 & ~w26527;
assign w32233 = ~w26571 & w32430;
assign w32234 = w26341 & a_29;
assign w32235 = ~w26341 & ~a_29;
assign w32236 = ~w5017 & w26636;
assign w32237 = ~w26803 & ~w26798;
assign w32238 = w26551 & w26829;
assign w32239 = w26677 & w26651;
assign w32240 = w26613 & ~w26888;
assign w32241 = w26894 & w7269;
assign w32242 = (~w7268 & w26894) | (~w7268 & w32431) | (w26894 & w32431);
assign w32243 = ~w26628 & ~w26359;
assign w32244 = w27104 & ~w27103;
assign w32245 = ~w27166 & ~w26928;
assign w32246 = w26922 & ~w26921;
assign w32247 = (w1226 & ~w22663) | (w1226 & w32432) | (~w22663 & w32432);
assign w32248 = w23309 & w27233;
assign w32249 = w26870 & ~w27164;
assign w32250 = ~w27283 & ~w27387;
assign w32251 = (w27274 & w27249) | (w27274 & w32433) | (w27249 & w32433);
assign w32252 = ~w27250 & ~w27417;
assign w32253 = ~w27424 & ~w27192;
assign w32254 = ~w27428 & w32434;
assign w32255 = w27198 & ~w26928;
assign w32256 = ~w27473 & ~w27212;
assign w32257 = ~w1226 & w27479;
assign w32258 = ~w27654 & ~w27656;
assign w32259 = ~w27678 & ~w27672;
assign w32260 = ~w1478 & w27698;
assign w32261 = ~w27866 & ~w27789;
assign w32262 = ~w27866 & ~w27874;
assign w32263 = ~w22904 & w4070;
assign w32264 = ~w1478 & w27943;
assign w32265 = ~w28115 & ~w28114;
assign w32266 = w27895 & ~w28010;
assign w32267 = w28132 & ~w28131;
assign w32268 = ~w28134 & w28158;
assign w32269 = w28134 & ~w28158;
assign w32270 = ~w28162 & w27988;
assign w32271 = ~w1478 & w28190;
assign w32272 = ~w4070 & w28202;
assign w32273 = ~w1226 & w28214;
assign w32274 = ~w27717 & ~w27971;
assign w32275 = ~w28275 & w28283;
assign w32276 = ~w27849 & w28054;
assign w32277 = w27849 & ~w28054;
assign w32278 = ~w28309 & w28305;
assign w32279 = w28309 & ~w28305;
assign w32280 = w28309 & ~w28304;
assign w32281 = ~w28102 & ~w28269;
assign w32282 = w28163 & ~w28370;
assign w32283 = w28206 & ~w28195;
assign w32284 = w28223 & ~w28219;
assign w32285 = ~w28371 & ~w28458;
assign w32286 = w28371 & w28458;
assign w32287 = w28480 & ~w28479;
assign w32288 = ~w28263 & ~w28497;
assign w32289 = ~w6447 & w28542;
assign w32290 = ~w28698 & ~w28735;
assign w32291 = w28698 & w28735;
assign w32292 = w28668 & w28550;
assign w32293 = w28537 & ~w28682;
assign w32294 = ~w28907 & ~w28715;
assign w32295 = ~w4070 & w29004;
assign w32296 = ~w23030 & w1478;
assign w32297 = ~w28914 & w29115;
assign w32298 = ~w29108 & ~w29106;
assign w32299 = w29110 & ~w29306;
assign w32300 = ~w29110 & w29306;
assign w32301 = ~w28907 & w29478;
assign w32302 = ~w29483 & w29487;
assign w32303 = ~w1478 & w29572;
assign w32304 = ~w29124 & w29641;
assign w32305 = ~w29656 & ~w29652;
assign w32306 = w29482 & ~w29649;
assign w32307 = ~w29659 & ~w29658;
assign w32308 = ~w28907 & w29667;
assign w32309 = ~w6063 & w29696;
assign w32310 = ~w8391 & ~w29698;
assign w32311 = ~w4070 & w29727;
assign w32312 = ~w29669 & ~w29817;
assign w32313 = w29669 & w29817;
assign w32314 = ~w1478 & w29888;
assign w32315 = ~w29982 & ~w29981;
assign w32316 = ~w29986 & ~w29985;
assign w32317 = w29994 & w29980;
assign w32318 = ~w6063 & w30115;
assign w32319 = ~w8391 & ~w30117;
assign w32320 = w29989 & ~w30139;
assign w32321 = ~w5017 & w30215;
assign w32322 = w29994 & ~w30131;
assign w32323 = w30270 & ~w30269;
assign w32324 = w29820 & w30280;
assign w32325 = ~w29668 & w30410;
assign w32326 = ~w29668 & w30532;
assign w32327 = ~w30550 & w30663;
assign w32328 = ~w30667 & ~w30668;
assign w32329 = w30666 & w30774;
assign w32330 = ~w30667 & w30780;
assign w32331 = w30670 & w30783;
assign w32332 = ~w29668 & w30884;
assign w32333 = w30415 & w30889;
assign w32334 = ~w30785 & w30896;
assign w32335 = ~w30903 & w30997;
assign w32336 = w30902 & ~w30993;
assign w32337 = w30902 & ~w31096;
assign w32338 = w30902 & w31104;
assign w32339 = w30902 & w31195;
assign w32340 = ~w31198 & ~w31194;
assign w32341 = ~w31206 & w31202;
assign w32342 = ~w31198 & ~w31283;
assign w32343 = w31198 & ~w31280;
assign w32344 = ~w31204 & w31286;
assign w32345 = w31204 & ~w31286;
assign w32346 = ~w31357 & ~w31360;
assign w32347 = ~w31363 & w31364;
assign w32348 = ~w31204 & w31366;
assign w32349 = w31204 & w31370;
assign w32350 = ~w31447 & w31448;
assign w32351 = ~w2584 & w1399;
assign w32352 = ~w6678 & ~w1478;
assign w32353 = w21607 & ~w21907;
assign w32354 = ~w21607 & w21907;
assign w32355 = w21635 & ~w21670;
assign w32356 = ~w21916 & w21670;
assign w32357 = ~w21916 & ~w32005;
assign w32358 = w21370 & w6063;
assign w32359 = w21813 & w5309;
assign w32360 = ~w32021 & ~a_20;
assign w32361 = w21821 & w5309;
assign w32362 = w32028 & a_20;
assign w32363 = ~w32028 & ~a_20;
assign w32364 = ~w6061 & ~w6304;
assign w32365 = w22334 & a_17;
assign w32366 = w32041 & a_17;
assign w32367 = w21792 & w6447;
assign w32368 = w32049 & a_14;
assign w32369 = ~w32049 & ~a_14;
assign w32370 = w21813 & w6447;
assign w32371 = ~w6998 & ~w6996;
assign w32372 = w22468 & a_14;
assign w32373 = w32060 & a_14;
assign w32374 = ~w32056 & ~a_14;
assign w32375 = w21821 & w6447;
assign w32376 = w32063 & a_14;
assign w32377 = ~w32063 & ~a_14;
assign w32378 = w21902 & ~w21914;
assign w32379 = w21792 & w6063;
assign w32380 = w32070 & a_17;
assign w32381 = ~w32070 & ~a_17;
assign w32382 = w21792 & w7193;
assign w32383 = ~w32081 & ~a_11;
assign w32384 = w32081 & a_11;
assign w32385 = w21813 & w7193;
assign w32386 = ~w7489 & ~w7511;
assign w32387 = w22787 & a_11;
assign w32388 = w32091 & a_11;
assign w32389 = ~w32087 & ~a_11;
assign w32390 = w21821 & w7193;
assign w32391 = w32094 & a_11;
assign w32392 = ~w32094 & ~a_11;
assign w32393 = w21370 & w8278;
assign w32394 = w21813 & w8278;
assign w32395 = ~w8298 & ~w8295;
assign w32396 = w23177 & a_8;
assign w32397 = w32119 & a_8;
assign w32398 = ~w32115 & ~a_8;
assign w32399 = w21821 & w8278;
assign w32400 = w32122 & a_8;
assign w32401 = ~w32122 & ~a_8;
assign w32402 = w22903 & w9456;
assign w32403 = w21370 & w5309;
assign w32404 = w23734 & ~w9790;
assign w32405 = ~w23741 & ~w23738;
assign w32406 = w21792 & w5309;
assign w32407 = w32137 & a_20;
assign w32408 = ~w32137 & ~a_20;
assign w32409 = w21370 & w5017;
assign w32410 = w22903 & w8419;
assign w32411 = w21792 & w5017;
assign w32412 = ~w32160 & ~a_23;
assign w32413 = w32160 & a_23;
assign w32414 = w21821 & w4070;
assign w32415 = ~w32178 & ~a_29;
assign w32416 = w32178 & a_29;
assign w32417 = w21370 & w1226;
assign w32418 = w22903 & w5309;
assign w32419 = ~w23308 & w8419;
assign w32420 = w25141 & ~w24987;
assign w32421 = w21792 & w1226;
assign w32422 = w32203 & a_26;
assign w32423 = ~w32203 & ~a_26;
assign w32424 = ~a_26 & ~w4403;
assign w32425 = ~w25831 & ~w10837;
assign w32426 = ~w26172 & ~w25706;
assign w32427 = ~w4070 & a_29;
assign w32428 = w4070 & ~a_29;
assign w32429 = w21370 & w4070;
assign w32430 = w26572 & ~w4070;
assign w32431 = ~a_29 & ~w7268;
assign w32432 = w22903 & w1226;
assign w32433 = w27164 & w27274;
assign w32434 = w27429 & ~w1478;
assign w32435 = w6187 & ~w6199;
assign w32436 = w6187 & ~w31571;
assign w32437 = ~w1478 & w6786;
assign w32438 = ~w6792 & ~w6551;
assign w32439 = w6782 & w5017;
assign w32440 = ~w8021 & ~a_23;
assign w32441 = w8021 & a_23;
assign w32442 = ~w11894 & ~w11892;
assign w32443 = ~w12153 & ~w12152;
assign w32444 = ~w12268 & ~w12267;
assign w32445 = w12403 & w12391;
assign w32446 = w12644 & ~w12642;
assign w32447 = w12644 & ~w31763;
assign w32448 = ~w12641 & w12433;
assign w32449 = ~w12641 & ~w31764;
assign w32450 = ~w12100 & ~w12776;
assign w32451 = ~w12405 & ~w12407;
assign w32452 = ~w12798 & ~w12826;
assign w32453 = ~w12652 & ~w12648;
assign w32454 = w12658 & ~w12648;
assign w32455 = ~w21636 & w21672;
assign w32456 = ~w21673 & w21680;
assign w32457 = ~w21636 & w21917;
assign w32458 = ~w21932 & ~w21929;
assign w32459 = ~w21673 & w21931;
assign w32460 = w32008 & ~w21930;
assign w32461 = (~w21930 & w32008) | (~w21930 & w21673) | (w32008 & w21673);
assign w32462 = ~w21918 & w21948;
assign w32463 = ~w21673 & ~w21676;
assign w32464 = w22077 & w22080;
assign w32465 = ~w22077 & ~w22080;
assign w32466 = a_14 & ~w22101;
assign w32467 = a_14 & ~w32016;
assign w32468 = ~a_14 & w22101;
assign w32469 = ~a_14 & w32016;
assign w32470 = w22129 & ~a_20;
assign w32471 = w22129 & ~w32026;
assign w32472 = w22159 & ~w22129;
assign w32473 = ~w22319 & ~w22288;
assign w32474 = w22153 & ~a_17;
assign w32475 = w22153 & ~w32042;
assign w32476 = w22368 & ~w22320;
assign w32477 = ~w22153 & a_17;
assign w32478 = ~w22153 & w32042;
assign w32479 = w8564 & ~w22443;
assign w32480 = w22333 & ~a_14;
assign w32481 = w22333 & ~w32061;
assign w32482 = w22473 & ~w22333;
assign w32483 = ~w8564 & w22443;
assign w32484 = w22577 & ~w21914;
assign w32485 = w22577 & w32069;
assign w32486 = ~w22577 & w21914;
assign w32487 = ~w22577 & ~w32069;
assign w32488 = w22240 & ~w22239;
assign w32489 = a_11 & ~w22680;
assign w32490 = a_11 & ~w32080;
assign w32491 = ~a_11 & w22680;
assign w32492 = ~a_11 & w32080;
assign w32493 = w22467 & ~a_11;
assign w32494 = w22467 & ~w32092;
assign w32495 = w22792 & ~w22467;
assign w32496 = w22767 & ~w22772;
assign w32497 = w22421 & ~w22549;
assign w32498 = ~w22688 & ~w22891;
assign w32499 = ~w22670 & ~w22893;
assign w32500 = w22077 & ~w21952;
assign w32501 = w22570 & ~w22572;
assign w32502 = w22089 & ~w22918;
assign w32503 = ~w22380 & ~w22649;
assign w32504 = w23028 & ~w23027;
assign w32505 = a_8 & ~w23070;
assign w32506 = a_8 & ~w32111;
assign w32507 = ~a_8 & w23070;
assign w32508 = ~a_8 & w32111;
assign w32509 = ~w8278 & w23081;
assign w32510 = w23135 & ~w23134;
assign w32511 = w23151 & ~w23148;
assign w32512 = w22786 & ~a_8;
assign w32513 = w22786 & ~w32120;
assign w32514 = w23180 & ~w22786;
assign w32515 = w22703 & ~w22871;
assign w32516 = w22901 & w23285;
assign w32517 = ~w23029 & w23308;
assign w32518 = ~w23361 & ~w23385;
assign w32519 = w23386 & w23049;
assign w32520 = w22952 & ~w22648;
assign w32521 = w23013 & ~w23014;
assign w32522 = ~w23498 & ~w23468;
assign w32523 = a_17 & ~w23518;
assign w32524 = a_17 & ~w32132;
assign w32525 = ~a_17 & w23518;
assign w32526 = ~a_17 & w32132;
assign w32527 = ~w9790 & w23668;
assign w32528 = ~w9790 & w23702;
assign w32529 = ~w23717 & w23716;
assign w32530 = ~w32134 & a_5;
assign w32531 = w23745 & a_5;
assign w32532 = ~a_5 & w32133;
assign w32533 = ~a_5 & w23735;
assign w32534 = ~a_5 & w23770;
assign w32535 = ~a_5 & w32135;
assign w32536 = a_5 & ~w23770;
assign w32537 = a_5 & ~w32135;
assign w32538 = ~w23787 & ~w23789;
assign w32539 = w23089 & ~w23221;
assign w32540 = ~w23854 & ~w23841;
assign w32541 = ~w23890 & ~w23878;
assign w32542 = ~w23619 & ~w23916;
assign w32543 = ~w23921 & ~w23620;
assign w32544 = w23386 & w23936;
assign w32545 = ~w23348 & ~w23354;
assign w32546 = w23457 & ~w23499;
assign w32547 = w24076 & ~w23980;
assign w32548 = w24244 & ~w24338;
assign w32549 = ~w24244 & w24338;
assign w32550 = w24239 & ~w24238;
assign w32551 = ~w24389 & ~w24402;
assign w32552 = a_20 & ~w24424;
assign w32553 = a_20 & ~w32158;
assign w32554 = ~a_20 & w24424;
assign w32555 = ~a_20 & w32158;
assign w32556 = w24407 & ~w24403;
assign w32557 = w24623 & ~a_26;
assign w32558 = w24623 & w7680;
assign w32559 = ~w5017 & w24784;
assign w32560 = ~w24770 & w24930;
assign w32561 = w24770 & ~w24930;
assign w32562 = a_23 & ~w25009;
assign w32563 = a_23 & ~w32187;
assign w32564 = ~a_23 & w25009;
assign w32565 = ~a_23 & w32187;
assign w32566 = ~w4070 & w25032;
assign w32567 = w25228 & ~w25227;
assign w32568 = w25079 & ~w25078;
assign w32569 = ~w25066 & w25071;
assign w32570 = w25087 & ~w25324;
assign w32571 = ~w25495 & w25516;
assign w32572 = ~w25301 & ~w25486;
assign w32573 = ~a_2 & ~w25804;
assign w32574 = ~a_2 & ~w32218;
assign w32575 = a_2 & w25804;
assign w32576 = a_2 & w32218;
assign w32577 = ~w10837 & w25812;
assign w32578 = ~a_2 & ~w32219;
assign w32579 = ~a_2 & ~w25832;
assign w32580 = a_2 & w32219;
assign w32581 = a_2 & w25832;
assign w32582 = ~w10837 & w25895;
assign w32583 = ~w10837 & w25909;
assign w32584 = ~w23880 & ~w23878;
assign w32585 = ~w23897 & ~w23899;
assign w32586 = ~w25758 & ~w26030;
assign w32587 = ~w23918 & ~w23916;
assign w32588 = w26195 & w25656;
assign w32589 = a_26 & ~w26274;
assign w32590 = a_26 & ~w32225;
assign w32591 = ~a_26 & w26274;
assign w32592 = ~a_26 & w32225;
assign w32593 = ~w25485 & ~w25325;
assign w32594 = ~w26227 & w26215;
assign w32595 = ~w26436 & w26517;
assign w32596 = w26381 & ~w26378;
assign w32597 = w25533 & ~w26354;
assign w32598 = ~w1478 & w26580;
assign w32599 = ~w26678 & ~w26691;
assign w32600 = w26678 & w26691;
assign w32601 = w26498 & w26788;
assign w32602 = ~w26789 & ~w26796;
assign w32603 = ~w26737 & w26541;
assign w32604 = ~w26697 & w26691;
assign w32605 = w26838 & ~w26840;
assign w32606 = ~a_29 & ~w32233;
assign w32607 = ~a_29 & ~w26573;
assign w32608 = a_29 & w32233;
assign w32609 = a_29 & w26573;
assign w32610 = w26602 & ~w26600;
assign w32611 = ~w1478 & w26905;
assign w32612 = ~w27007 & w27122;
assign w32613 = ~w26972 & w26651;
assign w32614 = ~w26972 & ~w26857;
assign w32615 = ~w27188 & ~w27187;
assign w32616 = ~w27208 & w27198;
assign w32617 = w27208 & ~w27198;
assign w32618 = w27289 & ~w27374;
assign w32619 = ~w27453 & ~w32254;
assign w32620 = ~w27453 & ~w27430;
assign w32621 = w27453 & w32254;
assign w32622 = w27453 & w27430;
assign w32623 = ~w27318 & w27572;
assign w32624 = w27471 & ~w27470;
assign w32625 = ~w4070 & w27688;
assign w32626 = w27585 & w27825;
assign w32627 = ~w27585 & ~w27825;
assign w32628 = w27847 & w28060;
assign w32629 = ~w28082 & ~w27864;
assign w32630 = ~w29480 & ~w29477;
assign w32631 = ~w30776 & ~w30775;
assign w32632 = w30889 & w31368;
assign w32633 = ~w31440 & w31443;
assign w32634 = w25141 & w24987;
assign w32635 = ~w7961 & ~w24783;
assign w32636 = ~w86 & ~w85;
assign w32637 = w78 & w92;
assign w32638 = ~w183 & ~w188;
assign w32639 = ~w206 & ~w205;
assign w32640 = w204 & ~w142;
assign w32641 = ~a_23 & ~w510;
assign w32642 = w511 & ~w501;
assign w32643 = w526 & ~w252;
assign w32644 = w847 & w851;
assign w32645 = w898 & ~w97;
assign w32646 = a_26 & ~w1183;
assign w32647 = ~w518 & w122;
assign w32648 = w521 & ~w264;
assign w32649 = ~w1322 & w668;
assign w32650 = ~w188 & ~w590;
assign w32651 = w1463 & w1474;
assign w32652 = ~w206 & ~w34;
assign w32653 = a_26 & w21;
assign w32654 = w894 & w2032;
assign w32655 = ~w834 & ~w420;
assign w32656 = w2200 & ~w559;
assign w32657 = ~w732 & ~w626;
assign w32658 = ~w3198 & ~w3197;
assign w32659 = w3304 & w2215;
assign w32660 = ~w3327 & w3272;
assign w32661 = ~w3327 & w31570;
assign w32662 = w3341 & w3362;
assign w32663 = w3441 & w3454;
assign w32664 = w3416 & w3455;
assign w32665 = ~w3326 & ~w3268;
assign w32666 = ~w3541 & ~w3548;
assign w32667 = ~w3553 & ~w3554;
assign w32668 = w3558 & w3554;
assign w32669 = w3558 & ~w32667;
assign w32670 = ~w2394 & w3618;
assign w32671 = ~w32670 & w3626;
assign w32672 = w2238 & ~w3626;
assign w32673 = w2238 & ~w32671;
assign w32674 = w3717 & w32672;
assign w32675 = w3717 & w32673;
assign w32676 = ~w3713 & ~w2006;
assign w32677 = ~w3722 & ~w32674;
assign w32678 = ~w3722 & ~w32675;
assign w32679 = ~w3725 & ~w2007;
assign w32680 = w1917 & ~w2007;
assign w32681 = w1917 & w32679;
assign w32682 = w3730 & ~w32680;
assign w32683 = w3730 & ~w32681;
assign w32684 = ~w1809 & ~w32682;
assign w32685 = ~w1809 & ~w32683;
assign w32686 = ~w896 & ~w369;
assign w32687 = w3816 & ~w32684;
assign w32688 = w3816 & ~w32685;
assign w32689 = w3819 & ~w32687;
assign w32690 = w3819 & ~w32688;
assign w32691 = w3821 & w32689;
assign w32692 = w3821 & w32690;
assign w32693 = ~w1630 & ~w3823;
assign w32694 = ~w32693 & w3827;
assign w32695 = w1479 & w3831;
assign w32696 = ~w1479 & ~w3831;
assign w32697 = ~w1478 & w3836;
assign w32698 = ~w1190 & ~w1188;
assign w32699 = w3840 & w1188;
assign w32700 = w3840 & ~w32698;
assign w32701 = ~w933 & ~w32699;
assign w32702 = ~w933 & ~w32700;
assign w32703 = w1354 & w3848;
assign w32704 = w1278 & w528;
assign w32705 = w3860 & a_29;
assign w32706 = ~w3860 & ~a_29;
assign w32707 = ~w3863 & w32701;
assign w32708 = ~w3863 & w32702;
assign w32709 = w3863 & ~w32701;
assign w32710 = w3863 & ~w32702;
assign w32711 = w3896 & ~w3891;
assign w32712 = w3902 & ~w16;
assign w32713 = ~w3905 & w1327;
assign w32714 = ~w1322 & w1399;
assign w32715 = w3923 & ~w265;
assign w32716 = w3905 & ~w3934;
assign w32717 = ~w3829 & ~w3831;
assign w32718 = ~w3829 & ~w32695;
assign w32719 = w3939 & ~w32717;
assign w32720 = w3939 & ~w32718;
assign w32721 = ~w3937 & ~w32719;
assign w32722 = ~w3937 & ~w32720;
assign w32723 = ~w3936 & ~w32721;
assign w32724 = ~w3936 & ~w32722;
assign w32725 = w3936 & w32721;
assign w32726 = w3936 & w32722;
assign w32727 = ~w1478 & w3944;
assign w32728 = w3909 & w3876;
assign w32729 = ~w3957 & ~a_29;
assign w32730 = ~w3905 & w668;
assign w32731 = ~w3939 & w32717;
assign w32732 = ~w3939 & w32718;
assign w32733 = ~w3962 & ~w3961;
assign w32734 = w3966 & w3959;
assign w32735 = ~w3840 & ~w1188;
assign w32736 = ~w3840 & w32698;
assign w32737 = ~w3966 & ~w3959;
assign w32738 = w1927 & w3998;
assign w32739 = ~w1561 & w1399;
assign w32740 = ~w1522 & w1327;
assign w32741 = w1630 & w4038;
assign w32742 = ~w1630 & ~w4038;
assign w32743 = ~w1478 & w4043;
assign w32744 = ~w4034 & ~w4032;
assign w32745 = w4047 & w4032;
assign w32746 = w4047 & ~w32744;
assign w32747 = ~w4047 & ~w4032;
assign w32748 = ~w4047 & w32744;
assign w32749 = ~w1522 & w1399;
assign w32750 = w4054 & ~w4038;
assign w32751 = w4054 & ~w32741;
assign w32752 = ~w1478 & w4058;
assign w32753 = w4059 & ~w4048;
assign w32754 = ~w1190 & w3836;
assign w32755 = ~w1190 & w32697;
assign w32756 = ~w3905 & w3957;
assign w32757 = w3906 & ~w32723;
assign w32758 = w3906 & ~w32724;
assign w32759 = ~w3958 & ~w32757;
assign w32760 = ~w3958 & ~w32758;
assign w32761 = w3934 & ~w32723;
assign w32762 = w3934 & ~w32724;
assign w32763 = ~w4070 & w4074;
assign w32764 = a_29 & ~w4074;
assign w32765 = a_29 & ~w32763;
assign w32766 = ~w4078 & ~w4064;
assign w32767 = a_23 & ~w4212;
assign w32768 = ~w1522 & w668;
assign w32769 = ~w1561 & w1327;
assign w32770 = ~w3821 & ~w32689;
assign w32771 = ~w3821 & ~w32690;
assign w32772 = ~w4221 & ~w4222;
assign w32773 = ~w4226 & w4219;
assign w32774 = ~w4217 & ~w4219;
assign w32775 = ~w4217 & ~w32773;
assign w32776 = ~w4034 & w4043;
assign w32777 = ~w4034 & w32743;
assign w32778 = ~w4229 & ~w4228;
assign w32779 = w4229 & w4228;
assign w32780 = ~w1561 & w668;
assign w32781 = ~w1794 & w1399;
assign w32782 = ~w3815 & w32689;
assign w32783 = ~w3815 & w32690;
assign w32784 = w4239 & w32684;
assign w32785 = w4239 & w32685;
assign w32786 = w4242 & ~w32784;
assign w32787 = w4242 & ~w32785;
assign w32788 = ~w4236 & ~w4237;
assign w32789 = ~w4246 & w4234;
assign w32790 = ~w125 & ~w279;
assign w32791 = a_20 & ~w4416;
assign w32792 = ~w1887 & w1399;
assign w32793 = ~w1794 & w668;
assign w32794 = ~w1915 & ~w32680;
assign w32795 = ~w1915 & ~w32681;
assign w32796 = ~w3729 & ~w32794;
assign w32797 = ~w3729 & ~w32795;
assign w32798 = ~w1478 & w4430;
assign w32799 = ~w4423 & ~w4421;
assign w32800 = w4434 & w4421;
assign w32801 = w4434 & ~w32799;
assign w32802 = ~w4289 & ~w32800;
assign w32803 = ~w4289 & ~w32801;
assign w32804 = w4246 & ~w4234;
assign w32805 = w4436 & ~w4247;
assign w32806 = w4226 & ~w4219;
assign w32807 = ~w1322 & w4446;
assign w32808 = ~w4070 & w4451;
assign w32809 = a_29 & ~w4451;
assign w32810 = a_29 & ~w32808;
assign w32811 = ~w4455 & ~w4443;
assign w32812 = ~w4232 & ~w4230;
assign w32813 = w4460 & w4230;
assign w32814 = w4460 & ~w32812;
assign w32815 = ~w4460 & ~w4230;
assign w32816 = ~w4460 & w32812;
assign w32817 = ~w3905 & w4068;
assign w32818 = ~w1322 & w3957;
assign w32819 = ~w4070 & w4468;
assign w32820 = ~a_29 & w4468;
assign w32821 = ~a_29 & w32819;
assign w32822 = ~w4472 & ~w4461;
assign w32823 = ~w1322 & w4068;
assign w32824 = ~w3905 & w4446;
assign w32825 = ~w4070 & w4482;
assign w32826 = ~a_29 & w4482;
assign w32827 = ~a_29 & w32825;
assign w32828 = w1226 & ~w32757;
assign w32829 = w1226 & ~w32758;
assign w32830 = w518 & ~w32828;
assign w32831 = w518 & ~w32829;
assign w32832 = ~w3958 & ~a_26;
assign w32833 = w3958 & a_26;
assign w32834 = ~w4485 & ~w4489;
assign w32835 = w4485 & w4489;
assign w32836 = ~w4494 & ~w4490;
assign w32837 = ~w4434 & ~w4421;
assign w32838 = ~w4434 & w32799;
assign w32839 = ~w1794 & w1327;
assign w32840 = ~w4239 & ~w32684;
assign w32841 = ~w4239 & ~w32685;
assign w32842 = ~w1478 & w4510;
assign w32843 = ~w3646 & w1399;
assign w32844 = ~w1985 & w1327;
assign w32845 = ~w1887 & w668;
assign w32846 = ~w1478 & w4580;
assign w32847 = ~w4573 & ~w4571;
assign w32848 = w4584 & w4571;
assign w32849 = w4584 & ~w32847;
assign w32850 = ~w4584 & ~w4571;
assign w32851 = ~w4584 & w32847;
assign w32852 = ~w1887 & w1327;
assign w32853 = ~w1985 & w1399;
assign w32854 = ~w1917 & w2007;
assign w32855 = ~w1917 & ~w32679;
assign w32856 = ~w1478 & w4594;
assign w32857 = w4595 & ~w4585;
assign w32858 = ~w4423 & w4430;
assign w32859 = ~w4423 & w32798;
assign w32860 = ~w1522 & w4446;
assign w32861 = ~w1561 & w4068;
assign w32862 = ~w4604 & ~w4605;
assign w32863 = w4607 & a_29;
assign w32864 = ~w4607 & ~a_29;
assign w32865 = w4610 & ~w4600;
assign w32866 = ~w4614 & ~w4512;
assign w32867 = w4617 & w4512;
assign w32868 = w4617 & ~w32866;
assign w32869 = ~w4617 & ~w4512;
assign w32870 = ~w4617 & w32866;
assign w32871 = ~w1522 & w3957;
assign w32872 = ~w4070 & w4625;
assign w32873 = ~a_29 & w4625;
assign w32874 = ~a_29 & w32872;
assign w32875 = ~w4629 & ~w4618;
assign w32876 = ~w3905 & ~w518;
assign w32877 = ~w1226 & w4640;
assign w32878 = ~a_26 & ~w4640;
assign w32879 = ~a_26 & ~w32877;
assign w32880 = w4644 & ~w4634;
assign w32881 = ~w1561 & w3957;
assign w32882 = ~w1522 & w4068;
assign w32883 = ~w4070 & w4657;
assign w32884 = ~a_29 & ~w4657;
assign w32885 = ~a_29 & ~w32883;
assign w32886 = ~w1322 & w4638;
assign w32887 = ~w3905 & w4666;
assign w32888 = ~w1226 & w4670;
assign w32889 = a_26 & ~w4670;
assign w32890 = a_26 & ~w32888;
assign w32891 = ~w4674 & ~w4662;
assign w32892 = ~w3905 & w4638;
assign w32893 = ~w1322 & ~w518;
assign w32894 = ~w1226 & w4681;
assign w32895 = ~a_26 & w4681;
assign w32896 = ~a_26 & w32894;
assign w32897 = ~w4688 & ~w4686;
assign w32898 = ~w1561 & w4446;
assign w32899 = ~w1794 & w3957;
assign w32900 = ~w4070 & w4704;
assign w32901 = ~a_29 & w4704;
assign w32902 = ~a_29 & w32900;
assign w32903 = a_17 & ~w4773;
assign w32904 = ~w3646 & w1327;
assign w32905 = ~w3699 & w1399;
assign w32906 = ~w1985 & w668;
assign w32907 = ~w3619 & ~w3718;
assign w32908 = ~w32670 & w4787;
assign w32909 = ~w4786 & ~w4787;
assign w32910 = ~w4786 & ~w32908;
assign w32911 = ~w3716 & ~w3720;
assign w32912 = ~w4785 & ~w3720;
assign w32913 = ~w4785 & w32911;
assign w32914 = w4791 & w1478;
assign w32915 = ~w4794 & w4780;
assign w32916 = ~w4778 & ~w4780;
assign w32917 = ~w4778 & ~w32915;
assign w32918 = ~w4573 & w4580;
assign w32919 = ~w4573 & w32846;
assign w32920 = ~w3646 & w668;
assign w32921 = ~w3699 & w1327;
assign w32922 = ~w2215 & w1399;
assign w32923 = ~w3714 & w32909;
assign w32924 = ~w3714 & w32910;
assign w32925 = w4807 & ~w32923;
assign w32926 = w4807 & ~w32924;
assign w32927 = ~w4807 & w32923;
assign w32928 = ~w4807 & w32924;
assign w32929 = ~w1478 & w4812;
assign w32930 = a_14 & ~w4947;
assign w32931 = ~w2215 & w668;
assign w32932 = ~w32670 & w3625;
assign w32933 = w2149 & w4959;
assign w32934 = ~w2149 & ~w4959;
assign w32935 = ~w1478 & w4964;
assign w32936 = ~w4954 & ~w4952;
assign w32937 = w4968 & w4952;
assign w32938 = w4968 & ~w32936;
assign w32939 = ~w4846 & ~w32937;
assign w32940 = ~w4846 & ~w32938;
assign w32941 = ~w4803 & w4812;
assign w32942 = ~w4803 & w32929;
assign w32943 = w4794 & ~w4780;
assign w32944 = ~w1887 & w3957;
assign w32945 = ~w1794 & w4446;
assign w32946 = ~w4070 & w4984;
assign w32947 = ~a_29 & w4984;
assign w32948 = ~a_29 & w32946;
assign w32949 = ~w4988 & ~w4977;
assign w32950 = ~w4801 & ~w4799;
assign w32951 = ~w4994 & ~w4709;
assign w32952 = ~w1322 & w4666;
assign w32953 = ~w1226 & w5006;
assign w32954 = ~a_26 & w5006;
assign w32955 = ~a_26 & w32953;
assign w32956 = ~w5010 & ~w4999;
assign w32957 = w5017 & ~w32757;
assign w32958 = w5017 & ~w32758;
assign w32959 = ~w5016 & ~w32957;
assign w32960 = ~w5016 & ~w32958;
assign w32961 = ~w3958 & ~a_23;
assign w32962 = w3958 & a_23;
assign w32963 = ~w5024 & ~w5022;
assign w32964 = ~w1522 & ~w518;
assign w32965 = ~w1226 & w5040;
assign w32966 = ~a_26 & w5040;
assign w32967 = ~a_26 & w32965;
assign w32968 = ~w1794 & w4068;
assign w32969 = ~w5049 & ~w5050;
assign w32970 = ~w5052 & a_29;
assign w32971 = w5052 & ~a_29;
assign w32972 = ~w1522 & w4638;
assign w32973 = ~w1561 & ~w518;
assign w32974 = ~w1226 & w5063;
assign w32975 = ~a_26 & w5063;
assign w32976 = ~a_26 & w32974;
assign w32977 = ~w5067 & ~w5056;
assign w32978 = ~w3905 & w5016;
assign w32979 = ~w5017 & w5082;
assign w32980 = ~a_23 & ~w5082;
assign w32981 = ~a_23 & ~w32979;
assign w32982 = w5086 & ~w5076;
assign w32983 = ~w4968 & ~w4952;
assign w32984 = ~w4968 & w32936;
assign w32985 = ~w3699 & w668;
assign w32986 = ~w2215 & w1327;
assign w32987 = w5100 & ~w32672;
assign w32988 = w5100 & ~w32673;
assign w32989 = ~w5100 & w32672;
assign w32990 = ~w5100 & w32673;
assign w32991 = ~w5097 & ~w5099;
assign w32992 = ~w3646 & w3957;
assign w32993 = ~w1985 & w4068;
assign w32994 = ~w1887 & w4446;
assign w32995 = ~w4070 & w5114;
assign w32996 = ~a_29 & w5114;
assign w32997 = ~a_29 & w32995;
assign w32998 = ~w5118 & ~w5107;
assign w32999 = ~w1887 & w4068;
assign w33000 = ~w1985 & w3957;
assign w33001 = ~w4070 & w5130;
assign w33002 = ~a_29 & w5130;
assign w33003 = ~a_29 & w33001;
assign w33004 = w5134 & ~w5123;
assign w33005 = ~w1522 & w4666;
assign w33006 = ~w1561 & w4638;
assign w33007 = ~w5141 & ~w5142;
assign w33008 = ~w5144 & a_26;
assign w33009 = w5144 & ~a_26;
assign w33010 = ~w1794 & ~w518;
assign w33011 = ~w1561 & w4666;
assign w33012 = ~w1226 & w5157;
assign w33013 = ~a_26 & w5157;
assign w33014 = ~a_26 & w33012;
assign w33015 = w2394 & w5223;
assign w33016 = ~w3616 & ~w5223;
assign w33017 = ~w3616 & ~w33015;
assign w33018 = w5222 & ~w33016;
assign w33019 = w5222 & ~w33017;
assign w33020 = ~w5222 & w33016;
assign w33021 = ~w5222 & w33017;
assign w33022 = ~w1478 & w5229;
assign w33023 = ~w5218 & ~w5216;
assign w33024 = w5233 & w5216;
assign w33025 = w5233 & ~w33023;
assign w33026 = ~w5233 & ~w5216;
assign w33027 = ~w5233 & w33023;
assign w33028 = w5240 & ~w33018;
assign w33029 = w5240 & ~w33019;
assign w33030 = ~w1478 & w5244;
assign w33031 = w5245 & ~w5234;
assign w33032 = ~w4954 & w4964;
assign w33033 = ~w4954 & w32935;
assign w33034 = ~w3646 & w4068;
assign w33035 = ~w1985 & w4446;
assign w33036 = ~w3699 & w3957;
assign w33037 = w4791 & w4070;
assign w33038 = ~w5258 & a_29;
assign w33039 = w5258 & ~a_29;
assign w33040 = ~w5261 & ~w5250;
assign w33041 = ~w1794 & w4638;
assign w33042 = ~w5270 & ~w5271;
assign w33043 = ~w5273 & a_26;
assign w33044 = w5273 & ~a_26;
assign w33045 = ~w5276 & ~w5266;
assign w33046 = w5278 & ~w5162;
assign w33047 = ~w1322 & w5286;
assign w33048 = ~w5017 & w5289;
assign w33049 = ~a_23 & w5289;
assign w33050 = ~a_23 & w33048;
assign w33051 = w5293 & ~w5283;
assign w33052 = w5309 & ~w32757;
assign w33053 = w5309 & ~w32758;
assign w33054 = ~w5308 & ~w33052;
assign w33055 = ~w5308 & ~w33053;
assign w33056 = ~w3958 & ~a_20;
assign w33057 = w3958 & a_20;
assign w33058 = w5147 & ~w5137;
assign w33059 = ~w3905 & w5286;
assign w33060 = ~w1322 & w5080;
assign w33061 = ~w5017 & w5327;
assign w33062 = ~a_23 & w5327;
assign w33063 = ~a_23 & w33061;
assign w33064 = ~w5334 & ~w5314;
assign w33065 = ~w5331 & ~w5320;
assign w33066 = ~w3905 & w5080;
assign w33067 = ~w1322 & w5016;
assign w33068 = ~w5017 & w5344;
assign w33069 = ~a_23 & w5344;
assign w33070 = ~a_23 & w33068;
assign w33071 = ~w3646 & ~w518;
assign w33072 = ~w1985 & w4638;
assign w33073 = ~w1887 & w4666;
assign w33074 = ~w1226 & w5360;
assign w33075 = ~a_26 & w5360;
assign w33076 = ~a_26 & w33074;
assign w33077 = a_11 & ~w5451;
assign w33078 = ~w2394 & ~w5223;
assign w33079 = ~w1478 & w5465;
assign w33080 = ~w5458 & ~w5456;
assign w33081 = ~w5218 & w5229;
assign w33082 = ~w5218 & w33022;
assign w33083 = ~w3515 & w1399;
assign w33084 = w3553 & w5479;
assign w33085 = ~w33084 & w5481;
assign w33086 = ~w1478 & w5485;
assign w33087 = a_8 & ~w5637;
assign w33088 = ~w3515 & w668;
assign w33089 = ~w3545 & w3552;
assign w33090 = w3476 & w5648;
assign w33091 = ~w3476 & ~w5648;
assign w33092 = ~w1478 & w5654;
assign w33093 = ~w5644 & ~w5642;
assign w33094 = w5658 & w5642;
assign w33095 = w5658 & ~w33093;
assign w33096 = ~w5511 & ~w33094;
assign w33097 = ~w5511 & ~w33095;
assign w33098 = ~w5475 & w5485;
assign w33099 = ~w5475 & w33086;
assign w33100 = w5660 & ~w5487;
assign w33101 = ~w5458 & w5465;
assign w33102 = ~w5458 & w33079;
assign w33103 = ~w2215 & w4446;
assign w33104 = ~w4070 & w5674;
assign w33105 = ~a_29 & w5674;
assign w33106 = ~a_29 & w33104;
assign w33107 = ~w5678 & ~w5667;
assign w33108 = ~w2215 & w4068;
assign w33109 = ~w3699 & w4446;
assign w33110 = ~w5684 & ~w5686;
assign w33111 = ~w5688 & a_29;
assign w33112 = w5688 & ~a_29;
assign w33113 = ~w5658 & ~w5642;
assign w33114 = ~w5658 & w33093;
assign w33115 = ~w3515 & w1327;
assign w33116 = ~w3553 & ~w5479;
assign w33117 = ~w1478 & w5708;
assign w33118 = ~w4070 & w5717;
assign w33119 = ~a_29 & ~w5717;
assign w33120 = ~a_29 & ~w33118;
assign w33121 = w5721 & ~w5710;
assign w33122 = ~w4070 & w5733;
assign w33123 = ~a_29 & w5733;
assign w33124 = ~a_29 & w33122;
assign w33125 = w5737 & ~w5726;
assign w33126 = ~w3646 & w4638;
assign w33127 = ~w1985 & w4666;
assign w33128 = ~w3699 & ~w518;
assign w33129 = w4791 & w1226;
assign w33130 = ~w5746 & a_26;
assign w33131 = w5746 & ~a_26;
assign w33132 = w5749 & ~w5740;
assign w33133 = ~w1561 & w5016;
assign w33134 = ~w1794 & w5080;
assign w33135 = ~w5758 & ~w5759;
assign w33136 = w5761 & a_23;
assign w33137 = ~w5761 & ~a_23;
assign w33138 = w5764 & ~w5754;
assign w33139 = ~w5364 & ~w5692;
assign w33140 = ~w5473 & ~w5471;
assign w33141 = ~w3646 & w4446;
assign w33142 = ~w3699 & w4068;
assign w33143 = ~w2215 & w3957;
assign w33144 = ~w4070 & w5775;
assign w33145 = ~a_29 & w5775;
assign w33146 = ~a_29 & w33144;
assign w33147 = ~w1887 & w4638;
assign w33148 = ~w1985 & ~w518;
assign w33149 = ~w1226 & w5790;
assign w33150 = ~a_26 & w5790;
assign w33151 = ~a_26 & w33149;
assign w33152 = ~w1794 & w5016;
assign w33153 = ~w1561 & w5286;
assign w33154 = ~w5017 & w5805;
assign w33155 = ~a_23 & w5805;
assign w33156 = ~a_23 & w33154;
assign w33157 = ~w1522 & w5308;
assign w33158 = ~w5309 & w5822;
assign w33159 = ~a_20 & ~w5822;
assign w33160 = ~a_20 & ~w33158;
assign w33161 = ~w3646 & w4666;
assign w33162 = ~w3699 & w4638;
assign w33163 = ~w2215 & ~w518;
assign w33164 = ~w1226 & w5838;
assign w33165 = ~a_26 & w5838;
assign w33166 = ~a_26 & w33164;
assign w33167 = a_5 & ~w5888;
assign w33168 = ~w3206 & w1327;
assign w33169 = ~w5900 & ~w3272;
assign w33170 = ~w5900 & ~w31570;
assign w33171 = w5900 & w3272;
assign w33172 = w5900 & w31570;
assign w33173 = ~w1478 & w5905;
assign w33174 = ~w5895 & ~w5893;
assign w33175 = w5909 & w5893;
assign w33176 = w5909 & ~w33174;
assign w33177 = ~w5871 & ~w33175;
assign w33178 = ~w5871 & ~w33176;
assign w33179 = ~w5920 & ~w5921;
assign w33180 = ~w1478 & w5925;
assign w33181 = w5926 & ~w5914;
assign w33182 = ~w5644 & w5654;
assign w33183 = ~w5644 & w33092;
assign w33184 = ~w4070 & w5938;
assign w33185 = ~a_29 & w5938;
assign w33186 = ~a_29 & w33184;
assign w33187 = ~w5942 & ~w5931;
assign w33188 = ~w3699 & w4666;
assign w33189 = ~w2215 & w4638;
assign w33190 = ~w1226 & w5954;
assign w33191 = ~a_26 & w5954;
assign w33192 = ~a_26 & w33190;
assign w33193 = ~w5958 & ~w5947;
assign w33194 = w5960 & ~w5843;
assign w33195 = ~w1887 & w5016;
assign w33196 = ~w1561 & w5080;
assign w33197 = ~w1794 & w5286;
assign w33198 = ~w5017 & w5972;
assign w33199 = ~a_23 & ~w5972;
assign w33200 = ~a_23 & ~w33198;
assign w33201 = ~w5976 & ~w5965;
assign w33202 = ~w1561 & w5308;
assign w33203 = ~w1522 & w5818;
assign w33204 = ~w5309 & w5984;
assign w33205 = ~a_20 & w5984;
assign w33206 = ~a_20 & w33204;
assign w33207 = ~w5988 & ~w5979;
assign w33208 = ~w1322 & w5816;
assign w33209 = ~w5309 & w6001;
assign w33210 = ~a_20 & w6001;
assign w33211 = ~a_20 & w33209;
assign w33212 = ~w1522 & w5286;
assign w33213 = ~w6007 & ~w6008;
assign w33214 = ~w6010 & a_23;
assign w33215 = w6010 & ~a_23;
assign w33216 = ~w1887 & ~w518;
assign w33217 = ~w1794 & w4666;
assign w33218 = ~w1226 & w6024;
assign w33219 = ~a_26 & w6024;
assign w33220 = ~a_26 & w33218;
assign w33221 = ~w3905 & w6059;
assign w33222 = ~w6063 & w6064;
assign w33223 = ~a_17 & w6064;
assign w33224 = ~a_17 & w33222;
assign w33225 = ~w1887 & w5080;
assign w33226 = ~w1985 & w5016;
assign w33227 = ~w5017 & w6080;
assign w33228 = ~a_23 & ~w6080;
assign w33229 = ~a_23 & ~w33227;
assign w33230 = ~w3515 & w3957;
assign w33231 = ~w4070 & w6094;
assign w33232 = ~a_29 & w6094;
assign w33233 = ~a_29 & w33231;
assign w33234 = ~w5909 & ~w5893;
assign w33235 = ~w5909 & w33174;
assign w33236 = ~w3206 & w1399;
assign w33237 = w3544 & w6105;
assign w33238 = ~w3544 & ~w6105;
assign w33239 = ~w1478 & w6110;
assign w33240 = ~w6185 & ~w32435;
assign w33241 = ~w6185 & ~w32436;
assign w33242 = w6202 & ~w33240;
assign w33243 = w6202 & ~w33241;
assign w33244 = w6154 & w6205;
assign w33245 = ~w6137 & ~w6205;
assign w33246 = ~w6137 & ~w33244;
assign w33247 = w6208 & ~w33245;
assign w33248 = w6208 & ~w33246;
assign w33249 = ~w6208 & w33245;
assign w33250 = ~w6208 & w33246;
assign w33251 = ~w3206 & w668;
assign w33252 = ~w3273 & w1478;
assign w33253 = w6226 & ~w6209;
assign w33254 = ~w5895 & w5905;
assign w33255 = ~w5895 & w33173;
assign w33256 = ~w3515 & w4446;
assign w33257 = ~w4070 & w6238;
assign w33258 = ~a_29 & ~w6238;
assign w33259 = ~a_29 & ~w33257;
assign w33260 = w6242 & ~w6231;
assign w33261 = ~w6114 & ~w6112;
assign w33262 = ~w2215 & w4666;
assign w33263 = ~w1226 & w6260;
assign w33264 = ~a_26 & w6260;
assign w33265 = ~a_26 & w33263;
assign w33266 = w6264 & ~w6253;
assign w33267 = ~w3646 & w5016;
assign w33268 = ~w1985 & w5080;
assign w33269 = ~w1887 & w5286;
assign w33270 = ~w5017 & w6272;
assign w33271 = ~a_23 & w6272;
assign w33272 = ~a_23 & w33270;
assign w33273 = ~w6276 & ~w6267;
assign w33274 = w6280 & ~w6085;
assign w33275 = ~w1522 & w5816;
assign w33276 = ~w1561 & w5818;
assign w33277 = ~w6289 & ~w6290;
assign w33278 = ~w6292 & a_20;
assign w33279 = w6292 & ~a_20;
assign w33280 = ~w6295 & ~w6285;
assign w33281 = ~w3905 & w6304;
assign w33282 = ~w1322 & w6061;
assign w33283 = ~w6063 & w6308;
assign w33284 = ~a_17 & w6308;
assign w33285 = ~a_17 & w33283;
assign w33286 = ~w6312 & ~w6300;
assign w33287 = ~w3905 & w6061;
assign w33288 = ~w1322 & w6059;
assign w33289 = ~w6063 & w6319;
assign w33290 = ~a_17 & w6319;
assign w33291 = ~a_17 & w33289;
assign w33292 = ~w6326 & ~w6324;
assign w33293 = ~w1794 & w5308;
assign w33294 = ~w1561 & w5816;
assign w33295 = ~w5309 & w6338;
assign w33296 = ~a_20 & w6338;
assign w33297 = ~a_20 & w33295;
assign w33298 = ~w1226 & w6354;
assign w33299 = ~a_26 & w6354;
assign w33300 = ~a_26 & w33298;
assign w33301 = ~w3515 & w4068;
assign w33302 = ~w4070 & w6366;
assign w33303 = ~a_29 & ~w6366;
assign w33304 = ~a_29 & ~w33302;
assign w33305 = ~w1226 & w6376;
assign w33306 = ~a_26 & w6376;
assign w33307 = ~a_26 & w33305;
assign w33308 = ~w6380 & ~w6371;
assign w33309 = ~w3646 & w5080;
assign w33310 = ~w1985 & w5286;
assign w33311 = ~w3699 & w5016;
assign w33312 = w4791 & w5017;
assign w33313 = ~w6397 & a_23;
assign w33314 = w6397 & ~a_23;
assign w33315 = w6400 & ~w6389;
assign w33316 = ~w1794 & w5818;
assign w33317 = ~w6405 & ~w6406;
assign w33318 = ~w6408 & a_20;
assign w33319 = w6408 & ~a_20;
assign w33320 = ~w6411 & ~w6403;
assign w33321 = w6415 & ~w6343;
assign w33322 = ~w1322 & w6304;
assign w33323 = ~w6063 & w6429;
assign w33324 = ~a_17 & w6429;
assign w33325 = ~a_17 & w33323;
assign w33326 = w6433 & ~w6422;
assign w33327 = w6447 & ~w32757;
assign w33328 = w6447 & ~w32758;
assign w33329 = ~w6446 & ~w33327;
assign w33330 = ~w6446 & ~w33328;
assign w33331 = ~w3958 & ~a_14;
assign w33332 = w3958 & a_14;
assign w33333 = ~w6456 & ~w6452;
assign w33334 = ~w3646 & w5286;
assign w33335 = ~w2215 & w5016;
assign w33336 = ~w3699 & w5080;
assign w33337 = ~w5017 & w6470;
assign w33338 = ~a_23 & ~w6470;
assign w33339 = ~a_23 & ~w33337;
assign w33340 = ~w6154 & ~w6205;
assign w33341 = ~w1478 & w6493;
assign w33342 = ~w6202 & w33240;
assign w33343 = ~w6202 & w33241;
assign w33344 = ~w1478 & w6507;
assign w33345 = ~w1478 & w6549;
assign w33346 = ~w2736 & w668;
assign w33347 = ~w46 & ~w62;
assign w33348 = ~w2465 & w1399;
assign w33349 = ~w2736 & w1327;
assign w33350 = w6723 & ~w6720;
assign w33351 = ~w6723 & w6720;
assign w33352 = ~w2736 & w1399;
assign w33353 = ~w6773 & ~w6786;
assign w33354 = ~w6773 & ~w32437;
assign w33355 = w6773 & w6786;
assign w33356 = w6773 & w32437;
assign w33357 = ~w6740 & w6789;
assign w33358 = ~w6539 & ~w6549;
assign w33359 = ~w6539 & ~w33345;
assign w33360 = ~w6187 & w6199;
assign w33361 = ~w6187 & w31571;
assign w33362 = ~w6794 & w6551;
assign w33363 = ~w6794 & ~w32438;
assign w33364 = w6794 & ~w6551;
assign w33365 = w6794 & w32438;
assign w33366 = ~w3273 & w4070;
assign w33367 = ~w6802 & a_29;
assign w33368 = w6802 & ~a_29;
assign w33369 = ~w6795 & w6511;
assign w33370 = w6509 & w6809;
assign w33371 = w6495 & w6812;
assign w33372 = ~w4070 & w6818;
assign w33373 = ~a_29 & w6818;
assign w33374 = ~a_29 & w33372;
assign w33375 = ~w6495 & ~w6812;
assign w33376 = ~w6822 & ~w6813;
assign w33377 = ~w1226 & w6832;
assign w33378 = ~a_26 & w6832;
assign w33379 = ~a_26 & w33377;
assign w33380 = w6836 & ~w6827;
assign w33381 = ~w3699 & w5286;
assign w33382 = ~w2215 & w5080;
assign w33383 = ~w6842 & ~w6844;
assign w33384 = ~w6846 & a_23;
assign w33385 = w6846 & ~a_23;
assign w33386 = w6849 & ~w6841;
assign w33387 = ~w1887 & w5308;
assign w33388 = ~w1794 & w5816;
assign w33389 = ~w5309 & w6863;
assign w33390 = ~a_20 & w6863;
assign w33391 = ~a_20 & w33389;
assign w33392 = ~w6867 & ~w6858;
assign w33393 = ~w1561 & w6059;
assign w33394 = ~w1522 & w6061;
assign w33395 = ~w6063 & w6881;
assign w33396 = ~a_17 & ~w6881;
assign w33397 = ~a_17 & ~w33395;
assign w33398 = ~w1887 & w5818;
assign w33399 = ~w1985 & w5308;
assign w33400 = ~w5309 & w6895;
assign w33401 = ~a_20 & w6895;
assign w33402 = ~a_20 & w33400;
assign w33403 = ~w3515 & ~w518;
assign w33404 = ~w1226 & w6907;
assign w33405 = ~a_26 & w6907;
assign w33406 = ~a_26 & w33404;
assign w33407 = ~w6509 & ~w6809;
assign w33408 = ~w3206 & w3957;
assign w33409 = ~w4070 & w6922;
assign w33410 = ~a_29 & w6922;
assign w33411 = ~a_29 & w33409;
assign w33412 = ~w3515 & w4638;
assign w33413 = ~w1226 & w6932;
assign w33414 = ~a_26 & w6932;
assign w33415 = ~a_26 & w33413;
assign w33416 = w6936 & ~w6927;
assign w33417 = ~w2215 & w5286;
assign w33418 = ~w5017 & w6948;
assign w33419 = ~a_23 & w6948;
assign w33420 = ~a_23 & w33418;
assign w33421 = w6952 & ~w6943;
assign w33422 = ~w3646 & w5308;
assign w33423 = ~w1985 & w5818;
assign w33424 = ~w1887 & w5816;
assign w33425 = ~w5309 & w6964;
assign w33426 = ~a_20 & w6964;
assign w33427 = ~a_20 & w33425;
assign w33428 = ~w6968 & ~w6959;
assign w33429 = ~w1522 & w6304;
assign w33430 = ~w1561 & w6061;
assign w33431 = ~w6983 & ~w6984;
assign w33432 = w6986 & a_17;
assign w33433 = ~w6986 & ~a_17;
assign w33434 = ~w6989 & ~w6979;
assign w33435 = ~w3905 & w6996;
assign w33436 = ~w1322 & w6998;
assign w33437 = ~w6447 & w7001;
assign w33438 = ~a_14 & w7001;
assign w33439 = ~a_14 & w33437;
assign w33440 = ~w7005 & ~w6992;
assign w33441 = ~w3905 & w6998;
assign w33442 = ~w1322 & w6446;
assign w33443 = ~w6447 & w7012;
assign w33444 = ~a_14 & w7012;
assign w33445 = ~a_14 & w33443;
assign w33446 = w6885 & ~w6874;
assign w33447 = ~w1522 & w6059;
assign w33448 = ~w6063 & w7025;
assign w33449 = ~a_17 & ~w7025;
assign w33450 = ~a_17 & ~w33448;
assign w33451 = ~w7035 & ~w7017;
assign w33452 = w7018 & ~w7030;
assign w33453 = ~w3905 & w6446;
assign w33454 = ~w6447 & w7045;
assign w33455 = ~a_14 & w7045;
assign w33456 = ~a_14 & w33454;
assign w33457 = ~w1794 & w6059;
assign w33458 = ~w1561 & w6304;
assign w33459 = ~w6063 & w7067;
assign w33460 = ~a_17 & w7067;
assign w33461 = ~a_17 & w33459;
assign w33462 = w6795 & ~w6511;
assign w33463 = ~w3206 & w4068;
assign w33464 = ~w4070 & w7079;
assign w33465 = ~a_29 & ~w7079;
assign w33466 = ~a_29 & ~w33464;
assign w33467 = ~w3515 & w4666;
assign w33468 = ~w1226 & w7091;
assign w33469 = ~a_26 & ~w7091;
assign w33470 = ~a_26 & ~w33468;
assign w33471 = w7095 & ~w7084;
assign w33472 = ~w5017 & w7102;
assign w33473 = ~a_23 & ~w7102;
assign w33474 = ~a_23 & ~w33472;
assign w33475 = ~w5017 & w7119;
assign w33476 = ~a_23 & w7119;
assign w33477 = ~a_23 & w33475;
assign w33478 = ~w3646 & w5818;
assign w33479 = ~w1985 & w5816;
assign w33480 = ~w3699 & w5308;
assign w33481 = w4791 & w5309;
assign w33482 = ~w7138 & a_20;
assign w33483 = w7138 & ~a_20;
assign w33484 = w7144 & ~w7142;
assign w33485 = ~w1794 & w6061;
assign w33486 = ~w7150 & ~w7151;
assign w33487 = ~w7153 & a_17;
assign w33488 = w7153 & ~a_17;
assign w33489 = ~w7159 & ~w7157;
assign w33490 = w7163 & ~w7072;
assign w33491 = ~w1322 & w6996;
assign w33492 = ~w6447 & w7173;
assign w33493 = ~a_14 & w7173;
assign w33494 = ~a_14 & w33492;
assign w33495 = ~w7177 & ~w7168;
assign w33496 = w7193 & ~w32757;
assign w33497 = w7193 & ~w32758;
assign w33498 = ~w7192 & ~w33496;
assign w33499 = ~w7192 & ~w33497;
assign w33500 = ~w3958 & ~a_11;
assign w33501 = w3958 & a_11;
assign w33502 = ~w7200 & ~w7198;
assign w33503 = ~w1522 & w6446;
assign w33504 = ~w6447 & w7214;
assign w33505 = ~a_14 & w7214;
assign w33506 = ~a_14 & w33504;
assign w33507 = ~w3646 & w5816;
assign w33508 = ~w2215 & w5308;
assign w33509 = ~w3699 & w5818;
assign w33510 = ~w5309 & w7224;
assign w33511 = ~a_20 & ~w7224;
assign w33512 = ~a_20 & ~w33510;
assign w33513 = ~w2215 & w5818;
assign w33514 = ~w3699 & w5816;
assign w33515 = ~w7229 & ~w7231;
assign w33516 = ~w7233 & a_20;
assign w33517 = w7233 & ~a_20;
assign w33518 = ~w1226 & w7243;
assign w33519 = a_26 & ~w7243;
assign w33520 = a_26 & ~w33518;
assign w33521 = w6740 & ~w6789;
assign w33522 = ~w4070 & w7262;
assign w33523 = a_29 & ~w7262;
assign w33524 = a_29 & ~w33522;
assign w33525 = ~w2736 & w3957;
assign w33526 = ~w7272 & w7269;
assign w33527 = w7272 & a_29;
assign w33528 = ~w7272 & ~a_29;
assign w33529 = ~w2465 & w668;
assign w33530 = ~w2588 & w1327;
assign w33531 = ~w1478 & w7291;
assign w33532 = ~w2736 & w4446;
assign w33533 = ~w2465 & w3957;
assign w33534 = ~w7312 & ~a_29;
assign w33535 = ~w4070 & w7314;
assign w33536 = w7312 & a_29;
assign w33537 = ~w2588 & ~w1477;
assign w33538 = w6604 & w6629;
assign w33539 = ~w7348 & ~a_29;
assign w33540 = ~w7348 & w7269;
assign w33541 = a_29 & ~w7389;
assign w33542 = a_29 & ~w31600;
assign w33543 = ~a_29 & w7389;
assign w33544 = ~a_29 & w31600;
assign w33545 = ~w7392 & ~w7381;
assign w33546 = ~w7402 & ~w7267;
assign w33547 = w7408 & a_29;
assign w33548 = ~w7408 & ~a_29;
assign w33549 = ~w7268 & ~w7410;
assign w33550 = ~w7420 & w7425;
assign w33551 = ~w5017 & w7435;
assign w33552 = ~a_23 & w7435;
assign w33553 = ~a_23 & w33551;
assign w33554 = w7429 & w7236;
assign w33555 = ~w7429 & ~w7236;
assign w33556 = w7441 & ~w7228;
assign w33557 = ~w7441 & w7228;
assign w33558 = ~w1887 & w6059;
assign w33559 = ~w1794 & w6304;
assign w33560 = ~w6063 & w7456;
assign w33561 = ~a_17 & ~w7456;
assign w33562 = ~a_17 & ~w33560;
assign w33563 = w7446 & ~w7460;
assign w33564 = ~w7446 & w7460;
assign w33565 = ~w7465 & ~w7461;
assign w33566 = ~w1561 & w6446;
assign w33567 = ~w1522 & w6998;
assign w33568 = ~w6447 & w7477;
assign w33569 = ~a_14 & w7477;
assign w33570 = ~a_14 & w33568;
assign w33571 = ~w7481 & ~w7470;
assign w33572 = w7483 & ~w7219;
assign w33573 = ~w3905 & w7192;
assign w33574 = ~w7193 & w7491;
assign w33575 = ~a_11 & w7491;
assign w33576 = ~a_11 & w33574;
assign w33577 = ~w7498 & ~w7496;
assign w33578 = ~w7207 & w7058;
assign w33579 = ~w1322 & w7489;
assign w33580 = ~w3905 & w7511;
assign w33581 = ~w7193 & w7515;
assign w33582 = ~a_11 & w7515;
assign w33583 = ~a_11 & w33581;
assign w33584 = ~w1522 & w6996;
assign w33585 = ~w1561 & w6998;
assign w33586 = ~w7523 & ~w7524;
assign w33587 = ~w7526 & a_14;
assign w33588 = w7526 & ~a_14;
assign w33589 = ~w3515 & w5016;
assign w33590 = ~w5017 & w7541;
assign w33591 = ~a_23 & w7541;
assign w33592 = ~a_23 & w33590;
assign w33593 = ~w3206 & ~w518;
assign w33594 = ~w1226 & w7551;
assign w33595 = ~a_26 & w7551;
assign w33596 = ~a_26 & w33594;
assign w33597 = ~w1226 & w7570;
assign w33598 = ~a_26 & w7570;
assign w33599 = ~a_26 & w33597;
assign w33600 = ~w2465 & ~w518;
assign w33601 = ~w7596 & ~a_26;
assign w33602 = ~w1226 & w7598;
assign w33603 = w7596 & a_26;
assign w33604 = ~w2465 & w4638;
assign w33605 = ~w7608 & ~w7609;
assign w33606 = ~w2736 & w4666;
assign w33607 = ~w7637 & ~a_26;
assign w33608 = ~w2736 & ~w518;
assign w33609 = ~w7633 & a_29;
assign w33610 = ~w7674 & ~a_26;
assign w33611 = ~w7674 & w7680;
assign w33612 = w31574 & w1226;
assign w33613 = w7708 & ~w7703;
assign w33614 = w7708 & ~w31616;
assign w33615 = w7727 & a_26;
assign w33616 = ~w7727 & ~a_26;
assign w33617 = ~w4403 & ~w7729;
assign w33618 = ~w7383 & ~w7381;
assign w33619 = ~w3206 & w4666;
assign w33620 = ~w7747 & ~a_26;
assign w33621 = ~w3273 & w4403;
assign w33622 = ~w7747 & w7680;
assign w33623 = w7747 & a_26;
assign w33624 = ~w7398 & ~w7400;
assign w33625 = w7772 & ~w3272;
assign w33626 = w7772 & ~w31570;
assign w33627 = ~w3206 & w4638;
assign w33628 = ~w7768 & w7792;
assign w33629 = ~w7799 & ~w7546;
assign w33630 = ~w2215 & w5816;
assign w33631 = ~w5309 & w7811;
assign w33632 = ~a_20 & w7811;
assign w33633 = ~a_20 & w33631;
assign w33634 = w7815 & ~w7806;
assign w33635 = ~w3646 & w6059;
assign w33636 = ~w1985 & w6061;
assign w33637 = ~w1887 & w6304;
assign w33638 = ~w6063 & w7829;
assign w33639 = ~a_17 & w7829;
assign w33640 = ~a_17 & w33638;
assign w33641 = ~w7833 & ~w7824;
assign w33642 = ~w1887 & w6061;
assign w33643 = ~w1985 & w6059;
assign w33644 = ~w6063 & w7845;
assign w33645 = ~a_17 & w7845;
assign w33646 = ~a_17 & w33644;
assign w33647 = ~w7849 & ~w7838;
assign w33648 = w7851 & ~w7530;
assign w33649 = ~w3905 & w7489;
assign w33650 = ~w1322 & w7192;
assign w33651 = ~w7193 & w7864;
assign w33652 = ~a_11 & w7864;
assign w33653 = ~a_11 & w33651;
assign w33654 = ~w7854 & w7868;
assign w33655 = w7854 & ~w7868;
assign w33656 = ~w7871 & ~w7869;
assign w33657 = ~w1794 & w6446;
assign w33658 = ~w1561 & w6996;
assign w33659 = ~w6447 & w7887;
assign w33660 = ~a_14 & w7887;
assign w33661 = ~a_14 & w33659;
assign w33662 = ~w5309 & w7900;
assign w33663 = ~a_20 & w7900;
assign w33664 = ~a_20 & w33662;
assign w33665 = ~w3206 & w5286;
assign w33666 = ~w3273 & w5017;
assign w33667 = ~w7915 & a_23;
assign w33668 = w7915 & ~a_23;
assign w33669 = ~w7947 & a_26;
assign w33670 = ~w2736 & w5080;
assign w33671 = ~w7955 & ~a_23;
assign w33672 = ~w7955 & w7962;
assign w33673 = ~w2465 & w5080;
assign w33674 = ~w2588 & w5016;
assign w33675 = ~w7972 & ~w7974;
assign w33676 = ~w2465 & w5016;
assign w33677 = w7989 & a_23;
assign w33678 = ~w7989 & ~a_23;
assign w33679 = ~w7961 & ~w7991;
assign w33680 = ~w2736 & w5286;
assign w33681 = w8006 & a_23;
assign w33682 = ~w2736 & w5016;
assign w33683 = w31574 & w5017;
assign w33684 = w8055 & ~w8050;
assign w33685 = w8055 & ~w31631;
assign w33686 = ~w8068 & ~a_23;
assign w33687 = ~w8068 & w7962;
assign w33688 = w8068 & a_23;
assign w33689 = w8099 & a_23;
assign w33690 = ~w8099 & ~a_23;
assign w33691 = ~w7961 & ~w8101;
assign w33692 = ~w3206 & w5080;
assign w33693 = ~w5017 & w8123;
assign w33694 = ~a_23 & w8123;
assign w33695 = ~a_23 & w33693;
assign w33696 = ~w3206 & w5016;
assign w33697 = ~w5017 & w8144;
assign w33698 = a_23 & ~w8144;
assign w33699 = a_23 & ~w33697;
assign w33700 = ~w5017 & w8164;
assign w33701 = ~a_23 & w8164;
assign w33702 = ~a_23 & w33700;
assign w33703 = ~w3515 & w5286;
assign w33704 = ~w5017 & w8184;
assign w33705 = ~a_23 & w8184;
assign w33706 = ~a_23 & w33704;
assign w33707 = ~w3515 & w5080;
assign w33708 = ~w5017 & w8204;
assign w33709 = ~a_23 & ~w8204;
assign w33710 = ~a_23 & ~w33708;
assign w33711 = w8214 & ~w8215;
assign w33712 = ~w3646 & w6061;
assign w33713 = ~w3699 & w6059;
assign w33714 = ~w1985 & w6304;
assign w33715 = w4791 & w6063;
assign w33716 = w8229 & a_17;
assign w33717 = ~w8229 & ~a_17;
assign w33718 = w8232 & ~w8221;
assign w33719 = ~w1794 & w6998;
assign w33720 = ~w8238 & ~w8239;
assign w33721 = ~w8241 & a_14;
assign w33722 = w8241 & ~a_14;
assign w33723 = w7893 & w8244;
assign w33724 = ~w1322 & w7511;
assign w33725 = ~w7193 & w8260;
assign w33726 = ~a_11 & w8260;
assign w33727 = ~a_11 & w33725;
assign w33728 = ~w8264 & ~w8253;
assign w33729 = w8278 & ~w32757;
assign w33730 = w8278 & ~w32758;
assign w33731 = ~w8277 & ~w33729;
assign w33732 = ~w8277 & ~w33730;
assign w33733 = ~w3958 & ~a_8;
assign w33734 = w3958 & a_8;
assign w33735 = ~w8285 & ~w8283;
assign w33736 = ~w3699 & w8295;
assign w33737 = ~w2215 & w8298;
assign w33738 = ~w8296 & ~w8299;
assign w33739 = ~w8301 & a_8;
assign w33740 = w8301 & ~a_8;
assign w33741 = ~w2736 & w5818;
assign w33742 = ~w8307 & ~a_20;
assign w33743 = w8307 & a_20;
assign w33744 = ~w7983 & a_23;
assign w33745 = ~w2465 & w5818;
assign w33746 = ~w2588 & w5308;
assign w33747 = ~w8323 & ~w8325;
assign w33748 = ~w2465 & w5308;
assign w33749 = ~w8343 & a_20;
assign w33750 = w8343 & ~a_20;
assign w33751 = ~w2736 & w5816;
assign w33752 = ~w6063 & w8377;
assign w33753 = ~a_17 & ~w8377;
assign w33754 = ~a_17 & ~w33752;
assign w33755 = ~w2736 & w6061;
assign w33756 = ~w8387 & ~a_17;
assign w33757 = w8387 & a_17;
assign w33758 = ~w8334 & a_20;
assign w33759 = ~w2465 & w6061;
assign w33760 = ~w2588 & w6059;
assign w33761 = ~w8403 & ~w8405;
assign w33762 = ~w2465 & w6059;
assign w33763 = ~w8423 & a_17;
assign w33764 = w8423 & ~a_17;
assign w33765 = ~w2736 & w6304;
assign w33766 = ~w2736 & w6059;
assign w33767 = a_17 & ~w8456;
assign w33768 = a_17 & ~w31655;
assign w33769 = ~a_17 & w8456;
assign w33770 = ~a_17 & w31655;
assign w33771 = ~w3206 & w6998;
assign w33772 = ~w6447 & w8496;
assign w33773 = ~a_14 & w8496;
assign w33774 = ~a_14 & w33772;
assign w33775 = ~w2736 & w5308;
assign w33776 = a_20 & ~w8506;
assign w33777 = a_20 & ~w31658;
assign w33778 = ~a_20 & w8506;
assign w33779 = ~a_20 & w31658;
assign w33780 = ~w6063 & w8522;
assign w33781 = a_17 & ~w8522;
assign w33782 = a_17 & ~w33780;
assign w33783 = ~w6447 & w8550;
assign w33784 = ~a_14 & w8550;
assign w33785 = ~a_14 & w33783;
assign w33786 = ~w2736 & w6998;
assign w33787 = ~w8560 & ~a_14;
assign w33788 = w8560 & a_14;
assign w33789 = ~w8414 & a_17;
assign w33790 = ~w2465 & w6998;
assign w33791 = ~w2588 & w6446;
assign w33792 = ~w8576 & ~w8578;
assign w33793 = ~w2465 & w6446;
assign w33794 = ~w8596 & a_14;
assign w33795 = w8596 & ~a_14;
assign w33796 = ~w2736 & w6996;
assign w33797 = ~w2736 & w6446;
assign w33798 = a_14 & ~w8645;
assign w33799 = a_14 & ~w31671;
assign w33800 = ~a_14 & w8645;
assign w33801 = ~a_14 & w31671;
assign w33802 = ~w6447 & w8668;
assign w33803 = ~a_14 & w8668;
assign w33804 = ~a_14 & w33802;
assign w33805 = ~w6486 & w8592;
assign w33806 = ~w6485 & w8689;
assign w33807 = w8693 & ~a_14;
assign w33808 = ~w8693 & a_14;
assign w33809 = ~w3206 & w6996;
assign w33810 = ~w3273 & w6447;
assign w33811 = ~w8720 & a_14;
assign w33812 = w8720 & ~a_14;
assign w33813 = w8724 & ~w8726;
assign w33814 = ~w6486 & w8419;
assign w33815 = ~w6485 & w8750;
assign w33816 = w8754 & ~a_17;
assign w33817 = ~w8754 & a_17;
assign w33818 = ~w6447 & w8778;
assign w33819 = ~a_14 & ~w8778;
assign w33820 = ~a_14 & ~w33818;
assign w33821 = w8793 & ~a_20;
assign w33822 = ~w8793 & a_20;
assign w33823 = ~w3273 & w8391;
assign w33824 = ~w3206 & w6304;
assign w33825 = w8814 & a_17;
assign w33826 = ~w3273 & w6063;
assign w33827 = ~w8814 & ~a_17;
assign w33828 = w8537 & w8500;
assign w33829 = ~w8531 & ~w8769;
assign w33830 = ~w3206 & w6446;
assign w33831 = ~w6447 & w8841;
assign w33832 = ~a_14 & w8841;
assign w33833 = ~a_14 & w33831;
assign w33834 = w8848 & ~w8728;
assign w33835 = ~w7193 & w8866;
assign w33836 = ~a_11 & w8866;
assign w33837 = ~a_11 & w33835;
assign w33838 = w31574 & w5309;
assign w33839 = w8887 & ~w8882;
assign w33840 = w8887 & ~w31678;
assign w33841 = ~w3206 & w6061;
assign w33842 = ~w6063 & w8908;
assign w33843 = ~a_17 & ~w8908;
assign w33844 = ~a_17 & ~w33842;
assign w33845 = ~w3515 & w6996;
assign w33846 = ~w6447 & w8923;
assign w33847 = ~a_14 & w8923;
assign w33848 = ~a_14 & w33846;
assign w33849 = ~w3515 & w7192;
assign w33850 = ~w7193 & w8949;
assign w33851 = ~a_11 & ~w8949;
assign w33852 = ~a_11 & ~w33850;
assign w33853 = ~w8537 & ~w8500;
assign w33854 = ~w3515 & w7489;
assign w33855 = ~w7193 & w8970;
assign w33856 = ~a_11 & ~w8970;
assign w33857 = ~a_11 & ~w33855;
assign w33858 = ~w8965 & ~w8974;
assign w33859 = ~w3206 & w7192;
assign w33860 = ~w7193 & w8992;
assign w33861 = ~a_11 & w8992;
assign w33862 = ~a_11 & w33860;
assign w33863 = ~w8684 & w8708;
assign w33864 = ~w3206 & w7489;
assign w33865 = ~w7193 & w9009;
assign w33866 = ~a_11 & ~w9009;
assign w33867 = ~a_11 & ~w33865;
assign w33868 = ~w3206 & w7511;
assign w33869 = ~w3273 & w7193;
assign w33870 = ~w9035 & a_11;
assign w33871 = w9035 & ~a_11;
assign w33872 = ~w7193 & w9047;
assign w33873 = ~a_11 & w9047;
assign w33874 = ~a_11 & w33872;
assign w33875 = ~w2736 & w7489;
assign w33876 = ~w9057 & ~a_11;
assign w33877 = w9057 & a_11;
assign w33878 = ~w8587 & a_14;
assign w33879 = ~w2465 & w7489;
assign w33880 = ~w2588 & w7192;
assign w33881 = ~w9073 & ~w9075;
assign w33882 = ~w2465 & w7192;
assign w33883 = ~w9093 & a_11;
assign w33884 = w9093 & ~a_11;
assign w33885 = ~w2736 & w7511;
assign w33886 = ~w2736 & w7192;
assign w33887 = a_11 & ~w9142;
assign w33888 = a_11 & ~w31690;
assign w33889 = ~a_11 & w9142;
assign w33890 = ~a_11 & w31690;
assign w33891 = ~w7193 & w9165;
assign w33892 = ~a_11 & w9165;
assign w33893 = ~a_11 & w33891;
assign w33894 = ~w6486 & w9089;
assign w33895 = ~w6485 & w9186;
assign w33896 = w9190 & ~a_11;
assign w33897 = ~w9190 & a_11;
assign w33898 = w9040 & ~w9039;
assign w33899 = ~w7193 & w9218;
assign w33900 = ~a_11 & ~w9218;
assign w33901 = ~a_11 & ~w33899;
assign w33902 = ~w3515 & w7511;
assign w33903 = ~w7193 & w9238;
assign w33904 = ~a_11 & w9238;
assign w33905 = ~a_11 & w33903;
assign w33906 = ~w6486 & w8339;
assign w33907 = ~w6485 & w9272;
assign w33908 = w9276 & ~a_20;
assign w33909 = ~w9276 & a_20;
assign w33910 = ~w3206 & w6059;
assign w33911 = ~w6063 & w9298;
assign w33912 = ~a_17 & w9298;
assign w33913 = ~a_17 & w33911;
assign w33914 = ~w8897 & ~w9291;
assign w33915 = ~w3515 & w6998;
assign w33916 = ~w6447 & w9316;
assign w33917 = ~a_14 & ~w9316;
assign w33918 = ~a_14 & ~w33916;
assign w33919 = ~w7193 & w9331;
assign w33920 = ~a_11 & w9331;
assign w33921 = ~a_11 & w33919;
assign w33922 = ~w3515 & w8277;
assign w33923 = ~w8278 & w9356;
assign w33924 = ~a_8 & w9356;
assign w33925 = ~a_8 & w33923;
assign w33926 = ~w3515 & w8298;
assign w33927 = ~w8278 & w9373;
assign w33928 = ~a_8 & w9373;
assign w33929 = ~a_8 & w33927;
assign w33930 = ~w3206 & w8277;
assign w33931 = ~w8278 & w9394;
assign w33932 = ~a_8 & w9394;
assign w33933 = ~a_8 & w33931;
assign w33934 = ~w9181 & w9205;
assign w33935 = ~w3206 & w8298;
assign w33936 = ~w8278 & w9411;
assign w33937 = ~a_8 & w9411;
assign w33938 = ~a_8 & w33936;
assign w33939 = ~w3206 & w8295;
assign w33940 = ~w3273 & w8278;
assign w33941 = w9431 & a_8;
assign w33942 = ~w9431 & ~a_8;
assign w33943 = ~w8278 & w9442;
assign w33944 = ~a_8 & w9442;
assign w33945 = ~a_8 & w33943;
assign w33946 = ~w2736 & w8298;
assign w33947 = ~w9452 & ~a_8;
assign w33948 = w9452 & a_8;
assign w33949 = ~w9084 & a_11;
assign w33950 = ~w2465 & w8298;
assign w33951 = ~w2588 & w8277;
assign w33952 = ~w9468 & ~w9470;
assign w33953 = ~w2465 & w8277;
assign w33954 = ~w9488 & a_8;
assign w33955 = w9488 & ~a_8;
assign w33956 = ~w2736 & w8295;
assign w33957 = ~w2736 & w8277;
assign w33958 = a_8 & ~w9537;
assign w33959 = a_8 & ~w31708;
assign w33960 = ~a_8 & w9537;
assign w33961 = ~a_8 & w31708;
assign w33962 = ~w8278 & w9560;
assign w33963 = ~a_8 & w9560;
assign w33964 = ~a_8 & w33962;
assign w33965 = ~w6486 & w9484;
assign w33966 = ~w6485 & w9581;
assign w33967 = w9585 & ~a_8;
assign w33968 = ~w9585 & a_8;
assign w33969 = ~w8278 & w9622;
assign w33970 = ~a_8 & w9622;
assign w33971 = ~a_8 & w33969;
assign w33972 = ~w3515 & w8295;
assign w33973 = ~w8278 & w9642;
assign w33974 = ~a_8 & w9642;
assign w33975 = ~a_8 & w33973;
assign w33976 = ~w9231 & ~w9233;
assign w33977 = w9672 & a_8;
assign w33978 = ~w9672 & ~a_8;
assign w33979 = ~w9456 & ~w9674;
assign w33980 = ~w8278 & w9694;
assign w33981 = ~a_8 & w9694;
assign w33982 = ~a_8 & w33980;
assign w33983 = w8965 & w8974;
assign w33984 = w9724 & a_8;
assign w33985 = ~w9724 & ~a_8;
assign w33986 = ~w9456 & ~w9726;
assign w33987 = ~w2215 & w8295;
assign w33988 = ~w8278 & w9749;
assign w33989 = ~a_8 & w9749;
assign w33990 = ~a_8 & w33988;
assign w33991 = ~w1887 & w9780;
assign w33992 = ~w1985 & w9786;
assign w33993 = ~w1561 & w9788;
assign w33994 = ~w9790 & w9792;
assign w33995 = ~a_5 & ~w9792;
assign w33996 = ~a_5 & ~w33994;
assign w33997 = ~w2215 & w8277;
assign w33998 = ~w3699 & w8298;
assign w33999 = ~w3646 & w8295;
assign w34000 = ~w8278 & w9816;
assign w34001 = ~w6063 & w9837;
assign w34002 = ~a_17 & ~w9837;
assign w34003 = ~a_17 & ~w34001;
assign w34004 = ~w3206 & w5816;
assign w34005 = ~w3273 & w5309;
assign w34006 = ~w9847 & a_20;
assign w34007 = w9847 & ~a_20;
assign w34008 = ~w3515 & w6446;
assign w34009 = ~w6447 & w9875;
assign w34010 = ~a_14 & w9875;
assign w34011 = ~a_14 & w34009;
assign w34012 = w9882 & a_11;
assign w34013 = ~w9882 & ~a_11;
assign w34014 = ~w9061 & ~w9884;
assign w34015 = ~w3515 & w9786;
assign w34016 = ~w9790 & w9914;
assign w34017 = ~a_5 & w9914;
assign w34018 = ~a_5 & w34016;
assign w34019 = w9614 & ~w9421;
assign w34020 = ~w3515 & w9780;
assign w34021 = ~w9790 & w9930;
assign w34022 = ~a_5 & w9930;
assign w34023 = ~a_5 & w34021;
assign w34024 = ~w3515 & w9788;
assign w34025 = ~w9790 & w9951;
assign w34026 = ~a_5 & w9951;
assign w34027 = ~a_5 & w34025;
assign w34028 = ~w3206 & w9786;
assign w34029 = ~w9790 & w9971;
assign w34030 = ~a_5 & w9971;
assign w34031 = ~a_5 & w34029;
assign w34032 = ~w9576 & w9600;
assign w34033 = ~w3206 & w9780;
assign w34034 = ~w9790 & w9988;
assign w34035 = ~a_5 & w9988;
assign w34036 = ~a_5 & w34034;
assign w34037 = ~w3206 & w9788;
assign w34038 = ~w3273 & w9790;
assign w34039 = w10008 & a_5;
assign w34040 = ~w10008 & ~a_5;
assign w34041 = ~w9790 & w10019;
assign w34042 = ~a_5 & ~w10019;
assign w34043 = ~a_5 & ~w34041;
assign w34044 = ~w2736 & w9780;
assign w34045 = ~w10029 & ~a_5;
assign w34046 = w10029 & a_5;
assign w34047 = ~w9479 & a_8;
assign w34048 = ~w2588 & w9776;
assign w34049 = ~w2588 & w9780;
assign w34050 = ~w2465 & w9788;
assign w34051 = ~w9790 & w10049;
assign w34052 = ~w2588 & w9786;
assign w34053 = ~w2465 & w9780;
assign w34054 = ~w10053 & ~w10054;
assign w34055 = w31714 & a_5;
assign w34056 = ~w10058 & ~w9477;
assign w34057 = ~w2465 & w9786;
assign w34058 = ~w10065 & a_5;
assign w34059 = w10065 & ~a_5;
assign w34060 = ~w2736 & w9788;
assign w34061 = ~w9790 & w10100;
assign w34062 = ~a_5 & w10100;
assign w34063 = ~a_5 & w34061;
assign w34064 = ~w2736 & w9786;
assign w34065 = ~a_5 & w10110;
assign w34066 = ~a_5 & w31718;
assign w34067 = a_5 & ~w10110;
assign w34068 = a_5 & ~w31718;
assign w34069 = ~w9790 & w10133;
assign w34070 = a_5 & ~w10133;
assign w34071 = a_5 & ~w34069;
assign w34072 = ~w6486 & w10061;
assign w34073 = ~w6485 & w10149;
assign w34074 = w10153 & ~a_5;
assign w34075 = ~w10153 & a_5;
assign w34076 = ~w9790 & w10196;
assign w34077 = ~a_5 & ~w10196;
assign w34078 = ~a_5 & ~w34076;
assign w34079 = w9635 & ~w9637;
assign w34080 = ~w9790 & w10221;
assign w34081 = ~a_5 & w10221;
assign w34082 = ~a_5 & w34080;
assign w34083 = ~w9790 & w10237;
assign w34084 = ~a_5 & w10237;
assign w34085 = ~a_5 & w34083;
assign w34086 = ~w2215 & w9788;
assign w34087 = ~w9790 & w10263;
assign w34088 = ~a_5 & w10263;
assign w34089 = ~a_5 & w34087;
assign w34090 = w9664 & w9382;
assign w34091 = ~w9790 & w10279;
assign w34092 = ~a_5 & ~w10279;
assign w34093 = ~a_5 & ~w34091;
assign w34094 = w9688 & ~w9708;
assign w34095 = ~w3699 & w9788;
assign w34096 = ~w2215 & w9780;
assign w34097 = ~w10306 & ~w10308;
assign w34098 = ~w10310 & a_5;
assign w34099 = w10310 & ~a_5;
assign w34100 = ~w3646 & w9788;
assign w34101 = ~w3699 & w9780;
assign w34102 = ~w2215 & w9786;
assign w34103 = ~w9790 & w10326;
assign w34104 = ~a_5 & w10326;
assign w34105 = ~a_5 & w34103;
assign w34106 = ~w3646 & w9780;
assign w34107 = ~w1985 & w9788;
assign w34108 = ~w3699 & w9786;
assign w34109 = w4791 & w9790;
assign w34110 = ~w10359 & a_5;
assign w34111 = w10359 & ~a_5;
assign w34112 = ~w3646 & w9786;
assign w34113 = ~w1985 & w9780;
assign w34114 = ~w1887 & w9788;
assign w34115 = ~w9790 & w10380;
assign w34116 = ~a_5 & w10380;
assign w34117 = ~a_5 & w34115;
assign w34118 = ~w1887 & w9786;
assign w34119 = ~w1561 & w9780;
assign w34120 = ~w1794 & w9788;
assign w34121 = ~w9790 & w10423;
assign w34122 = ~a_5 & ~w10423;
assign w34123 = ~a_5 & ~w34121;
assign w34124 = ~w2215 & w7511;
assign w34125 = ~w7193 & w10436;
assign w34126 = ~a_11 & w10436;
assign w34127 = ~a_11 & w34125;
assign w34128 = ~w3515 & w6304;
assign w34129 = ~w6063 & w10456;
assign w34130 = ~a_17 & ~w10456;
assign w34131 = ~a_17 & ~w34129;
assign w34132 = ~w3206 & w5818;
assign w34133 = ~w5309 & w10468;
assign w34134 = ~a_20 & ~w10468;
assign w34135 = ~a_20 & ~w34133;
assign w34136 = ~w6447 & w10494;
assign w34137 = ~a_14 & w10494;
assign w34138 = ~a_14 & w34136;
assign w34139 = ~w3646 & w8298;
assign w34140 = ~w3699 & w8277;
assign w34141 = ~w1985 & w8295;
assign w34142 = w4791 & w8278;
assign w34143 = w10513 & a_8;
assign w34144 = ~w10513 & ~a_8;
assign w34145 = ~w3646 & w8277;
assign w34146 = ~w1985 & w8298;
assign w34147 = ~w1887 & w8295;
assign w34148 = ~w8278 & w10571;
assign w34149 = ~a_8 & w10571;
assign w34150 = ~a_8 & w34148;
assign w34151 = ~w3515 & w6061;
assign w34152 = ~w6063 & w10591;
assign w34153 = ~a_17 & ~w10591;
assign w34154 = ~a_17 & ~w34152;
assign w34155 = ~w3206 & w5308;
assign w34156 = ~w5309 & w10603;
assign w34157 = ~a_20 & ~w10603;
assign w34158 = ~a_20 & ~w34156;
assign w34159 = ~w6447 & w10621;
assign w34160 = ~a_14 & ~w10621;
assign w34161 = ~a_14 & ~w34159;
assign w34162 = ~w3699 & w7511;
assign w34163 = ~w2215 & w7489;
assign w34164 = ~w10627 & ~w10629;
assign w34165 = ~w9089 & w10633;
assign w34166 = ~w1561 & w9786;
assign w34167 = ~w1794 & w9780;
assign w34168 = ~w10655 & ~w10656;
assign w34169 = w10658 & a_5;
assign w34170 = ~w10658 & ~a_5;
assign w34171 = ~w1887 & w8298;
assign w34172 = ~w1985 & w8277;
assign w34173 = ~w1561 & w8295;
assign w34174 = ~w10706 & a_8;
assign w34175 = w10706 & ~a_8;
assign w34176 = ~w9484 & w10710;
assign w34177 = ~w3646 & w7511;
assign w34178 = ~w2215 & w7192;
assign w34179 = ~w3699 & w7489;
assign w34180 = ~w7193 & w10720;
assign w34181 = ~a_11 & w10720;
assign w34182 = ~a_11 & w34180;
assign w34183 = ~w5309 & w10736;
assign w34184 = ~a_20 & w10736;
assign w34185 = ~a_20 & w34183;
assign w34186 = ~w3515 & w6059;
assign w34187 = ~w6063 & w10745;
assign w34188 = ~a_17 & w10745;
assign w34189 = ~a_17 & w34187;
assign w34190 = ~w10792 & a_14;
assign w34191 = w10792 & ~a_14;
assign w34192 = ~w8592 & w10796;
assign w34193 = ~w1794 & w9786;
assign w34194 = ~w9790 & w10820;
assign w34195 = ~a_5 & w10820;
assign w34196 = ~a_5 & w34194;
assign w34197 = ~w10837 & w10838;
assign w34198 = ~w1522 & w10839;
assign w34199 = ~w10841 & w10838;
assign w34200 = ~w10841 & w34197;
assign w34201 = a_2 & ~w10838;
assign w34202 = a_2 & ~w34197;
assign w34203 = w10289 & w10300;
assign w34204 = ~w3646 & w10835;
assign w34205 = ~w1985 & w3;
assign w34206 = w4791 & w10837;
assign w34207 = ~w3699 & w10839;
assign w34208 = w10858 & ~w10860;
assign w34209 = ~w10858 & a_2;
assign w34210 = ~w10837 & w10870;
assign w34211 = ~w10839 & a_2;
assign w34212 = a_2 & ~w10870;
assign w34213 = a_2 & ~w34210;
assign w34214 = w10186 & ~w9998;
assign w34215 = ~w3515 & w10835;
assign w34216 = ~w10837 & w10885;
assign w34217 = a_2 & ~w10885;
assign w34218 = a_2 & ~w34216;
assign w34219 = ~w31714 & a_5;
assign w34220 = ~w2736 & w10835;
assign w34221 = a_2 & ~w10898;
assign w34222 = a_2 & ~w31730;
assign w34223 = ~w10900 & w10895;
assign w34224 = w10058 & w9477;
assign w34225 = ~w2736 & w10909;
assign w34226 = ~a_2 & ~w10913;
assign w34227 = ~a_2 & ~w31731;
assign w34228 = a_2 & w10913;
assign w34229 = a_2 & w31731;
assign w34230 = ~w10837 & w10923;
assign w34231 = ~w2465 & w10839;
assign w34232 = ~w10927 & w10923;
assign w34233 = ~w10927 & w34230;
assign w34234 = ~w2465 & ~w10839;
assign w34235 = w2588 & a_2;
assign w34236 = w10932 & ~w10930;
assign w34237 = ~w10933 & ~w10044;
assign w34238 = ~w10934 & ~w10928;
assign w34239 = w10900 & ~w10895;
assign w34240 = ~w2736 & w3;
assign w34241 = ~w10837 & w10942;
assign w34242 = ~a_2 & w10942;
assign w34243 = ~a_2 & w34241;
assign w34244 = ~a_2 & ~w10939;
assign w34245 = ~w10837 & w10958;
assign w34246 = a_2 & w10958;
assign w34247 = a_2 & w34245;
assign w34248 = w10961 & ~w10955;
assign w34249 = ~w10837 & w10972;
assign w34250 = a_2 & ~w10972;
assign w34251 = a_2 & ~w34249;
assign w34252 = ~w10837 & w10986;
assign w34253 = a_2 & ~w10986;
assign w34254 = a_2 & ~w34252;
assign w34255 = ~w10991 & ~w10980;
assign w34256 = ~w10837 & w10997;
assign w34257 = a_2 & ~w10997;
assign w34258 = a_2 & ~w34256;
assign w34259 = ~w10121 & ~w10119;
assign w34260 = ~w3206 & w3;
assign w34261 = ~w3273 & w10837;
assign w34262 = ~w11017 & a_2;
assign w34263 = ~w3206 & w10835;
assign w34264 = ~w10837 & w11034;
assign w34265 = a_2 & ~w11034;
assign w34266 = a_2 & ~w34264;
assign w34267 = w11039 & ~w11026;
assign w34268 = w10172 & w10168;
assign w34269 = ~w10837 & w11047;
assign w34270 = a_2 & ~w11047;
assign w34271 = a_2 & ~w34269;
assign w34272 = ~w10837 & w11061;
assign w34273 = a_2 & ~w11061;
assign w34274 = a_2 & ~w34272;
assign w34275 = w11066 & ~w11056;
assign w34276 = ~w3515 & w3;
assign w34277 = ~w10837 & w11071;
assign w34278 = a_2 & ~w11071;
assign w34279 = a_2 & ~w34277;
assign w34280 = ~w10837 & w11093;
assign w34281 = a_2 & ~w11093;
assign w34282 = a_2 & ~w34280;
assign w34283 = w10201 & ~w10203;
assign w34284 = ~w10837 & w11110;
assign w34285 = a_2 & ~w11110;
assign w34286 = a_2 & ~w34284;
assign w34287 = w10211 & w9939;
assign w34288 = ~w10837 & w11132;
assign w34289 = a_2 & ~w11132;
assign w34290 = a_2 & ~w34288;
assign w34291 = ~w11129 & w11137;
assign w34292 = ~w11140 & ~w11138;
assign w34293 = ~w2215 & w3;
assign w34294 = ~w10837 & w11148;
assign w34295 = a_2 & ~w11148;
assign w34296 = a_2 & ~w34294;
assign w34297 = w11129 & ~w11137;
assign w34298 = w11153 & ~w11156;
assign w34299 = ~w3699 & w3;
assign w34300 = ~w2215 & w10835;
assign w34301 = ~w10837 & w11163;
assign w34302 = a_2 & ~w11163;
assign w34303 = a_2 & ~w34301;
assign w34304 = ~w11160 & w11168;
assign w34305 = ~w3646 & w3;
assign w34306 = ~w3699 & w10835;
assign w34307 = ~w10837 & w11178;
assign w34308 = a_2 & ~w11178;
assign w34309 = a_2 & ~w34307;
assign w34310 = w11160 & ~w11168;
assign w34311 = w10289 & w11183;
assign w34312 = ~w1887 & w3;
assign w34313 = ~w1985 & w10835;
assign w34314 = ~w10837 & w11204;
assign w34315 = a_2 & ~w11204;
assign w34316 = a_2 & ~w34314;
assign w34317 = ~w1887 & w10835;
assign w34318 = ~w1561 & w3;
assign w34319 = ~w10837 & w11217;
assign w34320 = a_2 & ~w11217;
assign w34321 = a_2 & ~w34319;
assign w34322 = ~w11214 & w11222;
assign w34323 = ~w1794 & w3;
assign w34324 = ~w1561 & w10835;
assign w34325 = ~w10837 & w11232;
assign w34326 = a_2 & ~w11232;
assign w34327 = a_2 & ~w34325;
assign w34328 = w11214 & ~w11222;
assign w34329 = ~w1794 & w10835;
assign w34330 = ~w10837 & w11252;
assign w34331 = a_2 & ~w11252;
assign w34332 = a_2 & ~w34330;
assign w34333 = w10341 & w11237;
assign w34334 = ~w10837 & w11272;
assign w34335 = a_2 & ~w11272;
assign w34336 = a_2 & ~w34334;
assign w34337 = ~w1522 & w3;
assign w34338 = ~w10837 & w11291;
assign w34339 = a_2 & ~w11291;
assign w34340 = a_2 & ~w34338;
assign w34341 = ~w1522 & w10835;
assign w34342 = ~w10837 & w11310;
assign w34343 = a_2 & ~w11310;
assign w34344 = a_2 & ~w34342;
assign w34345 = ~w1522 & w9788;
assign w34346 = ~w11357 & ~w11358;
assign w34347 = w11360 & a_5;
assign w34348 = ~w11360 & ~a_5;
assign w34349 = ~w1887 & w8277;
assign w34350 = ~w1561 & w8298;
assign w34351 = ~w1794 & w8295;
assign w34352 = ~w8278 & w11391;
assign w34353 = ~a_8 & ~w11391;
assign w34354 = ~a_8 & ~w34352;
assign w34355 = ~w6063 & w11412;
assign w34356 = ~a_17 & w11412;
assign w34357 = ~a_17 & w34355;
assign w34358 = ~w5306 & ~a_20;
assign w34359 = ~w3515 & w5816;
assign w34360 = ~w11420 & ~w11417;
assign w34361 = w11420 & ~a_20;
assign w34362 = ~w11420 & ~a_20;
assign w34363 = ~w11425 & ~w11424;
assign w34364 = ~w2215 & w6996;
assign w34365 = ~w6447 & w11448;
assign w34366 = ~a_14 & w11448;
assign w34367 = ~a_14 & w34365;
assign w34368 = w4791 & w7193;
assign w34369 = ~w1985 & w7511;
assign w34370 = ~w3699 & w7192;
assign w34371 = ~w3646 & w7489;
assign w34372 = ~w11458 & a_11;
assign w34373 = w11458 & ~a_11;
assign w34374 = ~w1322 & w3;
assign w34375 = ~w10837 & w11488;
assign w34376 = a_2 & ~w11488;
assign w34377 = a_2 & ~w34375;
assign w34378 = ~w11451 & w10798;
assign w34379 = ~w2215 & w6998;
assign w34380 = ~w3699 & w6996;
assign w34381 = ~w11561 & ~w11563;
assign w34382 = ~w11565 & a_14;
assign w34383 = w11565 & ~a_14;
assign w34384 = ~w3515 & w5818;
assign w34385 = ~w5309 & w11577;
assign w34386 = ~a_20 & ~w11577;
assign w34387 = ~a_20 & ~w34385;
assign w34388 = ~w6063 & w11596;
assign w34389 = ~a_17 & w11596;
assign w34390 = ~a_17 & w34388;
assign w34391 = ~w3646 & w7192;
assign w34392 = ~w1985 & w7489;
assign w34393 = ~w1887 & w7511;
assign w34394 = ~w7193 & w11617;
assign w34395 = ~a_11 & w11617;
assign w34396 = ~a_11 & w34394;
assign w34397 = ~w1794 & w8298;
assign w34398 = ~w1561 & w8277;
assign w34399 = ~w9484 & w11630;
assign w34400 = ~w1522 & w9780;
assign w34401 = ~w9790 & w11648;
assign w34402 = ~a_5 & ~w11648;
assign w34403 = ~a_5 & ~w34401;
assign w34404 = ~w3905 & w3;
assign w34405 = ~w1322 & w10835;
assign w34406 = ~w10837 & w11666;
assign w34407 = a_2 & ~w11666;
assign w34408 = a_2 & ~w34406;
assign w34409 = ~w3905 & w10835;
assign w34410 = ~w10837 & w11691;
assign w34411 = a_2 & ~w11691;
assign w34412 = a_2 & ~w34410;
assign w34413 = ~w1522 & w9786;
assign w34414 = w11701 & a_5;
assign w34415 = ~w11701 & ~a_5;
assign w34416 = ~w10033 & ~w11703;
assign w34417 = ~w1887 & w7489;
assign w34418 = ~w1985 & w7192;
assign w34419 = ~w1561 & w7511;
assign w34420 = ~w7193 & w11740;
assign w34421 = ~a_11 & ~w11740;
assign w34422 = ~a_11 & ~w34420;
assign w34423 = ~w3646 & w6996;
assign w34424 = ~w3699 & w6998;
assign w34425 = ~w2215 & w6446;
assign w34426 = ~w6447 & w11752;
assign w34427 = ~a_14 & w11752;
assign w34428 = ~a_14 & w34426;
assign w34429 = ~w3515 & w5308;
assign w34430 = ~w5309 & w11764;
assign w34431 = ~a_20 & w11764;
assign w34432 = ~a_20 & w34430;
assign w34433 = ~w11772 & a_17;
assign w34434 = w11772 & ~a_17;
assign w34435 = ~w8419 & w11776;
assign w34436 = ~w1794 & w8277;
assign w34437 = ~w11796 & ~w11797;
assign w34438 = w11798 & ~a_8;
assign w34439 = ~w11798 & a_8;
assign w34440 = ~w10837 & ~w11831;
assign w34441 = a_2 & w11831;
assign w34442 = a_2 & ~w34440;
assign w34443 = ~w1322 & w9788;
assign w34444 = ~w9790 & w11856;
assign w34445 = ~a_5 & w11856;
assign w34446 = ~a_5 & w34444;
assign w34447 = w11790 & ~w11756;
assign w34448 = ~w5309 & w11887;
assign w34449 = ~a_20 & w11887;
assign w34450 = ~a_20 & w34448;
assign w34451 = ~w2215 & w6304;
assign w34452 = ~w6063 & w11899;
assign w34453 = ~a_17 & w11899;
assign w34454 = ~a_17 & w34452;
assign w34455 = ~w3646 & w6998;
assign w34456 = ~w1985 & w6996;
assign w34457 = ~w3699 & w6446;
assign w34458 = w4791 & w6447;
assign w34459 = ~w11909 & a_14;
assign w34460 = w11909 & ~a_14;
assign w34461 = ~w1794 & w7511;
assign w34462 = ~w1561 & w7489;
assign w34463 = ~w1887 & w7192;
assign w34464 = ~w7193 & w11932;
assign w34465 = ~a_11 & w11932;
assign w34466 = ~a_11 & w34464;
assign w34467 = ~w1522 & w8295;
assign w34468 = ~w11938 & ~w11939;
assign w34469 = ~w11941 & a_8;
assign w34470 = w11941 & ~a_8;
assign w34471 = ~w1322 & w9780;
assign w34472 = ~w3905 & w9788;
assign w34473 = ~w9790 & w11991;
assign w34474 = ~a_5 & w11991;
assign w34475 = ~a_5 & w34473;
assign w34476 = a_0 & w32759;
assign w34477 = a_0 & w32760;
assign w34478 = ~w11994 & ~w11999;
assign w34479 = w11994 & w11999;
assign w34480 = ~w1522 & w8298;
assign w34481 = ~w8278 & w12018;
assign w34482 = ~a_8 & ~w12018;
assign w34483 = ~a_8 & ~w34481;
assign w34484 = ~w1561 & w7192;
assign w34485 = ~w1794 & w7489;
assign w34486 = ~w12031 & ~w12032;
assign w34487 = ~w12034 & a_11;
assign w34488 = w12034 & ~a_11;
assign w34489 = ~w5309 & w12042;
assign w34490 = ~a_20 & w12042;
assign w34491 = ~a_20 & w34489;
assign w34492 = ~w2215 & w6061;
assign w34493 = ~w3699 & w6304;
assign w34494 = ~w12053 & ~w12055;
assign w34495 = ~w12057 & a_17;
assign w34496 = w12057 & ~a_17;
assign w34497 = ~w3646 & w6446;
assign w34498 = ~w1985 & w6998;
assign w34499 = ~w1887 & w6996;
assign w34500 = ~w6447 & w12065;
assign w34501 = ~a_14 & w12065;
assign w34502 = ~a_14 & w34500;
assign w34503 = ~w12012 & ~w12084;
assign w34504 = w12012 & w12084;
assign w34505 = w12114 & ~w12119;
assign w34506 = ~w3905 & w9780;
assign w34507 = ~w1322 & w9786;
assign w34508 = ~w9790 & w12125;
assign w34509 = ~a_5 & ~w12125;
assign w34510 = ~a_5 & ~w34508;
assign w34511 = ~w12135 & ~w12141;
assign w34512 = ~w1522 & w8277;
assign w34513 = ~w8278 & w12147;
assign w34514 = a_8 & ~w12147;
assign w34515 = a_8 & ~w34513;
assign w34516 = ~w1794 & w7192;
assign w34517 = ~w12157 & ~w12158;
assign w34518 = ~w12159 & a_11;
assign w34519 = w12159 & ~a_11;
assign w34520 = ~w3646 & w6304;
assign w34521 = ~w3699 & w6061;
assign w34522 = ~w2215 & w6059;
assign w34523 = ~w6063 & w12169;
assign w34524 = ~a_17 & w12169;
assign w34525 = ~a_17 & w34523;
assign w34526 = ~w1887 & w6998;
assign w34527 = ~w1985 & w6446;
assign w34528 = ~w12177 & a_14;
assign w34529 = w12177 & ~a_14;
assign w34530 = ~w8592 & w12181;
assign w34531 = ~w3905 & w9786;
assign w34532 = ~w9790 & w12223;
assign w34533 = ~a_5 & w12223;
assign w34534 = ~a_5 & w34532;
assign w34535 = w12151 & ~w12227;
assign w34536 = ~w12151 & w12227;
assign w34537 = ~w1322 & w8295;
assign w34538 = ~w8278 & w12238;
assign w34539 = ~a_8 & w12238;
assign w34540 = ~a_8 & w34538;
assign w34541 = ~w12164 & w12152;
assign w34542 = ~w12164 & ~w32443;
assign w34543 = w12164 & ~w12152;
assign w34544 = w12164 & w32443;
assign w34545 = ~w1887 & w6446;
assign w34546 = ~w1794 & w6996;
assign w34547 = ~w6447 & w12256;
assign w34548 = ~a_14 & ~w12256;
assign w34549 = ~a_14 & ~w34547;
assign w34550 = ~w1522 & w7511;
assign w34551 = ~w12271 & ~w12272;
assign w34552 = ~w12274 & a_11;
assign w34553 = w12274 & ~a_11;
assign w34554 = ~w12139 & ~w12286;
assign w34555 = ~w1522 & w7192;
assign w34556 = ~w7193 & w12307;
assign w34557 = ~a_11 & w12307;
assign w34558 = ~a_11 & w34556;
assign w34559 = w12260 & ~w12249;
assign w34560 = ~w1522 & w7489;
assign w34561 = ~w7193 & w12324;
assign w34562 = ~a_11 & ~w12324;
assign w34563 = ~a_11 & ~w34561;
assign w34564 = w12328 & ~w12317;
assign w34565 = ~w12263 & ~w12278;
assign w34566 = ~w3905 & w8295;
assign w34567 = ~w1322 & w8298;
assign w34568 = ~w8278 & w12346;
assign w34569 = ~a_8 & w12346;
assign w34570 = ~a_8 & w34568;
assign w34571 = w12355 & ~w12351;
assign w34572 = ~w3905 & w8298;
assign w34573 = ~w1322 & w8277;
assign w34574 = ~w8278 & w12362;
assign w34575 = ~a_8 & ~w12362;
assign w34576 = ~a_8 & ~w34574;
assign w34577 = w9790 & ~w32757;
assign w34578 = w9790 & ~w32758;
assign w34579 = ~w9786 & ~w34577;
assign w34580 = ~w9786 & ~w34578;
assign w34581 = ~w3958 & ~a_5;
assign w34582 = w3958 & a_5;
assign w34583 = ~w12231 & w12227;
assign w34584 = w12295 & ~w12398;
assign w34585 = w12298 & ~w12402;
assign w34586 = ~w3905 & w8277;
assign w34587 = ~w8278 & w12412;
assign w34588 = ~a_8 & w12412;
assign w34589 = ~a_8 & w34587;
assign w34590 = ~w12337 & ~w12332;
assign w34591 = ~w12340 & ~w12367;
assign w34592 = ~w12425 & ~w12429;
assign w34593 = ~w12405 & w12431;
assign w34594 = w12425 & ~w12436;
assign w34595 = w12435 & ~w7878;
assign w34596 = ~w12439 & w31760;
assign w34597 = ~w33578 & ~w7056;
assign w34598 = w12443 & ~w31760;
assign w34599 = w12443 & ~w34596;
assign w34600 = ~w12447 & ~w34598;
assign w34601 = ~w12447 & ~w34599;
assign w34602 = w12451 & ~w34600;
assign w34603 = w12451 & ~w34601;
assign w34604 = w6461 & ~w6331;
assign w34605 = ~w1522 & w5080;
assign w34606 = ~w5017 & w12459;
assign w34607 = ~a_23 & w12459;
assign w34608 = ~a_23 & w34606;
assign w34609 = w6028 & ~w6017;
assign w34610 = w6013 & ~w6033;
assign w34611 = ~w3905 & w5816;
assign w34612 = ~w1322 & w5818;
assign w34613 = ~w5309 & w12481;
assign w34614 = ~a_20 & w12481;
assign w34615 = ~a_20 & w34613;
assign w34616 = ~w6005 & ~w6040;
assign w34617 = w6063 & ~w32757;
assign w34618 = w6063 & ~w32758;
assign w34619 = w6059 & ~w3958;
assign w34620 = a_17 & w3958;
assign w34621 = a_17 & ~w34619;
assign w34622 = w6068 & ~w6046;
assign w34623 = w6071 & ~w12502;
assign w34624 = w12503 & w6331;
assign w34625 = w12503 & ~w34604;
assign w34626 = ~w12488 & ~w12495;
assign w34627 = ~w12463 & ~w12467;
assign w34628 = ~w1522 & w5016;
assign w34629 = ~w5017 & w12513;
assign w34630 = ~a_23 & w12513;
assign w34631 = ~a_23 & w34629;
assign w34632 = ~w12485 & ~w12474;
assign w34633 = ~w3905 & w5818;
assign w34634 = ~w1322 & w5308;
assign w34635 = ~w5309 & w12529;
assign w34636 = ~a_20 & ~w12529;
assign w34637 = ~a_20 & ~w34635;
assign w34638 = ~w12523 & ~w12534;
assign w34639 = w12506 & ~w12518;
assign w34640 = ~w3905 & w5308;
assign w34641 = ~w5309 & w12553;
assign w34642 = ~a_20 & ~w12553;
assign w34643 = ~a_20 & ~w34641;
assign w34644 = w12557 & ~w12548;
assign w34645 = w12570 & ~w34624;
assign w34646 = w12570 & ~w34625;
assign w34647 = w12576 & ~w34645;
assign w34648 = w12576 & ~w34646;
assign w34649 = ~w5338 & ~w5350;
assign w34650 = ~w5355 & ~w12581;
assign w34651 = w12580 & ~w12583;
assign w34652 = ~w34650 & w12585;
assign w34653 = w12586 & ~w12585;
assign w34654 = w12586 & ~w34652;
assign w34655 = w4697 & ~w34653;
assign w34656 = w4697 & ~w34654;
assign w34657 = ~w4695 & ~w4650;
assign w34658 = ~w34657 & ~w4649;
assign w34659 = ~w4501 & ~w4499;
assign w34660 = w12591 & w4499;
assign w34661 = w12591 & ~w34659;
assign w34662 = ~w4477 & ~w34660;
assign w34663 = ~w4477 & ~w34661;
assign w34664 = w12594 & ~w34662;
assign w34665 = w12594 & ~w34663;
assign w34666 = ~w4083 & ~w34664;
assign w34667 = ~w4083 & ~w34665;
assign w34668 = w3976 & ~w34666;
assign w34669 = w3976 & ~w34667;
assign w34670 = ~w3976 & w34666;
assign w34671 = ~w3976 & w34667;
assign w34672 = ~w12594 & w34662;
assign w34673 = ~w12594 & w34663;
assign w34674 = ~w12591 & ~w4499;
assign w34675 = ~w12591 & w34659;
assign w34676 = ~w4501 & w4649;
assign w34677 = ~w4501 & ~w34658;
assign w34678 = ~w12609 & ~w34655;
assign w34679 = ~w12609 & ~w34656;
assign w34680 = ~w5092 & ~w12585;
assign w34681 = ~w5092 & ~w34652;
assign w34682 = w4695 & w4650;
assign w34683 = ~w4695 & w4649;
assign w34684 = ~w12619 & ~w34598;
assign w34685 = ~w12619 & ~w34599;
assign w34686 = w12619 & w34598;
assign w34687 = w12619 & w34599;
assign w34688 = ~w12439 & w31761;
assign w34689 = w7507 & w31761;
assign w34690 = w7507 & w34688;
assign w34691 = w7207 & ~w7058;
assign w34692 = ~w12627 & ~w34689;
assign w34693 = ~w12627 & ~w34690;
assign w34694 = w7058 & w34689;
assign w34695 = w7058 & w34690;
assign w34696 = w31762 & w12438;
assign w34697 = (w12438 & w31762) | (w12438 & w12405) | (w31762 & w12405);
assign w34698 = w31763 & w12642;
assign w34699 = (w12642 & w31763) | (w12642 & w12405) | (w31763 & w12405);
assign w34700 = w32447 | w32446;
assign w34701 = (w32446 & w32447) | (w32446 & ~w12405) | (w32447 & ~w12405);
assign w34702 = w32449 | w32448;
assign w34703 = (w32448 & w32449) | (w32448 & ~w12405) | (w32449 & ~w12405);
assign w34704 = w31765 & ~w12623;
assign w34705 = (~w12623 & w31765) | (~w12623 & w12439) | (w31765 & w12439);
assign w34706 = w12666 & ~w31761;
assign w34707 = w12666 & ~w34688;
assign w34708 = w12666 & w34704;
assign w34709 = w12666 & w34705;
assign w34710 = ~w12666 & ~w34704;
assign w34711 = ~w12666 & ~w34705;
assign w34712 = w12217 & w12299;
assign w34713 = ~w12651 & ~w12652;
assign w34714 = w32453 & ~w12662;
assign w34715 = ~w12833 & w12837;
assign w34716 = ~w12850 & w34684;
assign w34717 = ~w12850 & w34685;
assign w34718 = w12850 & ~w34684;
assign w34719 = w12850 & ~w34685;
assign w34720 = w12853 & ~w12631;
assign w34721 = w12853 & w31782;
assign w34722 = w12848 & ~w34686;
assign w34723 = w12848 & ~w34687;
assign w34724 = ~w12454 & w6331;
assign w34725 = ~w12454 & ~w34604;
assign w34726 = w6461 & w12454;
assign w34727 = ~w12857 & ~w12859;
assign w34728 = ~w12861 & w34720;
assign w34729 = ~w12861 & w34721;
assign w34730 = ~w12856 & ~w12863;
assign w34731 = w12866 & ~w34724;
assign w34732 = w12866 & ~w34725;
assign w34733 = ~w12866 & w34724;
assign w34734 = ~w12866 & w34725;
assign w34735 = w12865 & ~w12870;
assign w34736 = w12543 & ~w34624;
assign w34737 = w12543 & ~w34625;
assign w34738 = w12872 & ~w34731;
assign w34739 = w12872 & ~w34732;
assign w34740 = ~w12540 & ~w34736;
assign w34741 = ~w12540 & ~w34737;
assign w34742 = w12875 & w34740;
assign w34743 = w12875 & w34741;
assign w34744 = ~w12875 & ~w34740;
assign w34745 = ~w12875 & ~w34741;
assign w34746 = w12881 & w34733;
assign w34747 = w12881 & w34734;
assign w34748 = ~w12881 & ~w34733;
assign w34749 = ~w12881 & ~w34734;
assign w34750 = w12869 & ~w12884;
assign w34751 = ~w34735 & w12886;
assign w34752 = w12574 & ~w34736;
assign w34753 = w12574 & ~w34737;
assign w34754 = ~w12561 & ~w34752;
assign w34755 = ~w12561 & ~w34753;
assign w34756 = ~w12890 & ~w34754;
assign w34757 = ~w12890 & ~w34755;
assign w34758 = w12896 & ~w12886;
assign w34759 = w12896 & ~w34751;
assign w34760 = w12899 & w34756;
assign w34761 = w12899 & w34757;
assign w34762 = ~w12899 & ~w34756;
assign w34763 = ~w12899 & ~w34757;
assign w34764 = ~w12878 & ~w12902;
assign w34765 = w12903 & ~w34758;
assign w34766 = w12903 & ~w34759;
assign w34767 = ~w12890 & w12898;
assign w34768 = w5355 & ~w12907;
assign w34769 = ~w5355 & w12907;
assign w34770 = ~w34650 & ~w12582;
assign w34771 = ~w12912 & w12582;
assign w34772 = ~w12912 & ~w34770;
assign w34773 = w12911 & w12921;
assign w34774 = w12924 & w34771;
assign w34775 = w12924 & w34772;
assign w34776 = ~w12924 & ~w34771;
assign w34777 = ~w12924 & ~w34772;
assign w34778 = ~w12910 & ~w12927;
assign w34779 = w12928 & ~w12921;
assign w34780 = w12928 & ~w34773;
assign w34781 = ~w12912 & w12923;
assign w34782 = ~w12932 & w34779;
assign w34783 = ~w12932 & w34780;
assign w34784 = w12611 & w12610;
assign w34785 = ~w12936 & w12938;
assign w34786 = ~w12618 & ~w12938;
assign w34787 = ~w12618 & ~w34785;
assign w34788 = ~w12943 & ~w34786;
assign w34789 = ~w12943 & ~w34787;
assign w34790 = ~w12947 & ~w12608;
assign w34791 = w12950 & w12608;
assign w34792 = w12950 & ~w34790;
assign w34793 = w4083 & ~w34662;
assign w34794 = w4083 & ~w34663;
assign w34795 = w12593 & w34662;
assign w34796 = w12593 & w34663;
assign w34797 = w12958 & ~w34791;
assign w34798 = w12958 & ~w34792;
assign w34799 = ~w12948 & ~w34791;
assign w34800 = ~w12948 & ~w34792;
assign w34801 = ~w12957 & ~w34799;
assign w34802 = ~w12957 & ~w34800;
assign w34803 = ~w1478 & w12963;
assign w34804 = ~w666 & ~w664;
assign w34805 = w1463 & w12976;
assign w34806 = w3945 & ~w3865;
assign w34807 = ~w3859 & ~w12993;
assign w34808 = w3859 & w12993;
assign w34809 = ~w1478 & ~w12997;
assign w34810 = ~w12996 & ~w12997;
assign w34811 = ~w12996 & w34809;
assign w34812 = w13007 & w34670;
assign w34813 = w13007 & w34671;
assign w34814 = ~w13007 & ~w34670;
assign w34815 = ~w13007 & ~w34671;
assign w34816 = w13007 & ~w34668;
assign w34817 = w13007 & ~w34669;
assign w34818 = ~w13012 & w668;
assign w34819 = ~w13017 & ~w34797;
assign w34820 = ~w13017 & ~w34798;
assign w34821 = ~w1478 & w13023;
assign w34822 = ~w12981 & w13023;
assign w34823 = ~w12981 & w34821;
assign w34824 = ~w13026 & ~w12966;
assign w34825 = w13026 & w12966;
assign w34826 = w13047 & w3999;
assign w34827 = ~a_20 & ~w13110;
assign w34828 = w13111 & ~w13108;
assign w34829 = w12614 & w1327;
assign w34830 = w12610 & w1399;
assign w34831 = ~w12606 & w668;
assign w34832 = w12943 & w34786;
assign w34833 = w12943 & w34787;
assign w34834 = ~w1478 & w13125;
assign w34835 = ~w13118 & ~w13116;
assign w34836 = w13129 & w13116;
assign w34837 = w13129 & ~w34835;
assign w34838 = ~w13049 & ~w34836;
assign w34839 = ~w13049 & ~w34837;
assign w34840 = w13132 & ~w34838;
assign w34841 = w13132 & ~w34839;
assign w34842 = ~w13132 & w34838;
assign w34843 = ~w13132 & w34839;
assign w34844 = ~w12606 & w1399;
assign w34845 = ~w12950 & ~w12608;
assign w34846 = ~w12950 & w34790;
assign w34847 = ~w1478 & w13142;
assign w34848 = w13143 & ~w13133;
assign w34849 = ~w666 & w12963;
assign w34850 = ~w666 & w34803;
assign w34851 = ~w12996 & ~w12995;
assign w34852 = w13169 & w12995;
assign w34853 = w13169 & ~w34851;
assign w34854 = ~w13169 & ~w12995;
assign w34855 = ~w13169 & w34851;
assign w34856 = ~w3974 & ~w34668;
assign w34857 = ~w3974 & ~w34669;
assign w34858 = ~w13002 & w34856;
assign w34859 = ~w13002 & w34857;
assign w34860 = ~w13003 & ~w34858;
assign w34861 = ~w13003 & ~w34859;
assign w34862 = ~w13172 & ~w13170;
assign w34863 = w13167 & w13170;
assign w34864 = w13167 & ~w34862;
assign w34865 = ~w13167 & w34862;
assign w34866 = ~w13172 & ~w34860;
assign w34867 = ~w13172 & ~w34861;
assign w34868 = ~w13179 & w4068;
assign w34869 = ~w13012 & w3957;
assign w34870 = w13167 & ~w34854;
assign w34871 = w13167 & ~w34855;
assign w34872 = ~w13167 & w34854;
assign w34873 = ~w13167 & w34855;
assign w34874 = ~w13185 & ~w34860;
assign w34875 = ~w13185 & ~w34861;
assign w34876 = w13166 & w34852;
assign w34877 = w13166 & w34853;
assign w34878 = ~w13167 & ~w34852;
assign w34879 = ~w13167 & ~w34853;
assign w34880 = w13189 & w34860;
assign w34881 = w13189 & w34861;
assign w34882 = w13180 & w13191;
assign w34883 = ~w13003 & w34856;
assign w34884 = ~w13003 & w34857;
assign w34885 = ~w13002 & ~w34856;
assign w34886 = ~w13002 & ~w34857;
assign w34887 = ~w13011 & w34797;
assign w34888 = ~w13011 & w34798;
assign w34889 = w13200 & w13203;
assign w34890 = ~w13192 & ~w13203;
assign w34891 = ~w13192 & ~w34889;
assign w34892 = ~w13180 & ~w13191;
assign w34893 = ~w13206 & w13204;
assign w34894 = ~w4070 & w13209;
assign w34895 = ~a_29 & w13209;
assign w34896 = ~a_29 & w34894;
assign w34897 = w13148 & w13029;
assign w34898 = ~w12981 & ~w12978;
assign w34899 = w3901 & w3909;
assign w34900 = w1214 & w13222;
assign w34901 = w13223 & w13219;
assign w34902 = ~w13230 & ~w12978;
assign w34903 = ~w13230 & w34898;
assign w34904 = w13230 & w12978;
assign w34905 = w13230 & ~w34898;
assign w34906 = ~w13179 & w668;
assign w34907 = ~w13012 & w1327;
assign w34908 = ~w13200 & w13198;
assign w34909 = ~w13237 & w1478;
assign w34910 = ~w13236 & ~w13234;
assign w34911 = ~w13244 & w34890;
assign w34912 = ~w13244 & w34891;
assign w34913 = w4070 & ~w34911;
assign w34914 = w4070 & ~w34912;
assign w34915 = ~w3957 & w13246;
assign w34916 = w13247 & ~a_29;
assign w34917 = ~w13247 & a_29;
assign w34918 = ~w13179 & w3957;
assign w34919 = w13183 & ~w13170;
assign w34920 = w13183 & w34862;
assign w34921 = ~w13261 & w34890;
assign w34922 = ~w13261 & w34891;
assign w34923 = w13244 & ~w34921;
assign w34924 = w13244 & ~w34922;
assign w34925 = ~w13244 & w34921;
assign w34926 = ~w13244 & w34922;
assign w34927 = ~w4070 & w13266;
assign w34928 = a_29 & ~w13266;
assign w34929 = a_29 & ~w34927;
assign w34930 = ~w13269 & ~w13218;
assign w34931 = ~w13148 & ~w13029;
assign w34932 = w13269 & w13218;
assign w34933 = ~w13274 & ~w13270;
assign w34934 = ~w13129 & ~w13116;
assign w34935 = ~w13129 & w34835;
assign w34936 = ~w12606 & w1327;
assign w34937 = w12614 & w1399;
assign w34938 = ~w12945 & w13285;
assign w34939 = w12945 & ~w13285;
assign w34940 = ~w1478 & w13290;
assign w34941 = ~w13012 & w4446;
assign w34942 = ~w4070 & w13299;
assign w34943 = ~a_29 & w13299;
assign w34944 = ~a_29 & w34942;
assign w34945 = w13292 & w13306;
assign w34946 = ~w13292 & ~w13306;
assign w34947 = ~w13179 & w4446;
assign w34948 = ~w13012 & w4068;
assign w34949 = ~w13237 & w4070;
assign w34950 = ~w13312 & ~w13310;
assign w34951 = ~w13314 & a_29;
assign w34952 = w13314 & ~a_29;
assign w34953 = ~w13317 & ~w13307;
assign w34954 = ~w518 & ~w34919;
assign w34955 = ~w518 & ~w34920;
assign w34956 = w3890 & ~w34954;
assign w34957 = w3890 & ~w34955;
assign w34958 = a_26 & ~w34956;
assign w34959 = a_26 & ~w34957;
assign w34960 = ~w13328 & ~w13322;
assign w34961 = ~w13118 & w13125;
assign w34962 = ~w13118 & w34834;
assign w34963 = w12610 & w668;
assign w34964 = ~w12915 & w1399;
assign w34965 = w12611 & w1327;
assign w34966 = ~w12934 & ~w34779;
assign w34967 = ~w12934 & ~w34780;
assign w34968 = ~w1478 & w13377;
assign w34969 = ~w13367 & ~w13365;
assign w34970 = ~w13381 & ~w13365;
assign w34971 = ~w13381 & w34969;
assign w34972 = w13381 & w13365;
assign w34973 = w13381 & ~w34969;
assign w34974 = w12614 & w668;
assign w34975 = w12610 & w1327;
assign w34976 = w12611 & w1399;
assign w34977 = w12936 & ~w12938;
assign w34978 = ~w1478 & w13391;
assign w34979 = ~w13392 & ~w13382;
assign w34980 = ~w4070 & w13402;
assign w34981 = a_29 & ~w13402;
assign w34982 = a_29 & ~w34980;
assign w34983 = ~w13406 & ~w13395;
assign w34984 = ~w13179 & ~w518;
assign w34985 = w4666 & ~w34919;
assign w34986 = w4666 & ~w34920;
assign w34987 = ~w1226 & w13418;
assign w34988 = ~a_26 & w13418;
assign w34989 = ~a_26 & w34987;
assign w34990 = ~w13422 & ~w13411;
assign w34991 = w4638 & ~w34919;
assign w34992 = w4638 & ~w34920;
assign w34993 = w1226 & ~w34911;
assign w34994 = w1226 & ~w34912;
assign w34995 = ~w4666 & ~w34991;
assign w34996 = ~w4666 & ~w34992;
assign w34997 = ~w13428 & a_26;
assign w34998 = w13428 & ~a_26;
assign w34999 = ~w13434 & ~w13432;
assign w35000 = ~a_17 & ~w13488;
assign w35001 = w13489 & ~w13486;
assign w35002 = w12611 & w668;
assign w35003 = ~w12915 & w1327;
assign w35004 = ~w12922 & ~w12921;
assign w35005 = ~w12922 & ~w34773;
assign w35006 = ~w12929 & w1478;
assign w35007 = ~w13504 & w13496;
assign w35008 = ~w13494 & ~w13496;
assign w35009 = ~w13494 & ~w35007;
assign w35010 = ~w13367 & w13377;
assign w35011 = ~w13367 & w34968;
assign w35012 = ~w13507 & ~w13506;
assign w35013 = w13507 & w13506;
assign w35014 = ~w12915 & w668;
assign w35015 = w12577 & w1399;
assign w35016 = w12911 & w12920;
assign w35017 = ~w13516 & ~w12920;
assign w35018 = ~w13516 & ~w35016;
assign w35019 = w13519 & w1478;
assign w35020 = ~w13522 & w13512;
assign w35021 = ~a_14 & ~w13585;
assign w35022 = w13586 & ~w13583;
assign w35023 = w12577 & w668;
assign w35024 = ~w12893 & w1327;
assign w35025 = ~w12897 & ~w34758;
assign w35026 = ~w12897 & ~w34759;
assign w35027 = ~w12904 & w1478;
assign w35028 = ~w13601 & w13593;
assign w35029 = ~w13591 & ~w13593;
assign w35030 = ~w13591 & ~w35028;
assign w35031 = w13604 & ~w35029;
assign w35032 = w13604 & ~w35030;
assign w35033 = ~w13546 & ~w35031;
assign w35034 = ~w13546 & ~w35032;
assign w35035 = w13522 & ~w13512;
assign w35036 = w13606 & ~w13523;
assign w35037 = w13504 & ~w13496;
assign w35038 = w12614 & w4068;
assign w35039 = w12610 & w3957;
assign w35040 = ~w12606 & w4446;
assign w35041 = ~w4070 & w13620;
assign w35042 = ~a_29 & w13620;
assign w35043 = ~a_29 & w35041;
assign w35044 = ~w13624 & ~w13613;
assign w35045 = ~w13510 & ~w13508;
assign w35046 = w13447 & ~w13508;
assign w35047 = w13447 & w35045;
assign w35048 = ~w13447 & w13508;
assign w35049 = ~w13447 & ~w35045;
assign w35050 = ~w12606 & w3957;
assign w35051 = ~w4070 & w13635;
assign w35052 = a_29 & ~w13635;
assign w35053 = a_29 & ~w35051;
assign w35054 = w13639 & ~w13628;
assign w35055 = ~w13012 & ~w518;
assign w35056 = ~w13179 & w4638;
assign w35057 = ~w1226 & w13649;
assign w35058 = a_26 & ~w13649;
assign w35059 = a_26 & ~w35057;
assign w35060 = w13653 & ~w13642;
assign w35061 = ~w13658 & ~w13656;
assign w35062 = ~w13179 & w4666;
assign w35063 = ~w13012 & w4638;
assign w35064 = ~w13237 & w1226;
assign w35065 = ~w13675 & ~w13674;
assign w35066 = w13678 & a_26;
assign w35067 = ~w13678 & ~a_26;
assign w35068 = ~w12606 & w4068;
assign w35069 = w12614 & w3957;
assign w35070 = ~w4070 & w13689;
assign w35071 = a_29 & ~w13689;
assign w35072 = a_29 & ~w35070;
assign w35073 = ~w13012 & w4666;
assign w35074 = ~w1226 & w13701;
assign w35075 = a_26 & ~w13701;
assign w35076 = a_26 & ~w35074;
assign w35077 = ~w13705 & ~w13694;
assign w35078 = w13707 & ~w13682;
assign w35079 = a_22 & ~w34919;
assign w35080 = a_22 & ~w34920;
assign w35081 = a_23 & w34919;
assign w35082 = a_23 & w34920;
assign w35083 = w508 & ~w35079;
assign w35084 = w508 & ~w35080;
assign w35085 = w13718 & ~w13712;
assign w35086 = w13601 & ~w13593;
assign w35087 = ~w34735 & w12885;
assign w35088 = w12888 & w13767;
assign w35089 = ~w12888 & ~w13767;
assign w35090 = ~w1478 & w13773;
assign w35091 = ~w13763 & ~w13761;
assign w35092 = ~w13777 & ~w13761;
assign w35093 = ~w13777 & w35091;
assign w35094 = w13777 & w13761;
assign w35095 = w13777 & ~w35091;
assign w35096 = ~w12893 & w668;
assign w35097 = w12889 & ~w12886;
assign w35098 = w12889 & ~w34751;
assign w35099 = w13784 & ~w35097;
assign w35100 = w13784 & ~w35098;
assign w35101 = ~w13784 & w35097;
assign w35102 = ~w13784 & w35098;
assign w35103 = ~w1478 & w13789;
assign w35104 = ~w13790 & ~w13778;
assign w35105 = w12611 & w4446;
assign w35106 = ~w12915 & w4068;
assign w35107 = ~w12929 & w4070;
assign w35108 = w13801 & ~a_29;
assign w35109 = ~w13801 & a_29;
assign w35110 = ~w13804 & ~w13793;
assign w35111 = ~w13604 & w35029;
assign w35112 = ~w13604 & w35030;
assign w35113 = w12577 & w1327;
assign w35114 = ~w12893 & w1399;
assign w35115 = w12919 & w13812;
assign w35116 = ~w12919 & ~w13812;
assign w35117 = ~w13811 & ~w13809;
assign w35118 = w12610 & w4446;
assign w35119 = ~w12915 & w3957;
assign w35120 = w12611 & w4068;
assign w35121 = ~w4070 & w13826;
assign w35122 = a_29 & ~w13826;
assign w35123 = a_29 & ~w35121;
assign w35124 = w12614 & ~w518;
assign w35125 = ~w12606 & w4638;
assign w35126 = ~w1226 & w13841;
assign w35127 = ~a_26 & w13841;
assign w35128 = ~a_26 & w35126;
assign w35129 = ~w13845 & ~w13834;
assign w35130 = w12614 & w4446;
assign w35131 = w12610 & w4068;
assign w35132 = w12611 & w3957;
assign w35133 = ~w4070 & w13858;
assign w35134 = a_29 & ~w13858;
assign w35135 = a_29 & ~w35133;
assign w35136 = ~w12606 & ~w518;
assign w35137 = ~w1226 & w13870;
assign w35138 = ~a_26 & ~w13870;
assign w35139 = ~a_26 & ~w35137;
assign w35140 = ~w13179 & w5286;
assign w35141 = ~w13012 & w5080;
assign w35142 = ~w13237 & w5017;
assign w35143 = ~w13882 & ~w13881;
assign w35144 = w13885 & a_23;
assign w35145 = ~w13885 & ~a_23;
assign w35146 = ~w12915 & w4446;
assign w35147 = w12577 & w3957;
assign w35148 = w13519 & w4070;
assign w35149 = ~w13897 & a_29;
assign w35150 = w13897 & ~a_29;
assign w35151 = ~a_11 & ~w13947;
assign w35152 = w13948 & ~w13945;
assign w35153 = ~w12859 & ~w12866;
assign w35154 = w12859 & w12866;
assign w35155 = ~w12865 & ~w13961;
assign w35156 = ~w12869 & w12884;
assign w35157 = w13963 & w13961;
assign w35158 = w13963 & ~w35155;
assign w35159 = ~w13958 & ~w13956;
assign w35160 = ~w13967 & w13955;
assign w35161 = ~w13953 & ~w13955;
assign w35162 = ~w13953 & ~w35160;
assign w35163 = ~w13763 & w13773;
assign w35164 = ~w13763 & w35090;
assign w35165 = ~w13970 & ~w13969;
assign w35166 = w13970 & w13969;
assign w35167 = w12865 & w13961;
assign w35168 = ~w1327 & ~w13976;
assign w35169 = ~w1478 & w13981;
assign w35170 = ~w562 & ~w710;
assign w35171 = w3170 & w14030;
assign w35172 = ~a_8 & ~w14078;
assign w35173 = w14079 & ~w14076;
assign w35174 = ~w12853 & w12631;
assign w35175 = ~w12853 & ~w31782;
assign w35176 = ~w1478 & w14093;
assign w35177 = ~w14086 & ~w14084;
assign w35178 = w14097 & w14084;
assign w35179 = w14097 & ~w35177;
assign w35180 = ~w14019 & ~w35178;
assign w35181 = ~w14019 & ~w35179;
assign w35182 = ~w13975 & w13981;
assign w35183 = ~w13975 & w35169;
assign w35184 = ~w14100 & ~w14099;
assign w35185 = w13967 & ~w13955;
assign w35186 = w12577 & w4446;
assign w35187 = ~w12893 & w4068;
assign w35188 = ~w12904 & w4070;
assign w35189 = w14113 & ~a_29;
assign w35190 = ~w14113 & a_29;
assign w35191 = ~w14116 & ~w14105;
assign w35192 = ~w13973 & ~w13971;
assign w35193 = ~w12606 & w4666;
assign w35194 = w12610 & ~w518;
assign w35195 = w12614 & w4638;
assign w35196 = ~w1226 & w14134;
assign w35197 = ~a_26 & w14134;
assign w35198 = ~a_26 & w35196;
assign w35199 = ~w14138 & ~w14127;
assign w35200 = ~w13012 & w5286;
assign w35201 = ~w5017 & w14150;
assign w35202 = a_23 & ~w14150;
assign w35203 = a_23 & ~w35201;
assign w35204 = ~w14154 & ~w14143;
assign w35205 = w14156 & ~w13889;
assign w35206 = w13847 & ~w13875;
assign w35207 = ~w13862 & ~w13852;
assign w35208 = ~w1226 & w14172;
assign w35209 = a_26 & ~w14172;
assign w35210 = a_26 & ~w35208;
assign w35211 = ~w13012 & w5016;
assign w35212 = ~w13179 & w5080;
assign w35213 = ~w5017 & w14187;
assign w35214 = a_23 & ~w14187;
assign w35215 = a_23 & ~w35213;
assign w35216 = a_19 & ~w34919;
assign w35217 = a_19 & ~w34920;
assign w35218 = a_20 & w34919;
assign w35219 = a_20 & w34920;
assign w35220 = w5304 & ~w35216;
assign w35221 = w5304 & ~w35217;
assign w35222 = ~w14201 & ~w14195;
assign w35223 = ~w14191 & ~w14180;
assign w35224 = ~w14176 & ~w14166;
assign w35225 = ~w13179 & w5016;
assign w35226 = w5286 & ~w34919;
assign w35227 = w5286 & ~w34920;
assign w35228 = ~w5017 & w14218;
assign w35229 = a_23 & ~w14218;
assign w35230 = a_23 & ~w35228;
assign w35231 = w12614 & w4666;
assign w35232 = w12611 & ~w518;
assign w35233 = w12610 & w4638;
assign w35234 = ~w1226 & w14236;
assign w35235 = ~a_26 & w14236;
assign w35236 = ~a_26 & w35234;
assign w35237 = w12577 & w4068;
assign w35238 = ~w12893 & w3957;
assign w35239 = ~w14246 & ~w14244;
assign w35240 = w14248 & ~a_29;
assign w35241 = ~w14248 & a_29;
assign w35242 = w12610 & w4666;
assign w35243 = ~w12915 & ~w518;
assign w35244 = w12611 & w4638;
assign w35245 = ~w1226 & w14259;
assign w35246 = ~a_26 & w14259;
assign w35247 = ~a_26 & w35245;
assign w35248 = ~w14263 & ~w14252;
assign w35249 = ~w5017 & w14279;
assign w35250 = a_23 & ~w14279;
assign w35251 = a_23 & ~w35249;
assign w35252 = ~w14283 & ~w14272;
assign w35253 = ~w13179 & w5308;
assign w35254 = w5816 & ~w34919;
assign w35255 = w5816 & ~w34920;
assign w35256 = ~w5309 & w14295;
assign w35257 = ~a_20 & w14295;
assign w35258 = ~a_20 & w35256;
assign w35259 = ~w14299 & ~w14288;
assign w35260 = w5818 & ~w34919;
assign w35261 = w5818 & ~w34920;
assign w35262 = w5309 & ~w34911;
assign w35263 = w5309 & ~w34912;
assign w35264 = ~w5816 & ~w35260;
assign w35265 = ~w5816 & ~w35261;
assign w35266 = ~w14305 & a_20;
assign w35267 = w14305 & ~a_20;
assign w35268 = ~w14311 & ~w14309;
assign w35269 = ~w14320 & ~w14229;
assign w35270 = ~w429 & ~w249;
assign w35271 = ~a_5 & ~w14378;
assign w35272 = w14379 & ~w14376;
assign w35273 = ~w12663 & ~w12670;
assign w35274 = ~w14390 & ~w12673;
assign w35275 = ~w1478 & w14395;
assign w35276 = ~w14386 & ~w14384;
assign w35277 = w14399 & w14384;
assign w35278 = w14399 & ~w35276;
assign w35279 = ~w14338 & ~w35277;
assign w35280 = ~w14338 & ~w35278;
assign w35281 = w14402 & ~w35279;
assign w35282 = w14402 & ~w35280;
assign w35283 = ~w14402 & w35279;
assign w35284 = ~w14402 & w35280;
assign w35285 = w12846 & w14409;
assign w35286 = ~w12846 & ~w14409;
assign w35287 = ~w1478 & w14414;
assign w35288 = w14415 & ~w14403;
assign w35289 = ~w14086 & w14093;
assign w35290 = ~w14086 & w35176;
assign w35291 = ~w14425 & ~w14423;
assign w35292 = w14427 & ~a_29;
assign w35293 = ~w14427 & a_29;
assign w35294 = ~w14430 & ~w14420;
assign w35295 = ~w14097 & ~w14084;
assign w35296 = ~w14097 & w35177;
assign w35297 = ~w12863 & ~w34720;
assign w35298 = ~w12863 & ~w34721;
assign w35299 = ~w1478 & w14444;
assign w35300 = ~w4070 & w14453;
assign w35301 = ~a_29 & w14453;
assign w35302 = ~a_29 & w35300;
assign w35303 = w12577 & w4638;
assign w35304 = ~w12893 & ~w518;
assign w35305 = ~w14466 & ~w14464;
assign w35306 = w14468 & ~a_26;
assign w35307 = ~w14468 & a_26;
assign w35308 = ~w14471 & ~w14461;
assign w35309 = w14100 & w14099;
assign w35310 = w14446 & w14475;
assign w35311 = ~w14446 & ~w14475;
assign w35312 = ~w12893 & w4446;
assign w35313 = ~w4070 & w14483;
assign w35314 = a_29 & ~w14483;
assign w35315 = a_29 & ~w35313;
assign w35316 = ~w12915 & w4666;
assign w35317 = w12577 & ~w518;
assign w35318 = w13519 & w1226;
assign w35319 = w14496 & ~a_26;
assign w35320 = ~w14496 & a_26;
assign w35321 = w12614 & w5286;
assign w35322 = w12610 & w5080;
assign w35323 = w12611 & w5016;
assign w35324 = ~w5017 & w14510;
assign w35325 = ~a_23 & w14510;
assign w35326 = ~a_23 & w35324;
assign w35327 = ~w4068 & ~w14518;
assign w35328 = ~w4070 & w14521;
assign w35329 = ~a_29 & w14521;
assign w35330 = ~a_29 & w35328;
assign w35331 = ~w14399 & ~w14384;
assign w35332 = ~w14399 & w35276;
assign w35333 = w12844 & ~w14532;
assign w35334 = ~w12844 & w14532;
assign w35335 = ~w1478 & w14537;
assign w35336 = ~w14386 & w14395;
assign w35337 = ~w14386 & w35275;
assign w35338 = w14582 & w14596;
assign w35339 = w14597 & ~w14339;
assign w35340 = ~w14597 & w14339;
assign w35341 = w14612 & w14619;
assign w35342 = w14612 & w31784;
assign w35343 = ~w14610 & ~w35341;
assign w35344 = ~w14610 & ~w35342;
assign w35345 = ~w14623 & ~w14575;
assign w35346 = w14559 & ~w14575;
assign w35347 = w14559 & w35345;
assign w35348 = ~w14557 & ~w35346;
assign w35349 = ~w14557 & ~w35347;
assign w35350 = w14627 & ~w35348;
assign w35351 = w14627 & ~w35349;
assign w35352 = ~w14627 & w35348;
assign w35353 = ~w14627 & w35349;
assign w35354 = ~w14638 & ~w14639;
assign w35355 = ~w1478 & w14643;
assign w35356 = ~w4070 & w14653;
assign w35357 = a_29 & ~w14653;
assign w35358 = a_29 & ~w35356;
assign w35359 = ~w14541 & ~w14539;
assign w35360 = w12577 & w4666;
assign w35361 = ~w12893 & w4638;
assign w35362 = ~w12904 & w1226;
assign w35363 = w14676 & ~a_26;
assign w35364 = ~w14676 & a_26;
assign w35365 = ~w14679 & ~w14668;
assign w35366 = w12610 & w5286;
assign w35367 = ~w12915 & w5016;
assign w35368 = w12611 & w5080;
assign w35369 = ~w5017 & w14691;
assign w35370 = ~a_23 & ~w14691;
assign w35371 = ~a_23 & ~w35369;
assign w35372 = w14695 & ~w14684;
assign w35373 = w14697 & ~w14515;
assign w35374 = w14473 & ~w14500;
assign w35375 = ~w14487 & ~w14476;
assign w35376 = w12611 & w4666;
assign w35377 = ~w12915 & w4638;
assign w35378 = ~w12929 & w1226;
assign w35379 = ~w14714 & a_26;
assign w35380 = w14714 & ~a_26;
assign w35381 = w12614 & w5080;
assign w35382 = w12610 & w5016;
assign w35383 = ~w12606 & w5286;
assign w35384 = ~w5017 & w14728;
assign w35385 = a_23 & ~w14728;
assign w35386 = a_23 & ~w35384;
assign w35387 = ~w5309 & w14743;
assign w35388 = ~a_20 & w14743;
assign w35389 = ~a_20 & w35387;
assign w35390 = ~w14747 & ~w14736;
assign w35391 = ~w14732 & ~w14722;
assign w35392 = ~w14717 & ~w14706;
assign w35393 = w12614 & w5016;
assign w35394 = ~w12606 & w5080;
assign w35395 = ~w5017 & w14761;
assign w35396 = a_23 & ~w14761;
assign w35397 = a_23 & ~w35395;
assign w35398 = ~w13012 & w5816;
assign w35399 = ~w5309 & w14776;
assign w35400 = a_20 & ~w14776;
assign w35401 = a_20 & ~w35399;
assign w35402 = ~w13179 & w6059;
assign w35403 = w6304 & ~w34919;
assign w35404 = w6304 & ~w34920;
assign w35405 = ~w6063 & w14791;
assign w35406 = a_17 & ~w14791;
assign w35407 = a_17 & ~w35405;
assign w35408 = ~w14795 & ~w14784;
assign w35409 = w6061 & ~w34919;
assign w35410 = w6061 & ~w34920;
assign w35411 = w6063 & ~w34911;
assign w35412 = w6063 & ~w34912;
assign w35413 = ~w6304 & ~w35409;
assign w35414 = ~w6304 & ~w35410;
assign w35415 = ~w14801 & a_17;
assign w35416 = w14801 & ~a_17;
assign w35417 = ~w14780 & ~w14770;
assign w35418 = ~w14765 & ~w14754;
assign w35419 = ~w12606 & w5016;
assign w35420 = ~w5017 & w14814;
assign w35421 = ~a_23 & ~w14814;
assign w35422 = ~a_23 & ~w35420;
assign w35423 = ~w13179 & w5816;
assign w35424 = ~w13012 & w5818;
assign w35425 = ~w13237 & w5309;
assign w35426 = ~w14827 & ~w14825;
assign w35427 = ~w14829 & a_20;
assign w35428 = w14829 & ~a_20;
assign w35429 = ~w14838 & ~w14805;
assign w35430 = ~w13179 & w5818;
assign w35431 = ~w13012 & w5308;
assign w35432 = ~w5309 & w14854;
assign w35433 = ~a_20 & w14854;
assign w35434 = ~a_20 & w35432;
assign w35435 = a_16 & ~w34919;
assign w35436 = a_16 & ~w34920;
assign w35437 = a_17 & w34919;
assign w35438 = a_17 & w34920;
assign w35439 = w6058 & ~w35435;
assign w35440 = w6058 & ~w35436;
assign w35441 = ~w14858 & ~w14847;
assign w35442 = ~w14878 & ~w14874;
assign w35443 = ~w14868 & ~w14862;
assign w35444 = ~w12893 & w4666;
assign w35445 = ~w1226 & w14898;
assign w35446 = ~a_26 & w14898;
assign w35447 = ~a_26 & w35445;
assign w35448 = ~w4070 & w14910;
assign w35449 = ~a_29 & w14910;
assign w35450 = ~a_29 & w35448;
assign w35451 = ~w1226 & w14922;
assign w35452 = a_26 & ~w14922;
assign w35453 = a_26 & ~w35451;
assign w35454 = ~w14926 & ~w14915;
assign w35455 = w12611 & w5286;
assign w35456 = ~w12915 & w5080;
assign w35457 = ~w12929 & w5017;
assign w35458 = w14943 & a_23;
assign w35459 = ~w14943 & ~a_23;
assign w35460 = w14946 & ~w14935;
assign w35461 = ~w12606 & w5818;
assign w35462 = w12614 & w5308;
assign w35463 = ~w5309 & w14958;
assign w35464 = ~a_20 & w14958;
assign w35465 = ~a_20 & w35463;
assign w35466 = ~w14962 & ~w14951;
assign w35467 = ~w12606 & w5308;
assign w35468 = ~w5309 & w14971;
assign w35469 = a_20 & ~w14971;
assign w35470 = a_20 & ~w35468;
assign w35471 = ~w13179 & w6304;
assign w35472 = ~w13012 & w6061;
assign w35473 = ~w13237 & w6063;
assign w35474 = ~w14984 & ~w14982;
assign w35475 = ~w14986 & a_17;
assign w35476 = w14986 & ~a_17;
assign w35477 = ~w12915 & w5286;
assign w35478 = w12577 & w5016;
assign w35479 = w13519 & w5017;
assign w35480 = ~w14998 & a_23;
assign w35481 = w14998 & ~a_23;
assign w35482 = ~w4070 & w15009;
assign w35483 = ~a_29 & w15009;
assign w35484 = ~a_29 & w35482;
assign w35485 = ~w14559 & w14575;
assign w35486 = ~w14559 & ~w35345;
assign w35487 = ~w12658 & ~w12649;
assign w35488 = w12658 & w12649;
assign w35489 = ~w15021 & ~w15023;
assign w35490 = w12657 & ~w12831;
assign w35491 = w12657 & w12800;
assign w35492 = w12651 & ~w12826;
assign w35493 = ~w15039 & w1478;
assign w35494 = ~w1399 & ~w15036;
assign w35495 = ~w14612 & ~w14619;
assign w35496 = ~w14612 & ~w31784;
assign w35497 = w15058 & ~w4070;
assign w35498 = w15058 & w14640;
assign w35499 = ~w12781 & ~w12820;
assign w35500 = ~w12794 & ~w15064;
assign w35501 = w12794 & w15064;
assign w35502 = ~w1478 & w15076;
assign w35503 = w15096 & w15076;
assign w35504 = w15096 & w35502;
assign w35505 = ~w12781 & ~w15098;
assign w35506 = w12781 & w15098;
assign w35507 = ~w12764 & w1399;
assign w35508 = ~w1478 & w15106;
assign w35509 = w15119 & w15106;
assign w35510 = w15119 & w35508;
assign w35511 = ~w12764 & w1327;
assign w35512 = ~w15131 & ~w15132;
assign w35513 = ~w15133 & ~w15145;
assign w35514 = w15133 & w15145;
assign w35515 = ~w1478 & w15162;
assign w35516 = w15198 & w15162;
assign w35517 = w15198 & w35515;
assign w35518 = ~w1327 & ~w15201;
assign w35519 = ~w15200 & w15206;
assign w35520 = ~w15275 & ~w15271;
assign w35521 = ~w15279 & ~w15276;
assign w35522 = w15275 & w15271;
assign w35523 = ~w15198 & ~w15162;
assign w35524 = ~w15198 & ~w35515;
assign w35525 = ~w12764 & w668;
assign w35526 = w15429 & ~w15426;
assign w35527 = ~w15436 & ~w15431;
assign w35528 = ~w15429 & w15426;
assign w35529 = ~w15438 & ~w15441;
assign w35530 = ~w15119 & ~w15106;
assign w35531 = ~w15119 & ~w35508;
assign w35532 = ~w15445 & ~w15120;
assign w35533 = ~w15448 & ~w15097;
assign w35534 = w15450 & ~w15063;
assign w35535 = w15051 & ~w15050;
assign w35536 = ~w15033 & ~w15031;
assign w35537 = w15458 & w15031;
assign w35538 = w15458 & ~w35536;
assign w35539 = ~w15018 & ~w15463;
assign w35540 = w15018 & w15463;
assign w35541 = ~w15468 & ~w15467;
assign w35542 = w15471 & a_26;
assign w35543 = ~w15471 & ~a_26;
assign w35544 = ~w15474 & ~w15464;
assign w35545 = w12577 & w5080;
assign w35546 = ~w12893 & w5016;
assign w35547 = ~w15481 & ~w15480;
assign w35548 = w15484 & ~a_23;
assign w35549 = ~w15484 & a_23;
assign w35550 = ~w15487 & ~w15477;
assign w35551 = ~w12606 & w5816;
assign w35552 = w12610 & w5308;
assign w35553 = w12614 & w5818;
assign w35554 = ~w5309 & w15503;
assign w35555 = ~a_20 & w15503;
assign w35556 = ~a_20 & w35554;
assign w35557 = ~w15507 & ~w15496;
assign w35558 = ~w13012 & w6304;
assign w35559 = ~w6063 & w15519;
assign w35560 = a_17 & ~w15519;
assign w35561 = a_17 & ~w35559;
assign w35562 = ~w15523 & ~w15512;
assign w35563 = w15525 & ~w14990;
assign w35564 = w14964 & ~w14976;
assign w35565 = ~w13179 & w6061;
assign w35566 = ~w13012 & w6059;
assign w35567 = ~w6063 & w15540;
assign w35568 = ~a_17 & w15540;
assign w35569 = ~a_17 & w35567;
assign w35570 = a_12 & ~w34919;
assign w35571 = a_12 & ~w34920;
assign w35572 = a_14 & w34919;
assign w35573 = a_14 & w34920;
assign w35574 = w6445 & ~w35570;
assign w35575 = w6445 & ~w35571;
assign w35576 = ~w15554 & ~w15548;
assign w35577 = ~w15544 & ~w15533;
assign w35578 = w12614 & w5816;
assign w35579 = w12610 & w5818;
assign w35580 = w12611 & w5308;
assign w35581 = ~w5309 & w15573;
assign w35582 = ~a_20 & w15573;
assign w35583 = ~a_20 & w35581;
assign w35584 = ~w15458 & ~w15031;
assign w35585 = ~w15458 & w35536;
assign w35586 = ~w4638 & ~w15583;
assign w35587 = ~w1226 & w15586;
assign w35588 = a_26 & ~w15586;
assign w35589 = a_26 & ~w35587;
assign w35590 = ~w15033 & w15050;
assign w35591 = ~w15033 & ~w35535;
assign w35592 = ~w4070 & w15597;
assign w35593 = ~a_29 & ~w15597;
assign w35594 = ~a_29 & ~w35592;
assign w35595 = ~w15592 & ~w15601;
assign w35596 = w15592 & w15601;
assign w35597 = ~w1226 & w15609;
assign w35598 = a_26 & ~w15609;
assign w35599 = a_26 & ~w35597;
assign w35600 = ~w15613 & ~w15602;
assign w35601 = w12577 & w5286;
assign w35602 = ~w12893 & w5080;
assign w35603 = ~w12904 & w5017;
assign w35604 = w15630 & ~a_23;
assign w35605 = ~w15630 & a_23;
assign w35606 = ~w15633 & ~w15622;
assign w35607 = w12610 & w5816;
assign w35608 = ~w12915 & w5308;
assign w35609 = w12611 & w5818;
assign w35610 = ~w5309 & w15643;
assign w35611 = a_20 & ~w15643;
assign w35612 = a_20 & ~w35610;
assign w35613 = ~w15647 & ~w15636;
assign w35614 = ~w6063 & w15663;
assign w35615 = a_17 & ~w15663;
assign w35616 = a_17 & ~w35614;
assign w35617 = ~w15667 & ~w15656;
assign w35618 = ~w13179 & w6446;
assign w35619 = w6996 & ~w34919;
assign w35620 = w6996 & ~w34920;
assign w35621 = ~w6447 & w15679;
assign w35622 = a_14 & ~w15679;
assign w35623 = a_14 & ~w35621;
assign w35624 = ~w15683 & ~w15672;
assign w35625 = w6998 & ~w34919;
assign w35626 = w6998 & ~w34920;
assign w35627 = w6447 & ~w34911;
assign w35628 = w6447 & ~w34912;
assign w35629 = ~w6996 & ~w35625;
assign w35630 = ~w6996 & ~w35626;
assign w35631 = ~w15689 & a_14;
assign w35632 = w15689 & ~a_14;
assign w35633 = ~w15695 & ~w15693;
assign w35634 = ~w12606 & w6059;
assign w35635 = ~w6063 & w15710;
assign w35636 = a_17 & ~w15710;
assign w35637 = a_17 & ~w35635;
assign w35638 = w12611 & w5816;
assign w35639 = ~w12915 & w5818;
assign w35640 = ~w12929 & w5309;
assign w35641 = w15723 & ~a_20;
assign w35642 = ~w15723 & a_20;
assign w35643 = ~w12893 & w5286;
assign w35644 = ~w5017 & w15733;
assign w35645 = ~a_23 & ~w15733;
assign w35646 = ~a_23 & ~w35644;
assign w35647 = ~w1226 & w15744;
assign w35648 = a_26 & ~w15744;
assign w35649 = a_26 & ~w35647;
assign w35650 = ~w4070 & w15754;
assign w35651 = a_29 & ~w15754;
assign w35652 = a_29 & ~w35650;
assign w35653 = ~w5017 & w15772;
assign w35654 = ~a_23 & ~w15772;
assign w35655 = ~a_23 & ~w35653;
assign w35656 = w15738 & w15726;
assign w35657 = ~w15738 & ~w15726;
assign w35658 = ~w12606 & w6061;
assign w35659 = w12614 & w6059;
assign w35660 = ~w6063 & w15799;
assign w35661 = ~a_17 & w15799;
assign w35662 = ~a_17 & w35660;
assign w35663 = w15803 & ~w15792;
assign w35664 = ~w13179 & w6998;
assign w35665 = ~w13012 & w6446;
assign w35666 = ~w6447 & w15819;
assign w35667 = ~a_14 & w15819;
assign w35668 = ~a_14 & w35666;
assign w35669 = ~w15823 & ~w15812;
assign w35670 = ~w15830 & ~w15826;
assign w35671 = ~w1226 & w15859;
assign w35672 = ~a_26 & w15859;
assign w35673 = ~a_26 & w35671;
assign w35674 = ~w15870 & ~w15872;
assign w35675 = w15873 & ~a_29;
assign w35676 = ~w15873 & a_29;
assign w35677 = ~w15039 & w4070;
assign w35678 = ~w3957 & ~w15878;
assign w35679 = w15882 & ~a_29;
assign w35680 = ~w15882 & a_29;
assign w35681 = ~w15146 & ~w15886;
assign w35682 = w15146 & w15886;
assign w35683 = ~w15896 & a_29;
assign w35684 = w15896 & ~a_29;
assign w35685 = ~w7268 & ~w15897;
assign w35686 = ~w12764 & w3957;
assign w35687 = ~w15905 & w15910;
assign w35688 = ~w11501 & w4446;
assign w35689 = ~w3954 & a_29;
assign w35690 = ~w16013 & w16015;
assign w35691 = w16049 & ~a_29;
assign w35692 = ~w12764 & w4446;
assign w35693 = ~w16069 & a_29;
assign w35694 = w15945 & ~w16081;
assign w35695 = ~w16083 & ~w15946;
assign w35696 = w15199 & ~w15413;
assign w35697 = ~w16097 & a_29;
assign w35698 = w16097 & ~a_29;
assign w35699 = w16097 & w7269;
assign w35700 = ~w16111 & ~w15903;
assign w35701 = ~w16114 & ~w15890;
assign w35702 = w16117 & ~w15877;
assign w35703 = w16118 & ~w15864;
assign w35704 = ~w16126 & ~w16124;
assign w35705 = w16128 & ~a_23;
assign w35706 = ~w16128 & a_23;
assign w35707 = ~w16131 & ~w16121;
assign w35708 = ~w12893 & w5308;
assign w35709 = w12577 & w5818;
assign w35710 = ~w16135 & ~w16137;
assign w35711 = ~w8339 & w16140;
assign w35712 = w16146 & ~w16144;
assign w35713 = ~w12915 & w5816;
assign w35714 = w12577 & w5308;
assign w35715 = w13519 & w5309;
assign w35716 = ~w16157 & a_20;
assign w35717 = w16157 & ~a_20;
assign w35718 = ~w15777 & ~w16160;
assign w35719 = w15777 & w16160;
assign w35720 = ~w12606 & w6304;
assign w35721 = w12610 & w6059;
assign w35722 = w12614 & w6061;
assign w35723 = ~w6063 & w16174;
assign w35724 = ~a_17 & w16174;
assign w35725 = ~a_17 & w35723;
assign w35726 = w16187 & a_14;
assign w35727 = ~w16187 & ~a_14;
assign w35728 = ~w8564 & ~w16189;
assign w35729 = w12614 & w6304;
assign w35730 = w12610 & w6061;
assign w35731 = w12611 & w6059;
assign w35732 = ~w6063 & w16201;
assign w35733 = ~a_17 & ~w16201;
assign w35734 = ~a_17 & ~w35732;
assign w35735 = w12610 & w6304;
assign w35736 = ~w12915 & w6059;
assign w35737 = w12611 & w6061;
assign w35738 = ~w6063 & w16214;
assign w35739 = ~a_17 & w16214;
assign w35740 = ~a_17 & w35738;
assign w35741 = w12577 & w5816;
assign w35742 = ~w12893 & w5818;
assign w35743 = ~w12904 & w5309;
assign w35744 = w16227 & ~a_20;
assign w35745 = ~w16227 & a_20;
assign w35746 = ~w1226 & w16242;
assign w35747 = a_26 & ~w16242;
assign w35748 = a_26 & ~w35746;
assign w35749 = w16253 & ~w1226;
assign w35750 = w16253 & w14640;
assign w35751 = w16107 & ~w16109;
assign w35752 = ~a_26 & w16271;
assign w35753 = ~a_26 & w31818;
assign w35754 = a_26 & ~w16271;
assign w35755 = a_26 & ~w31818;
assign w35756 = ~w16078 & ~w16081;
assign w35757 = ~w12764 & ~w518;
assign w35758 = ~w16284 & w16289;
assign w35759 = ~w12732 & w1226;
assign w35760 = ~w12764 & w4666;
assign w35761 = ~w16304 & a_26;
assign w35762 = w16304 & ~a_26;
assign w35763 = w3954 & a_29;
assign w35764 = ~w16013 & ~w16331;
assign w35765 = w16013 & w16331;
assign w35766 = ~w1222 & a_26;
assign w35767 = ~w16381 & ~w16380;
assign w35768 = w16382 & a_26;
assign w35769 = ~w16384 & ~w16011;
assign w35770 = w16392 & ~a_26;
assign w35771 = ~w1226 & w16408;
assign w35772 = ~w12764 & w4638;
assign w35773 = ~w16425 & ~w16426;
assign w35774 = ~w15966 & ~w16445;
assign w35775 = w15966 & w16445;
assign w35776 = w16452 & ~a_26;
assign w35777 = w16452 & w7680;
assign w35778 = ~w16452 & a_26;
assign w35779 = ~w16453 & w16457;
assign w35780 = ~w16465 & ~w16280;
assign w35781 = ~w15039 & w1226;
assign w35782 = w16475 & ~a_26;
assign w35783 = ~w16475 & a_26;
assign w35784 = ~w16484 & ~w16485;
assign w35785 = w16266 & ~w16248;
assign w35786 = ~w1226 & w16520;
assign w35787 = a_26 & ~w16520;
assign w35788 = a_26 & ~w35786;
assign w35789 = w16247 & ~w16530;
assign w35790 = w16532 & w16235;
assign w35791 = ~w16532 & ~w16235;
assign w35792 = ~w5080 & ~w16535;
assign w35793 = ~w5017 & w16538;
assign w35794 = ~a_23 & ~w16538;
assign w35795 = ~a_23 & ~w35793;
assign w35796 = w16544 & ~w16231;
assign w35797 = w16546 & ~w16219;
assign w35798 = w16206 & ~w16194;
assign w35799 = ~w16206 & w16194;
assign w35800 = ~w12606 & w6446;
assign w35801 = ~w6447 & w16562;
assign w35802 = a_14 & ~w16562;
assign w35803 = a_14 & ~w35801;
assign w35804 = ~w12893 & w5816;
assign w35805 = ~w5309 & w16582;
assign w35806 = ~a_20 & w16582;
assign w35807 = ~a_20 & w35805;
assign w35808 = ~w5017 & w16597;
assign w35809 = ~a_23 & w16597;
assign w35810 = ~a_23 & w35808;
assign w35811 = w16618 & ~a_23;
assign w35812 = w16618 & w7962;
assign w35813 = ~w16618 & a_23;
assign w35814 = ~w16619 & w16623;
assign w35815 = ~w12764 & w5016;
assign w35816 = ~w16630 & w16635;
assign w35817 = ~w12732 & w5017;
assign w35818 = ~w16652 & ~a_23;
assign w35819 = w16652 & a_23;
assign w35820 = ~w16382 & a_26;
assign w35821 = ~w5080 & ~w16665;
assign w35822 = ~a_23 & ~w16668;
assign w35823 = a_23 & w16668;
assign w35824 = ~w16670 & ~w16669;
assign w35825 = ~a_23 & w16668;
assign w35826 = a_23 & ~w16668;
assign w35827 = ~w16377 & w16380;
assign w35828 = ~w504 & a_23;
assign w35829 = ~w5017 & w16753;
assign w35830 = ~w12764 & w5080;
assign w35831 = ~w16776 & ~w16777;
assign w35832 = w16774 & a_23;
assign w35833 = ~w16774 & ~a_23;
assign w35834 = w16804 & w7962;
assign w35835 = ~w16804 & a_23;
assign w35836 = w16804 & ~a_23;
assign w35837 = ~w15039 & w7961;
assign w35838 = ~w5016 & ~w16820;
assign w35839 = ~w16821 & w7962;
assign w35840 = w16821 & a_23;
assign w35841 = ~w16821 & ~a_23;
assign w35842 = ~w16854 & ~w16855;
assign w35843 = ~w5017 & w16858;
assign w35844 = ~w16462 & ~w16460;
assign w35845 = w16868 & a_23;
assign w35846 = ~w16868 & ~a_23;
assign w35847 = ~w16868 & w7962;
assign w35848 = ~w5017 & w16895;
assign w35849 = ~a_23 & ~w16895;
assign w35850 = ~a_23 & ~w35848;
assign w35851 = ~w16907 & ~w16479;
assign w35852 = w16913 & a_23;
assign w35853 = ~w16913 & ~a_23;
assign w35854 = ~w7961 & ~w16915;
assign w35855 = w31850 & ~w16920;
assign w35856 = ~w31850 & w16920;
assign w35857 = ~w16935 & ~w16612;
assign w35858 = ~w5017 & w16941;
assign w35859 = a_23 & ~w16941;
assign w35860 = a_23 & ~w35858;
assign w35861 = w16954 & ~w16955;
assign w35862 = ~w5017 & w16961;
assign w35863 = a_23 & ~w16961;
assign w35864 = a_23 & ~w35862;
assign w35865 = ~w16971 & ~w16972;
assign w35866 = w12611 & w6304;
assign w35867 = ~w12915 & w6061;
assign w35868 = ~w12929 & w6063;
assign w35869 = w16985 & ~a_17;
assign w35870 = ~w16985 & a_17;
assign w35871 = ~w16988 & ~w16977;
assign w35872 = ~w12606 & w6998;
assign w35873 = w12614 & w6446;
assign w35874 = ~w6447 & w16998;
assign w35875 = ~a_14 & w16998;
assign w35876 = ~a_14 & w35874;
assign w35877 = w17002 & ~w16991;
assign w35878 = w16572 & ~w16571;
assign w35879 = ~w13179 & w7489;
assign w35880 = ~w13012 & w7192;
assign w35881 = ~w7193 & w17013;
assign w35882 = ~a_11 & ~w17013;
assign w35883 = ~a_11 & ~w35881;
assign w35884 = w17017 & ~w17006;
assign w35885 = ~w15850 & ~w16179;
assign w35886 = ~w13012 & w6996;
assign w35887 = ~w6447 & w17033;
assign w35888 = a_14 & ~w17033;
assign w35889 = a_14 & ~w35887;
assign w35890 = ~w13179 & w7192;
assign w35891 = w7511 & ~w34919;
assign w35892 = w7511 & ~w34920;
assign w35893 = ~w7193 & w17049;
assign w35894 = a_11 & ~w17049;
assign w35895 = a_11 & ~w35893;
assign w35896 = ~w17022 & ~w17020;
assign w35897 = ~w17037 & ~w17026;
assign w35898 = ~w13179 & w6996;
assign w35899 = ~w13012 & w6998;
assign w35900 = ~w13237 & w6447;
assign w35901 = ~w17064 & ~w17062;
assign w35902 = ~w17066 & a_14;
assign w35903 = w17066 & ~a_14;
assign w35904 = w17053 & ~w17043;
assign w35905 = w7489 & ~w34919;
assign w35906 = w7489 & ~w34920;
assign w35907 = w7193 & ~w34911;
assign w35908 = w7193 & ~w34912;
assign w35909 = ~w7511 & ~w35905;
assign w35910 = ~w7511 & ~w35906;
assign w35911 = ~w17080 & a_11;
assign w35912 = w17080 & ~a_11;
assign w35913 = ~w13179 & w7511;
assign w35914 = ~w13012 & w7489;
assign w35915 = ~w13237 & w7193;
assign w35916 = ~w17095 & ~w17093;
assign w35917 = ~w17097 & a_11;
assign w35918 = w17097 & ~a_11;
assign w35919 = ~w12915 & w6304;
assign w35920 = w12577 & w6059;
assign w35921 = w13519 & w6063;
assign w35922 = ~w17114 & a_17;
assign w35923 = w17114 & ~a_17;
assign w35924 = ~w17123 & ~w17121;
assign w35925 = ~w17125 & a_20;
assign w35926 = w17125 & ~a_20;
assign w35927 = ~w5818 & ~w17139;
assign w35928 = ~w5309 & w17142;
assign w35929 = a_20 & ~w17142;
assign w35930 = a_20 & ~w35928;
assign w35931 = ~w16930 & ~w16934;
assign w35932 = ~w16905 & w16926;
assign w35933 = w17160 & a_20;
assign w35934 = ~w17160 & ~a_20;
assign w35935 = ~w8339 & w17163;
assign w35936 = ~w16888 & ~w16890;
assign w35937 = ~w5309 & w17187;
assign w35938 = a_20 & ~w17187;
assign w35939 = a_20 & ~w35937;
assign w35940 = ~w5309 & w17209;
assign w35941 = ~a_20 & w17209;
assign w35942 = ~a_20 & w35940;
assign w35943 = w16888 & ~w17213;
assign w35944 = ~w5309 & w17227;
assign w35945 = a_20 & ~w17227;
assign w35946 = a_20 & ~w35944;
assign w35947 = ~w5309 & w17242;
assign w35948 = ~a_20 & ~w17242;
assign w35949 = ~a_20 & ~w35947;
assign w35950 = w17266 & a_20;
assign w35951 = ~w17266 & ~a_20;
assign w35952 = ~w8339 & w17269;
assign w35953 = ~w12764 & w5308;
assign w35954 = w17278 & ~a_20;
assign w35955 = ~w17278 & a_20;
assign w35956 = ~w8339 & w17282;
assign w35957 = w17288 & ~a_20;
assign w35958 = ~w17288 & a_20;
assign w35959 = ~w17288 & w17294;
assign w35960 = w504 & a_23;
assign w35961 = w17304 & a_23;
assign w35962 = ~w5818 & ~w17310;
assign w35963 = ~w5309 & w17315;
assign w35964 = ~w17317 & ~w17319;
assign w35965 = ~w5309 & w17323;
assign w35966 = ~w17325 & ~w17327;
assign w35967 = ~w5300 & a_20;
assign w35968 = ~w5309 & w17402;
assign w35969 = ~w12764 & w5818;
assign w35970 = ~w17423 & ~w17425;
assign w35971 = ~w17449 & ~a_20;
assign w35972 = w17449 & a_20;
assign w35973 = ~w8339 & w17452;
assign w35974 = ~w15039 & w8311;
assign w35975 = ~w15039 & w8339;
assign w35976 = ~w5308 & ~w17471;
assign w35977 = w17472 & ~a_20;
assign w35978 = ~w17472 & a_20;
assign w35979 = ~w17491 & ~w17492;
assign w35980 = ~w5309 & w17495;
assign w35981 = w35334 & w8339;
assign w35982 = w12844 & w17511;
assign w35983 = w17514 & a_20;
assign w35984 = ~w17514 & ~a_20;
assign w35985 = ~w17518 & ~w17511;
assign w35986 = ~w17518 & ~w35982;
assign w35987 = ~w17138 & w17133;
assign w35988 = ~w5309 & w17551;
assign w35989 = ~a_20 & w17551;
assign w35990 = ~a_20 & w35988;
assign w35991 = ~w17561 & ~w17133;
assign w35992 = ~w17561 & ~w35987;
assign w35993 = w12614 & w6998;
assign w35994 = w12610 & w6446;
assign w35995 = ~w12606 & w6996;
assign w35996 = ~w6447 & w17576;
assign w35997 = ~a_14 & ~w17576;
assign w35998 = ~a_14 & ~w35996;
assign w35999 = ~w17580 & ~w17569;
assign w36000 = ~w13012 & w7511;
assign w36001 = ~w7193 & w17592;
assign w36002 = a_11 & ~w17592;
assign w36003 = a_11 & ~w36001;
assign w36004 = w17596 & ~w17585;
assign w36005 = w17106 & ~w17105;
assign w36006 = a_5 & ~w34919;
assign w36007 = a_5 & ~w34920;
assign w36008 = a_8 & w34919;
assign w36009 = a_8 & w34920;
assign w36010 = w8276 & ~w36006;
assign w36011 = w8276 & ~w36007;
assign w36012 = ~w17606 & ~w17600;
assign w36013 = a_9 & ~w34919;
assign w36014 = a_9 & ~w34920;
assign w36015 = a_11 & w34919;
assign w36016 = a_11 & w34920;
assign w36017 = w7191 & ~w36013;
assign w36018 = w7191 & ~w36014;
assign w36019 = ~w17083 & ~w17075;
assign w36020 = ~w17623 & ~w17618;
assign w36021 = ~w12915 & w8295;
assign w36022 = w12577 & w8277;
assign w36023 = w13519 & w8278;
assign w36024 = w17643 & ~a_8;
assign w36025 = ~w17643 & a_8;
assign w36026 = ~w7193 & w17651;
assign w36027 = ~a_11 & w17651;
assign w36028 = ~a_11 & w36026;
assign w36029 = w17662 & a_17;
assign w36030 = ~w17662 & ~a_17;
assign w36031 = ~w8419 & w17665;
assign w36032 = ~w12764 & w6059;
assign w36033 = w17674 & ~a_17;
assign w36034 = ~w17674 & a_17;
assign w36035 = ~w8419 & w17678;
assign w36036 = w17688 & ~a_17;
assign w36037 = ~w17688 & a_17;
assign w36038 = ~w17688 & w17695;
assign w36039 = w5300 & a_20;
assign w36040 = w17701 & a_20;
assign w36041 = ~w6061 & ~w17707;
assign w36042 = ~w6063 & w17712;
assign w36043 = ~w17714 & ~w17716;
assign w36044 = ~w6063 & w17720;
assign w36045 = ~w17722 & ~w17724;
assign w36046 = ~w6054 & a_17;
assign w36047 = ~w6063 & w17799;
assign w36048 = ~w12764 & w6061;
assign w36049 = ~w17820 & ~w17822;
assign w36050 = ~w17680 & ~w17834;
assign w36051 = ~w17846 & ~a_17;
assign w36052 = w17846 & a_17;
assign w36053 = ~w8419 & w17849;
assign w36054 = ~w17422 & ~w17437;
assign w36055 = ~w15039 & w8391;
assign w36056 = ~w15039 & w8419;
assign w36057 = ~w6059 & ~w17867;
assign w36058 = w17868 & ~a_17;
assign w36059 = ~w17868 & a_17;
assign w36060 = ~w17887 & a_14;
assign w36061 = w17887 & ~a_14;
assign w36062 = ~w8592 & w17891;
assign w36063 = w17901 & a_14;
assign w36064 = ~w17901 & ~a_14;
assign w36065 = ~w8592 & w17904;
assign w36066 = ~w12764 & w6446;
assign w36067 = w17913 & ~a_14;
assign w36068 = ~w17913 & a_14;
assign w36069 = ~w8592 & w17917;
assign w36070 = w17927 & ~a_14;
assign w36071 = ~w17927 & a_14;
assign w36072 = ~w6437 & ~a_14;
assign w36073 = ~w17927 & w17934;
assign w36074 = w6054 & a_17;
assign w36075 = w17940 & a_17;
assign w36076 = ~w6998 & ~w17946;
assign w36077 = ~w6447 & w17951;
assign w36078 = ~w17953 & ~w17955;
assign w36079 = ~w6447 & w17959;
assign w36080 = ~w17961 & ~w17963;
assign w36081 = ~w6441 & a_14;
assign w36082 = ~w6447 & w18038;
assign w36083 = ~w12764 & w6998;
assign w36084 = ~w18059 & ~w18061;
assign w36085 = ~w17919 & ~w18073;
assign w36086 = ~w18085 & ~a_14;
assign w36087 = w18085 & a_14;
assign w36088 = ~w8592 & w18088;
assign w36089 = ~w15039 & w8564;
assign w36090 = ~w15039 & w8592;
assign w36091 = ~w6446 & ~w18106;
assign w36092 = w18107 & ~a_14;
assign w36093 = ~w18107 & a_14;
assign w36094 = ~w18126 & ~w18127;
assign w36095 = ~w8592 & w18131;
assign w36096 = ~w6447 & w18144;
assign w36097 = a_14 & ~w18144;
assign w36098 = a_14 & ~w36096;
assign w36099 = ~w18175 & ~w18176;
assign w36100 = ~w8419 & w18180;
assign w36101 = w18189 & ~a_14;
assign w36102 = ~w18189 & a_14;
assign w36103 = ~w8592 & w18193;
assign w36104 = ~w6063 & w18215;
assign w36105 = a_17 & ~w18215;
assign w36106 = a_17 & ~w36104;
assign w36107 = ~w18229 & a_14;
assign w36108 = w18229 & ~a_14;
assign w36109 = ~w8592 & w18233;
assign w36110 = ~w6447 & w18260;
assign w36111 = ~a_14 & w18260;
assign w36112 = ~a_14 & w36110;
assign w36113 = ~w18268 & a_17;
assign w36114 = w18268 & ~a_17;
assign w36115 = ~w8419 & w18272;
assign w36116 = w18306 & a_14;
assign w36117 = ~w18306 & ~a_14;
assign w36118 = ~w8592 & w18309;
assign w36119 = w35334 & w8419;
assign w36120 = w12844 & w18321;
assign w36121 = w18324 & a_17;
assign w36122 = ~w18324 & ~a_17;
assign w36123 = ~w18328 & ~w18321;
assign w36124 = ~w18328 & ~w36120;
assign w36125 = w18365 & a_11;
assign w36126 = ~w18365 & ~a_11;
assign w36127 = ~w9089 & w18368;
assign w36128 = ~w12764 & w7192;
assign w36129 = w18377 & ~a_11;
assign w36130 = ~w18377 & a_11;
assign w36131 = ~w9089 & w18381;
assign w36132 = w18391 & ~a_11;
assign w36133 = ~w18391 & a_11;
assign w36134 = ~w7183 & ~a_11;
assign w36135 = ~w18391 & w18398;
assign w36136 = w6441 & a_14;
assign w36137 = w18404 & a_14;
assign w36138 = ~w7489 & ~w18410;
assign w36139 = ~w7193 & w18415;
assign w36140 = ~w18417 & ~w18419;
assign w36141 = ~w7193 & w18423;
assign w36142 = ~w18425 & ~w18427;
assign w36143 = ~w7187 & a_11;
assign w36144 = ~w11501 & w7192;
assign w36145 = ~w7193 & w18502;
assign w36146 = ~w12764 & w7489;
assign w36147 = ~w18523 & ~w18525;
assign w36148 = ~w18383 & ~w18537;
assign w36149 = ~w18549 & ~a_11;
assign w36150 = w18549 & a_11;
assign w36151 = ~w9089 & w18552;
assign w36152 = ~w15039 & w9061;
assign w36153 = ~w15039 & w9089;
assign w36154 = ~w7192 & ~w18570;
assign w36155 = w18571 & ~a_11;
assign w36156 = ~w18571 & a_11;
assign w36157 = ~w18590 & ~w18591;
assign w36158 = ~w9089 & w18595;
assign w36159 = ~w7193 & w18608;
assign w36160 = a_11 & ~w18608;
assign w36161 = a_11 & ~w36159;
assign w36162 = ~w18628 & a_11;
assign w36163 = w18628 & ~a_11;
assign w36164 = ~w9089 & w18632;
assign w36165 = w18653 & ~a_11;
assign w36166 = ~w18653 & a_11;
assign w36167 = ~w9089 & w18657;
assign w36168 = w18649 & w18659;
assign w36169 = ~w18674 & a_11;
assign w36170 = w18674 & ~a_11;
assign w36171 = ~w9089 & w18678;
assign w36172 = w18695 & a_11;
assign w36173 = ~w18695 & ~a_11;
assign w36174 = ~w9061 & ~w18697;
assign w36175 = ~w18701 & w17893;
assign w36176 = w18701 & ~w17893;
assign w36177 = w18718 & a_11;
assign w36178 = ~w18718 & ~a_11;
assign w36179 = ~w9089 & w18721;
assign w36180 = ~w7193 & w18762;
assign w36181 = w18763 & w18235;
assign w36182 = ~w18763 & ~w18235;
assign w36183 = ~w18780 & ~w18778;
assign w36184 = ~w18782 & a_11;
assign w36185 = w18782 & ~a_11;
assign w36186 = ~w6063 & w18816;
assign w36187 = ~a_17 & w18816;
assign w36188 = ~a_17 & w36186;
assign w36189 = ~w6998 & ~w18840;
assign w36190 = ~w6447 & w18843;
assign w36191 = ~a_14 & ~w18843;
assign w36192 = ~a_14 & ~w36190;
assign w36193 = ~w12893 & w7511;
assign w36194 = ~w7193 & w18861;
assign w36195 = ~a_11 & w18861;
assign w36196 = ~a_11 & w36194;
assign w36197 = w12577 & w8298;
assign w36198 = ~w12893 & w8277;
assign w36199 = ~w18880 & ~w18879;
assign w36200 = w18883 & ~a_8;
assign w36201 = ~w18883 & a_8;
assign w36202 = ~w8278 & w18893;
assign w36203 = ~a_8 & w18893;
assign w36204 = ~a_8 & w36202;
assign w36205 = ~w12893 & w8295;
assign w36206 = ~w8278 & w18909;
assign w36207 = ~a_8 & w18909;
assign w36208 = ~a_8 & w36206;
assign w36209 = ~w18928 & ~w18926;
assign w36210 = w18930 & ~a_8;
assign w36211 = ~w18930 & a_8;
assign w36212 = w18943 & a_8;
assign w36213 = ~w18943 & ~a_8;
assign w36214 = ~w9484 & w18946;
assign w36215 = ~w8278 & w18964;
assign w36216 = ~a_8 & w18964;
assign w36217 = ~a_8 & w36215;
assign w36218 = ~w18618 & w18624;
assign w36219 = ~w18996 & a_8;
assign w36220 = w18996 & ~a_8;
assign w36221 = ~w9484 & w19000;
assign w36222 = ~w19007 & a_8;
assign w36223 = w19007 & ~a_8;
assign w36224 = ~w9484 & w19011;
assign w36225 = w19031 & a_8;
assign w36226 = ~w19031 & ~a_8;
assign w36227 = ~w9484 & w19034;
assign w36228 = ~w12764 & w8277;
assign w36229 = w19043 & ~a_8;
assign w36230 = ~w19043 & a_8;
assign w36231 = ~w9484 & w19047;
assign w36232 = w19057 & ~a_8;
assign w36233 = ~w19057 & a_8;
assign w36234 = ~w8267 & ~a_8;
assign w36235 = ~w19057 & w19064;
assign w36236 = w7187 & a_11;
assign w36237 = w19070 & a_11;
assign w36238 = ~w8298 & ~w19076;
assign w36239 = ~w8278 & w19081;
assign w36240 = ~w19083 & ~w19085;
assign w36241 = ~w8278 & w19166;
assign w36242 = ~w19168 & ~w19170;
assign w36243 = ~w19172 & w19087;
assign w36244 = ~w8278 & w19178;
assign w36245 = ~w12764 & w8298;
assign w36246 = ~w19049 & ~w19214;
assign w36247 = ~w19226 & ~a_8;
assign w36248 = w19226 & a_8;
assign w36249 = ~w9484 & w19229;
assign w36250 = ~w15039 & w9456;
assign w36251 = ~w15039 & w9484;
assign w36252 = ~w8277 & ~w19247;
assign w36253 = w19248 & ~a_8;
assign w36254 = ~w19248 & a_8;
assign w36255 = ~w19267 & ~w19268;
assign w36256 = ~w9484 & w19272;
assign w36257 = ~w8278 & w19285;
assign w36258 = ~a_8 & w19285;
assign w36259 = ~a_8 & w36257;
assign w36260 = w19310 & ~a_8;
assign w36261 = ~w19310 & a_8;
assign w36262 = ~w9484 & w19314;
assign w36263 = ~w18989 & w19002;
assign w36264 = w18597 & w19316;
assign w36265 = ~w18584 & w19327;
assign w36266 = ~w19332 & ~w19003;
assign w36267 = w18665 & ~w18668;
assign w36268 = ~w8278 & w19351;
assign w36269 = w19352 & w18680;
assign w36270 = ~w19352 & ~w18680;
assign w36271 = w12577 & w8295;
assign w36272 = ~w12893 & w8298;
assign w36273 = ~w12904 & w8278;
assign w36274 = ~w19390 & a_8;
assign w36275 = w19390 & ~a_8;
assign w36276 = w12614 & w9788;
assign w36277 = w12610 & w9780;
assign w36278 = w12611 & w9786;
assign w36279 = ~w9790 & w19419;
assign w36280 = ~a_5 & w19419;
assign w36281 = ~a_5 & w36279;
assign w36282 = w12610 & w9788;
assign w36283 = ~w12915 & w9786;
assign w36284 = w12611 & w9780;
assign w36285 = ~w9790 & w19429;
assign w36286 = ~a_5 & ~w19429;
assign w36287 = ~a_5 & ~w36285;
assign w36288 = ~w12893 & w9788;
assign w36289 = ~w9790 & w19449;
assign w36290 = ~a_5 & w19449;
assign w36291 = ~a_5 & w36289;
assign w36292 = ~w9790 & w19466;
assign w36293 = ~a_5 & ~w19466;
assign w36294 = ~a_5 & ~w36292;
assign w36295 = ~w19487 & ~w19485;
assign w36296 = w19489 & ~a_5;
assign w36297 = ~w19489 & a_5;
assign w36298 = ~w9790 & w19498;
assign w36299 = ~a_5 & w19498;
assign w36300 = ~a_5 & w36298;
assign w36301 = ~w19295 & w19301;
assign w36302 = ~w19514 & ~w19515;
assign w36303 = ~w10061 & w19519;
assign w36304 = w19529 & a_5;
assign w36305 = ~w19529 & ~a_5;
assign w36306 = ~w10061 & w19532;
assign w36307 = ~w12764 & w9786;
assign w36308 = w19541 & ~a_5;
assign w36309 = ~w19541 & a_5;
assign w36310 = ~w10061 & w19545;
assign w36311 = ~w12764 & w9788;
assign w36312 = w19555 & ~a_5;
assign w36313 = ~w19555 & a_5;
assign w36314 = ~w9783 & ~a_5;
assign w36315 = ~w19555 & w19562;
assign w36316 = ~w9780 & ~w19568;
assign w36317 = a_5 & ~w31949;
assign w36318 = w19577 & ~w19573;
assign w36319 = w19577 & ~w31950;
assign w36320 = ~w9790 & w19580;
assign w36321 = ~w19582 & ~w19584;
assign w36322 = w19107 & w19106;
assign w36323 = ~w11501 & w9786;
assign w36324 = ~w9780 & ~w19591;
assign w36325 = ~w9790 & w19594;
assign w36326 = ~w11501 & w9788;
assign w36327 = ~w9776 & a_5;
assign w36328 = ~w19600 & w19607;
assign w36329 = ~w19620 & ~w19588;
assign w36330 = w19620 & w19588;
assign w36331 = w19622 & ~w19621;
assign w36332 = ~w9790 & w19647;
assign w36333 = ~w12764 & w9780;
assign w36334 = ~w19666 & ~w19668;
assign w36335 = ~w19547 & ~w19680;
assign w36336 = ~w19685 & ~w19548;
assign w36337 = ~w19691 & ~a_5;
assign w36338 = w19691 & a_5;
assign w36339 = ~w10061 & w19694;
assign w36340 = ~w15039 & w10033;
assign w36341 = ~w15039 & w10061;
assign w36342 = ~w9786 & ~w19710;
assign w36343 = ~w19711 & a_5;
assign w36344 = w19711 & ~a_5;
assign w36345 = ~w19734 & a_5;
assign w36346 = w19734 & ~a_5;
assign w36347 = ~w10061 & w19738;
assign w36348 = ~w9790 & w19752;
assign w36349 = ~a_5 & w19752;
assign w36350 = ~a_5 & w36348;
assign w36351 = w19782 & ~a_5;
assign w36352 = ~w19782 & a_5;
assign w36353 = ~w10061 & w19786;
assign w36354 = w19801 & ~a_5;
assign w36355 = ~w19801 & a_5;
assign w36356 = ~w10061 & w19805;
assign w36357 = w19274 & w19788;
assign w36358 = ~w19261 & w19814;
assign w36359 = ~w19817 & ~w19821;
assign w36360 = w19830 & a_5;
assign w36361 = ~w19830 & ~a_5;
assign w36362 = ~w10061 & w19833;
assign w36363 = ~w19835 & ~w19507;
assign w36364 = w19322 & w19330;
assign w36365 = ~w9790 & w19848;
assign w36366 = w19849 & w19002;
assign w36367 = ~w19849 & ~w19002;
assign w36368 = w19862 & ~w19493;
assign w36369 = w19365 & ~w19883;
assign w36370 = w12577 & w9788;
assign w36371 = ~w12893 & w9780;
assign w36372 = ~w12904 & w9790;
assign w36373 = w19891 & a_5;
assign w36374 = ~w19891 & ~a_5;
assign w36375 = w12577 & w9780;
assign w36376 = ~w12893 & w9786;
assign w36377 = ~w19903 & ~w19902;
assign w36378 = w19906 & ~a_5;
assign w36379 = ~w19906 & a_5;
assign w36380 = ~w12915 & w9788;
assign w36381 = w12577 & w9786;
assign w36382 = w13519 & w9790;
assign w36383 = w19938 & ~a_5;
assign w36384 = ~w19938 & a_5;
assign w36385 = w12611 & w9788;
assign w36386 = ~w12915 & w9780;
assign w36387 = ~w12929 & w9790;
assign w36388 = w19955 & ~a_5;
assign w36389 = ~w19955 & a_5;
assign w36390 = ~w19991 & ~w19989;
assign w36391 = ~w19993 & a_14;
assign w36392 = w19993 & ~a_14;
assign w36393 = ~w6063 & w20008;
assign w36394 = ~a_17 & w20008;
assign w36395 = ~a_17 & w36393;
assign w36396 = w12577 & w7511;
assign w36397 = ~w12893 & w7489;
assign w36398 = ~w12904 & w7193;
assign w36399 = ~w20035 & a_11;
assign w36400 = w20035 & ~a_11;
assign w36401 = w12611 & w8295;
assign w36402 = ~w12915 & w8298;
assign w36403 = ~w12929 & w8278;
assign w36404 = w20050 & a_8;
assign w36405 = ~w20050 & ~a_8;
assign w36406 = w12610 & w8295;
assign w36407 = ~w12915 & w8277;
assign w36408 = w12611 & w8298;
assign w36409 = ~w8278 & w20080;
assign w36410 = ~a_8 & w20080;
assign w36411 = ~a_8 & w36409;
assign w36412 = w12577 & w7489;
assign w36413 = ~w12893 & w7192;
assign w36414 = ~w20090 & ~w20088;
assign w36415 = ~w20092 & a_11;
assign w36416 = w20092 & ~a_11;
assign w36417 = ~w20108 & ~a_14;
assign w36418 = ~w6447 & w20110;
assign w36419 = w20108 & a_14;
assign w36420 = w20120 & a_17;
assign w36421 = ~w20120 & ~a_17;
assign w36422 = ~w8419 & w20123;
assign w36423 = ~w20111 & ~w20125;
assign w36424 = w20111 & w20125;
assign w36425 = w12614 & w9786;
assign w36426 = ~w12606 & w9780;
assign w36427 = ~w9790 & w20151;
assign w36428 = ~a_5 & ~w20151;
assign w36429 = ~a_5 & ~w36427;
assign w36430 = w12614 & w9780;
assign w36431 = w12610 & w9786;
assign w36432 = ~w12606 & w9788;
assign w36433 = ~w9790 & w20167;
assign w36434 = ~a_5 & ~w20167;
assign w36435 = ~a_5 & ~w36433;
assign w36436 = w12614 & w8295;
assign w36437 = w12610 & w8298;
assign w36438 = w12611 & w8277;
assign w36439 = ~w8278 & w20205;
assign w36440 = ~a_8 & ~w20205;
assign w36441 = ~a_8 & ~w36439;
assign w36442 = ~w6061 & ~w20227;
assign w36443 = ~w6063 & w20230;
assign w36444 = ~a_17 & w20230;
assign w36445 = ~a_17 & w36443;
assign w36446 = ~w12893 & w6996;
assign w36447 = ~w6447 & w20248;
assign w36448 = ~a_14 & w20248;
assign w36449 = ~a_14 & w36447;
assign w36450 = w13519 & w9061;
assign w36451 = w12577 & w7192;
assign w36452 = ~w12915 & w7511;
assign w36453 = w20256 & a_11;
assign w36454 = w13519 & w7193;
assign w36455 = ~w20256 & ~a_11;
assign w36456 = w17538 & w20291;
assign w36457 = ~w20298 & ~w20296;
assign w36458 = w20300 & ~a_17;
assign w36459 = ~w20300 & a_17;
assign w36460 = ~w12904 & w8564;
assign w36461 = ~w12893 & w6998;
assign w36462 = w12577 & w6996;
assign w36463 = w20313 & a_14;
assign w36464 = ~w12904 & w8592;
assign w36465 = ~w20313 & ~a_14;
assign w36466 = ~w12606 & w8295;
assign w36467 = w12610 & w8277;
assign w36468 = w12614 & w8298;
assign w36469 = ~w20329 & ~a_8;
assign w36470 = ~w8278 & w20331;
assign w36471 = w20329 & a_8;
assign w36472 = w12611 & w7511;
assign w36473 = ~w12915 & w7489;
assign w36474 = ~w12929 & w7193;
assign w36475 = w20342 & ~a_11;
assign w36476 = ~w20342 & a_11;
assign w36477 = ~w20286 & w20354;
assign w36478 = w20286 & ~w20354;
assign w36479 = ~w9790 & w20364;
assign w36480 = a_5 & ~w20364;
assign w36481 = a_5 & ~w36479;
assign w36482 = w20285 & w20370;
assign w36483 = ~w12606 & w9786;
assign w36484 = ~w9790 & w20378;
assign w36485 = a_5 & ~w20378;
assign w36486 = a_5 & ~w36484;
assign w36487 = ~w20285 & w20392;
assign w36488 = w20285 & w20394;
assign w36489 = w20402 & ~w20345;
assign w36490 = ~w20263 & ~w20345;
assign w36491 = ~w20402 & ~w20416;
assign w36492 = ~w20422 & ~w20418;
assign w36493 = ~w12893 & w6446;
assign w36494 = ~w6447 & w20428;
assign w36495 = a_14 & ~w20428;
assign w36496 = a_14 & ~w36494;
assign w36497 = w20435 & ~w17202;
assign w36498 = ~w6063 & w20442;
assign w36499 = ~a_17 & w20442;
assign w36500 = ~a_17 & w36498;
assign w36501 = w12610 & w7511;
assign w36502 = ~w12915 & w7192;
assign w36503 = w12611 & w7489;
assign w36504 = ~w7193 & w20468;
assign w36505 = a_11 & ~w20468;
assign w36506 = a_11 & ~w36504;
assign w36507 = ~w13012 & w9788;
assign w36508 = ~w9790 & w20483;
assign w36509 = ~w12606 & w8298;
assign w36510 = w12614 & w8277;
assign w36511 = ~w8278 & w20489;
assign w36512 = ~a_8 & w20489;
assign w36513 = ~a_8 & w36511;
assign w36514 = w20492 & a_5;
assign w36515 = ~w20492 & ~a_5;
assign w36516 = a_5 & ~w20483;
assign w36517 = a_5 & ~w36508;
assign w36518 = ~a_5 & w20483;
assign w36519 = ~a_5 & w36508;
assign w36520 = ~w13179 & w9788;
assign w36521 = ~w13012 & w9780;
assign w36522 = ~w13237 & w9790;
assign w36523 = ~w20523 & ~w20522;
assign w36524 = w20526 & a_5;
assign w36525 = ~w20526 & ~a_5;
assign w36526 = ~w20538 & w20457;
assign w36527 = ~w12893 & w6304;
assign w36528 = ~w6063 & w20550;
assign w36529 = ~a_17 & ~w20550;
assign w36530 = ~a_17 & ~w36528;
assign w36531 = ~w12915 & w6996;
assign w36532 = w12577 & w6446;
assign w36533 = w13519 & w6447;
assign w36534 = w20563 & ~a_14;
assign w36535 = ~w20563 & a_14;
assign w36536 = ~w12606 & w8277;
assign w36537 = ~w8278 & w20583;
assign w36538 = a_8 & ~w20583;
assign w36539 = a_8 & ~w36537;
assign w36540 = w12614 & w7511;
assign w36541 = w12610 & w7489;
assign w36542 = w12611 & w7192;
assign w36543 = ~w7193 & w20592;
assign w36544 = a_11 & ~w20592;
assign w36545 = a_11 & ~w36543;
assign w36546 = w10835 & ~w34919;
assign w36547 = w10835 & ~w34920;
assign w36548 = w10837 & ~w34911;
assign w36549 = w10837 & ~w34912;
assign w36550 = ~w3 & ~w36546;
assign w36551 = ~w3 & ~w36547;
assign w36552 = ~w20613 & a_2;
assign w36553 = w3 & ~w34919;
assign w36554 = w3 & ~w34920;
assign w36555 = ~w10835 & ~w20624;
assign w36556 = ~w13179 & w10839;
assign w36557 = w20626 & ~w20628;
assign w36558 = ~w20626 & a_2;
assign w36559 = ~w10835 & ~w20647;
assign w36560 = ~w20649 & a_2;
assign w36561 = ~w15039 & w10837;
assign w36562 = ~w20659 & a_2;
assign w36563 = ~w19682 & ~w19680;
assign w36564 = ~w3 & ~w20672;
assign w36565 = ~w20674 & ~a_2;
assign w36566 = w20674 & a_2;
assign w36567 = w19642 & ~w19662;
assign w36568 = ~w12764 & w10909;
assign w36569 = ~w10837 & w20691;
assign w36570 = a_2 & w20691;
assign w36571 = a_2 & w36569;
assign w36572 = w20694 & ~w20688;
assign w36573 = ~w12764 & w10835;
assign w36574 = ~w10837 & w20699;
assign w36575 = a_2 & ~w20699;
assign w36576 = a_2 & ~w36574;
assign w36577 = ~w12764 & w3;
assign w36578 = ~w10837 & w20711;
assign w36579 = a_2 & w20711;
assign w36580 = a_2 & w36578;
assign w36581 = w20714 & ~w20708;
assign w36582 = ~w19596 & a_5;
assign w36583 = ~w19619 & w19595;
assign w36584 = w19619 & ~w19595;
assign w36585 = ~w10837 & w20729;
assign w36586 = a_2 & w20729;
assign w36587 = a_2 & w36585;
assign w36588 = w20732 & ~w20726;
assign w36589 = w9776 & a_5;
assign w36590 = ~w19604 & ~w20736;
assign w36591 = w20739 & ~w20738;
assign w36592 = ~w20739 & w20738;
assign w36593 = ~w10837 & w20746;
assign w36594 = a_2 & ~w20746;
assign w36595 = a_2 & ~w36593;
assign w36596 = ~w20749 & w20742;
assign w36597 = w19604 & w20736;
assign w36598 = ~w11501 & w10909;
assign w36599 = ~w10837 & w20756;
assign w36600 = w9776 & ~a_2;
assign w36601 = ~w11501 & a_1;
assign w36602 = ~a_0 & w20764;
assign w36603 = w19602 & ~w20753;
assign w36604 = w20760 & ~w20752;
assign w36605 = ~w20760 & w20752;
assign w36606 = ~w3 & ~w20771;
assign w36607 = ~w20773 & a_2;
assign w36608 = w20773 & ~a_2;
assign w36609 = w20775 & ~w20769;
assign w36610 = w20749 & ~w20742;
assign w36611 = w20720 & w20707;
assign w36612 = w20785 & ~w20707;
assign w36613 = w20785 & ~w36611;
assign w36614 = ~w20720 & ~w20707;
assign w36615 = ~w20654 & ~w20684;
assign w36616 = ~w10837 & w20803;
assign w36617 = a_2 & w20803;
assign w36618 = a_2 & w36616;
assign w36619 = w20806 & ~w20800;
assign w36620 = ~w10837 & w20819;
assign w36621 = a_2 & ~w20819;
assign w36622 = a_2 & ~w36620;
assign w36623 = w20824 & ~w20811;
assign w36624 = ~w10837 & w20832;
assign w36625 = a_2 & ~w20832;
assign w36626 = a_2 & ~w36624;
assign w36627 = ~w10837 & w20849;
assign w36628 = a_2 & ~w20849;
assign w36629 = a_2 & ~w36627;
assign w36630 = w20854 & ~w20841;
assign w36631 = ~w10837 & w20863;
assign w36632 = a_2 & ~w20863;
assign w36633 = a_2 & ~w36631;
assign w36634 = w19762 & ~w19773;
assign w36635 = ~w10837 & w20879;
assign w36636 = a_2 & ~w20879;
assign w36637 = a_2 & ~w36635;
assign w36638 = w20856 & ~w20871;
assign w36639 = ~w3 & ~w20891;
assign w36640 = ~w20893 & a_2;
assign w36641 = ~w20898 & ~w20888;
assign w36642 = w19794 & w19816;
assign w36643 = ~w10837 & w20909;
assign w36644 = a_2 & ~w20909;
assign w36645 = a_2 & ~w36643;
assign w36646 = ~w10837 & w20922;
assign w36647 = a_2 & ~w20922;
assign w36648 = a_2 & ~w36646;
assign w36649 = ~w10837 & w20938;
assign w36650 = a_2 & ~w20938;
assign w36651 = a_2 & ~w36649;
assign w36652 = ~w12893 & w3;
assign w36653 = ~w10837 & w20952;
assign w36654 = a_2 & ~w20952;
assign w36655 = a_2 & ~w36653;
assign w36656 = w12577 & w3;
assign w36657 = ~w12893 & w10835;
assign w36658 = ~w12904 & w10837;
assign w36659 = ~w20970 & a_2;
assign w36660 = w12577 & w10835;
assign w36661 = ~w10837 & w20984;
assign w36662 = a_2 & ~w20984;
assign w36663 = a_2 & ~w36661;
assign w36664 = ~w12915 & w3;
assign w36665 = w13519 & w10837;
assign w36666 = w12577 & w10839;
assign w36667 = w20998 & ~w21000;
assign w36668 = ~w20998 & a_2;
assign w36669 = ~w20994 & ~w21003;
assign w36670 = w12611 & w3;
assign w36671 = ~w12915 & w10835;
assign w36672 = ~w12929 & w10837;
assign w36673 = ~w21016 & a_2;
assign w36674 = w20994 & w21003;
assign w36675 = ~w21021 & ~w21024;
assign w36676 = w12610 & w3;
assign w36677 = w12611 & w10835;
assign w36678 = ~w10837 & w21031;
assign w36679 = a_2 & ~w21031;
assign w36680 = a_2 & ~w36678;
assign w36681 = w12614 & w3;
assign w36682 = w12610 & w10835;
assign w36683 = ~w10837 & w21046;
assign w36684 = a_2 & ~w21046;
assign w36685 = a_2 & ~w36683;
assign w36686 = w12614 & w10835;
assign w36687 = ~w12606 & w3;
assign w36688 = ~w10837 & w21073;
assign w36689 = a_2 & ~w21073;
assign w36690 = a_2 & ~w36688;
assign w36691 = ~w12606 & w10835;
assign w36692 = ~w10837 & w21101;
assign w36693 = a_2 & ~w21101;
assign w36694 = a_2 & ~w36692;
assign w36695 = ~w10837 & w21117;
assign w36696 = a_2 & ~w21117;
assign w36697 = a_2 & ~w36695;
assign w36698 = ~w10837 & w21144;
assign w36699 = a_2 & ~w21144;
assign w36700 = a_2 & ~w36698;
assign w36701 = ~w13012 & w3;
assign w36702 = ~w10837 & w21163;
assign w36703 = a_2 & ~w21163;
assign w36704 = a_2 & ~w36702;
assign w36705 = ~w13179 & w3;
assign w36706 = ~w13012 & w10835;
assign w36707 = ~w13237 & w10837;
assign w36708 = ~w21189 & a_2;
assign w36709 = ~w13179 & w10835;
assign w36710 = ~w10837 & w21213;
assign w36711 = a_2 & ~w21213;
assign w36712 = a_2 & ~w36710;
assign w36713 = w20396 & ~w21218;
assign w36714 = ~w20396 & w21218;
assign w36715 = ~w21206 & ~w21224;
assign w36716 = w10909 & w34919;
assign w36717 = w10909 & w34920;
assign w36718 = ~w14339 & ~w36716;
assign w36719 = ~w14339 & ~w36717;
assign w36720 = ~w31979 & w21268;
assign w36721 = w12611 & w6996;
assign w36722 = ~w12915 & w6998;
assign w36723 = ~w12929 & w6447;
assign w36724 = w21288 & ~a_14;
assign w36725 = ~w21288 & a_14;
assign w36726 = w12577 & w6304;
assign w36727 = ~w12893 & w6061;
assign w36728 = ~w12904 & w6063;
assign w36729 = w21298 & ~a_17;
assign w36730 = ~w21298 & a_17;
assign w36731 = w12614 & w7489;
assign w36732 = w12610 & w7192;
assign w36733 = ~w12606 & w7511;
assign w36734 = ~w7193 & w21323;
assign w36735 = a_11 & ~w21323;
assign w36736 = a_11 & ~w36734;
assign w36737 = ~w8278 & w21341;
assign w36738 = a_8 & ~w21341;
assign w36739 = a_8 & ~w36737;
assign w36740 = ~w13179 & w9780;
assign w36741 = ~w13012 & w9786;
assign w36742 = w21348 & a_5;
assign w36743 = ~w21348 & ~a_5;
assign w36744 = ~w10033 & ~w21350;
assign w36745 = ~w21354 & w21345;
assign w36746 = w21354 & ~w21345;
assign w36747 = w9788 & ~w34919;
assign w36748 = w9788 & ~w34920;
assign w36749 = ~w13179 & w9786;
assign w36750 = ~w10061 & w21394;
assign w36751 = w12610 & w6996;
assign w36752 = ~w12915 & w6446;
assign w36753 = w12611 & w6998;
assign w36754 = ~w6447 & w21409;
assign w36755 = a_14 & ~w21409;
assign w36756 = a_14 & ~w36754;
assign w36757 = w12577 & w6061;
assign w36758 = ~w12893 & w6059;
assign w36759 = ~w21416 & ~w21414;
assign w36760 = w21418 & ~a_17;
assign w36761 = ~w21418 & a_17;
assign w36762 = ~w12606 & w7489;
assign w36763 = w12614 & w7192;
assign w36764 = ~w7193 & w21441;
assign w36765 = ~a_11 & w21441;
assign w36766 = ~a_11 & w36764;
assign w36767 = ~w13012 & w8295;
assign w36768 = ~w8278 & w21450;
assign w36769 = ~a_8 & w21450;
assign w36770 = ~a_8 & w36768;
assign w36771 = w12610 & w6998;
assign w36772 = w12611 & w6446;
assign w36773 = w12614 & w6996;
assign w36774 = ~w8592 & w21498;
assign w36775 = ~w21403 & w21427;
assign w36776 = w21488 & ~w21510;
assign w36777 = ~w21488 & w21510;
assign w36778 = ~w13179 & w8295;
assign w36779 = ~w13012 & w8298;
assign w36780 = ~w13237 & w8278;
assign w36781 = ~w21516 & ~w21514;
assign w36782 = ~w21518 & a_8;
assign w36783 = w21518 & ~a_8;
assign w36784 = ~w12606 & w7192;
assign w36785 = ~w7193 & w21526;
assign w36786 = ~a_11 & w21526;
assign w36787 = ~a_11 & w36785;
assign w36788 = w9780 & ~w34919;
assign w36789 = w9780 & ~w34920;
assign w36790 = w9790 & ~w34911;
assign w36791 = w9790 & ~w34912;
assign w36792 = ~w9788 & ~w36788;
assign w36793 = ~w9788 & ~w36789;
assign w36794 = ~w21543 & a_5;
assign w36795 = w21543 & ~a_5;
assign w36796 = ~w21375 & w21552;
assign w36797 = ~w21504 & ~w21502;
assign w36798 = ~w7193 & w21571;
assign w36799 = ~a_11 & w21571;
assign w36800 = ~a_11 & w36798;
assign w36801 = ~w13179 & w8298;
assign w36802 = ~w13012 & w8277;
assign w36803 = ~w8278 & w21580;
assign w36804 = ~a_8 & w21580;
assign w36805 = ~a_8 & w36803;
assign w36806 = w21583 & w21575;
assign w36807 = ~w21583 & ~w21575;
assign w36808 = ~w21560 & ~w21595;
assign w36809 = w21560 & w21595;
assign w36810 = a_3 & ~w34919;
assign w36811 = a_3 & ~w34920;
assign w36812 = a_5 & w34919;
assign w36813 = a_5 & w34920;
assign w36814 = w9785 & ~w36810;
assign w36815 = w9785 & ~w36811;
assign w36816 = ~w13179 & w8277;
assign w36817 = w8295 & ~w34919;
assign w36818 = w8295 & ~w34920;
assign w36819 = ~w8278 & w21619;
assign w36820 = ~a_8 & w21619;
assign w36821 = ~a_8 & w36819;
assign w36822 = w21627 & w14379;
assign w36823 = ~w21627 & ~w14379;
assign w36824 = w21605 & ~w21635;
assign w36825 = ~w21626 & ~w21628;
assign w36826 = ~w21623 & ~w21613;
assign w36827 = w8298 & ~w34919;
assign w36828 = w8298 & ~w34920;
assign w36829 = w8278 & ~w34911;
assign w36830 = w8278 & ~w34912;
assign w36831 = ~w8295 & ~w36827;
assign w36832 = ~w8295 & ~w36828;
assign w36833 = ~w21649 & a_8;
assign w36834 = w21649 & ~a_8;
assign w36835 = w21657 & ~w21658;
assign w36836 = w21633 & ~w21663;
assign w36837 = w21475 & w21673;
assign w36838 = ~w21669 & ~w21667;
assign w36839 = w17637 & ~w21682;
assign w36840 = (w21687 & w31993) | (w21687 & w21680) | (w31993 & w21680);
assign w36841 = (w21687 & w31993) | (w21687 & w32456) | (w31993 & w32456);
assign w36842 = w15847 & ~w14891;
assign w36843 = ~w15703 & w21689;
assign w36844 = w21692 & ~w21689;
assign w36845 = w21692 & ~w36843;
assign w36846 = ~w21693 & w21700;
assign w36847 = w21701 & ~w36844;
assign w36848 = w21701 & ~w36845;
assign w36849 = ~w14322 & ~w36847;
assign w36850 = ~w14322 & ~w36848;
assign w36851 = ~w14222 & ~w14212;
assign w36852 = w5080 & ~w34919;
assign w36853 = w5080 & ~w34920;
assign w36854 = w5017 & ~w34911;
assign w36855 = w5017 & ~w34912;
assign w36856 = ~w21710 & a_23;
assign w36857 = w21710 & ~a_23;
assign w36858 = ~w21720 & w36849;
assign w36859 = ~w21720 & w36850;
assign w36860 = ~w21704 & ~w21715;
assign w36861 = w21728 & ~w36858;
assign w36862 = w21728 & ~w36859;
assign w36863 = ~w21733 & ~w36861;
assign w36864 = ~w21733 & ~w36862;
assign w36865 = ~w13722 & ~w36863;
assign w36866 = ~w13722 & ~w36864;
assign w36867 = ~w13721 & ~w36865;
assign w36868 = ~w13721 & ~w36866;
assign w36869 = ~w13667 & ~w13665;
assign w36870 = w13443 & w13665;
assign w36871 = w13443 & ~w36869;
assign w36872 = ~w13441 & ~w36870;
assign w36873 = ~w13441 & ~w36871;
assign w36874 = w21739 & ~w36872;
assign w36875 = w21739 & ~w36873;
assign w36876 = ~w13333 & ~w36874;
assign w36877 = ~w13333 & ~w36875;
assign w36878 = ~w13279 & ~w36876;
assign w36879 = ~w13279 & ~w36877;
assign w36880 = w13279 & w36876;
assign w36881 = w13279 & w36877;
assign w36882 = ~w21739 & w36872;
assign w36883 = ~w21739 & w36873;
assign w36884 = ~w13443 & ~w13665;
assign w36885 = ~w13443 & w36869;
assign w36886 = ~w13667 & w36867;
assign w36887 = ~w13667 & w36868;
assign w36888 = w21733 & w36861;
assign w36889 = w21733 & w36862;
assign w36890 = w21697 & ~w36844;
assign w36891 = w21697 & ~w36845;
assign w36892 = w21699 & w36890;
assign w36893 = w21699 & w36891;
assign w36894 = ~w15703 & w15848;
assign w36895 = ~w14884 & ~w21690;
assign w36896 = ~w14884 & ~w21691;
assign w36897 = w21763 & w36895;
assign w36898 = w21763 & w36896;
assign w36899 = ~w21695 & w36897;
assign w36900 = ~w21695 & w36898;
assign w36901 = w21769 & ~w36897;
assign w36902 = w21769 & ~w36898;
assign w36903 = ~w21763 & ~w36895;
assign w36904 = ~w21763 & ~w36896;
assign w36905 = ~w21699 & w21777;
assign w36906 = w21699 & ~w21777;
assign w36907 = ~w21774 & w21780;
assign w36908 = w21206 & w21224;
assign w36909 = ~w20396 & ~w21218;
assign w36910 = w21475 & w32002;
assign w36911 = w32003 & w21907;
assign w36912 = (w21907 & w32003) | (w21907 & ~w21475) | (w32003 & ~w21475);
assign w36913 = w21475 & w21918;
assign w36914 = w32006 & ~w21916;
assign w36915 = (~w21916 & w32006) | (~w21916 & ~w21475) | (w32006 & ~w21475);
assign w36916 = w21930 & w21926;
assign w36917 = w21936 & ~w21931;
assign w36918 = w21936 & ~w32459;
assign w36919 = ~w21936 & w21931;
assign w36920 = ~w21936 & w32459;
assign w36921 = w21965 & w17633;
assign w36922 = w21965 & w32007;
assign w36923 = ~w21965 & ~w17633;
assign w36924 = ~w21965 & ~w32007;
assign w36925 = (~w21686 & w32011) | (~w21686 & w21680) | (w32011 & w21680);
assign w36926 = (~w21686 & w32011) | (~w21686 & w32456) | (w32011 & w32456);
assign w36927 = ~w15837 & ~w21682;
assign w36928 = ~w15837 & w36839;
assign w36929 = (w21982 & w32012) | (w21982 & w21680) | (w32012 & w21680);
assign w36930 = (w21982 & w32012) | (w21982 & w32456) | (w32012 & w32456);
assign w36931 = ~w15702 & ~w21682;
assign w36932 = ~w15702 & w36839;
assign w36933 = (w21987 & w32013) | (w21987 & w21680) | (w32013 & w21680);
assign w36934 = (w21987 & w32013) | (w21987 & w32456) | (w32013 & w32456);
assign w36935 = w21989 & w21986;
assign w36936 = ~w21989 & ~w21986;
assign w36937 = ~w21978 & w22001;
assign w36938 = ~w15838 & w22004;
assign w36939 = ~w22003 & ~w15848;
assign w36940 = ~w22003 & ~w36894;
assign w36941 = ~w15844 & ~w21690;
assign w36942 = ~w22012 & w22018;
assign w36943 = ~w22012 & w32014;
assign w36944 = w22024 & w22028;
assign w36945 = ~w36944 & ~w21783;
assign w36946 = w22029 & ~w36849;
assign w36947 = w22029 & ~w36850;
assign w36948 = ~w22029 & w36849;
assign w36949 = ~w22029 & w36850;
assign w36950 = ~w14320 & w36892;
assign w36951 = ~w14320 & w36893;
assign w36952 = ~w21777 & ~w36892;
assign w36953 = ~w21777 & ~w36893;
assign w36954 = w22037 & ~w36946;
assign w36955 = w22037 & ~w36947;
assign w36956 = w22041 & w21783;
assign w36957 = w22041 & ~w36945;
assign w36958 = ~w22045 & w22051;
assign w36959 = ~w22052 & ~w22051;
assign w36960 = ~w22052 & ~w36958;
assign w36961 = ~w21758 & w22056;
assign w36962 = ~w36961 & w22060;
assign w36963 = ~w21753 & ~w22060;
assign w36964 = ~w21753 & ~w36962;
assign w36965 = w21750 & w36963;
assign w36966 = w21750 & w36964;
assign w36967 = ~w21750 & ~w36963;
assign w36968 = ~w21750 & ~w36964;
assign w36969 = ~w10837 & w22066;
assign w36970 = a_2 & ~w22066;
assign w36971 = a_2 & ~w36969;
assign w36972 = w21905 & w22078;
assign w36973 = ~w7193 & w22085;
assign w36974 = ~a_11 & w22085;
assign w36975 = ~a_11 & w36973;
assign w36976 = ~w21893 & w6446;
assign w36977 = ~w5818 & ~w22163;
assign w36978 = ~w21797 & w5818;
assign w36979 = ~w5080 & ~w22194;
assign w36980 = ~w6061 & ~w22250;
assign w36981 = ~w22129 & a_20;
assign w36982 = ~w22129 & w32026;
assign w36983 = ~w22273 & a_17;
assign w36984 = w22273 & ~a_17;
assign w36985 = w22273 & ~w17695;
assign w36986 = ~w22334 & w32040;
assign w36987 = ~w22334 & ~w22335;
assign w36988 = ~w6063 & w22337;
assign w36989 = ~w6061 & ~w22341;
assign w36990 = w22339 & ~w22153;
assign w36991 = ~w21797 & w6061;
assign w36992 = ~w6998 & ~w22424;
assign w36993 = w22449 & ~a_14;
assign w36994 = ~w22449 & a_14;
assign w36995 = ~w22468 & w32059;
assign w36996 = ~w22468 & ~w22469;
assign w36997 = ~w6447 & w22471;
assign w36998 = ~w6998 & ~w22475;
assign w36999 = ~w6063 & w22336;
assign w37000 = ~w21797 & w6998;
assign w37001 = ~w8592 & ~w22452;
assign w37002 = ~w21893 & w6998;
assign w37003 = ~w6996 & ~w22557;
assign w37004 = ~w8592 & w22563;
assign w37005 = ~w22584 & a_14;
assign w37006 = w22584 & ~a_14;
assign w37007 = ~w8592 & w22588;
assign w37008 = w21818 & w5017;
assign w37009 = ~w22625 & a_20;
assign w37010 = w22625 & ~a_20;
assign w37011 = w22625 & ~w17294;
assign w37012 = ~w7193 & w22666;
assign w37013 = ~a_11 & ~w22666;
assign w37014 = ~a_11 & ~w37012;
assign w37015 = ~w21893 & w7192;
assign w37016 = ~w21893 & w7489;
assign w37017 = ~w7511 & ~w22690;
assign w37018 = ~w9089 & w22696;
assign w37019 = ~w7489 & ~w22744;
assign w37020 = w22762 & ~a_11;
assign w37021 = ~w22762 & a_11;
assign w37022 = ~w9089 & ~w22765;
assign w37023 = ~w22333 & a_14;
assign w37024 = ~w22333 & w32061;
assign w37025 = ~w9061 & w22772;
assign w37026 = ~w22787 & w32090;
assign w37027 = ~w22787 & ~w22788;
assign w37028 = ~w7193 & w22790;
assign w37029 = ~w7489 & ~w22794;
assign w37030 = ~w6447 & w22470;
assign w37031 = ~w21797 & w7489;
assign w37032 = w22879 & ~a_11;
assign w37033 = ~w22879 & a_11;
assign w37034 = ~w9089 & w22883;
assign w37035 = w21921 & w21910;
assign w37036 = ~w22903 & ~w22661;
assign w37037 = ~w22903 & w32079;
assign w37038 = ~w22904 & w7193;
assign w37039 = ~w22899 & ~w22900;
assign w37040 = w22907 & a_11;
assign w37041 = ~w22907 & ~a_11;
assign w37042 = ~w21958 & ~w21963;
assign w37043 = ~w32100 & ~w22924;
assign w37044 = w32100 & w22924;
assign w37045 = ~w9484 & w22939;
assign w37046 = ~w6447 & w22948;
assign w37047 = ~a_14 & w22948;
assign w37048 = ~a_14 & w37046;
assign w37049 = ~w21893 & w6061;
assign w37050 = ~w6304 & ~w22957;
assign w37051 = ~w8419 & w22963;
assign w37052 = ~w5818 & ~w22968;
assign w37053 = ~w4666 & ~w22979;
assign w37054 = ~w22980 & w22977;
assign w37055 = ~w22604 & ~a_23;
assign w37056 = ~w21797 & w5080;
assign w37057 = ~w7193 & w23034;
assign w37058 = ~a_11 & w23034;
assign w37059 = ~a_11 & w37057;
assign w37060 = ~w8278 & w23054;
assign w37061 = ~a_8 & w23054;
assign w37062 = ~a_8 & w37060;
assign w37063 = ~w21893 & w8277;
assign w37064 = ~w21893 & w8295;
assign w37065 = a_8 & ~w23081;
assign w37066 = a_8 & ~w32509;
assign w37067 = ~a_8 & w23081;
assign w37068 = ~a_8 & w32509;
assign w37069 = ~w8298 & ~w23114;
assign w37070 = ~w22467 & a_11;
assign w37071 = ~w22467 & w32092;
assign w37072 = ~w23139 & ~a_8;
assign w37073 = w23139 & a_8;
assign w37074 = ~w9484 & w23142;
assign w37075 = ~w21797 & w8277;
assign w37076 = ~w8298 & ~w23153;
assign w37077 = ~w23151 & w23148;
assign w37078 = ~w23177 & w32118;
assign w37079 = ~w23177 & ~w23174;
assign w37080 = ~w8278 & w23178;
assign w37081 = ~w8298 & ~w23182;
assign w37082 = ~w7193 & w22789;
assign w37083 = ~w21797 & w8298;
assign w37084 = w23162 & ~w23161;
assign w37085 = w23111 & ~w23089;
assign w37086 = ~w21893 & w8298;
assign w37087 = ~w8295 & ~w23223;
assign w37088 = ~w9484 & w23229;
assign w37089 = ~w23231 & ~w23221;
assign w37090 = w23238 & ~w23074;
assign w37091 = ~w23246 & a_8;
assign w37092 = w23246 & ~a_8;
assign w37093 = ~w9484 & w23250;
assign w37094 = ~w8278 & w23266;
assign w37095 = ~a_8 & w23266;
assign w37096 = ~a_8 & w37094;
assign w37097 = w23313 & a_8;
assign w37098 = ~w23313 & ~a_8;
assign w37099 = ~w9456 & ~w23315;
assign w37100 = ~w8278 & w23338;
assign w37101 = a_8 & ~w23338;
assign w37102 = a_8 & ~w37100;
assign w37103 = w22916 & ~w22918;
assign w37104 = ~w32100 & ~w23363;
assign w37105 = w23370 & ~a_8;
assign w37106 = ~w23370 & a_8;
assign w37107 = ~w9484 & w23374;
assign w37108 = w22010 & ~w22011;
assign w37109 = w22010 & ~w32128;
assign w37110 = ~w22019 & w10033;
assign w37111 = ~w22019 & w10061;
assign w37112 = ~w22904 & w6447;
assign w37113 = ~w23420 & ~w23422;
assign w37114 = w23424 & ~a_14;
assign w37115 = ~w23424 & a_14;
assign w37116 = w23430 & a_11;
assign w37117 = ~w23430 & ~a_11;
assign w37118 = ~w9061 & ~w23432;
assign w37119 = ~w32102 & a_26;
assign w37120 = ~w4638 & ~w23461;
assign w37121 = ~w21893 & w6059;
assign w37122 = ~w21978 & ~w21999;
assign w37123 = ~w21978 & w22000;
assign w37124 = ~w23552 & w9456;
assign w37125 = ~w23552 & w9484;
assign w37126 = ~w23558 & a_8;
assign w37127 = w23558 & ~a_8;
assign w37128 = ~w22010 & w22011;
assign w37129 = ~w22010 & w32128;
assign w37130 = ~w9790 & w23582;
assign w37131 = ~a_5 & w23582;
assign w37132 = ~a_5 & w37130;
assign w37133 = ~w10061 & w23617;
assign w37134 = ~w9790 & w23625;
assign w37135 = ~a_5 & w23625;
assign w37136 = ~a_5 & w37134;
assign w37137 = ~w23639 & a_5;
assign w37138 = w23639 & ~a_5;
assign w37139 = ~w10061 & w23643;
assign w37140 = ~w21893 & w9780;
assign w37141 = ~w9788 & ~w23654;
assign w37142 = ~w10061 & w23660;
assign w37143 = ~w21893 & w9788;
assign w37144 = a_5 & ~w23668;
assign w37145 = a_5 & ~w32527;
assign w37146 = ~a_5 & w23668;
assign w37147 = ~a_5 & w32527;
assign w37148 = ~w9790 & w23686;
assign w37149 = ~w9788 & ~w23699;
assign w37150 = a_5 & ~w23702;
assign w37151 = a_5 & ~w32528;
assign w37152 = ~a_5 & w23702;
assign w37153 = ~a_5 & w32528;
assign w37154 = ~w22786 & a_8;
assign w37155 = ~w22786 & w32120;
assign w37156 = ~w23721 & ~a_5;
assign w37157 = w23721 & a_5;
assign w37158 = ~w10061 & w23724;
assign w37159 = ~w21797 & w9788;
assign w37160 = ~w9788 & ~w23741;
assign w37161 = ~w9790 & w23742;
assign w37162 = ~w9780 & ~w23747;
assign w37163 = w23745 & ~w23176;
assign w37164 = ~w8278 & w23175;
assign w37165 = ~w21797 & w9780;
assign w37166 = ~w21797 & w9786;
assign w37167 = ~w9780 & ~w23779;
assign w37168 = w10033 & ~w23777;
assign w37169 = ~w10033 & w23777;
assign w37170 = w23711 & ~w23710;
assign w37171 = w23797 & ~w23694;
assign w37172 = ~w23662 & ~w23676;
assign w37173 = ~w21893 & w9786;
assign w37174 = ~w9790 & w23809;
assign w37175 = ~a_5 & ~w23809;
assign w37176 = ~a_5 & ~w37174;
assign w37177 = ~w23214 & ~w23127;
assign w37178 = ~w23645 & ~w23819;
assign w37179 = ~w9790 & w23831;
assign w37180 = ~a_5 & ~w23831;
assign w37181 = ~a_5 & ~w37179;
assign w37182 = ~w22904 & w10033;
assign w37183 = ~w23845 & ~w23847;
assign w37184 = ~w22904 & w10061;
assign w37185 = ~w9790 & w23873;
assign w37186 = ~a_5 & w23873;
assign w37187 = ~a_5 & w37185;
assign w37188 = ~w9790 & w23886;
assign w37189 = ~a_5 & w23886;
assign w37190 = ~a_5 & w37188;
assign w37191 = ~w23242 & ~w23258;
assign w37192 = w23629 & ~w23899;
assign w37193 = w23908 & a_5;
assign w37194 = ~w23908 & ~a_5;
assign w37195 = ~w10033 & ~w23910;
assign w37196 = w23361 & w23385;
assign w37197 = ~w21996 & w21995;
assign w37198 = w21996 & ~w21995;
assign w37199 = ~w9790 & w23932;
assign w37200 = ~a_5 & ~w23932;
assign w37201 = ~a_5 & ~w37199;
assign w37202 = ~w23552 & w9790;
assign w37203 = w23945 & ~a_5;
assign w37204 = ~w23945 & a_5;
assign w37205 = ~w23331 & w23948;
assign w37206 = w23331 & ~w23948;
assign w37207 = w23570 & w23971;
assign w37208 = w23978 & ~w23980;
assign w37209 = ~w23985 & a_8;
assign w37210 = w23985 & ~a_8;
assign w37211 = ~w9484 & w23989;
assign w37212 = ~w23999 & a_17;
assign w37213 = w23999 & ~a_17;
assign w37214 = ~w8419 & w24003;
assign w37215 = w23459 & a_26;
assign w37216 = ~w24039 & a_23;
assign w37217 = w24039 & ~a_23;
assign w37218 = w24039 & ~w24044;
assign w37219 = ~w6447 & w24072;
assign w37220 = ~a_14 & w24072;
assign w37221 = ~a_14 & w37219;
assign w37222 = ~w24083 & a_11;
assign w37223 = w24083 & ~a_11;
assign w37224 = ~w9089 & w24087;
assign w37225 = ~w22015 & ~w22018;
assign w37226 = ~w22015 & ~w36942;
assign w37227 = ~w9790 & w24124;
assign w37228 = a_5 & ~w24124;
assign w37229 = a_5 & ~w37227;
assign w37230 = ~w23981 & w24089;
assign w37231 = ~w9089 & w24160;
assign w37232 = ~w6063 & w24168;
assign w37233 = a_17 & ~w24168;
assign w37234 = a_17 & ~w37232;
assign w37235 = ~w21893 & w5818;
assign w37236 = ~w5816 & ~w24177;
assign w37237 = ~w8339 & w24183;
assign w37238 = ~w5080 & ~w24188;
assign w37239 = ~w4446 & ~w24208;
assign w37240 = ~w24209 & w24201;
assign w37241 = w24209 & ~w24201;
assign w37242 = ~w21797 & w4638;
assign w37243 = ~w6447 & w24251;
assign w37244 = ~a_14 & ~w24251;
assign w37245 = ~a_14 & ~w37243;
assign w37246 = ~w24276 & a_8;
assign w37247 = w24276 & ~a_8;
assign w37248 = ~w9484 & w24280;
assign w37249 = w22024 & ~w24292;
assign w37250 = ~w22024 & w24292;
assign w37251 = ~w24299 & a_5;
assign w37252 = w24299 & ~a_5;
assign w37253 = ~w10061 & w24303;
assign w37254 = ~w23552 & w9061;
assign w37255 = ~w23552 & w9089;
assign w37256 = ~w24332 & a_11;
assign w37257 = w24332 & ~a_11;
assign w37258 = w3956 & a_29;
assign w37259 = ~w21893 & w5308;
assign w37260 = ~w22904 & w8391;
assign w37261 = ~w24433 & ~w24435;
assign w37262 = w24455 & a_14;
assign w37263 = ~w24455 & ~a_14;
assign w37264 = ~w8564 & ~w24457;
assign w37265 = ~w22019 & w9456;
assign w37266 = ~w22019 & w9484;
assign w37267 = w22024 & w22027;
assign w37268 = w21775 & ~w22026;
assign w37269 = w24500 & ~w24292;
assign w37270 = w24500 & ~w37250;
assign w37271 = ~w24501 & w10033;
assign w37272 = ~w24501 & w10061;
assign w37273 = ~w21761 & w9788;
assign w37274 = ~w24507 & a_5;
assign w37275 = w24507 & ~a_5;
assign w37276 = ~w21761 & w9780;
assign w37277 = w21775 & w21780;
assign w37278 = ~w21775 & ~w21780;
assign w37279 = ~w9790 & w24531;
assign w37280 = ~a_5 & w24531;
assign w37281 = ~a_5 & w37279;
assign w37282 = ~w24558 & a_11;
assign w37283 = w24558 & ~a_11;
assign w37284 = ~w9089 & w24562;
assign w37285 = ~w24244 & w24451;
assign w37286 = ~w24570 & a_14;
assign w37287 = w24570 & ~a_14;
assign w37288 = ~w8592 & w24574;
assign w37289 = ~w21225 & w4666;
assign w37290 = ~w4403 & w24624;
assign w37291 = w24643 & w21914;
assign w37292 = w24643 & ~w32069;
assign w37293 = ~w21905 & w24646;
assign w37294 = ~w24648 & ~a_20;
assign w37295 = w24648 & a_20;
assign w37296 = w24657 & ~w21914;
assign w37297 = w24657 & w32069;
assign w37298 = w24659 & w21914;
assign w37299 = w24659 & ~w32069;
assign w37300 = ~a_17 & w24678;
assign w37301 = ~a_17 & w32170;
assign w37302 = a_17 & ~w24678;
assign w37303 = a_17 & ~w32170;
assign w37304 = ~w24708 & a_8;
assign w37305 = w24708 & ~a_8;
assign w37306 = ~w9484 & w24712;
assign w37307 = ~w24746 & a_8;
assign w37308 = w24746 & ~a_8;
assign w37309 = ~w9484 & w24750;
assign w37310 = w24753 & ~w21783;
assign w37311 = w24753 & w36945;
assign w37312 = ~w24753 & w21783;
assign w37313 = ~w24753 & ~w36945;
assign w37314 = ~w21761 & w9786;
assign w37315 = w24760 & ~a_5;
assign w37316 = ~w24760 & a_5;
assign w37317 = ~w10061 & w24764;
assign w37318 = ~w21893 & w5080;
assign w37319 = ~w5286 & ~w24779;
assign w37320 = ~w4638 & ~w24790;
assign w37321 = a_26 & w4;
assign w37322 = ~w21797 & w4068;
assign w37323 = ~w5309 & w24877;
assign w37324 = ~a_20 & ~w24877;
assign w37325 = ~a_20 & ~w37323;
assign w37326 = w24891 & ~a_11;
assign w37327 = ~w24891 & a_11;
assign w37328 = ~w9089 & w24895;
assign w37329 = ~w21974 & w8592;
assign w37330 = w32100 & w24900;
assign w37331 = ~w6063 & w24917;
assign w37332 = a_17 & ~w24917;
assign w37333 = a_17 & ~w37331;
assign w37334 = w22045 & ~w22040;
assign w37335 = ~w9790 & w24964;
assign w37336 = a_5 & ~w24964;
assign w37337 = a_5 & ~w37335;
assign w37338 = w24741 & w24933;
assign w37339 = ~w21761 & w8295;
assign w37340 = ~w24501 & w8278;
assign w37341 = w24983 & ~a_8;
assign w37342 = ~w24983 & a_8;
assign w37343 = ~w21893 & w5016;
assign w37344 = ~w21797 & w3957;
assign w37345 = ~w4068 & ~w25029;
assign w37346 = ~w24839 & ~w25049;
assign w37347 = w24839 & w25049;
assign w37348 = ~w1327 & ~w25054;
assign w37349 = ~w25098 & a_20;
assign w37350 = w25098 & ~a_20;
assign w37351 = w25105 & ~a_17;
assign w37352 = ~w25105 & a_17;
assign w37353 = ~w22925 & w25109;
assign w37354 = ~w22019 & w7193;
assign w37355 = w25129 & a_11;
assign w37356 = ~w25129 & ~a_11;
assign w37357 = ~w23552 & w6447;
assign w37358 = ~w25138 & a_14;
assign w37359 = w25138 & ~a_14;
assign w37360 = ~w24975 & ~w24703;
assign w37361 = ~w24975 & w24737;
assign w37362 = ~w21761 & w8298;
assign w37363 = ~w8278 & w25195;
assign w37364 = a_8 & ~w25195;
assign w37365 = a_8 & ~w37363;
assign w37366 = ~w22045 & w22048;
assign w37367 = w22045 & ~w22048;
assign w37368 = ~w9790 & w25207;
assign w37369 = ~a_5 & w25207;
assign w37370 = ~a_5 & w37368;
assign w37371 = w25212 & w25183;
assign w37372 = w25212 & ~w24996;
assign w37373 = w25214 & ~w25183;
assign w37374 = w25214 & w24996;
assign w37375 = ~w5309 & w25235;
assign w37376 = ~a_20 & w25235;
assign w37377 = ~a_20 & w37375;
assign w37378 = w25242 & a_23;
assign w37379 = ~w25242 & ~a_23;
assign w37380 = ~w7961 & ~w25244;
assign w37381 = ~w25255 & a_29;
assign w37382 = w25255 & ~a_29;
assign w37383 = w25255 & ~w25260;
assign w37384 = ~w6063 & w25340;
assign w37385 = ~a_17 & w25340;
assign w37386 = ~a_17 & w37384;
assign w37387 = w25347 & a_14;
assign w37388 = ~w25347 & ~a_14;
assign w37389 = ~w8564 & ~w25349;
assign w37390 = ~w25393 & a_11;
assign w37391 = w25393 & ~a_11;
assign w37392 = ~w9089 & w25397;
assign w37393 = ~w25214 & w25183;
assign w37394 = ~w25214 & ~w24996;
assign w37395 = ~w25212 & ~w25183;
assign w37396 = ~w25212 & w24996;
assign w37397 = w25425 & w25179;
assign w37398 = w25425 & ~w25170;
assign w37399 = w25122 & ~w25470;
assign w37400 = ~w5017 & w25481;
assign w37401 = ~a_23 & ~w25481;
assign w37402 = ~a_23 & ~w37400;
assign w37403 = ~w4446 & ~w25489;
assign w37404 = ~w22245 & w25492;
assign w37405 = ~w21797 & w1327;
assign w37406 = ~w21893 & w4638;
assign w37407 = ~w4666 & ~w25537;
assign w37408 = ~w5309 & w25565;
assign w37409 = ~a_20 & w25565;
assign w37410 = ~a_20 & w37408;
assign w37411 = ~w8419 & w25578;
assign w37412 = ~w6447 & w25608;
assign w37413 = ~a_14 & w25608;
assign w37414 = ~a_14 & w37412;
assign w37415 = ~w25616 & a_11;
assign w37416 = w25616 & ~a_11;
assign w37417 = ~w9089 & w25620;
assign w37418 = ~w21761 & w8277;
assign w37419 = ~w8278 & w25652;
assign w37420 = ~a_8 & w25652;
assign w37421 = ~a_8 & w37419;
assign w37422 = ~w25656 & w25388;
assign w37423 = ~w25656 & w25189;
assign w37424 = w25656 & ~w25388;
assign w37425 = w25656 & ~w25189;
assign w37426 = w25665 & ~w25448;
assign w37427 = w25665 & ~w25178;
assign w37428 = ~w21754 & w9788;
assign w37429 = w25673 & ~w22048;
assign w37430 = w25673 & ~w37366;
assign w37431 = ~w9790 & w25677;
assign w37432 = a_5 & ~w25677;
assign w37433 = a_5 & ~w37431;
assign w37434 = ~w36961 & ~w22054;
assign w37435 = ~w22059 & w22054;
assign w37436 = ~w22059 & ~w37434;
assign w37437 = ~w10837 & w25701;
assign w37438 = a_2 & ~w25701;
assign w37439 = a_2 & ~w37437;
assign w37440 = ~w10837 & w25715;
assign w37441 = a_2 & ~w25715;
assign w37442 = a_2 & ~w37440;
assign w37443 = ~w10837 & w25727;
assign w37444 = a_2 & ~w25727;
assign w37445 = a_2 & ~w37443;
assign w37446 = ~w10837 & w25736;
assign w37447 = a_2 & ~w25736;
assign w37448 = a_2 & ~w37446;
assign w37449 = ~w23954 & ~w23620;
assign w37450 = ~w23954 & w23919;
assign w37451 = ~w10837 & w25753;
assign w37452 = a_2 & ~w25753;
assign w37453 = a_2 & ~w37451;
assign w37454 = ~w22904 & w10837;
assign w37455 = ~w25765 & a_2;
assign w37456 = ~w10837 & w25774;
assign w37457 = a_2 & ~w25774;
assign w37458 = a_2 & ~w37456;
assign w37459 = ~w10837 & w25791;
assign w37460 = a_2 & ~w25791;
assign w37461 = a_2 & ~w37459;
assign w37462 = ~w21893 & w10909;
assign w37463 = ~w21893 & w10835;
assign w37464 = a_2 & ~w25812;
assign w37465 = a_2 & ~w32577;
assign w37466 = ~w21893 & w3;
assign w37467 = ~w10837 & w25840;
assign w37468 = ~w10837 & w25855;
assign w37469 = a_2 & w25855;
assign w37470 = a_2 & w37468;
assign w37471 = w25858 & ~w25852;
assign w37472 = ~w3 & ~w25870;
assign w37473 = ~w25872 & a_2;
assign w37474 = w25874 & ~w25869;
assign w37475 = ~w25874 & w25869;
assign w37476 = ~w21797 & w10839;
assign w37477 = ~w10837 & w25885;
assign w37478 = a_2 & ~w25885;
assign w37479 = a_2 & ~w37477;
assign w37480 = w25888 & ~w25880;
assign w37481 = ~w25888 & w25880;
assign w37482 = ~w21797 & w3;
assign w37483 = a_2 & ~w25895;
assign w37484 = a_2 & ~w32582;
assign w37485 = w10839 & w25901;
assign w37486 = ~w25902 & ~w23737;
assign w37487 = ~w21797 & w10835;
assign w37488 = ~w3 & ~w25908;
assign w37489 = ~a_2 & ~w25909;
assign w37490 = ~a_2 & ~w32583;
assign w37491 = w25907 & ~w25906;
assign w37492 = w25890 & ~w25889;
assign w37493 = ~w25828 & ~w25851;
assign w37494 = w25809 & ~w25798;
assign w37495 = ~w10837 & w25935;
assign w37496 = a_2 & w25935;
assign w37497 = a_2 & w37495;
assign w37498 = w25938 & ~w25932;
assign w37499 = ~w25797 & w25939;
assign w37500 = ~w37499 & w25945;
assign w37501 = ~w25786 & ~w25946;
assign w37502 = ~w10837 & w25956;
assign w37503 = a_2 & ~w25956;
assign w37504 = a_2 & ~w37502;
assign w37505 = ~w10837 & w25973;
assign w37506 = a_2 & ~w25973;
assign w37507 = a_2 & ~w37505;
assign w37508 = ~w10837 & w25987;
assign w37509 = a_2 & ~w25987;
assign w37510 = a_2 & ~w37508;
assign w37511 = ~w10837 & w25999;
assign w37512 = a_2 & ~w25999;
assign w37513 = a_2 & ~w37511;
assign w37514 = ~w26004 & ~w25996;
assign w37515 = ~w23552 & w10837;
assign w37516 = ~w26016 & a_2;
assign w37517 = ~w22019 & w10837;
assign w37518 = ~w26036 & a_2;
assign w37519 = ~w10837 & w26049;
assign w37520 = a_2 & ~w26049;
assign w37521 = a_2 & ~w37519;
assign w37522 = w23954 & w23620;
assign w37523 = w23954 & ~w23919;
assign w37524 = ~w21761 & w10835;
assign w37525 = ~w10837 & w26081;
assign w37526 = a_2 & ~w26081;
assign w37527 = a_2 & ~w37525;
assign w37528 = ~w23592 & ~w26087;
assign w37529 = w23592 & w26087;
assign w37530 = ~w21761 & w3;
assign w37531 = ~w24501 & w10837;
assign w37532 = ~w26094 & a_2;
assign w37533 = w26086 & ~w26100;
assign w37534 = w26086 & w26104;
assign w37535 = ~w10837 & w26117;
assign w37536 = a_2 & ~w26117;
assign w37537 = a_2 & ~w37535;
assign w37538 = ~w10837 & w26134;
assign w37539 = a_2 & ~w26134;
assign w37540 = a_2 & ~w37538;
assign w37541 = ~w24948 & w24951;
assign w37542 = ~w24948 & w24730;
assign w37543 = ~w21754 & w3;
assign w37544 = ~w10837 & w26148;
assign w37545 = a_2 & ~w26148;
assign w37546 = a_2 & ~w37544;
assign w37547 = ~w21754 & w10835;
assign w37548 = w21758 & ~w22056;
assign w37549 = ~w10837 & w26167;
assign w37550 = a_2 & ~w26167;
assign w37551 = a_2 & ~w37549;
assign w37552 = w26172 & ~w26157;
assign w37553 = ~w26176 & ~w25707;
assign w37554 = ~w21754 & w9780;
assign w37555 = ~w9790 & w26212;
assign w37556 = ~w8278 & w26223;
assign w37557 = a_8 & ~w26223;
assign w37558 = a_8 & ~w37556;
assign w37559 = w26232 & ~w26231;
assign w37560 = ~w21761 & w7511;
assign w37561 = ~w24501 & w7193;
assign w37562 = w26240 & ~a_11;
assign w37563 = ~w7268 & ~w7316;
assign w37564 = ~w4403 & ~w7600;
assign w37565 = ~w5017 & w16671;
assign w37566 = ~w5017 & w16675;
assign w37567 = ~w16677 & ~w16678;
assign w37568 = w16384 & w16011;
assign w37569 = ~w17284 & ~w17437;
assign w37570 = ~w18154 & w18160;
assign w37571 = w18201 & ~w18205;
assign w37572 = w18752 & ~w18774;
assign w37573 = w18775 & w18802;
assign w37574 = ~w18712 & ~w18739;
assign w37575 = w18712 & ~w18933;
assign w37576 = ~w18686 & ~w18691;
assign w37577 = ~w19371 & w18938;
assign w37578 = w19382 & ~w18776;
assign w37579 = ~w19900 & ~w19917;
assign w37580 = ~w27102 & ~w27103;
assign w37581 = ~w27102 & w26813;
assign w37582 = w27102 & w27103;
assign w37583 = w27102 & ~w26813;
assign one = 1;
assign result_0 = w26506;// level 167
assign result_1 = w26795;// level 168
assign result_2 = w27085;// level 169
assign result_3 = w27335;// level 170
assign result_4 = w27592;// level 172
assign result_5 = w27831;// level 173
assign result_6 = w28080;// level 174
assign result_7 = w28316;// level 175
assign result_8 = w28533;// level 176
assign result_9 = w28725;// level 177
assign result_10 = w28921;// level 178
assign result_11 = w29123;// level 179
assign result_12 = w29313;// level 179
assign result_13 = w29493;// level 179
assign result_14 = w29666;// level 180
assign result_15 = w29823;// level 179
assign result_16 = w29992;// level 180
assign result_17 = w30142;// level 180
assign result_18 = w30282;// level 180
assign result_19 = w30420;// level 180
assign result_20 = w30544;// level 180
assign result_21 = w30673;// level 180
assign result_22 = w30787;// level 180
assign result_23 = w30898;// level 180
assign result_24 = ~w31007;// level 180
assign result_25 = ~w31115;// level 180
assign result_26 = w31208;// level 180
assign result_27 = ~w31289;// level 180
assign result_28 = ~w31372;// level 180
assign result_29 = w31445;// level 180
assign result_30 = w31512;// level 181
assign result_31 = ~w31559;// level 181
endmodule

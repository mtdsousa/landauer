//Written by the Majority Logic Package Thu Jun 18 12:07:41 2015
module top (
            in0_0, in0_1, in0_2, in0_3, in0_4, in0_5, in0_6, in0_7, in0_8, in0_9, in0_10, in0_11, in0_12, in0_13, in0_14, in0_15, in0_16, in0_17, in0_18, in0_19, in0_20, in0_21, in0_22, in0_23, in0_24, in0_25, in0_26, in0_27, in0_28, in0_29, in0_30, in0_31, in0_32, in0_33, in0_34, in0_35, in0_36, in0_37, in0_38, in0_39, in0_40, in0_41, in0_42, in0_43, in0_44, in0_45, in0_46, in0_47, in0_48, in0_49, in0_50, in0_51, in0_52, in0_53, in0_54, in0_55, in0_56, in0_57, in0_58, in0_59, in0_60, in0_61, in0_62, in0_63, in0_64, in0_65, in0_66, in0_67, in0_68, in0_69, in0_70, in0_71, in0_72, in0_73, in0_74, in0_75, in0_76, in0_77, in0_78, in0_79, in0_80, in0_81, in0_82, in0_83, in0_84, in0_85, in0_86, in0_87, in0_88, in0_89, in0_90, in0_91, in0_92, in0_93, in0_94, in0_95, in0_96, in0_97, in0_98, in0_99, in0_100, in0_101, in0_102, in0_103, in0_104, in0_105, in0_106, in0_107, in0_108, in0_109, in0_110, in0_111, in0_112, in0_113, in0_114, in0_115, in0_116, in0_117, in0_118, in0_119, in0_120, in0_121, in0_122, in0_123, in0_124, in0_125, in0_126, in0_127, in1_0, in1_1, in1_2, in1_3, in1_4, in1_5, in1_6, in1_7, in1_8, in1_9, in1_10, in1_11, in1_12, in1_13, in1_14, in1_15, in1_16, in1_17, in1_18, in1_19, in1_20, in1_21, in1_22, in1_23, in1_24, in1_25, in1_26, in1_27, in1_28, in1_29, in1_30, in1_31, in1_32, in1_33, in1_34, in1_35, in1_36, in1_37, in1_38, in1_39, in1_40, in1_41, in1_42, in1_43, in1_44, in1_45, in1_46, in1_47, in1_48, in1_49, in1_50, in1_51, in1_52, in1_53, in1_54, in1_55, in1_56, in1_57, in1_58, in1_59, in1_60, in1_61, in1_62, in1_63, in1_64, in1_65, in1_66, in1_67, in1_68, in1_69, in1_70, in1_71, in1_72, in1_73, in1_74, in1_75, in1_76, in1_77, in1_78, in1_79, in1_80, in1_81, in1_82, in1_83, in1_84, in1_85, in1_86, in1_87, in1_88, in1_89, in1_90, in1_91, in1_92, in1_93, in1_94, in1_95, in1_96, in1_97, in1_98, in1_99, in1_100, in1_101, in1_102, in1_103, in1_104, in1_105, in1_106, in1_107, in1_108, in1_109, in1_110, in1_111, in1_112, in1_113, in1_114, in1_115, in1_116, in1_117, in1_118, in1_119, in1_120, in1_121, in1_122, in1_123, in1_124, in1_125, in1_126, in1_127, in2_0, in2_1, in2_2, in2_3, in2_4, in2_5, in2_6, in2_7, in2_8, in2_9, in2_10, in2_11, in2_12, in2_13, in2_14, in2_15, in2_16, in2_17, in2_18, in2_19, in2_20, in2_21, in2_22, in2_23, in2_24, in2_25, in2_26, in2_27, in2_28, in2_29, in2_30, in2_31, in2_32, in2_33, in2_34, in2_35, in2_36, in2_37, in2_38, in2_39, in2_40, in2_41, in2_42, in2_43, in2_44, in2_45, in2_46, in2_47, in2_48, in2_49, in2_50, in2_51, in2_52, in2_53, in2_54, in2_55, in2_56, in2_57, in2_58, in2_59, in2_60, in2_61, in2_62, in2_63, in2_64, in2_65, in2_66, in2_67, in2_68, in2_69, in2_70, in2_71, in2_72, in2_73, in2_74, in2_75, in2_76, in2_77, in2_78, in2_79, in2_80, in2_81, in2_82, in2_83, in2_84, in2_85, in2_86, in2_87, in2_88, in2_89, in2_90, in2_91, in2_92, in2_93, in2_94, in2_95, in2_96, in2_97, in2_98, in2_99, in2_100, in2_101, in2_102, in2_103, in2_104, in2_105, in2_106, in2_107, in2_108, in2_109, in2_110, in2_111, in2_112, in2_113, in2_114, in2_115, in2_116, in2_117, in2_118, in2_119, in2_120, in2_121, in2_122, in2_123, in2_124, in2_125, in2_126, in2_127, in3_0, in3_1, in3_2, in3_3, in3_4, in3_5, in3_6, in3_7, in3_8, in3_9, in3_10, in3_11, in3_12, in3_13, in3_14, in3_15, in3_16, in3_17, in3_18, in3_19, in3_20, in3_21, in3_22, in3_23, in3_24, in3_25, in3_26, in3_27, in3_28, in3_29, in3_30, in3_31, in3_32, in3_33, in3_34, in3_35, in3_36, in3_37, in3_38, in3_39, in3_40, in3_41, in3_42, in3_43, in3_44, in3_45, in3_46, in3_47, in3_48, in3_49, in3_50, in3_51, in3_52, in3_53, in3_54, in3_55, in3_56, in3_57, in3_58, in3_59, in3_60, in3_61, in3_62, in3_63, in3_64, in3_65, in3_66, in3_67, in3_68, in3_69, in3_70, in3_71, in3_72, in3_73, in3_74, in3_75, in3_76, in3_77, in3_78, in3_79, in3_80, in3_81, in3_82, in3_83, in3_84, in3_85, in3_86, in3_87, in3_88, in3_89, in3_90, in3_91, in3_92, in3_93, in3_94, in3_95, in3_96, in3_97, in3_98, in3_99, in3_100, in3_101, in3_102, in3_103, in3_104, in3_105, in3_106, in3_107, in3_108, in3_109, in3_110, in3_111, in3_112, in3_113, in3_114, in3_115, in3_116, in3_117, in3_118, in3_119, in3_120, in3_121, in3_122, in3_123, in3_124, in3_125, in3_126, in3_127, 
            result_0, result_1, result_2, result_3, result_4, result_5, result_6, result_7, result_8, result_9, result_10, result_11, result_12, result_13, result_14, result_15, result_16, result_17, result_18, result_19, result_20, result_21, result_22, result_23, result_24, result_25, result_26, result_27, result_28, result_29, result_30, result_31, result_32, result_33, result_34, result_35, result_36, result_37, result_38, result_39, result_40, result_41, result_42, result_43, result_44, result_45, result_46, result_47, result_48, result_49, result_50, result_51, result_52, result_53, result_54, result_55, result_56, result_57, result_58, result_59, result_60, result_61, result_62, result_63, result_64, result_65, result_66, result_67, result_68, result_69, result_70, result_71, result_72, result_73, result_74, result_75, result_76, result_77, result_78, result_79, result_80, result_81, result_82, result_83, result_84, result_85, result_86, result_87, result_88, result_89, result_90, result_91, result_92, result_93, result_94, result_95, result_96, result_97, result_98, result_99, result_100, result_101, result_102, result_103, result_104, result_105, result_106, result_107, result_108, result_109, result_110, result_111, result_112, result_113, result_114, result_115, result_116, result_117, result_118, result_119, result_120, result_121, result_122, result_123, result_124, result_125, result_126, result_127, address_0, address_1);
input in0_0, in0_1, in0_2, in0_3, in0_4, in0_5, in0_6, in0_7, in0_8, in0_9, in0_10, in0_11, in0_12, in0_13, in0_14, in0_15, in0_16, in0_17, in0_18, in0_19, in0_20, in0_21, in0_22, in0_23, in0_24, in0_25, in0_26, in0_27, in0_28, in0_29, in0_30, in0_31, in0_32, in0_33, in0_34, in0_35, in0_36, in0_37, in0_38, in0_39, in0_40, in0_41, in0_42, in0_43, in0_44, in0_45, in0_46, in0_47, in0_48, in0_49, in0_50, in0_51, in0_52, in0_53, in0_54, in0_55, in0_56, in0_57, in0_58, in0_59, in0_60, in0_61, in0_62, in0_63, in0_64, in0_65, in0_66, in0_67, in0_68, in0_69, in0_70, in0_71, in0_72, in0_73, in0_74, in0_75, in0_76, in0_77, in0_78, in0_79, in0_80, in0_81, in0_82, in0_83, in0_84, in0_85, in0_86, in0_87, in0_88, in0_89, in0_90, in0_91, in0_92, in0_93, in0_94, in0_95, in0_96, in0_97, in0_98, in0_99, in0_100, in0_101, in0_102, in0_103, in0_104, in0_105, in0_106, in0_107, in0_108, in0_109, in0_110, in0_111, in0_112, in0_113, in0_114, in0_115, in0_116, in0_117, in0_118, in0_119, in0_120, in0_121, in0_122, in0_123, in0_124, in0_125, in0_126, in0_127, in1_0, in1_1, in1_2, in1_3, in1_4, in1_5, in1_6, in1_7, in1_8, in1_9, in1_10, in1_11, in1_12, in1_13, in1_14, in1_15, in1_16, in1_17, in1_18, in1_19, in1_20, in1_21, in1_22, in1_23, in1_24, in1_25, in1_26, in1_27, in1_28, in1_29, in1_30, in1_31, in1_32, in1_33, in1_34, in1_35, in1_36, in1_37, in1_38, in1_39, in1_40, in1_41, in1_42, in1_43, in1_44, in1_45, in1_46, in1_47, in1_48, in1_49, in1_50, in1_51, in1_52, in1_53, in1_54, in1_55, in1_56, in1_57, in1_58, in1_59, in1_60, in1_61, in1_62, in1_63, in1_64, in1_65, in1_66, in1_67, in1_68, in1_69, in1_70, in1_71, in1_72, in1_73, in1_74, in1_75, in1_76, in1_77, in1_78, in1_79, in1_80, in1_81, in1_82, in1_83, in1_84, in1_85, in1_86, in1_87, in1_88, in1_89, in1_90, in1_91, in1_92, in1_93, in1_94, in1_95, in1_96, in1_97, in1_98, in1_99, in1_100, in1_101, in1_102, in1_103, in1_104, in1_105, in1_106, in1_107, in1_108, in1_109, in1_110, in1_111, in1_112, in1_113, in1_114, in1_115, in1_116, in1_117, in1_118, in1_119, in1_120, in1_121, in1_122, in1_123, in1_124, in1_125, in1_126, in1_127, in2_0, in2_1, in2_2, in2_3, in2_4, in2_5, in2_6, in2_7, in2_8, in2_9, in2_10, in2_11, in2_12, in2_13, in2_14, in2_15, in2_16, in2_17, in2_18, in2_19, in2_20, in2_21, in2_22, in2_23, in2_24, in2_25, in2_26, in2_27, in2_28, in2_29, in2_30, in2_31, in2_32, in2_33, in2_34, in2_35, in2_36, in2_37, in2_38, in2_39, in2_40, in2_41, in2_42, in2_43, in2_44, in2_45, in2_46, in2_47, in2_48, in2_49, in2_50, in2_51, in2_52, in2_53, in2_54, in2_55, in2_56, in2_57, in2_58, in2_59, in2_60, in2_61, in2_62, in2_63, in2_64, in2_65, in2_66, in2_67, in2_68, in2_69, in2_70, in2_71, in2_72, in2_73, in2_74, in2_75, in2_76, in2_77, in2_78, in2_79, in2_80, in2_81, in2_82, in2_83, in2_84, in2_85, in2_86, in2_87, in2_88, in2_89, in2_90, in2_91, in2_92, in2_93, in2_94, in2_95, in2_96, in2_97, in2_98, in2_99, in2_100, in2_101, in2_102, in2_103, in2_104, in2_105, in2_106, in2_107, in2_108, in2_109, in2_110, in2_111, in2_112, in2_113, in2_114, in2_115, in2_116, in2_117, in2_118, in2_119, in2_120, in2_121, in2_122, in2_123, in2_124, in2_125, in2_126, in2_127, in3_0, in3_1, in3_2, in3_3, in3_4, in3_5, in3_6, in3_7, in3_8, in3_9, in3_10, in3_11, in3_12, in3_13, in3_14, in3_15, in3_16, in3_17, in3_18, in3_19, in3_20, in3_21, in3_22, in3_23, in3_24, in3_25, in3_26, in3_27, in3_28, in3_29, in3_30, in3_31, in3_32, in3_33, in3_34, in3_35, in3_36, in3_37, in3_38, in3_39, in3_40, in3_41, in3_42, in3_43, in3_44, in3_45, in3_46, in3_47, in3_48, in3_49, in3_50, in3_51, in3_52, in3_53, in3_54, in3_55, in3_56, in3_57, in3_58, in3_59, in3_60, in3_61, in3_62, in3_63, in3_64, in3_65, in3_66, in3_67, in3_68, in3_69, in3_70, in3_71, in3_72, in3_73, in3_74, in3_75, in3_76, in3_77, in3_78, in3_79, in3_80, in3_81, in3_82, in3_83, in3_84, in3_85, in3_86, in3_87, in3_88, in3_89, in3_90, in3_91, in3_92, in3_93, in3_94, in3_95, in3_96, in3_97, in3_98, in3_99, in3_100, in3_101, in3_102, in3_103, in3_104, in3_105, in3_106, in3_107, in3_108, in3_109, in3_110, in3_111, in3_112, in3_113, in3_114, in3_115, in3_116, in3_117, in3_118, in3_119, in3_120, in3_121, in3_122, in3_123, in3_124, in3_125, in3_126, in3_127;
output result_0, result_1, result_2, result_3, result_4, result_5, result_6, result_7, result_8, result_9, result_10, result_11, result_12, result_13, result_14, result_15, result_16, result_17, result_18, result_19, result_20, result_21, result_22, result_23, result_24, result_25, result_26, result_27, result_28, result_29, result_30, result_31, result_32, result_33, result_34, result_35, result_36, result_37, result_38, result_39, result_40, result_41, result_42, result_43, result_44, result_45, result_46, result_47, result_48, result_49, result_50, result_51, result_52, result_53, result_54, result_55, result_56, result_57, result_58, result_59, result_60, result_61, result_62, result_63, result_64, result_65, result_66, result_67, result_68, result_69, result_70, result_71, result_72, result_73, result_74, result_75, result_76, result_77, result_78, result_79, result_80, result_81, result_82, result_83, result_84, result_85, result_86, result_87, result_88, result_89, result_90, result_91, result_92, result_93, result_94, result_95, result_96, result_97, result_98, result_99, result_100, result_101, result_102, result_103, result_104, result_105, result_106, result_107, result_108, result_109, result_110, result_111, result_112, result_113, result_114, result_115, result_116, result_117, result_118, result_119, result_120, result_121, result_122, result_123, result_124, result_125, result_126, result_127, address_0, address_1;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201;
assign w0 = in0_1 & ~in1_1;
assign w1 = in0_0 & ~in1_0;
assign w2 = ~w0 & ~w1;
assign w3 = ~in0_2 & in1_2;
assign w4 = ~in0_1 & in1_1;
assign w5 = ~w3 & ~w4;
assign w6 = ~w2 & w5;
assign w7 = in0_5 & ~in1_5;
assign w8 = in0_4 & ~in1_4;
assign w9 = ~w7 & ~w8;
assign w10 = in0_3 & ~in1_3;
assign w11 = in0_2 & ~in1_2;
assign w12 = ~w10 & ~w11;
assign w13 = w9 & w12;
assign w14 = ~w6 & w13;
assign w15 = ~in0_4 & in1_4;
assign w16 = ~in0_3 & in1_3;
assign w17 = ~w15 & ~w16;
assign w18 = w9 & ~w17;
assign w19 = ~in0_8 & in1_8;
assign w20 = ~in0_7 & in1_7;
assign w21 = ~w19 & ~w20;
assign w22 = ~in0_6 & in1_6;
assign w23 = ~in0_5 & in1_5;
assign w24 = ~w22 & ~w23;
assign w25 = w21 & w24;
assign w26 = ~w18 & w25;
assign w27 = ~w14 & w26;
assign w28 = in0_9 & ~in1_9;
assign w29 = in0_7 & ~in1_7;
assign w30 = in0_6 & ~in1_6;
assign w31 = ~w29 & ~w30;
assign w32 = w21 & ~w31;
assign w33 = in0_11 & ~in1_11;
assign w34 = in0_10 & ~in1_10;
assign w35 = ~w33 & ~w34;
assign w36 = in0_8 & ~in1_8;
assign w37 = ~w28 & ~w36;
assign w38 = w35 & w37;
assign w39 = ~w32 & w38;
assign w40 = ~in0_12 & in1_12;
assign w41 = ~in0_10 & in1_10;
assign w42 = ~in0_9 & in1_9;
assign w43 = ~w41 & ~w42;
assign w44 = w35 & ~w43;
assign w45 = ~in0_14 & in1_14;
assign w46 = ~in0_13 & in1_13;
assign w47 = ~w45 & ~w46;
assign w48 = ~in0_11 & in1_11;
assign w49 = ~w40 & ~w48;
assign w50 = w47 & w49;
assign w51 = ~w44 & w50;
assign w52 = (w51 & w27) | (w51 & w3672) | (w27 & w3672);
assign w53 = in0_14 & ~in1_14;
assign w54 = in0_21 & ~in1_21;
assign w55 = ~in0_20 & in1_20;
assign w56 = ~in0_19 & in1_19;
assign w57 = ~w55 & ~w56;
assign w58 = in0_19 & ~in1_19;
assign w59 = in0_18 & ~in1_18;
assign w60 = ~w58 & ~w59;
assign w61 = w57 & ~w60;
assign w62 = in0_23 & ~in1_23;
assign w63 = in0_22 & ~in1_22;
assign w64 = ~w62 & ~w63;
assign w65 = in0_20 & ~in1_20;
assign w66 = ~w54 & ~w65;
assign w67 = w64 & w66;
assign w68 = ~w61 & w67;
assign w69 = in0_13 & ~in1_13;
assign w70 = in0_12 & ~in1_12;
assign w71 = ~w69 & ~w70;
assign w72 = w47 & ~w71;
assign w73 = in0_17 & ~in1_17;
assign w74 = in0_16 & ~in1_16;
assign w75 = ~w73 & ~w74;
assign w76 = in0_15 & ~in1_15;
assign w77 = ~w53 & ~w76;
assign w78 = w75 & w77;
assign w79 = ~w72 & w78;
assign w80 = w68 & w79;
assign w81 = ~w52 & w80;
assign w82 = ~in0_17 & in1_17;
assign w83 = ~in0_16 & in1_16;
assign w84 = ~in0_15 & in1_15;
assign w85 = ~w83 & ~w84;
assign w86 = w75 & ~w85;
assign w87 = ~in0_18 & in1_18;
assign w88 = ~w82 & ~w87;
assign w89 = w57 & w88;
assign w90 = ~w86 & w89;
assign w91 = w68 & ~w90;
assign w92 = ~in0_32 & in1_32;
assign w93 = ~in0_35 & in1_35;
assign w94 = ~in0_36 & in1_36;
assign w95 = ~in0_34 & in1_34;
assign w96 = ~in0_37 & in1_37;
assign w97 = ~in0_39 & in1_39;
assign w98 = ~in0_38 & in1_38;
assign w99 = ~w96 & ~w97;
assign w100 = ~w98 & w99;
assign w101 = ~w93 & ~w94;
assign w102 = ~w95 & w101;
assign w103 = w100 & w102;
assign w104 = ~w92 & w103;
assign w105 = ~in0_23 & in1_23;
assign w106 = in0_29 & ~in1_29;
assign w107 = in0_28 & ~in1_28;
assign w108 = ~w106 & ~w107;
assign w109 = ~in0_28 & in1_28;
assign w110 = ~in0_27 & in1_27;
assign w111 = ~w109 & ~w110;
assign w112 = w108 & ~w111;
assign w113 = ~in0_33 & in1_33;
assign w114 = ~in0_31 & in1_31;
assign w115 = ~w113 & ~w114;
assign w116 = ~in0_30 & in1_30;
assign w117 = ~in0_29 & in1_29;
assign w118 = ~w116 & ~w117;
assign w119 = w115 & w118;
assign w120 = ~w112 & w119;
assign w121 = ~in0_22 & in1_22;
assign w122 = ~in0_21 & in1_21;
assign w123 = ~w121 & ~w122;
assign w124 = w64 & ~w123;
assign w125 = ~in0_26 & in1_26;
assign w126 = ~in0_25 & in1_25;
assign w127 = ~w125 & ~w126;
assign w128 = ~in0_24 & in1_24;
assign w129 = ~w105 & ~w128;
assign w130 = w127 & w129;
assign w131 = ~w124 & w130;
assign w132 = w120 & w131;
assign w133 = ~w91 & w132;
assign w134 = w104 & w133;
assign w135 = ~w81 & w134;
assign w136 = in0_25 & ~in1_25;
assign w137 = in0_24 & ~in1_24;
assign w138 = ~w136 & ~w137;
assign w139 = w127 & ~w138;
assign w140 = in0_26 & ~in1_26;
assign w141 = in0_27 & ~in1_27;
assign w142 = ~w140 & ~w141;
assign w143 = w108 & w142;
assign w144 = ~w139 & w143;
assign w145 = w120 & ~w144;
assign w146 = in0_31 & ~in1_31;
assign w147 = in0_30 & ~in1_30;
assign w148 = ~w146 & ~w147;
assign w149 = w115 & ~w148;
assign w150 = ~w145 & ~w149;
assign w151 = w104 & ~w150;
assign w152 = ~in0_41 & in1_41;
assign w153 = in0_40 & ~in1_40;
assign w154 = ~w152 & w153;
assign w155 = in0_42 & ~in1_42;
assign w156 = in0_41 & ~in1_41;
assign w157 = ~w155 & ~w156;
assign w158 = ~w154 & w157;
assign w159 = ~in0_43 & in1_43;
assign w160 = ~in0_44 & in1_44;
assign w161 = ~in0_42 & in1_42;
assign w162 = ~w159 & ~w160;
assign w163 = ~w161 & w162;
assign w164 = ~w158 & w163;
assign w165 = in0_44 & ~in1_44;
assign w166 = in0_45 & ~in1_45;
assign w167 = in0_43 & ~in1_43;
assign w168 = ~w160 & w167;
assign w169 = ~w165 & ~w166;
assign w170 = ~w168 & w169;
assign w171 = ~in0_45 & in1_45;
assign w172 = ~in0_47 & in1_47;
assign w173 = ~in0_46 & in1_46;
assign w174 = ~w171 & ~w172;
assign w175 = ~w173 & w174;
assign w176 = (w175 & w164) | (w175 & w3673) | (w164 & w3673);
assign w177 = in0_47 & ~in1_47;
assign w178 = in0_46 & ~in1_46;
assign w179 = ~w172 & w178;
assign w180 = ~w177 & ~w179;
assign w181 = ~w176 & w180;
assign w182 = in0_34 & ~in1_34;
assign w183 = in0_33 & ~in1_33;
assign w184 = in0_32 & ~in1_32;
assign w185 = ~w113 & w184;
assign w186 = ~w182 & ~w183;
assign w187 = ~w185 & w186;
assign w188 = w103 & ~w187;
assign w189 = in0_37 & ~in1_37;
assign w190 = in0_36 & ~in1_36;
assign w191 = in0_35 & ~in1_35;
assign w192 = ~w94 & w191;
assign w193 = ~w189 & ~w190;
assign w194 = ~w192 & w193;
assign w195 = w100 & ~w194;
assign w196 = in0_39 & ~in1_39;
assign w197 = in0_38 & ~in1_38;
assign w198 = ~w97 & w197;
assign w199 = ~w196 & ~w198;
assign w200 = ~w195 & w199;
assign w201 = ~w188 & w200;
assign w202 = ~w151 & w3674;
assign w203 = ~w135 & w202;
assign w204 = ~in0_40 & in1_40;
assign w205 = ~w152 & ~w204;
assign w206 = w163 & w205;
assign w207 = w175 & w206;
assign w208 = ~in0_51 & in1_51;
assign w209 = ~in0_53 & in1_53;
assign w210 = ~in0_52 & in1_52;
assign w211 = ~w209 & ~w210;
assign w212 = ~in0_50 & in1_50;
assign w213 = ~w208 & ~w212;
assign w214 = w211 & w213;
assign w215 = ~in0_55 & in1_55;
assign w216 = ~in0_54 & in1_54;
assign w217 = ~w215 & ~w216;
assign w218 = ~in0_49 & in1_49;
assign w219 = ~in0_56 & in1_56;
assign w220 = ~in0_60 & in1_60;
assign w221 = ~in0_61 & in1_61;
assign w222 = ~in0_63 & in1_63;
assign w223 = ~in0_62 & in1_62;
assign w224 = ~w221 & ~w222;
assign w225 = ~w223 & w224;
assign w226 = w224 & w4919;
assign w227 = ~in0_59 & in1_59;
assign w228 = ~in0_58 & in1_58;
assign w229 = ~w227 & ~w228;
assign w230 = ~in0_57 & in1_57;
assign w231 = ~w219 & ~w230;
assign w232 = w229 & w231;
assign w233 = w226 & w232;
assign w234 = ~in0_48 & in1_48;
assign w235 = ~in0_70 & in1_70;
assign w236 = ~in0_71 & in1_71;
assign w237 = ~in0_69 & in1_69;
assign w238 = ~w235 & ~w236;
assign w239 = ~w237 & w238;
assign w240 = ~in0_68 & in1_68;
assign w241 = ~in0_72 & in1_72;
assign w242 = ~in0_75 & in1_75;
assign w243 = ~in0_74 & in1_74;
assign w244 = ~w242 & ~w243;
assign w245 = ~in0_73 & in1_73;
assign w246 = ~w241 & ~w245;
assign w247 = w244 & w246;
assign w248 = ~in0_76 & in1_76;
assign w249 = ~in0_78 & in1_78;
assign w250 = ~in0_79 & in1_79;
assign w251 = ~in0_77 & in1_77;
assign w252 = ~w249 & ~w250;
assign w253 = ~w251 & w252;
assign w254 = w252 & w4920;
assign w255 = in0_77 & ~in1_77;
assign w256 = in0_76 & ~in1_76;
assign w257 = ~w255 & ~w256;
assign w258 = w253 & ~w257;
assign w259 = in0_79 & ~in1_79;
assign w260 = in0_78 & ~in1_78;
assign w261 = ~w250 & w260;
assign w262 = ~w259 & ~w261;
assign w263 = ~w258 & w262;
assign w264 = ~w258 & w4921;
assign w265 = ~in0_81 & in1_81;
assign w266 = ~in0_87 & in1_87;
assign w267 = ~in0_85 & in1_85;
assign w268 = ~w266 & ~w267;
assign w269 = ~in0_86 & in1_86;
assign w270 = ~in0_84 & in1_84;
assign w271 = ~w269 & ~w270;
assign w272 = w268 & w271;
assign w273 = ~in0_83 & in1_83;
assign w274 = ~in0_82 & in1_82;
assign w275 = ~w273 & ~w274;
assign w276 = w272 & w275;
assign w277 = ~in0_80 & in1_80;
assign w278 = ~w265 & ~w277;
assign w279 = w272 & w4922;
assign w280 = ~w264 & w279;
assign w281 = in0_67 & ~in1_67;
assign w282 = ~in0_67 & in1_67;
assign w283 = ~in0_66 & in1_66;
assign w284 = ~w282 & ~w283;
assign w285 = in0_66 & ~in1_66;
assign w286 = in0_65 & ~in1_65;
assign w287 = ~in0_65 & in1_65;
assign w288 = in0_64 & ~in1_64;
assign w289 = ~w287 & w288;
assign w290 = ~w285 & ~w286;
assign w291 = ~w289 & w290;
assign w292 = (~w281 & w291) | (~w281 & w4923) | (w291 & w4923);
assign w293 = ~in0_64 & in1_64;
assign w294 = ~w287 & ~w293;
assign w295 = w284 & w294;
assign w296 = w292 & ~w295;
assign w297 = w238 & w4924;
assign w298 = w247 & w297;
assign w299 = ~w296 & w298;
assign w300 = w280 & w299;
assign w301 = ~w218 & ~w234;
assign w302 = w217 & w301;
assign w303 = w214 & w302;
assign w304 = w233 & w303;
assign w305 = (w304 & ~w181) | (w304 & w4925) | (~w181 & w4925);
assign w306 = w300 & w305;
assign w307 = ~w203 & w306;
assign w308 = in0_55 & ~in1_55;
assign w309 = ~w217 & ~w308;
assign w310 = in0_50 & ~in1_50;
assign w311 = in0_49 & ~in1_49;
assign w312 = in0_48 & ~in1_48;
assign w313 = ~w218 & w312;
assign w314 = ~w310 & ~w311;
assign w315 = ~w313 & w314;
assign w316 = w214 & ~w315;
assign w317 = in0_52 & ~in1_52;
assign w318 = in0_51 & ~in1_51;
assign w319 = ~w317 & ~w318;
assign w320 = w211 & ~w319;
assign w321 = in0_53 & ~in1_53;
assign w322 = in0_54 & ~in1_54;
assign w323 = ~w308 & ~w321;
assign w324 = ~w322 & w323;
assign w325 = ~w320 & w324;
assign w326 = ~w316 & w325;
assign w327 = w233 & ~w309;
assign w328 = ~w326 & w327;
assign w329 = in0_59 & ~in1_59;
assign w330 = in0_58 & ~in1_58;
assign w331 = in0_57 & ~in1_57;
assign w332 = in0_56 & ~in1_56;
assign w333 = ~w230 & w332;
assign w334 = ~w330 & ~w331;
assign w335 = ~w333 & w334;
assign w336 = (~w329 & w335) | (~w329 & w4926) | (w335 & w4926);
assign w337 = w226 & ~w336;
assign w338 = in0_63 & ~in1_63;
assign w339 = in0_61 & ~in1_61;
assign w340 = in0_60 & ~in1_60;
assign w341 = ~w339 & ~w340;
assign w342 = w225 & ~w341;
assign w343 = in0_62 & ~in1_62;
assign w344 = ~w222 & w343;
assign w345 = ~w338 & ~w344;
assign w346 = ~w342 & w345;
assign w347 = w292 & w346;
assign w348 = ~w337 & w347;
assign w349 = ~w328 & w348;
assign w350 = w300 & ~w349;
assign w351 = ~in0_108 & in1_108;
assign w352 = ~in0_109 & in1_109;
assign w353 = ~in0_111 & in1_111;
assign w354 = ~in0_110 & in1_110;
assign w355 = ~w352 & ~w353;
assign w356 = ~w354 & w355;
assign w357 = w355 & w4927;
assign w358 = in0_107 & ~in1_107;
assign w359 = ~in0_107 & in1_107;
assign w360 = ~in0_106 & in1_106;
assign w361 = ~w359 & ~w360;
assign w362 = in0_106 & ~in1_106;
assign w363 = in0_105 & ~in1_105;
assign w364 = ~in0_105 & in1_105;
assign w365 = in0_104 & ~in1_104;
assign w366 = ~w364 & w365;
assign w367 = ~w362 & ~w363;
assign w368 = ~w366 & w367;
assign w369 = (~w358 & w368) | (~w358 & w3675) | (w368 & w3675);
assign w370 = w357 & ~w369;
assign w371 = in0_111 & ~in1_111;
assign w372 = in0_115 & ~in1_115;
assign w373 = ~in0_115 & in1_115;
assign w374 = ~in0_114 & in1_114;
assign w375 = ~w373 & ~w374;
assign w376 = ~in0_113 & in1_113;
assign w377 = in0_112 & ~in1_112;
assign w378 = ~w376 & w377;
assign w379 = in0_114 & ~in1_114;
assign w380 = in0_113 & ~in1_113;
assign w381 = ~w379 & ~w380;
assign w382 = ~w378 & w381;
assign w383 = (~w372 & w382) | (~w372 & w3676) | (w382 & w3676);
assign w384 = in0_109 & ~in1_109;
assign w385 = in0_108 & ~in1_108;
assign w386 = ~w384 & ~w385;
assign w387 = w356 & ~w386;
assign w388 = in0_110 & ~in1_110;
assign w389 = ~w353 & w388;
assign w390 = ~w371 & ~w389;
assign w391 = ~w387 & w390;
assign w392 = w383 & w391;
assign w393 = ~w370 & w392;
assign w394 = ~in0_112 & in1_112;
assign w395 = ~w376 & ~w394;
assign w396 = w375 & w395;
assign w397 = w383 & ~w396;
assign w398 = ~in0_119 & in1_119;
assign w399 = ~in0_121 & in1_121;
assign w400 = ~in0_123 & in1_123;
assign w401 = ~in0_122 & in1_122;
assign w402 = ~w400 & ~w401;
assign w403 = ~in0_120 & in1_120;
assign w404 = ~w399 & ~w403;
assign w405 = w402 & w404;
assign w406 = ~in0_118 & in1_118;
assign w407 = ~in0_117 & in1_117;
assign w408 = ~w406 & ~w407;
assign w409 = ~in0_116 & in1_116;
assign w410 = ~w398 & ~w409;
assign w411 = w408 & w410;
assign w412 = w405 & w411;
assign w413 = ~w397 & w412;
assign w414 = ~w393 & w413;
assign w415 = in0_69 & ~in1_69;
assign w416 = in0_68 & ~in1_68;
assign w417 = ~w415 & ~w416;
assign w418 = w239 & ~w417;
assign w419 = in0_71 & ~in1_71;
assign w420 = in0_70 & ~in1_70;
assign w421 = ~w236 & w420;
assign w422 = ~w419 & ~w421;
assign w423 = (w247 & w418) | (w247 & w4928) | (w418 & w4928);
assign w424 = in0_72 & ~in1_72;
assign w425 = ~w245 & w424;
assign w426 = in0_74 & ~in1_74;
assign w427 = in0_73 & ~in1_73;
assign w428 = ~w426 & ~w427;
assign w429 = ~w425 & w428;
assign w430 = in0_75 & ~in1_75;
assign w431 = (~w430 & w429) | (~w430 & w4929) | (w429 & w4929);
assign w432 = w263 & w431;
assign w433 = ~w423 & w432;
assign w434 = w280 & ~w433;
assign w435 = in0_93 & ~in1_93;
assign w436 = in0_92 & ~in1_92;
assign w437 = ~w435 & ~w436;
assign w438 = ~in0_94 & in1_94;
assign w439 = ~in0_95 & in1_95;
assign w440 = ~in0_93 & in1_93;
assign w441 = ~w438 & ~w439;
assign w442 = ~w440 & w441;
assign w443 = ~w437 & w442;
assign w444 = in0_95 & ~in1_95;
assign w445 = in0_94 & ~in1_94;
assign w446 = ~w439 & w445;
assign w447 = ~w444 & ~w446;
assign w448 = ~in0_96 & in1_96;
assign w449 = ~in0_99 & in1_99;
assign w450 = ~in0_98 & in1_98;
assign w451 = ~w449 & ~w450;
assign w452 = ~in0_97 & in1_97;
assign w453 = ~w448 & ~w452;
assign w454 = w451 & w453;
assign w455 = (w454 & w443) | (w454 & w3677) | (w443 & w3677);
assign w456 = in0_101 & ~in1_101;
assign w457 = in0_100 & ~in1_100;
assign w458 = ~w456 & ~w457;
assign w459 = ~in0_102 & in1_102;
assign w460 = ~in0_103 & in1_103;
assign w461 = ~in0_101 & in1_101;
assign w462 = ~w459 & ~w460;
assign w463 = ~w461 & w462;
assign w464 = ~w458 & w463;
assign w465 = in0_103 & ~in1_103;
assign w466 = in0_102 & ~in1_102;
assign w467 = ~w460 & w466;
assign w468 = ~w465 & ~w467;
assign w469 = ~w464 & w468;
assign w470 = in0_99 & ~in1_99;
assign w471 = in0_96 & ~in1_96;
assign w472 = ~w452 & w471;
assign w473 = in0_98 & ~in1_98;
assign w474 = in0_97 & ~in1_97;
assign w475 = ~w473 & ~w474;
assign w476 = ~w472 & w475;
assign w477 = (~w470 & w476) | (~w470 & w3678) | (w476 & w3678);
assign w478 = w469 & w477;
assign w479 = ~w455 & w478;
assign w480 = in0_82 & ~in1_82;
assign w481 = in0_81 & ~in1_81;
assign w482 = in0_80 & ~in1_80;
assign w483 = ~w265 & w482;
assign w484 = ~w480 & ~w481;
assign w485 = ~w483 & w484;
assign w486 = w276 & ~w485;
assign w487 = in0_91 & ~in1_91;
assign w488 = ~in0_91 & in1_91;
assign w489 = ~in0_90 & in1_90;
assign w490 = ~w488 & ~w489;
assign w491 = ~in0_89 & in1_89;
assign w492 = in0_88 & ~in1_88;
assign w493 = ~w491 & w492;
assign w494 = in0_90 & ~in1_90;
assign w495 = in0_89 & ~in1_89;
assign w496 = ~w494 & ~w495;
assign w497 = ~w493 & w496;
assign w498 = (~w487 & w497) | (~w487 & w3679) | (w497 & w3679);
assign w499 = in0_83 & ~in1_83;
assign w500 = w272 & w499;
assign w501 = in0_87 & ~in1_87;
assign w502 = in0_86 & ~in1_86;
assign w503 = ~w266 & w502;
assign w504 = in0_85 & ~in1_85;
assign w505 = in0_84 & ~in1_84;
assign w506 = ~w504 & ~w505;
assign w507 = w268 & ~w269;
assign w508 = ~w506 & w507;
assign w509 = ~w501 & ~w503;
assign w510 = ~w500 & w509;
assign w511 = ~w508 & w510;
assign w512 = ~w486 & w498;
assign w513 = w511 & w512;
assign w514 = w479 & w513;
assign w515 = ~w414 & w514;
assign w516 = ~w434 & w515;
assign w517 = ~w350 & w516;
assign w518 = ~w307 & w517;
assign w519 = ~in0_88 & in1_88;
assign w520 = ~w491 & ~w519;
assign w521 = w490 & w520;
assign w522 = w498 & ~w521;
assign w523 = ~in0_92 & in1_92;
assign w524 = w441 & w4930;
assign w525 = w454 & w524;
assign w526 = ~w522 & w525;
assign w527 = w479 & ~w526;
assign w528 = ~in0_100 & in1_100;
assign w529 = w462 & w4931;
assign w530 = ~w464 & w4932;
assign w531 = ~in0_104 & in1_104;
assign w532 = ~w364 & ~w531;
assign w533 = w361 & w532;
assign w534 = w357 & w533;
assign w535 = ~w530 & w534;
assign w536 = w413 & w535;
assign w537 = ~w527 & w536;
assign w538 = ~in0_124 & in1_124;
assign w539 = ~in0_125 & in1_125;
assign w540 = in0_127 & ~in1_127;
assign w541 = ~in0_126 & in1_126;
assign w542 = ~w539 & ~w540;
assign w543 = ~w541 & w542;
assign w544 = w542 & w4933;
assign w545 = (w544 & w537) | (w544 & w3680) | (w537 & w3680);
assign w546 = (w545 & ~w517) | (w545 & w4934) | (~w517 & w4934);
assign w547 = in0_123 & ~in1_123;
assign w548 = in0_119 & ~in1_119;
assign w549 = in0_118 & ~in1_118;
assign w550 = in0_117 & ~in1_117;
assign w551 = in0_116 & ~in1_116;
assign w552 = ~w550 & ~w551;
assign w553 = w408 & ~w552;
assign w554 = in0_120 & ~in1_120;
assign w555 = ~w548 & ~w554;
assign w556 = w555 & w7147;
assign w557 = w405 & ~w556;
assign w558 = in0_122 & ~in1_122;
assign w559 = in0_121 & ~in1_121;
assign w560 = ~w558 & ~w559;
assign w561 = w402 & ~w560;
assign w562 = ~w547 & ~w561;
assign w563 = (w544 & w557) | (w544 & w4935) | (w557 & w4935);
assign w564 = ~in0_127 & in1_127;
assign w565 = in0_125 & ~in1_125;
assign w566 = in0_124 & ~in1_124;
assign w567 = ~w565 & ~w566;
assign w568 = w543 & ~w567;
assign w569 = in0_126 & ~in1_126;
assign w570 = ~w540 & w569;
assign w571 = ~w564 & ~w570;
assign w572 = ~w568 & w571;
assign w573 = ~w563 & w572;
assign w574 = ~w563 & w4936;
assign w575 = (w517 & w5447) | (w517 & w5448) | (w5447 & w5448);
assign w576 = (in0_0 & w563) | (in0_0 & w4937) | (w563 & w4937);
assign w577 = (w517 & w6864) | (w517 & w6865) | (w6864 & w6865);
assign w578 = ~w575 & w577;
assign w579 = in2_1 & ~in3_1;
assign w580 = in2_0 & ~in3_0;
assign w581 = ~w579 & ~w580;
assign w582 = ~in2_2 & in3_2;
assign w583 = ~in2_1 & in3_1;
assign w584 = ~w582 & ~w583;
assign w585 = ~w581 & w584;
assign w586 = in2_5 & ~in3_5;
assign w587 = in2_4 & ~in3_4;
assign w588 = ~w586 & ~w587;
assign w589 = in2_3 & ~in3_3;
assign w590 = in2_2 & ~in3_2;
assign w591 = ~w589 & ~w590;
assign w592 = w588 & w591;
assign w593 = ~w585 & w592;
assign w594 = ~in2_4 & in3_4;
assign w595 = ~in2_3 & in3_3;
assign w596 = ~w594 & ~w595;
assign w597 = w588 & ~w596;
assign w598 = ~in2_8 & in3_8;
assign w599 = ~in2_7 & in3_7;
assign w600 = ~w598 & ~w599;
assign w601 = ~in2_6 & in3_6;
assign w602 = ~in2_5 & in3_5;
assign w603 = ~w601 & ~w602;
assign w604 = w600 & w603;
assign w605 = ~w597 & w604;
assign w606 = ~w593 & w605;
assign w607 = in2_9 & ~in3_9;
assign w608 = in2_7 & ~in3_7;
assign w609 = in2_6 & ~in3_6;
assign w610 = ~w608 & ~w609;
assign w611 = w600 & ~w610;
assign w612 = in2_11 & ~in3_11;
assign w613 = in2_10 & ~in3_10;
assign w614 = ~w612 & ~w613;
assign w615 = in2_8 & ~in3_8;
assign w616 = ~w607 & ~w615;
assign w617 = w614 & w616;
assign w618 = ~w611 & w617;
assign w619 = ~in2_12 & in3_12;
assign w620 = ~in2_10 & in3_10;
assign w621 = ~in2_9 & in3_9;
assign w622 = ~w620 & ~w621;
assign w623 = w614 & ~w622;
assign w624 = ~in2_14 & in3_14;
assign w625 = ~in2_13 & in3_13;
assign w626 = ~w624 & ~w625;
assign w627 = ~in2_11 & in3_11;
assign w628 = ~w619 & ~w627;
assign w629 = w626 & w628;
assign w630 = ~w623 & w629;
assign w631 = (w630 & w606) | (w630 & w3683) | (w606 & w3683);
assign w632 = in2_14 & ~in3_14;
assign w633 = in2_21 & ~in3_21;
assign w634 = ~in2_20 & in3_20;
assign w635 = ~in2_19 & in3_19;
assign w636 = ~w634 & ~w635;
assign w637 = in2_19 & ~in3_19;
assign w638 = in2_18 & ~in3_18;
assign w639 = ~w637 & ~w638;
assign w640 = w636 & ~w639;
assign w641 = in2_23 & ~in3_23;
assign w642 = in2_22 & ~in3_22;
assign w643 = ~w641 & ~w642;
assign w644 = in2_20 & ~in3_20;
assign w645 = ~w633 & ~w644;
assign w646 = w643 & w645;
assign w647 = ~w640 & w646;
assign w648 = in2_13 & ~in3_13;
assign w649 = in2_12 & ~in3_12;
assign w650 = ~w648 & ~w649;
assign w651 = w626 & ~w650;
assign w652 = in2_17 & ~in3_17;
assign w653 = in2_16 & ~in3_16;
assign w654 = ~w652 & ~w653;
assign w655 = in2_15 & ~in3_15;
assign w656 = ~w632 & ~w655;
assign w657 = w654 & w656;
assign w658 = ~w651 & w657;
assign w659 = w647 & w658;
assign w660 = ~w631 & w659;
assign w661 = ~in2_18 & in3_18;
assign w662 = ~in2_16 & in3_16;
assign w663 = ~in2_15 & in3_15;
assign w664 = ~w662 & ~w663;
assign w665 = w654 & ~w664;
assign w666 = ~in2_17 & in3_17;
assign w667 = ~w661 & ~w666;
assign w668 = w636 & w667;
assign w669 = ~w665 & w668;
assign w670 = w647 & ~w669;
assign w671 = ~in2_32 & in3_32;
assign w672 = ~in2_35 & in3_35;
assign w673 = ~in2_36 & in3_36;
assign w674 = ~in2_34 & in3_34;
assign w675 = ~in2_37 & in3_37;
assign w676 = ~in2_39 & in3_39;
assign w677 = ~in2_38 & in3_38;
assign w678 = ~w675 & ~w676;
assign w679 = ~w677 & w678;
assign w680 = ~w672 & ~w673;
assign w681 = ~w674 & w680;
assign w682 = w679 & w681;
assign w683 = ~w671 & w682;
assign w684 = ~in2_23 & in3_23;
assign w685 = in2_29 & ~in3_29;
assign w686 = in2_28 & ~in3_28;
assign w687 = ~w685 & ~w686;
assign w688 = ~in2_28 & in3_28;
assign w689 = ~in2_27 & in3_27;
assign w690 = ~w688 & ~w689;
assign w691 = w687 & ~w690;
assign w692 = ~in2_33 & in3_33;
assign w693 = ~in2_31 & in3_31;
assign w694 = ~w692 & ~w693;
assign w695 = ~in2_30 & in3_30;
assign w696 = ~in2_29 & in3_29;
assign w697 = ~w695 & ~w696;
assign w698 = w694 & w697;
assign w699 = ~w691 & w698;
assign w700 = ~in2_22 & in3_22;
assign w701 = ~in2_21 & in3_21;
assign w702 = ~w700 & ~w701;
assign w703 = w643 & ~w702;
assign w704 = ~in2_26 & in3_26;
assign w705 = ~in2_25 & in3_25;
assign w706 = ~w704 & ~w705;
assign w707 = ~in2_24 & in3_24;
assign w708 = ~w684 & ~w707;
assign w709 = w706 & w708;
assign w710 = ~w703 & w709;
assign w711 = w699 & w710;
assign w712 = ~w670 & w711;
assign w713 = w683 & w712;
assign w714 = ~w660 & w713;
assign w715 = in2_25 & ~in3_25;
assign w716 = in2_24 & ~in3_24;
assign w717 = ~w715 & ~w716;
assign w718 = w706 & ~w717;
assign w719 = in2_26 & ~in3_26;
assign w720 = in2_27 & ~in3_27;
assign w721 = ~w719 & ~w720;
assign w722 = w687 & w721;
assign w723 = ~w718 & w722;
assign w724 = w699 & ~w723;
assign w725 = in2_31 & ~in3_31;
assign w726 = in2_30 & ~in3_30;
assign w727 = ~w725 & ~w726;
assign w728 = w694 & ~w727;
assign w729 = ~w724 & ~w728;
assign w730 = w683 & ~w729;
assign w731 = ~in2_41 & in3_41;
assign w732 = in2_40 & ~in3_40;
assign w733 = ~w731 & w732;
assign w734 = in2_42 & ~in3_42;
assign w735 = in2_41 & ~in3_41;
assign w736 = ~w734 & ~w735;
assign w737 = ~w733 & w736;
assign w738 = ~in2_43 & in3_43;
assign w739 = ~in2_44 & in3_44;
assign w740 = ~in2_42 & in3_42;
assign w741 = ~w738 & ~w739;
assign w742 = ~w740 & w741;
assign w743 = ~w737 & w742;
assign w744 = in2_44 & ~in3_44;
assign w745 = in2_45 & ~in3_45;
assign w746 = in2_43 & ~in3_43;
assign w747 = ~w739 & w746;
assign w748 = ~w744 & ~w745;
assign w749 = ~w747 & w748;
assign w750 = ~in2_45 & in3_45;
assign w751 = ~in2_47 & in3_47;
assign w752 = ~in2_46 & in3_46;
assign w753 = ~w750 & ~w751;
assign w754 = ~w752 & w753;
assign w755 = (w754 & w743) | (w754 & w3684) | (w743 & w3684);
assign w756 = in2_47 & ~in3_47;
assign w757 = in2_46 & ~in3_46;
assign w758 = ~w751 & w757;
assign w759 = ~w756 & ~w758;
assign w760 = ~w755 & w759;
assign w761 = in2_34 & ~in3_34;
assign w762 = in2_33 & ~in3_33;
assign w763 = in2_32 & ~in3_32;
assign w764 = ~w692 & w763;
assign w765 = ~w761 & ~w762;
assign w766 = ~w764 & w765;
assign w767 = w682 & ~w766;
assign w768 = in2_37 & ~in3_37;
assign w769 = in2_36 & ~in3_36;
assign w770 = in2_35 & ~in3_35;
assign w771 = ~w673 & w770;
assign w772 = ~w768 & ~w769;
assign w773 = ~w771 & w772;
assign w774 = w679 & ~w773;
assign w775 = in2_39 & ~in3_39;
assign w776 = in2_38 & ~in3_38;
assign w777 = ~w676 & w776;
assign w778 = ~w775 & ~w777;
assign w779 = ~w774 & w778;
assign w780 = ~w767 & w779;
assign w781 = ~w730 & w3685;
assign w782 = ~w714 & w781;
assign w783 = ~in2_40 & in3_40;
assign w784 = ~w731 & ~w783;
assign w785 = w742 & w784;
assign w786 = w754 & w785;
assign w787 = ~in2_51 & in3_51;
assign w788 = ~in2_53 & in3_53;
assign w789 = ~in2_52 & in3_52;
assign w790 = ~w788 & ~w789;
assign w791 = ~in2_50 & in3_50;
assign w792 = ~w787 & ~w791;
assign w793 = w790 & w792;
assign w794 = ~in2_55 & in3_55;
assign w795 = ~in2_54 & in3_54;
assign w796 = ~w794 & ~w795;
assign w797 = ~in2_49 & in3_49;
assign w798 = ~in2_56 & in3_56;
assign w799 = ~in2_60 & in3_60;
assign w800 = ~in2_61 & in3_61;
assign w801 = ~in2_63 & in3_63;
assign w802 = ~in2_62 & in3_62;
assign w803 = ~w800 & ~w801;
assign w804 = ~w802 & w803;
assign w805 = w803 & w4938;
assign w806 = ~in2_59 & in3_59;
assign w807 = ~in2_58 & in3_58;
assign w808 = ~w806 & ~w807;
assign w809 = ~in2_57 & in3_57;
assign w810 = ~w798 & ~w809;
assign w811 = w808 & w810;
assign w812 = w805 & w811;
assign w813 = ~in2_48 & in3_48;
assign w814 = ~in2_70 & in3_70;
assign w815 = ~in2_71 & in3_71;
assign w816 = ~in2_69 & in3_69;
assign w817 = ~w814 & ~w815;
assign w818 = ~w816 & w817;
assign w819 = ~in2_68 & in3_68;
assign w820 = ~in2_72 & in3_72;
assign w821 = ~in2_75 & in3_75;
assign w822 = ~in2_74 & in3_74;
assign w823 = ~w821 & ~w822;
assign w824 = ~in2_73 & in3_73;
assign w825 = ~w820 & ~w824;
assign w826 = w823 & w825;
assign w827 = ~in2_76 & in3_76;
assign w828 = ~in2_78 & in3_78;
assign w829 = ~in2_79 & in3_79;
assign w830 = ~in2_77 & in3_77;
assign w831 = ~w828 & ~w829;
assign w832 = ~w830 & w831;
assign w833 = w831 & w4939;
assign w834 = in2_77 & ~in3_77;
assign w835 = in2_76 & ~in3_76;
assign w836 = ~w834 & ~w835;
assign w837 = w832 & ~w836;
assign w838 = in2_79 & ~in3_79;
assign w839 = in2_78 & ~in3_78;
assign w840 = ~w829 & w839;
assign w841 = ~w838 & ~w840;
assign w842 = ~w837 & w841;
assign w843 = ~w837 & w4940;
assign w844 = ~in2_81 & in3_81;
assign w845 = ~in2_87 & in3_87;
assign w846 = ~in2_85 & in3_85;
assign w847 = ~w845 & ~w846;
assign w848 = ~in2_86 & in3_86;
assign w849 = ~in2_84 & in3_84;
assign w850 = ~w848 & ~w849;
assign w851 = w847 & w850;
assign w852 = ~in2_83 & in3_83;
assign w853 = ~in2_82 & in3_82;
assign w854 = ~w852 & ~w853;
assign w855 = w851 & w854;
assign w856 = ~in2_80 & in3_80;
assign w857 = ~w844 & ~w856;
assign w858 = w851 & w4941;
assign w859 = ~w843 & w858;
assign w860 = in2_67 & ~in3_67;
assign w861 = ~in2_67 & in3_67;
assign w862 = ~in2_66 & in3_66;
assign w863 = ~w861 & ~w862;
assign w864 = in2_66 & ~in3_66;
assign w865 = in2_65 & ~in3_65;
assign w866 = ~in2_65 & in3_65;
assign w867 = in2_64 & ~in3_64;
assign w868 = ~w866 & w867;
assign w869 = ~w864 & ~w865;
assign w870 = ~w868 & w869;
assign w871 = (~w860 & w870) | (~w860 & w4942) | (w870 & w4942);
assign w872 = ~in2_64 & in3_64;
assign w873 = ~w866 & ~w872;
assign w874 = w863 & w873;
assign w875 = w871 & ~w874;
assign w876 = w817 & w4943;
assign w877 = w826 & w876;
assign w878 = ~w875 & w877;
assign w879 = w859 & w878;
assign w880 = ~w797 & ~w813;
assign w881 = w796 & w880;
assign w882 = w793 & w881;
assign w883 = w812 & w882;
assign w884 = (w883 & ~w760) | (w883 & w4944) | (~w760 & w4944);
assign w885 = w879 & w884;
assign w886 = ~w782 & w885;
assign w887 = in2_55 & ~in3_55;
assign w888 = ~w796 & ~w887;
assign w889 = in2_50 & ~in3_50;
assign w890 = in2_49 & ~in3_49;
assign w891 = in2_48 & ~in3_48;
assign w892 = ~w797 & w891;
assign w893 = ~w889 & ~w890;
assign w894 = ~w892 & w893;
assign w895 = w793 & ~w894;
assign w896 = in2_52 & ~in3_52;
assign w897 = in2_51 & ~in3_51;
assign w898 = ~w896 & ~w897;
assign w899 = w790 & ~w898;
assign w900 = in2_53 & ~in3_53;
assign w901 = in2_54 & ~in3_54;
assign w902 = ~w887 & ~w900;
assign w903 = ~w901 & w902;
assign w904 = ~w899 & w903;
assign w905 = ~w895 & w904;
assign w906 = w812 & ~w888;
assign w907 = ~w905 & w906;
assign w908 = in2_59 & ~in3_59;
assign w909 = in2_58 & ~in3_58;
assign w910 = in2_57 & ~in3_57;
assign w911 = in2_56 & ~in3_56;
assign w912 = ~w809 & w911;
assign w913 = ~w909 & ~w910;
assign w914 = ~w912 & w913;
assign w915 = (~w908 & w914) | (~w908 & w4945) | (w914 & w4945);
assign w916 = w805 & ~w915;
assign w917 = in2_63 & ~in3_63;
assign w918 = in2_61 & ~in3_61;
assign w919 = in2_60 & ~in3_60;
assign w920 = ~w918 & ~w919;
assign w921 = w804 & ~w920;
assign w922 = in2_62 & ~in3_62;
assign w923 = ~w801 & w922;
assign w924 = ~w917 & ~w923;
assign w925 = ~w921 & w924;
assign w926 = w871 & w925;
assign w927 = ~w916 & w926;
assign w928 = ~w907 & w927;
assign w929 = w879 & ~w928;
assign w930 = ~in2_108 & in3_108;
assign w931 = ~in2_109 & in3_109;
assign w932 = ~in2_111 & in3_111;
assign w933 = ~in2_110 & in3_110;
assign w934 = ~w931 & ~w932;
assign w935 = ~w933 & w934;
assign w936 = w934 & w4946;
assign w937 = in2_107 & ~in3_107;
assign w938 = ~in2_107 & in3_107;
assign w939 = ~in2_106 & in3_106;
assign w940 = ~w938 & ~w939;
assign w941 = in2_106 & ~in3_106;
assign w942 = in2_105 & ~in3_105;
assign w943 = ~in2_105 & in3_105;
assign w944 = in2_104 & ~in3_104;
assign w945 = ~w943 & w944;
assign w946 = ~w941 & ~w942;
assign w947 = ~w945 & w946;
assign w948 = (~w937 & w947) | (~w937 & w3686) | (w947 & w3686);
assign w949 = w936 & ~w948;
assign w950 = in2_111 & ~in3_111;
assign w951 = in2_115 & ~in3_115;
assign w952 = ~in2_115 & in3_115;
assign w953 = ~in2_114 & in3_114;
assign w954 = ~w952 & ~w953;
assign w955 = ~in2_113 & in3_113;
assign w956 = in2_112 & ~in3_112;
assign w957 = ~w955 & w956;
assign w958 = in2_114 & ~in3_114;
assign w959 = in2_113 & ~in3_113;
assign w960 = ~w958 & ~w959;
assign w961 = ~w957 & w960;
assign w962 = (~w951 & w961) | (~w951 & w3687) | (w961 & w3687);
assign w963 = in2_109 & ~in3_109;
assign w964 = in2_108 & ~in3_108;
assign w965 = ~w963 & ~w964;
assign w966 = w935 & ~w965;
assign w967 = in2_110 & ~in3_110;
assign w968 = ~w932 & w967;
assign w969 = ~w950 & ~w968;
assign w970 = ~w966 & w969;
assign w971 = w962 & w970;
assign w972 = ~w949 & w971;
assign w973 = ~in2_112 & in3_112;
assign w974 = ~w955 & ~w973;
assign w975 = w954 & w974;
assign w976 = w962 & ~w975;
assign w977 = ~in2_119 & in3_119;
assign w978 = ~in2_121 & in3_121;
assign w979 = ~in2_123 & in3_123;
assign w980 = ~in2_122 & in3_122;
assign w981 = ~w979 & ~w980;
assign w982 = ~in2_120 & in3_120;
assign w983 = ~w978 & ~w982;
assign w984 = w981 & w983;
assign w985 = ~in2_118 & in3_118;
assign w986 = ~in2_117 & in3_117;
assign w987 = ~w985 & ~w986;
assign w988 = ~in2_116 & in3_116;
assign w989 = ~w977 & ~w988;
assign w990 = w987 & w989;
assign w991 = w984 & w990;
assign w992 = ~w976 & w991;
assign w993 = ~w972 & w992;
assign w994 = in2_69 & ~in3_69;
assign w995 = in2_68 & ~in3_68;
assign w996 = ~w994 & ~w995;
assign w997 = w818 & ~w996;
assign w998 = in2_71 & ~in3_71;
assign w999 = in2_70 & ~in3_70;
assign w1000 = ~w815 & w999;
assign w1001 = ~w998 & ~w1000;
assign w1002 = (w826 & w997) | (w826 & w4947) | (w997 & w4947);
assign w1003 = in2_72 & ~in3_72;
assign w1004 = ~w824 & w1003;
assign w1005 = in2_74 & ~in3_74;
assign w1006 = in2_73 & ~in3_73;
assign w1007 = ~w1005 & ~w1006;
assign w1008 = ~w1004 & w1007;
assign w1009 = in2_75 & ~in3_75;
assign w1010 = (~w1009 & w1008) | (~w1009 & w4948) | (w1008 & w4948);
assign w1011 = w842 & w1010;
assign w1012 = ~w1002 & w1011;
assign w1013 = w859 & ~w1012;
assign w1014 = in2_93 & ~in3_93;
assign w1015 = in2_92 & ~in3_92;
assign w1016 = ~w1014 & ~w1015;
assign w1017 = ~in2_94 & in3_94;
assign w1018 = ~in2_95 & in3_95;
assign w1019 = ~in2_93 & in3_93;
assign w1020 = ~w1017 & ~w1018;
assign w1021 = ~w1019 & w1020;
assign w1022 = ~w1016 & w1021;
assign w1023 = in2_95 & ~in3_95;
assign w1024 = in2_94 & ~in3_94;
assign w1025 = ~w1018 & w1024;
assign w1026 = ~w1023 & ~w1025;
assign w1027 = ~in2_96 & in3_96;
assign w1028 = ~in2_99 & in3_99;
assign w1029 = ~in2_98 & in3_98;
assign w1030 = ~w1028 & ~w1029;
assign w1031 = ~in2_97 & in3_97;
assign w1032 = ~w1027 & ~w1031;
assign w1033 = w1030 & w1032;
assign w1034 = (w1033 & w1022) | (w1033 & w3688) | (w1022 & w3688);
assign w1035 = in2_101 & ~in3_101;
assign w1036 = in2_100 & ~in3_100;
assign w1037 = ~w1035 & ~w1036;
assign w1038 = ~in2_102 & in3_102;
assign w1039 = ~in2_103 & in3_103;
assign w1040 = ~in2_101 & in3_101;
assign w1041 = ~w1038 & ~w1039;
assign w1042 = ~w1040 & w1041;
assign w1043 = ~w1037 & w1042;
assign w1044 = in2_103 & ~in3_103;
assign w1045 = in2_102 & ~in3_102;
assign w1046 = ~w1039 & w1045;
assign w1047 = ~w1044 & ~w1046;
assign w1048 = ~w1043 & w1047;
assign w1049 = in2_99 & ~in3_99;
assign w1050 = in2_96 & ~in3_96;
assign w1051 = ~w1031 & w1050;
assign w1052 = in2_98 & ~in3_98;
assign w1053 = in2_97 & ~in3_97;
assign w1054 = ~w1052 & ~w1053;
assign w1055 = ~w1051 & w1054;
assign w1056 = (~w1049 & w1055) | (~w1049 & w3689) | (w1055 & w3689);
assign w1057 = w1048 & w1056;
assign w1058 = ~w1034 & w1057;
assign w1059 = in2_82 & ~in3_82;
assign w1060 = in2_81 & ~in3_81;
assign w1061 = in2_80 & ~in3_80;
assign w1062 = ~w844 & w1061;
assign w1063 = ~w1059 & ~w1060;
assign w1064 = ~w1062 & w1063;
assign w1065 = w855 & ~w1064;
assign w1066 = in2_91 & ~in3_91;
assign w1067 = ~in2_91 & in3_91;
assign w1068 = ~in2_90 & in3_90;
assign w1069 = ~w1067 & ~w1068;
assign w1070 = ~in2_89 & in3_89;
assign w1071 = in2_88 & ~in3_88;
assign w1072 = ~w1070 & w1071;
assign w1073 = in2_90 & ~in3_90;
assign w1074 = in2_89 & ~in3_89;
assign w1075 = ~w1073 & ~w1074;
assign w1076 = ~w1072 & w1075;
assign w1077 = (~w1066 & w1076) | (~w1066 & w3690) | (w1076 & w3690);
assign w1078 = in2_83 & ~in3_83;
assign w1079 = w851 & w1078;
assign w1080 = in2_87 & ~in3_87;
assign w1081 = in2_86 & ~in3_86;
assign w1082 = ~w845 & w1081;
assign w1083 = in2_85 & ~in3_85;
assign w1084 = in2_84 & ~in3_84;
assign w1085 = ~w1083 & ~w1084;
assign w1086 = w847 & ~w848;
assign w1087 = ~w1085 & w1086;
assign w1088 = ~w1080 & ~w1082;
assign w1089 = ~w1079 & w1088;
assign w1090 = ~w1087 & w1089;
assign w1091 = ~w1065 & w1077;
assign w1092 = w1090 & w1091;
assign w1093 = w1058 & w1092;
assign w1094 = ~w993 & w1093;
assign w1095 = ~w1013 & w1094;
assign w1096 = ~w929 & w1095;
assign w1097 = ~w886 & w1096;
assign w1098 = ~in2_124 & in3_124;
assign w1099 = ~in2_125 & in3_125;
assign w1100 = in2_127 & ~in3_127;
assign w1101 = ~in2_126 & in3_126;
assign w1102 = ~w1099 & ~w1100;
assign w1103 = ~w1101 & w1102;
assign w1104 = w1102 & w4949;
assign w1105 = ~in2_88 & in3_88;
assign w1106 = ~w1070 & ~w1105;
assign w1107 = w1069 & w1106;
assign w1108 = w1077 & ~w1107;
assign w1109 = ~in2_92 & in3_92;
assign w1110 = w1020 & w4950;
assign w1111 = w1033 & w1110;
assign w1112 = ~w1108 & w1111;
assign w1113 = w1058 & ~w1112;
assign w1114 = ~in2_100 & in3_100;
assign w1115 = w1041 & w4951;
assign w1116 = ~w1043 & w4952;
assign w1117 = ~in2_104 & in3_104;
assign w1118 = ~w943 & ~w1117;
assign w1119 = w940 & w1118;
assign w1120 = w936 & w1119;
assign w1121 = ~w1116 & w1120;
assign w1122 = w992 & w1121;
assign w1123 = ~w1113 & w1122;
assign w1124 = (w1104 & w1123) | (w1104 & w3691) | (w1123 & w3691);
assign w1125 = (w1124 & ~w1096) | (w1124 & w4953) | (~w1096 & w4953);
assign w1126 = in2_123 & ~in3_123;
assign w1127 = in2_119 & ~in3_119;
assign w1128 = in2_118 & ~in3_118;
assign w1129 = in2_117 & ~in3_117;
assign w1130 = in2_116 & ~in3_116;
assign w1131 = ~w1129 & ~w1130;
assign w1132 = w987 & ~w1131;
assign w1133 = in2_120 & ~in3_120;
assign w1134 = ~w1127 & ~w1133;
assign w1135 = w1134 & w7148;
assign w1136 = w984 & ~w1135;
assign w1137 = in2_122 & ~in3_122;
assign w1138 = in2_121 & ~in3_121;
assign w1139 = ~w1137 & ~w1138;
assign w1140 = w981 & ~w1139;
assign w1141 = ~w1126 & ~w1140;
assign w1142 = (w1104 & w1136) | (w1104 & w4954) | (w1136 & w4954);
assign w1143 = ~in2_127 & in3_127;
assign w1144 = in2_125 & ~in3_125;
assign w1145 = in2_124 & ~in3_124;
assign w1146 = ~w1144 & ~w1145;
assign w1147 = w1103 & ~w1146;
assign w1148 = in2_126 & ~in3_126;
assign w1149 = ~w1100 & w1148;
assign w1150 = ~w1143 & ~w1149;
assign w1151 = ~w1147 & w1150;
assign w1152 = ~w1142 & w1151;
assign w1153 = ~w1142 & w4955;
assign w1154 = (w1096 & w5449) | (w1096 & w5450) | (w5449 & w5450);
assign w1155 = (in2_0 & w1142) | (in2_0 & w4956) | (w1142 & w4956);
assign w1156 = (w1096 & w6866) | (w1096 & w6867) | (w6866 & w6867);
assign w1157 = ~w1154 & w1156;
assign w1158 = ~w578 & w1157;
assign w1159 = ~w1142 & w4957;
assign w1160 = (w1096 & w5451) | (w1096 & w5452) | (w5451 & w5452);
assign w1161 = (in2_1 & w1142) | (in2_1 & w4958) | (w1142 & w4958);
assign w1162 = (w1096 & w6868) | (w1096 & w6869) | (w6868 & w6869);
assign w1163 = ~w1160 & w1162;
assign w1164 = ~w563 & w4959;
assign w1165 = (w517 & w5453) | (w517 & w5454) | (w5453 & w5454);
assign w1166 = (in0_1 & w563) | (in0_1 & w4960) | (w563 & w4960);
assign w1167 = (w517 & w6870) | (w517 & w6871) | (w6870 & w6871);
assign w1168 = ~w1165 & w1167;
assign w1169 = w1163 & ~w1168;
assign w1170 = ~w1158 & ~w1169;
assign w1171 = ~w1163 & w1168;
assign w1172 = ~w563 & w4961;
assign w1173 = (w517 & w5455) | (w517 & w5456) | (w5455 & w5456);
assign w1174 = (in0_2 & w563) | (in0_2 & w4962) | (w563 & w4962);
assign w1175 = (w517 & w6872) | (w517 & w6873) | (w6872 & w6873);
assign w1176 = ~w1173 & w1175;
assign w1177 = ~w1142 & w4963;
assign w1178 = (w1096 & w5457) | (w1096 & w5458) | (w5457 & w5458);
assign w1179 = (in2_2 & w1142) | (in2_2 & w4964) | (w1142 & w4964);
assign w1180 = (w1096 & w6874) | (w1096 & w6875) | (w6874 & w6875);
assign w1181 = ~w1178 & w1180;
assign w1182 = w1176 & ~w1181;
assign w1183 = ~w1171 & ~w1182;
assign w1184 = ~w1170 & w1183;
assign w1185 = (w517 & w5551) | (w517 & w5552) | (w5551 & w5552);
assign w1186 = (~w518 & w4244) | (~w518 & w4245) | (w4244 & w4245);
assign w1187 = (w518 & w4246) | (w518 & w4247) | (w4246 & w4247);
assign w1188 = ~w1186 & ~w1187;
assign w1189 = (w1096 & w5553) | (w1096 & w5554) | (w5553 & w5554);
assign w1190 = (~w1097 & w4248) | (~w1097 & w4249) | (w4248 & w4249);
assign w1191 = (w1097 & w4250) | (w1097 & w4251) | (w4250 & w4251);
assign w1192 = ~w1190 & ~w1191;
assign w1193 = ~w1188 & w1192;
assign w1194 = ~w563 & w4965;
assign w1195 = (w517 & w5459) | (w517 & w5460) | (w5459 & w5460);
assign w1196 = (in0_4 & w563) | (in0_4 & w4966) | (w563 & w4966);
assign w1197 = (w517 & w6876) | (w517 & w6877) | (w6876 & w6877);
assign w1198 = ~w1195 & w1197;
assign w1199 = ~w1142 & w4967;
assign w1200 = (w1096 & w5461) | (w1096 & w5462) | (w5461 & w5462);
assign w1201 = (in2_4 & w1142) | (in2_4 & w4968) | (w1142 & w4968);
assign w1202 = (w1096 & w6878) | (w1096 & w6879) | (w6878 & w6879);
assign w1203 = ~w1200 & w1202;
assign w1204 = ~w1198 & w1203;
assign w1205 = ~w1176 & w1181;
assign w1206 = ~w1204 & ~w1205;
assign w1207 = ~w1193 & w1206;
assign w1208 = ~w1184 & w1207;
assign w1209 = (~w518 & w4256) | (~w518 & w4257) | (w4256 & w4257);
assign w1210 = (w518 & w4258) | (w518 & w4259) | (w4258 & w4259);
assign w1211 = ~w1209 & ~w1210;
assign w1212 = (~w1097 & w4260) | (~w1097 & w4261) | (w4260 & w4261);
assign w1213 = (w1097 & w4262) | (w1097 & w4263) | (w4262 & w4263);
assign w1214 = ~w1212 & ~w1213;
assign w1215 = w1211 & ~w1214;
assign w1216 = ~w563 & w4969;
assign w1217 = (w517 & w5463) | (w517 & w5464) | (w5463 & w5464);
assign w1218 = (in0_6 & w563) | (in0_6 & w4970) | (w563 & w4970);
assign w1219 = (w517 & w6880) | (w517 & w6881) | (w6880 & w6881);
assign w1220 = ~w1217 & w1219;
assign w1221 = ~w1142 & w4971;
assign w1222 = (w1096 & w5465) | (w1096 & w5466) | (w5465 & w5466);
assign w1223 = (in2_6 & w1142) | (in2_6 & w4972) | (w1142 & w4972);
assign w1224 = (w1096 & w6882) | (w1096 & w6883) | (w6882 & w6883);
assign w1225 = ~w1222 & w1224;
assign w1226 = w1220 & ~w1225;
assign w1227 = w1198 & ~w1203;
assign w1228 = w1188 & ~w1192;
assign w1229 = ~w1204 & w1228;
assign w1230 = ~w1226 & ~w1227;
assign w1231 = ~w1215 & w1230;
assign w1232 = ~w1229 & w1231;
assign w1233 = ~w1208 & w1232;
assign w1234 = ~w563 & w4973;
assign w1235 = (w517 & w5467) | (w517 & w5468) | (w5467 & w5468);
assign w1236 = (in0_11 & w563) | (in0_11 & w4974) | (w563 & w4974);
assign w1237 = (w517 & w6884) | (w517 & w6885) | (w6884 & w6885);
assign w1238 = ~w1235 & w1237;
assign w1239 = ~w1142 & w4975;
assign w1240 = (w1096 & w5469) | (w1096 & w5470) | (w5469 & w5470);
assign w1241 = (in2_11 & w1142) | (in2_11 & w4976) | (w1142 & w4976);
assign w1242 = (w1096 & w6886) | (w1096 & w6887) | (w6886 & w6887);
assign w1243 = ~w1240 & w1242;
assign w1244 = w1238 & ~w1243;
assign w1245 = ~w563 & w4977;
assign w1246 = (w517 & w5471) | (w517 & w5472) | (w5471 & w5472);
assign w1247 = (in0_12 & w563) | (in0_12 & w4978) | (w563 & w4978);
assign w1248 = (w517 & w6888) | (w517 & w6889) | (w6888 & w6889);
assign w1249 = ~w1246 & w1248;
assign w1250 = ~w1142 & w4979;
assign w1251 = (w1096 & w5473) | (w1096 & w5474) | (w5473 & w5474);
assign w1252 = (in2_12 & w1142) | (in2_12 & w4980) | (w1142 & w4980);
assign w1253 = (w1096 & w6890) | (w1096 & w6891) | (w6890 & w6891);
assign w1254 = ~w1251 & w1253;
assign w1255 = w1249 & ~w1254;
assign w1256 = ~w1244 & ~w1255;
assign w1257 = ~w1238 & w1243;
assign w1258 = ~w563 & w4981;
assign w1259 = (w517 & w5475) | (w517 & w5476) | (w5475 & w5476);
assign w1260 = (in0_10 & w563) | (in0_10 & w4982) | (w563 & w4982);
assign w1261 = (w517 & w6892) | (w517 & w6893) | (w6892 & w6893);
assign w1262 = ~w1259 & w1261;
assign w1263 = ~w1142 & w4983;
assign w1264 = (w1096 & w5477) | (w1096 & w5478) | (w5477 & w5478);
assign w1265 = (in2_10 & w1142) | (in2_10 & w4984) | (w1142 & w4984);
assign w1266 = (w1096 & w6894) | (w1096 & w6895) | (w6894 & w6895);
assign w1267 = ~w1264 & w1266;
assign w1268 = ~w1262 & w1267;
assign w1269 = ~w1257 & ~w1268;
assign w1270 = w1256 & ~w1269;
assign w1271 = ~w563 & w4985;
assign w1272 = (w517 & w5479) | (w517 & w5480) | (w5479 & w5480);
assign w1273 = (in0_14 & w563) | (in0_14 & w4986) | (w563 & w4986);
assign w1274 = (w517 & w6896) | (w517 & w6897) | (w6896 & w6897);
assign w1275 = ~w1272 & w1274;
assign w1276 = ~w1142 & w4987;
assign w1277 = (w1096 & w5481) | (w1096 & w5482) | (w5481 & w5482);
assign w1278 = (in2_14 & w1142) | (in2_14 & w4988) | (w1142 & w4988);
assign w1279 = (w1096 & w6898) | (w1096 & w6899) | (w6898 & w6899);
assign w1280 = ~w1277 & w1279;
assign w1281 = ~w1275 & w1280;
assign w1282 = ~w563 & w4989;
assign w1283 = (w517 & w5483) | (w517 & w5484) | (w5483 & w5484);
assign w1284 = (in0_15 & w563) | (in0_15 & w4990) | (w563 & w4990);
assign w1285 = (w517 & w6900) | (w517 & w6901) | (w6900 & w6901);
assign w1286 = ~w1283 & w1285;
assign w1287 = ~w1142 & w4991;
assign w1288 = (w1096 & w5485) | (w1096 & w5486) | (w5485 & w5486);
assign w1289 = (in2_15 & w1142) | (in2_15 & w4992) | (w1142 & w4992);
assign w1290 = (w1096 & w6902) | (w1096 & w6903) | (w6902 & w6903);
assign w1291 = ~w1288 & w1290;
assign w1292 = ~w1286 & w1291;
assign w1293 = ~w1281 & ~w1292;
assign w1294 = ~w1249 & w1254;
assign w1295 = ~w563 & w4993;
assign w1296 = (w517 & w5487) | (w517 & w5488) | (w5487 & w5488);
assign w1297 = (in0_13 & w563) | (in0_13 & w4994) | (w563 & w4994);
assign w1298 = (w517 & w6904) | (w517 & w6905) | (w6904 & w6905);
assign w1299 = ~w1296 & w1298;
assign w1300 = ~w1142 & w4995;
assign w1301 = (w1096 & w5489) | (w1096 & w5490) | (w5489 & w5490);
assign w1302 = (in2_13 & w1142) | (in2_13 & w4996) | (w1142 & w4996);
assign w1303 = (w1096 & w6906) | (w1096 & w6907) | (w6906 & w6907);
assign w1304 = ~w1301 & w1303;
assign w1305 = ~w1299 & w1304;
assign w1306 = ~w1294 & ~w1305;
assign w1307 = w1293 & w1306;
assign w1308 = ~w1270 & w1307;
assign w1309 = ~w1142 & w4997;
assign w1310 = (w1096 & w5491) | (w1096 & w5492) | (w5491 & w5492);
assign w1311 = (in2_8 & w1142) | (in2_8 & w4998) | (w1142 & w4998);
assign w1312 = (w1096 & w6908) | (w1096 & w6909) | (w6908 & w6909);
assign w1313 = ~w1310 & w1312;
assign w1314 = ~w563 & w4999;
assign w1315 = (w517 & w5493) | (w517 & w5494) | (w5493 & w5494);
assign w1316 = (in0_8 & w563) | (in0_8 & w5000) | (w563 & w5000);
assign w1317 = (w517 & w6910) | (w517 & w6911) | (w6910 & w6911);
assign w1318 = ~w1315 & w1317;
assign w1319 = w1313 & ~w1318;
assign w1320 = ~w563 & w5001;
assign w1321 = (w517 & w5495) | (w517 & w5496) | (w5495 & w5496);
assign w1322 = (in0_9 & w563) | (in0_9 & w5002) | (w563 & w5002);
assign w1323 = (w517 & w6912) | (w517 & w6913) | (w6912 & w6913);
assign w1324 = ~w1321 & w1323;
assign w1325 = ~w1142 & w5003;
assign w1326 = (w1096 & w5497) | (w1096 & w5498) | (w5497 & w5498);
assign w1327 = (in2_9 & w1142) | (in2_9 & w5004) | (w1142 & w5004);
assign w1328 = (w1096 & w6914) | (w1096 & w6915) | (w6914 & w6915);
assign w1329 = ~w1326 & w1328;
assign w1330 = ~w1324 & w1329;
assign w1331 = ~w1319 & ~w1330;
assign w1332 = ~w1220 & w1225;
assign w1333 = ~w563 & w5005;
assign w1334 = (w517 & w5499) | (w517 & w5500) | (w5499 & w5500);
assign w1335 = (in0_7 & w563) | (in0_7 & w5006) | (w563 & w5006);
assign w1336 = (w517 & w6916) | (w517 & w6917) | (w6916 & w6917);
assign w1337 = ~w1334 & w1336;
assign w1338 = ~w1142 & w5007;
assign w1339 = (w1096 & w5501) | (w1096 & w5502) | (w5501 & w5502);
assign w1340 = (in2_7 & w1142) | (in2_7 & w5008) | (w1142 & w5008);
assign w1341 = (w1096 & w6918) | (w1096 & w6919) | (w6918 & w6919);
assign w1342 = ~w1339 & w1341;
assign w1343 = ~w1337 & w1342;
assign w1344 = ~w1211 & w1214;
assign w1345 = ~w1226 & w1344;
assign w1346 = ~w1332 & ~w1343;
assign w1347 = w1331 & w1346;
assign w1348 = ~w1345 & w1347;
assign w1349 = w1308 & w1348;
assign w1350 = ~w1233 & w1349;
assign w1351 = ~w1313 & w1318;
assign w1352 = w1337 & ~w1342;
assign w1353 = ~w1351 & ~w1352;
assign w1354 = w1331 & ~w1353;
assign w1355 = w1262 & ~w1267;
assign w1356 = w1324 & ~w1329;
assign w1357 = ~w1355 & ~w1356;
assign w1358 = w1256 & w1357;
assign w1359 = ~w1354 & w1358;
assign w1360 = w1308 & ~w1359;
assign w1361 = ~w563 & w5009;
assign w1362 = (w517 & w5503) | (w517 & w5504) | (w5503 & w5504);
assign w1363 = (in0_19 & w563) | (in0_19 & w5010) | (w563 & w5010);
assign w1364 = (w517 & w6920) | (w517 & w6921) | (w6920 & w6921);
assign w1365 = ~w1362 & w1364;
assign w1366 = ~w1142 & w5011;
assign w1367 = (w1096 & w5505) | (w1096 & w5506) | (w5505 & w5506);
assign w1368 = (in2_19 & w1142) | (in2_19 & w5012) | (w1142 & w5012);
assign w1369 = (w1096 & w6922) | (w1096 & w6923) | (w6922 & w6923);
assign w1370 = ~w1367 & w1369;
assign w1371 = w1365 & ~w1370;
assign w1372 = ~w563 & w5013;
assign w1373 = (w517 & w5507) | (w517 & w5508) | (w5507 & w5508);
assign w1374 = (in0_18 & w563) | (in0_18 & w5014) | (w563 & w5014);
assign w1375 = (w517 & w6924) | (w517 & w6925) | (w6924 & w6925);
assign w1376 = ~w1373 & w1375;
assign w1377 = ~w1142 & w5015;
assign w1378 = (w1096 & w5509) | (w1096 & w5510) | (w5509 & w5510);
assign w1379 = (in2_18 & w1142) | (in2_18 & w5016) | (w1142 & w5016);
assign w1380 = (w1096 & w6926) | (w1096 & w6927) | (w6926 & w6927);
assign w1381 = ~w1378 & w1380;
assign w1382 = w1376 & ~w1381;
assign w1383 = ~w1371 & ~w1382;
assign w1384 = ~w1365 & w1370;
assign w1385 = ~w563 & w5017;
assign w1386 = (w517 & w5511) | (w517 & w5512) | (w5511 & w5512);
assign w1387 = (in0_20 & w563) | (in0_20 & w5018) | (w563 & w5018);
assign w1388 = (w517 & w6928) | (w517 & w6929) | (w6928 & w6929);
assign w1389 = ~w1386 & w1388;
assign w1390 = ~w1142 & w5019;
assign w1391 = (w1096 & w5513) | (w1096 & w5514) | (w5513 & w5514);
assign w1392 = (in2_20 & w1142) | (in2_20 & w5020) | (w1142 & w5020);
assign w1393 = (w1096 & w6930) | (w1096 & w6931) | (w6930 & w6931);
assign w1394 = ~w1391 & w1393;
assign w1395 = ~w1389 & w1394;
assign w1396 = ~w1384 & ~w1395;
assign w1397 = ~w1383 & w1396;
assign w1398 = (~w518 & w4316) | (~w518 & w4317) | (w4316 & w4317);
assign w1399 = (w518 & w4318) | (w518 & w4319) | (w4318 & w4319);
assign w1400 = ~w1398 & ~w1399;
assign w1401 = (~w1097 & w4320) | (~w1097 & w4321) | (w4320 & w4321);
assign w1402 = (w1097 & w4322) | (w1097 & w4323) | (w4322 & w4323);
assign w1403 = ~w1401 & ~w1402;
assign w1404 = w1400 & ~w1403;
assign w1405 = ~w563 & w5021;
assign w1406 = (w517 & w5515) | (w517 & w5516) | (w5515 & w5516);
assign w1407 = (in0_22 & w563) | (in0_22 & w5022) | (w563 & w5022);
assign w1408 = (w517 & w6932) | (w517 & w6933) | (w6932 & w6933);
assign w1409 = ~w1406 & w1408;
assign w1410 = ~w1142 & w5023;
assign w1411 = (w1096 & w5517) | (w1096 & w5518) | (w5517 & w5518);
assign w1412 = (in2_22 & w1142) | (in2_22 & w5024) | (w1142 & w5024);
assign w1413 = (w1096 & w6934) | (w1096 & w6935) | (w6934 & w6935);
assign w1414 = ~w1411 & w1413;
assign w1415 = w1409 & ~w1414;
assign w1416 = w1389 & ~w1394;
assign w1417 = ~w1415 & ~w1416;
assign w1418 = ~w1404 & w1417;
assign w1419 = ~w1397 & w1418;
assign w1420 = w1275 & ~w1280;
assign w1421 = w1299 & ~w1304;
assign w1422 = ~w1420 & ~w1421;
assign w1423 = w1293 & ~w1422;
assign w1424 = (~w518 & w4328) | (~w518 & w4329) | (w4328 & w4329);
assign w1425 = (w518 & w4330) | (w518 & w4331) | (w4330 & w4331);
assign w1426 = ~w1424 & ~w1425;
assign w1427 = (~w1097 & w4332) | (~w1097 & w4333) | (w4332 & w4333);
assign w1428 = (w1097 & w4334) | (w1097 & w4335) | (w4334 & w4335);
assign w1429 = ~w1427 & ~w1428;
assign w1430 = w1426 & ~w1429;
assign w1431 = ~w1142 & w5025;
assign w1432 = (w1096 & w5519) | (w1096 & w5520) | (w5519 & w5520);
assign w1433 = (in2_17 & w1142) | (in2_17 & w5026) | (w1142 & w5026);
assign w1434 = (w1096 & w6936) | (w1096 & w6937) | (w6936 & w6937);
assign w1435 = ~w1432 & w1434;
assign w1436 = ~w563 & w5027;
assign w1437 = (w517 & w5521) | (w517 & w5522) | (w5521 & w5522);
assign w1438 = (in0_17 & w563) | (in0_17 & w5028) | (w563 & w5028);
assign w1439 = (w517 & w6938) | (w517 & w6939) | (w6938 & w6939);
assign w1440 = ~w1437 & w1439;
assign w1441 = ~w1435 & w1440;
assign w1442 = w1286 & ~w1291;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = ~w1430 & w1443;
assign w1445 = ~w1423 & w1444;
assign w1446 = w1419 & w1445;
assign w1447 = ~w1360 & w1446;
assign w1448 = ~w1350 & w1447;
assign w1449 = w1435 & ~w1440;
assign w1450 = ~w1376 & w1381;
assign w1451 = ~w1426 & w1429;
assign w1452 = ~w1441 & w1451;
assign w1453 = ~w1449 & ~w1450;
assign w1454 = w1396 & w1453;
assign w1455 = ~w1452 & w1454;
assign w1456 = w1419 & ~w1455;
assign w1457 = (~w518 & w4340) | (~w518 & w4341) | (w4340 & w4341);
assign w1458 = (w518 & w4342) | (w518 & w4343) | (w4342 & w4343);
assign w1459 = ~w1457 & ~w1458;
assign w1460 = (~w1097 & w4344) | (~w1097 & w4345) | (w4344 & w4345);
assign w1461 = (w1097 & w4346) | (w1097 & w4347) | (w4346 & w4347);
assign w1462 = ~w1460 & ~w1461;
assign w1463 = w1459 & ~w1462;
assign w1464 = (~w518 & w4348) | (~w518 & w4349) | (w4348 & w4349);
assign w1465 = (w518 & w4350) | (w518 & w4351) | (w4350 & w4351);
assign w1466 = ~w1464 & ~w1465;
assign w1467 = (~w1097 & w4352) | (~w1097 & w4353) | (w4352 & w4353);
assign w1468 = (w1097 & w4354) | (w1097 & w4355) | (w4354 & w4355);
assign w1469 = ~w1467 & ~w1468;
assign w1470 = w1466 & ~w1469;
assign w1471 = ~w1463 & ~w1470;
assign w1472 = ~w1459 & w1462;
assign w1473 = (~w518 & w4356) | (~w518 & w4357) | (w4356 & w4357);
assign w1474 = (w518 & w4358) | (w518 & w4359) | (w4358 & w4359);
assign w1475 = ~w1473 & ~w1474;
assign w1476 = (~w1097 & w4360) | (~w1097 & w4361) | (w4360 & w4361);
assign w1477 = (w1097 & w4362) | (w1097 & w4363) | (w4362 & w4363);
assign w1478 = ~w1476 & ~w1477;
assign w1479 = ~w1475 & w1478;
assign w1480 = ~w1472 & ~w1479;
assign w1481 = w1471 & ~w1480;
assign w1482 = (~w518 & w4364) | (~w518 & w4365) | (w4364 & w4365);
assign w1483 = (w518 & w4366) | (w518 & w4367) | (w4366 & w4367);
assign w1484 = ~w1482 & ~w1483;
assign w1485 = (~w1097 & w4368) | (~w1097 & w4369) | (w4368 & w4369);
assign w1486 = (w1097 & w4370) | (w1097 & w4371) | (w4370 & w4371);
assign w1487 = ~w1485 & ~w1486;
assign w1488 = ~w1484 & w1487;
assign w1489 = (~w518 & w4372) | (~w518 & w4373) | (w4372 & w4373);
assign w1490 = (w518 & w4374) | (w518 & w4375) | (w4374 & w4375);
assign w1491 = ~w1489 & ~w1490;
assign w1492 = (~w1097 & w4376) | (~w1097 & w4377) | (w4376 & w4377);
assign w1493 = (w1097 & w4378) | (w1097 & w4379) | (w4378 & w4379);
assign w1494 = ~w1492 & ~w1493;
assign w1495 = ~w1491 & w1494;
assign w1496 = ~w1488 & ~w1495;
assign w1497 = ~w1466 & w1469;
assign w1498 = (~w518 & w4380) | (~w518 & w4381) | (w4380 & w4381);
assign w1499 = (w518 & w4382) | (w518 & w4383) | (w4382 & w4383);
assign w1500 = ~w1498 & ~w1499;
assign w1501 = (~w1097 & w4384) | (~w1097 & w4385) | (w4384 & w4385);
assign w1502 = (w1097 & w4386) | (w1097 & w4387) | (w4386 & w4387);
assign w1503 = ~w1501 & ~w1502;
assign w1504 = ~w1500 & w1503;
assign w1505 = ~w1497 & ~w1504;
assign w1506 = w1496 & w1505;
assign w1507 = ~w1481 & w1506;
assign w1508 = (~w518 & w4388) | (~w518 & w4389) | (w4388 & w4389);
assign w1509 = (w518 & w4390) | (w518 & w4391) | (w4390 & w4391);
assign w1510 = ~w1508 & ~w1509;
assign w1511 = (~w1097 & w4392) | (~w1097 & w4393) | (w4392 & w4393);
assign w1512 = (w1097 & w4394) | (w1097 & w4395) | (w4394 & w4395);
assign w1513 = ~w1511 & ~w1512;
assign w1514 = ~w1510 & w1513;
assign w1515 = (~w518 & w4396) | (~w518 & w4397) | (w4396 & w4397);
assign w1516 = (w518 & w4398) | (w518 & w4399) | (w4398 & w4399);
assign w1517 = ~w1515 & ~w1516;
assign w1518 = (~w1097 & w4400) | (~w1097 & w4401) | (w4400 & w4401);
assign w1519 = (w1097 & w4402) | (w1097 & w4403) | (w4402 & w4403);
assign w1520 = ~w1518 & ~w1519;
assign w1521 = ~w1517 & w1520;
assign w1522 = ~w1514 & ~w1521;
assign w1523 = ~w1409 & w1414;
assign w1524 = (~w518 & w4404) | (~w518 & w4405) | (w4404 & w4405);
assign w1525 = (w518 & w4406) | (w518 & w4407) | (w4406 & w4407);
assign w1526 = ~w1524 & ~w1525;
assign w1527 = (~w1097 & w4408) | (~w1097 & w4409) | (w4408 & w4409);
assign w1528 = (w1097 & w4410) | (w1097 & w4411) | (w4410 & w4411);
assign w1529 = ~w1527 & ~w1528;
assign w1530 = ~w1526 & w1529;
assign w1531 = ~w1400 & w1403;
assign w1532 = ~w1415 & w1531;
assign w1533 = ~w1523 & ~w1530;
assign w1534 = w1522 & w1533;
assign w1535 = ~w1532 & w1534;
assign w1536 = ~w1456 & w4412;
assign w1537 = ~w1448 & w1536;
assign w1538 = w1510 & ~w1513;
assign w1539 = w1526 & ~w1529;
assign w1540 = ~w1538 & ~w1539;
assign w1541 = w1522 & ~w1540;
assign w1542 = w1475 & ~w1478;
assign w1543 = w1517 & ~w1520;
assign w1544 = ~w1542 & ~w1543;
assign w1545 = w1471 & w1544;
assign w1546 = ~w1541 & w1545;
assign w1547 = w1507 & ~w1546;
assign w1548 = (~w518 & w4413) | (~w518 & w4414) | (w4413 & w4414);
assign w1549 = (w518 & w4415) | (w518 & w4416) | (w4415 & w4416);
assign w1550 = ~w1548 & ~w1549;
assign w1551 = (~w1097 & w4417) | (~w1097 & w4418) | (w4417 & w4418);
assign w1552 = (w1097 & w4419) | (w1097 & w4420) | (w4419 & w4420);
assign w1553 = ~w1551 & ~w1552;
assign w1554 = w1550 & ~w1553;
assign w1555 = (~w518 & w4421) | (~w518 & w4422) | (w4421 & w4422);
assign w1556 = (w518 & w4423) | (w518 & w4424) | (w4423 & w4424);
assign w1557 = ~w1555 & ~w1556;
assign w1558 = (~w1097 & w4425) | (~w1097 & w4426) | (w4425 & w4426);
assign w1559 = (w1097 & w4427) | (w1097 & w4428) | (w4427 & w4428);
assign w1560 = ~w1558 & ~w1559;
assign w1561 = w1557 & ~w1560;
assign w1562 = (~w518 & w4429) | (~w518 & w4430) | (w4429 & w4430);
assign w1563 = (w518 & w4431) | (w518 & w4432) | (w4431 & w4432);
assign w1564 = ~w1562 & ~w1563;
assign w1565 = (~w1097 & w4433) | (~w1097 & w4434) | (w4433 & w4434);
assign w1566 = (w1097 & w4435) | (w1097 & w4436) | (w4435 & w4436);
assign w1567 = ~w1565 & ~w1566;
assign w1568 = w1564 & ~w1567;
assign w1569 = (~w518 & w4437) | (~w518 & w4438) | (w4437 & w4438);
assign w1570 = (w518 & w4439) | (w518 & w4440) | (w4439 & w4440);
assign w1571 = ~w1569 & ~w1570;
assign w1572 = (~w1097 & w4441) | (~w1097 & w4442) | (w4441 & w4442);
assign w1573 = (w1097 & w4443) | (w1097 & w4444) | (w4443 & w4444);
assign w1574 = ~w1572 & ~w1573;
assign w1575 = w1571 & ~w1574;
assign w1576 = (~w1097 & w4445) | (~w1097 & w4446) | (w4445 & w4446);
assign w1577 = (w1097 & w4447) | (w1097 & w4448) | (w4447 & w4448);
assign w1578 = ~w1576 & ~w1577;
assign w1579 = (~w518 & w4449) | (~w518 & w4450) | (w4449 & w4450);
assign w1580 = (w518 & w4451) | (w518 & w4452) | (w4451 & w4452);
assign w1581 = ~w1579 & ~w1580;
assign w1582 = ~w1578 & w1581;
assign w1583 = (~w518 & w4453) | (~w518 & w4454) | (w4453 & w4454);
assign w1584 = (w518 & w4455) | (w518 & w4456) | (w4455 & w4456);
assign w1585 = ~w1583 & ~w1584;
assign w1586 = (~w1097 & w4457) | (~w1097 & w4458) | (w4457 & w4458);
assign w1587 = (w1097 & w4459) | (w1097 & w4460) | (w4459 & w4460);
assign w1588 = ~w1586 & ~w1587;
assign w1589 = w1585 & ~w1588;
assign w1590 = ~w1582 & ~w1589;
assign w1591 = (~w518 & w4461) | (~w518 & w4462) | (w4461 & w4462);
assign w1592 = (w518 & w4463) | (w518 & w4464) | (w4463 & w4464);
assign w1593 = ~w1591 & ~w1592;
assign w1594 = (~w1097 & w4465) | (~w1097 & w4466) | (w4465 & w4466);
assign w1595 = (w1097 & w4467) | (w1097 & w4468) | (w4467 & w4468);
assign w1596 = ~w1594 & ~w1595;
assign w1597 = w1593 & ~w1596;
assign w1598 = (~w518 & w4469) | (~w518 & w4470) | (w4469 & w4470);
assign w1599 = (w518 & w4471) | (w518 & w4472) | (w4471 & w4472);
assign w1600 = ~w1598 & ~w1599;
assign w1601 = (~w1097 & w4473) | (~w1097 & w4474) | (w4473 & w4474);
assign w1602 = (w1097 & w4475) | (w1097 & w4476) | (w4475 & w4476);
assign w1603 = ~w1601 & ~w1602;
assign w1604 = w1600 & ~w1603;
assign w1605 = (~w518 & w4477) | (~w518 & w4478) | (w4477 & w4478);
assign w1606 = (w518 & w4479) | (w518 & w4480) | (w4479 & w4480);
assign w1607 = ~w1605 & ~w1606;
assign w1608 = (~w1097 & w4481) | (~w1097 & w4482) | (w4481 & w4482);
assign w1609 = (w1097 & w4483) | (w1097 & w4484) | (w4483 & w4484);
assign w1610 = ~w1608 & ~w1609;
assign w1611 = w1607 & ~w1610;
assign w1612 = ~w1597 & ~w1604;
assign w1613 = ~w1611 & w1612;
assign w1614 = ~w1554 & ~w1561;
assign w1615 = ~w1568 & ~w1575;
assign w1616 = w1614 & w1615;
assign w1617 = w1590 & w1616;
assign w1618 = w1613 & w1617;
assign w1619 = ~w1142 & w5029;
assign w1620 = (w1096 & w5523) | (w1096 & w5524) | (w5523 & w5524);
assign w1621 = (in2_32 & w1142) | (in2_32 & w5030) | (w1142 & w5030);
assign w1622 = (w1096 & w6940) | (w1096 & w6941) | (w6940 & w6941);
assign w1623 = ~w1620 & w1622;
assign w1624 = ~w563 & w5031;
assign w1625 = (w517 & w5525) | (w517 & w5526) | (w5525 & w5526);
assign w1626 = (in0_32 & w563) | (in0_32 & w5032) | (w563 & w5032);
assign w1627 = (w517 & w6942) | (w517 & w6943) | (w6942 & w6943);
assign w1628 = ~w1625 & w1627;
assign w1629 = ~w1623 & w1628;
assign w1630 = ~w563 & w5033;
assign w1631 = (w517 & w5527) | (w517 & w5528) | (w5527 & w5528);
assign w1632 = (in0_33 & w563) | (in0_33 & w5034) | (w563 & w5034);
assign w1633 = (w517 & w6944) | (w517 & w6945) | (w6944 & w6945);
assign w1634 = ~w1631 & w1633;
assign w1635 = ~w1142 & w5035;
assign w1636 = (w1096 & w5529) | (w1096 & w5530) | (w5529 & w5530);
assign w1637 = (in2_33 & w1142) | (in2_33 & w5036) | (w1142 & w5036);
assign w1638 = (w1096 & w6946) | (w1096 & w6947) | (w6946 & w6947);
assign w1639 = ~w1636 & w1638;
assign w1640 = w1634 & ~w1639;
assign w1641 = ~w1142 & w5037;
assign w1642 = (w1096 & w5531) | (w1096 & w5532) | (w5531 & w5532);
assign w1643 = (in2_34 & w1142) | (in2_34 & w5038) | (w1142 & w5038);
assign w1644 = (w1096 & w6948) | (w1096 & w6949) | (w6948 & w6949);
assign w1645 = ~w1642 & w1644;
assign w1646 = ~w563 & w5039;
assign w1647 = (w517 & w5533) | (w517 & w5534) | (w5533 & w5534);
assign w1648 = (in0_34 & w563) | (in0_34 & w5040) | (w563 & w5040);
assign w1649 = (w517 & w6950) | (w517 & w6951) | (w6950 & w6951);
assign w1650 = ~w1647 & w1649;
assign w1651 = ~w1645 & w1650;
assign w1652 = ~w1640 & ~w1651;
assign w1653 = w1491 & ~w1494;
assign w1654 = w1484 & ~w1487;
assign w1655 = w1500 & ~w1503;
assign w1656 = ~w1654 & ~w1655;
assign w1657 = w1496 & ~w1656;
assign w1658 = (~w518 & w4497) | (~w518 & w4498) | (w4497 & w4498);
assign w1659 = (w518 & w4499) | (w518 & w4500) | (w4499 & w4500);
assign w1660 = ~w1658 & ~w1659;
assign w1661 = (~w1097 & w4501) | (~w1097 & w4502) | (w4501 & w4502);
assign w1662 = (w1097 & w4503) | (w1097 & w4504) | (w4503 & w4504);
assign w1663 = ~w1661 & ~w1662;
assign w1664 = w1660 & ~w1663;
assign w1665 = (~w1097 & w4505) | (~w1097 & w4506) | (w4505 & w4506);
assign w1666 = (w1097 & w4507) | (w1097 & w4508) | (w4507 & w4508);
assign w1667 = ~w1665 & ~w1666;
assign w1668 = (~w518 & w4509) | (~w518 & w4510) | (w4509 & w4510);
assign w1669 = (w518 & w4511) | (w518 & w4512) | (w4511 & w4512);
assign w1670 = ~w1668 & ~w1669;
assign w1671 = ~w1667 & w1670;
assign w1672 = ~w1664 & ~w1671;
assign w1673 = (~w518 & w4513) | (~w518 & w4514) | (w4513 & w4514);
assign w1674 = (w518 & w4515) | (w518 & w4516) | (w4515 & w4516);
assign w1675 = ~w1673 & ~w1674;
assign w1676 = (~w1097 & w4517) | (~w1097 & w4518) | (w4517 & w4518);
assign w1677 = (w1097 & w4519) | (w1097 & w4520) | (w4519 & w4520);
assign w1678 = ~w1676 & ~w1677;
assign w1679 = w1675 & ~w1678;
assign w1680 = (~w518 & w4521) | (~w518 & w4522) | (w4521 & w4522);
assign w1681 = (w518 & w4523) | (w518 & w4524) | (w4523 & w4524);
assign w1682 = ~w1680 & ~w1681;
assign w1683 = (~w1097 & w4525) | (~w1097 & w4526) | (w4525 & w4526);
assign w1684 = (w1097 & w4527) | (w1097 & w4528) | (w4527 & w4528);
assign w1685 = ~w1683 & ~w1684;
assign w1686 = w1682 & ~w1685;
assign w1687 = ~w1679 & ~w1686;
assign w1688 = w1672 & w1687;
assign w1689 = w1652 & w4529;
assign w1690 = ~w1657 & w1689;
assign w1691 = w1688 & w1690;
assign w1692 = ~w1547 & w1691;
assign w1693 = w1618 & w1692;
assign w1694 = ~w1537 & w1693;
assign w1695 = ~w563 & w5041;
assign w1696 = (w517 & w5555) | (w517 & w5556) | (w5555 & w5556);
assign w1697 = (in0_55 & w563) | (in0_55 & w5042) | (w563 & w5042);
assign w1698 = (w517 & w7079) | (w517 & w7080) | (w7079 & w7080);
assign w1699 = ~w1696 & w1698;
assign w1700 = ~w1142 & w5043;
assign w1701 = (w1096 & w5557) | (w1096 & w5558) | (w5557 & w5558);
assign w1702 = (in2_55 & w1142) | (in2_55 & w5044) | (w1142 & w5044);
assign w1703 = (w1096 & w7081) | (w1096 & w7082) | (w7081 & w7082);
assign w1704 = ~w1701 & w1703;
assign w1705 = ~w1699 & w1704;
assign w1706 = w1699 & ~w1704;
assign w1707 = ~w1142 & w5045;
assign w1708 = (w1096 & w5559) | (w1096 & w5560) | (w5559 & w5560);
assign w1709 = (in2_54 & w1142) | (in2_54 & w5046) | (w1142 & w5046);
assign w1710 = (w1096 & w7083) | (w1096 & w7084) | (w7083 & w7084);
assign w1711 = ~w1708 & w1710;
assign w1712 = ~w563 & w5047;
assign w1713 = (w517 & w5561) | (w517 & w5562) | (w5561 & w5562);
assign w1714 = (in0_54 & w563) | (in0_54 & w5048) | (w563 & w5048);
assign w1715 = (w517 & w7085) | (w517 & w7086) | (w7085 & w7086);
assign w1716 = ~w1713 & w1715;
assign w1717 = ~w1711 & w1716;
assign w1718 = ~w1706 & ~w1717;
assign w1719 = ~w1705 & ~w1718;
assign w1720 = ~w563 & w5049;
assign w1721 = (w517 & w5563) | (w517 & w5564) | (w5563 & w5564);
assign w1722 = (in0_52 & w563) | (in0_52 & w5050) | (w563 & w5050);
assign w1723 = (w517 & w7087) | (w517 & w7088) | (w7087 & w7088);
assign w1724 = ~w1721 & w1723;
assign w1725 = ~w1142 & w5051;
assign w1726 = (w1096 & w5565) | (w1096 & w5566) | (w5565 & w5566);
assign w1727 = (in2_52 & w1142) | (in2_52 & w5052) | (w1142 & w5052);
assign w1728 = (w1096 & w7089) | (w1096 & w7090) | (w7089 & w7090);
assign w1729 = ~w1726 & w1728;
assign w1730 = ~w1724 & w1729;
assign w1731 = ~w563 & w5053;
assign w1732 = (w517 & w5567) | (w517 & w5568) | (w5567 & w5568);
assign w1733 = (in0_51 & w563) | (in0_51 & w5054) | (w563 & w5054);
assign w1734 = (w517 & w7091) | (w517 & w7092) | (w7091 & w7092);
assign w1735 = ~w1732 & w1734;
assign w1736 = ~w1142 & w5055;
assign w1737 = (w1096 & w5569) | (w1096 & w5570) | (w5569 & w5570);
assign w1738 = (in2_51 & w1142) | (in2_51 & w5056) | (w1142 & w5056);
assign w1739 = (w1096 & w7093) | (w1096 & w7094) | (w7093 & w7094);
assign w1740 = ~w1737 & w1739;
assign w1741 = w1735 & ~w1740;
assign w1742 = ~w1730 & w1741;
assign w1743 = w1724 & ~w1729;
assign w1744 = ~w563 & w5057;
assign w1745 = (w517 & w5571) | (w517 & w5572) | (w5571 & w5572);
assign w1746 = (in0_53 & w563) | (in0_53 & w5058) | (w563 & w5058);
assign w1747 = (w517 & w7095) | (w517 & w7096) | (w7095 & w7096);
assign w1748 = ~w1745 & w1747;
assign w1749 = ~w1142 & w5059;
assign w1750 = (w1096 & w5573) | (w1096 & w5574) | (w5573 & w5574);
assign w1751 = (in2_53 & w1142) | (in2_53 & w5060) | (w1142 & w5060);
assign w1752 = (w1096 & w7097) | (w1096 & w7098) | (w7097 & w7098);
assign w1753 = ~w1750 & w1752;
assign w1754 = w1748 & ~w1753;
assign w1755 = ~w1743 & ~w1754;
assign w1756 = ~w1742 & w1755;
assign w1757 = ~w1719 & w1756;
assign w1758 = ~w563 & w5061;
assign w1759 = (w517 & w5575) | (w517 & w5576) | (w5575 & w5576);
assign w1760 = (in0_49 & w563) | (in0_49 & w5062) | (w563 & w5062);
assign w1761 = (w517 & w7099) | (w517 & w7100) | (w7099 & w7100);
assign w1762 = ~w1759 & w1761;
assign w1763 = ~w1142 & w5063;
assign w1764 = (w1096 & w5577) | (w1096 & w5578) | (w5577 & w5578);
assign w1765 = (in2_49 & w1142) | (in2_49 & w5064) | (w1142 & w5064);
assign w1766 = (w1096 & w7101) | (w1096 & w7102) | (w7101 & w7102);
assign w1767 = ~w1764 & w1766;
assign w1768 = ~w1762 & w1767;
assign w1769 = ~w1142 & w5065;
assign w1770 = (w1096 & w5579) | (w1096 & w5580) | (w5579 & w5580);
assign w1771 = (in2_48 & w1142) | (in2_48 & w5066) | (w1142 & w5066);
assign w1772 = (w1096 & w7103) | (w1096 & w7104) | (w7103 & w7104);
assign w1773 = ~w1770 & w1772;
assign w1774 = ~w563 & w5067;
assign w1775 = (w517 & w5581) | (w517 & w5582) | (w5581 & w5582);
assign w1776 = (in0_48 & w563) | (in0_48 & w5068) | (w563 & w5068);
assign w1777 = (w517 & w7105) | (w517 & w7106) | (w7105 & w7106);
assign w1778 = ~w1775 & w1777;
assign w1779 = w1773 & ~w1778;
assign w1780 = ~w1768 & ~w1779;
assign w1781 = w1762 & ~w1767;
assign w1782 = ~w1142 & w5069;
assign w1783 = (w1096 & w5583) | (w1096 & w5584) | (w5583 & w5584);
assign w1784 = (in2_50 & w1142) | (in2_50 & w5070) | (w1142 & w5070);
assign w1785 = (w1096 & w7107) | (w1096 & w7108) | (w7107 & w7108);
assign w1786 = ~w1783 & w1785;
assign w1787 = ~w563 & w5071;
assign w1788 = (w517 & w5585) | (w517 & w5586) | (w5585 & w5586);
assign w1789 = (in0_50 & w563) | (in0_50 & w5072) | (w563 & w5072);
assign w1790 = (w517 & w7109) | (w517 & w7110) | (w7109 & w7110);
assign w1791 = ~w1788 & w1790;
assign w1792 = ~w1786 & w1791;
assign w1793 = ~w1781 & ~w1792;
assign w1794 = ~w1780 & w1793;
assign w1795 = ~w1735 & w1740;
assign w1796 = w1786 & ~w1791;
assign w1797 = ~w1730 & ~w1795;
assign w1798 = ~w1796 & w1797;
assign w1799 = ~w1794 & w1798;
assign w1800 = w1757 & ~w1799;
assign w1801 = w1711 & ~w1716;
assign w1802 = ~w1748 & w1753;
assign w1803 = ~w1705 & ~w1801;
assign w1804 = ~w1802 & w1803;
assign w1805 = ~w1719 & ~w1804;
assign w1806 = ~w1800 & ~w1805;
assign w1807 = w1623 & ~w1628;
assign w1808 = ~w1634 & w1639;
assign w1809 = ~w1807 & ~w1808;
assign w1810 = w1652 & ~w1809;
assign w1811 = ~w1682 & w1685;
assign w1812 = w1645 & ~w1650;
assign w1813 = ~w1811 & ~w1812;
assign w1814 = ~w1810 & w1813;
assign w1815 = w1688 & ~w1814;
assign w1816 = ~w1660 & w1663;
assign w1817 = ~w1675 & w1678;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = w1672 & ~w1818;
assign w1820 = ~w1550 & w1553;
assign w1821 = w1667 & ~w1670;
assign w1822 = ~w1820 & ~w1821;
assign w1823 = ~w1819 & w1822;
assign w1824 = ~w1815 & w1823;
assign w1825 = w1618 & ~w1824;
assign w1826 = ~w1564 & w1567;
assign w1827 = ~w1575 & w1826;
assign w1828 = ~w1607 & w1610;
assign w1829 = ~w1571 & w1574;
assign w1830 = ~w1828 & ~w1829;
assign w1831 = ~w1827 & w1830;
assign w1832 = w1613 & ~w1831;
assign w1833 = ~w1600 & w1603;
assign w1834 = w1578 & ~w1581;
assign w1835 = ~w1585 & w1588;
assign w1836 = ~w1557 & w1560;
assign w1837 = ~w1593 & w1596;
assign w1838 = ~w1604 & w1837;
assign w1839 = ~w1833 & ~w1834;
assign w1840 = ~w1835 & ~w1836;
assign w1841 = w1839 & w1840;
assign w1842 = ~w1838 & w1841;
assign w1843 = ~w1832 & w1842;
assign w1844 = w1561 & ~w1834;
assign w1845 = w1590 & ~w1844;
assign w1846 = ~w1835 & ~w1845;
assign w1847 = ~w1843 & ~w1846;
assign w1848 = ~w563 & w5073;
assign w1849 = (w517 & w5535) | (w517 & w5536) | (w5535 & w5536);
assign w1850 = (in0_57 & w563) | (in0_57 & w5074) | (w563 & w5074);
assign w1851 = (w517 & w6952) | (w517 & w6953) | (w6952 & w6953);
assign w1852 = ~w1849 & w1851;
assign w1853 = ~w1142 & w5075;
assign w1854 = (w1096 & w5537) | (w1096 & w5538) | (w5537 & w5538);
assign w1855 = (in2_57 & w1142) | (in2_57 & w5076) | (w1142 & w5076);
assign w1856 = (w1096 & w6954) | (w1096 & w6955) | (w6954 & w6955);
assign w1857 = ~w1854 & w1856;
assign w1858 = w1852 & ~w1857;
assign w1859 = ~w563 & w5077;
assign w1860 = (w517 & w5539) | (w517 & w5540) | (w5539 & w5540);
assign w1861 = (in0_56 & w563) | (in0_56 & w5078) | (w563 & w5078);
assign w1862 = (w517 & w6956) | (w517 & w6957) | (w6956 & w6957);
assign w1863 = ~w1860 & w1862;
assign w1864 = ~w1142 & w5079;
assign w1865 = (w1096 & w5541) | (w1096 & w5542) | (w5541 & w5542);
assign w1866 = (in2_56 & w1142) | (in2_56 & w5080) | (w1142 & w5080);
assign w1867 = (w1096 & w6958) | (w1096 & w6959) | (w6958 & w6959);
assign w1868 = ~w1865 & w1867;
assign w1869 = ~w1863 & w1868;
assign w1870 = ~w1858 & w1869;
assign w1871 = ~w1852 & w1857;
assign w1872 = ~w563 & w5081;
assign w1873 = (w517 & w5543) | (w517 & w5544) | (w5543 & w5544);
assign w1874 = (in0_58 & w563) | (in0_58 & w5082) | (w563 & w5082);
assign w1875 = (w517 & w6960) | (w517 & w6961) | (w6960 & w6961);
assign w1876 = ~w1873 & w1875;
assign w1877 = ~w1142 & w5083;
assign w1878 = (w1096 & w5545) | (w1096 & w5546) | (w5545 & w5546);
assign w1879 = (in2_58 & w1142) | (in2_58 & w5084) | (w1142 & w5084);
assign w1880 = (w1096 & w6962) | (w1096 & w6963) | (w6962 & w6963);
assign w1881 = ~w1878 & w1880;
assign w1882 = ~w1876 & w1881;
assign w1883 = ~w1871 & ~w1882;
assign w1884 = ~w1870 & w1883;
assign w1885 = w1876 & ~w1881;
assign w1886 = ~w563 & w5085;
assign w1887 = (w517 & w5547) | (w517 & w5548) | (w5547 & w5548);
assign w1888 = (in0_60 & w563) | (in0_60 & w5086) | (w563 & w5086);
assign w1889 = (w517 & w6964) | (w517 & w6965) | (w6964 & w6965);
assign w1890 = ~w1887 & w1889;
assign w1891 = ~w1142 & w5087;
assign w1892 = (w1096 & w5549) | (w1096 & w5550) | (w5549 & w5550);
assign w1893 = (in2_60 & w1142) | (in2_60 & w5088) | (w1142 & w5088);
assign w1894 = (w1096 & w6966) | (w1096 & w6967) | (w6966 & w6967);
assign w1895 = ~w1892 & w1894;
assign w1896 = w1890 & ~w1895;
assign w1897 = ~w563 & w5089;
assign w1898 = (w517 & w6121) | (w517 & w6122) | (w6121 & w6122);
assign w1899 = (in0_59 & w563) | (in0_59 & w5090) | (w563 & w5090);
assign w1900 = (w517 & w6968) | (w517 & w6969) | (w6968 & w6969);
assign w1901 = ~w1898 & w1900;
assign w1902 = ~w1142 & w5091;
assign w1903 = (w1096 & w6123) | (w1096 & w6124) | (w6123 & w6124);
assign w1904 = (in2_59 & w1142) | (in2_59 & w5092) | (w1142 & w5092);
assign w1905 = (w1096 & w6970) | (w1096 & w6971) | (w6970 & w6971);
assign w1906 = ~w1903 & w1905;
assign w1907 = w1901 & ~w1906;
assign w1908 = ~w1885 & ~w1896;
assign w1909 = ~w1907 & w1908;
assign w1910 = ~w1884 & w1909;
assign w1911 = (~w1097 & w4582) | (~w1097 & w4583) | (w4582 & w4583);
assign w1912 = (w1097 & w4584) | (w1097 & w4585) | (w4584 & w4585);
assign w1913 = ~w1911 & ~w1912;
assign w1914 = (~w518 & w4586) | (~w518 & w4587) | (w4586 & w4587);
assign w1915 = (w518 & w4588) | (w518 & w4589) | (w4588 & w4589);
assign w1916 = ~w1914 & ~w1915;
assign w1917 = w1913 & ~w1916;
assign w1918 = (~w518 & w4590) | (~w518 & w4591) | (w4590 & w4591);
assign w1919 = (w518 & w4592) | (w518 & w4593) | (w4592 & w4593);
assign w1920 = ~w1918 & ~w1919;
assign w1921 = (~w1097 & w4594) | (~w1097 & w4595) | (w4594 & w4595);
assign w1922 = (w1097 & w4596) | (w1097 & w4597) | (w4596 & w4597);
assign w1923 = ~w1921 & ~w1922;
assign w1924 = ~w1920 & w1923;
assign w1925 = ~w1917 & ~w1924;
assign w1926 = ~w1901 & w1906;
assign w1927 = ~w1896 & w1926;
assign w1928 = ~w1890 & w1895;
assign w1929 = ~w563 & w5093;
assign w1930 = (w517 & w6125) | (w517 & w6126) | (w6125 & w6126);
assign w1931 = (in0_61 & w563) | (in0_61 & w5094) | (w563 & w5094);
assign w1932 = (w517 & w6972) | (w517 & w6973) | (w6972 & w6973);
assign w1933 = ~w1930 & w1932;
assign w1934 = ~w1142 & w5095;
assign w1935 = (w1096 & w6127) | (w1096 & w6128) | (w6127 & w6128);
assign w1936 = (in2_61 & w1142) | (in2_61 & w5096) | (w1142 & w5096);
assign w1937 = (w1096 & w6974) | (w1096 & w6975) | (w6974 & w6975);
assign w1938 = ~w1935 & w1937;
assign w1939 = ~w1933 & w1938;
assign w1940 = ~w1928 & ~w1939;
assign w1941 = ~w1927 & w1940;
assign w1942 = w1925 & w1941;
assign w1943 = ~w1910 & w1942;
assign w1944 = (~w518 & w4602) | (~w518 & w4603) | (w4602 & w4603);
assign w1945 = (w518 & w4604) | (w518 & w4605) | (w4604 & w4605);
assign w1946 = ~w1944 & ~w1945;
assign w1947 = (~w1097 & w4606) | (~w1097 & w4607) | (w4606 & w4607);
assign w1948 = (w1097 & w4608) | (w1097 & w4609) | (w4608 & w4609);
assign w1949 = ~w1947 & ~w1948;
assign w1950 = w1946 & ~w1949;
assign w1951 = ~w1142 & w5097;
assign w1952 = (w1096 & w6193) | (w1096 & w6194) | (w6193 & w6194);
assign w1953 = (in2_66 & w1142) | (in2_66 & w5098) | (w1142 & w5098);
assign w1954 = (w1096 & w7111) | (w1096 & w7112) | (w7111 & w7112);
assign w1955 = ~w1952 & w1954;
assign w1956 = ~w563 & w5099;
assign w1957 = (w517 & w6195) | (w517 & w6196) | (w6195 & w6196);
assign w1958 = (in0_66 & w563) | (in0_66 & w5100) | (w563 & w5100);
assign w1959 = (w517 & w7113) | (w517 & w7114) | (w7113 & w7114);
assign w1960 = ~w1957 & w1959;
assign w1961 = ~w1955 & w1960;
assign w1962 = ~w1950 & ~w1961;
assign w1963 = w1920 & ~w1923;
assign w1964 = ~w563 & w5101;
assign w1965 = (w517 & w6129) | (w517 & w6130) | (w6129 & w6130);
assign w1966 = (in0_65 & w563) | (in0_65 & w5102) | (w563 & w5102);
assign w1967 = (w517 & w6976) | (w517 & w6977) | (w6976 & w6977);
assign w1968 = ~w1965 & w1967;
assign w1969 = ~w1142 & w5103;
assign w1970 = (w1096 & w6131) | (w1096 & w6132) | (w6131 & w6132);
assign w1971 = (in2_65 & w1142) | (in2_65 & w5104) | (w1142 & w5104);
assign w1972 = (w1096 & w6978) | (w1096 & w6979) | (w6978 & w6979);
assign w1973 = ~w1970 & w1972;
assign w1974 = w1968 & ~w1973;
assign w1975 = ~w1142 & w5105;
assign w1976 = (w1096 & w6133) | (w1096 & w6134) | (w6133 & w6134);
assign w1977 = (in2_64 & w1142) | (in2_64 & w5106) | (w1142 & w5106);
assign w1978 = (w1096 & w6980) | (w1096 & w6981) | (w6980 & w6981);
assign w1979 = ~w1976 & w1978;
assign w1980 = ~w563 & w5107;
assign w1981 = (w517 & w6135) | (w517 & w6136) | (w6135 & w6136);
assign w1982 = (in0_64 & w563) | (in0_64 & w5108) | (w563 & w5108);
assign w1983 = (w517 & w6982) | (w517 & w6983) | (w6982 & w6983);
assign w1984 = ~w1981 & w1983;
assign w1985 = ~w1979 & w1984;
assign w1986 = ~w1974 & ~w1985;
assign w1987 = ~w1963 & w1986;
assign w1988 = w1962 & w1987;
assign w1989 = ~w1913 & w1916;
assign w1990 = w1933 & ~w1938;
assign w1991 = ~w1989 & ~w1990;
assign w1992 = w1925 & ~w1991;
assign w1993 = w1988 & ~w1992;
assign w1994 = ~w1943 & w1993;
assign w1995 = ~w1946 & w1949;
assign w1996 = w1979 & ~w1984;
assign w1997 = ~w1974 & w1996;
assign w1998 = w1955 & ~w1960;
assign w1999 = ~w1968 & w1973;
assign w2000 = ~w1998 & ~w1999;
assign w2001 = ~w1997 & w2000;
assign w2002 = (~w518 & w4622) | (~w518 & w4623) | (w4622 & w4623);
assign w2003 = (w518 & w4624) | (w518 & w4625) | (w4624 & w4625);
assign w2004 = ~w2002 & ~w2003;
assign w2005 = (~w1097 & w4626) | (~w1097 & w4627) | (w4626 & w4627);
assign w2006 = (w1097 & w4628) | (w1097 & w4629) | (w4628 & w4629);
assign w2007 = ~w2005 & ~w2006;
assign w2008 = ~w2004 & w2007;
assign w2009 = ~w563 & w5109;
assign w2010 = (w517 & w6137) | (w517 & w6138) | (w6137 & w6138);
assign w2011 = (in0_69 & w563) | (in0_69 & w5110) | (w563 & w5110);
assign w2012 = (w517 & w6984) | (w517 & w6985) | (w6984 & w6985);
assign w2013 = ~w2010 & w2012;
assign w2014 = ~w1142 & w5111;
assign w2015 = (w1096 & w6139) | (w1096 & w6140) | (w6139 & w6140);
assign w2016 = (in2_69 & w1142) | (in2_69 & w5112) | (w1142 & w5112);
assign w2017 = (w1096 & w6986) | (w1096 & w6987) | (w6986 & w6987);
assign w2018 = ~w2015 & w2017;
assign w2019 = ~w2013 & w2018;
assign w2020 = ~w2008 & ~w2019;
assign w2021 = (~w518 & w4634) | (~w518 & w4635) | (w4634 & w4635);
assign w2022 = (w518 & w4636) | (w518 & w4637) | (w4636 & w4637);
assign w2023 = ~w2021 & ~w2022;
assign w2024 = (~w1097 & w4638) | (~w1097 & w4639) | (w4638 & w4639);
assign w2025 = (w1097 & w4640) | (w1097 & w4641) | (w4640 & w4641);
assign w2026 = ~w2024 & ~w2025;
assign w2027 = w2023 & ~w2026;
assign w2028 = w2013 & ~w2018;
assign w2029 = ~w1142 & w5113;
assign w2030 = (w1096 & w6141) | (w1096 & w6142) | (w6141 & w6142);
assign w2031 = (in2_70 & w1142) | (in2_70 & w5114) | (w1142 & w5114);
assign w2032 = (w1096 & w6988) | (w1096 & w6989) | (w6988 & w6989);
assign w2033 = ~w2030 & w2032;
assign w2034 = ~w563 & w5115;
assign w2035 = (w517 & w6143) | (w517 & w6144) | (w6143 & w6144);
assign w2036 = (in0_70 & w563) | (in0_70 & w5116) | (w563 & w5116);
assign w2037 = (w517 & w6990) | (w517 & w6991) | (w6990 & w6991);
assign w2038 = ~w2035 & w2037;
assign w2039 = ~w2033 & w2038;
assign w2040 = ~w2028 & ~w2039;
assign w2041 = ~w2027 & w2040;
assign w2042 = ~w2020 & w2041;
assign w2043 = ~w2023 & w2026;
assign w2044 = w2033 & ~w2038;
assign w2045 = ~w2027 & w2044;
assign w2046 = ~w2043 & ~w2045;
assign w2047 = ~w2042 & w2046;
assign w2048 = (~w1995 & w2001) | (~w1995 & w4646) | (w2001 & w4646);
assign w2049 = w2047 & w2048;
assign w2050 = ~w1994 & w2049;
assign w2051 = w1806 & ~w1825;
assign w2052 = ~w1847 & w2050;
assign w2053 = w2051 & w2052;
assign w2054 = ~w1694 & w2053;
assign w2055 = ~w1773 & w1778;
assign w2056 = w1793 & ~w2055;
assign w2057 = w1757 & w2056;
assign w2058 = w1863 & ~w1868;
assign w2059 = ~w1858 & ~w2058;
assign w2060 = w1909 & w5117;
assign w2061 = w1988 & w2060;
assign w2062 = (w2061 & ~w1806) | (w2061 & w5118) | (~w1806 & w5118);
assign w2063 = w2050 & ~w2062;
assign w2064 = w2004 & ~w2007;
assign w2065 = w2040 & w5119;
assign w2066 = ~w2042 & w5120;
assign w2067 = (~w518 & w5121) | (~w518 & w5122) | (w5121 & w5122);
assign w2068 = (w518 & w5123) | (w518 & w5124) | (w5123 & w5124);
assign w2069 = ~w2067 & ~w2068;
assign w2070 = (~w518 & w4647) | (~w518 & w4648) | (w4647 & w4648);
assign w2071 = (w518 & w4649) | (w518 & w4650) | (w4649 & w4650);
assign w2072 = ~w2070 & ~w2071;
assign w2073 = (~w1097 & w4651) | (~w1097 & w4652) | (w4651 & w4652);
assign w2074 = (w1097 & w4653) | (w1097 & w4654) | (w4653 & w4654);
assign w2075 = ~w2073 & ~w2074;
assign w2076 = ~w2072 & w2075;
assign w2077 = (~w1097 & w5125) | (~w1097 & w5126) | (w5125 & w5126);
assign w2078 = (w1097 & w5127) | (w1097 & w5128) | (w5127 & w5128);
assign w2079 = ~w2077 & ~w2078;
assign w2080 = w2069 & ~w2079;
assign w2081 = ~w2076 & w2080;
assign w2082 = (~w1097 & w4655) | (~w1097 & w4656) | (w4655 & w4656);
assign w2083 = (w1097 & w4657) | (w1097 & w4658) | (w4657 & w4658);
assign w2084 = ~w2082 & ~w2083;
assign w2085 = (~w518 & w4659) | (~w518 & w4660) | (w4659 & w4660);
assign w2086 = (w518 & w4661) | (w518 & w4662) | (w4661 & w4662);
assign w2087 = ~w2085 & ~w2086;
assign w2088 = ~w2084 & w2087;
assign w2089 = (~w518 & w4663) | (~w518 & w4664) | (w4663 & w4664);
assign w2090 = (w518 & w4665) | (w518 & w4666) | (w4665 & w4666);
assign w2091 = ~w2089 & ~w2090;
assign w2092 = (~w1097 & w4667) | (~w1097 & w4668) | (w4667 & w4668);
assign w2093 = (w1097 & w4669) | (w1097 & w4670) | (w4669 & w4670);
assign w2094 = ~w2092 & ~w2093;
assign w2095 = w2091 & ~w2094;
assign w2096 = (~w518 & w4671) | (~w518 & w4672) | (w4671 & w4672);
assign w2097 = (w518 & w4673) | (w518 & w4674) | (w4673 & w4674);
assign w2098 = ~w2096 & ~w2097;
assign w2099 = (~w1097 & w4675) | (~w1097 & w4676) | (w4675 & w4676);
assign w2100 = (w1097 & w4677) | (w1097 & w4678) | (w4677 & w4678);
assign w2101 = ~w2099 & ~w2100;
assign w2102 = w2098 & ~w2101;
assign w2103 = ~w563 & w5129;
assign w2104 = (w517 & w6145) | (w517 & w6146) | (w6145 & w6146);
assign w2105 = (in0_91 & w563) | (in0_91 & w5130) | (w563 & w5130);
assign w2106 = (w517 & w6992) | (w517 & w6993) | (w6992 & w6993);
assign w2107 = ~w2104 & w2106;
assign w2108 = ~w1142 & w5131;
assign w2109 = (w1096 & w6147) | (w1096 & w6148) | (w6147 & w6148);
assign w2110 = (in2_91 & w1142) | (in2_91 & w5132) | (w1142 & w5132);
assign w2111 = (w1096 & w6994) | (w1096 & w6995) | (w6994 & w6995);
assign w2112 = ~w2109 & w2111;
assign w2113 = w2107 & ~w2112;
assign w2114 = ~w1142 & w5133;
assign w2115 = (w1096 & w6149) | (w1096 & w6150) | (w6149 & w6150);
assign w2116 = (in2_90 & w1142) | (in2_90 & w5134) | (w1142 & w5134);
assign w2117 = (w1096 & w6996) | (w1096 & w6997) | (w6996 & w6997);
assign w2118 = ~w2115 & w2117;
assign w2119 = ~w563 & w5135;
assign w2120 = (w517 & w6151) | (w517 & w6152) | (w6151 & w6152);
assign w2121 = (in0_90 & w563) | (in0_90 & w5136) | (w563 & w5136);
assign w2122 = (w517 & w6998) | (w517 & w6999) | (w6998 & w6999);
assign w2123 = ~w2120 & w2122;
assign w2124 = ~w2118 & w2123;
assign w2125 = ~w2113 & ~w2124;
assign w2126 = ~w2088 & ~w2095;
assign w2127 = ~w2102 & w2125;
assign w2128 = w2126 & w2127;
assign w2129 = w2072 & ~w2075;
assign w2130 = ~w1142 & w5137;
assign w2131 = (w1096 & w6153) | (w1096 & w6154) | (w6153 & w6154);
assign w2132 = (in2_86 & w1142) | (in2_86 & w5138) | (w1142 & w5138);
assign w2133 = (w1096 & w7000) | (w1096 & w7001) | (w7000 & w7001);
assign w2134 = ~w2131 & w2133;
assign w2135 = ~w563 & w5139;
assign w2136 = (w517 & w6155) | (w517 & w6156) | (w6155 & w6156);
assign w2137 = (in0_86 & w563) | (in0_86 & w5140) | (w563 & w5140);
assign w2138 = (w517 & w7002) | (w517 & w7003) | (w7002 & w7003);
assign w2139 = ~w2136 & w2138;
assign w2140 = ~w2134 & w2139;
assign w2141 = ~w563 & w5141;
assign w2142 = (w517 & w6157) | (w517 & w6158) | (w6157 & w6158);
assign w2143 = (in0_85 & w563) | (in0_85 & w5142) | (w563 & w5142);
assign w2144 = (w517 & w7004) | (w517 & w7005) | (w7004 & w7005);
assign w2145 = ~w2142 & w2144;
assign w2146 = ~w1142 & w5143;
assign w2147 = (w1096 & w6159) | (w1096 & w6160) | (w6159 & w6160);
assign w2148 = (in2_85 & w1142) | (in2_85 & w5144) | (w1142 & w5144);
assign w2149 = (w1096 & w7006) | (w1096 & w7007) | (w7006 & w7007);
assign w2150 = ~w2147 & w2149;
assign w2151 = w2145 & ~w2150;
assign w2152 = ~w2140 & ~w2151;
assign w2153 = ~w563 & w5145;
assign w2154 = (w517 & w6161) | (w517 & w6162) | (w6161 & w6162);
assign w2155 = (in0_84 & w563) | (in0_84 & w5146) | (w563 & w5146);
assign w2156 = (w517 & w7008) | (w517 & w7009) | (w7008 & w7009);
assign w2157 = ~w2154 & w2156;
assign w2158 = ~w1142 & w5147;
assign w2159 = (w1096 & w6163) | (w1096 & w6164) | (w6163 & w6164);
assign w2160 = (in2_84 & w1142) | (in2_84 & w5148) | (w1142 & w5148);
assign w2161 = (w1096 & w7010) | (w1096 & w7011) | (w7010 & w7011);
assign w2162 = ~w2159 & w2161;
assign w2163 = w2157 & ~w2162;
assign w2164 = (~w518 & w5149) | (~w518 & w5150) | (w5149 & w5150);
assign w2165 = (w518 & w5151) | (w518 & w5152) | (w5151 & w5152);
assign w2166 = ~w2164 & ~w2165;
assign w2167 = (~w1097 & w5153) | (~w1097 & w5154) | (w5153 & w5154);
assign w2168 = (w1097 & w5155) | (w1097 & w5156) | (w5155 & w5156);
assign w2169 = ~w2167 & ~w2168;
assign w2170 = ~w2166 & w2169;
assign w2171 = ~w2069 & w2079;
assign w2172 = ~w2076 & ~w2170;
assign w2173 = ~w2171 & w2172;
assign w2174 = w2166 & ~w2169;
assign w2175 = (~w518 & w5157) | (~w518 & w5158) | (w5157 & w5158);
assign w2176 = (w518 & w5159) | (w518 & w5160) | (w5159 & w5160);
assign w2177 = ~w2175 & ~w2176;
assign w2178 = ~w2174 & ~w2177;
assign w2179 = (~w1097 & w5161) | (~w1097 & w5162) | (w5161 & w5162);
assign w2180 = (w1097 & w5163) | (w1097 & w5164) | (w5163 & w5164);
assign w2181 = ~w2179 & ~w2180;
assign w2182 = ~w2174 & w2181;
assign w2183 = ~w2178 & ~w2182;
assign w2184 = w2173 & w2183;
assign w2185 = ~w2129 & ~w2163;
assign w2186 = w2152 & w2185;
assign w2187 = ~w2081 & w2186;
assign w2188 = w2128 & w2187;
assign w2189 = ~w2184 & w2188;
assign w2190 = (~w1097 & w4699) | (~w1097 & w4700) | (w4699 & w4700);
assign w2191 = (w1097 & w4701) | (w1097 & w4702) | (w4701 & w4702);
assign w2192 = ~w2190 & ~w2191;
assign w2193 = (~w518 & w4703) | (~w518 & w4704) | (w4703 & w4704);
assign w2194 = (w518 & w4705) | (w518 & w4706) | (w4705 & w4706);
assign w2195 = ~w2193 & ~w2194;
assign w2196 = ~w2192 & w2195;
assign w2197 = ~w563 & w5165;
assign w2198 = (w517 & w6197) | (w517 & w6198) | (w6197 & w6198);
assign w2199 = (in0_77 & w563) | (in0_77 & w5166) | (w563 & w5166);
assign w2200 = (w517 & w7115) | (w517 & w7116) | (w7115 & w7116);
assign w2201 = ~w2198 & w2200;
assign w2202 = ~w1142 & w5167;
assign w2203 = (w1096 & w6199) | (w1096 & w6200) | (w6199 & w6200);
assign w2204 = (in2_77 & w1142) | (in2_77 & w5168) | (w1142 & w5168);
assign w2205 = (w1096 & w7117) | (w1096 & w7118) | (w7117 & w7118);
assign w2206 = ~w2203 & w2205;
assign w2207 = w2201 & ~w2206;
assign w2208 = ~w2196 & ~w2207;
assign w2209 = ~w1142 & w5169;
assign w2210 = (w1096 & w6201) | (w1096 & w6202) | (w6201 & w6202);
assign w2211 = (in2_72 & w1142) | (in2_72 & w5170) | (w1142 & w5170);
assign w2212 = (w1096 & w7119) | (w1096 & w7120) | (w7119 & w7120);
assign w2213 = ~w2210 & w2212;
assign w2214 = ~w563 & w5171;
assign w2215 = (w517 & w6203) | (w517 & w6204) | (w6203 & w6204);
assign w2216 = (in0_72 & w563) | (in0_72 & w5172) | (w563 & w5172);
assign w2217 = (w517 & w7121) | (w517 & w7122) | (w7121 & w7122);
assign w2218 = ~w2215 & w2217;
assign w2219 = ~w2213 & w2218;
assign w2220 = ~w563 & w5173;
assign w2221 = (w517 & w6205) | (w517 & w6206) | (w6205 & w6206);
assign w2222 = (in0_73 & w563) | (in0_73 & w5174) | (w563 & w5174);
assign w2223 = (w517 & w7123) | (w517 & w7124) | (w7123 & w7124);
assign w2224 = ~w2221 & w2223;
assign w2225 = ~w1142 & w5175;
assign w2226 = (w1096 & w6207) | (w1096 & w6208) | (w6207 & w6208);
assign w2227 = (in2_73 & w1142) | (in2_73 & w5176) | (w1142 & w5176);
assign w2228 = (w1096 & w7125) | (w1096 & w7126) | (w7125 & w7126);
assign w2229 = ~w2226 & w2228;
assign w2230 = w2224 & ~w2229;
assign w2231 = (~w518 & w4719) | (~w518 & w4720) | (w4719 & w4720);
assign w2232 = (w518 & w4721) | (w518 & w4722) | (w4721 & w4722);
assign w2233 = ~w2231 & ~w2232;
assign w2234 = (~w1097 & w4723) | (~w1097 & w4724) | (w4723 & w4724);
assign w2235 = (w1097 & w4725) | (w1097 & w4726) | (w4725 & w4726);
assign w2236 = ~w2234 & ~w2235;
assign w2237 = w2233 & ~w2236;
assign w2238 = ~w563 & w5177;
assign w2239 = (w517 & w6209) | (w517 & w6210) | (w6209 & w6210);
assign w2240 = (in0_75 & w563) | (in0_75 & w5178) | (w563 & w5178);
assign w2241 = (w517 & w7127) | (w517 & w7128) | (w7127 & w7128);
assign w2242 = ~w2239 & w2241;
assign w2243 = ~w1142 & w5179;
assign w2244 = (w1096 & w6211) | (w1096 & w6212) | (w6211 & w6212);
assign w2245 = (in2_75 & w1142) | (in2_75 & w5180) | (w1142 & w5180);
assign w2246 = (w1096 & w7129) | (w1096 & w7130) | (w7129 & w7130);
assign w2247 = ~w2244 & w2246;
assign w2248 = w2242 & ~w2247;
assign w2249 = ~w563 & w5181;
assign w2250 = (w517 & w6213) | (w517 & w6214) | (w6213 & w6214);
assign w2251 = (in0_76 & w563) | (in0_76 & w5182) | (w563 & w5182);
assign w2252 = (w517 & w7131) | (w517 & w7132) | (w7131 & w7132);
assign w2253 = ~w2250 & w2252;
assign w2254 = ~w1142 & w5183;
assign w2255 = (w1096 & w6215) | (w1096 & w6216) | (w6215 & w6216);
assign w2256 = (in2_76 & w1142) | (in2_76 & w5184) | (w1142 & w5184);
assign w2257 = (w1096 & w7133) | (w1096 & w7134) | (w7133 & w7134);
assign w2258 = ~w2255 & w2257;
assign w2259 = w2253 & ~w2258;
assign w2260 = ~w1142 & w5185;
assign w2261 = (w1096 & w6217) | (w1096 & w6218) | (w6217 & w6218);
assign w2262 = (in2_74 & w1142) | (in2_74 & w5186) | (w1142 & w5186);
assign w2263 = (w1096 & w7135) | (w1096 & w7136) | (w7135 & w7136);
assign w2264 = ~w2261 & w2263;
assign w2265 = ~w563 & w5187;
assign w2266 = (w517 & w6219) | (w517 & w6220) | (w6219 & w6220);
assign w2267 = (in0_74 & w563) | (in0_74 & w5188) | (w563 & w5188);
assign w2268 = (w517 & w7137) | (w517 & w7138) | (w7137 & w7138);
assign w2269 = ~w2266 & w2268;
assign w2270 = ~w2264 & w2269;
assign w2271 = ~w2248 & ~w2259;
assign w2272 = ~w2270 & w2271;
assign w2273 = ~w2219 & ~w2230;
assign w2274 = ~w2237 & w2273;
assign w2275 = w2208 & w2274;
assign w2276 = w2272 & w2275;
assign w2277 = ~w2066 & w2276;
assign w2278 = w2189 & w2277;
assign w2279 = ~w2063 & w2278;
assign w2280 = ~w2054 & w2279;
assign w2281 = (~w518 & w4739) | (~w518 & w4740) | (w4739 & w4740);
assign w2282 = (w518 & w4741) | (w518 & w4742) | (w4741 & w4742);
assign w2283 = ~w2281 & ~w2282;
assign w2284 = (~w1097 & w4743) | (~w1097 & w4744) | (w4743 & w4744);
assign w2285 = (w1097 & w4745) | (w1097 & w4746) | (w4745 & w4746);
assign w2286 = ~w2284 & ~w2285;
assign w2287 = w2283 & ~w2286;
assign w2288 = ~w1142 & w5189;
assign w2289 = (w1096 & w6221) | (w1096 & w6222) | (w6221 & w6222);
assign w2290 = (in2_118 & w1142) | (in2_118 & w5190) | (w1142 & w5190);
assign w2291 = (w1096 & w7139) | (w1096 & w7140) | (w7139 & w7140);
assign w2292 = ~w2289 & w2291;
assign w2293 = ~w563 & w5191;
assign w2294 = (w517 & w6223) | (w517 & w6224) | (w6223 & w6224);
assign w2295 = (in0_118 & w563) | (in0_118 & w5192) | (w563 & w5192);
assign w2296 = (w517 & w7141) | (w517 & w7142) | (w7141 & w7142);
assign w2297 = ~w2294 & w2296;
assign w2298 = ~w2292 & w2297;
assign w2299 = ~w563 & w5193;
assign w2300 = (w517 & w6225) | (w517 & w6226) | (w6225 & w6226);
assign w2301 = (in0_117 & w563) | (in0_117 & w5194) | (w563 & w5194);
assign w2302 = (w517 & w7143) | (w517 & w7144) | (w7143 & w7144);
assign w2303 = ~w2300 & w2302;
assign w2304 = ~w1142 & w5195;
assign w2305 = (w1096 & w6227) | (w1096 & w6228) | (w6227 & w6228);
assign w2306 = (in2_117 & w1142) | (in2_117 & w5196) | (w1142 & w5196);
assign w2307 = (w1096 & w7145) | (w1096 & w7146) | (w7145 & w7146);
assign w2308 = ~w2305 & w2307;
assign w2309 = w2303 & ~w2308;
assign w2310 = ~w2298 & ~w2309;
assign w2311 = ~w2287 & w2310;
assign w2312 = (~w518 & w4755) | (~w518 & w4756) | (w4755 & w4756);
assign w2313 = (w518 & w4757) | (w518 & w4758) | (w4757 & w4758);
assign w2314 = ~w2312 & ~w2313;
assign w2315 = (~w1097 & w4759) | (~w1097 & w4760) | (w4759 & w4760);
assign w2316 = (w1097 & w4761) | (w1097 & w4762) | (w4761 & w4762);
assign w2317 = ~w2315 & ~w2316;
assign w2318 = w2314 & ~w2317;
assign w2319 = w2310 & w5197;
assign w2320 = ~w2303 & w2308;
assign w2321 = ~w2314 & w2317;
assign w2322 = ~w2320 & ~w2321;
assign w2323 = w2311 & ~w2322;
assign w2324 = ~w2283 & w2286;
assign w2325 = w2292 & ~w2297;
assign w2326 = ~w2287 & w2325;
assign w2327 = ~w2324 & ~w2326;
assign w2328 = ~w2323 & w5198;
assign w2329 = (~w518 & w4763) | (~w518 & w4764) | (w4763 & w4764);
assign w2330 = (w518 & w4765) | (w518 & w4766) | (w4765 & w4766);
assign w2331 = ~w2329 & ~w2330;
assign w2332 = (~w1097 & w4767) | (~w1097 & w4768) | (w4767 & w4768);
assign w2333 = (w1097 & w4769) | (w1097 & w4770) | (w4769 & w4770);
assign w2334 = ~w2332 & ~w2333;
assign w2335 = w2331 & ~w2334;
assign w2336 = (~w518 & w4771) | (~w518 & w4772) | (w4771 & w4772);
assign w2337 = (w518 & w4773) | (w518 & w4774) | (w4773 & w4774);
assign w2338 = ~w2336 & ~w2337;
assign w2339 = (~w1097 & w4775) | (~w1097 & w4776) | (w4775 & w4776);
assign w2340 = (w1097 & w4777) | (w1097 & w4778) | (w4777 & w4778);
assign w2341 = ~w2339 & ~w2340;
assign w2342 = w2338 & ~w2341;
assign w2343 = ~w2335 & ~w2342;
assign w2344 = (~w518 & w4779) | (~w518 & w4780) | (w4779 & w4780);
assign w2345 = (w518 & w4781) | (w518 & w4782) | (w4781 & w4782);
assign w2346 = ~w2344 & ~w2345;
assign w2347 = (~w1097 & w4783) | (~w1097 & w4784) | (w4783 & w4784);
assign w2348 = (w1097 & w4785) | (w1097 & w4786) | (w4785 & w4786);
assign w2349 = ~w2347 & ~w2348;
assign w2350 = w2346 & ~w2349;
assign w2351 = w2343 & ~w2350;
assign w2352 = (~w518 & w5199) | (~w518 & w5200) | (w5199 & w5200);
assign w2353 = (w518 & w5201) | (w518 & w5202) | (w5201 & w5202);
assign w2354 = ~w2352 & ~w2353;
assign w2355 = (~w1097 & w5203) | (~w1097 & w5204) | (w5203 & w5204);
assign w2356 = (w1097 & w5205) | (w1097 & w5206) | (w5205 & w5206);
assign w2357 = ~w2355 & ~w2356;
assign w2358 = w2354 & ~w2357;
assign w2359 = (~w1097 & w5207) | (~w1097 & w5208) | (w5207 & w5208);
assign w2360 = (w1097 & w5209) | (w1097 & w5210) | (w5209 & w5210);
assign w2361 = ~w2359 & ~w2360;
assign w2362 = (~w518 & w5211) | (~w518 & w5212) | (w5211 & w5212);
assign w2363 = (w518 & w5213) | (w518 & w5214) | (w5213 & w5214);
assign w2364 = ~w2362 & ~w2363;
assign w2365 = ~w2361 & w2364;
assign w2366 = ~w2358 & ~w2365;
assign w2367 = w2351 & w2366;
assign w2368 = (~w518 & w5215) | (~w518 & w5216) | (w5215 & w5216);
assign w2369 = (w518 & w5217) | (w518 & w5218) | (w5217 & w5218);
assign w2370 = ~w2368 & ~w2369;
assign w2371 = (~w1097 & w5219) | (~w1097 & w5220) | (w5219 & w5220);
assign w2372 = (w1097 & w5221) | (w1097 & w5222) | (w5221 & w5222);
assign w2373 = ~w2371 & ~w2372;
assign w2374 = w2370 & ~w2373;
assign w2375 = (~w1097 & w5223) | (~w1097 & w5224) | (w5223 & w5224);
assign w2376 = (w1097 & w5225) | (w1097 & w5226) | (w5225 & w5226);
assign w2377 = ~w2375 & ~w2376;
assign w2378 = (~w518 & w5227) | (~w518 & w5228) | (w5227 & w5228);
assign w2379 = (w518 & w5229) | (w518 & w5230) | (w5229 & w5230);
assign w2380 = ~w2378 & ~w2379;
assign w2381 = ~w2377 & w2380;
assign w2382 = ~w2374 & ~w2381;
assign w2383 = w2351 & w5231;
assign w2384 = ~w2328 & w2383;
assign w2385 = ~w563 & w5232;
assign w2386 = (w517 & w6165) | (w517 & w6166) | (w6165 & w6166);
assign w2387 = (in0_115 & w563) | (in0_115 & w5233) | (w563 & w5233);
assign w2388 = (w517 & w7012) | (w517 & w7013) | (w7012 & w7013);
assign w2389 = ~w2386 & w2388;
assign w2390 = ~w1142 & w5234;
assign w2391 = (w1096 & w6167) | (w1096 & w6168) | (w6167 & w6168);
assign w2392 = (in2_115 & w1142) | (in2_115 & w5235) | (w1142 & w5235);
assign w2393 = (w1096 & w7014) | (w1096 & w7015) | (w7014 & w7015);
assign w2394 = ~w2391 & w2393;
assign w2395 = ~w2389 & w2394;
assign w2396 = w2389 & ~w2394;
assign w2397 = ~w1142 & w5236;
assign w2398 = (w1096 & w6169) | (w1096 & w6170) | (w6169 & w6170);
assign w2399 = (in2_114 & w1142) | (in2_114 & w5237) | (w1142 & w5237);
assign w2400 = (w1096 & w7016) | (w1096 & w7017) | (w7016 & w7017);
assign w2401 = ~w2398 & w2400;
assign w2402 = ~w563 & w5238;
assign w2403 = (w517 & w6171) | (w517 & w6172) | (w6171 & w6172);
assign w2404 = (in0_114 & w563) | (in0_114 & w5239) | (w563 & w5239);
assign w2405 = (w517 & w7018) | (w517 & w7019) | (w7018 & w7019);
assign w2406 = ~w2403 & w2405;
assign w2407 = ~w2401 & w2406;
assign w2408 = ~w2396 & ~w2407;
assign w2409 = (~w518 & w4795) | (~w518 & w4796) | (w4795 & w4796);
assign w2410 = (w518 & w4797) | (w518 & w4798) | (w4797 & w4798);
assign w2411 = ~w2409 & ~w2410;
assign w2412 = (~w1097 & w4799) | (~w1097 & w4800) | (w4799 & w4800);
assign w2413 = (w1097 & w4801) | (w1097 & w4802) | (w4801 & w4802);
assign w2414 = ~w2412 & ~w2413;
assign w2415 = w2411 & ~w2414;
assign w2416 = (~w1097 & w4803) | (~w1097 & w4804) | (w4803 & w4804);
assign w2417 = (w1097 & w4805) | (w1097 & w4806) | (w4805 & w4806);
assign w2418 = ~w2416 & ~w2417;
assign w2419 = (~w518 & w4807) | (~w518 & w4808) | (w4807 & w4808);
assign w2420 = (w518 & w4809) | (w518 & w4810) | (w4809 & w4810);
assign w2421 = ~w2419 & ~w2420;
assign w2422 = w2418 & ~w2421;
assign w2423 = ~w2415 & w2422;
assign w2424 = w2401 & ~w2406;
assign w2425 = ~w2411 & w2414;
assign w2426 = ~w2424 & ~w2425;
assign w2427 = ~w2423 & w2426;
assign w2428 = w2408 & ~w2427;
assign w2429 = ~w563 & w5240;
assign w2430 = (w517 & w6173) | (w517 & w6174) | (w6173 & w6174);
assign w2431 = (in0_109 & w563) | (in0_109 & w5241) | (w563 & w5241);
assign w2432 = (w517 & w7020) | (w517 & w7021) | (w7020 & w7021);
assign w2433 = ~w2430 & w2432;
assign w2434 = ~w1142 & w5242;
assign w2435 = (w1096 & w6175) | (w1096 & w6176) | (w6175 & w6176);
assign w2436 = (in2_109 & w1142) | (in2_109 & w5243) | (w1142 & w5243);
assign w2437 = (w1096 & w7022) | (w1096 & w7023) | (w7022 & w7023);
assign w2438 = ~w2435 & w2437;
assign w2439 = w2433 & ~w2438;
assign w2440 = ~w1142 & w5244;
assign w2441 = (w1096 & w6177) | (w1096 & w6178) | (w6177 & w6178);
assign w2442 = (in2_110 & w1142) | (in2_110 & w5245) | (w1142 & w5245);
assign w2443 = (w1096 & w7024) | (w1096 & w7025) | (w7024 & w7025);
assign w2444 = ~w2441 & w2443;
assign w2445 = ~w563 & w5246;
assign w2446 = (w517 & w6179) | (w517 & w6180) | (w6179 & w6180);
assign w2447 = (in0_110 & w563) | (in0_110 & w5247) | (w563 & w5247);
assign w2448 = (w517 & w7026) | (w517 & w7027) | (w7026 & w7027);
assign w2449 = ~w2446 & w2448;
assign w2450 = ~w2444 & w2449;
assign w2451 = ~w2439 & ~w2450;
assign w2452 = ~w2433 & w2438;
assign w2453 = ~w563 & w5248;
assign w2454 = (w517 & w6181) | (w517 & w6182) | (w6181 & w6182);
assign w2455 = (in0_108 & w563) | (in0_108 & w5249) | (w563 & w5249);
assign w2456 = (w517 & w7028) | (w517 & w7029) | (w7028 & w7029);
assign w2457 = ~w2454 & w2456;
assign w2458 = ~w1142 & w5250;
assign w2459 = (w1096 & w6183) | (w1096 & w6184) | (w6183 & w6184);
assign w2460 = (in2_108 & w1142) | (in2_108 & w5251) | (w1142 & w5251);
assign w2461 = (w1096 & w7030) | (w1096 & w7031) | (w7030 & w7031);
assign w2462 = ~w2459 & w2461;
assign w2463 = ~w2457 & w2462;
assign w2464 = ~w2452 & ~w2463;
assign w2465 = w2451 & ~w2464;
assign w2466 = w2444 & ~w2449;
assign w2467 = (~w518 & w4823) | (~w518 & w4824) | (w4823 & w4824);
assign w2468 = (w518 & w4825) | (w518 & w4826) | (w4825 & w4826);
assign w2469 = ~w2467 & ~w2468;
assign w2470 = (~w1097 & w4827) | (~w1097 & w4828) | (w4827 & w4828);
assign w2471 = (w1097 & w4829) | (w1097 & w4830) | (w4829 & w4830);
assign w2472 = ~w2470 & ~w2471;
assign w2473 = ~w2469 & w2472;
assign w2474 = ~w2466 & ~w2473;
assign w2475 = ~w2465 & w2474;
assign w2476 = ~w2418 & w2421;
assign w2477 = w2469 & ~w2472;
assign w2478 = w2408 & ~w2415;
assign w2479 = ~w2476 & ~w2477;
assign w2480 = w2478 & w2479;
assign w2481 = ~w2475 & w2480;
assign w2482 = ~w2323 & w4831;
assign w2483 = ~w2428 & ~w2481;
assign w2484 = w2482 & w2483;
assign w2485 = w2384 & ~w2484;
assign w2486 = w2361 & ~w2364;
assign w2487 = ~w2370 & w2373;
assign w2488 = w2377 & ~w2380;
assign w2489 = ~w2374 & w2488;
assign w2490 = ~w2486 & ~w2487;
assign w2491 = ~w2489 & w2490;
assign w2492 = w2367 & ~w2491;
assign w2493 = ~w2354 & w2357;
assign w2494 = w2343 & w5252;
assign w2495 = ~w2338 & w2341;
assign w2496 = ~w2346 & w2349;
assign w2497 = ~w2495 & ~w2496;
assign w2498 = w2343 & ~w2497;
assign w2499 = (in2_127 & w1125) | (in2_127 & w5253) | (w1125 & w5253);
assign w2500 = ~in1_127 & ~w563;
assign w2501 = (in0_127 & w546) | (in0_127 & w5254) | (w546 & w5254);
assign w2502 = w2499 & ~w2501;
assign w2503 = ~w2498 & ~w2502;
assign w2504 = ~w2494 & w2503;
assign w2505 = ~w2492 & w2504;
assign w2506 = ~w2331 & w2334;
assign w2507 = w2505 & ~w2506;
assign w2508 = ~w2485 & w2507;
assign w2509 = w2213 & ~w2218;
assign w2510 = ~w2230 & w2509;
assign w2511 = w2264 & ~w2269;
assign w2512 = ~w2224 & w2229;
assign w2513 = ~w2511 & ~w2512;
assign w2514 = ~w2510 & w2513;
assign w2515 = w2272 & ~w2514;
assign w2516 = w2192 & ~w2195;
assign w2517 = ~w2233 & w2236;
assign w2518 = ~w2516 & ~w2517;
assign w2519 = ~w2242 & w2247;
assign w2520 = ~w2259 & w2519;
assign w2521 = ~w2253 & w2258;
assign w2522 = ~w2201 & w2206;
assign w2523 = ~w2521 & ~w2522;
assign w2524 = ~w2520 & w2523;
assign w2525 = w2518 & w2524;
assign w2526 = ~w2515 & w2525;
assign w2527 = ~w2208 & w2518;
assign w2528 = ~w2237 & ~w2527;
assign w2529 = ~w2174 & w5255;
assign w2530 = w2173 & ~w2529;
assign w2531 = (w2530 & w2526) | (w2530 & w5256) | (w2526 & w5256);
assign w2532 = w2189 & ~w2531;
assign w2533 = (~w518 & w4832) | (~w518 & w4833) | (w4832 & w4833);
assign w2534 = (w518 & w4834) | (w518 & w4835) | (w4834 & w4835);
assign w2535 = ~w2533 & ~w2534;
assign w2536 = (~w1097 & w4836) | (~w1097 & w4837) | (w4836 & w4837);
assign w2537 = (w1097 & w4838) | (w1097 & w4839) | (w4838 & w4839);
assign w2538 = ~w2536 & ~w2537;
assign w2539 = w2535 & ~w2538;
assign w2540 = ~w1142 & w5257;
assign w2541 = (w1096 & w6185) | (w1096 & w6186) | (w6185 & w6186);
assign w2542 = (in2_102 & w1142) | (in2_102 & w5258) | (w1142 & w5258);
assign w2543 = (w1096 & w7032) | (w1096 & w7033) | (w7032 & w7033);
assign w2544 = ~w2541 & w2543;
assign w2545 = ~w563 & w5259;
assign w2546 = (w517 & w6187) | (w517 & w6188) | (w6187 & w6188);
assign w2547 = (in0_102 & w563) | (in0_102 & w5260) | (w563 & w5260);
assign w2548 = (w517 & w7034) | (w517 & w7035) | (w7034 & w7035);
assign w2549 = ~w2546 & w2548;
assign w2550 = ~w2544 & w2549;
assign w2551 = ~w563 & w5261;
assign w2552 = (w517 & w6189) | (w517 & w6190) | (w6189 & w6190);
assign w2553 = (in0_101 & w563) | (in0_101 & w5262) | (w563 & w5262);
assign w2554 = (w517 & w7036) | (w517 & w7037) | (w7036 & w7037);
assign w2555 = ~w2552 & w2554;
assign w2556 = ~w1142 & w5263;
assign w2557 = (w1096 & w6191) | (w1096 & w6192) | (w6191 & w6192);
assign w2558 = (in2_101 & w1142) | (in2_101 & w5264) | (w1142 & w5264);
assign w2559 = (w1096 & w7038) | (w1096 & w7039) | (w7038 & w7039);
assign w2560 = ~w2557 & w2559;
assign w2561 = w2555 & ~w2560;
assign w2562 = ~w2550 & ~w2561;
assign w2563 = ~w2539 & w2562;
assign w2564 = (~w518 & w4848) | (~w518 & w4849) | (w4848 & w4849);
assign w2565 = (w518 & w4850) | (w518 & w4851) | (w4850 & w4851);
assign w2566 = ~w2564 & ~w2565;
assign w2567 = (~w1097 & w4852) | (~w1097 & w4853) | (w4852 & w4853);
assign w2568 = (w1097 & w4854) | (w1097 & w4855) | (w4854 & w4855);
assign w2569 = ~w2567 & ~w2568;
assign w2570 = w2566 & ~w2569;
assign w2571 = w2562 & w5265;
assign w2572 = (~w518 & w4856) | (~w518 & w4857) | (w4856 & w4857);
assign w2573 = (w518 & w4858) | (w518 & w4859) | (w4858 & w4859);
assign w2574 = ~w2572 & ~w2573;
assign w2575 = (~w1097 & w4860) | (~w1097 & w4861) | (w4860 & w4861);
assign w2576 = (w1097 & w4862) | (w1097 & w4863) | (w4862 & w4863);
assign w2577 = ~w2575 & ~w2576;
assign w2578 = ~w2574 & w2577;
assign w2579 = w2574 & ~w2577;
assign w2580 = ~w1142 & w5266;
assign w2581 = (w1096 & w6229) | (w1096 & w6230) | (w6229 & w6230);
assign w2582 = (in2_98 & w1142) | (in2_98 & w5267) | (w1142 & w5267);
assign w2583 = (w1096 & w7040) | (w1096 & w7041) | (w7040 & w7041);
assign w2584 = ~w2581 & w2583;
assign w2585 = ~w563 & w5268;
assign w2586 = (w517 & w6231) | (w517 & w6232) | (w6231 & w6232);
assign w2587 = (in0_98 & w563) | (in0_98 & w5269) | (w563 & w5269);
assign w2588 = (w517 & w7042) | (w517 & w7043) | (w7042 & w7043);
assign w2589 = ~w2586 & w2588;
assign w2590 = ~w2584 & w2589;
assign w2591 = ~w2579 & ~w2590;
assign w2592 = ~w563 & w5270;
assign w2593 = (w517 & w6233) | (w517 & w6234) | (w6233 & w6234);
assign w2594 = (in0_97 & w563) | (in0_97 & w5271) | (w563 & w5271);
assign w2595 = (w517 & w7044) | (w517 & w7045) | (w7044 & w7045);
assign w2596 = ~w2593 & w2595;
assign w2597 = ~w1142 & w5272;
assign w2598 = (w1096 & w6235) | (w1096 & w6236) | (w6235 & w6236);
assign w2599 = (in2_97 & w1142) | (in2_97 & w5273) | (w1142 & w5273);
assign w2600 = (w1096 & w7046) | (w1096 & w7047) | (w7046 & w7047);
assign w2601 = ~w2598 & w2600;
assign w2602 = w2596 & ~w2601;
assign w2603 = ~w1142 & w5274;
assign w2604 = (w1096 & w6237) | (w1096 & w6238) | (w6237 & w6238);
assign w2605 = (in2_96 & w1142) | (in2_96 & w5275) | (w1142 & w5275);
assign w2606 = (w1096 & w7048) | (w1096 & w7049) | (w7048 & w7049);
assign w2607 = ~w2604 & w2606;
assign w2608 = ~w563 & w5276;
assign w2609 = (w517 & w6239) | (w517 & w6240) | (w6239 & w6240);
assign w2610 = (in0_96 & w563) | (in0_96 & w5277) | (w563 & w5277);
assign w2611 = (w517 & w7050) | (w517 & w7051) | (w7050 & w7051);
assign w2612 = ~w2609 & w2611;
assign w2613 = w2607 & ~w2612;
assign w2614 = ~w2602 & w2613;
assign w2615 = w2584 & ~w2589;
assign w2616 = ~w2596 & w2601;
assign w2617 = ~w2615 & ~w2616;
assign w2618 = ~w2614 & w2617;
assign w2619 = (~w2578 & w2618) | (~w2578 & w4876) | (w2618 & w4876);
assign w2620 = w2571 & ~w2619;
assign w2621 = (~w518 & w4877) | (~w518 & w4878) | (w4877 & w4878);
assign w2622 = (w518 & w4879) | (w518 & w4880) | (w4879 & w4880);
assign w2623 = ~w2621 & ~w2622;
assign w2624 = (~w1097 & w4881) | (~w1097 & w4882) | (w4881 & w4882);
assign w2625 = (w1097 & w4883) | (w1097 & w4884) | (w4883 & w4884);
assign w2626 = ~w2624 & ~w2625;
assign w2627 = ~w2623 & w2626;
assign w2628 = w2623 & ~w2626;
assign w2629 = ~w1142 & w5278;
assign w2630 = (w1096 & w6241) | (w1096 & w6242) | (w6241 & w6242);
assign w2631 = (in2_106 & w1142) | (in2_106 & w5279) | (w1142 & w5279);
assign w2632 = (w1096 & w7052) | (w1096 & w7053) | (w7052 & w7053);
assign w2633 = ~w2630 & w2632;
assign w2634 = ~w563 & w5280;
assign w2635 = (w517 & w6243) | (w517 & w6244) | (w6243 & w6244);
assign w2636 = (in0_106 & w563) | (in0_106 & w5281) | (w563 & w5281);
assign w2637 = (w517 & w7054) | (w517 & w7055) | (w7054 & w7055);
assign w2638 = ~w2635 & w2637;
assign w2639 = ~w2633 & w2638;
assign w2640 = ~w2628 & ~w2639;
assign w2641 = ~w563 & w5282;
assign w2642 = (w517 & w6245) | (w517 & w6246) | (w6245 & w6246);
assign w2643 = (in0_105 & w563) | (in0_105 & w5283) | (w563 & w5283);
assign w2644 = (w517 & w7056) | (w517 & w7057) | (w7056 & w7057);
assign w2645 = ~w2642 & w2644;
assign w2646 = ~w1142 & w5284;
assign w2647 = (w1096 & w6247) | (w1096 & w6248) | (w6247 & w6248);
assign w2648 = (in2_105 & w1142) | (in2_105 & w5285) | (w1142 & w5285);
assign w2649 = (w1096 & w7058) | (w1096 & w7059) | (w7058 & w7059);
assign w2650 = ~w2647 & w2649;
assign w2651 = w2645 & ~w2650;
assign w2652 = ~w1142 & w5286;
assign w2653 = (w1096 & w6249) | (w1096 & w6250) | (w6249 & w6250);
assign w2654 = (in2_104 & w1142) | (in2_104 & w5287) | (w1142 & w5287);
assign w2655 = (w1096 & w7060) | (w1096 & w7061) | (w7060 & w7061);
assign w2656 = ~w2653 & w2655;
assign w2657 = ~w563 & w5288;
assign w2658 = (w517 & w6251) | (w517 & w6252) | (w6251 & w6252);
assign w2659 = (in0_104 & w563) | (in0_104 & w5289) | (w563 & w5289);
assign w2660 = (w517 & w7062) | (w517 & w7063) | (w7062 & w7063);
assign w2661 = ~w2658 & w2660;
assign w2662 = w2656 & ~w2661;
assign w2663 = ~w2651 & w2662;
assign w2664 = w2633 & ~w2638;
assign w2665 = ~w2645 & w2650;
assign w2666 = ~w2664 & ~w2665;
assign w2667 = ~w2663 & w2666;
assign w2668 = (~w2627 & w2667) | (~w2627 & w4897) | (w2667 & w4897);
assign w2669 = ~w2555 & w2560;
assign w2670 = ~w2566 & w2569;
assign w2671 = ~w2669 & ~w2670;
assign w2672 = w2563 & ~w2671;
assign w2673 = ~w2535 & w2538;
assign w2674 = w2544 & ~w2549;
assign w2675 = ~w2539 & w2674;
assign w2676 = ~w2673 & ~w2675;
assign w2677 = ~w2672 & w2676;
assign w2678 = w2668 & w2677;
assign w2679 = ~w2620 & w2678;
assign w2680 = ~w2107 & w2112;
assign w2681 = ~w2157 & w2162;
assign w2682 = ~w2145 & w2150;
assign w2683 = ~w2681 & ~w2682;
assign w2684 = w2152 & ~w2683;
assign w2685 = ~w2098 & w2101;
assign w2686 = w2134 & ~w2139;
assign w2687 = ~w2685 & ~w2686;
assign w2688 = ~w2684 & w2687;
assign w2689 = w2128 & ~w2688;
assign w2690 = (~w518 & w4898) | (~w518 & w4899) | (w4898 & w4899);
assign w2691 = (w518 & w4900) | (w518 & w4901) | (w4900 & w4901);
assign w2692 = ~w2690 & ~w2691;
assign w2693 = (~w1097 & w4902) | (~w1097 & w4903) | (w4902 & w4903);
assign w2694 = (w1097 & w4904) | (w1097 & w4905) | (w4904 & w4905);
assign w2695 = ~w2693 & ~w2694;
assign w2696 = w2692 & ~w2695;
assign w2697 = ~w563 & w5290;
assign w2698 = (w517 & w6253) | (w517 & w6254) | (w6253 & w6254);
assign w2699 = (in0_92 & w563) | (in0_92 & w5291) | (w563 & w5291);
assign w2700 = (w517 & w7064) | (w517 & w7065) | (w7064 & w7065);
assign w2701 = ~w2698 & w2700;
assign w2702 = ~w1142 & w5292;
assign w2703 = (w1096 & w6255) | (w1096 & w6256) | (w6255 & w6256);
assign w2704 = (in2_92 & w1142) | (in2_92 & w5293) | (w1142 & w5293);
assign w2705 = (w1096 & w7066) | (w1096 & w7067) | (w7066 & w7067);
assign w2706 = ~w2703 & w2705;
assign w2707 = ~w2701 & w2706;
assign w2708 = ~w563 & w5294;
assign w2709 = (w517 & w6257) | (w517 & w6258) | (w6257 & w6258);
assign w2710 = (in0_93 & w563) | (in0_93 & w5295) | (w563 & w5295);
assign w2711 = (w517 & w7068) | (w517 & w7069) | (w7068 & w7069);
assign w2712 = ~w2709 & w2711;
assign w2713 = ~w1142 & w5296;
assign w2714 = (w1096 & w6259) | (w1096 & w6260) | (w6259 & w6260);
assign w2715 = (in2_93 & w1142) | (in2_93 & w5297) | (w1142 & w5297);
assign w2716 = (w1096 & w7070) | (w1096 & w7071) | (w7070 & w7071);
assign w2717 = ~w2714 & w2716;
assign w2718 = ~w2712 & w2717;
assign w2719 = ~w2707 & ~w2718;
assign w2720 = w2712 & ~w2717;
assign w2721 = ~w1142 & w5298;
assign w2722 = (w1096 & w6261) | (w1096 & w6262) | (w6261 & w6262);
assign w2723 = (in2_94 & w1142) | (in2_94 & w5299) | (w1142 & w5299);
assign w2724 = (w1096 & w7072) | (w1096 & w7073) | (w7072 & w7073);
assign w2725 = ~w2722 & w2724;
assign w2726 = ~w563 & w5300;
assign w2727 = (w517 & w6263) | (w517 & w6264) | (w6263 & w6264);
assign w2728 = (in0_94 & w563) | (in0_94 & w5301) | (w563 & w5301);
assign w2729 = (w517 & w7074) | (w517 & w7075) | (w7074 & w7075);
assign w2730 = ~w2727 & w2729;
assign w2731 = ~w2725 & w2730;
assign w2732 = ~w2720 & ~w2731;
assign w2733 = ~w2719 & w2732;
assign w2734 = ~w2692 & w2695;
assign w2735 = w2725 & ~w2730;
assign w2736 = ~w2734 & ~w2735;
assign w2737 = (~w2696 & w2733) | (~w2696 & w4918) | (w2733 & w4918);
assign w2738 = w2084 & ~w2087;
assign w2739 = ~w2095 & w2738;
assign w2740 = ~w2091 & w2094;
assign w2741 = w2118 & ~w2123;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = ~w2739 & w2742;
assign w2744 = w2125 & ~w2743;
assign w2745 = ~w2680 & ~w2689;
assign w2746 = ~w2737 & ~w2744;
assign w2747 = w2745 & w2746;
assign w2748 = w2679 & w2747;
assign w2749 = ~w2532 & w2748;
assign w2750 = w2508 & w2749;
assign w2751 = ~w2280 & w2750;
assign w2752 = ~w2499 & w2501;
assign w2753 = w2701 & ~w2706;
assign w2754 = ~w2696 & ~w2753;
assign w2755 = w2732 & w2754;
assign w2756 = ~w2737 & ~w2755;
assign w2757 = ~w2607 & w2612;
assign w2758 = ~w2602 & ~w2757;
assign w2759 = w2591 & w2758;
assign w2760 = w2571 & w2759;
assign w2761 = ~w2756 & w2760;
assign w2762 = w2679 & ~w2761;
assign w2763 = ~w2656 & w2661;
assign w2764 = ~w2651 & ~w2763;
assign w2765 = w2640 & w2764;
assign w2766 = w2668 & ~w2765;
assign w2767 = w2457 & ~w2462;
assign w2768 = w2451 & ~w2767;
assign w2769 = w2480 & w2768;
assign w2770 = ~w2766 & w2769;
assign w2771 = w2384 & w2770;
assign w2772 = ~w2762 & w2771;
assign w2773 = w2508 & ~w2772;
assign w2774 = ~w2752 & ~w2773;
assign w2775 = ~w2773 & w3972;
assign w2776 = ~w2751 & w2775;
assign w2777 = (~w1157 & w2773) | (~w1157 & w3973) | (w2773 & w3973);
assign w2778 = ~w1157 & w2750;
assign w2779 = ~w2280 & w2778;
assign w2780 = ~w2777 & ~w2779;
assign w2781 = ~w2776 & w2780;
assign w2782 = ~w2773 & w3974;
assign w2783 = ~w2751 & w2782;
assign w2784 = (w1163 & w2773) | (w1163 & w3975) | (w2773 & w3975);
assign w2785 = w1163 & w2750;
assign w2786 = ~w2280 & w2785;
assign w2787 = ~w2784 & ~w2786;
assign w2788 = ~w2783 & w2787;
assign w2789 = ~w2773 & w3976;
assign w2790 = ~w2751 & w2789;
assign w2791 = (~w1181 & w2773) | (~w1181 & w3977) | (w2773 & w3977);
assign w2792 = ~w1181 & w2750;
assign w2793 = ~w2280 & w2792;
assign w2794 = ~w2791 & ~w2793;
assign w2795 = ~w2790 & w2794;
assign w2796 = ~w2773 & w3978;
assign w2797 = ~w2751 & w2796;
assign w2798 = (~w1192 & w2773) | (~w1192 & w3979) | (w2773 & w3979);
assign w2799 = ~w1192 & w2750;
assign w2800 = ~w2280 & w2799;
assign w2801 = ~w2798 & ~w2800;
assign w2802 = ~w2797 & w2801;
assign w2803 = ~w2773 & w3980;
assign w2804 = ~w2751 & w2803;
assign w2805 = (~w1203 & w2773) | (~w1203 & w3981) | (w2773 & w3981);
assign w2806 = ~w1203 & w2750;
assign w2807 = ~w2280 & w2806;
assign w2808 = ~w2805 & ~w2807;
assign w2809 = ~w2804 & w2808;
assign w2810 = ~w2773 & w3982;
assign w2811 = ~w2751 & w2810;
assign w2812 = (~w1214 & w2773) | (~w1214 & w3983) | (w2773 & w3983);
assign w2813 = ~w1214 & w2750;
assign w2814 = ~w2280 & w2813;
assign w2815 = ~w2812 & ~w2814;
assign w2816 = ~w2811 & w2815;
assign w2817 = ~w2773 & w3984;
assign w2818 = ~w2751 & w2817;
assign w2819 = (~w1225 & w2773) | (~w1225 & w3985) | (w2773 & w3985);
assign w2820 = ~w1225 & w2750;
assign w2821 = ~w2280 & w2820;
assign w2822 = ~w2819 & ~w2821;
assign w2823 = ~w2818 & w2822;
assign w2824 = ~w2773 & w3986;
assign w2825 = ~w2751 & w2824;
assign w2826 = (~w1342 & w2773) | (~w1342 & w3987) | (w2773 & w3987);
assign w2827 = ~w1342 & w2750;
assign w2828 = ~w2280 & w2827;
assign w2829 = ~w2826 & ~w2828;
assign w2830 = ~w2825 & w2829;
assign w2831 = ~w2773 & w3988;
assign w2832 = ~w2751 & w2831;
assign w2833 = (~w1313 & w2773) | (~w1313 & w3989) | (w2773 & w3989);
assign w2834 = ~w1313 & w2750;
assign w2835 = ~w2280 & w2834;
assign w2836 = ~w2833 & ~w2835;
assign w2837 = ~w2832 & w2836;
assign w2838 = ~w2773 & w3990;
assign w2839 = ~w2751 & w2838;
assign w2840 = (~w1329 & w2773) | (~w1329 & w3991) | (w2773 & w3991);
assign w2841 = ~w1329 & w2750;
assign w2842 = ~w2280 & w2841;
assign w2843 = ~w2840 & ~w2842;
assign w2844 = ~w2839 & w2843;
assign w2845 = ~w2773 & w3992;
assign w2846 = ~w2751 & w2845;
assign w2847 = (~w1267 & w2773) | (~w1267 & w3993) | (w2773 & w3993);
assign w2848 = ~w1267 & w2750;
assign w2849 = ~w2280 & w2848;
assign w2850 = ~w2847 & ~w2849;
assign w2851 = ~w2846 & w2850;
assign w2852 = ~w2773 & w3994;
assign w2853 = ~w2751 & w2852;
assign w2854 = (~w1243 & w2773) | (~w1243 & w3995) | (w2773 & w3995);
assign w2855 = ~w1243 & w2750;
assign w2856 = ~w2280 & w2855;
assign w2857 = ~w2854 & ~w2856;
assign w2858 = ~w2853 & w2857;
assign w2859 = ~w2773 & w3996;
assign w2860 = ~w2751 & w2859;
assign w2861 = (~w1254 & w2773) | (~w1254 & w3997) | (w2773 & w3997);
assign w2862 = ~w1254 & w2750;
assign w2863 = ~w2280 & w2862;
assign w2864 = ~w2861 & ~w2863;
assign w2865 = ~w2860 & w2864;
assign w2866 = ~w2773 & w3998;
assign w2867 = ~w2751 & w2866;
assign w2868 = (~w1304 & w2773) | (~w1304 & w3999) | (w2773 & w3999);
assign w2869 = ~w1304 & w2750;
assign w2870 = ~w2280 & w2869;
assign w2871 = ~w2868 & ~w2870;
assign w2872 = ~w2867 & w2871;
assign w2873 = ~w2773 & w4000;
assign w2874 = ~w2751 & w2873;
assign w2875 = (~w1280 & w2773) | (~w1280 & w4001) | (w2773 & w4001);
assign w2876 = ~w1280 & w2750;
assign w2877 = ~w2280 & w2876;
assign w2878 = ~w2875 & ~w2877;
assign w2879 = ~w2874 & w2878;
assign w2880 = ~w2773 & w4002;
assign w2881 = ~w2751 & w2880;
assign w2882 = (~w1291 & w2773) | (~w1291 & w4003) | (w2773 & w4003);
assign w2883 = ~w1291 & w2750;
assign w2884 = ~w2280 & w2883;
assign w2885 = ~w2882 & ~w2884;
assign w2886 = ~w2881 & w2885;
assign w2887 = ~w2773 & w4004;
assign w2888 = ~w2751 & w2887;
assign w2889 = (~w1429 & w2773) | (~w1429 & w4005) | (w2773 & w4005);
assign w2890 = ~w1429 & w2750;
assign w2891 = ~w2280 & w2890;
assign w2892 = ~w2889 & ~w2891;
assign w2893 = ~w2888 & w2892;
assign w2894 = ~w2773 & w4006;
assign w2895 = ~w2751 & w2894;
assign w2896 = (w1435 & w2773) | (w1435 & w4007) | (w2773 & w4007);
assign w2897 = w1435 & w2750;
assign w2898 = ~w2280 & w2897;
assign w2899 = ~w2896 & ~w2898;
assign w2900 = ~w2895 & w2899;
assign w2901 = ~w2773 & w4008;
assign w2902 = ~w2751 & w2901;
assign w2903 = (~w1381 & w2773) | (~w1381 & w4009) | (w2773 & w4009);
assign w2904 = ~w1381 & w2750;
assign w2905 = ~w2280 & w2904;
assign w2906 = ~w2903 & ~w2905;
assign w2907 = ~w2902 & w2906;
assign w2908 = ~w2773 & w4010;
assign w2909 = ~w2751 & w2908;
assign w2910 = (~w1370 & w2773) | (~w1370 & w4011) | (w2773 & w4011);
assign w2911 = ~w1370 & w2750;
assign w2912 = ~w2280 & w2911;
assign w2913 = ~w2910 & ~w2912;
assign w2914 = ~w2909 & w2913;
assign w2915 = ~w2773 & w4012;
assign w2916 = ~w2751 & w2915;
assign w2917 = (~w1394 & w2773) | (~w1394 & w4013) | (w2773 & w4013);
assign w2918 = ~w1394 & w2750;
assign w2919 = ~w2280 & w2918;
assign w2920 = ~w2917 & ~w2919;
assign w2921 = ~w2916 & w2920;
assign w2922 = ~w2773 & w4014;
assign w2923 = ~w2751 & w2922;
assign w2924 = (~w1403 & w2773) | (~w1403 & w4015) | (w2773 & w4015);
assign w2925 = ~w1403 & w2750;
assign w2926 = ~w2280 & w2925;
assign w2927 = ~w2924 & ~w2926;
assign w2928 = ~w2923 & w2927;
assign w2929 = ~w2773 & w4016;
assign w2930 = ~w2751 & w2929;
assign w2931 = (~w1414 & w2773) | (~w1414 & w4017) | (w2773 & w4017);
assign w2932 = ~w1414 & w2750;
assign w2933 = ~w2280 & w2932;
assign w2934 = ~w2931 & ~w2933;
assign w2935 = ~w2930 & w2934;
assign w2936 = ~w2773 & w4018;
assign w2937 = ~w2751 & w2936;
assign w2938 = (~w1529 & w2773) | (~w1529 & w4019) | (w2773 & w4019);
assign w2939 = ~w1529 & w2750;
assign w2940 = ~w2280 & w2939;
assign w2941 = ~w2938 & ~w2940;
assign w2942 = ~w2937 & w2941;
assign w2943 = ~w2773 & w4020;
assign w2944 = ~w2751 & w2943;
assign w2945 = (~w1513 & w2773) | (~w1513 & w4021) | (w2773 & w4021);
assign w2946 = ~w1513 & w2750;
assign w2947 = ~w2280 & w2946;
assign w2948 = ~w2945 & ~w2947;
assign w2949 = ~w2944 & w2948;
assign w2950 = ~w2773 & w4022;
assign w2951 = ~w2751 & w2950;
assign w2952 = (~w1520 & w2773) | (~w1520 & w4023) | (w2773 & w4023);
assign w2953 = ~w1520 & w2750;
assign w2954 = ~w2280 & w2953;
assign w2955 = ~w2952 & ~w2954;
assign w2956 = ~w2951 & w2955;
assign w2957 = ~w2773 & w4024;
assign w2958 = ~w2751 & w2957;
assign w2959 = (~w1478 & w2773) | (~w1478 & w4025) | (w2773 & w4025);
assign w2960 = ~w1478 & w2750;
assign w2961 = ~w2280 & w2960;
assign w2962 = ~w2959 & ~w2961;
assign w2963 = ~w2958 & w2962;
assign w2964 = ~w2773 & w4026;
assign w2965 = ~w2751 & w2964;
assign w2966 = (~w1462 & w2773) | (~w1462 & w4027) | (w2773 & w4027);
assign w2967 = ~w1462 & w2750;
assign w2968 = ~w2280 & w2967;
assign w2969 = ~w2966 & ~w2968;
assign w2970 = ~w2965 & w2969;
assign w2971 = ~w2773 & w4028;
assign w2972 = ~w2751 & w2971;
assign w2973 = (~w1469 & w2773) | (~w1469 & w4029) | (w2773 & w4029);
assign w2974 = ~w1469 & w2750;
assign w2975 = ~w2280 & w2974;
assign w2976 = ~w2973 & ~w2975;
assign w2977 = ~w2972 & w2976;
assign w2978 = ~w2773 & w4030;
assign w2979 = ~w2751 & w2978;
assign w2980 = (~w1503 & w2773) | (~w1503 & w4031) | (w2773 & w4031);
assign w2981 = ~w1503 & w2750;
assign w2982 = ~w2280 & w2981;
assign w2983 = ~w2980 & ~w2982;
assign w2984 = ~w2979 & w2983;
assign w2985 = ~w2773 & w4032;
assign w2986 = ~w2751 & w2985;
assign w2987 = (~w1487 & w2773) | (~w1487 & w4033) | (w2773 & w4033);
assign w2988 = ~w1487 & w2750;
assign w2989 = ~w2280 & w2988;
assign w2990 = ~w2987 & ~w2989;
assign w2991 = ~w2986 & w2990;
assign w2992 = ~w2773 & w4034;
assign w2993 = ~w2751 & w2992;
assign w2994 = (~w1494 & w2773) | (~w1494 & w4035) | (w2773 & w4035);
assign w2995 = ~w1494 & w2750;
assign w2996 = ~w2280 & w2995;
assign w2997 = ~w2994 & ~w2996;
assign w2998 = ~w2993 & w2997;
assign w2999 = ~w2773 & w4036;
assign w3000 = ~w2751 & w2999;
assign w3001 = (w1623 & w2773) | (w1623 & w4037) | (w2773 & w4037);
assign w3002 = w1623 & w2750;
assign w3003 = ~w2280 & w3002;
assign w3004 = ~w3001 & ~w3003;
assign w3005 = ~w3000 & w3004;
assign w3006 = ~w2773 & w4038;
assign w3007 = ~w2751 & w3006;
assign w3008 = (~w1639 & w2773) | (~w1639 & w4039) | (w2773 & w4039);
assign w3009 = ~w1639 & w2750;
assign w3010 = ~w2280 & w3009;
assign w3011 = ~w3008 & ~w3010;
assign w3012 = ~w3007 & w3011;
assign w3013 = ~w2773 & w4040;
assign w3014 = ~w2751 & w3013;
assign w3015 = (w1645 & w2773) | (w1645 & w4041) | (w2773 & w4041);
assign w3016 = w1645 & w2750;
assign w3017 = ~w2280 & w3016;
assign w3018 = ~w3015 & ~w3017;
assign w3019 = ~w3014 & w3018;
assign w3020 = ~w2773 & w4042;
assign w3021 = ~w2751 & w3020;
assign w3022 = (~w1685 & w2773) | (~w1685 & w4043) | (w2773 & w4043);
assign w3023 = ~w1685 & w2750;
assign w3024 = ~w2280 & w3023;
assign w3025 = ~w3022 & ~w3024;
assign w3026 = ~w3021 & w3025;
assign w3027 = ~w2773 & w4044;
assign w3028 = ~w2751 & w3027;
assign w3029 = (~w1678 & w2773) | (~w1678 & w4045) | (w2773 & w4045);
assign w3030 = ~w1678 & w2750;
assign w3031 = ~w2280 & w3030;
assign w3032 = ~w3029 & ~w3031;
assign w3033 = ~w3028 & w3032;
assign w3034 = ~w2773 & w4046;
assign w3035 = ~w2751 & w3034;
assign w3036 = (~w1663 & w2773) | (~w1663 & w4047) | (w2773 & w4047);
assign w3037 = ~w1663 & w2750;
assign w3038 = ~w2280 & w3037;
assign w3039 = ~w3036 & ~w3038;
assign w3040 = ~w3035 & w3039;
assign w3041 = ~w2773 & w4048;
assign w3042 = ~w2751 & w3041;
assign w3043 = (w1667 & w2773) | (w1667 & w4049) | (w2773 & w4049);
assign w3044 = w1667 & w2750;
assign w3045 = ~w2280 & w3044;
assign w3046 = ~w3043 & ~w3045;
assign w3047 = ~w3042 & w3046;
assign w3048 = ~w2773 & w4050;
assign w3049 = ~w2751 & w3048;
assign w3050 = (~w1553 & w2773) | (~w1553 & w4051) | (w2773 & w4051);
assign w3051 = ~w1553 & w2750;
assign w3052 = ~w2280 & w3051;
assign w3053 = ~w3050 & ~w3052;
assign w3054 = ~w3049 & w3053;
assign w3055 = ~w2773 & w4052;
assign w3056 = ~w2751 & w3055;
assign w3057 = (~w1567 & w2773) | (~w1567 & w4053) | (w2773 & w4053);
assign w3058 = ~w1567 & w2750;
assign w3059 = ~w2280 & w3058;
assign w3060 = ~w3057 & ~w3059;
assign w3061 = ~w3056 & w3060;
assign w3062 = ~w2773 & w4054;
assign w3063 = ~w2751 & w3062;
assign w3064 = (~w1574 & w2773) | (~w1574 & w4055) | (w2773 & w4055);
assign w3065 = ~w1574 & w2750;
assign w3066 = ~w2280 & w3065;
assign w3067 = ~w3064 & ~w3066;
assign w3068 = ~w3063 & w3067;
assign w3069 = ~w2773 & w4056;
assign w3070 = ~w2751 & w3069;
assign w3071 = (~w1610 & w2773) | (~w1610 & w4057) | (w2773 & w4057);
assign w3072 = ~w1610 & w2750;
assign w3073 = ~w2280 & w3072;
assign w3074 = ~w3071 & ~w3073;
assign w3075 = ~w3070 & w3074;
assign w3076 = ~w2773 & w4058;
assign w3077 = ~w2751 & w3076;
assign w3078 = (~w1596 & w2773) | (~w1596 & w4059) | (w2773 & w4059);
assign w3079 = ~w1596 & w2750;
assign w3080 = ~w2280 & w3079;
assign w3081 = ~w3078 & ~w3080;
assign w3082 = ~w3077 & w3081;
assign w3083 = ~w2773 & w4060;
assign w3084 = ~w2751 & w3083;
assign w3085 = (~w1603 & w2773) | (~w1603 & w4061) | (w2773 & w4061);
assign w3086 = ~w1603 & w2750;
assign w3087 = ~w2280 & w3086;
assign w3088 = ~w3085 & ~w3087;
assign w3089 = ~w3084 & w3088;
assign w3090 = ~w2773 & w4062;
assign w3091 = ~w2751 & w3090;
assign w3092 = (~w1560 & w2773) | (~w1560 & w4063) | (w2773 & w4063);
assign w3093 = ~w1560 & w2750;
assign w3094 = ~w2280 & w3093;
assign w3095 = ~w3092 & ~w3094;
assign w3096 = ~w3091 & w3095;
assign w3097 = ~w2773 & w4064;
assign w3098 = ~w2751 & w3097;
assign w3099 = (w1578 & w2773) | (w1578 & w4065) | (w2773 & w4065);
assign w3100 = w1578 & w2750;
assign w3101 = ~w2280 & w3100;
assign w3102 = ~w3099 & ~w3101;
assign w3103 = ~w3098 & w3102;
assign w3104 = ~w2773 & w4066;
assign w3105 = ~w2751 & w3104;
assign w3106 = (~w1588 & w2773) | (~w1588 & w4067) | (w2773 & w4067);
assign w3107 = ~w1588 & w2750;
assign w3108 = ~w2280 & w3107;
assign w3109 = ~w3106 & ~w3108;
assign w3110 = ~w3105 & w3109;
assign w3111 = ~w2773 & w4068;
assign w3112 = ~w2751 & w3111;
assign w3113 = (w1773 & w2773) | (w1773 & w4069) | (w2773 & w4069);
assign w3114 = w1773 & w2750;
assign w3115 = ~w2280 & w3114;
assign w3116 = ~w3113 & ~w3115;
assign w3117 = ~w3112 & w3116;
assign w3118 = ~w2773 & w4070;
assign w3119 = ~w2751 & w3118;
assign w3120 = (~w1767 & w2773) | (~w1767 & w4071) | (w2773 & w4071);
assign w3121 = ~w1767 & w2750;
assign w3122 = ~w2280 & w3121;
assign w3123 = ~w3120 & ~w3122;
assign w3124 = ~w3119 & w3123;
assign w3125 = ~w2773 & w4072;
assign w3126 = ~w2751 & w3125;
assign w3127 = (w1786 & w2773) | (w1786 & w4073) | (w2773 & w4073);
assign w3128 = w1786 & w2750;
assign w3129 = ~w2280 & w3128;
assign w3130 = ~w3127 & ~w3129;
assign w3131 = ~w3126 & w3130;
assign w3132 = ~w2773 & w4074;
assign w3133 = ~w2751 & w3132;
assign w3134 = (~w1740 & w2773) | (~w1740 & w4075) | (w2773 & w4075);
assign w3135 = ~w1740 & w2750;
assign w3136 = ~w2280 & w3135;
assign w3137 = ~w3134 & ~w3136;
assign w3138 = ~w3133 & w3137;
assign w3139 = ~w2773 & w4076;
assign w3140 = ~w2751 & w3139;
assign w3141 = (~w1729 & w2773) | (~w1729 & w4077) | (w2773 & w4077);
assign w3142 = ~w1729 & w2750;
assign w3143 = ~w2280 & w3142;
assign w3144 = ~w3141 & ~w3143;
assign w3145 = ~w3140 & w3144;
assign w3146 = ~w2773 & w4078;
assign w3147 = ~w2751 & w3146;
assign w3148 = (~w1753 & w2773) | (~w1753 & w4079) | (w2773 & w4079);
assign w3149 = ~w1753 & w2750;
assign w3150 = ~w2280 & w3149;
assign w3151 = ~w3148 & ~w3150;
assign w3152 = ~w3147 & w3151;
assign w3153 = ~w2773 & w4080;
assign w3154 = ~w2751 & w3153;
assign w3155 = (w1711 & w2773) | (w1711 & w4081) | (w2773 & w4081);
assign w3156 = w1711 & w2750;
assign w3157 = ~w2280 & w3156;
assign w3158 = ~w3155 & ~w3157;
assign w3159 = ~w3154 & w3158;
assign w3160 = ~w2773 & w4082;
assign w3161 = ~w2751 & w3160;
assign w3162 = (~w1704 & w2773) | (~w1704 & w4083) | (w2773 & w4083);
assign w3163 = ~w1704 & w2750;
assign w3164 = ~w2280 & w3163;
assign w3165 = ~w3162 & ~w3164;
assign w3166 = ~w3161 & w3165;
assign w3167 = ~w2773 & w4084;
assign w3168 = ~w2751 & w3167;
assign w3169 = (~w1868 & w2773) | (~w1868 & w4085) | (w2773 & w4085);
assign w3170 = ~w1868 & w2750;
assign w3171 = ~w2280 & w3170;
assign w3172 = ~w3169 & ~w3171;
assign w3173 = ~w3168 & w3172;
assign w3174 = ~w2773 & w4086;
assign w3175 = ~w2751 & w3174;
assign w3176 = (~w1857 & w2773) | (~w1857 & w4087) | (w2773 & w4087);
assign w3177 = ~w1857 & w2750;
assign w3178 = ~w2280 & w3177;
assign w3179 = ~w3176 & ~w3178;
assign w3180 = ~w3175 & w3179;
assign w3181 = ~w2773 & w4088;
assign w3182 = ~w2751 & w3181;
assign w3183 = (~w1881 & w2773) | (~w1881 & w4089) | (w2773 & w4089);
assign w3184 = ~w1881 & w2750;
assign w3185 = ~w2280 & w3184;
assign w3186 = ~w3183 & ~w3185;
assign w3187 = ~w3182 & w3186;
assign w3188 = ~w2773 & w4090;
assign w3189 = ~w2751 & w3188;
assign w3190 = (~w1906 & w2773) | (~w1906 & w4091) | (w2773 & w4091);
assign w3191 = ~w1906 & w2750;
assign w3192 = ~w2280 & w3191;
assign w3193 = ~w3190 & ~w3192;
assign w3194 = ~w3189 & w3193;
assign w3195 = ~w2773 & w4092;
assign w3196 = ~w2751 & w3195;
assign w3197 = (~w1895 & w2773) | (~w1895 & w4093) | (w2773 & w4093);
assign w3198 = ~w1895 & w2750;
assign w3199 = ~w2280 & w3198;
assign w3200 = ~w3197 & ~w3199;
assign w3201 = ~w3196 & w3200;
assign w3202 = ~w2773 & w4094;
assign w3203 = ~w2751 & w3202;
assign w3204 = (~w1938 & w2773) | (~w1938 & w4095) | (w2773 & w4095);
assign w3205 = ~w1938 & w2750;
assign w3206 = ~w2280 & w3205;
assign w3207 = ~w3204 & ~w3206;
assign w3208 = ~w3203 & w3207;
assign w3209 = ~w2773 & w4096;
assign w3210 = ~w2751 & w3209;
assign w3211 = (w1913 & w2773) | (w1913 & w4097) | (w2773 & w4097);
assign w3212 = w1913 & w2750;
assign w3213 = ~w2280 & w3212;
assign w3214 = ~w3211 & ~w3213;
assign w3215 = ~w3210 & w3214;
assign w3216 = ~w2773 & w4098;
assign w3217 = ~w2751 & w3216;
assign w3218 = (~w1923 & w2773) | (~w1923 & w4099) | (w2773 & w4099);
assign w3219 = ~w1923 & w2750;
assign w3220 = ~w2280 & w3219;
assign w3221 = ~w3218 & ~w3220;
assign w3222 = ~w3217 & w3221;
assign w3223 = ~w2773 & w4100;
assign w3224 = ~w2751 & w3223;
assign w3225 = (w1979 & w2773) | (w1979 & w4101) | (w2773 & w4101);
assign w3226 = w1979 & w2750;
assign w3227 = ~w2280 & w3226;
assign w3228 = ~w3225 & ~w3227;
assign w3229 = ~w3224 & w3228;
assign w3230 = ~w2773 & w4102;
assign w3231 = ~w2751 & w3230;
assign w3232 = (~w1973 & w2773) | (~w1973 & w4103) | (w2773 & w4103);
assign w3233 = ~w1973 & w2750;
assign w3234 = ~w2280 & w3233;
assign w3235 = ~w3232 & ~w3234;
assign w3236 = ~w3231 & w3235;
assign w3237 = ~w2773 & w4104;
assign w3238 = ~w2751 & w3237;
assign w3239 = (w1955 & w2773) | (w1955 & w4105) | (w2773 & w4105);
assign w3240 = w1955 & w2750;
assign w3241 = ~w2280 & w3240;
assign w3242 = ~w3239 & ~w3241;
assign w3243 = ~w3238 & w3242;
assign w3244 = ~w2773 & w4106;
assign w3245 = ~w2751 & w3244;
assign w3246 = (~w1949 & w2773) | (~w1949 & w4107) | (w2773 & w4107);
assign w3247 = ~w1949 & w2750;
assign w3248 = ~w2280 & w3247;
assign w3249 = ~w3246 & ~w3248;
assign w3250 = ~w3245 & w3249;
assign w3251 = ~w2773 & w4108;
assign w3252 = ~w2751 & w3251;
assign w3253 = (~w2007 & w2773) | (~w2007 & w4109) | (w2773 & w4109);
assign w3254 = ~w2007 & w2750;
assign w3255 = ~w2280 & w3254;
assign w3256 = ~w3253 & ~w3255;
assign w3257 = ~w3252 & w3256;
assign w3258 = ~w2773 & w4110;
assign w3259 = ~w2751 & w3258;
assign w3260 = (~w2018 & w2773) | (~w2018 & w4111) | (w2773 & w4111);
assign w3261 = ~w2018 & w2750;
assign w3262 = ~w2280 & w3261;
assign w3263 = ~w3260 & ~w3262;
assign w3264 = ~w3259 & w3263;
assign w3265 = ~w2773 & w4112;
assign w3266 = ~w2751 & w3265;
assign w3267 = (w2033 & w2773) | (w2033 & w4113) | (w2773 & w4113);
assign w3268 = w2033 & w2750;
assign w3269 = ~w2280 & w3268;
assign w3270 = ~w3267 & ~w3269;
assign w3271 = ~w3266 & w3270;
assign w3272 = ~w2773 & w4114;
assign w3273 = ~w2751 & w3272;
assign w3274 = (~w2026 & w2773) | (~w2026 & w4115) | (w2773 & w4115);
assign w3275 = ~w2026 & w2750;
assign w3276 = ~w2280 & w3275;
assign w3277 = ~w3274 & ~w3276;
assign w3278 = ~w3273 & w3277;
assign w3279 = ~w2773 & w4116;
assign w3280 = ~w2751 & w3279;
assign w3281 = (w2213 & w2773) | (w2213 & w4117) | (w2773 & w4117);
assign w3282 = w2213 & w2750;
assign w3283 = ~w2280 & w3282;
assign w3284 = ~w3281 & ~w3283;
assign w3285 = ~w3280 & w3284;
assign w3286 = ~w2773 & w4118;
assign w3287 = ~w2751 & w3286;
assign w3288 = (~w2229 & w2773) | (~w2229 & w4119) | (w2773 & w4119);
assign w3289 = ~w2229 & w2750;
assign w3290 = ~w2280 & w3289;
assign w3291 = ~w3288 & ~w3290;
assign w3292 = ~w3287 & w3291;
assign w3293 = ~w2773 & w4120;
assign w3294 = ~w2751 & w3293;
assign w3295 = (w2264 & w2773) | (w2264 & w4121) | (w2773 & w4121);
assign w3296 = w2264 & w2750;
assign w3297 = ~w2280 & w3296;
assign w3298 = ~w3295 & ~w3297;
assign w3299 = ~w3294 & w3298;
assign w3300 = ~w2773 & w4122;
assign w3301 = ~w2751 & w3300;
assign w3302 = (~w2247 & w2773) | (~w2247 & w4123) | (w2773 & w4123);
assign w3303 = ~w2247 & w2750;
assign w3304 = ~w2280 & w3303;
assign w3305 = ~w3302 & ~w3304;
assign w3306 = ~w3301 & w3305;
assign w3307 = ~w2773 & w4124;
assign w3308 = ~w2751 & w3307;
assign w3309 = (~w2258 & w2773) | (~w2258 & w4125) | (w2773 & w4125);
assign w3310 = ~w2258 & w2750;
assign w3311 = ~w2280 & w3310;
assign w3312 = ~w3309 & ~w3311;
assign w3313 = ~w3308 & w3312;
assign w3314 = ~w2773 & w4126;
assign w3315 = ~w2751 & w3314;
assign w3316 = (~w2206 & w2773) | (~w2206 & w4127) | (w2773 & w4127);
assign w3317 = ~w2206 & w2750;
assign w3318 = ~w2280 & w3317;
assign w3319 = ~w3316 & ~w3318;
assign w3320 = ~w3315 & w3319;
assign w3321 = ~w2773 & w4128;
assign w3322 = ~w2751 & w3321;
assign w3323 = (w2192 & w2773) | (w2192 & w4129) | (w2773 & w4129);
assign w3324 = w2192 & w2750;
assign w3325 = ~w2280 & w3324;
assign w3326 = ~w3323 & ~w3325;
assign w3327 = ~w3322 & w3326;
assign w3328 = ~w2773 & w4130;
assign w3329 = ~w2751 & w3328;
assign w3330 = (~w2236 & w2773) | (~w2236 & w4131) | (w2773 & w4131);
assign w3331 = ~w2236 & w2750;
assign w3332 = ~w2280 & w3331;
assign w3333 = ~w3330 & ~w3332;
assign w3334 = ~w3329 & w3333;
assign w3335 = ~w2773 & w4132;
assign w3336 = ~w2751 & w3335;
assign w3337 = (w2181 & w2773) | (w2181 & w4133) | (w2773 & w4133);
assign w3338 = w2181 & w2750;
assign w3339 = ~w2280 & w3338;
assign w3340 = ~w3337 & ~w3339;
assign w3341 = ~w3336 & w3340;
assign w3342 = ~w2773 & w4134;
assign w3343 = ~w2751 & w3342;
assign w3344 = (~w2169 & w2773) | (~w2169 & w4135) | (w2773 & w4135);
assign w3345 = ~w2169 & w2750;
assign w3346 = ~w2280 & w3345;
assign w3347 = ~w3344 & ~w3346;
assign w3348 = ~w3343 & w3347;
assign w3349 = ~w2773 & w4136;
assign w3350 = ~w2751 & w3349;
assign w3351 = (w2079 & w2773) | (w2079 & w4137) | (w2773 & w4137);
assign w3352 = w2079 & w2750;
assign w3353 = ~w2280 & w3352;
assign w3354 = ~w3351 & ~w3353;
assign w3355 = ~w3350 & w3354;
assign w3356 = ~w2773 & w4138;
assign w3357 = ~w2751 & w3356;
assign w3358 = (~w2075 & w2773) | (~w2075 & w4139) | (w2773 & w4139);
assign w3359 = ~w2075 & w2750;
assign w3360 = ~w2280 & w3359;
assign w3361 = ~w3358 & ~w3360;
assign w3362 = ~w3357 & w3361;
assign w3363 = ~w2773 & w4140;
assign w3364 = ~w2751 & w3363;
assign w3365 = (~w2162 & w2773) | (~w2162 & w4141) | (w2773 & w4141);
assign w3366 = ~w2162 & w2750;
assign w3367 = ~w2280 & w3366;
assign w3368 = ~w3365 & ~w3367;
assign w3369 = ~w3364 & w3368;
assign w3370 = ~w2773 & w4142;
assign w3371 = ~w2751 & w3370;
assign w3372 = (~w2150 & w2773) | (~w2150 & w4143) | (w2773 & w4143);
assign w3373 = ~w2150 & w2750;
assign w3374 = ~w2280 & w3373;
assign w3375 = ~w3372 & ~w3374;
assign w3376 = ~w3371 & w3375;
assign w3377 = ~w2773 & w4144;
assign w3378 = ~w2751 & w3377;
assign w3379 = (w2134 & w2773) | (w2134 & w4145) | (w2773 & w4145);
assign w3380 = w2134 & w2750;
assign w3381 = ~w2280 & w3380;
assign w3382 = ~w3379 & ~w3381;
assign w3383 = ~w3378 & w3382;
assign w3384 = ~w2773 & w4146;
assign w3385 = ~w2751 & w3384;
assign w3386 = (~w2101 & w2773) | (~w2101 & w4147) | (w2773 & w4147);
assign w3387 = ~w2101 & w2750;
assign w3388 = ~w2280 & w3387;
assign w3389 = ~w3386 & ~w3388;
assign w3390 = ~w3385 & w3389;
assign w3391 = ~w2773 & w4148;
assign w3392 = ~w2751 & w3391;
assign w3393 = (w2084 & w2773) | (w2084 & w4149) | (w2773 & w4149);
assign w3394 = w2084 & w2750;
assign w3395 = ~w2280 & w3394;
assign w3396 = ~w3393 & ~w3395;
assign w3397 = ~w3392 & w3396;
assign w3398 = ~w2773 & w4150;
assign w3399 = ~w2751 & w3398;
assign w3400 = (~w2094 & w2773) | (~w2094 & w4151) | (w2773 & w4151);
assign w3401 = ~w2094 & w2750;
assign w3402 = ~w2280 & w3401;
assign w3403 = ~w3400 & ~w3402;
assign w3404 = ~w3399 & w3403;
assign w3405 = ~w2773 & w4152;
assign w3406 = ~w2751 & w3405;
assign w3407 = (w2118 & w2773) | (w2118 & w4153) | (w2773 & w4153);
assign w3408 = w2118 & w2750;
assign w3409 = ~w2280 & w3408;
assign w3410 = ~w3407 & ~w3409;
assign w3411 = ~w3406 & w3410;
assign w3412 = ~w2773 & w4154;
assign w3413 = ~w2751 & w3412;
assign w3414 = (~w2112 & w2773) | (~w2112 & w4155) | (w2773 & w4155);
assign w3415 = ~w2112 & w2750;
assign w3416 = ~w2280 & w3415;
assign w3417 = ~w3414 & ~w3416;
assign w3418 = ~w3413 & w3417;
assign w3419 = ~w2773 & w4156;
assign w3420 = ~w2751 & w3419;
assign w3421 = ~w2706 & w2750;
assign w3422 = ~w2280 & w3421;
assign w3423 = (~w2706 & w2773) | (~w2706 & w4157) | (w2773 & w4157);
assign w3424 = ~w3422 & ~w3423;
assign w3425 = ~w3420 & w3424;
assign w3426 = ~w2773 & w4158;
assign w3427 = ~w2751 & w3426;
assign w3428 = ~w2717 & w2750;
assign w3429 = ~w2280 & w3428;
assign w3430 = (~w2717 & w2773) | (~w2717 & w4159) | (w2773 & w4159);
assign w3431 = ~w3429 & ~w3430;
assign w3432 = ~w3427 & w3431;
assign w3433 = ~w2773 & w4160;
assign w3434 = ~w2751 & w3433;
assign w3435 = (w2725 & w2773) | (w2725 & w4161) | (w2773 & w4161);
assign w3436 = w2725 & w2750;
assign w3437 = ~w2280 & w3436;
assign w3438 = ~w3435 & ~w3437;
assign w3439 = ~w3434 & w3438;
assign w3440 = ~w2773 & w4162;
assign w3441 = ~w2751 & w3440;
assign w3442 = ~w2695 & w2750;
assign w3443 = ~w2280 & w3442;
assign w3444 = (~w2695 & w2773) | (~w2695 & w4163) | (w2773 & w4163);
assign w3445 = ~w3443 & ~w3444;
assign w3446 = ~w3441 & w3445;
assign w3447 = ~w2773 & w4164;
assign w3448 = ~w2751 & w3447;
assign w3449 = (w2607 & w2773) | (w2607 & w4165) | (w2773 & w4165);
assign w3450 = w2607 & w2750;
assign w3451 = ~w2280 & w3450;
assign w3452 = ~w3449 & ~w3451;
assign w3453 = ~w3448 & w3452;
assign w3454 = ~w2773 & w4166;
assign w3455 = ~w2751 & w3454;
assign w3456 = ~w2601 & w2750;
assign w3457 = ~w2280 & w3456;
assign w3458 = (~w2601 & w2773) | (~w2601 & w4167) | (w2773 & w4167);
assign w3459 = ~w3457 & ~w3458;
assign w3460 = ~w3455 & w3459;
assign w3461 = ~w2773 & w4168;
assign w3462 = ~w2751 & w3461;
assign w3463 = (w2584 & w2773) | (w2584 & w4169) | (w2773 & w4169);
assign w3464 = w2584 & w2750;
assign w3465 = ~w2280 & w3464;
assign w3466 = ~w3463 & ~w3465;
assign w3467 = ~w3462 & w3466;
assign w3468 = ~w2773 & w4170;
assign w3469 = ~w2751 & w3468;
assign w3470 = ~w2577 & w2750;
assign w3471 = ~w2280 & w3470;
assign w3472 = (~w2577 & w2773) | (~w2577 & w4171) | (w2773 & w4171);
assign w3473 = ~w3471 & ~w3472;
assign w3474 = ~w3469 & w3473;
assign w3475 = ~w2773 & w4172;
assign w3476 = ~w2751 & w3475;
assign w3477 = ~w2569 & w2750;
assign w3478 = ~w2280 & w3477;
assign w3479 = (~w2569 & w2773) | (~w2569 & w4173) | (w2773 & w4173);
assign w3480 = ~w3478 & ~w3479;
assign w3481 = ~w3476 & w3480;
assign w3482 = ~w2773 & w4174;
assign w3483 = ~w2751 & w3482;
assign w3484 = ~w2560 & w2750;
assign w3485 = ~w2280 & w3484;
assign w3486 = (~w2560 & w2773) | (~w2560 & w4175) | (w2773 & w4175);
assign w3487 = ~w3485 & ~w3486;
assign w3488 = ~w3483 & w3487;
assign w3489 = ~w2773 & w4176;
assign w3490 = ~w2751 & w3489;
assign w3491 = (w2544 & w2773) | (w2544 & w4177) | (w2773 & w4177);
assign w3492 = w2544 & w2750;
assign w3493 = ~w2280 & w3492;
assign w3494 = ~w3491 & ~w3493;
assign w3495 = ~w3490 & w3494;
assign w3496 = ~w2773 & w4178;
assign w3497 = ~w2751 & w3496;
assign w3498 = ~w2538 & w2750;
assign w3499 = ~w2280 & w3498;
assign w3500 = (~w2538 & w2773) | (~w2538 & w4179) | (w2773 & w4179);
assign w3501 = ~w3499 & ~w3500;
assign w3502 = ~w3497 & w3501;
assign w3503 = ~w2773 & w4180;
assign w3504 = ~w2751 & w3503;
assign w3505 = (w2656 & w2773) | (w2656 & w4181) | (w2773 & w4181);
assign w3506 = w2656 & w2750;
assign w3507 = ~w2280 & w3506;
assign w3508 = ~w3505 & ~w3507;
assign w3509 = ~w3504 & w3508;
assign w3510 = ~w2773 & w4182;
assign w3511 = ~w2751 & w3510;
assign w3512 = ~w2650 & w2750;
assign w3513 = ~w2280 & w3512;
assign w3514 = (~w2650 & w2773) | (~w2650 & w4183) | (w2773 & w4183);
assign w3515 = ~w3513 & ~w3514;
assign w3516 = ~w3511 & w3515;
assign w3517 = ~w2773 & w4184;
assign w3518 = ~w2751 & w3517;
assign w3519 = (w2633 & w2773) | (w2633 & w4185) | (w2773 & w4185);
assign w3520 = w2633 & w2750;
assign w3521 = ~w2280 & w3520;
assign w3522 = ~w3519 & ~w3521;
assign w3523 = ~w3518 & w3522;
assign w3524 = ~w2773 & w4186;
assign w3525 = ~w2751 & w3524;
assign w3526 = ~w2626 & w2750;
assign w3527 = ~w2280 & w3526;
assign w3528 = (~w2626 & w2773) | (~w2626 & w4187) | (w2773 & w4187);
assign w3529 = ~w3527 & ~w3528;
assign w3530 = ~w3525 & w3529;
assign w3531 = ~w2773 & w4188;
assign w3532 = ~w2751 & w3531;
assign w3533 = ~w2462 & w2750;
assign w3534 = ~w2280 & w3533;
assign w3535 = (~w2462 & w2773) | (~w2462 & w4189) | (w2773 & w4189);
assign w3536 = ~w3534 & ~w3535;
assign w3537 = ~w3532 & w3536;
assign w3538 = ~w2773 & w4190;
assign w3539 = ~w2751 & w3538;
assign w3540 = ~w2438 & w2750;
assign w3541 = ~w2280 & w3540;
assign w3542 = (~w2438 & w2773) | (~w2438 & w4191) | (w2773 & w4191);
assign w3543 = ~w3541 & ~w3542;
assign w3544 = ~w3539 & w3543;
assign w3545 = ~w2773 & w4192;
assign w3546 = ~w2751 & w3545;
assign w3547 = (w2444 & w2773) | (w2444 & w4193) | (w2773 & w4193);
assign w3548 = w2444 & w2750;
assign w3549 = ~w2280 & w3548;
assign w3550 = ~w3547 & ~w3549;
assign w3551 = ~w3546 & w3550;
assign w3552 = ~w2773 & w4194;
assign w3553 = ~w2751 & w3552;
assign w3554 = ~w2472 & w2750;
assign w3555 = ~w2280 & w3554;
assign w3556 = (~w2472 & w2773) | (~w2472 & w4195) | (w2773 & w4195);
assign w3557 = ~w3555 & ~w3556;
assign w3558 = ~w3553 & w3557;
assign w3559 = ~w2773 & w4196;
assign w3560 = ~w2751 & w3559;
assign w3561 = (w2418 & w2773) | (w2418 & w4197) | (w2773 & w4197);
assign w3562 = w2418 & w2750;
assign w3563 = ~w2280 & w3562;
assign w3564 = ~w3561 & ~w3563;
assign w3565 = ~w3560 & w3564;
assign w3566 = ~w2773 & w4198;
assign w3567 = ~w2751 & w3566;
assign w3568 = ~w2414 & w2750;
assign w3569 = ~w2280 & w3568;
assign w3570 = (~w2414 & w2773) | (~w2414 & w4199) | (w2773 & w4199);
assign w3571 = ~w3569 & ~w3570;
assign w3572 = ~w3567 & w3571;
assign w3573 = ~w2773 & w4200;
assign w3574 = ~w2751 & w3573;
assign w3575 = (w2401 & w2773) | (w2401 & w4201) | (w2773 & w4201);
assign w3576 = w2401 & w2750;
assign w3577 = ~w2280 & w3576;
assign w3578 = ~w3575 & ~w3577;
assign w3579 = ~w3574 & w3578;
assign w3580 = ~w2773 & w4202;
assign w3581 = ~w2751 & w3580;
assign w3582 = ~w2394 & w2750;
assign w3583 = ~w2280 & w3582;
assign w3584 = (~w2394 & w2773) | (~w2394 & w4203) | (w2773 & w4203);
assign w3585 = ~w3583 & ~w3584;
assign w3586 = ~w3581 & w3585;
assign w3587 = ~w2773 & w4204;
assign w3588 = ~w2751 & w3587;
assign w3589 = ~w2317 & w2750;
assign w3590 = ~w2280 & w3589;
assign w3591 = (~w2317 & w2773) | (~w2317 & w4205) | (w2773 & w4205);
assign w3592 = ~w3590 & ~w3591;
assign w3593 = ~w3588 & w3592;
assign w3594 = ~w2773 & w4206;
assign w3595 = ~w2751 & w3594;
assign w3596 = ~w2308 & w2750;
assign w3597 = ~w2280 & w3596;
assign w3598 = (~w2308 & w2773) | (~w2308 & w4207) | (w2773 & w4207);
assign w3599 = ~w3597 & ~w3598;
assign w3600 = ~w3595 & w3599;
assign w3601 = ~w2773 & w4208;
assign w3602 = ~w2751 & w3601;
assign w3603 = (w2292 & w2773) | (w2292 & w4209) | (w2773 & w4209);
assign w3604 = w2292 & w2750;
assign w3605 = ~w2280 & w3604;
assign w3606 = ~w3603 & ~w3605;
assign w3607 = ~w3602 & w3606;
assign w3608 = ~w2773 & w4210;
assign w3609 = ~w2751 & w3608;
assign w3610 = ~w2286 & w2750;
assign w3611 = ~w2280 & w3610;
assign w3612 = (~w2286 & w2773) | (~w2286 & w4211) | (w2773 & w4211);
assign w3613 = ~w3611 & ~w3612;
assign w3614 = ~w3609 & w3613;
assign w3615 = ~w2773 & w4212;
assign w3616 = ~w2751 & w3615;
assign w3617 = (w2377 & w2773) | (w2377 & w4213) | (w2773 & w4213);
assign w3618 = w2377 & w2750;
assign w3619 = ~w2280 & w3618;
assign w3620 = ~w3617 & ~w3619;
assign w3621 = ~w3616 & w3620;
assign w3622 = ~w2773 & w4214;
assign w3623 = ~w2751 & w3622;
assign w3624 = ~w2373 & w2750;
assign w3625 = ~w2280 & w3624;
assign w3626 = (~w2373 & w2773) | (~w2373 & w4215) | (w2773 & w4215);
assign w3627 = ~w3625 & ~w3626;
assign w3628 = ~w3623 & w3627;
assign w3629 = ~w2773 & w4216;
assign w3630 = ~w2751 & w3629;
assign w3631 = (w2361 & w2773) | (w2361 & w4217) | (w2773 & w4217);
assign w3632 = w2361 & w2750;
assign w3633 = ~w2280 & w3632;
assign w3634 = ~w3631 & ~w3633;
assign w3635 = ~w3630 & w3634;
assign w3636 = ~w2773 & w4218;
assign w3637 = ~w2751 & w3636;
assign w3638 = ~w2357 & w2750;
assign w3639 = ~w2280 & w3638;
assign w3640 = (~w2357 & w2773) | (~w2357 & w4219) | (w2773 & w4219);
assign w3641 = ~w3639 & ~w3640;
assign w3642 = ~w3637 & w3641;
assign w3643 = ~w2773 & w4220;
assign w3644 = ~w2751 & w3643;
assign w3645 = ~w2349 & w2750;
assign w3646 = ~w2280 & w3645;
assign w3647 = (~w2349 & w2773) | (~w2349 & w4221) | (w2773 & w4221);
assign w3648 = ~w3646 & ~w3647;
assign w3649 = ~w3644 & w3648;
assign w3650 = ~w2773 & w4222;
assign w3651 = ~w2751 & w3650;
assign w3652 = ~w2341 & w2750;
assign w3653 = ~w2280 & w3652;
assign w3654 = (~w2341 & w2773) | (~w2341 & w4223) | (w2773 & w4223);
assign w3655 = ~w3653 & ~w3654;
assign w3656 = ~w3651 & w3655;
assign w3657 = ~w2773 & w4224;
assign w3658 = ~w2751 & w3657;
assign w3659 = (~w2772 & w5303) | (~w2772 & w5304) | (w5303 & w5304);
assign w3660 = w2749 & w5305;
assign w3661 = (~w3659 & w2280) | (~w3659 & w5306) | (w2280 & w5306);
assign w3662 = ~w3658 & w3661;
assign w3663 = w2499 & w2501;
assign w3664 = ~w2773 & w4226;
assign w3665 = ~w2751 & w3664;
assign w3666 = (~w1189 & w2773) | (~w1189 & w4227) | (w2773 & w4227);
assign w3667 = ~w1189 & w2750;
assign w3668 = ~w2280 & w3667;
assign w3669 = ~w3666 & ~w3668;
assign w3670 = ~w3665 & w3669;
assign w3671 = ~w2751 & w2774;
assign w3672 = ~w39 & w51;
assign w3673 = ~w170 & w175;
assign w3674 = w201 & w181;
assign w3675 = ~w361 & ~w358;
assign w3676 = ~w375 & ~w372;
assign w3677 = ~w447 & w454;
assign w3678 = ~w451 & ~w470;
assign w3679 = ~w490 & ~w487;
assign w3680 = ~w393 & w4228;
assign w3681 = (~w537 & w5307) | (~w537 & w5308) | (w5307 & w5308);
assign w3682 = (~w537 & w6265) | (~w537 & w6266) | (w6265 & w6266);
assign w3683 = ~w618 & w630;
assign w3684 = ~w749 & w754;
assign w3685 = w780 & w760;
assign w3686 = ~w940 & ~w937;
assign w3687 = ~w954 & ~w951;
assign w3688 = ~w1026 & w1033;
assign w3689 = ~w1030 & ~w1049;
assign w3690 = ~w1069 & ~w1066;
assign w3691 = ~w972 & w4229;
assign w3692 = (~w1123 & w5309) | (~w1123 & w5310) | (w5309 & w5310);
assign w3693 = (~w1123 & w6267) | (~w1123 & w6268) | (w6267 & w6268);
assign w3694 = (~w1123 & w5311) | (~w1123 & w5312) | (w5311 & w5312);
assign w3695 = (~w1123 & w6269) | (~w1123 & w6270) | (w6269 & w6270);
assign w3696 = (~w537 & w5313) | (~w537 & w5314) | (w5313 & w5314);
assign w3697 = (~w537 & w6271) | (~w537 & w6272) | (w6271 & w6272);
assign w3698 = (~w537 & w5315) | (~w537 & w5316) | (w5315 & w5316);
assign w3699 = (~w537 & w6273) | (~w537 & w6274) | (w6273 & w6274);
assign w3700 = (~w1123 & w5317) | (~w1123 & w5318) | (w5317 & w5318);
assign w3701 = (~w1123 & w6275) | (~w1123 & w6276) | (w6275 & w6276);
assign w3702 = (~w537 & w5319) | (~w537 & w5320) | (w5319 & w5320);
assign w3703 = (~w1123 & w5321) | (~w1123 & w5322) | (w5321 & w5322);
assign w3704 = (~w537 & w5323) | (~w537 & w5324) | (w5323 & w5324);
assign w3705 = (~w537 & w6277) | (~w537 & w6278) | (w6277 & w6278);
assign w3706 = (~w1123 & w5325) | (~w1123 & w5326) | (w5325 & w5326);
assign w3707 = (~w1123 & w6279) | (~w1123 & w6280) | (w6279 & w6280);
assign w3708 = (~w537 & w5327) | (~w537 & w5328) | (w5327 & w5328);
assign w3709 = (~w537 & w6281) | (~w537 & w6282) | (w6281 & w6282);
assign w3710 = (~w1123 & w5329) | (~w1123 & w5330) | (w5329 & w5330);
assign w3711 = (~w1123 & w6283) | (~w1123 & w6284) | (w6283 & w6284);
assign w3712 = (~w537 & w5331) | (~w537 & w5332) | (w5331 & w5332);
assign w3713 = (~w537 & w6285) | (~w537 & w6286) | (w6285 & w6286);
assign w3714 = (~w1123 & w5333) | (~w1123 & w5334) | (w5333 & w5334);
assign w3715 = (~w1123 & w6287) | (~w1123 & w6288) | (w6287 & w6288);
assign w3716 = (~w537 & w5335) | (~w537 & w5336) | (w5335 & w5336);
assign w3717 = (~w537 & w6289) | (~w537 & w6290) | (w6289 & w6290);
assign w3718 = (~w1123 & w5337) | (~w1123 & w5338) | (w5337 & w5338);
assign w3719 = (~w1123 & w6291) | (~w1123 & w6292) | (w6291 & w6292);
assign w3720 = (~w537 & w5339) | (~w537 & w5340) | (w5339 & w5340);
assign w3721 = (~w537 & w6293) | (~w537 & w6294) | (w6293 & w6294);
assign w3722 = (~w1123 & w5341) | (~w1123 & w5342) | (w5341 & w5342);
assign w3723 = (~w1123 & w6295) | (~w1123 & w6296) | (w6295 & w6296);
assign w3724 = (~w537 & w5343) | (~w537 & w5344) | (w5343 & w5344);
assign w3725 = (~w537 & w6297) | (~w537 & w6298) | (w6297 & w6298);
assign w3726 = (~w1123 & w5345) | (~w1123 & w5346) | (w5345 & w5346);
assign w3727 = (~w1123 & w6299) | (~w1123 & w6300) | (w6299 & w6300);
assign w3728 = (~w537 & w5347) | (~w537 & w5348) | (w5347 & w5348);
assign w3729 = (~w537 & w6301) | (~w537 & w6302) | (w6301 & w6302);
assign w3730 = (~w1123 & w5349) | (~w1123 & w5350) | (w5349 & w5350);
assign w3731 = (~w1123 & w6303) | (~w1123 & w6304) | (w6303 & w6304);
assign w3732 = (~w537 & w5351) | (~w537 & w5352) | (w5351 & w5352);
assign w3733 = (~w537 & w6305) | (~w537 & w6306) | (w6305 & w6306);
assign w3734 = (~w1123 & w5353) | (~w1123 & w5354) | (w5353 & w5354);
assign w3735 = (~w1123 & w6307) | (~w1123 & w6308) | (w6307 & w6308);
assign w3736 = (~w1123 & w5355) | (~w1123 & w5356) | (w5355 & w5356);
assign w3737 = (~w1123 & w6309) | (~w1123 & w6310) | (w6309 & w6310);
assign w3738 = (~w537 & w5357) | (~w537 & w5358) | (w5357 & w5358);
assign w3739 = (~w537 & w6311) | (~w537 & w6312) | (w6311 & w6312);
assign w3740 = (~w537 & w5359) | (~w537 & w5360) | (w5359 & w5360);
assign w3741 = (~w537 & w6313) | (~w537 & w6314) | (w6313 & w6314);
assign w3742 = (~w1123 & w5361) | (~w1123 & w5362) | (w5361 & w5362);
assign w3743 = (~w1123 & w6315) | (~w1123 & w6316) | (w6315 & w6316);
assign w3744 = (~w537 & w5363) | (~w537 & w5364) | (w5363 & w5364);
assign w3745 = (~w537 & w6317) | (~w537 & w6318) | (w6317 & w6318);
assign w3746 = (~w1123 & w5365) | (~w1123 & w5366) | (w5365 & w5366);
assign w3747 = (~w1123 & w6319) | (~w1123 & w6320) | (w6319 & w6320);
assign w3748 = (~w537 & w5367) | (~w537 & w5368) | (w5367 & w5368);
assign w3749 = (~w537 & w6321) | (~w537 & w6322) | (w6321 & w6322);
assign w3750 = (~w1123 & w5369) | (~w1123 & w5370) | (w5369 & w5370);
assign w3751 = (~w1123 & w6323) | (~w1123 & w6324) | (w6323 & w6324);
assign w3752 = (~w537 & w5371) | (~w537 & w5372) | (w5371 & w5372);
assign w3753 = (~w537 & w6325) | (~w537 & w6326) | (w6325 & w6326);
assign w3754 = (~w1123 & w5373) | (~w1123 & w5374) | (w5373 & w5374);
assign w3755 = (~w1123 & w6327) | (~w1123 & w6328) | (w6327 & w6328);
assign w3756 = (~w537 & w5375) | (~w537 & w5376) | (w5375 & w5376);
assign w3757 = (~w537 & w6329) | (~w537 & w6330) | (w6329 & w6330);
assign w3758 = (~w1123 & w5377) | (~w1123 & w5378) | (w5377 & w5378);
assign w3759 = (~w1123 & w6331) | (~w1123 & w6332) | (w6331 & w6332);
assign w3760 = (~w537 & w5379) | (~w537 & w5380) | (w5379 & w5380);
assign w3761 = (~w537 & w6333) | (~w537 & w6334) | (w6333 & w6334);
assign w3762 = (~w1123 & w5381) | (~w1123 & w5382) | (w5381 & w5382);
assign w3763 = (~w1123 & w6335) | (~w1123 & w6336) | (w6335 & w6336);
assign w3764 = (~w1123 & w5383) | (~w1123 & w5384) | (w5383 & w5384);
assign w3765 = (~w1123 & w6337) | (~w1123 & w6338) | (w6337 & w6338);
assign w3766 = (~w537 & w5385) | (~w537 & w5386) | (w5385 & w5386);
assign w3767 = (~w537 & w6339) | (~w537 & w6340) | (w6339 & w6340);
assign w3768 = (~w1123 & w5387) | (~w1123 & w5388) | (w5387 & w5388);
assign w3769 = (~w1123 & w6341) | (~w1123 & w6342) | (w6341 & w6342);
assign w3770 = (~w537 & w5389) | (~w537 & w5390) | (w5389 & w5390);
assign w3771 = (~w537 & w6343) | (~w537 & w6344) | (w6343 & w6344);
assign w3772 = (~w537 & w5391) | (~w537 & w5392) | (w5391 & w5392);
assign w3773 = (~w537 & w6345) | (~w537 & w6346) | (w6345 & w6346);
assign w3774 = (~w1123 & w5393) | (~w1123 & w5394) | (w5393 & w5394);
assign w3775 = (~w1123 & w6347) | (~w1123 & w6348) | (w6347 & w6348);
assign w3776 = (~w1123 & w5395) | (~w1123 & w5396) | (w5395 & w5396);
assign w3777 = (~w1123 & w6349) | (~w1123 & w6350) | (w6349 & w6350);
assign w3778 = (~w537 & w5397) | (~w537 & w5398) | (w5397 & w5398);
assign w3779 = (~w537 & w6351) | (~w537 & w6352) | (w6351 & w6352);
assign w3780 = (~w537 & w5399) | (~w537 & w5400) | (w5399 & w5400);
assign w3781 = ~w1697 & w7149;
assign w3782 = (~w1123 & w5401) | (~w1123 & w5402) | (w5401 & w5402);
assign w3783 = ~w1702 & w7150;
assign w3784 = (~w1123 & w5403) | (~w1123 & w5404) | (w5403 & w5404);
assign w3785 = ~w1709 & w7151;
assign w3786 = (~w537 & w5405) | (~w537 & w5406) | (w5405 & w5406);
assign w3787 = ~w1714 & w7152;
assign w3788 = (~w537 & w5407) | (~w537 & w5408) | (w5407 & w5408);
assign w3789 = ~w1722 & w7153;
assign w3790 = (~w1123 & w5409) | (~w1123 & w5410) | (w5409 & w5410);
assign w3791 = ~w1727 & w7154;
assign w3792 = (~w537 & w5411) | (~w537 & w5412) | (w5411 & w5412);
assign w3793 = ~w1733 & w7155;
assign w3794 = (~w1123 & w5413) | (~w1123 & w5414) | (w5413 & w5414);
assign w3795 = ~w1738 & w7156;
assign w3796 = (~w537 & w5415) | (~w537 & w5416) | (w5415 & w5416);
assign w3797 = ~w1746 & w7157;
assign w3798 = (~w1123 & w5417) | (~w1123 & w5418) | (w5417 & w5418);
assign w3799 = ~w1751 & w7158;
assign w3800 = (~w537 & w5419) | (~w537 & w5420) | (w5419 & w5420);
assign w3801 = ~w1760 & w7159;
assign w3802 = (~w1123 & w5421) | (~w1123 & w5422) | (w5421 & w5422);
assign w3803 = ~w1765 & w7160;
assign w3804 = (~w1123 & w5423) | (~w1123 & w5424) | (w5423 & w5424);
assign w3805 = ~w1771 & w7161;
assign w3806 = (~w537 & w5425) | (~w537 & w5426) | (w5425 & w5426);
assign w3807 = ~w1776 & w7162;
assign w3808 = (~w1123 & w5427) | (~w1123 & w5428) | (w5427 & w5428);
assign w3809 = ~w1784 & w7163;
assign w3810 = (~w537 & w5429) | (~w537 & w5430) | (w5429 & w5430);
assign w3811 = ~w1789 & w7164;
assign w3812 = (~w537 & w5431) | (~w537 & w5432) | (w5431 & w5432);
assign w3813 = (~w537 & w6353) | (~w537 & w6354) | (w6353 & w6354);
assign w3814 = (~w1123 & w5433) | (~w1123 & w5434) | (w5433 & w5434);
assign w3815 = (~w1123 & w6355) | (~w1123 & w6356) | (w6355 & w6356);
assign w3816 = (~w537 & w5435) | (~w537 & w5436) | (w5435 & w5436);
assign w3817 = (~w537 & w6357) | (~w537 & w6358) | (w6357 & w6358);
assign w3818 = (~w1123 & w5437) | (~w1123 & w5438) | (w5437 & w5438);
assign w3819 = (~w1123 & w6359) | (~w1123 & w6360) | (w6359 & w6360);
assign w3820 = (~w537 & w5439) | (~w537 & w5440) | (w5439 & w5440);
assign w3821 = (~w537 & w6361) | (~w537 & w6362) | (w6361 & w6362);
assign w3822 = (~w1123 & w5441) | (~w1123 & w5442) | (w5441 & w5442);
assign w3823 = (~w1123 & w6363) | (~w1123 & w6364) | (w6363 & w6364);
assign w3824 = (~w537 & w5443) | (~w537 & w5444) | (w5443 & w5444);
assign w3825 = (~w537 & w6365) | (~w537 & w6366) | (w6365 & w6366);
assign w3826 = (~w1123 & w5445) | (~w1123 & w5446) | (w5445 & w5446);
assign w3827 = (~w1123 & w6367) | (~w1123 & w6368) | (w6367 & w6368);
assign w3828 = (~w537 & w5587) | (~w537 & w5588) | (w5587 & w5588);
assign w3829 = (~w537 & w6369) | (~w537 & w6370) | (w6369 & w6370);
assign w3830 = (~w1123 & w5589) | (~w1123 & w5590) | (w5589 & w5590);
assign w3831 = (~w1123 & w6371) | (~w1123 & w6372) | (w6371 & w6372);
assign w3832 = (~w537 & w5591) | (~w537 & w5592) | (w5591 & w5592);
assign w3833 = (~w537 & w6373) | (~w537 & w6374) | (w6373 & w6374);
assign w3834 = (~w1123 & w5593) | (~w1123 & w5594) | (w5593 & w5594);
assign w3835 = (~w1123 & w6375) | (~w1123 & w6376) | (w6375 & w6376);
assign w3836 = (~w1123 & w5595) | (~w1123 & w5596) | (w5595 & w5596);
assign w3837 = ~w1953 & w7165;
assign w3838 = (~w537 & w5597) | (~w537 & w5598) | (w5597 & w5598);
assign w3839 = ~w1958 & w7166;
assign w3840 = (~w537 & w5599) | (~w537 & w5600) | (w5599 & w5600);
assign w3841 = (~w537 & w6377) | (~w537 & w6378) | (w6377 & w6378);
assign w3842 = (~w1123 & w5601) | (~w1123 & w5602) | (w5601 & w5602);
assign w3843 = (~w1123 & w6379) | (~w1123 & w6380) | (w6379 & w6380);
assign w3844 = (~w1123 & w5603) | (~w1123 & w5604) | (w5603 & w5604);
assign w3845 = (~w1123 & w6381) | (~w1123 & w6382) | (w6381 & w6382);
assign w3846 = (~w537 & w5605) | (~w537 & w5606) | (w5605 & w5606);
assign w3847 = (~w537 & w6383) | (~w537 & w6384) | (w6383 & w6384);
assign w3848 = (~w537 & w5607) | (~w537 & w5608) | (w5607 & w5608);
assign w3849 = (~w537 & w6385) | (~w537 & w6386) | (w6385 & w6386);
assign w3850 = (~w1123 & w5609) | (~w1123 & w5610) | (w5609 & w5610);
assign w3851 = (~w1123 & w6387) | (~w1123 & w6388) | (w6387 & w6388);
assign w3852 = (~w1123 & w5611) | (~w1123 & w5612) | (w5611 & w5612);
assign w3853 = (~w1123 & w6389) | (~w1123 & w6390) | (w6389 & w6390);
assign w3854 = (~w537 & w5613) | (~w537 & w5614) | (w5613 & w5614);
assign w3855 = (~w537 & w6391) | (~w537 & w6392) | (w6391 & w6392);
assign w3856 = (~w537 & w5615) | (~w537 & w5616) | (w5615 & w5616);
assign w3857 = (~w537 & w6393) | (~w537 & w6394) | (w6393 & w6394);
assign w3858 = (~w1123 & w5617) | (~w1123 & w5618) | (w5617 & w5618);
assign w3859 = (~w1123 & w6395) | (~w1123 & w6396) | (w6395 & w6396);
assign w3860 = (~w1123 & w5619) | (~w1123 & w5620) | (w5619 & w5620);
assign w3861 = (~w1123 & w6397) | (~w1123 & w6398) | (w6397 & w6398);
assign w3862 = (~w537 & w5621) | (~w537 & w5622) | (w5621 & w5622);
assign w3863 = (~w537 & w6399) | (~w537 & w6400) | (w6399 & w6400);
assign w3864 = (~w1123 & w5623) | (~w1123 & w5624) | (w5623 & w5624);
assign w3865 = (~w1123 & w6401) | (~w1123 & w6402) | (w6401 & w6402);
assign w3866 = (~w537 & w5625) | (~w537 & w5626) | (w5625 & w5626);
assign w3867 = (~w537 & w6403) | (~w537 & w6404) | (w6403 & w6404);
assign w3868 = (~w537 & w5627) | (~w537 & w5628) | (w5627 & w5628);
assign w3869 = (~w537 & w6405) | (~w537 & w6406) | (w6405 & w6406);
assign w3870 = (~w1123 & w5629) | (~w1123 & w5630) | (w5629 & w5630);
assign w3871 = (~w1123 & w6407) | (~w1123 & w6408) | (w6407 & w6408);
assign w3872 = (~w537 & w5631) | (~w537 & w5632) | (w5631 & w5632);
assign w3873 = (~w537 & w6409) | (~w537 & w6410) | (w6409 & w6410);
assign w3874 = (~w1123 & w5633) | (~w1123 & w5634) | (w5633 & w5634);
assign w3875 = (~w1123 & w6411) | (~w1123 & w6412) | (w6411 & w6412);
assign w3876 = (~w537 & w5635) | (~w537 & w5636) | (w5635 & w5636);
assign w3877 = ~w2199 & w7167;
assign w3878 = (~w1123 & w5637) | (~w1123 & w5638) | (w5637 & w5638);
assign w3879 = ~w2204 & w7168;
assign w3880 = (~w1123 & w5639) | (~w1123 & w5640) | (w5639 & w5640);
assign w3881 = ~w2211 & w7169;
assign w3882 = (~w537 & w5641) | (~w537 & w5642) | (w5641 & w5642);
assign w3883 = ~w2216 & w7170;
assign w3884 = (~w537 & w5643) | (~w537 & w5644) | (w5643 & w5644);
assign w3885 = ~w2222 & w7171;
assign w3886 = (~w1123 & w5645) | (~w1123 & w5646) | (w5645 & w5646);
assign w3887 = ~w2227 & w7172;
assign w3888 = (~w537 & w5647) | (~w537 & w5648) | (w5647 & w5648);
assign w3889 = ~w2240 & w7173;
assign w3890 = (~w1123 & w5649) | (~w1123 & w5650) | (w5649 & w5650);
assign w3891 = ~w2245 & w7174;
assign w3892 = (~w537 & w5651) | (~w537 & w5652) | (w5651 & w5652);
assign w3893 = ~w2251 & w7175;
assign w3894 = (~w1123 & w5653) | (~w1123 & w5654) | (w5653 & w5654);
assign w3895 = ~w2256 & w7176;
assign w3896 = (~w1123 & w5655) | (~w1123 & w5656) | (w5655 & w5656);
assign w3897 = ~w2262 & w7177;
assign w3898 = (~w537 & w5657) | (~w537 & w5658) | (w5657 & w5658);
assign w3899 = ~w2267 & w7178;
assign w3900 = (~w1123 & w5659) | (~w1123 & w5660) | (w5659 & w5660);
assign w3901 = ~w2290 & w7179;
assign w3902 = (~w537 & w5661) | (~w537 & w5662) | (w5661 & w5662);
assign w3903 = ~w2295 & w7180;
assign w3904 = (~w537 & w5663) | (~w537 & w5664) | (w5663 & w5664);
assign w3905 = ~w2301 & w7181;
assign w3906 = (~w1123 & w5665) | (~w1123 & w5666) | (w5665 & w5666);
assign w3907 = ~w2306 & w7182;
assign w3908 = (~w537 & w5667) | (~w537 & w5668) | (w5667 & w5668);
assign w3909 = (~w537 & w6413) | (~w537 & w6414) | (w6413 & w6414);
assign w3910 = (~w1123 & w5669) | (~w1123 & w5670) | (w5669 & w5670);
assign w3911 = (~w1123 & w6415) | (~w1123 & w6416) | (w6415 & w6416);
assign w3912 = (~w1123 & w5671) | (~w1123 & w5672) | (w5671 & w5672);
assign w3913 = (~w1123 & w6417) | (~w1123 & w6418) | (w6417 & w6418);
assign w3914 = (~w537 & w5673) | (~w537 & w5674) | (w5673 & w5674);
assign w3915 = (~w537 & w6419) | (~w537 & w6420) | (w6419 & w6420);
assign w3916 = (~w537 & w5675) | (~w537 & w5676) | (w5675 & w5676);
assign w3917 = (~w537 & w6421) | (~w537 & w6422) | (w6421 & w6422);
assign w3918 = (~w1123 & w5677) | (~w1123 & w5678) | (w5677 & w5678);
assign w3919 = (~w1123 & w6423) | (~w1123 & w6424) | (w6423 & w6424);
assign w3920 = (~w1123 & w5679) | (~w1123 & w5680) | (w5679 & w5680);
assign w3921 = (~w1123 & w6425) | (~w1123 & w6426) | (w6425 & w6426);
assign w3922 = (~w537 & w5681) | (~w537 & w5682) | (w5681 & w5682);
assign w3923 = (~w537 & w6427) | (~w537 & w6428) | (w6427 & w6428);
assign w3924 = (~w537 & w5683) | (~w537 & w5684) | (w5683 & w5684);
assign w3925 = (~w537 & w6429) | (~w537 & w6430) | (w6429 & w6430);
assign w3926 = (~w1123 & w5685) | (~w1123 & w5686) | (w5685 & w5686);
assign w3927 = (~w1123 & w6431) | (~w1123 & w6432) | (w6431 & w6432);
assign w3928 = (~w1123 & w5687) | (~w1123 & w5688) | (w5687 & w5688);
assign w3929 = (~w1123 & w6433) | (~w1123 & w6434) | (w6433 & w6434);
assign w3930 = (~w537 & w5689) | (~w537 & w5690) | (w5689 & w5690);
assign w3931 = (~w537 & w6435) | (~w537 & w6436) | (w6435 & w6436);
assign w3932 = (~w537 & w5691) | (~w537 & w5692) | (w5691 & w5692);
assign w3933 = (~w537 & w6437) | (~w537 & w6438) | (w6437 & w6438);
assign w3934 = (~w1123 & w5693) | (~w1123 & w5694) | (w5693 & w5694);
assign w3935 = (~w1123 & w6439) | (~w1123 & w6440) | (w6439 & w6440);
assign w3936 = (~w1123 & w5695) | (~w1123 & w5696) | (w5695 & w5696);
assign w3937 = ~w2582 & w7183;
assign w3938 = (~w537 & w5697) | (~w537 & w5698) | (w5697 & w5698);
assign w3939 = ~w2587 & w7184;
assign w3940 = (~w537 & w5699) | (~w537 & w5700) | (w5699 & w5700);
assign w3941 = ~w2594 & w7185;
assign w3942 = (~w1123 & w5701) | (~w1123 & w5702) | (w5701 & w5702);
assign w3943 = ~w2599 & w7186;
assign w3944 = (~w1123 & w5703) | (~w1123 & w5704) | (w5703 & w5704);
assign w3945 = ~w2605 & w7187;
assign w3946 = (~w537 & w5705) | (~w537 & w5706) | (w5705 & w5706);
assign w3947 = ~w2610 & w7188;
assign w3948 = (~w1123 & w5707) | (~w1123 & w5708) | (w5707 & w5708);
assign w3949 = ~w2631 & w7189;
assign w3950 = (~w537 & w5709) | (~w537 & w5710) | (w5709 & w5710);
assign w3951 = ~w2636 & w7190;
assign w3952 = (~w537 & w5711) | (~w537 & w5712) | (w5711 & w5712);
assign w3953 = ~w2643 & w7191;
assign w3954 = (~w1123 & w5713) | (~w1123 & w5714) | (w5713 & w5714);
assign w3955 = ~w2648 & w7192;
assign w3956 = (~w1123 & w5715) | (~w1123 & w5716) | (w5715 & w5716);
assign w3957 = ~w2654 & w7193;
assign w3958 = (~w537 & w5717) | (~w537 & w5718) | (w5717 & w5718);
assign w3959 = ~w2659 & w7194;
assign w3960 = (~w537 & w5719) | (~w537 & w5720) | (w5719 & w5720);
assign w3961 = ~w2699 & w7195;
assign w3962 = (~w1123 & w5721) | (~w1123 & w5722) | (w5721 & w5722);
assign w3963 = ~w2704 & w7196;
assign w3964 = (~w537 & w5723) | (~w537 & w5724) | (w5723 & w5724);
assign w3965 = ~w2710 & w7197;
assign w3966 = (~w1123 & w5725) | (~w1123 & w5726) | (w5725 & w5726);
assign w3967 = ~w2715 & w7198;
assign w3968 = (~w1123 & w5727) | (~w1123 & w5728) | (w5727 & w5728);
assign w3969 = ~w2723 & w7199;
assign w3970 = (~w537 & w5729) | (~w537 & w5730) | (w5729 & w5730);
assign w3971 = ~w2728 & w7200;
assign w3972 = ~w2752 & ~w578;
assign w3973 = w2752 & ~w1157;
assign w3974 = ~w2752 & w1168;
assign w3975 = w2752 & w1163;
assign w3976 = ~w2752 & ~w1176;
assign w3977 = w2752 & ~w1181;
assign w3978 = ~w2752 & ~w1188;
assign w3979 = w2752 & ~w1192;
assign w3980 = ~w2752 & ~w1198;
assign w3981 = w2752 & ~w1203;
assign w3982 = ~w2752 & ~w1211;
assign w3983 = w2752 & ~w1214;
assign w3984 = ~w2752 & ~w1220;
assign w3985 = w2752 & ~w1225;
assign w3986 = ~w2752 & ~w1337;
assign w3987 = w2752 & ~w1342;
assign w3988 = ~w2752 & ~w1318;
assign w3989 = w2752 & ~w1313;
assign w3990 = ~w2752 & ~w1324;
assign w3991 = w2752 & ~w1329;
assign w3992 = ~w2752 & ~w1262;
assign w3993 = w2752 & ~w1267;
assign w3994 = ~w2752 & ~w1238;
assign w3995 = w2752 & ~w1243;
assign w3996 = ~w2752 & ~w1249;
assign w3997 = w2752 & ~w1254;
assign w3998 = ~w2752 & ~w1299;
assign w3999 = w2752 & ~w1304;
assign w4000 = ~w2752 & ~w1275;
assign w4001 = w2752 & ~w1280;
assign w4002 = ~w2752 & ~w1286;
assign w4003 = w2752 & ~w1291;
assign w4004 = ~w2752 & ~w1426;
assign w4005 = w2752 & ~w1429;
assign w4006 = ~w2752 & w1440;
assign w4007 = w2752 & w1435;
assign w4008 = ~w2752 & ~w1376;
assign w4009 = w2752 & ~w1381;
assign w4010 = ~w2752 & ~w1365;
assign w4011 = w2752 & ~w1370;
assign w4012 = ~w2752 & ~w1389;
assign w4013 = w2752 & ~w1394;
assign w4014 = ~w2752 & ~w1400;
assign w4015 = w2752 & ~w1403;
assign w4016 = ~w2752 & ~w1409;
assign w4017 = w2752 & ~w1414;
assign w4018 = ~w2752 & ~w1526;
assign w4019 = w2752 & ~w1529;
assign w4020 = ~w2752 & ~w1510;
assign w4021 = w2752 & ~w1513;
assign w4022 = ~w2752 & ~w1517;
assign w4023 = w2752 & ~w1520;
assign w4024 = ~w2752 & ~w1475;
assign w4025 = w2752 & ~w1478;
assign w4026 = ~w2752 & ~w1459;
assign w4027 = w2752 & ~w1462;
assign w4028 = ~w2752 & ~w1466;
assign w4029 = w2752 & ~w1469;
assign w4030 = ~w2752 & ~w1500;
assign w4031 = w2752 & ~w1503;
assign w4032 = ~w2752 & ~w1484;
assign w4033 = w2752 & ~w1487;
assign w4034 = ~w2752 & ~w1491;
assign w4035 = w2752 & ~w1494;
assign w4036 = ~w2752 & w1628;
assign w4037 = w2752 & w1623;
assign w4038 = ~w2752 & ~w1634;
assign w4039 = w2752 & ~w1639;
assign w4040 = ~w2752 & w1650;
assign w4041 = w2752 & w1645;
assign w4042 = ~w2752 & ~w1682;
assign w4043 = w2752 & ~w1685;
assign w4044 = ~w2752 & ~w1675;
assign w4045 = w2752 & ~w1678;
assign w4046 = ~w2752 & ~w1660;
assign w4047 = w2752 & ~w1663;
assign w4048 = ~w2752 & w1670;
assign w4049 = w2752 & w1667;
assign w4050 = ~w2752 & ~w1550;
assign w4051 = w2752 & ~w1553;
assign w4052 = ~w2752 & ~w1564;
assign w4053 = w2752 & ~w1567;
assign w4054 = ~w2752 & ~w1571;
assign w4055 = w2752 & ~w1574;
assign w4056 = ~w2752 & ~w1607;
assign w4057 = w2752 & ~w1610;
assign w4058 = ~w2752 & ~w1593;
assign w4059 = w2752 & ~w1596;
assign w4060 = ~w2752 & ~w1600;
assign w4061 = w2752 & ~w1603;
assign w4062 = ~w2752 & ~w1557;
assign w4063 = w2752 & ~w1560;
assign w4064 = ~w2752 & w1581;
assign w4065 = w2752 & w1578;
assign w4066 = ~w2752 & ~w1585;
assign w4067 = w2752 & ~w1588;
assign w4068 = ~w2752 & w1778;
assign w4069 = w2752 & w1773;
assign w4070 = ~w2752 & ~w1762;
assign w4071 = w2752 & ~w1767;
assign w4072 = ~w2752 & w1791;
assign w4073 = w2752 & w1786;
assign w4074 = ~w2752 & ~w1735;
assign w4075 = w2752 & ~w1740;
assign w4076 = ~w2752 & ~w1724;
assign w4077 = w2752 & ~w1729;
assign w4078 = ~w2752 & ~w1748;
assign w4079 = w2752 & ~w1753;
assign w4080 = ~w2752 & w1716;
assign w4081 = w2752 & w1711;
assign w4082 = ~w2752 & ~w1699;
assign w4083 = w2752 & ~w1704;
assign w4084 = ~w2752 & ~w1863;
assign w4085 = w2752 & ~w1868;
assign w4086 = ~w2752 & ~w1852;
assign w4087 = w2752 & ~w1857;
assign w4088 = ~w2752 & ~w1876;
assign w4089 = w2752 & ~w1881;
assign w4090 = ~w2752 & ~w1901;
assign w4091 = w2752 & ~w1906;
assign w4092 = ~w2752 & ~w1890;
assign w4093 = w2752 & ~w1895;
assign w4094 = ~w2752 & ~w1933;
assign w4095 = w2752 & ~w1938;
assign w4096 = ~w2752 & w1916;
assign w4097 = w2752 & w1913;
assign w4098 = ~w2752 & ~w1920;
assign w4099 = w2752 & ~w1923;
assign w4100 = ~w2752 & w1984;
assign w4101 = w2752 & w1979;
assign w4102 = ~w2752 & ~w1968;
assign w4103 = w2752 & ~w1973;
assign w4104 = ~w2752 & w1960;
assign w4105 = w2752 & w1955;
assign w4106 = ~w2752 & ~w1946;
assign w4107 = w2752 & ~w1949;
assign w4108 = ~w2752 & ~w2004;
assign w4109 = w2752 & ~w2007;
assign w4110 = ~w2752 & ~w2013;
assign w4111 = w2752 & ~w2018;
assign w4112 = ~w2752 & w2038;
assign w4113 = w2752 & w2033;
assign w4114 = ~w2752 & ~w2023;
assign w4115 = w2752 & ~w2026;
assign w4116 = ~w2752 & w2218;
assign w4117 = w2752 & w2213;
assign w4118 = ~w2752 & ~w2224;
assign w4119 = w2752 & ~w2229;
assign w4120 = ~w2752 & w2269;
assign w4121 = w2752 & w2264;
assign w4122 = ~w2752 & ~w2242;
assign w4123 = w2752 & ~w2247;
assign w4124 = ~w2752 & ~w2253;
assign w4125 = w2752 & ~w2258;
assign w4126 = ~w2752 & ~w2201;
assign w4127 = w2752 & ~w2206;
assign w4128 = ~w2752 & w2195;
assign w4129 = w2752 & w2192;
assign w4130 = ~w2752 & ~w2233;
assign w4131 = w2752 & ~w2236;
assign w4132 = ~w2752 & w2177;
assign w4133 = w2752 & w2181;
assign w4134 = ~w2752 & ~w2166;
assign w4135 = w2752 & ~w2169;
assign w4136 = ~w2752 & w2069;
assign w4137 = w2752 & w2079;
assign w4138 = ~w2752 & ~w2072;
assign w4139 = w2752 & ~w2075;
assign w4140 = ~w2752 & ~w2157;
assign w4141 = w2752 & ~w2162;
assign w4142 = ~w2752 & ~w2145;
assign w4143 = w2752 & ~w2150;
assign w4144 = ~w2752 & w2139;
assign w4145 = w2752 & w2134;
assign w4146 = ~w2752 & ~w2098;
assign w4147 = w2752 & ~w2101;
assign w4148 = ~w2752 & w2087;
assign w4149 = w2752 & w2084;
assign w4150 = ~w2752 & ~w2091;
assign w4151 = w2752 & ~w2094;
assign w4152 = ~w2752 & w2123;
assign w4153 = w2752 & w2118;
assign w4154 = ~w2752 & ~w2107;
assign w4155 = w2752 & ~w2112;
assign w4156 = ~w2752 & ~w2701;
assign w4157 = w2752 & ~w2706;
assign w4158 = ~w2752 & ~w2712;
assign w4159 = w2752 & ~w2717;
assign w4160 = ~w2752 & w2730;
assign w4161 = w2752 & w2725;
assign w4162 = ~w2752 & ~w2692;
assign w4163 = w2752 & ~w2695;
assign w4164 = ~w2752 & w2612;
assign w4165 = w2752 & w2607;
assign w4166 = ~w2752 & ~w2596;
assign w4167 = w2752 & ~w2601;
assign w4168 = ~w2752 & w2589;
assign w4169 = w2752 & w2584;
assign w4170 = ~w2752 & ~w2574;
assign w4171 = w2752 & ~w2577;
assign w4172 = ~w2752 & ~w2566;
assign w4173 = w2752 & ~w2569;
assign w4174 = ~w2752 & ~w2555;
assign w4175 = w2752 & ~w2560;
assign w4176 = ~w2752 & w2549;
assign w4177 = w2752 & w2544;
assign w4178 = ~w2752 & ~w2535;
assign w4179 = w2752 & ~w2538;
assign w4180 = ~w2752 & w2661;
assign w4181 = w2752 & w2656;
assign w4182 = ~w2752 & ~w2645;
assign w4183 = w2752 & ~w2650;
assign w4184 = ~w2752 & w2638;
assign w4185 = w2752 & w2633;
assign w4186 = ~w2752 & ~w2623;
assign w4187 = w2752 & ~w2626;
assign w4188 = ~w2752 & ~w2457;
assign w4189 = w2752 & ~w2462;
assign w4190 = ~w2752 & ~w2433;
assign w4191 = w2752 & ~w2438;
assign w4192 = ~w2752 & w2449;
assign w4193 = w2752 & w2444;
assign w4194 = ~w2752 & ~w2469;
assign w4195 = w2752 & ~w2472;
assign w4196 = ~w2752 & w2421;
assign w4197 = w2752 & w2418;
assign w4198 = ~w2752 & ~w2411;
assign w4199 = w2752 & ~w2414;
assign w4200 = ~w2752 & w2406;
assign w4201 = w2752 & w2401;
assign w4202 = ~w2752 & ~w2389;
assign w4203 = w2752 & ~w2394;
assign w4204 = ~w2752 & ~w2314;
assign w4205 = w2752 & ~w2317;
assign w4206 = ~w2752 & ~w2303;
assign w4207 = w2752 & ~w2308;
assign w4208 = ~w2752 & w2297;
assign w4209 = w2752 & w2292;
assign w4210 = ~w2752 & ~w2283;
assign w4211 = w2752 & ~w2286;
assign w4212 = ~w2752 & w2380;
assign w4213 = w2752 & w2377;
assign w4214 = ~w2752 & ~w2370;
assign w4215 = w2752 & ~w2373;
assign w4216 = ~w2752 & w2364;
assign w4217 = w2752 & w2361;
assign w4218 = ~w2752 & ~w2354;
assign w4219 = w2752 & ~w2357;
assign w4220 = ~w2752 & ~w2346;
assign w4221 = w2752 & ~w2349;
assign w4222 = ~w2752 & ~w2338;
assign w4223 = w2752 & ~w2341;
assign w4224 = ~w2752 & ~w2331;
assign w4225 = w2752 & ~w2334;
assign w4226 = ~w2752 & ~w1185;
assign w4227 = w2752 & ~w1189;
assign w4228 = ~w397 & w5731;
assign w4229 = ~w976 & w5732;
assign w4230 = w549 & ~w398;
assign w4231 = in0_0 & w544;
assign w4232 = ~w393 & w5733;
assign w4233 = w1128 & ~w977;
assign w4234 = in2_0 & w1104;
assign w4235 = ~w972 & w5734;
assign w4236 = in2_1 & w1104;
assign w4237 = ~w972 & w5735;
assign w4238 = in0_1 & w544;
assign w4239 = ~w393 & w5736;
assign w4240 = in0_2 & w544;
assign w4241 = ~w393 & w5737;
assign w4242 = in2_2 & w1104;
assign w4243 = ~w972 & w5738;
assign w4244 = (in0_3 & w563) | (in0_3 & w5739) | (w563 & w5739);
assign w4245 = in0_3 & ~w3702;
assign w4246 = ~w563 & w5740;
assign w4247 = in1_3 & w3702;
assign w4248 = (in2_3 & w1142) | (in2_3 & w5741) | (w1142 & w5741);
assign w4249 = in2_3 & ~w3703;
assign w4250 = ~w1142 & w5742;
assign w4251 = in3_3 & w3703;
assign w4252 = in0_4 & w544;
assign w4253 = ~w393 & w5743;
assign w4254 = in2_4 & w1104;
assign w4255 = ~w972 & w5744;
assign w4256 = (in0_5 & w563) | (in0_5 & w5745) | (w563 & w5745);
assign w4257 = in0_5 & ~w3702;
assign w4258 = ~w563 & w5746;
assign w4259 = in1_5 & w3702;
assign w4260 = (in2_5 & w1142) | (in2_5 & w5747) | (w1142 & w5747);
assign w4261 = in2_5 & ~w3703;
assign w4262 = ~w1142 & w5748;
assign w4263 = in3_5 & w3703;
assign w4264 = in0_6 & w544;
assign w4265 = ~w393 & w5749;
assign w4266 = in2_6 & w1104;
assign w4267 = ~w972 & w5750;
assign w4268 = in0_11 & w544;
assign w4269 = ~w393 & w5751;
assign w4270 = in2_11 & w1104;
assign w4271 = ~w972 & w5752;
assign w4272 = in0_12 & w544;
assign w4273 = ~w393 & w5753;
assign w4274 = in2_12 & w1104;
assign w4275 = ~w972 & w5754;
assign w4276 = in0_10 & w544;
assign w4277 = ~w393 & w5755;
assign w4278 = in2_10 & w1104;
assign w4279 = ~w972 & w5756;
assign w4280 = in0_14 & w544;
assign w4281 = ~w393 & w5757;
assign w4282 = in2_14 & w1104;
assign w4283 = ~w972 & w5758;
assign w4284 = in0_15 & w544;
assign w4285 = ~w393 & w5759;
assign w4286 = in2_15 & w1104;
assign w4287 = ~w972 & w5760;
assign w4288 = in0_13 & w544;
assign w4289 = ~w393 & w5761;
assign w4290 = in2_13 & w1104;
assign w4291 = ~w972 & w5762;
assign w4292 = in2_8 & w1104;
assign w4293 = ~w972 & w5763;
assign w4294 = in0_8 & w544;
assign w4295 = ~w393 & w5764;
assign w4296 = in0_9 & w544;
assign w4297 = ~w393 & w5765;
assign w4298 = in2_9 & w1104;
assign w4299 = ~w972 & w5766;
assign w4300 = in0_7 & w544;
assign w4301 = ~w393 & w5767;
assign w4302 = in2_7 & w1104;
assign w4303 = ~w972 & w5768;
assign w4304 = in0_19 & w544;
assign w4305 = ~w393 & w5769;
assign w4306 = in2_19 & w1104;
assign w4307 = ~w972 & w5770;
assign w4308 = in0_18 & w544;
assign w4309 = ~w393 & w5771;
assign w4310 = in2_18 & w1104;
assign w4311 = ~w972 & w5772;
assign w4312 = in0_20 & w544;
assign w4313 = ~w393 & w5773;
assign w4314 = in2_20 & w1104;
assign w4315 = ~w972 & w5774;
assign w4316 = (in0_21 & w563) | (in0_21 & w5775) | (w563 & w5775);
assign w4317 = in0_21 & ~w3702;
assign w4318 = ~w563 & w5776;
assign w4319 = in1_21 & w3702;
assign w4320 = (in2_21 & w1142) | (in2_21 & w5777) | (w1142 & w5777);
assign w4321 = in2_21 & ~w3703;
assign w4322 = ~w1142 & w5778;
assign w4323 = in3_21 & w3703;
assign w4324 = in0_22 & w544;
assign w4325 = ~w393 & w5779;
assign w4326 = in2_22 & w1104;
assign w4327 = ~w972 & w5780;
assign w4328 = (in0_16 & w563) | (in0_16 & w5781) | (w563 & w5781);
assign w4329 = in0_16 & ~w3702;
assign w4330 = ~w563 & w5782;
assign w4331 = in1_16 & w3702;
assign w4332 = (in2_16 & w1142) | (in2_16 & w5783) | (w1142 & w5783);
assign w4333 = in2_16 & ~w3703;
assign w4334 = ~w1142 & w5784;
assign w4335 = in3_16 & w3703;
assign w4336 = in2_17 & w1104;
assign w4337 = ~w972 & w5785;
assign w4338 = in0_17 & w544;
assign w4339 = ~w393 & w5786;
assign w4340 = (in0_27 & w563) | (in0_27 & w5787) | (w563 & w5787);
assign w4341 = in0_27 & ~w3702;
assign w4342 = ~w563 & w5788;
assign w4343 = in1_27 & w3702;
assign w4344 = (in2_27 & w1142) | (in2_27 & w5789) | (w1142 & w5789);
assign w4345 = in2_27 & ~w3703;
assign w4346 = ~w1142 & w5790;
assign w4347 = in3_27 & w3703;
assign w4348 = (in0_28 & w563) | (in0_28 & w5791) | (w563 & w5791);
assign w4349 = in0_28 & ~w3702;
assign w4350 = ~w563 & w5792;
assign w4351 = in1_28 & w3702;
assign w4352 = (in2_28 & w1142) | (in2_28 & w5793) | (w1142 & w5793);
assign w4353 = in2_28 & ~w3703;
assign w4354 = ~w1142 & w5794;
assign w4355 = in3_28 & w3703;
assign w4356 = (in0_26 & w563) | (in0_26 & w5795) | (w563 & w5795);
assign w4357 = in0_26 & ~w3702;
assign w4358 = ~w563 & w5796;
assign w4359 = in1_26 & w3702;
assign w4360 = (in2_26 & w1142) | (in2_26 & w5797) | (w1142 & w5797);
assign w4361 = in2_26 & ~w3703;
assign w4362 = ~w1142 & w5798;
assign w4363 = in3_26 & w3703;
assign w4364 = (in0_30 & w563) | (in0_30 & w5799) | (w563 & w5799);
assign w4365 = in0_30 & ~w3702;
assign w4366 = ~w563 & w5800;
assign w4367 = in1_30 & w3702;
assign w4368 = (in2_30 & w1142) | (in2_30 & w5801) | (w1142 & w5801);
assign w4369 = in2_30 & ~w3703;
assign w4370 = ~w1142 & w5802;
assign w4371 = in3_30 & w3703;
assign w4372 = (in0_31 & w563) | (in0_31 & w5803) | (w563 & w5803);
assign w4373 = in0_31 & ~w3702;
assign w4374 = ~w563 & w5804;
assign w4375 = in1_31 & w3702;
assign w4376 = (in2_31 & w1142) | (in2_31 & w5805) | (w1142 & w5805);
assign w4377 = in2_31 & ~w3703;
assign w4378 = ~w1142 & w5806;
assign w4379 = in3_31 & w3703;
assign w4380 = (in0_29 & w563) | (in0_29 & w5807) | (w563 & w5807);
assign w4381 = in0_29 & ~w3702;
assign w4382 = ~w563 & w5808;
assign w4383 = in1_29 & w3702;
assign w4384 = (in2_29 & w1142) | (in2_29 & w5809) | (w1142 & w5809);
assign w4385 = in2_29 & ~w3703;
assign w4386 = ~w1142 & w5810;
assign w4387 = in3_29 & w3703;
assign w4388 = (in0_24 & w563) | (in0_24 & w5811) | (w563 & w5811);
assign w4389 = in0_24 & ~w3702;
assign w4390 = ~w563 & w5812;
assign w4391 = in1_24 & w3702;
assign w4392 = (in2_24 & w1142) | (in2_24 & w5813) | (w1142 & w5813);
assign w4393 = in2_24 & ~w3703;
assign w4394 = ~w1142 & w5814;
assign w4395 = in3_24 & w3703;
assign w4396 = (in0_25 & w563) | (in0_25 & w5815) | (w563 & w5815);
assign w4397 = in0_25 & ~w3702;
assign w4398 = ~w563 & w5816;
assign w4399 = in1_25 & w3702;
assign w4400 = (in2_25 & w1142) | (in2_25 & w5817) | (w1142 & w5817);
assign w4401 = in2_25 & ~w3703;
assign w4402 = ~w1142 & w5818;
assign w4403 = in3_25 & w3703;
assign w4404 = (in0_23 & w563) | (in0_23 & w5819) | (w563 & w5819);
assign w4405 = in0_23 & ~w3702;
assign w4406 = ~w563 & w5820;
assign w4407 = in1_23 & w3702;
assign w4408 = (in2_23 & w1142) | (in2_23 & w5821) | (w1142 & w5821);
assign w4409 = in2_23 & ~w3703;
assign w4410 = ~w1142 & w5822;
assign w4411 = in3_23 & w3703;
assign w4412 = w1535 & w1507;
assign w4413 = (in0_39 & w563) | (in0_39 & w5823) | (w563 & w5823);
assign w4414 = in0_39 & ~w3702;
assign w4415 = ~w563 & w5824;
assign w4416 = in1_39 & w3702;
assign w4417 = (in2_39 & w1142) | (in2_39 & w5825) | (w1142 & w5825);
assign w4418 = in2_39 & ~w3703;
assign w4419 = ~w1142 & w5826;
assign w4420 = in3_39 & w3703;
assign w4421 = (in0_45 & w563) | (in0_45 & w5827) | (w563 & w5827);
assign w4422 = in0_45 & ~w3702;
assign w4423 = ~w563 & w5828;
assign w4424 = in1_45 & w3702;
assign w4425 = (in2_45 & w1142) | (in2_45 & w5829) | (w1142 & w5829);
assign w4426 = in2_45 & ~w3703;
assign w4427 = ~w1142 & w5830;
assign w4428 = in3_45 & w3703;
assign w4429 = (in0_40 & w563) | (in0_40 & w5831) | (w563 & w5831);
assign w4430 = in0_40 & ~w3702;
assign w4431 = ~w563 & w5832;
assign w4432 = in1_40 & w3702;
assign w4433 = (in2_40 & w1142) | (in2_40 & w5833) | (w1142 & w5833);
assign w4434 = in2_40 & ~w3703;
assign w4435 = ~w1142 & w5834;
assign w4436 = in3_40 & w3703;
assign w4437 = (in0_41 & w563) | (in0_41 & w5835) | (w563 & w5835);
assign w4438 = in0_41 & ~w3702;
assign w4439 = ~w563 & w5836;
assign w4440 = in1_41 & w3702;
assign w4441 = (in2_41 & w1142) | (in2_41 & w5837) | (w1142 & w5837);
assign w4442 = in2_41 & ~w3703;
assign w4443 = ~w1142 & w5838;
assign w4444 = in3_41 & w3703;
assign w4445 = (in2_46 & w1142) | (in2_46 & w5839) | (w1142 & w5839);
assign w4446 = in2_46 & ~w3703;
assign w4447 = ~w1142 & w5840;
assign w4448 = in3_46 & w3703;
assign w4449 = (in0_46 & w563) | (in0_46 & w5841) | (w563 & w5841);
assign w4450 = in0_46 & ~w3702;
assign w4451 = ~w563 & w5842;
assign w4452 = in1_46 & w3702;
assign w4453 = (in0_47 & w563) | (in0_47 & w5843) | (w563 & w5843);
assign w4454 = in0_47 & ~w3702;
assign w4455 = ~w563 & w5844;
assign w4456 = in1_47 & w3702;
assign w4457 = (in2_47 & w1142) | (in2_47 & w5845) | (w1142 & w5845);
assign w4458 = in2_47 & ~w3703;
assign w4459 = ~w1142 & w5846;
assign w4460 = in3_47 & w3703;
assign w4461 = (in0_43 & w563) | (in0_43 & w5847) | (w563 & w5847);
assign w4462 = in0_43 & ~w3702;
assign w4463 = ~w563 & w5848;
assign w4464 = in1_43 & w3702;
assign w4465 = (in2_43 & w1142) | (in2_43 & w5849) | (w1142 & w5849);
assign w4466 = in2_43 & ~w3703;
assign w4467 = ~w1142 & w5850;
assign w4468 = in3_43 & w3703;
assign w4469 = (in0_44 & w563) | (in0_44 & w5851) | (w563 & w5851);
assign w4470 = in0_44 & ~w3702;
assign w4471 = ~w563 & w5852;
assign w4472 = in1_44 & w3702;
assign w4473 = (in2_44 & w1142) | (in2_44 & w5853) | (w1142 & w5853);
assign w4474 = in2_44 & ~w3703;
assign w4475 = ~w1142 & w5854;
assign w4476 = in3_44 & w3703;
assign w4477 = (in0_42 & w563) | (in0_42 & w5855) | (w563 & w5855);
assign w4478 = in0_42 & ~w3702;
assign w4479 = ~w563 & w5856;
assign w4480 = in1_42 & w3702;
assign w4481 = (in2_42 & w1142) | (in2_42 & w5857) | (w1142 & w5857);
assign w4482 = in2_42 & ~w3703;
assign w4483 = ~w1142 & w5858;
assign w4484 = in3_42 & w3703;
assign w4485 = in2_32 & w1104;
assign w4486 = ~w972 & w5859;
assign w4487 = in0_32 & w544;
assign w4488 = ~w393 & w5860;
assign w4489 = in0_33 & w544;
assign w4490 = ~w393 & w5861;
assign w4491 = in2_33 & w1104;
assign w4492 = ~w972 & w5862;
assign w4493 = in2_34 & w1104;
assign w4494 = ~w972 & w5863;
assign w4495 = in0_34 & w544;
assign w4496 = ~w393 & w5864;
assign w4497 = (in0_37 & w563) | (in0_37 & w5865) | (w563 & w5865);
assign w4498 = in0_37 & ~w3702;
assign w4499 = ~w563 & w5866;
assign w4500 = in1_37 & w3702;
assign w4501 = (in2_37 & w1142) | (in2_37 & w5867) | (w1142 & w5867);
assign w4502 = in2_37 & ~w3703;
assign w4503 = ~w1142 & w5868;
assign w4504 = in3_37 & w3703;
assign w4505 = (in2_38 & w1142) | (in2_38 & w5869) | (w1142 & w5869);
assign w4506 = in2_38 & ~w3703;
assign w4507 = ~w1142 & w5870;
assign w4508 = in3_38 & w3703;
assign w4509 = (in0_38 & w563) | (in0_38 & w5871) | (w563 & w5871);
assign w4510 = in0_38 & ~w3702;
assign w4511 = ~w563 & w5872;
assign w4512 = in1_38 & w3702;
assign w4513 = (in0_36 & w563) | (in0_36 & w5873) | (w563 & w5873);
assign w4514 = in0_36 & ~w3702;
assign w4515 = ~w563 & w5874;
assign w4516 = in1_36 & w3702;
assign w4517 = (in2_36 & w1142) | (in2_36 & w5875) | (w1142 & w5875);
assign w4518 = in2_36 & ~w3703;
assign w4519 = ~w1142 & w5876;
assign w4520 = in3_36 & w3703;
assign w4521 = (in0_35 & w563) | (in0_35 & w5877) | (w563 & w5877);
assign w4522 = in0_35 & ~w3702;
assign w4523 = ~w563 & w5878;
assign w4524 = in1_35 & w3702;
assign w4525 = (in2_35 & w1142) | (in2_35 & w5879) | (w1142 & w5879);
assign w4526 = in2_35 & ~w3703;
assign w4527 = ~w1142 & w5880;
assign w4528 = in3_35 & w3703;
assign w4529 = ~w1629 & ~w1653;
assign w4530 = in0_55 & w544;
assign w4531 = ~w393 & w5881;
assign w4532 = in2_55 & w1104;
assign w4533 = ~w972 & w5882;
assign w4534 = in2_54 & w1104;
assign w4535 = ~w972 & w5883;
assign w4536 = in0_54 & w544;
assign w4537 = ~w393 & w5884;
assign w4538 = in0_52 & w544;
assign w4539 = ~w393 & w5885;
assign w4540 = in2_52 & w1104;
assign w4541 = ~w972 & w5886;
assign w4542 = in0_51 & w544;
assign w4543 = ~w393 & w5887;
assign w4544 = in2_51 & w1104;
assign w4545 = ~w972 & w5888;
assign w4546 = in0_53 & w544;
assign w4547 = ~w393 & w5889;
assign w4548 = in2_53 & w1104;
assign w4549 = ~w972 & w5890;
assign w4550 = in0_49 & w544;
assign w4551 = ~w393 & w5891;
assign w4552 = in2_49 & w1104;
assign w4553 = ~w972 & w5892;
assign w4554 = in2_48 & w1104;
assign w4555 = ~w972 & w5893;
assign w4556 = in0_48 & w544;
assign w4557 = ~w393 & w5894;
assign w4558 = in2_50 & w1104;
assign w4559 = ~w972 & w5895;
assign w4560 = in0_50 & w544;
assign w4561 = ~w393 & w5896;
assign w4562 = in0_57 & w544;
assign w4563 = ~w393 & w5897;
assign w4564 = in2_57 & w1104;
assign w4565 = ~w972 & w5898;
assign w4566 = in0_56 & w544;
assign w4567 = ~w393 & w5899;
assign w4568 = in2_56 & w1104;
assign w4569 = ~w972 & w5900;
assign w4570 = in0_58 & w544;
assign w4571 = ~w393 & w5901;
assign w4572 = in2_58 & w1104;
assign w4573 = ~w972 & w5902;
assign w4574 = in0_60 & w544;
assign w4575 = ~w393 & w5903;
assign w4576 = in2_60 & w1104;
assign w4577 = ~w972 & w5904;
assign w4578 = in0_59 & w544;
assign w4579 = ~w393 & w5905;
assign w4580 = in2_59 & w1104;
assign w4581 = ~w972 & w5906;
assign w4582 = (in2_62 & w1142) | (in2_62 & w5907) | (w1142 & w5907);
assign w4583 = in2_62 & ~w3703;
assign w4584 = ~w1142 & w5908;
assign w4585 = in3_62 & w3703;
assign w4586 = (in0_62 & w563) | (in0_62 & w5909) | (w563 & w5909);
assign w4587 = in0_62 & ~w3702;
assign w4588 = ~w563 & w5910;
assign w4589 = in1_62 & w3702;
assign w4590 = (in0_63 & w563) | (in0_63 & w5911) | (w563 & w5911);
assign w4591 = in0_63 & ~w3702;
assign w4592 = ~w563 & w5912;
assign w4593 = in1_63 & w3702;
assign w4594 = (in2_63 & w1142) | (in2_63 & w5913) | (w1142 & w5913);
assign w4595 = in2_63 & ~w3703;
assign w4596 = ~w1142 & w5914;
assign w4597 = in3_63 & w3703;
assign w4598 = in0_61 & w544;
assign w4599 = ~w393 & w5915;
assign w4600 = in2_61 & w1104;
assign w4601 = ~w972 & w5916;
assign w4602 = (in0_67 & w563) | (in0_67 & w5917) | (w563 & w5917);
assign w4603 = in0_67 & ~w3702;
assign w4604 = ~w563 & w5918;
assign w4605 = in1_67 & w3702;
assign w4606 = (in2_67 & w1142) | (in2_67 & w5919) | (w1142 & w5919);
assign w4607 = in2_67 & ~w3703;
assign w4608 = ~w1142 & w5920;
assign w4609 = in3_67 & w3703;
assign w4610 = in2_66 & w1104;
assign w4611 = ~w972 & w5921;
assign w4612 = in0_66 & w544;
assign w4613 = ~w393 & w5922;
assign w4614 = in0_65 & w544;
assign w4615 = ~w393 & w5923;
assign w4616 = in2_65 & w1104;
assign w4617 = ~w972 & w5924;
assign w4618 = in2_64 & w1104;
assign w4619 = ~w972 & w5925;
assign w4620 = in0_64 & w544;
assign w4621 = ~w393 & w5926;
assign w4622 = (in0_68 & w563) | (in0_68 & w5927) | (w563 & w5927);
assign w4623 = in0_68 & ~w3702;
assign w4624 = ~w563 & w5928;
assign w4625 = in1_68 & w3702;
assign w4626 = (in2_68 & w1142) | (in2_68 & w5929) | (w1142 & w5929);
assign w4627 = in2_68 & ~w3703;
assign w4628 = ~w1142 & w5930;
assign w4629 = in3_68 & w3703;
assign w4630 = in0_69 & w544;
assign w4631 = ~w393 & w5931;
assign w4632 = in2_69 & w1104;
assign w4633 = ~w972 & w5932;
assign w4634 = (in0_71 & w563) | (in0_71 & w5933) | (w563 & w5933);
assign w4635 = in0_71 & ~w3702;
assign w4636 = ~w563 & w5934;
assign w4637 = in1_71 & w3702;
assign w4638 = (in2_71 & w1142) | (in2_71 & w5935) | (w1142 & w5935);
assign w4639 = in2_71 & ~w3703;
assign w4640 = ~w1142 & w5936;
assign w4641 = in3_71 & w3703;
assign w4642 = in2_70 & w1104;
assign w4643 = ~w972 & w5937;
assign w4644 = in0_70 & w544;
assign w4645 = ~w393 & w5938;
assign w4646 = ~w1962 & ~w1995;
assign w4647 = (in0_83 & w563) | (in0_83 & w5939) | (w563 & w5939);
assign w4648 = in0_83 & ~w3702;
assign w4649 = ~w563 & w5940;
assign w4650 = in1_83 & w3702;
assign w4651 = (in2_83 & w1142) | (in2_83 & w5941) | (w1142 & w5941);
assign w4652 = in2_83 & ~w3703;
assign w4653 = ~w1142 & w5942;
assign w4654 = in3_83 & w3703;
assign w4655 = (in2_88 & w1142) | (in2_88 & w5943) | (w1142 & w5943);
assign w4656 = in2_88 & ~w3703;
assign w4657 = ~w1142 & w5944;
assign w4658 = in3_88 & w3703;
assign w4659 = (in0_88 & w563) | (in0_88 & w5945) | (w563 & w5945);
assign w4660 = in0_88 & ~w3702;
assign w4661 = ~w563 & w5946;
assign w4662 = in1_88 & w3702;
assign w4663 = (in0_89 & w563) | (in0_89 & w5947) | (w563 & w5947);
assign w4664 = in0_89 & ~w3702;
assign w4665 = ~w563 & w5948;
assign w4666 = in1_89 & w3702;
assign w4667 = (in2_89 & w1142) | (in2_89 & w5949) | (w1142 & w5949);
assign w4668 = in2_89 & ~w3703;
assign w4669 = ~w1142 & w5950;
assign w4670 = in3_89 & w3703;
assign w4671 = (in0_87 & w563) | (in0_87 & w5951) | (w563 & w5951);
assign w4672 = in0_87 & ~w3702;
assign w4673 = ~w563 & w5952;
assign w4674 = in1_87 & w3702;
assign w4675 = (in2_87 & w1142) | (in2_87 & w5953) | (w1142 & w5953);
assign w4676 = in2_87 & ~w3703;
assign w4677 = ~w1142 & w5954;
assign w4678 = in3_87 & w3703;
assign w4679 = in0_91 & w544;
assign w4680 = ~w393 & w5955;
assign w4681 = in2_91 & w1104;
assign w4682 = ~w972 & w5956;
assign w4683 = in2_90 & w1104;
assign w4684 = ~w972 & w5957;
assign w4685 = in0_90 & w544;
assign w4686 = ~w393 & w5958;
assign w4687 = in2_86 & w1104;
assign w4688 = ~w972 & w5959;
assign w4689 = in0_86 & w544;
assign w4690 = ~w393 & w5960;
assign w4691 = in0_85 & w544;
assign w4692 = ~w393 & w5961;
assign w4693 = in2_85 & w1104;
assign w4694 = ~w972 & w5962;
assign w4695 = in0_84 & w544;
assign w4696 = ~w393 & w5963;
assign w4697 = in2_84 & w1104;
assign w4698 = ~w972 & w5964;
assign w4699 = (in2_78 & w1142) | (in2_78 & w5965) | (w1142 & w5965);
assign w4700 = in2_78 & ~w3703;
assign w4701 = ~w1142 & w5966;
assign w4702 = in3_78 & w3703;
assign w4703 = (in0_78 & w563) | (in0_78 & w5967) | (w563 & w5967);
assign w4704 = in0_78 & ~w3702;
assign w4705 = ~w563 & w5968;
assign w4706 = in1_78 & w3702;
assign w4707 = in0_77 & w544;
assign w4708 = ~w393 & w5969;
assign w4709 = in2_77 & w1104;
assign w4710 = ~w972 & w5970;
assign w4711 = in2_72 & w1104;
assign w4712 = ~w972 & w5971;
assign w4713 = in0_72 & w544;
assign w4714 = ~w393 & w5972;
assign w4715 = in0_73 & w544;
assign w4716 = ~w393 & w5973;
assign w4717 = in2_73 & w1104;
assign w4718 = ~w972 & w5974;
assign w4719 = (in0_79 & w563) | (in0_79 & w5975) | (w563 & w5975);
assign w4720 = in0_79 & ~w3702;
assign w4721 = ~w563 & w5976;
assign w4722 = in1_79 & w3702;
assign w4723 = (in2_79 & w1142) | (in2_79 & w5977) | (w1142 & w5977);
assign w4724 = in2_79 & ~w3703;
assign w4725 = ~w1142 & w5978;
assign w4726 = in3_79 & w3703;
assign w4727 = in0_75 & w544;
assign w4728 = ~w393 & w5979;
assign w4729 = in2_75 & w1104;
assign w4730 = ~w972 & w5980;
assign w4731 = in0_76 & w544;
assign w4732 = ~w393 & w5981;
assign w4733 = in2_76 & w1104;
assign w4734 = ~w972 & w5982;
assign w4735 = in2_74 & w1104;
assign w4736 = ~w972 & w5983;
assign w4737 = in0_74 & w544;
assign w4738 = ~w393 & w5984;
assign w4739 = (in0_119 & w563) | (in0_119 & w5985) | (w563 & w5985);
assign w4740 = in0_119 & ~w3702;
assign w4741 = ~w563 & w5986;
assign w4742 = in1_119 & w3702;
assign w4743 = (in2_119 & w1142) | (in2_119 & w5987) | (w1142 & w5987);
assign w4744 = in2_119 & ~w3703;
assign w4745 = ~w1142 & w5988;
assign w4746 = in3_119 & w3703;
assign w4747 = in2_118 & w1104;
assign w4748 = ~w972 & w5989;
assign w4749 = in0_118 & w544;
assign w4750 = ~w393 & w5990;
assign w4751 = in0_117 & w544;
assign w4752 = ~w393 & w5991;
assign w4753 = in2_117 & w1104;
assign w4754 = ~w972 & w5992;
assign w4755 = (in0_116 & w563) | (in0_116 & w5993) | (w563 & w5993);
assign w4756 = in0_116 & ~w3702;
assign w4757 = ~w563 & w5994;
assign w4758 = in1_116 & w3702;
assign w4759 = (in2_116 & w1142) | (in2_116 & w5995) | (w1142 & w5995);
assign w4760 = in2_116 & ~w3703;
assign w4761 = ~w1142 & w5996;
assign w4762 = in3_116 & w3703;
assign w4763 = (in0_126 & w563) | (in0_126 & w5997) | (w563 & w5997);
assign w4764 = in0_126 & ~w3702;
assign w4765 = ~w563 & w5998;
assign w4766 = in1_126 & w3702;
assign w4767 = (in2_126 & w1142) | (in2_126 & w5999) | (w1142 & w5999);
assign w4768 = in2_126 & ~w3703;
assign w4769 = ~w1142 & w6000;
assign w4770 = in3_126 & w3703;
assign w4771 = (in0_125 & w563) | (in0_125 & w6001) | (w563 & w6001);
assign w4772 = in0_125 & ~w3702;
assign w4773 = ~w563 & w6002;
assign w4774 = in1_125 & w3702;
assign w4775 = (in2_125 & w1142) | (in2_125 & w6003) | (w1142 & w6003);
assign w4776 = in2_125 & ~w3703;
assign w4777 = ~w1142 & w6004;
assign w4778 = in3_125 & w3703;
assign w4779 = (in0_124 & w563) | (in0_124 & w6005) | (w563 & w6005);
assign w4780 = in0_124 & ~w3702;
assign w4781 = ~w563 & w6006;
assign w4782 = in1_124 & w3702;
assign w4783 = (in2_124 & w1142) | (in2_124 & w6007) | (w1142 & w6007);
assign w4784 = in2_124 & ~w3703;
assign w4785 = ~w1142 & w6008;
assign w4786 = in3_124 & w3703;
assign w4787 = in0_115 & w544;
assign w4788 = ~w393 & w6009;
assign w4789 = in2_115 & w1104;
assign w4790 = ~w972 & w6010;
assign w4791 = in2_114 & w1104;
assign w4792 = ~w972 & w6011;
assign w4793 = in0_114 & w544;
assign w4794 = ~w393 & w6012;
assign w4795 = (in0_113 & w563) | (in0_113 & w6013) | (w563 & w6013);
assign w4796 = in0_113 & ~w3702;
assign w4797 = ~w563 & w6014;
assign w4798 = in1_113 & w3702;
assign w4799 = (in2_113 & w1142) | (in2_113 & w6015) | (w1142 & w6015);
assign w4800 = in2_113 & ~w3703;
assign w4801 = ~w1142 & w6016;
assign w4802 = in3_113 & w3703;
assign w4803 = (in2_112 & w1142) | (in2_112 & w6017) | (w1142 & w6017);
assign w4804 = in2_112 & ~w3703;
assign w4805 = ~w1142 & w6018;
assign w4806 = in3_112 & w3703;
assign w4807 = (in0_112 & w563) | (in0_112 & w6019) | (w563 & w6019);
assign w4808 = in0_112 & ~w3702;
assign w4809 = ~w563 & w6020;
assign w4810 = in1_112 & w3702;
assign w4811 = in0_109 & w544;
assign w4812 = ~w393 & w6021;
assign w4813 = in2_109 & w1104;
assign w4814 = ~w972 & w6022;
assign w4815 = in2_110 & w1104;
assign w4816 = ~w972 & w6023;
assign w4817 = in0_110 & w544;
assign w4818 = ~w393 & w6024;
assign w4819 = in0_108 & w544;
assign w4820 = ~w393 & w6025;
assign w4821 = in2_108 & w1104;
assign w4822 = ~w972 & w6026;
assign w4823 = (in0_111 & w563) | (in0_111 & w6027) | (w563 & w6027);
assign w4824 = in0_111 & ~w3702;
assign w4825 = ~w563 & w6028;
assign w4826 = in1_111 & w3702;
assign w4827 = (in2_111 & w1142) | (in2_111 & w6029) | (w1142 & w6029);
assign w4828 = in2_111 & ~w3703;
assign w4829 = ~w1142 & w6030;
assign w4830 = in3_111 & w3703;
assign w4831 = ~w2326 & w6031;
assign w4832 = (in0_103 & w563) | (in0_103 & w6032) | (w563 & w6032);
assign w4833 = in0_103 & ~w3702;
assign w4834 = ~w563 & w6033;
assign w4835 = in1_103 & w3702;
assign w4836 = (in2_103 & w1142) | (in2_103 & w6034) | (w1142 & w6034);
assign w4837 = in2_103 & ~w3703;
assign w4838 = ~w1142 & w6035;
assign w4839 = in3_103 & w3703;
assign w4840 = in2_102 & w1104;
assign w4841 = ~w972 & w6036;
assign w4842 = in0_102 & w544;
assign w4843 = ~w393 & w6037;
assign w4844 = in0_101 & w544;
assign w4845 = ~w393 & w6038;
assign w4846 = in2_101 & w1104;
assign w4847 = ~w972 & w6039;
assign w4848 = (in0_100 & w563) | (in0_100 & w6040) | (w563 & w6040);
assign w4849 = in0_100 & ~w3702;
assign w4850 = ~w563 & w6041;
assign w4851 = in1_100 & w3702;
assign w4852 = (in2_100 & w1142) | (in2_100 & w6042) | (w1142 & w6042);
assign w4853 = in2_100 & ~w3703;
assign w4854 = ~w1142 & w6043;
assign w4855 = in3_100 & w3703;
assign w4856 = (in0_99 & w563) | (in0_99 & w6044) | (w563 & w6044);
assign w4857 = in0_99 & ~w3702;
assign w4858 = ~w563 & w6045;
assign w4859 = in1_99 & w3702;
assign w4860 = (in2_99 & w1142) | (in2_99 & w6046) | (w1142 & w6046);
assign w4861 = in2_99 & ~w3703;
assign w4862 = ~w1142 & w6047;
assign w4863 = in3_99 & w3703;
assign w4864 = in2_98 & w1104;
assign w4865 = ~w972 & w6048;
assign w4866 = in0_98 & w544;
assign w4867 = ~w393 & w6049;
assign w4868 = in0_97 & w544;
assign w4869 = ~w393 & w6050;
assign w4870 = in2_97 & w1104;
assign w4871 = ~w972 & w6051;
assign w4872 = in2_96 & w1104;
assign w4873 = ~w972 & w6052;
assign w4874 = in0_96 & w544;
assign w4875 = ~w393 & w6053;
assign w4876 = ~w2591 & ~w2578;
assign w4877 = (in0_107 & w563) | (in0_107 & w6054) | (w563 & w6054);
assign w4878 = in0_107 & ~w3702;
assign w4879 = ~w563 & w6055;
assign w4880 = in1_107 & w3702;
assign w4881 = (in2_107 & w1142) | (in2_107 & w6056) | (w1142 & w6056);
assign w4882 = in2_107 & ~w3703;
assign w4883 = ~w1142 & w6057;
assign w4884 = in3_107 & w3703;
assign w4885 = in2_106 & w1104;
assign w4886 = ~w972 & w6058;
assign w4887 = in0_106 & w544;
assign w4888 = ~w393 & w6059;
assign w4889 = in0_105 & w544;
assign w4890 = ~w393 & w6060;
assign w4891 = in2_105 & w1104;
assign w4892 = ~w972 & w6061;
assign w4893 = in2_104 & w1104;
assign w4894 = ~w972 & w6062;
assign w4895 = in0_104 & w544;
assign w4896 = ~w393 & w6063;
assign w4897 = ~w2640 & ~w2627;
assign w4898 = (in0_95 & w563) | (in0_95 & w6064) | (w563 & w6064);
assign w4899 = in0_95 & ~w3702;
assign w4900 = ~w563 & w6065;
assign w4901 = in1_95 & w3702;
assign w4902 = (in2_95 & w1142) | (in2_95 & w6066) | (w1142 & w6066);
assign w4903 = in2_95 & ~w3703;
assign w4904 = ~w1142 & w6067;
assign w4905 = in3_95 & w3703;
assign w4906 = in0_92 & w544;
assign w4907 = ~w393 & w6068;
assign w4908 = in2_92 & w1104;
assign w4909 = ~w972 & w6069;
assign w4910 = in0_93 & w544;
assign w4911 = ~w393 & w6070;
assign w4912 = in2_93 & w1104;
assign w4913 = ~w972 & w6071;
assign w4914 = in2_94 & w1104;
assign w4915 = ~w972 & w6072;
assign w4916 = in0_94 & w544;
assign w4917 = ~w393 & w6073;
assign w4918 = ~w2736 & ~w2696;
assign w4919 = ~w223 & ~w220;
assign w4920 = ~w251 & ~w248;
assign w4921 = w262 & ~w254;
assign w4922 = w275 & w278;
assign w4923 = ~w284 & ~w281;
assign w4924 = ~w237 & ~w240;
assign w4925 = w207 & w304;
assign w4926 = ~w229 & ~w329;
assign w4927 = ~w354 & ~w351;
assign w4928 = ~w422 & w247;
assign w4929 = ~w244 & ~w430;
assign w4930 = ~w440 & ~w523;
assign w4931 = ~w461 & ~w528;
assign w4932 = w468 & ~w529;
assign w4933 = ~w541 & ~w538;
assign w4934 = w307 & w545;
assign w4935 = ~w562 & w544;
assign w4936 = ~w568 & w6074;
assign w4937 = (in0_0 & w568) | (in0_0 & w6075) | (w568 & w6075);
assign w4938 = ~w802 & ~w799;
assign w4939 = ~w830 & ~w827;
assign w4940 = w841 & ~w833;
assign w4941 = w854 & w857;
assign w4942 = ~w863 & ~w860;
assign w4943 = ~w816 & ~w819;
assign w4944 = w786 & w883;
assign w4945 = ~w808 & ~w908;
assign w4946 = ~w933 & ~w930;
assign w4947 = ~w1001 & w826;
assign w4948 = ~w823 & ~w1009;
assign w4949 = ~w1101 & ~w1098;
assign w4950 = ~w1019 & ~w1109;
assign w4951 = ~w1040 & ~w1114;
assign w4952 = w1047 & ~w1115;
assign w4953 = w886 & w1124;
assign w4954 = ~w1141 & w1104;
assign w4955 = ~w1147 & w6076;
assign w4956 = (in2_0 & w1147) | (in2_0 & w6077) | (w1147 & w6077);
assign w4957 = ~w1147 & w6078;
assign w4958 = (in2_1 & w1147) | (in2_1 & w6079) | (w1147 & w6079);
assign w4959 = ~w568 & w6080;
assign w4960 = (in0_1 & w568) | (in0_1 & w6081) | (w568 & w6081);
assign w4961 = ~w568 & w6082;
assign w4962 = (in0_2 & w568) | (in0_2 & w6083) | (w568 & w6083);
assign w4963 = ~w1147 & w6084;
assign w4964 = (in2_2 & w1147) | (in2_2 & w6085) | (w1147 & w6085);
assign w4965 = ~w568 & w6086;
assign w4966 = (in0_4 & w568) | (in0_4 & w6087) | (w568 & w6087);
assign w4967 = ~w1147 & w6088;
assign w4968 = (in2_4 & w1147) | (in2_4 & w6089) | (w1147 & w6089);
assign w4969 = ~w568 & w6090;
assign w4970 = (in0_6 & w568) | (in0_6 & w6091) | (w568 & w6091);
assign w4971 = ~w1147 & w6092;
assign w4972 = (in2_6 & w1147) | (in2_6 & w6093) | (w1147 & w6093);
assign w4973 = ~w568 & w6094;
assign w4974 = (in0_11 & w568) | (in0_11 & w6095) | (w568 & w6095);
assign w4975 = ~w1147 & w6096;
assign w4976 = (in2_11 & w1147) | (in2_11 & w6097) | (w1147 & w6097);
assign w4977 = ~w568 & w6098;
assign w4978 = (in0_12 & w568) | (in0_12 & w6099) | (w568 & w6099);
assign w4979 = ~w1147 & w6100;
assign w4980 = (in2_12 & w1147) | (in2_12 & w6101) | (w1147 & w6101);
assign w4981 = ~w568 & w6102;
assign w4982 = (in0_10 & w568) | (in0_10 & w6103) | (w568 & w6103);
assign w4983 = ~w1147 & w6104;
assign w4984 = (in2_10 & w1147) | (in2_10 & w6105) | (w1147 & w6105);
assign w4985 = ~w568 & w6106;
assign w4986 = (in0_14 & w568) | (in0_14 & w6107) | (w568 & w6107);
assign w4987 = ~w1147 & w6108;
assign w4988 = (in2_14 & w1147) | (in2_14 & w6109) | (w1147 & w6109);
assign w4989 = ~w568 & w6110;
assign w4990 = (in0_15 & w568) | (in0_15 & w6111) | (w568 & w6111);
assign w4991 = ~w1147 & w6112;
assign w4992 = (in2_15 & w1147) | (in2_15 & w6113) | (w1147 & w6113);
assign w4993 = ~w568 & w6114;
assign w4994 = (in0_13 & w568) | (in0_13 & w6115) | (w568 & w6115);
assign w4995 = ~w1147 & w6116;
assign w4996 = (in2_13 & w1147) | (in2_13 & w6117) | (w1147 & w6117);
assign w4997 = ~w1147 & w6118;
assign w4998 = (in2_8 & w1147) | (in2_8 & w6119) | (w1147 & w6119);
assign w4999 = ~w568 & w6120;
assign w5000 = (in0_8 & w568) | (in0_8 & w6441) | (w568 & w6441);
assign w5001 = ~w568 & w6442;
assign w5002 = (in0_9 & w568) | (in0_9 & w6443) | (w568 & w6443);
assign w5003 = ~w1147 & w6444;
assign w5004 = (in2_9 & w1147) | (in2_9 & w6445) | (w1147 & w6445);
assign w5005 = ~w568 & w6446;
assign w5006 = (in0_7 & w568) | (in0_7 & w6447) | (w568 & w6447);
assign w5007 = ~w1147 & w6448;
assign w5008 = (in2_7 & w1147) | (in2_7 & w6449) | (w1147 & w6449);
assign w5009 = ~w568 & w6450;
assign w5010 = (in0_19 & w568) | (in0_19 & w6451) | (w568 & w6451);
assign w5011 = ~w1147 & w6452;
assign w5012 = (in2_19 & w1147) | (in2_19 & w6453) | (w1147 & w6453);
assign w5013 = ~w568 & w6454;
assign w5014 = (in0_18 & w568) | (in0_18 & w6455) | (w568 & w6455);
assign w5015 = ~w1147 & w6456;
assign w5016 = (in2_18 & w1147) | (in2_18 & w6457) | (w1147 & w6457);
assign w5017 = ~w568 & w6458;
assign w5018 = (in0_20 & w568) | (in0_20 & w6459) | (w568 & w6459);
assign w5019 = ~w1147 & w6460;
assign w5020 = (in2_20 & w1147) | (in2_20 & w6461) | (w1147 & w6461);
assign w5021 = ~w568 & w6462;
assign w5022 = (in0_22 & w568) | (in0_22 & w6463) | (w568 & w6463);
assign w5023 = ~w1147 & w6464;
assign w5024 = (in2_22 & w1147) | (in2_22 & w6465) | (w1147 & w6465);
assign w5025 = ~w1147 & w6466;
assign w5026 = (in2_17 & w1147) | (in2_17 & w6467) | (w1147 & w6467);
assign w5027 = ~w568 & w6468;
assign w5028 = (in0_17 & w568) | (in0_17 & w6469) | (w568 & w6469);
assign w5029 = ~w1147 & w6470;
assign w5030 = (in2_32 & w1147) | (in2_32 & w6471) | (w1147 & w6471);
assign w5031 = ~w568 & w6472;
assign w5032 = (in0_32 & w568) | (in0_32 & w6473) | (w568 & w6473);
assign w5033 = ~w568 & w6474;
assign w5034 = (in0_33 & w568) | (in0_33 & w6475) | (w568 & w6475);
assign w5035 = ~w1147 & w6476;
assign w5036 = (in2_33 & w1147) | (in2_33 & w6477) | (w1147 & w6477);
assign w5037 = ~w1147 & w6478;
assign w5038 = (in2_34 & w1147) | (in2_34 & w6479) | (w1147 & w6479);
assign w5039 = ~w568 & w6480;
assign w5040 = (in0_34 & w568) | (in0_34 & w6481) | (w568 & w6481);
assign w5041 = ~w568 & w6482;
assign w5042 = (in0_55 & w568) | (in0_55 & w6483) | (w568 & w6483);
assign w5043 = ~w1147 & w6484;
assign w5044 = (in2_55 & w1147) | (in2_55 & w6485) | (w1147 & w6485);
assign w5045 = ~w1147 & w6486;
assign w5046 = (in2_54 & w1147) | (in2_54 & w6487) | (w1147 & w6487);
assign w5047 = ~w568 & w6488;
assign w5048 = (in0_54 & w568) | (in0_54 & w6489) | (w568 & w6489);
assign w5049 = ~w568 & w6490;
assign w5050 = (in0_52 & w568) | (in0_52 & w6491) | (w568 & w6491);
assign w5051 = ~w1147 & w6492;
assign w5052 = (in2_52 & w1147) | (in2_52 & w6493) | (w1147 & w6493);
assign w5053 = ~w568 & w6494;
assign w5054 = (in0_51 & w568) | (in0_51 & w6495) | (w568 & w6495);
assign w5055 = ~w1147 & w6496;
assign w5056 = (in2_51 & w1147) | (in2_51 & w6497) | (w1147 & w6497);
assign w5057 = ~w568 & w6498;
assign w5058 = (in0_53 & w568) | (in0_53 & w6499) | (w568 & w6499);
assign w5059 = ~w1147 & w6500;
assign w5060 = (in2_53 & w1147) | (in2_53 & w6501) | (w1147 & w6501);
assign w5061 = ~w568 & w6502;
assign w5062 = (in0_49 & w568) | (in0_49 & w6503) | (w568 & w6503);
assign w5063 = ~w1147 & w6504;
assign w5064 = (in2_49 & w1147) | (in2_49 & w6505) | (w1147 & w6505);
assign w5065 = ~w1147 & w6506;
assign w5066 = (in2_48 & w1147) | (in2_48 & w6507) | (w1147 & w6507);
assign w5067 = ~w568 & w6508;
assign w5068 = (in0_48 & w568) | (in0_48 & w6509) | (w568 & w6509);
assign w5069 = ~w1147 & w6510;
assign w5070 = (in2_50 & w1147) | (in2_50 & w6511) | (w1147 & w6511);
assign w5071 = ~w568 & w6512;
assign w5072 = (in0_50 & w568) | (in0_50 & w6513) | (w568 & w6513);
assign w5073 = ~w568 & w6514;
assign w5074 = (in0_57 & w568) | (in0_57 & w6515) | (w568 & w6515);
assign w5075 = ~w1147 & w6516;
assign w5076 = (in2_57 & w1147) | (in2_57 & w6517) | (w1147 & w6517);
assign w5077 = ~w568 & w6518;
assign w5078 = (in0_56 & w568) | (in0_56 & w6519) | (w568 & w6519);
assign w5079 = ~w1147 & w6520;
assign w5080 = (in2_56 & w1147) | (in2_56 & w6521) | (w1147 & w6521);
assign w5081 = ~w568 & w6522;
assign w5082 = (in0_58 & w568) | (in0_58 & w6523) | (w568 & w6523);
assign w5083 = ~w1147 & w6524;
assign w5084 = (in2_58 & w1147) | (in2_58 & w6525) | (w1147 & w6525);
assign w5085 = ~w568 & w6526;
assign w5086 = (in0_60 & w568) | (in0_60 & w6527) | (w568 & w6527);
assign w5087 = ~w1147 & w6528;
assign w5088 = (in2_60 & w1147) | (in2_60 & w6529) | (w1147 & w6529);
assign w5089 = ~w568 & w6530;
assign w5090 = (in0_59 & w568) | (in0_59 & w6531) | (w568 & w6531);
assign w5091 = ~w1147 & w6532;
assign w5092 = (in2_59 & w1147) | (in2_59 & w6533) | (w1147 & w6533);
assign w5093 = ~w568 & w6534;
assign w5094 = (in0_61 & w568) | (in0_61 & w6535) | (w568 & w6535);
assign w5095 = ~w1147 & w6536;
assign w5096 = (in2_61 & w1147) | (in2_61 & w6537) | (w1147 & w6537);
assign w5097 = ~w1147 & w6538;
assign w5098 = (in2_66 & w1147) | (in2_66 & w6539) | (w1147 & w6539);
assign w5099 = ~w568 & w6540;
assign w5100 = (in0_66 & w568) | (in0_66 & w6541) | (w568 & w6541);
assign w5101 = ~w568 & w6542;
assign w5102 = (in0_65 & w568) | (in0_65 & w6543) | (w568 & w6543);
assign w5103 = ~w1147 & w6544;
assign w5104 = (in2_65 & w1147) | (in2_65 & w6545) | (w1147 & w6545);
assign w5105 = ~w1147 & w6546;
assign w5106 = (in2_64 & w1147) | (in2_64 & w6547) | (w1147 & w6547);
assign w5107 = ~w568 & w6548;
assign w5108 = (in0_64 & w568) | (in0_64 & w6549) | (w568 & w6549);
assign w5109 = ~w568 & w6550;
assign w5110 = (in0_69 & w568) | (in0_69 & w6551) | (w568 & w6551);
assign w5111 = ~w1147 & w6552;
assign w5112 = (in2_69 & w1147) | (in2_69 & w6553) | (w1147 & w6553);
assign w5113 = ~w1147 & w6554;
assign w5114 = (in2_70 & w1147) | (in2_70 & w6555) | (w1147 & w6555);
assign w5115 = ~w568 & w6556;
assign w5116 = (in0_70 & w568) | (in0_70 & w6557) | (w568 & w6557);
assign w5117 = w2059 & w1991;
assign w5118 = w2057 & w2061;
assign w5119 = ~w2027 & ~w2064;
assign w5120 = w2046 & ~w2065;
assign w5121 = (in0_82 & w563) | (in0_82 & w6558) | (w563 & w6558);
assign w5122 = in0_82 & ~w3702;
assign w5123 = ~w563 & w6559;
assign w5124 = in1_82 & w3702;
assign w5125 = (in2_82 & w1142) | (in2_82 & w6560) | (w1142 & w6560);
assign w5126 = in2_82 & ~w3703;
assign w5127 = ~w1142 & w6561;
assign w5128 = in3_82 & w3703;
assign w5129 = ~w568 & w6562;
assign w5130 = (in0_91 & w568) | (in0_91 & w6563) | (w568 & w6563);
assign w5131 = ~w1147 & w6564;
assign w5132 = (in2_91 & w1147) | (in2_91 & w6565) | (w1147 & w6565);
assign w5133 = ~w1147 & w6566;
assign w5134 = (in2_90 & w1147) | (in2_90 & w6567) | (w1147 & w6567);
assign w5135 = ~w568 & w6568;
assign w5136 = (in0_90 & w568) | (in0_90 & w6569) | (w568 & w6569);
assign w5137 = ~w1147 & w6570;
assign w5138 = (in2_86 & w1147) | (in2_86 & w6571) | (w1147 & w6571);
assign w5139 = ~w568 & w6572;
assign w5140 = (in0_86 & w568) | (in0_86 & w6573) | (w568 & w6573);
assign w5141 = ~w568 & w6574;
assign w5142 = (in0_85 & w568) | (in0_85 & w6575) | (w568 & w6575);
assign w5143 = ~w1147 & w6576;
assign w5144 = (in2_85 & w1147) | (in2_85 & w6577) | (w1147 & w6577);
assign w5145 = ~w568 & w6578;
assign w5146 = (in0_84 & w568) | (in0_84 & w6579) | (w568 & w6579);
assign w5147 = ~w1147 & w6580;
assign w5148 = (in2_84 & w1147) | (in2_84 & w6581) | (w1147 & w6581);
assign w5149 = (in0_81 & w563) | (in0_81 & w6582) | (w563 & w6582);
assign w5150 = in0_81 & ~w3702;
assign w5151 = ~w563 & w6583;
assign w5152 = in1_81 & w3702;
assign w5153 = (in2_81 & w1142) | (in2_81 & w6584) | (w1142 & w6584);
assign w5154 = in2_81 & ~w3703;
assign w5155 = ~w1142 & w6585;
assign w5156 = in3_81 & w3703;
assign w5157 = (in0_80 & w563) | (in0_80 & w6586) | (w563 & w6586);
assign w5158 = in0_80 & ~w3702;
assign w5159 = ~w563 & w6587;
assign w5160 = in1_80 & w3702;
assign w5161 = (in2_80 & w1142) | (in2_80 & w6588) | (w1142 & w6588);
assign w5162 = in2_80 & ~w3703;
assign w5163 = ~w1142 & w6589;
assign w5164 = in3_80 & w3703;
assign w5165 = ~w568 & w6590;
assign w5166 = (in0_77 & w568) | (in0_77 & w6591) | (w568 & w6591);
assign w5167 = ~w1147 & w6592;
assign w5168 = (in2_77 & w1147) | (in2_77 & w6593) | (w1147 & w6593);
assign w5169 = ~w1147 & w6594;
assign w5170 = (in2_72 & w1147) | (in2_72 & w6595) | (w1147 & w6595);
assign w5171 = ~w568 & w6596;
assign w5172 = (in0_72 & w568) | (in0_72 & w6597) | (w568 & w6597);
assign w5173 = ~w568 & w6598;
assign w5174 = (in0_73 & w568) | (in0_73 & w6599) | (w568 & w6599);
assign w5175 = ~w1147 & w6600;
assign w5176 = (in2_73 & w1147) | (in2_73 & w6601) | (w1147 & w6601);
assign w5177 = ~w568 & w6602;
assign w5178 = (in0_75 & w568) | (in0_75 & w6603) | (w568 & w6603);
assign w5179 = ~w1147 & w6604;
assign w5180 = (in2_75 & w1147) | (in2_75 & w6605) | (w1147 & w6605);
assign w5181 = ~w568 & w6606;
assign w5182 = (in0_76 & w568) | (in0_76 & w6607) | (w568 & w6607);
assign w5183 = ~w1147 & w6608;
assign w5184 = (in2_76 & w1147) | (in2_76 & w6609) | (w1147 & w6609);
assign w5185 = ~w1147 & w6610;
assign w5186 = (in2_74 & w1147) | (in2_74 & w6611) | (w1147 & w6611);
assign w5187 = ~w568 & w6612;
assign w5188 = (in0_74 & w568) | (in0_74 & w6613) | (w568 & w6613);
assign w5189 = ~w1147 & w6614;
assign w5190 = (in2_118 & w1147) | (in2_118 & w6615) | (w1147 & w6615);
assign w5191 = ~w568 & w6616;
assign w5192 = (in0_118 & w568) | (in0_118 & w6617) | (w568 & w6617);
assign w5193 = ~w568 & w6618;
assign w5194 = (in0_117 & w568) | (in0_117 & w6619) | (w568 & w6619);
assign w5195 = ~w1147 & w6620;
assign w5196 = (in2_117 & w1147) | (in2_117 & w6621) | (w1147 & w6621);
assign w5197 = ~w2287 & ~w2318;
assign w5198 = w2327 & ~w2319;
assign w5199 = (in0_123 & w563) | (in0_123 & w6622) | (w563 & w6622);
assign w5200 = in0_123 & ~w3702;
assign w5201 = ~w563 & w6623;
assign w5202 = in1_123 & w3702;
assign w5203 = (in2_123 & w1142) | (in2_123 & w6624) | (w1142 & w6624);
assign w5204 = in2_123 & ~w3703;
assign w5205 = ~w1142 & w6625;
assign w5206 = in3_123 & w3703;
assign w5207 = (in2_122 & w1142) | (in2_122 & w6626) | (w1142 & w6626);
assign w5208 = in2_122 & ~w3703;
assign w5209 = ~w1142 & w6627;
assign w5210 = in3_122 & w3703;
assign w5211 = (in0_122 & w563) | (in0_122 & w6628) | (w563 & w6628);
assign w5212 = in0_122 & ~w3702;
assign w5213 = ~w563 & w6629;
assign w5214 = in1_122 & w3702;
assign w5215 = (in0_121 & w563) | (in0_121 & w6630) | (w563 & w6630);
assign w5216 = in0_121 & ~w3702;
assign w5217 = ~w563 & w6631;
assign w5218 = in1_121 & w3702;
assign w5219 = (in2_121 & w1142) | (in2_121 & w6632) | (w1142 & w6632);
assign w5220 = in2_121 & ~w3703;
assign w5221 = ~w1142 & w6633;
assign w5222 = in3_121 & w3703;
assign w5223 = (in2_120 & w1142) | (in2_120 & w6634) | (w1142 & w6634);
assign w5224 = in2_120 & ~w3703;
assign w5225 = ~w1142 & w6635;
assign w5226 = in3_120 & w3703;
assign w5227 = (in0_120 & w563) | (in0_120 & w6636) | (w563 & w6636);
assign w5228 = in0_120 & ~w3702;
assign w5229 = ~w563 & w6637;
assign w5230 = in1_120 & w3702;
assign w5231 = w2366 & w2382;
assign w5232 = ~w568 & w6638;
assign w5233 = (in0_115 & w568) | (in0_115 & w6639) | (w568 & w6639);
assign w5234 = ~w1147 & w6640;
assign w5235 = (in2_115 & w1147) | (in2_115 & w6641) | (w1147 & w6641);
assign w5236 = ~w1147 & w6642;
assign w5237 = (in2_114 & w1147) | (in2_114 & w6643) | (w1147 & w6643);
assign w5238 = ~w568 & w6644;
assign w5239 = (in0_114 & w568) | (in0_114 & w6645) | (w568 & w6645);
assign w5240 = ~w568 & w6646;
assign w5241 = (in0_109 & w568) | (in0_109 & w6647) | (w568 & w6647);
assign w5242 = ~w1147 & w6648;
assign w5243 = (in2_109 & w1147) | (in2_109 & w6649) | (w1147 & w6649);
assign w5244 = ~w1147 & w6650;
assign w5245 = (in2_110 & w1147) | (in2_110 & w6651) | (w1147 & w6651);
assign w5246 = ~w568 & w6652;
assign w5247 = (in0_110 & w568) | (in0_110 & w6653) | (w568 & w6653);
assign w5248 = ~w568 & w6654;
assign w5249 = (in0_108 & w568) | (in0_108 & w6655) | (w568 & w6655);
assign w5250 = ~w1147 & w6656;
assign w5251 = (in2_108 & w1147) | (in2_108 & w6657) | (w1147 & w6657);
assign w5252 = ~w2350 & w2493;
assign w5253 = (in2_127 & w1142) | (in2_127 & w6658) | (w1142 & w6658);
assign w5254 = ~w2500 & in0_127;
assign w5255 = ~w2177 & w2181;
assign w5256 = ~w2528 & w2530;
assign w5257 = ~w1147 & w6659;
assign w5258 = (in2_102 & w1147) | (in2_102 & w6660) | (w1147 & w6660);
assign w5259 = ~w568 & w6661;
assign w5260 = (in0_102 & w568) | (in0_102 & w6662) | (w568 & w6662);
assign w5261 = ~w568 & w6663;
assign w5262 = (in0_101 & w568) | (in0_101 & w6664) | (w568 & w6664);
assign w5263 = ~w1147 & w6665;
assign w5264 = (in2_101 & w1147) | (in2_101 & w6666) | (w1147 & w6666);
assign w5265 = ~w2539 & ~w2570;
assign w5266 = ~w1147 & w6667;
assign w5267 = (in2_98 & w1147) | (in2_98 & w6668) | (w1147 & w6668);
assign w5268 = ~w568 & w6669;
assign w5269 = (in0_98 & w568) | (in0_98 & w6670) | (w568 & w6670);
assign w5270 = ~w568 & w6671;
assign w5271 = (in0_97 & w568) | (in0_97 & w6672) | (w568 & w6672);
assign w5272 = ~w1147 & w6673;
assign w5273 = (in2_97 & w1147) | (in2_97 & w6674) | (w1147 & w6674);
assign w5274 = ~w1147 & w6675;
assign w5275 = (in2_96 & w1147) | (in2_96 & w6676) | (w1147 & w6676);
assign w5276 = ~w568 & w6677;
assign w5277 = (in0_96 & w568) | (in0_96 & w6678) | (w568 & w6678);
assign w5278 = ~w1147 & w6679;
assign w5279 = (in2_106 & w1147) | (in2_106 & w6680) | (w1147 & w6680);
assign w5280 = ~w568 & w6681;
assign w5281 = (in0_106 & w568) | (in0_106 & w6682) | (w568 & w6682);
assign w5282 = ~w568 & w6683;
assign w5283 = (in0_105 & w568) | (in0_105 & w6684) | (w568 & w6684);
assign w5284 = ~w1147 & w6685;
assign w5285 = (in2_105 & w1147) | (in2_105 & w6686) | (w1147 & w6686);
assign w5286 = ~w1147 & w6687;
assign w5287 = (in2_104 & w1147) | (in2_104 & w6688) | (w1147 & w6688);
assign w5288 = ~w568 & w6689;
assign w5289 = (in0_104 & w568) | (in0_104 & w6690) | (w568 & w6690);
assign w5290 = ~w568 & w6691;
assign w5291 = (in0_92 & w568) | (in0_92 & w6692) | (w568 & w6692);
assign w5292 = ~w1147 & w6693;
assign w5293 = (in2_92 & w1147) | (in2_92 & w6694) | (w1147 & w6694);
assign w5294 = ~w568 & w6695;
assign w5295 = (in0_93 & w568) | (in0_93 & w6696) | (w568 & w6696);
assign w5296 = ~w1147 & w6697;
assign w5297 = (in2_93 & w1147) | (in2_93 & w6698) | (w1147 & w6698);
assign w5298 = ~w1147 & w6699;
assign w5299 = (in2_94 & w1147) | (in2_94 & w6700) | (w1147 & w6700);
assign w5300 = ~w568 & w6701;
assign w5301 = (in0_94 & w568) | (in0_94 & w6702) | (w568 & w6702);
assign w5302 = ~w2384 & w2505;
assign w5303 = w4225 & ~w2334;
assign w5304 = (w5302 & w7076) | (w5302 & w7077) | (w7076 & w7077);
assign w5305 = w2505 & w7201;
assign w5306 = ~w3660 & ~w3659;
assign w5307 = ~w563 & w6703;
assign w5308 = w574 & ~w3680;
assign w5309 = ~w1142 & w6704;
assign w5310 = w1153 & ~w3691;
assign w5311 = ~w1142 & w6705;
assign w5312 = w1159 & ~w3691;
assign w5313 = ~w563 & w6706;
assign w5314 = w1164 & ~w3680;
assign w5315 = ~w563 & w6707;
assign w5316 = w1172 & ~w3680;
assign w5317 = ~w1142 & w6708;
assign w5318 = w1177 & ~w3691;
assign w5319 = ~w563 & w6709;
assign w5320 = w573 & ~w3680;
assign w5321 = ~w1142 & w6710;
assign w5322 = w1152 & ~w3691;
assign w5323 = ~w563 & w6711;
assign w5324 = w1194 & ~w3680;
assign w5325 = ~w1142 & w6712;
assign w5326 = w1199 & ~w3691;
assign w5327 = ~w563 & w6713;
assign w5328 = w1216 & ~w3680;
assign w5329 = ~w1142 & w6714;
assign w5330 = w1221 & ~w3691;
assign w5331 = ~w563 & w6715;
assign w5332 = w1234 & ~w3680;
assign w5333 = ~w1142 & w6716;
assign w5334 = w1239 & ~w3691;
assign w5335 = ~w563 & w6717;
assign w5336 = w1245 & ~w3680;
assign w5337 = ~w1142 & w6718;
assign w5338 = w1250 & ~w3691;
assign w5339 = ~w563 & w6719;
assign w5340 = w1258 & ~w3680;
assign w5341 = ~w1142 & w6720;
assign w5342 = w1263 & ~w3691;
assign w5343 = ~w563 & w6721;
assign w5344 = w1271 & ~w3680;
assign w5345 = ~w1142 & w6722;
assign w5346 = w1276 & ~w3691;
assign w5347 = ~w563 & w6723;
assign w5348 = w1282 & ~w3680;
assign w5349 = ~w1142 & w6724;
assign w5350 = w1287 & ~w3691;
assign w5351 = ~w563 & w6725;
assign w5352 = w1295 & ~w3680;
assign w5353 = ~w1142 & w6726;
assign w5354 = w1300 & ~w3691;
assign w5355 = ~w1142 & w6727;
assign w5356 = w1309 & ~w3691;
assign w5357 = ~w563 & w6728;
assign w5358 = w1314 & ~w3680;
assign w5359 = ~w563 & w6729;
assign w5360 = w1320 & ~w3680;
assign w5361 = ~w1142 & w6730;
assign w5362 = w1325 & ~w3691;
assign w5363 = ~w563 & w6731;
assign w5364 = w1333 & ~w3680;
assign w5365 = ~w1142 & w6732;
assign w5366 = w1338 & ~w3691;
assign w5367 = ~w563 & w6733;
assign w5368 = w1361 & ~w3680;
assign w5369 = ~w1142 & w6734;
assign w5370 = w1366 & ~w3691;
assign w5371 = ~w563 & w6735;
assign w5372 = w1372 & ~w3680;
assign w5373 = ~w1142 & w6736;
assign w5374 = w1377 & ~w3691;
assign w5375 = ~w563 & w6737;
assign w5376 = w1385 & ~w3680;
assign w5377 = ~w1142 & w6738;
assign w5378 = w1390 & ~w3691;
assign w5379 = ~w563 & w6739;
assign w5380 = w1405 & ~w3680;
assign w5381 = ~w1142 & w6740;
assign w5382 = w1410 & ~w3691;
assign w5383 = ~w1142 & w6741;
assign w5384 = w1431 & ~w3691;
assign w5385 = ~w563 & w6742;
assign w5386 = w1436 & ~w3680;
assign w5387 = ~w1142 & w6743;
assign w5388 = w1619 & ~w3691;
assign w5389 = ~w563 & w6744;
assign w5390 = w1624 & ~w3680;
assign w5391 = ~w563 & w6745;
assign w5392 = w1630 & ~w3680;
assign w5393 = ~w1142 & w6746;
assign w5394 = w1635 & ~w3691;
assign w5395 = ~w1142 & w6747;
assign w5396 = w1641 & ~w3691;
assign w5397 = ~w563 & w6748;
assign w5398 = w1646 & ~w3680;
assign w5399 = ~w563 & w6749;
assign w5400 = w1695 & ~w3680;
assign w5401 = ~w1142 & w6750;
assign w5402 = w1700 & ~w3691;
assign w5403 = ~w1142 & w6751;
assign w5404 = w1707 & ~w3691;
assign w5405 = ~w563 & w6752;
assign w5406 = w1712 & ~w3680;
assign w5407 = ~w563 & w6753;
assign w5408 = w1720 & ~w3680;
assign w5409 = ~w1142 & w6754;
assign w5410 = w1725 & ~w3691;
assign w5411 = ~w563 & w6755;
assign w5412 = w1731 & ~w3680;
assign w5413 = ~w1142 & w6756;
assign w5414 = w1736 & ~w3691;
assign w5415 = ~w563 & w6757;
assign w5416 = w1744 & ~w3680;
assign w5417 = ~w1142 & w6758;
assign w5418 = w1749 & ~w3691;
assign w5419 = ~w563 & w6759;
assign w5420 = w1758 & ~w3680;
assign w5421 = ~w1142 & w6760;
assign w5422 = w1763 & ~w3691;
assign w5423 = ~w1142 & w6761;
assign w5424 = w1769 & ~w3691;
assign w5425 = ~w563 & w6762;
assign w5426 = w1774 & ~w3680;
assign w5427 = ~w1142 & w6763;
assign w5428 = w1782 & ~w3691;
assign w5429 = ~w563 & w6764;
assign w5430 = w1787 & ~w3680;
assign w5431 = ~w563 & w6765;
assign w5432 = w1848 & ~w3680;
assign w5433 = ~w1142 & w6766;
assign w5434 = w1853 & ~w3691;
assign w5435 = ~w563 & w6767;
assign w5436 = w1859 & ~w3680;
assign w5437 = ~w1142 & w6768;
assign w5438 = w1864 & ~w3691;
assign w5439 = ~w563 & w6769;
assign w5440 = w1872 & ~w3680;
assign w5441 = ~w1142 & w6770;
assign w5442 = w1877 & ~w3691;
assign w5443 = ~w563 & w6771;
assign w5444 = w1886 & ~w3680;
assign w5445 = ~w1142 & w6772;
assign w5446 = w1891 & ~w3691;
assign w5447 = w3681 & w574;
assign w5448 = (w574 & w3681) | (w574 & ~w307) | (w3681 & ~w307);
assign w5449 = w3692 & w1153;
assign w5450 = (w1153 & w3692) | (w1153 & ~w886) | (w3692 & ~w886);
assign w5451 = w3694 & w1159;
assign w5452 = (w1159 & w3694) | (w1159 & ~w886) | (w3694 & ~w886);
assign w5453 = w3696 & w1164;
assign w5454 = (w1164 & w3696) | (w1164 & ~w307) | (w3696 & ~w307);
assign w5455 = w3698 & w1172;
assign w5456 = (w1172 & w3698) | (w1172 & ~w307) | (w3698 & ~w307);
assign w5457 = w3700 & w1177;
assign w5458 = (w1177 & w3700) | (w1177 & ~w886) | (w3700 & ~w886);
assign w5459 = w3704 & w1194;
assign w5460 = (w1194 & w3704) | (w1194 & ~w307) | (w3704 & ~w307);
assign w5461 = w3706 & w1199;
assign w5462 = (w1199 & w3706) | (w1199 & ~w886) | (w3706 & ~w886);
assign w5463 = w3708 & w1216;
assign w5464 = (w1216 & w3708) | (w1216 & ~w307) | (w3708 & ~w307);
assign w5465 = w3710 & w1221;
assign w5466 = (w1221 & w3710) | (w1221 & ~w886) | (w3710 & ~w886);
assign w5467 = w3712 & w1234;
assign w5468 = (w1234 & w3712) | (w1234 & ~w307) | (w3712 & ~w307);
assign w5469 = w3714 & w1239;
assign w5470 = (w1239 & w3714) | (w1239 & ~w886) | (w3714 & ~w886);
assign w5471 = w3716 & w1245;
assign w5472 = (w1245 & w3716) | (w1245 & ~w307) | (w3716 & ~w307);
assign w5473 = w3718 & w1250;
assign w5474 = (w1250 & w3718) | (w1250 & ~w886) | (w3718 & ~w886);
assign w5475 = w3720 & w1258;
assign w5476 = (w1258 & w3720) | (w1258 & ~w307) | (w3720 & ~w307);
assign w5477 = w3722 & w1263;
assign w5478 = (w1263 & w3722) | (w1263 & ~w886) | (w3722 & ~w886);
assign w5479 = w3724 & w1271;
assign w5480 = (w1271 & w3724) | (w1271 & ~w307) | (w3724 & ~w307);
assign w5481 = w3726 & w1276;
assign w5482 = (w1276 & w3726) | (w1276 & ~w886) | (w3726 & ~w886);
assign w5483 = w3728 & w1282;
assign w5484 = (w1282 & w3728) | (w1282 & ~w307) | (w3728 & ~w307);
assign w5485 = w3730 & w1287;
assign w5486 = (w1287 & w3730) | (w1287 & ~w886) | (w3730 & ~w886);
assign w5487 = w3732 & w1295;
assign w5488 = (w1295 & w3732) | (w1295 & ~w307) | (w3732 & ~w307);
assign w5489 = w3734 & w1300;
assign w5490 = (w1300 & w3734) | (w1300 & ~w886) | (w3734 & ~w886);
assign w5491 = w3736 & w1309;
assign w5492 = (w1309 & w3736) | (w1309 & ~w886) | (w3736 & ~w886);
assign w5493 = w3738 & w1314;
assign w5494 = (w1314 & w3738) | (w1314 & ~w307) | (w3738 & ~w307);
assign w5495 = w3740 & w1320;
assign w5496 = (w1320 & w3740) | (w1320 & ~w307) | (w3740 & ~w307);
assign w5497 = w3742 & w1325;
assign w5498 = (w1325 & w3742) | (w1325 & ~w886) | (w3742 & ~w886);
assign w5499 = w3744 & w1333;
assign w5500 = (w1333 & w3744) | (w1333 & ~w307) | (w3744 & ~w307);
assign w5501 = w3746 & w1338;
assign w5502 = (w1338 & w3746) | (w1338 & ~w886) | (w3746 & ~w886);
assign w5503 = w3748 & w1361;
assign w5504 = (w1361 & w3748) | (w1361 & ~w307) | (w3748 & ~w307);
assign w5505 = w3750 & w1366;
assign w5506 = (w1366 & w3750) | (w1366 & ~w886) | (w3750 & ~w886);
assign w5507 = w3752 & w1372;
assign w5508 = (w1372 & w3752) | (w1372 & ~w307) | (w3752 & ~w307);
assign w5509 = w3754 & w1377;
assign w5510 = (w1377 & w3754) | (w1377 & ~w886) | (w3754 & ~w886);
assign w5511 = w3756 & w1385;
assign w5512 = (w1385 & w3756) | (w1385 & ~w307) | (w3756 & ~w307);
assign w5513 = w3758 & w1390;
assign w5514 = (w1390 & w3758) | (w1390 & ~w886) | (w3758 & ~w886);
assign w5515 = w3760 & w1405;
assign w5516 = (w1405 & w3760) | (w1405 & ~w307) | (w3760 & ~w307);
assign w5517 = w3762 & w1410;
assign w5518 = (w1410 & w3762) | (w1410 & ~w886) | (w3762 & ~w886);
assign w5519 = w3764 & w1431;
assign w5520 = (w1431 & w3764) | (w1431 & ~w886) | (w3764 & ~w886);
assign w5521 = w3766 & w1436;
assign w5522 = (w1436 & w3766) | (w1436 & ~w307) | (w3766 & ~w307);
assign w5523 = w3768 & w1619;
assign w5524 = (w1619 & w3768) | (w1619 & ~w886) | (w3768 & ~w886);
assign w5525 = w3770 & w1624;
assign w5526 = (w1624 & w3770) | (w1624 & ~w307) | (w3770 & ~w307);
assign w5527 = w3772 & w1630;
assign w5528 = (w1630 & w3772) | (w1630 & ~w307) | (w3772 & ~w307);
assign w5529 = w3774 & w1635;
assign w5530 = (w1635 & w3774) | (w1635 & ~w886) | (w3774 & ~w886);
assign w5531 = w3776 & w1641;
assign w5532 = (w1641 & w3776) | (w1641 & ~w886) | (w3776 & ~w886);
assign w5533 = w3778 & w1646;
assign w5534 = (w1646 & w3778) | (w1646 & ~w307) | (w3778 & ~w307);
assign w5535 = w3812 & w1848;
assign w5536 = (w1848 & w3812) | (w1848 & ~w307) | (w3812 & ~w307);
assign w5537 = w3814 & w1853;
assign w5538 = (w1853 & w3814) | (w1853 & ~w886) | (w3814 & ~w886);
assign w5539 = w3816 & w1859;
assign w5540 = (w1859 & w3816) | (w1859 & ~w307) | (w3816 & ~w307);
assign w5541 = w3818 & w1864;
assign w5542 = (w1864 & w3818) | (w1864 & ~w886) | (w3818 & ~w886);
assign w5543 = w3820 & w1872;
assign w5544 = (w1872 & w3820) | (w1872 & ~w307) | (w3820 & ~w307);
assign w5545 = w3822 & w1877;
assign w5546 = (w1877 & w3822) | (w1877 & ~w886) | (w3822 & ~w886);
assign w5547 = w3824 & w1886;
assign w5548 = (w1886 & w3824) | (w1886 & ~w307) | (w3824 & ~w307);
assign w5549 = w3826 & w1891;
assign w5550 = (w1891 & w3826) | (w1891 & ~w886) | (w3826 & ~w886);
assign w5551 = w3702 & w573;
assign w5552 = (w573 & w3702) | (w573 & ~w307) | (w3702 & ~w307);
assign w5553 = w3703 & w1152;
assign w5554 = (w1152 & w3703) | (w1152 & ~w886) | (w3703 & ~w886);
assign w5555 = w3780 & w1695;
assign w5556 = (w1695 & w3780) | (w1695 & ~w307) | (w3780 & ~w307);
assign w5557 = w3782 & w1700;
assign w5558 = (w1700 & w3782) | (w1700 & ~w886) | (w3782 & ~w886);
assign w5559 = w3784 & w1707;
assign w5560 = (w1707 & w3784) | (w1707 & ~w886) | (w3784 & ~w886);
assign w5561 = w3786 & w1712;
assign w5562 = (w1712 & w3786) | (w1712 & ~w307) | (w3786 & ~w307);
assign w5563 = w3788 & w1720;
assign w5564 = (w1720 & w3788) | (w1720 & ~w307) | (w3788 & ~w307);
assign w5565 = w3790 & w1725;
assign w5566 = (w1725 & w3790) | (w1725 & ~w886) | (w3790 & ~w886);
assign w5567 = w3792 & w1731;
assign w5568 = (w1731 & w3792) | (w1731 & ~w307) | (w3792 & ~w307);
assign w5569 = w3794 & w1736;
assign w5570 = (w1736 & w3794) | (w1736 & ~w886) | (w3794 & ~w886);
assign w5571 = w3796 & w1744;
assign w5572 = (w1744 & w3796) | (w1744 & ~w307) | (w3796 & ~w307);
assign w5573 = w3798 & w1749;
assign w5574 = (w1749 & w3798) | (w1749 & ~w886) | (w3798 & ~w886);
assign w5575 = w3800 & w1758;
assign w5576 = (w1758 & w3800) | (w1758 & ~w307) | (w3800 & ~w307);
assign w5577 = w3802 & w1763;
assign w5578 = (w1763 & w3802) | (w1763 & ~w886) | (w3802 & ~w886);
assign w5579 = w3804 & w1769;
assign w5580 = (w1769 & w3804) | (w1769 & ~w886) | (w3804 & ~w886);
assign w5581 = w3806 & w1774;
assign w5582 = (w1774 & w3806) | (w1774 & ~w307) | (w3806 & ~w307);
assign w5583 = w3808 & w1782;
assign w5584 = (w1782 & w3808) | (w1782 & ~w886) | (w3808 & ~w886);
assign w5585 = w3810 & w1787;
assign w5586 = (w1787 & w3810) | (w1787 & ~w307) | (w3810 & ~w307);
assign w5587 = ~w563 & w6773;
assign w5588 = w1897 & ~w3680;
assign w5589 = ~w1142 & w6774;
assign w5590 = w1902 & ~w3691;
assign w5591 = ~w563 & w6775;
assign w5592 = w1929 & ~w3680;
assign w5593 = ~w1142 & w6776;
assign w5594 = w1934 & ~w3691;
assign w5595 = ~w1142 & w6777;
assign w5596 = w1951 & ~w3691;
assign w5597 = ~w563 & w6778;
assign w5598 = w1956 & ~w3680;
assign w5599 = ~w563 & w6779;
assign w5600 = w1964 & ~w3680;
assign w5601 = ~w1142 & w6780;
assign w5602 = w1969 & ~w3691;
assign w5603 = ~w1142 & w6781;
assign w5604 = w1975 & ~w3691;
assign w5605 = ~w563 & w6782;
assign w5606 = w1980 & ~w3680;
assign w5607 = ~w563 & w6783;
assign w5608 = w2009 & ~w3680;
assign w5609 = ~w1142 & w6784;
assign w5610 = w2014 & ~w3691;
assign w5611 = ~w1142 & w6785;
assign w5612 = w2029 & ~w3691;
assign w5613 = ~w563 & w6786;
assign w5614 = w2034 & ~w3680;
assign w5615 = ~w563 & w6787;
assign w5616 = w2103 & ~w3680;
assign w5617 = ~w1142 & w6788;
assign w5618 = w2108 & ~w3691;
assign w5619 = ~w1142 & w6789;
assign w5620 = w2114 & ~w3691;
assign w5621 = ~w563 & w6790;
assign w5622 = w2119 & ~w3680;
assign w5623 = ~w1142 & w6791;
assign w5624 = w2130 & ~w3691;
assign w5625 = ~w563 & w6792;
assign w5626 = w2135 & ~w3680;
assign w5627 = ~w563 & w6793;
assign w5628 = w2141 & ~w3680;
assign w5629 = ~w1142 & w6794;
assign w5630 = w2146 & ~w3691;
assign w5631 = ~w563 & w6795;
assign w5632 = w2153 & ~w3680;
assign w5633 = ~w1142 & w6796;
assign w5634 = w2158 & ~w3691;
assign w5635 = ~w563 & w6797;
assign w5636 = w2197 & ~w3680;
assign w5637 = ~w1142 & w6798;
assign w5638 = w2202 & ~w3691;
assign w5639 = ~w1142 & w6799;
assign w5640 = w2209 & ~w3691;
assign w5641 = ~w563 & w6800;
assign w5642 = w2214 & ~w3680;
assign w5643 = ~w563 & w6801;
assign w5644 = w2220 & ~w3680;
assign w5645 = ~w1142 & w6802;
assign w5646 = w2225 & ~w3691;
assign w5647 = ~w563 & w6803;
assign w5648 = w2238 & ~w3680;
assign w5649 = ~w1142 & w6804;
assign w5650 = w2243 & ~w3691;
assign w5651 = ~w563 & w6805;
assign w5652 = w2249 & ~w3680;
assign w5653 = ~w1142 & w6806;
assign w5654 = w2254 & ~w3691;
assign w5655 = ~w1142 & w6807;
assign w5656 = w2260 & ~w3691;
assign w5657 = ~w563 & w6808;
assign w5658 = w2265 & ~w3680;
assign w5659 = ~w1142 & w6809;
assign w5660 = w2288 & ~w3691;
assign w5661 = ~w563 & w6810;
assign w5662 = w2293 & ~w3680;
assign w5663 = ~w563 & w6811;
assign w5664 = w2299 & ~w3680;
assign w5665 = ~w1142 & w6812;
assign w5666 = w2304 & ~w3691;
assign w5667 = ~w563 & w6813;
assign w5668 = w2385 & ~w3680;
assign w5669 = ~w1142 & w6814;
assign w5670 = w2390 & ~w3691;
assign w5671 = ~w1142 & w6815;
assign w5672 = w2397 & ~w3691;
assign w5673 = ~w563 & w6816;
assign w5674 = w2402 & ~w3680;
assign w5675 = ~w563 & w6817;
assign w5676 = w2429 & ~w3680;
assign w5677 = ~w1142 & w6818;
assign w5678 = w2434 & ~w3691;
assign w5679 = ~w1142 & w6819;
assign w5680 = w2440 & ~w3691;
assign w5681 = ~w563 & w6820;
assign w5682 = w2445 & ~w3680;
assign w5683 = ~w563 & w6821;
assign w5684 = w2453 & ~w3680;
assign w5685 = ~w1142 & w6822;
assign w5686 = w2458 & ~w3691;
assign w5687 = ~w1142 & w6823;
assign w5688 = w2540 & ~w3691;
assign w5689 = ~w563 & w6824;
assign w5690 = w2545 & ~w3680;
assign w5691 = ~w563 & w6825;
assign w5692 = w2551 & ~w3680;
assign w5693 = ~w1142 & w6826;
assign w5694 = w2556 & ~w3691;
assign w5695 = ~w1142 & w6827;
assign w5696 = w2580 & ~w3691;
assign w5697 = ~w563 & w6828;
assign w5698 = w2585 & ~w3680;
assign w5699 = ~w563 & w6829;
assign w5700 = w2592 & ~w3680;
assign w5701 = ~w1142 & w6830;
assign w5702 = w2597 & ~w3691;
assign w5703 = ~w1142 & w6831;
assign w5704 = w2603 & ~w3691;
assign w5705 = ~w563 & w6832;
assign w5706 = w2608 & ~w3680;
assign w5707 = ~w1142 & w6833;
assign w5708 = w2629 & ~w3691;
assign w5709 = ~w563 & w6834;
assign w5710 = w2634 & ~w3680;
assign w5711 = ~w563 & w6835;
assign w5712 = w2641 & ~w3680;
assign w5713 = ~w1142 & w6836;
assign w5714 = w2646 & ~w3691;
assign w5715 = ~w1142 & w6837;
assign w5716 = w2652 & ~w3691;
assign w5717 = ~w563 & w6838;
assign w5718 = w2657 & ~w3680;
assign w5719 = ~w563 & w6839;
assign w5720 = w2697 & ~w3680;
assign w5721 = ~w1142 & w6840;
assign w5722 = w2702 & ~w3691;
assign w5723 = ~w563 & w6841;
assign w5724 = w2708 & ~w3680;
assign w5725 = ~w1142 & w6842;
assign w5726 = w2713 & ~w3691;
assign w5727 = ~w1142 & w6843;
assign w5728 = w2721 & ~w3691;
assign w5729 = ~w563 & w6844;
assign w5730 = w2726 & ~w3680;
assign w5731 = w412 & w544;
assign w5732 = w991 & w1104;
assign w5733 = w4228 & in0_0;
assign w5734 = w4229 & in2_0;
assign w5735 = w4229 & in2_1;
assign w5736 = w4228 & in0_1;
assign w5737 = w4228 & in0_2;
assign w5738 = w4229 & in2_2;
assign w5739 = (in0_3 & w568) | (in0_3 & w6845) | (w568 & w6845);
assign w5740 = ~w568 & w6846;
assign w5741 = (in2_3 & w1147) | (in2_3 & w6847) | (w1147 & w6847);
assign w5742 = ~w1147 & w6848;
assign w5743 = w4228 & in0_4;
assign w5744 = w4229 & in2_4;
assign w5745 = (in0_5 & w568) | (in0_5 & w6849) | (w568 & w6849);
assign w5746 = ~w568 & w6850;
assign w5747 = (in2_5 & w1147) | (in2_5 & w6851) | (w1147 & w6851);
assign w5748 = ~w1147 & w6852;
assign w5749 = w4228 & in0_6;
assign w5750 = w4229 & in2_6;
assign w5751 = w4228 & in0_11;
assign w5752 = w4229 & in2_11;
assign w5753 = w4228 & in0_12;
assign w5754 = w4229 & in2_12;
assign w5755 = w4228 & in0_10;
assign w5756 = w4229 & in2_10;
assign w5757 = w4228 & in0_14;
assign w5758 = w4229 & in2_14;
assign w5759 = w4228 & in0_15;
assign w5760 = w4229 & in2_15;
assign w5761 = w4228 & in0_13;
assign w5762 = w4229 & in2_13;
assign w5763 = w4229 & in2_8;
assign w5764 = w4228 & in0_8;
assign w5765 = w4228 & in0_9;
assign w5766 = w4229 & in2_9;
assign w5767 = w4228 & in0_7;
assign w5768 = w4229 & in2_7;
assign w5769 = w4228 & in0_19;
assign w5770 = w4229 & in2_19;
assign w5771 = w4228 & in0_18;
assign w5772 = w4229 & in2_18;
assign w5773 = w4228 & in0_20;
assign w5774 = w4229 & in2_20;
assign w5775 = (in0_21 & w568) | (in0_21 & w6853) | (w568 & w6853);
assign w5776 = ~w568 & w6854;
assign w5777 = (in2_21 & w1147) | (in2_21 & w6855) | (w1147 & w6855);
assign w5778 = ~w1147 & w6856;
assign w5779 = w4228 & in0_22;
assign w5780 = w4229 & in2_22;
assign w5781 = (in0_16 & w568) | (in0_16 & w6857) | (w568 & w6857);
assign w5782 = ~w568 & w6858;
assign w5783 = (in2_16 & w1147) | (in2_16 & w6859) | (w1147 & w6859);
assign w5784 = ~w1147 & w6860;
assign w5785 = w4229 & in2_17;
assign w5786 = w4228 & in0_17;
assign w5787 = (in0_27 & w568) | (in0_27 & w6861) | (w568 & w6861);
assign w5788 = ~w568 & w6862;
assign w5789 = (in2_27 & w1147) | (in2_27 & w6863) | (w1147 & w6863);
assign w5790 = w1151 & in3_27;
assign w5791 = ~w572 & in0_28;
assign w5792 = w572 & in1_28;
assign w5793 = ~w1151 & in2_28;
assign w5794 = w1151 & in3_28;
assign w5795 = ~w572 & in0_26;
assign w5796 = w572 & in1_26;
assign w5797 = ~w1151 & in2_26;
assign w5798 = w1151 & in3_26;
assign w5799 = ~w572 & in0_30;
assign w5800 = w572 & in1_30;
assign w5801 = ~w1151 & in2_30;
assign w5802 = w1151 & in3_30;
assign w5803 = ~w572 & in0_31;
assign w5804 = w572 & in1_31;
assign w5805 = ~w1151 & in2_31;
assign w5806 = w1151 & in3_31;
assign w5807 = ~w572 & in0_29;
assign w5808 = w572 & in1_29;
assign w5809 = ~w1151 & in2_29;
assign w5810 = w1151 & in3_29;
assign w5811 = ~w572 & in0_24;
assign w5812 = w572 & in1_24;
assign w5813 = ~w1151 & in2_24;
assign w5814 = w1151 & in3_24;
assign w5815 = ~w572 & in0_25;
assign w5816 = w572 & in1_25;
assign w5817 = ~w1151 & in2_25;
assign w5818 = w1151 & in3_25;
assign w5819 = ~w572 & in0_23;
assign w5820 = w572 & in1_23;
assign w5821 = ~w1151 & in2_23;
assign w5822 = w1151 & in3_23;
assign w5823 = ~w572 & in0_39;
assign w5824 = w572 & in1_39;
assign w5825 = ~w1151 & in2_39;
assign w5826 = w1151 & in3_39;
assign w5827 = ~w572 & in0_45;
assign w5828 = w572 & in1_45;
assign w5829 = ~w1151 & in2_45;
assign w5830 = w1151 & in3_45;
assign w5831 = ~w572 & in0_40;
assign w5832 = w572 & in1_40;
assign w5833 = ~w1151 & in2_40;
assign w5834 = w1151 & in3_40;
assign w5835 = ~w572 & in0_41;
assign w5836 = w572 & in1_41;
assign w5837 = ~w1151 & in2_41;
assign w5838 = w1151 & in3_41;
assign w5839 = ~w1151 & in2_46;
assign w5840 = w1151 & in3_46;
assign w5841 = ~w572 & in0_46;
assign w5842 = w572 & in1_46;
assign w5843 = ~w572 & in0_47;
assign w5844 = w572 & in1_47;
assign w5845 = ~w1151 & in2_47;
assign w5846 = w1151 & in3_47;
assign w5847 = ~w572 & in0_43;
assign w5848 = w572 & in1_43;
assign w5849 = ~w1151 & in2_43;
assign w5850 = w1151 & in3_43;
assign w5851 = ~w572 & in0_44;
assign w5852 = w572 & in1_44;
assign w5853 = ~w1151 & in2_44;
assign w5854 = w1151 & in3_44;
assign w5855 = ~w572 & in0_42;
assign w5856 = w572 & in1_42;
assign w5857 = ~w1151 & in2_42;
assign w5858 = w1151 & in3_42;
assign w5859 = w4229 & in2_32;
assign w5860 = w4228 & in0_32;
assign w5861 = w4228 & in0_33;
assign w5862 = w4229 & in2_33;
assign w5863 = w4229 & in2_34;
assign w5864 = w4228 & in0_34;
assign w5865 = ~w572 & in0_37;
assign w5866 = w572 & in1_37;
assign w5867 = ~w1151 & in2_37;
assign w5868 = w1151 & in3_37;
assign w5869 = ~w1151 & in2_38;
assign w5870 = w1151 & in3_38;
assign w5871 = ~w572 & in0_38;
assign w5872 = w572 & in1_38;
assign w5873 = ~w572 & in0_36;
assign w5874 = w572 & in1_36;
assign w5875 = ~w1151 & in2_36;
assign w5876 = w1151 & in3_36;
assign w5877 = ~w572 & in0_35;
assign w5878 = w572 & in1_35;
assign w5879 = ~w1151 & in2_35;
assign w5880 = w1151 & in3_35;
assign w5881 = w4228 & in0_55;
assign w5882 = w4229 & in2_55;
assign w5883 = w4229 & in2_54;
assign w5884 = w4228 & in0_54;
assign w5885 = w4228 & in0_52;
assign w5886 = w4229 & in2_52;
assign w5887 = w4228 & in0_51;
assign w5888 = w4229 & in2_51;
assign w5889 = w4228 & in0_53;
assign w5890 = w4229 & in2_53;
assign w5891 = w4228 & in0_49;
assign w5892 = w4229 & in2_49;
assign w5893 = w4229 & in2_48;
assign w5894 = w4228 & in0_48;
assign w5895 = w4229 & in2_50;
assign w5896 = w4228 & in0_50;
assign w5897 = w4228 & in0_57;
assign w5898 = w4229 & in2_57;
assign w5899 = w4228 & in0_56;
assign w5900 = w4229 & in2_56;
assign w5901 = w4228 & in0_58;
assign w5902 = w4229 & in2_58;
assign w5903 = w4228 & in0_60;
assign w5904 = w4229 & in2_60;
assign w5905 = w4228 & in0_59;
assign w5906 = w4229 & in2_59;
assign w5907 = ~w1151 & in2_62;
assign w5908 = w1151 & in3_62;
assign w5909 = ~w572 & in0_62;
assign w5910 = w572 & in1_62;
assign w5911 = ~w572 & in0_63;
assign w5912 = w572 & in1_63;
assign w5913 = ~w1151 & in2_63;
assign w5914 = w1151 & in3_63;
assign w5915 = w4228 & in0_61;
assign w5916 = w4229 & in2_61;
assign w5917 = ~w572 & in0_67;
assign w5918 = w572 & in1_67;
assign w5919 = ~w1151 & in2_67;
assign w5920 = w1151 & in3_67;
assign w5921 = w4229 & in2_66;
assign w5922 = w4228 & in0_66;
assign w5923 = w4228 & in0_65;
assign w5924 = w4229 & in2_65;
assign w5925 = w4229 & in2_64;
assign w5926 = w4228 & in0_64;
assign w5927 = ~w572 & in0_68;
assign w5928 = w572 & in1_68;
assign w5929 = ~w1151 & in2_68;
assign w5930 = w1151 & in3_68;
assign w5931 = w4228 & in0_69;
assign w5932 = w4229 & in2_69;
assign w5933 = ~w572 & in0_71;
assign w5934 = w572 & in1_71;
assign w5935 = ~w1151 & in2_71;
assign w5936 = w1151 & in3_71;
assign w5937 = w4229 & in2_70;
assign w5938 = w4228 & in0_70;
assign w5939 = ~w572 & in0_83;
assign w5940 = w572 & in1_83;
assign w5941 = ~w1151 & in2_83;
assign w5942 = w1151 & in3_83;
assign w5943 = ~w1151 & in2_88;
assign w5944 = w1151 & in3_88;
assign w5945 = ~w572 & in0_88;
assign w5946 = w572 & in1_88;
assign w5947 = ~w572 & in0_89;
assign w5948 = w572 & in1_89;
assign w5949 = ~w1151 & in2_89;
assign w5950 = w1151 & in3_89;
assign w5951 = ~w572 & in0_87;
assign w5952 = w572 & in1_87;
assign w5953 = ~w1151 & in2_87;
assign w5954 = w1151 & in3_87;
assign w5955 = w4228 & in0_91;
assign w5956 = w4229 & in2_91;
assign w5957 = w4229 & in2_90;
assign w5958 = w4228 & in0_90;
assign w5959 = w4229 & in2_86;
assign w5960 = w4228 & in0_86;
assign w5961 = w4228 & in0_85;
assign w5962 = w4229 & in2_85;
assign w5963 = w4228 & in0_84;
assign w5964 = w4229 & in2_84;
assign w5965 = ~w1151 & in2_78;
assign w5966 = w1151 & in3_78;
assign w5967 = ~w572 & in0_78;
assign w5968 = w572 & in1_78;
assign w5969 = w4228 & in0_77;
assign w5970 = w4229 & in2_77;
assign w5971 = w4229 & in2_72;
assign w5972 = w4228 & in0_72;
assign w5973 = w4228 & in0_73;
assign w5974 = w4229 & in2_73;
assign w5975 = ~w572 & in0_79;
assign w5976 = w572 & in1_79;
assign w5977 = ~w1151 & in2_79;
assign w5978 = w1151 & in3_79;
assign w5979 = w4228 & in0_75;
assign w5980 = w4229 & in2_75;
assign w5981 = w4228 & in0_76;
assign w5982 = w4229 & in2_76;
assign w5983 = w4229 & in2_74;
assign w5984 = w4228 & in0_74;
assign w5985 = ~w572 & in0_119;
assign w5986 = w572 & in1_119;
assign w5987 = ~w1151 & in2_119;
assign w5988 = w1151 & in3_119;
assign w5989 = w4229 & in2_118;
assign w5990 = w4228 & in0_118;
assign w5991 = w4228 & in0_117;
assign w5992 = w4229 & in2_117;
assign w5993 = ~w572 & in0_116;
assign w5994 = w572 & in1_116;
assign w5995 = ~w1151 & in2_116;
assign w5996 = w1151 & in3_116;
assign w5997 = ~w572 & in0_126;
assign w5998 = w572 & in1_126;
assign w5999 = ~w1151 & in2_126;
assign w6000 = w1151 & in3_126;
assign w6001 = ~w572 & in0_125;
assign w6002 = w572 & in1_125;
assign w6003 = ~w1151 & in2_125;
assign w6004 = w1151 & in3_125;
assign w6005 = ~w572 & in0_124;
assign w6006 = w572 & in1_124;
assign w6007 = ~w1151 & in2_124;
assign w6008 = w1151 & in3_124;
assign w6009 = w4228 & in0_115;
assign w6010 = w4229 & in2_115;
assign w6011 = w4229 & in2_114;
assign w6012 = w4228 & in0_114;
assign w6013 = ~w572 & in0_113;
assign w6014 = w572 & in1_113;
assign w6015 = ~w1151 & in2_113;
assign w6016 = w1151 & in3_113;
assign w6017 = ~w1151 & in2_112;
assign w6018 = w1151 & in3_112;
assign w6019 = ~w572 & in0_112;
assign w6020 = w572 & in1_112;
assign w6021 = w4228 & in0_109;
assign w6022 = w4229 & in2_109;
assign w6023 = w4229 & in2_110;
assign w6024 = w4228 & in0_110;
assign w6025 = w4228 & in0_108;
assign w6026 = w4229 & in2_108;
assign w6027 = ~w572 & in0_111;
assign w6028 = w572 & in1_111;
assign w6029 = ~w1151 & in2_111;
assign w6030 = w1151 & in3_111;
assign w6031 = ~w2324 & ~w2395;
assign w6032 = ~w572 & in0_103;
assign w6033 = w572 & in1_103;
assign w6034 = ~w1151 & in2_103;
assign w6035 = w1151 & in3_103;
assign w6036 = w4229 & in2_102;
assign w6037 = w4228 & in0_102;
assign w6038 = w4228 & in0_101;
assign w6039 = w4229 & in2_101;
assign w6040 = ~w572 & in0_100;
assign w6041 = w572 & in1_100;
assign w6042 = ~w1151 & in2_100;
assign w6043 = w1151 & in3_100;
assign w6044 = ~w572 & in0_99;
assign w6045 = w572 & in1_99;
assign w6046 = ~w1151 & in2_99;
assign w6047 = w1151 & in3_99;
assign w6048 = w4229 & in2_98;
assign w6049 = w4228 & in0_98;
assign w6050 = w4228 & in0_97;
assign w6051 = w4229 & in2_97;
assign w6052 = w4229 & in2_96;
assign w6053 = w4228 & in0_96;
assign w6054 = ~w572 & in0_107;
assign w6055 = w572 & in1_107;
assign w6056 = ~w1151 & in2_107;
assign w6057 = w1151 & in3_107;
assign w6058 = w4229 & in2_106;
assign w6059 = w4228 & in0_106;
assign w6060 = w4228 & in0_105;
assign w6061 = w4229 & in2_105;
assign w6062 = w4229 & in2_104;
assign w6063 = w4228 & in0_104;
assign w6064 = ~w572 & in0_95;
assign w6065 = w572 & in1_95;
assign w6066 = ~w1151 & in2_95;
assign w6067 = w1151 & in3_95;
assign w6068 = w4228 & in0_92;
assign w6069 = w4229 & in2_92;
assign w6070 = w4228 & in0_93;
assign w6071 = w4229 & in2_93;
assign w6072 = w4229 & in2_94;
assign w6073 = w4228 & in0_94;
assign w6074 = w571 & in1_0;
assign w6075 = ~w571 & in0_0;
assign w6076 = w1150 & in3_0;
assign w6077 = ~w1150 & in2_0;
assign w6078 = w1150 & in3_1;
assign w6079 = ~w1150 & in2_1;
assign w6080 = w571 & in1_1;
assign w6081 = ~w571 & in0_1;
assign w6082 = w571 & in1_2;
assign w6083 = ~w571 & in0_2;
assign w6084 = w1150 & in3_2;
assign w6085 = ~w1150 & in2_2;
assign w6086 = w571 & in1_4;
assign w6087 = ~w571 & in0_4;
assign w6088 = w1150 & in3_4;
assign w6089 = ~w1150 & in2_4;
assign w6090 = w571 & in1_6;
assign w6091 = ~w571 & in0_6;
assign w6092 = w1150 & in3_6;
assign w6093 = ~w1150 & in2_6;
assign w6094 = w571 & in1_11;
assign w6095 = ~w571 & in0_11;
assign w6096 = w1150 & in3_11;
assign w6097 = ~w1150 & in2_11;
assign w6098 = w571 & in1_12;
assign w6099 = ~w571 & in0_12;
assign w6100 = w1150 & in3_12;
assign w6101 = ~w1150 & in2_12;
assign w6102 = w571 & in1_10;
assign w6103 = ~w571 & in0_10;
assign w6104 = w1150 & in3_10;
assign w6105 = ~w1150 & in2_10;
assign w6106 = w571 & in1_14;
assign w6107 = ~w571 & in0_14;
assign w6108 = w1150 & in3_14;
assign w6109 = ~w1150 & in2_14;
assign w6110 = w571 & in1_15;
assign w6111 = ~w571 & in0_15;
assign w6112 = w1150 & in3_15;
assign w6113 = ~w1150 & in2_15;
assign w6114 = w571 & in1_13;
assign w6115 = ~w571 & in0_13;
assign w6116 = w1150 & in3_13;
assign w6117 = ~w1150 & in2_13;
assign w6118 = w1150 & in3_8;
assign w6119 = ~w1150 & in2_8;
assign w6120 = w571 & in1_8;
assign w6121 = w3828 & w1897;
assign w6122 = (w1897 & w3828) | (w1897 & ~w307) | (w3828 & ~w307);
assign w6123 = w3830 & w1902;
assign w6124 = (w1902 & w3830) | (w1902 & ~w886) | (w3830 & ~w886);
assign w6125 = w3832 & w1929;
assign w6126 = (w1929 & w3832) | (w1929 & ~w307) | (w3832 & ~w307);
assign w6127 = w3834 & w1934;
assign w6128 = (w1934 & w3834) | (w1934 & ~w886) | (w3834 & ~w886);
assign w6129 = w3840 & w1964;
assign w6130 = (w1964 & w3840) | (w1964 & ~w307) | (w3840 & ~w307);
assign w6131 = w3842 & w1969;
assign w6132 = (w1969 & w3842) | (w1969 & ~w886) | (w3842 & ~w886);
assign w6133 = w3844 & w1975;
assign w6134 = (w1975 & w3844) | (w1975 & ~w886) | (w3844 & ~w886);
assign w6135 = w3846 & w1980;
assign w6136 = (w1980 & w3846) | (w1980 & ~w307) | (w3846 & ~w307);
assign w6137 = w3848 & w2009;
assign w6138 = (w2009 & w3848) | (w2009 & ~w307) | (w3848 & ~w307);
assign w6139 = w3850 & w2014;
assign w6140 = (w2014 & w3850) | (w2014 & ~w886) | (w3850 & ~w886);
assign w6141 = w3852 & w2029;
assign w6142 = (w2029 & w3852) | (w2029 & ~w886) | (w3852 & ~w886);
assign w6143 = w3854 & w2034;
assign w6144 = (w2034 & w3854) | (w2034 & ~w307) | (w3854 & ~w307);
assign w6145 = w3856 & w2103;
assign w6146 = (w2103 & w3856) | (w2103 & ~w307) | (w3856 & ~w307);
assign w6147 = w3858 & w2108;
assign w6148 = (w2108 & w3858) | (w2108 & ~w886) | (w3858 & ~w886);
assign w6149 = w3860 & w2114;
assign w6150 = (w2114 & w3860) | (w2114 & ~w886) | (w3860 & ~w886);
assign w6151 = w3862 & w2119;
assign w6152 = (w2119 & w3862) | (w2119 & ~w307) | (w3862 & ~w307);
assign w6153 = w3864 & w2130;
assign w6154 = (w2130 & w3864) | (w2130 & ~w886) | (w3864 & ~w886);
assign w6155 = w3866 & w2135;
assign w6156 = (w2135 & w3866) | (w2135 & ~w307) | (w3866 & ~w307);
assign w6157 = w3868 & w2141;
assign w6158 = (w2141 & w3868) | (w2141 & ~w307) | (w3868 & ~w307);
assign w6159 = w3870 & w2146;
assign w6160 = (w2146 & w3870) | (w2146 & ~w886) | (w3870 & ~w886);
assign w6161 = w3872 & w2153;
assign w6162 = (w2153 & w3872) | (w2153 & ~w307) | (w3872 & ~w307);
assign w6163 = w3874 & w2158;
assign w6164 = (w2158 & w3874) | (w2158 & ~w886) | (w3874 & ~w886);
assign w6165 = w3908 & w2385;
assign w6166 = (w2385 & w3908) | (w2385 & ~w307) | (w3908 & ~w307);
assign w6167 = w3910 & w2390;
assign w6168 = (w2390 & w3910) | (w2390 & ~w886) | (w3910 & ~w886);
assign w6169 = w3912 & w2397;
assign w6170 = (w2397 & w3912) | (w2397 & ~w886) | (w3912 & ~w886);
assign w6171 = w3914 & w2402;
assign w6172 = (w2402 & w3914) | (w2402 & ~w307) | (w3914 & ~w307);
assign w6173 = w3916 & w2429;
assign w6174 = (w2429 & w3916) | (w2429 & ~w307) | (w3916 & ~w307);
assign w6175 = w3918 & w2434;
assign w6176 = (w2434 & w3918) | (w2434 & ~w886) | (w3918 & ~w886);
assign w6177 = w3920 & w2440;
assign w6178 = (w2440 & w3920) | (w2440 & ~w886) | (w3920 & ~w886);
assign w6179 = w3922 & w2445;
assign w6180 = (w2445 & w3922) | (w2445 & ~w307) | (w3922 & ~w307);
assign w6181 = w3924 & w2453;
assign w6182 = (w2453 & w3924) | (w2453 & ~w307) | (w3924 & ~w307);
assign w6183 = w3926 & w2458;
assign w6184 = (w2458 & w3926) | (w2458 & ~w886) | (w3926 & ~w886);
assign w6185 = w3928 & w2540;
assign w6186 = (w2540 & w3928) | (w2540 & ~w886) | (w3928 & ~w886);
assign w6187 = w3930 & w2545;
assign w6188 = (w2545 & w3930) | (w2545 & ~w307) | (w3930 & ~w307);
assign w6189 = w3932 & w2551;
assign w6190 = (w2551 & w3932) | (w2551 & ~w307) | (w3932 & ~w307);
assign w6191 = w3934 & w2556;
assign w6192 = (w2556 & w3934) | (w2556 & ~w886) | (w3934 & ~w886);
assign w6193 = w3836 & w1951;
assign w6194 = (w1951 & w3836) | (w1951 & ~w886) | (w3836 & ~w886);
assign w6195 = w3838 & w1956;
assign w6196 = (w1956 & w3838) | (w1956 & ~w307) | (w3838 & ~w307);
assign w6197 = w3876 & w2197;
assign w6198 = (w2197 & w3876) | (w2197 & ~w307) | (w3876 & ~w307);
assign w6199 = w3878 & w2202;
assign w6200 = (w2202 & w3878) | (w2202 & ~w886) | (w3878 & ~w886);
assign w6201 = w3880 & w2209;
assign w6202 = (w2209 & w3880) | (w2209 & ~w886) | (w3880 & ~w886);
assign w6203 = w3882 & w2214;
assign w6204 = (w2214 & w3882) | (w2214 & ~w307) | (w3882 & ~w307);
assign w6205 = w3884 & w2220;
assign w6206 = (w2220 & w3884) | (w2220 & ~w307) | (w3884 & ~w307);
assign w6207 = w3886 & w2225;
assign w6208 = (w2225 & w3886) | (w2225 & ~w886) | (w3886 & ~w886);
assign w6209 = w3888 & w2238;
assign w6210 = (w2238 & w3888) | (w2238 & ~w307) | (w3888 & ~w307);
assign w6211 = w3890 & w2243;
assign w6212 = (w2243 & w3890) | (w2243 & ~w886) | (w3890 & ~w886);
assign w6213 = w3892 & w2249;
assign w6214 = (w2249 & w3892) | (w2249 & ~w307) | (w3892 & ~w307);
assign w6215 = w3894 & w2254;
assign w6216 = (w2254 & w3894) | (w2254 & ~w886) | (w3894 & ~w886);
assign w6217 = w3896 & w2260;
assign w6218 = (w2260 & w3896) | (w2260 & ~w886) | (w3896 & ~w886);
assign w6219 = w3898 & w2265;
assign w6220 = (w2265 & w3898) | (w2265 & ~w307) | (w3898 & ~w307);
assign w6221 = w3900 & w2288;
assign w6222 = (w2288 & w3900) | (w2288 & ~w886) | (w3900 & ~w886);
assign w6223 = w3902 & w2293;
assign w6224 = (w2293 & w3902) | (w2293 & ~w307) | (w3902 & ~w307);
assign w6225 = w3904 & w2299;
assign w6226 = (w2299 & w3904) | (w2299 & ~w307) | (w3904 & ~w307);
assign w6227 = w3906 & w2304;
assign w6228 = (w2304 & w3906) | (w2304 & ~w886) | (w3906 & ~w886);
assign w6229 = w3936 & w2580;
assign w6230 = (w2580 & w3936) | (w2580 & ~w886) | (w3936 & ~w886);
assign w6231 = w3938 & w2585;
assign w6232 = (w2585 & w3938) | (w2585 & ~w307) | (w3938 & ~w307);
assign w6233 = w3940 & w2592;
assign w6234 = (w2592 & w3940) | (w2592 & ~w307) | (w3940 & ~w307);
assign w6235 = w3942 & w2597;
assign w6236 = (w2597 & w3942) | (w2597 & ~w886) | (w3942 & ~w886);
assign w6237 = w3944 & w2603;
assign w6238 = (w2603 & w3944) | (w2603 & ~w886) | (w3944 & ~w886);
assign w6239 = w3946 & w2608;
assign w6240 = (w2608 & w3946) | (w2608 & ~w307) | (w3946 & ~w307);
assign w6241 = w3948 & w2629;
assign w6242 = (w2629 & w3948) | (w2629 & ~w886) | (w3948 & ~w886);
assign w6243 = w3950 & w2634;
assign w6244 = (w2634 & w3950) | (w2634 & ~w307) | (w3950 & ~w307);
assign w6245 = w3952 & w2641;
assign w6246 = (w2641 & w3952) | (w2641 & ~w307) | (w3952 & ~w307);
assign w6247 = w3954 & w2646;
assign w6248 = (w2646 & w3954) | (w2646 & ~w886) | (w3954 & ~w886);
assign w6249 = w3956 & w2652;
assign w6250 = (w2652 & w3956) | (w2652 & ~w886) | (w3956 & ~w886);
assign w6251 = w3958 & w2657;
assign w6252 = (w2657 & w3958) | (w2657 & ~w307) | (w3958 & ~w307);
assign w6253 = w3960 & w2697;
assign w6254 = (w2697 & w3960) | (w2697 & ~w307) | (w3960 & ~w307);
assign w6255 = w3962 & w2702;
assign w6256 = (w2702 & w3962) | (w2702 & ~w886) | (w3962 & ~w886);
assign w6257 = w3964 & w2708;
assign w6258 = (w2708 & w3964) | (w2708 & ~w307) | (w3964 & ~w307);
assign w6259 = w3966 & w2713;
assign w6260 = (w2713 & w3966) | (w2713 & ~w886) | (w3966 & ~w886);
assign w6261 = w3968 & w2721;
assign w6262 = (w2721 & w3968) | (w2721 & ~w886) | (w3968 & ~w886);
assign w6263 = w3970 & w2726;
assign w6264 = (w2726 & w3970) | (w2726 & ~w307) | (w3970 & ~w307);
assign w6265 = ~w576 & ~w4231;
assign w6266 = ~w576 & ~w4232;
assign w6267 = ~w1155 & ~w4234;
assign w6268 = ~w1155 & ~w4235;
assign w6269 = ~w1161 & ~w4236;
assign w6270 = ~w1161 & ~w4237;
assign w6271 = ~w1166 & ~w4238;
assign w6272 = ~w1166 & ~w4239;
assign w6273 = ~w1174 & ~w4240;
assign w6274 = ~w1174 & ~w4241;
assign w6275 = ~w1179 & ~w4242;
assign w6276 = ~w1179 & ~w4243;
assign w6277 = ~w1196 & ~w4252;
assign w6278 = ~w1196 & ~w4253;
assign w6279 = ~w1201 & ~w4254;
assign w6280 = ~w1201 & ~w4255;
assign w6281 = ~w1218 & ~w4264;
assign w6282 = ~w1218 & ~w4265;
assign w6283 = ~w1223 & ~w4266;
assign w6284 = ~w1223 & ~w4267;
assign w6285 = ~w1236 & ~w4268;
assign w6286 = ~w1236 & ~w4269;
assign w6287 = ~w1241 & ~w4270;
assign w6288 = ~w1241 & ~w4271;
assign w6289 = ~w1247 & ~w4272;
assign w6290 = ~w1247 & ~w4273;
assign w6291 = ~w1252 & ~w4274;
assign w6292 = ~w1252 & ~w4275;
assign w6293 = ~w1260 & ~w4276;
assign w6294 = ~w1260 & ~w4277;
assign w6295 = ~w1265 & ~w4278;
assign w6296 = ~w1265 & ~w4279;
assign w6297 = ~w1273 & ~w4280;
assign w6298 = ~w1273 & ~w4281;
assign w6299 = ~w1278 & ~w4282;
assign w6300 = ~w1278 & ~w4283;
assign w6301 = ~w1284 & ~w4284;
assign w6302 = ~w1284 & ~w4285;
assign w6303 = ~w1289 & ~w4286;
assign w6304 = ~w1289 & ~w4287;
assign w6305 = ~w1297 & ~w4288;
assign w6306 = ~w1297 & ~w4289;
assign w6307 = ~w1302 & ~w4290;
assign w6308 = ~w1302 & ~w4291;
assign w6309 = ~w1311 & ~w4292;
assign w6310 = ~w1311 & ~w4293;
assign w6311 = ~w1316 & ~w4294;
assign w6312 = ~w1316 & ~w4295;
assign w6313 = ~w1322 & ~w4296;
assign w6314 = ~w1322 & ~w4297;
assign w6315 = ~w1327 & ~w4298;
assign w6316 = ~w1327 & ~w4299;
assign w6317 = ~w1335 & ~w4300;
assign w6318 = ~w1335 & ~w4301;
assign w6319 = ~w1340 & ~w4302;
assign w6320 = ~w1340 & ~w4303;
assign w6321 = ~w1363 & ~w4304;
assign w6322 = ~w1363 & ~w4305;
assign w6323 = ~w1368 & ~w4306;
assign w6324 = ~w1368 & ~w4307;
assign w6325 = ~w1374 & ~w4308;
assign w6326 = ~w1374 & ~w4309;
assign w6327 = ~w1379 & ~w4310;
assign w6328 = ~w1379 & ~w4311;
assign w6329 = ~w1387 & ~w4312;
assign w6330 = ~w1387 & ~w4313;
assign w6331 = ~w1392 & ~w4314;
assign w6332 = ~w1392 & ~w4315;
assign w6333 = ~w1407 & ~w4324;
assign w6334 = ~w1407 & ~w4325;
assign w6335 = ~w1412 & ~w4326;
assign w6336 = ~w1412 & ~w4327;
assign w6337 = ~w1433 & ~w4336;
assign w6338 = ~w1433 & ~w4337;
assign w6339 = ~w1438 & ~w4338;
assign w6340 = ~w1438 & ~w4339;
assign w6341 = ~w1621 & ~w4485;
assign w6342 = ~w1621 & ~w4486;
assign w6343 = ~w1626 & ~w4487;
assign w6344 = ~w1626 & ~w4488;
assign w6345 = ~w1632 & ~w4489;
assign w6346 = ~w1632 & ~w4490;
assign w6347 = ~w1637 & ~w4491;
assign w6348 = ~w1637 & ~w4492;
assign w6349 = ~w1643 & ~w4493;
assign w6350 = ~w1643 & ~w4494;
assign w6351 = ~w1648 & ~w4495;
assign w6352 = ~w1648 & ~w4496;
assign w6353 = ~w1850 & ~w4562;
assign w6354 = ~w1850 & ~w4563;
assign w6355 = ~w1855 & ~w4564;
assign w6356 = ~w1855 & ~w4565;
assign w6357 = ~w1861 & ~w4566;
assign w6358 = ~w1861 & ~w4567;
assign w6359 = ~w1866 & ~w4568;
assign w6360 = ~w1866 & ~w4569;
assign w6361 = ~w1874 & ~w4570;
assign w6362 = ~w1874 & ~w4571;
assign w6363 = ~w1879 & ~w4572;
assign w6364 = ~w1879 & ~w4573;
assign w6365 = ~w1888 & ~w4574;
assign w6366 = ~w1888 & ~w4575;
assign w6367 = ~w1893 & ~w4576;
assign w6368 = ~w1893 & ~w4577;
assign w6369 = ~w1899 & ~w4578;
assign w6370 = ~w1899 & ~w4579;
assign w6371 = ~w1904 & ~w4580;
assign w6372 = ~w1904 & ~w4581;
assign w6373 = ~w1931 & ~w4598;
assign w6374 = ~w1931 & ~w4599;
assign w6375 = ~w1936 & ~w4600;
assign w6376 = ~w1936 & ~w4601;
assign w6377 = ~w1966 & ~w4614;
assign w6378 = ~w1966 & ~w4615;
assign w6379 = ~w1971 & ~w4616;
assign w6380 = ~w1971 & ~w4617;
assign w6381 = ~w1977 & ~w4618;
assign w6382 = ~w1977 & ~w4619;
assign w6383 = ~w1982 & ~w4620;
assign w6384 = ~w1982 & ~w4621;
assign w6385 = ~w2011 & ~w4630;
assign w6386 = ~w2011 & ~w4631;
assign w6387 = ~w2016 & ~w4632;
assign w6388 = ~w2016 & ~w4633;
assign w6389 = ~w2031 & ~w4642;
assign w6390 = ~w2031 & ~w4643;
assign w6391 = ~w2036 & ~w4644;
assign w6392 = ~w2036 & ~w4645;
assign w6393 = ~w2105 & ~w4679;
assign w6394 = ~w2105 & ~w4680;
assign w6395 = ~w2110 & ~w4681;
assign w6396 = ~w2110 & ~w4682;
assign w6397 = ~w2116 & ~w4683;
assign w6398 = ~w2116 & ~w4684;
assign w6399 = ~w2121 & ~w4685;
assign w6400 = ~w2121 & ~w4686;
assign w6401 = ~w2132 & ~w4687;
assign w6402 = ~w2132 & ~w4688;
assign w6403 = ~w2137 & ~w4689;
assign w6404 = ~w2137 & ~w4690;
assign w6405 = ~w2143 & ~w4691;
assign w6406 = ~w2143 & ~w4692;
assign w6407 = ~w2148 & ~w4693;
assign w6408 = ~w2148 & ~w4694;
assign w6409 = ~w2155 & ~w4695;
assign w6410 = ~w2155 & ~w4696;
assign w6411 = ~w2160 & ~w4697;
assign w6412 = ~w2160 & ~w4698;
assign w6413 = ~w2387 & ~w4787;
assign w6414 = ~w2387 & ~w4788;
assign w6415 = ~w2392 & ~w4789;
assign w6416 = ~w2392 & ~w4790;
assign w6417 = ~w2399 & ~w4791;
assign w6418 = ~w2399 & ~w4792;
assign w6419 = ~w2404 & ~w4793;
assign w6420 = ~w2404 & ~w4794;
assign w6421 = ~w2431 & ~w4811;
assign w6422 = ~w2431 & ~w4812;
assign w6423 = ~w2436 & ~w4813;
assign w6424 = ~w2436 & ~w4814;
assign w6425 = ~w2442 & ~w4815;
assign w6426 = ~w2442 & ~w4816;
assign w6427 = ~w2447 & ~w4817;
assign w6428 = ~w2447 & ~w4818;
assign w6429 = ~w2455 & ~w4819;
assign w6430 = ~w2455 & ~w4820;
assign w6431 = ~w2460 & ~w4821;
assign w6432 = ~w2460 & ~w4822;
assign w6433 = ~w2542 & ~w4840;
assign w6434 = ~w2542 & ~w4841;
assign w6435 = ~w2547 & ~w4842;
assign w6436 = ~w2547 & ~w4843;
assign w6437 = ~w2553 & ~w4844;
assign w6438 = ~w2553 & ~w4845;
assign w6439 = ~w2558 & ~w4846;
assign w6440 = ~w2558 & ~w4847;
assign w6441 = ~w571 & in0_8;
assign w6442 = w571 & in1_9;
assign w6443 = ~w571 & in0_9;
assign w6444 = w1150 & in3_9;
assign w6445 = ~w1150 & in2_9;
assign w6446 = w571 & in1_7;
assign w6447 = ~w571 & in0_7;
assign w6448 = w1150 & in3_7;
assign w6449 = ~w1150 & in2_7;
assign w6450 = w571 & in1_19;
assign w6451 = ~w571 & in0_19;
assign w6452 = w1150 & in3_19;
assign w6453 = ~w1150 & in2_19;
assign w6454 = w571 & in1_18;
assign w6455 = ~w571 & in0_18;
assign w6456 = w1150 & in3_18;
assign w6457 = ~w1150 & in2_18;
assign w6458 = w571 & in1_20;
assign w6459 = ~w571 & in0_20;
assign w6460 = w1150 & in3_20;
assign w6461 = ~w1150 & in2_20;
assign w6462 = w571 & in1_22;
assign w6463 = ~w571 & in0_22;
assign w6464 = w1150 & in3_22;
assign w6465 = ~w1150 & in2_22;
assign w6466 = w1150 & in3_17;
assign w6467 = ~w1150 & in2_17;
assign w6468 = w571 & in1_17;
assign w6469 = ~w571 & in0_17;
assign w6470 = w1150 & in3_32;
assign w6471 = ~w1150 & in2_32;
assign w6472 = w571 & in1_32;
assign w6473 = ~w571 & in0_32;
assign w6474 = w571 & in1_33;
assign w6475 = ~w571 & in0_33;
assign w6476 = w1150 & in3_33;
assign w6477 = ~w1150 & in2_33;
assign w6478 = w1150 & in3_34;
assign w6479 = ~w1150 & in2_34;
assign w6480 = w571 & in1_34;
assign w6481 = ~w571 & in0_34;
assign w6482 = w571 & in1_55;
assign w6483 = ~w571 & in0_55;
assign w6484 = w1150 & in3_55;
assign w6485 = ~w1150 & in2_55;
assign w6486 = w1150 & in3_54;
assign w6487 = ~w1150 & in2_54;
assign w6488 = w571 & in1_54;
assign w6489 = ~w571 & in0_54;
assign w6490 = w571 & in1_52;
assign w6491 = ~w571 & in0_52;
assign w6492 = w1150 & in3_52;
assign w6493 = ~w1150 & in2_52;
assign w6494 = w571 & in1_51;
assign w6495 = ~w571 & in0_51;
assign w6496 = w1150 & in3_51;
assign w6497 = ~w1150 & in2_51;
assign w6498 = w571 & in1_53;
assign w6499 = ~w571 & in0_53;
assign w6500 = w1150 & in3_53;
assign w6501 = ~w1150 & in2_53;
assign w6502 = w571 & in1_49;
assign w6503 = ~w571 & in0_49;
assign w6504 = w1150 & in3_49;
assign w6505 = ~w1150 & in2_49;
assign w6506 = w1150 & in3_48;
assign w6507 = ~w1150 & in2_48;
assign w6508 = w571 & in1_48;
assign w6509 = ~w571 & in0_48;
assign w6510 = w1150 & in3_50;
assign w6511 = ~w1150 & in2_50;
assign w6512 = w571 & in1_50;
assign w6513 = ~w571 & in0_50;
assign w6514 = w571 & in1_57;
assign w6515 = ~w571 & in0_57;
assign w6516 = w1150 & in3_57;
assign w6517 = ~w1150 & in2_57;
assign w6518 = w571 & in1_56;
assign w6519 = ~w571 & in0_56;
assign w6520 = w1150 & in3_56;
assign w6521 = ~w1150 & in2_56;
assign w6522 = w571 & in1_58;
assign w6523 = ~w571 & in0_58;
assign w6524 = w1150 & in3_58;
assign w6525 = ~w1150 & in2_58;
assign w6526 = w571 & in1_60;
assign w6527 = ~w571 & in0_60;
assign w6528 = w1150 & in3_60;
assign w6529 = ~w1150 & in2_60;
assign w6530 = w571 & in1_59;
assign w6531 = ~w571 & in0_59;
assign w6532 = w1150 & in3_59;
assign w6533 = ~w1150 & in2_59;
assign w6534 = w571 & in1_61;
assign w6535 = ~w571 & in0_61;
assign w6536 = w1150 & in3_61;
assign w6537 = ~w1150 & in2_61;
assign w6538 = w1150 & in3_66;
assign w6539 = ~w1150 & in2_66;
assign w6540 = w571 & in1_66;
assign w6541 = ~w571 & in0_66;
assign w6542 = w571 & in1_65;
assign w6543 = ~w571 & in0_65;
assign w6544 = w1150 & in3_65;
assign w6545 = ~w1150 & in2_65;
assign w6546 = w1150 & in3_64;
assign w6547 = ~w1150 & in2_64;
assign w6548 = w571 & in1_64;
assign w6549 = ~w571 & in0_64;
assign w6550 = w571 & in1_69;
assign w6551 = ~w571 & in0_69;
assign w6552 = w1150 & in3_69;
assign w6553 = ~w1150 & in2_69;
assign w6554 = w1150 & in3_70;
assign w6555 = ~w1150 & in2_70;
assign w6556 = w571 & in1_70;
assign w6557 = ~w571 & in0_70;
assign w6558 = ~w572 & in0_82;
assign w6559 = w572 & in1_82;
assign w6560 = ~w1151 & in2_82;
assign w6561 = w1151 & in3_82;
assign w6562 = w571 & in1_91;
assign w6563 = ~w571 & in0_91;
assign w6564 = w1150 & in3_91;
assign w6565 = ~w1150 & in2_91;
assign w6566 = w1150 & in3_90;
assign w6567 = ~w1150 & in2_90;
assign w6568 = w571 & in1_90;
assign w6569 = ~w571 & in0_90;
assign w6570 = w1150 & in3_86;
assign w6571 = ~w1150 & in2_86;
assign w6572 = w571 & in1_86;
assign w6573 = ~w571 & in0_86;
assign w6574 = w571 & in1_85;
assign w6575 = ~w571 & in0_85;
assign w6576 = w1150 & in3_85;
assign w6577 = ~w1150 & in2_85;
assign w6578 = w571 & in1_84;
assign w6579 = ~w571 & in0_84;
assign w6580 = w1150 & in3_84;
assign w6581 = ~w1150 & in2_84;
assign w6582 = ~w572 & in0_81;
assign w6583 = w572 & in1_81;
assign w6584 = ~w1151 & in2_81;
assign w6585 = w1151 & in3_81;
assign w6586 = ~w572 & in0_80;
assign w6587 = w572 & in1_80;
assign w6588 = ~w1151 & in2_80;
assign w6589 = w1151 & in3_80;
assign w6590 = w571 & in1_77;
assign w6591 = ~w571 & in0_77;
assign w6592 = w1150 & in3_77;
assign w6593 = ~w1150 & in2_77;
assign w6594 = w1150 & in3_72;
assign w6595 = ~w1150 & in2_72;
assign w6596 = w571 & in1_72;
assign w6597 = ~w571 & in0_72;
assign w6598 = w571 & in1_73;
assign w6599 = ~w571 & in0_73;
assign w6600 = w1150 & in3_73;
assign w6601 = ~w1150 & in2_73;
assign w6602 = w571 & in1_75;
assign w6603 = ~w571 & in0_75;
assign w6604 = w1150 & in3_75;
assign w6605 = ~w1150 & in2_75;
assign w6606 = w571 & in1_76;
assign w6607 = ~w571 & in0_76;
assign w6608 = w1150 & in3_76;
assign w6609 = ~w1150 & in2_76;
assign w6610 = w1150 & in3_74;
assign w6611 = ~w1150 & in2_74;
assign w6612 = w571 & in1_74;
assign w6613 = ~w571 & in0_74;
assign w6614 = w1150 & in3_118;
assign w6615 = ~w1150 & in2_118;
assign w6616 = w571 & in1_118;
assign w6617 = ~w571 & in0_118;
assign w6618 = w571 & in1_117;
assign w6619 = ~w571 & in0_117;
assign w6620 = w1150 & in3_117;
assign w6621 = ~w1150 & in2_117;
assign w6622 = ~w572 & in0_123;
assign w6623 = w572 & in1_123;
assign w6624 = ~w1151 & in2_123;
assign w6625 = w1151 & in3_123;
assign w6626 = ~w1151 & in2_122;
assign w6627 = w1151 & in3_122;
assign w6628 = ~w572 & in0_122;
assign w6629 = w572 & in1_122;
assign w6630 = ~w572 & in0_121;
assign w6631 = w572 & in1_121;
assign w6632 = ~w1151 & in2_121;
assign w6633 = w1151 & in3_121;
assign w6634 = ~w1151 & in2_120;
assign w6635 = w1151 & in3_120;
assign w6636 = ~w572 & in0_120;
assign w6637 = w572 & in1_120;
assign w6638 = w571 & in1_115;
assign w6639 = ~w571 & in0_115;
assign w6640 = w1150 & in3_115;
assign w6641 = ~w1150 & in2_115;
assign w6642 = w1150 & in3_114;
assign w6643 = ~w1150 & in2_114;
assign w6644 = w571 & in1_114;
assign w6645 = ~w571 & in0_114;
assign w6646 = w571 & in1_109;
assign w6647 = ~w571 & in0_109;
assign w6648 = w1150 & in3_109;
assign w6649 = ~w1150 & in2_109;
assign w6650 = w1150 & in3_110;
assign w6651 = ~w1150 & in2_110;
assign w6652 = w571 & in1_110;
assign w6653 = ~w571 & in0_110;
assign w6654 = w571 & in1_108;
assign w6655 = ~w571 & in0_108;
assign w6656 = w1150 & in3_108;
assign w6657 = ~w1150 & in2_108;
assign w6658 = in3_127 & in2_127;
assign w6659 = w1150 & in3_102;
assign w6660 = ~w1150 & in2_102;
assign w6661 = w571 & in1_102;
assign w6662 = ~w571 & in0_102;
assign w6663 = w571 & in1_101;
assign w6664 = ~w571 & in0_101;
assign w6665 = w1150 & in3_101;
assign w6666 = ~w1150 & in2_101;
assign w6667 = w1150 & in3_98;
assign w6668 = ~w1150 & in2_98;
assign w6669 = w571 & in1_98;
assign w6670 = ~w571 & in0_98;
assign w6671 = w571 & in1_97;
assign w6672 = ~w571 & in0_97;
assign w6673 = w1150 & in3_97;
assign w6674 = ~w1150 & in2_97;
assign w6675 = w1150 & in3_96;
assign w6676 = ~w1150 & in2_96;
assign w6677 = w571 & in1_96;
assign w6678 = ~w571 & in0_96;
assign w6679 = w1150 & in3_106;
assign w6680 = ~w1150 & in2_106;
assign w6681 = w571 & in1_106;
assign w6682 = ~w571 & in0_106;
assign w6683 = w571 & in1_105;
assign w6684 = ~w571 & in0_105;
assign w6685 = w1150 & in3_105;
assign w6686 = ~w1150 & in2_105;
assign w6687 = w1150 & in3_104;
assign w6688 = ~w1150 & in2_104;
assign w6689 = w571 & in1_104;
assign w6690 = ~w571 & in0_104;
assign w6691 = w571 & in1_92;
assign w6692 = ~w571 & in0_92;
assign w6693 = w1150 & in3_92;
assign w6694 = ~w1150 & in2_92;
assign w6695 = w571 & in1_93;
assign w6696 = ~w571 & in0_93;
assign w6697 = w1150 & in3_93;
assign w6698 = ~w1150 & in2_93;
assign w6699 = w1150 & in3_94;
assign w6700 = ~w1150 & in2_94;
assign w6701 = w571 & in1_94;
assign w6702 = ~w571 & in0_94;
assign w6703 = w4936 & ~w544;
assign w6704 = w4955 & ~w1104;
assign w6705 = w4957 & ~w1104;
assign w6706 = w4959 & ~w544;
assign w6707 = w4961 & ~w544;
assign w6708 = w4963 & ~w1104;
assign w6709 = w572 & ~w544;
assign w6710 = w1151 & ~w1104;
assign w6711 = w4965 & ~w544;
assign w6712 = w4967 & ~w1104;
assign w6713 = w4969 & ~w544;
assign w6714 = w4971 & ~w1104;
assign w6715 = w4973 & ~w544;
assign w6716 = w4975 & ~w1104;
assign w6717 = w4977 & ~w544;
assign w6718 = w4979 & ~w1104;
assign w6719 = w4981 & ~w544;
assign w6720 = w4983 & ~w1104;
assign w6721 = w4985 & ~w544;
assign w6722 = w4987 & ~w1104;
assign w6723 = w4989 & ~w544;
assign w6724 = w4991 & ~w1104;
assign w6725 = w4993 & ~w544;
assign w6726 = w4995 & ~w1104;
assign w6727 = w4997 & ~w1104;
assign w6728 = w4999 & ~w544;
assign w6729 = w5001 & ~w544;
assign w6730 = w5003 & ~w1104;
assign w6731 = w5005 & ~w544;
assign w6732 = w5007 & ~w1104;
assign w6733 = w5009 & ~w544;
assign w6734 = w5011 & ~w1104;
assign w6735 = w5013 & ~w544;
assign w6736 = w5015 & ~w1104;
assign w6737 = w5017 & ~w544;
assign w6738 = w5019 & ~w1104;
assign w6739 = w5021 & ~w544;
assign w6740 = w5023 & ~w1104;
assign w6741 = w5025 & ~w1104;
assign w6742 = w5027 & ~w544;
assign w6743 = w5029 & ~w1104;
assign w6744 = w5031 & ~w544;
assign w6745 = w5033 & ~w544;
assign w6746 = w5035 & ~w1104;
assign w6747 = w5037 & ~w1104;
assign w6748 = w5039 & ~w544;
assign w6749 = w5041 & ~w544;
assign w6750 = w5043 & ~w1104;
assign w6751 = w5045 & ~w1104;
assign w6752 = w5047 & ~w544;
assign w6753 = w5049 & ~w544;
assign w6754 = w5051 & ~w1104;
assign w6755 = w5053 & ~w544;
assign w6756 = w5055 & ~w1104;
assign w6757 = w5057 & ~w544;
assign w6758 = w5059 & ~w1104;
assign w6759 = w5061 & ~w544;
assign w6760 = w5063 & ~w1104;
assign w6761 = w5065 & ~w1104;
assign w6762 = w5067 & ~w544;
assign w6763 = w5069 & ~w1104;
assign w6764 = w5071 & ~w544;
assign w6765 = w5073 & ~w544;
assign w6766 = w5075 & ~w1104;
assign w6767 = w5077 & ~w544;
assign w6768 = w5079 & ~w1104;
assign w6769 = w5081 & ~w544;
assign w6770 = w5083 & ~w1104;
assign w6771 = w5085 & ~w544;
assign w6772 = w5087 & ~w1104;
assign w6773 = w5089 & ~w544;
assign w6774 = w5091 & ~w1104;
assign w6775 = w5093 & ~w544;
assign w6776 = w5095 & ~w1104;
assign w6777 = w5097 & ~w1104;
assign w6778 = w5099 & ~w544;
assign w6779 = w5101 & ~w544;
assign w6780 = w5103 & ~w1104;
assign w6781 = w5105 & ~w1104;
assign w6782 = w5107 & ~w544;
assign w6783 = w5109 & ~w544;
assign w6784 = w5111 & ~w1104;
assign w6785 = w5113 & ~w1104;
assign w6786 = w5115 & ~w544;
assign w6787 = w5129 & ~w544;
assign w6788 = w5131 & ~w1104;
assign w6789 = w5133 & ~w1104;
assign w6790 = w5135 & ~w544;
assign w6791 = w5137 & ~w1104;
assign w6792 = w5139 & ~w544;
assign w6793 = w5141 & ~w544;
assign w6794 = w5143 & ~w1104;
assign w6795 = w5145 & ~w544;
assign w6796 = w5147 & ~w1104;
assign w6797 = w5165 & ~w544;
assign w6798 = w5167 & ~w1104;
assign w6799 = w5169 & ~w1104;
assign w6800 = w5171 & ~w544;
assign w6801 = w5173 & ~w544;
assign w6802 = w5175 & ~w1104;
assign w6803 = w5177 & ~w544;
assign w6804 = w5179 & ~w1104;
assign w6805 = w5181 & ~w544;
assign w6806 = w5183 & ~w1104;
assign w6807 = w5185 & ~w1104;
assign w6808 = w5187 & ~w544;
assign w6809 = w5189 & ~w1104;
assign w6810 = w5191 & ~w544;
assign w6811 = w5193 & ~w544;
assign w6812 = w5195 & ~w1104;
assign w6813 = w5232 & ~w544;
assign w6814 = w5234 & ~w1104;
assign w6815 = w5236 & ~w1104;
assign w6816 = w5238 & ~w544;
assign w6817 = w5240 & ~w544;
assign w6818 = w5242 & ~w1104;
assign w6819 = w5244 & ~w1104;
assign w6820 = w5246 & ~w544;
assign w6821 = w5248 & ~w544;
assign w6822 = w5250 & ~w1104;
assign w6823 = w5257 & ~w1104;
assign w6824 = w5259 & ~w544;
assign w6825 = w5261 & ~w544;
assign w6826 = w5263 & ~w1104;
assign w6827 = w5266 & ~w1104;
assign w6828 = w5268 & ~w544;
assign w6829 = w5270 & ~w544;
assign w6830 = w5272 & ~w1104;
assign w6831 = w5274 & ~w1104;
assign w6832 = w5276 & ~w544;
assign w6833 = w5278 & ~w1104;
assign w6834 = w5280 & ~w544;
assign w6835 = w5282 & ~w544;
assign w6836 = w5284 & ~w1104;
assign w6837 = w5286 & ~w1104;
assign w6838 = w5288 & ~w544;
assign w6839 = w5290 & ~w544;
assign w6840 = w5292 & ~w1104;
assign w6841 = w5294 & ~w544;
assign w6842 = w5296 & ~w1104;
assign w6843 = w5298 & ~w1104;
assign w6844 = w5300 & ~w544;
assign w6845 = ~w571 & in0_3;
assign w6846 = w571 & in1_3;
assign w6847 = ~w1150 & in2_3;
assign w6848 = w1150 & in3_3;
assign w6849 = ~w571 & in0_5;
assign w6850 = w571 & in1_5;
assign w6851 = ~w1150 & in2_5;
assign w6852 = w1150 & in3_5;
assign w6853 = ~w571 & in0_21;
assign w6854 = w571 & in1_21;
assign w6855 = ~w1150 & in2_21;
assign w6856 = w1150 & in3_21;
assign w6857 = ~w571 & in0_16;
assign w6858 = w571 & in1_16;
assign w6859 = ~w1150 & in2_16;
assign w6860 = w1150 & in3_16;
assign w6861 = ~w571 & in0_27;
assign w6862 = w571 & in1_27;
assign w6863 = ~w1150 & in2_27;
assign w6864 = w3682 & ~w576;
assign w6865 = (~w576 & w3682) | (~w576 & ~w307) | (w3682 & ~w307);
assign w6866 = w3693 & ~w1155;
assign w6867 = (~w1155 & w3693) | (~w1155 & ~w886) | (w3693 & ~w886);
assign w6868 = w3695 & ~w1161;
assign w6869 = (~w1161 & w3695) | (~w1161 & ~w886) | (w3695 & ~w886);
assign w6870 = w3697 & ~w1166;
assign w6871 = (~w1166 & w3697) | (~w1166 & ~w307) | (w3697 & ~w307);
assign w6872 = w3699 & ~w1174;
assign w6873 = (~w1174 & w3699) | (~w1174 & ~w307) | (w3699 & ~w307);
assign w6874 = w3701 & ~w1179;
assign w6875 = (~w1179 & w3701) | (~w1179 & ~w886) | (w3701 & ~w886);
assign w6876 = w3705 & ~w1196;
assign w6877 = (~w1196 & w3705) | (~w1196 & ~w307) | (w3705 & ~w307);
assign w6878 = w3707 & ~w1201;
assign w6879 = (~w1201 & w3707) | (~w1201 & ~w886) | (w3707 & ~w886);
assign w6880 = w3709 & ~w1218;
assign w6881 = (~w1218 & w3709) | (~w1218 & ~w307) | (w3709 & ~w307);
assign w6882 = w3711 & ~w1223;
assign w6883 = (~w1223 & w3711) | (~w1223 & ~w886) | (w3711 & ~w886);
assign w6884 = w3713 & ~w1236;
assign w6885 = (~w1236 & w3713) | (~w1236 & ~w307) | (w3713 & ~w307);
assign w6886 = w3715 & ~w1241;
assign w6887 = (~w1241 & w3715) | (~w1241 & ~w886) | (w3715 & ~w886);
assign w6888 = w3717 & ~w1247;
assign w6889 = (~w1247 & w3717) | (~w1247 & ~w307) | (w3717 & ~w307);
assign w6890 = w3719 & ~w1252;
assign w6891 = (~w1252 & w3719) | (~w1252 & ~w886) | (w3719 & ~w886);
assign w6892 = w3721 & ~w1260;
assign w6893 = (~w1260 & w3721) | (~w1260 & ~w307) | (w3721 & ~w307);
assign w6894 = w3723 & ~w1265;
assign w6895 = (~w1265 & w3723) | (~w1265 & ~w886) | (w3723 & ~w886);
assign w6896 = w3725 & ~w1273;
assign w6897 = (~w1273 & w3725) | (~w1273 & ~w307) | (w3725 & ~w307);
assign w6898 = w3727 & ~w1278;
assign w6899 = (~w1278 & w3727) | (~w1278 & ~w886) | (w3727 & ~w886);
assign w6900 = w3729 & ~w1284;
assign w6901 = (~w1284 & w3729) | (~w1284 & ~w307) | (w3729 & ~w307);
assign w6902 = w3731 & ~w1289;
assign w6903 = (~w1289 & w3731) | (~w1289 & ~w886) | (w3731 & ~w886);
assign w6904 = w3733 & ~w1297;
assign w6905 = (~w1297 & w3733) | (~w1297 & ~w307) | (w3733 & ~w307);
assign w6906 = w3735 & ~w1302;
assign w6907 = (~w1302 & w3735) | (~w1302 & ~w886) | (w3735 & ~w886);
assign w6908 = w3737 & ~w1311;
assign w6909 = (~w1311 & w3737) | (~w1311 & ~w886) | (w3737 & ~w886);
assign w6910 = w3739 & ~w1316;
assign w6911 = (~w1316 & w3739) | (~w1316 & ~w307) | (w3739 & ~w307);
assign w6912 = w3741 & ~w1322;
assign w6913 = (~w1322 & w3741) | (~w1322 & ~w307) | (w3741 & ~w307);
assign w6914 = w3743 & ~w1327;
assign w6915 = (~w1327 & w3743) | (~w1327 & ~w886) | (w3743 & ~w886);
assign w6916 = w3745 & ~w1335;
assign w6917 = (~w1335 & w3745) | (~w1335 & ~w307) | (w3745 & ~w307);
assign w6918 = w3747 & ~w1340;
assign w6919 = (~w1340 & w3747) | (~w1340 & ~w886) | (w3747 & ~w886);
assign w6920 = w3749 & ~w1363;
assign w6921 = (~w1363 & w3749) | (~w1363 & ~w307) | (w3749 & ~w307);
assign w6922 = w3751 & ~w1368;
assign w6923 = (~w1368 & w3751) | (~w1368 & ~w886) | (w3751 & ~w886);
assign w6924 = w3753 & ~w1374;
assign w6925 = (~w1374 & w3753) | (~w1374 & ~w307) | (w3753 & ~w307);
assign w6926 = w3755 & ~w1379;
assign w6927 = (~w1379 & w3755) | (~w1379 & ~w886) | (w3755 & ~w886);
assign w6928 = w3757 & ~w1387;
assign w6929 = (~w1387 & w3757) | (~w1387 & ~w307) | (w3757 & ~w307);
assign w6930 = w3759 & ~w1392;
assign w6931 = (~w1392 & w3759) | (~w1392 & ~w886) | (w3759 & ~w886);
assign w6932 = w3761 & ~w1407;
assign w6933 = (~w1407 & w3761) | (~w1407 & ~w307) | (w3761 & ~w307);
assign w6934 = w3763 & ~w1412;
assign w6935 = (~w1412 & w3763) | (~w1412 & ~w886) | (w3763 & ~w886);
assign w6936 = w3765 & ~w1433;
assign w6937 = (~w1433 & w3765) | (~w1433 & ~w886) | (w3765 & ~w886);
assign w6938 = w3767 & ~w1438;
assign w6939 = (~w1438 & w3767) | (~w1438 & ~w307) | (w3767 & ~w307);
assign w6940 = w3769 & ~w1621;
assign w6941 = (~w1621 & w3769) | (~w1621 & ~w886) | (w3769 & ~w886);
assign w6942 = w3771 & ~w1626;
assign w6943 = (~w1626 & w3771) | (~w1626 & ~w307) | (w3771 & ~w307);
assign w6944 = w3773 & ~w1632;
assign w6945 = (~w1632 & w3773) | (~w1632 & ~w307) | (w3773 & ~w307);
assign w6946 = w3775 & ~w1637;
assign w6947 = (~w1637 & w3775) | (~w1637 & ~w886) | (w3775 & ~w886);
assign w6948 = w3777 & ~w1643;
assign w6949 = (~w1643 & w3777) | (~w1643 & ~w886) | (w3777 & ~w886);
assign w6950 = w3779 & ~w1648;
assign w6951 = (~w1648 & w3779) | (~w1648 & ~w307) | (w3779 & ~w307);
assign w6952 = w3813 & ~w1850;
assign w6953 = (~w1850 & w3813) | (~w1850 & ~w307) | (w3813 & ~w307);
assign w6954 = w3815 & ~w1855;
assign w6955 = (~w1855 & w3815) | (~w1855 & ~w886) | (w3815 & ~w886);
assign w6956 = w3817 & ~w1861;
assign w6957 = (~w1861 & w3817) | (~w1861 & ~w307) | (w3817 & ~w307);
assign w6958 = w3819 & ~w1866;
assign w6959 = (~w1866 & w3819) | (~w1866 & ~w886) | (w3819 & ~w886);
assign w6960 = w3821 & ~w1874;
assign w6961 = (~w1874 & w3821) | (~w1874 & ~w307) | (w3821 & ~w307);
assign w6962 = w3823 & ~w1879;
assign w6963 = (~w1879 & w3823) | (~w1879 & ~w886) | (w3823 & ~w886);
assign w6964 = w3825 & ~w1888;
assign w6965 = (~w1888 & w3825) | (~w1888 & ~w307) | (w3825 & ~w307);
assign w6966 = w3827 & ~w1893;
assign w6967 = (~w1893 & w3827) | (~w1893 & ~w886) | (w3827 & ~w886);
assign w6968 = w3829 & ~w1899;
assign w6969 = (~w1899 & w3829) | (~w1899 & ~w307) | (w3829 & ~w307);
assign w6970 = w3831 & ~w1904;
assign w6971 = (~w1904 & w3831) | (~w1904 & ~w886) | (w3831 & ~w886);
assign w6972 = w3833 & ~w1931;
assign w6973 = (~w1931 & w3833) | (~w1931 & ~w307) | (w3833 & ~w307);
assign w6974 = w3835 & ~w1936;
assign w6975 = (~w1936 & w3835) | (~w1936 & ~w886) | (w3835 & ~w886);
assign w6976 = w3841 & ~w1966;
assign w6977 = (~w1966 & w3841) | (~w1966 & ~w307) | (w3841 & ~w307);
assign w6978 = w3843 & ~w1971;
assign w6979 = (~w1971 & w3843) | (~w1971 & ~w886) | (w3843 & ~w886);
assign w6980 = w3845 & ~w1977;
assign w6981 = (~w1977 & w3845) | (~w1977 & ~w886) | (w3845 & ~w886);
assign w6982 = w3847 & ~w1982;
assign w6983 = (~w1982 & w3847) | (~w1982 & ~w307) | (w3847 & ~w307);
assign w6984 = w3849 & ~w2011;
assign w6985 = (~w2011 & w3849) | (~w2011 & ~w307) | (w3849 & ~w307);
assign w6986 = w3851 & ~w2016;
assign w6987 = (~w2016 & w3851) | (~w2016 & ~w886) | (w3851 & ~w886);
assign w6988 = w3853 & ~w2031;
assign w6989 = (~w2031 & w3853) | (~w2031 & ~w886) | (w3853 & ~w886);
assign w6990 = w3855 & ~w2036;
assign w6991 = (~w2036 & w3855) | (~w2036 & ~w307) | (w3855 & ~w307);
assign w6992 = w3857 & ~w2105;
assign w6993 = (~w2105 & w3857) | (~w2105 & ~w307) | (w3857 & ~w307);
assign w6994 = w3859 & ~w2110;
assign w6995 = (~w2110 & w3859) | (~w2110 & ~w886) | (w3859 & ~w886);
assign w6996 = w3861 & ~w2116;
assign w6997 = (~w2116 & w3861) | (~w2116 & ~w886) | (w3861 & ~w886);
assign w6998 = w3863 & ~w2121;
assign w6999 = (~w2121 & w3863) | (~w2121 & ~w307) | (w3863 & ~w307);
assign w7000 = w3865 & ~w2132;
assign w7001 = (~w2132 & w3865) | (~w2132 & ~w886) | (w3865 & ~w886);
assign w7002 = w3867 & ~w2137;
assign w7003 = (~w2137 & w3867) | (~w2137 & ~w307) | (w3867 & ~w307);
assign w7004 = w3869 & ~w2143;
assign w7005 = (~w2143 & w3869) | (~w2143 & ~w307) | (w3869 & ~w307);
assign w7006 = w3871 & ~w2148;
assign w7007 = (~w2148 & w3871) | (~w2148 & ~w886) | (w3871 & ~w886);
assign w7008 = w3873 & ~w2155;
assign w7009 = (~w2155 & w3873) | (~w2155 & ~w307) | (w3873 & ~w307);
assign w7010 = w3875 & ~w2160;
assign w7011 = (~w2160 & w3875) | (~w2160 & ~w886) | (w3875 & ~w886);
assign w7012 = w3909 & ~w2387;
assign w7013 = (~w2387 & w3909) | (~w2387 & ~w307) | (w3909 & ~w307);
assign w7014 = w3911 & ~w2392;
assign w7015 = (~w2392 & w3911) | (~w2392 & ~w886) | (w3911 & ~w886);
assign w7016 = w3913 & ~w2399;
assign w7017 = (~w2399 & w3913) | (~w2399 & ~w886) | (w3913 & ~w886);
assign w7018 = w3915 & ~w2404;
assign w7019 = (~w2404 & w3915) | (~w2404 & ~w307) | (w3915 & ~w307);
assign w7020 = w3917 & ~w2431;
assign w7021 = (~w2431 & w3917) | (~w2431 & ~w307) | (w3917 & ~w307);
assign w7022 = w3919 & ~w2436;
assign w7023 = (~w2436 & w3919) | (~w2436 & ~w886) | (w3919 & ~w886);
assign w7024 = w3921 & ~w2442;
assign w7025 = (~w2442 & w3921) | (~w2442 & ~w886) | (w3921 & ~w886);
assign w7026 = w3923 & ~w2447;
assign w7027 = (~w2447 & w3923) | (~w2447 & ~w307) | (w3923 & ~w307);
assign w7028 = w3925 & ~w2455;
assign w7029 = (~w2455 & w3925) | (~w2455 & ~w307) | (w3925 & ~w307);
assign w7030 = w3927 & ~w2460;
assign w7031 = (~w2460 & w3927) | (~w2460 & ~w886) | (w3927 & ~w886);
assign w7032 = w3929 & ~w2542;
assign w7033 = (~w2542 & w3929) | (~w2542 & ~w886) | (w3929 & ~w886);
assign w7034 = w3931 & ~w2547;
assign w7035 = (~w2547 & w3931) | (~w2547 & ~w307) | (w3931 & ~w307);
assign w7036 = w3933 & ~w2553;
assign w7037 = (~w2553 & w3933) | (~w2553 & ~w307) | (w3933 & ~w307);
assign w7038 = w3935 & ~w2558;
assign w7039 = (~w2558 & w3935) | (~w2558 & ~w886) | (w3935 & ~w886);
assign w7040 = w3937 & ~w2582;
assign w7041 = (~w2582 & w3937) | (~w2582 & ~w886) | (w3937 & ~w886);
assign w7042 = w3939 & ~w2587;
assign w7043 = (~w2587 & w3939) | (~w2587 & ~w307) | (w3939 & ~w307);
assign w7044 = w3941 & ~w2594;
assign w7045 = (~w2594 & w3941) | (~w2594 & ~w307) | (w3941 & ~w307);
assign w7046 = w3943 & ~w2599;
assign w7047 = (~w2599 & w3943) | (~w2599 & ~w886) | (w3943 & ~w886);
assign w7048 = w3945 & ~w2605;
assign w7049 = (~w2605 & w3945) | (~w2605 & ~w886) | (w3945 & ~w886);
assign w7050 = w3947 & ~w2610;
assign w7051 = (~w2610 & w3947) | (~w2610 & ~w307) | (w3947 & ~w307);
assign w7052 = w3949 & ~w2631;
assign w7053 = (~w2631 & w3949) | (~w2631 & ~w886) | (w3949 & ~w886);
assign w7054 = w3951 & ~w2636;
assign w7055 = (~w2636 & w3951) | (~w2636 & ~w307) | (w3951 & ~w307);
assign w7056 = w3953 & ~w2643;
assign w7057 = (~w2643 & w3953) | (~w2643 & ~w307) | (w3953 & ~w307);
assign w7058 = w3955 & ~w2648;
assign w7059 = (~w2648 & w3955) | (~w2648 & ~w886) | (w3955 & ~w886);
assign w7060 = w3957 & ~w2654;
assign w7061 = (~w2654 & w3957) | (~w2654 & ~w886) | (w3957 & ~w886);
assign w7062 = w3959 & ~w2659;
assign w7063 = (~w2659 & w3959) | (~w2659 & ~w307) | (w3959 & ~w307);
assign w7064 = w3961 & ~w2699;
assign w7065 = (~w2699 & w3961) | (~w2699 & ~w307) | (w3961 & ~w307);
assign w7066 = w3963 & ~w2704;
assign w7067 = (~w2704 & w3963) | (~w2704 & ~w886) | (w3963 & ~w886);
assign w7068 = w3965 & ~w2710;
assign w7069 = (~w2710 & w3965) | (~w2710 & ~w307) | (w3965 & ~w307);
assign w7070 = w3967 & ~w2715;
assign w7071 = (~w2715 & w3967) | (~w2715 & ~w886) | (w3967 & ~w886);
assign w7072 = w3969 & ~w2723;
assign w7073 = (~w2723 & w3969) | (~w2723 & ~w886) | (w3969 & ~w886);
assign w7074 = w3971 & ~w2728;
assign w7075 = (~w2728 & w3971) | (~w2728 & ~w307) | (w3971 & ~w307);
assign w7076 = (~w2334 & w4225) | (~w2334 & w2505) | (w4225 & w2505);
assign w7077 = (~w2334 & w4225) | (~w2334 & w2484) | (w4225 & w2484);
assign w7078 = ~w2334 & w2484;
assign w7079 = w3781 & ~w1697;
assign w7080 = (~w1697 & w3781) | (~w1697 & ~w307) | (w3781 & ~w307);
assign w7081 = w3783 & ~w1702;
assign w7082 = (~w1702 & w3783) | (~w1702 & ~w886) | (w3783 & ~w886);
assign w7083 = w3785 & ~w1709;
assign w7084 = (~w1709 & w3785) | (~w1709 & ~w886) | (w3785 & ~w886);
assign w7085 = w3787 & ~w1714;
assign w7086 = (~w1714 & w3787) | (~w1714 & ~w307) | (w3787 & ~w307);
assign w7087 = w3789 & ~w1722;
assign w7088 = (~w1722 & w3789) | (~w1722 & ~w307) | (w3789 & ~w307);
assign w7089 = w3791 & ~w1727;
assign w7090 = (~w1727 & w3791) | (~w1727 & ~w886) | (w3791 & ~w886);
assign w7091 = w3793 & ~w1733;
assign w7092 = (~w1733 & w3793) | (~w1733 & ~w307) | (w3793 & ~w307);
assign w7093 = w3795 & ~w1738;
assign w7094 = (~w1738 & w3795) | (~w1738 & ~w886) | (w3795 & ~w886);
assign w7095 = w3797 & ~w1746;
assign w7096 = (~w1746 & w3797) | (~w1746 & ~w307) | (w3797 & ~w307);
assign w7097 = w3799 & ~w1751;
assign w7098 = (~w1751 & w3799) | (~w1751 & ~w886) | (w3799 & ~w886);
assign w7099 = w3801 & ~w1760;
assign w7100 = (~w1760 & w3801) | (~w1760 & ~w307) | (w3801 & ~w307);
assign w7101 = w3803 & ~w1765;
assign w7102 = (~w1765 & w3803) | (~w1765 & ~w886) | (w3803 & ~w886);
assign w7103 = w3805 & ~w1771;
assign w7104 = (~w1771 & w3805) | (~w1771 & ~w886) | (w3805 & ~w886);
assign w7105 = w3807 & ~w1776;
assign w7106 = (~w1776 & w3807) | (~w1776 & ~w307) | (w3807 & ~w307);
assign w7107 = w3809 & ~w1784;
assign w7108 = (~w1784 & w3809) | (~w1784 & ~w886) | (w3809 & ~w886);
assign w7109 = w3811 & ~w1789;
assign w7110 = (~w1789 & w3811) | (~w1789 & ~w307) | (w3811 & ~w307);
assign w7111 = w3837 & ~w1953;
assign w7112 = (~w1953 & w3837) | (~w1953 & ~w886) | (w3837 & ~w886);
assign w7113 = w3839 & ~w1958;
assign w7114 = (~w1958 & w3839) | (~w1958 & ~w307) | (w3839 & ~w307);
assign w7115 = w3877 & ~w2199;
assign w7116 = (~w2199 & w3877) | (~w2199 & ~w307) | (w3877 & ~w307);
assign w7117 = w3879 & ~w2204;
assign w7118 = (~w2204 & w3879) | (~w2204 & ~w886) | (w3879 & ~w886);
assign w7119 = w3881 & ~w2211;
assign w7120 = (~w2211 & w3881) | (~w2211 & ~w886) | (w3881 & ~w886);
assign w7121 = w3883 & ~w2216;
assign w7122 = (~w2216 & w3883) | (~w2216 & ~w307) | (w3883 & ~w307);
assign w7123 = w3885 & ~w2222;
assign w7124 = (~w2222 & w3885) | (~w2222 & ~w307) | (w3885 & ~w307);
assign w7125 = w3887 & ~w2227;
assign w7126 = (~w2227 & w3887) | (~w2227 & ~w886) | (w3887 & ~w886);
assign w7127 = w3889 & ~w2240;
assign w7128 = (~w2240 & w3889) | (~w2240 & ~w307) | (w3889 & ~w307);
assign w7129 = w3891 & ~w2245;
assign w7130 = (~w2245 & w3891) | (~w2245 & ~w886) | (w3891 & ~w886);
assign w7131 = w3893 & ~w2251;
assign w7132 = (~w2251 & w3893) | (~w2251 & ~w307) | (w3893 & ~w307);
assign w7133 = w3895 & ~w2256;
assign w7134 = (~w2256 & w3895) | (~w2256 & ~w886) | (w3895 & ~w886);
assign w7135 = w3897 & ~w2262;
assign w7136 = (~w2262 & w3897) | (~w2262 & ~w886) | (w3897 & ~w886);
assign w7137 = w3899 & ~w2267;
assign w7138 = (~w2267 & w3899) | (~w2267 & ~w307) | (w3899 & ~w307);
assign w7139 = w3901 & ~w2290;
assign w7140 = (~w2290 & w3901) | (~w2290 & ~w886) | (w3901 & ~w886);
assign w7141 = w3903 & ~w2295;
assign w7142 = (~w2295 & w3903) | (~w2295 & ~w307) | (w3903 & ~w307);
assign w7143 = w3905 & ~w2301;
assign w7144 = (~w2301 & w3905) | (~w2301 & ~w307) | (w3905 & ~w307);
assign w7145 = w3907 & ~w2306;
assign w7146 = (~w2306 & w3907) | (~w2306 & ~w886) | (w3907 & ~w886);
assign w7147 = (w398 & ~w4230) | (w398 & ~w553) | (~w4230 & ~w553);
assign w7148 = (w977 & ~w4233) | (w977 & ~w1132) | (~w4233 & ~w1132);
assign w7149 = (~w4530 & ~w4531) | (~w4530 & ~w537) | (~w4531 & ~w537);
assign w7150 = (~w4532 & ~w4533) | (~w4532 & ~w1123) | (~w4533 & ~w1123);
assign w7151 = (~w4534 & ~w4535) | (~w4534 & ~w1123) | (~w4535 & ~w1123);
assign w7152 = (~w4536 & ~w4537) | (~w4536 & ~w537) | (~w4537 & ~w537);
assign w7153 = (~w4538 & ~w4539) | (~w4538 & ~w537) | (~w4539 & ~w537);
assign w7154 = (~w4540 & ~w4541) | (~w4540 & ~w1123) | (~w4541 & ~w1123);
assign w7155 = (~w4542 & ~w4543) | (~w4542 & ~w537) | (~w4543 & ~w537);
assign w7156 = (~w4544 & ~w4545) | (~w4544 & ~w1123) | (~w4545 & ~w1123);
assign w7157 = (~w4546 & ~w4547) | (~w4546 & ~w537) | (~w4547 & ~w537);
assign w7158 = (~w4548 & ~w4549) | (~w4548 & ~w1123) | (~w4549 & ~w1123);
assign w7159 = (~w4550 & ~w4551) | (~w4550 & ~w537) | (~w4551 & ~w537);
assign w7160 = (~w4552 & ~w4553) | (~w4552 & ~w1123) | (~w4553 & ~w1123);
assign w7161 = (~w4554 & ~w4555) | (~w4554 & ~w1123) | (~w4555 & ~w1123);
assign w7162 = (~w4556 & ~w4557) | (~w4556 & ~w537) | (~w4557 & ~w537);
assign w7163 = (~w4558 & ~w4559) | (~w4558 & ~w1123) | (~w4559 & ~w1123);
assign w7164 = (~w4560 & ~w4561) | (~w4560 & ~w537) | (~w4561 & ~w537);
assign w7165 = (~w4610 & ~w4611) | (~w4610 & ~w1123) | (~w4611 & ~w1123);
assign w7166 = (~w4612 & ~w4613) | (~w4612 & ~w537) | (~w4613 & ~w537);
assign w7167 = (~w4707 & ~w4708) | (~w4707 & ~w537) | (~w4708 & ~w537);
assign w7168 = (~w4709 & ~w4710) | (~w4709 & ~w1123) | (~w4710 & ~w1123);
assign w7169 = (~w4711 & ~w4712) | (~w4711 & ~w1123) | (~w4712 & ~w1123);
assign w7170 = (~w4713 & ~w4714) | (~w4713 & ~w537) | (~w4714 & ~w537);
assign w7171 = (~w4715 & ~w4716) | (~w4715 & ~w537) | (~w4716 & ~w537);
assign w7172 = (~w4717 & ~w4718) | (~w4717 & ~w1123) | (~w4718 & ~w1123);
assign w7173 = (~w4727 & ~w4728) | (~w4727 & ~w537) | (~w4728 & ~w537);
assign w7174 = (~w4729 & ~w4730) | (~w4729 & ~w1123) | (~w4730 & ~w1123);
assign w7175 = (~w4731 & ~w4732) | (~w4731 & ~w537) | (~w4732 & ~w537);
assign w7176 = (~w4733 & ~w4734) | (~w4733 & ~w1123) | (~w4734 & ~w1123);
assign w7177 = (~w4735 & ~w4736) | (~w4735 & ~w1123) | (~w4736 & ~w1123);
assign w7178 = (~w4737 & ~w4738) | (~w4737 & ~w537) | (~w4738 & ~w537);
assign w7179 = (~w4747 & ~w4748) | (~w4747 & ~w1123) | (~w4748 & ~w1123);
assign w7180 = (~w4749 & ~w4750) | (~w4749 & ~w537) | (~w4750 & ~w537);
assign w7181 = (~w4751 & ~w4752) | (~w4751 & ~w537) | (~w4752 & ~w537);
assign w7182 = (~w4753 & ~w4754) | (~w4753 & ~w1123) | (~w4754 & ~w1123);
assign w7183 = (~w4864 & ~w4865) | (~w4864 & ~w1123) | (~w4865 & ~w1123);
assign w7184 = (~w4866 & ~w4867) | (~w4866 & ~w537) | (~w4867 & ~w537);
assign w7185 = (~w4868 & ~w4869) | (~w4868 & ~w537) | (~w4869 & ~w537);
assign w7186 = (~w4870 & ~w4871) | (~w4870 & ~w1123) | (~w4871 & ~w1123);
assign w7187 = (~w4872 & ~w4873) | (~w4872 & ~w1123) | (~w4873 & ~w1123);
assign w7188 = (~w4874 & ~w4875) | (~w4874 & ~w537) | (~w4875 & ~w537);
assign w7189 = (~w4885 & ~w4886) | (~w4885 & ~w1123) | (~w4886 & ~w1123);
assign w7190 = (~w4887 & ~w4888) | (~w4887 & ~w537) | (~w4888 & ~w537);
assign w7191 = (~w4889 & ~w4890) | (~w4889 & ~w537) | (~w4890 & ~w537);
assign w7192 = (~w4891 & ~w4892) | (~w4891 & ~w1123) | (~w4892 & ~w1123);
assign w7193 = (~w4893 & ~w4894) | (~w4893 & ~w1123) | (~w4894 & ~w1123);
assign w7194 = (~w4895 & ~w4896) | (~w4895 & ~w537) | (~w4896 & ~w537);
assign w7195 = (~w4906 & ~w4907) | (~w4906 & ~w537) | (~w4907 & ~w537);
assign w7196 = (~w4908 & ~w4909) | (~w4908 & ~w1123) | (~w4909 & ~w1123);
assign w7197 = (~w4910 & ~w4911) | (~w4910 & ~w537) | (~w4911 & ~w537);
assign w7198 = (~w4912 & ~w4913) | (~w4912 & ~w1123) | (~w4913 & ~w1123);
assign w7199 = (~w4914 & ~w4915) | (~w4914 & ~w1123) | (~w4915 & ~w1123);
assign w7200 = (~w4916 & ~w4917) | (~w4916 & ~w537) | (~w4917 & ~w537);
assign w7201 = (~w2384 & ~w2334) | (~w2384 & w7078) | (~w2334 & w7078);
assign one = 1;
assign result_0 = ~w2781;// level 27
assign result_1 = w2788;// level 27
assign result_2 = ~w2795;// level 27
assign result_3 = ~w2802;// level 27
assign result_4 = ~w2809;// level 27
assign result_5 = ~w2816;// level 27
assign result_6 = ~w2823;// level 27
assign result_7 = ~w2830;// level 27
assign result_8 = ~w2837;// level 27
assign result_9 = ~w2844;// level 27
assign result_10 = ~w2851;// level 27
assign result_11 = ~w2858;// level 27
assign result_12 = ~w2865;// level 27
assign result_13 = ~w2872;// level 27
assign result_14 = ~w2879;// level 27
assign result_15 = ~w2886;// level 27
assign result_16 = ~w2893;// level 27
assign result_17 = w2900;// level 27
assign result_18 = ~w2907;// level 27
assign result_19 = ~w2914;// level 27
assign result_20 = ~w2921;// level 27
assign result_21 = ~w2928;// level 27
assign result_22 = ~w2935;// level 27
assign result_23 = ~w2942;// level 27
assign result_24 = ~w2949;// level 27
assign result_25 = ~w2956;// level 27
assign result_26 = ~w2963;// level 27
assign result_27 = ~w2970;// level 27
assign result_28 = ~w2977;// level 27
assign result_29 = ~w2984;// level 27
assign result_30 = ~w2991;// level 27
assign result_31 = ~w2998;// level 27
assign result_32 = w3005;// level 27
assign result_33 = ~w3012;// level 27
assign result_34 = w3019;// level 27
assign result_35 = ~w3026;// level 27
assign result_36 = ~w3033;// level 27
assign result_37 = ~w3040;// level 27
assign result_38 = w3047;// level 27
assign result_39 = ~w3054;// level 27
assign result_40 = ~w3061;// level 27
assign result_41 = ~w3068;// level 27
assign result_42 = ~w3075;// level 27
assign result_43 = ~w3082;// level 27
assign result_44 = ~w3089;// level 27
assign result_45 = ~w3096;// level 27
assign result_46 = w3103;// level 27
assign result_47 = ~w3110;// level 27
assign result_48 = w3117;// level 27
assign result_49 = ~w3124;// level 27
assign result_50 = w3131;// level 27
assign result_51 = ~w3138;// level 27
assign result_52 = ~w3145;// level 27
assign result_53 = ~w3152;// level 27
assign result_54 = w3159;// level 27
assign result_55 = ~w3166;// level 27
assign result_56 = ~w3173;// level 27
assign result_57 = ~w3180;// level 27
assign result_58 = ~w3187;// level 27
assign result_59 = ~w3194;// level 27
assign result_60 = ~w3201;// level 27
assign result_61 = ~w3208;// level 27
assign result_62 = w3215;// level 27
assign result_63 = ~w3222;// level 27
assign result_64 = w3229;// level 27
assign result_65 = ~w3236;// level 27
assign result_66 = w3243;// level 27
assign result_67 = ~w3250;// level 27
assign result_68 = ~w3257;// level 27
assign result_69 = ~w3264;// level 27
assign result_70 = w3271;// level 27
assign result_71 = ~w3278;// level 27
assign result_72 = w3285;// level 27
assign result_73 = ~w3292;// level 27
assign result_74 = w3299;// level 27
assign result_75 = ~w3306;// level 27
assign result_76 = ~w3313;// level 27
assign result_77 = ~w3320;// level 27
assign result_78 = w3327;// level 27
assign result_79 = ~w3334;// level 27
assign result_80 = w3341;// level 27
assign result_81 = ~w3348;// level 27
assign result_82 = w3355;// level 27
assign result_83 = ~w3362;// level 27
assign result_84 = ~w3369;// level 27
assign result_85 = ~w3376;// level 27
assign result_86 = w3383;// level 27
assign result_87 = ~w3390;// level 27
assign result_88 = w3397;// level 27
assign result_89 = ~w3404;// level 27
assign result_90 = w3411;// level 27
assign result_91 = ~w3418;// level 27
assign result_92 = ~w3425;// level 27
assign result_93 = ~w3432;// level 27
assign result_94 = w3439;// level 27
assign result_95 = ~w3446;// level 27
assign result_96 = w3453;// level 27
assign result_97 = ~w3460;// level 27
assign result_98 = w3467;// level 27
assign result_99 = ~w3474;// level 27
assign result_100 = ~w3481;// level 27
assign result_101 = ~w3488;// level 27
assign result_102 = w3495;// level 27
assign result_103 = ~w3502;// level 27
assign result_104 = w3509;// level 27
assign result_105 = ~w3516;// level 27
assign result_106 = w3523;// level 27
assign result_107 = ~w3530;// level 27
assign result_108 = ~w3537;// level 27
assign result_109 = ~w3544;// level 27
assign result_110 = w3551;// level 27
assign result_111 = ~w3558;// level 27
assign result_112 = w3565;// level 27
assign result_113 = ~w3572;// level 27
assign result_114 = w3579;// level 27
assign result_115 = ~w3586;// level 27
assign result_116 = ~w3593;// level 27
assign result_117 = ~w3600;// level 27
assign result_118 = w3607;// level 27
assign result_119 = ~w3614;// level 27
assign result_120 = w3621;// level 27
assign result_121 = ~w3628;// level 27
assign result_122 = w3635;// level 27
assign result_123 = ~w3642;// level 27
assign result_124 = ~w3649;// level 27
assign result_125 = ~w3656;// level 27
assign result_126 = ~w3662;// level 27
assign result_127 = w3663;// level 14
assign address_0 = w3670;// level 27
assign address_1 = ~w3671;// level 26
endmodule

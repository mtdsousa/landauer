// Benchmark "i2" written by ABC on Sun Apr 22 21:43:04 2018

module i2 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200,
    po0  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200;
  output po0;
  wire n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433;
  assign n203 = pi196 & pi200;
  assign n204 = pi198 & pi199;
  assign n205 = pi196 & n204;
  assign n206 = ~pi192 & ~pi193;
  assign n207 = ~pi190 & ~pi191;
  assign n208 = n206 & n207;
  assign n209 = pi194 & ~n208;
  assign n210 = ~pi188 & ~pi189;
  assign n211 = ~pi186 & ~pi187;
  assign n212 = n210 & n211;
  assign n213 = pi195 & ~n212;
  assign n214 = pi194 & n213;
  assign n215 = ~pi178 & ~pi179;
  assign n216 = ~pi176 & ~pi177;
  assign n217 = n215 & n216;
  assign n218 = ~pi174 & ~pi175;
  assign n219 = ~pi172 & ~pi173;
  assign n220 = n218 & n219;
  assign n221 = n217 & n220;
  assign n222 = ~pi170 & ~pi171;
  assign n223 = ~pi168 & ~pi169;
  assign n224 = n222 & n223;
  assign n225 = ~pi166 & ~pi167;
  assign n226 = ~pi164 & ~pi165;
  assign n227 = n225 & n226;
  assign n228 = n224 & n227;
  assign n229 = n221 & n228;
  assign n230 = pi180 & ~n229;
  assign n231 = ~pi162 & ~pi163;
  assign n232 = ~pi160 & ~pi161;
  assign n233 = n231 & n232;
  assign n234 = ~pi158 & ~pi159;
  assign n235 = ~pi156 & ~pi157;
  assign n236 = n234 & n235;
  assign n237 = n233 & n236;
  assign n238 = ~pi154 & ~pi155;
  assign n239 = ~pi152 & ~pi153;
  assign n240 = n238 & n239;
  assign n241 = ~pi150 & ~pi151;
  assign n242 = ~pi148 & ~pi149;
  assign n243 = n241 & n242;
  assign n244 = n240 & n243;
  assign n245 = n237 & n244;
  assign n246 = pi181 & ~n245;
  assign n247 = pi180 & n246;
  assign n248 = ~pi126 & ~pi127;
  assign n249 = ~pi124 & ~pi125;
  assign n250 = n248 & n249;
  assign n251 = ~pi122 & ~pi123;
  assign n252 = ~pi120 & ~pi121;
  assign n253 = n251 & n252;
  assign n254 = n250 & n253;
  assign n255 = ~pi118 & ~pi119;
  assign n256 = ~pi116 & ~pi117;
  assign n257 = n255 & n256;
  assign n258 = ~pi114 & ~pi115;
  assign n259 = ~pi112 & ~pi113;
  assign n260 = n258 & n259;
  assign n261 = n257 & n260;
  assign n262 = n254 & n261;
  assign n263 = ~pi110 & ~pi111;
  assign n264 = ~pi108 & ~pi109;
  assign n265 = n263 & n264;
  assign n266 = ~pi106 & ~pi107;
  assign n267 = ~pi104 & ~pi105;
  assign n268 = n266 & n267;
  assign n269 = n265 & n268;
  assign n270 = ~pi102 & ~pi103;
  assign n271 = ~pi100 & ~pi101;
  assign n272 = n270 & n271;
  assign n273 = ~pi098 & ~pi099;
  assign n274 = ~pi096 & ~pi097;
  assign n275 = n273 & n274;
  assign n276 = n272 & n275;
  assign n277 = n269 & n276;
  assign n278 = n262 & n277;
  assign n279 = pi130 & ~n278;
  assign n280 = pi128 & n279;
  assign n281 = pi128 & pi131;
  assign n282 = ~pi030 & ~pi031;
  assign n283 = ~pi028 & ~pi029;
  assign n284 = n282 & n283;
  assign n285 = ~pi026 & ~pi027;
  assign n286 = ~pi024 & ~pi025;
  assign n287 = n285 & n286;
  assign n288 = n284 & n287;
  assign n289 = ~pi022 & ~pi023;
  assign n290 = ~pi020 & ~pi021;
  assign n291 = n289 & n290;
  assign n292 = ~pi018 & ~pi019;
  assign n293 = ~pi016 & ~pi017;
  assign n294 = n292 & n293;
  assign n295 = n291 & n294;
  assign n296 = n288 & n295;
  assign n297 = ~pi014 & ~pi015;
  assign n298 = ~pi012 & ~pi013;
  assign n299 = n297 & n298;
  assign n300 = ~pi010 & ~pi011;
  assign n301 = ~pi008 & ~pi009;
  assign n302 = n300 & n301;
  assign n303 = n299 & n302;
  assign n304 = ~pi006 & ~pi007;
  assign n305 = ~pi004 & ~pi005;
  assign n306 = n304 & n305;
  assign n307 = ~pi002 & ~pi003;
  assign n308 = ~pi000 & ~pi001;
  assign n309 = n307 & n308;
  assign n310 = n306 & n309;
  assign n311 = n303 & n310;
  assign n312 = n296 & n311;
  assign n313 = pi130 & ~n312;
  assign n314 = ~pi128 & n313;
  assign n315 = ~pi128 & pi129;
  assign n316 = ~pi062 & ~pi063;
  assign n317 = ~pi060 & ~pi061;
  assign n318 = n316 & n317;
  assign n319 = ~pi058 & ~pi059;
  assign n320 = ~pi056 & ~pi057;
  assign n321 = n319 & n320;
  assign n322 = n318 & n321;
  assign n323 = ~pi054 & ~pi055;
  assign n324 = ~pi052 & ~pi053;
  assign n325 = n323 & n324;
  assign n326 = ~pi050 & ~pi051;
  assign n327 = ~pi048 & ~pi049;
  assign n328 = n326 & n327;
  assign n329 = n325 & n328;
  assign n330 = n322 & n329;
  assign n331 = ~pi046 & ~pi047;
  assign n332 = ~pi044 & ~pi045;
  assign n333 = n331 & n332;
  assign n334 = ~pi042 & ~pi043;
  assign n335 = ~pi040 & ~pi041;
  assign n336 = n334 & n335;
  assign n337 = n333 & n336;
  assign n338 = ~pi038 & ~pi039;
  assign n339 = ~pi036 & ~pi037;
  assign n340 = n338 & n339;
  assign n341 = ~pi034 & ~pi035;
  assign n342 = ~pi032 & ~pi033;
  assign n343 = n341 & n342;
  assign n344 = n340 & n343;
  assign n345 = n337 & n344;
  assign n346 = n330 & n345;
  assign n347 = pi130 & ~n346;
  assign n348 = ~pi128 & n347;
  assign n349 = ~pi094 & ~pi095;
  assign n350 = ~pi092 & ~pi093;
  assign n351 = n349 & n350;
  assign n352 = ~pi090 & ~pi091;
  assign n353 = ~pi088 & ~pi089;
  assign n354 = n352 & n353;
  assign n355 = n351 & n354;
  assign n356 = ~pi086 & ~pi087;
  assign n357 = ~pi084 & ~pi085;
  assign n358 = n356 & n357;
  assign n359 = ~pi082 & ~pi083;
  assign n360 = ~pi080 & ~pi081;
  assign n361 = n359 & n360;
  assign n362 = n358 & n361;
  assign n363 = n355 & n362;
  assign n364 = ~pi078 & ~pi079;
  assign n365 = ~pi076 & ~pi077;
  assign n366 = n364 & n365;
  assign n367 = ~pi074 & ~pi075;
  assign n368 = ~pi072 & ~pi073;
  assign n369 = n367 & n368;
  assign n370 = n366 & n369;
  assign n371 = ~pi070 & ~pi071;
  assign n372 = ~pi068 & ~pi069;
  assign n373 = n371 & n372;
  assign n374 = ~pi066 & ~pi067;
  assign n375 = ~pi064 & ~pi065;
  assign n376 = n374 & n375;
  assign n377 = n373 & n376;
  assign n378 = n370 & n377;
  assign n379 = n363 & n378;
  assign n380 = pi130 & ~n379;
  assign n381 = pi128 & n380;
  assign n382 = ~pi146 & ~pi147;
  assign n383 = ~pi144 & ~pi145;
  assign n384 = n382 & n383;
  assign n385 = ~pi142 & ~pi143;
  assign n386 = ~pi140 & ~pi141;
  assign n387 = n385 & n386;
  assign n388 = n384 & n387;
  assign n389 = ~pi138 & ~pi139;
  assign n390 = ~pi136 & ~pi137;
  assign n391 = n389 & n390;
  assign n392 = ~pi134 & ~pi135;
  assign n393 = ~pi132 & ~pi133;
  assign n394 = n392 & n393;
  assign n395 = n391 & n394;
  assign n396 = n388 & n395;
  assign n397 = pi180 & ~n396;
  assign n398 = pi181 & n397;
  assign n399 = pi181 & ~n229;
  assign n400 = pi180 & n399;
  assign n401 = ~pi184 & ~pi185;
  assign n402 = ~pi182 & ~pi183;
  assign n403 = n401 & n402;
  assign n404 = pi194 & ~n403;
  assign n405 = pi195 & n404;
  assign n406 = pi195 & ~n208;
  assign n407 = pi194 & n406;
  assign n408 = pi196 & pi197;
  assign n409 = pi198 & n408;
  assign n410 = pi198 & pi200;
  assign n411 = pi196 & n410;
  assign n412 = ~n409 & ~n411;
  assign n413 = ~n410 & n412;
  assign n414 = ~n405 & ~n407;
  assign n415 = ~n406 & n414;
  assign n416 = n413 & n415;
  assign n417 = ~n398 & ~n400;
  assign n418 = ~n399 & n417;
  assign n419 = ~n315 & ~n348;
  assign n420 = ~n381 & n419;
  assign n421 = n418 & n420;
  assign n422 = n416 & n421;
  assign n423 = ~n280 & ~n281;
  assign n424 = ~n314 & n423;
  assign n425 = ~n230 & ~n246;
  assign n426 = ~n247 & n425;
  assign n427 = n424 & n426;
  assign n428 = ~n209 & ~n213;
  assign n429 = ~n214 & n428;
  assign n430 = ~n203 & ~n204;
  assign n431 = ~n205 & n430;
  assign n432 = n429 & n431;
  assign n433 = n427 & n432;
  assign po0 = ~n422 | ~n433;
endmodule



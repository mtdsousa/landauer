// Benchmark "i8" written by ABC on Sun Apr 22 21:43:05 2018

module i8 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79, po80;
  wire n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n563, n564, n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
    n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3041,
    n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
    n3437, n3438, n3439, n3440, n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3516, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523;
  assign n215 = ~pi001 & ~pi005;
  assign n216 = ~pi095 & n215;
  assign n217 = pi007 & n216;
  assign n218 = pi088 & n217;
  assign n219 = ~pi005 & ~pi095;
  assign n220 = ~pi002 & n219;
  assign n221 = pi007 & n220;
  assign n222 = pi088 & n221;
  assign n223 = ~n217 & n222;
  assign n224 = ~pi007 & n219;
  assign n225 = pi089 & ~n221;
  assign n226 = ~n217 & n225;
  assign n227 = n224 & n226;
  assign n228 = ~pi005 & pi095;
  assign n229 = pi090 & ~n224;
  assign n230 = ~n217 & n229;
  assign n231 = ~n221 & n230;
  assign n232 = n228 & n231;
  assign n233 = pi087 & ~n228;
  assign n234 = ~n221 & n233;
  assign n235 = ~n217 & n234;
  assign n236 = ~n224 & n235;
  assign n237 = pi005 & n236;
  assign n238 = ~pi005 & ~n224;
  assign n239 = ~n217 & n238;
  assign n240 = ~n221 & n239;
  assign n241 = ~n228 & n240;
  assign n242 = ~n218 & ~n223;
  assign n243 = ~n227 & n242;
  assign n244 = ~n232 & ~n237;
  assign n245 = ~n241 & n244;
  assign po00 = ~n243 | ~n245;
  assign n247 = pi001 & ~pi095;
  assign n248 = pi002 & n247;
  assign n249 = ~pi008 & n248;
  assign n250 = ~pi130 & n249;
  assign n251 = pi000 & pi001;
  assign n252 = pi002 & n251;
  assign n253 = ~pi005 & ~n252;
  assign n254 = pi038 & ~n253;
  assign n255 = ~pi002 & ~pi005;
  assign n256 = ~pi001 & n255;
  assign n257 = pi007 & n256;
  assign n258 = ~pi004 & ~pi005;
  assign n259 = ~pi001 & n258;
  assign n260 = ~pi002 & n259;
  assign n261 = ~pi006 & n260;
  assign n262 = ~n257 & ~n261;
  assign n263 = pi001 & ~pi005;
  assign n264 = pi008 & n263;
  assign n265 = pi001 & n258;
  assign n266 = ~pi002 & n265;
  assign n267 = ~pi006 & n266;
  assign n268 = ~pi003 & ~pi005;
  assign n269 = ~pi004 & n268;
  assign n270 = pi007 & n268;
  assign n271 = ~n264 & ~n267;
  assign n272 = ~n269 & ~n270;
  assign n273 = n271 & n272;
  assign n274 = pi002 & ~pi005;
  assign n275 = ~pi001 & n274;
  assign n276 = pi008 & n275;
  assign n277 = pi001 & n274;
  assign n278 = ~pi000 & n277;
  assign n279 = pi003 & n259;
  assign n280 = pi002 & n279;
  assign n281 = ~pi006 & n280;
  assign n282 = ~n276 & ~n278;
  assign n283 = ~n281 & n282;
  assign n284 = n262 & n273;
  assign n285 = n253 & n284;
  assign n286 = n283 & n285;
  assign n287 = pi050 & n273;
  assign n288 = n253 & n287;
  assign n289 = ~n283 & n288;
  assign n290 = pi065 & n283;
  assign n291 = n253 & n290;
  assign n292 = n273 & n291;
  assign n293 = ~n262 & n292;
  assign n294 = ~n254 & ~n286;
  assign n295 = ~n289 & ~n293;
  assign n296 = n294 & n295;
  assign n297 = n250 & ~n296;
  assign n298 = ~pi008 & ~pi095;
  assign n299 = pi007 & n298;
  assign n300 = ~n296 & n299;
  assign n301 = ~n250 & n300;
  assign n302 = ~n296 & ~n299;
  assign n303 = ~n250 & n302;
  assign n304 = pi005 & n303;
  assign n305 = ~pi007 & n220;
  assign n306 = pi008 & n219;
  assign n307 = ~pi007 & n216;
  assign n308 = pi094 & ~n305;
  assign n309 = ~n306 & n308;
  assign n310 = ~n299 & n309;
  assign n311 = ~n250 & n310;
  assign n312 = ~pi005 & n311;
  assign n313 = ~n307 & n312;
  assign n314 = pi095 & n313;
  assign n315 = ~pi005 & n314;
  assign n316 = pi092 & ~n306;
  assign n317 = ~n299 & n316;
  assign n318 = ~n250 & n317;
  assign n319 = ~pi005 & n318;
  assign n320 = n307 & n319;
  assign n321 = pi092 & ~n307;
  assign n322 = ~pi005 & n321;
  assign n323 = ~n250 & n322;
  assign n324 = ~n299 & n323;
  assign n325 = ~n306 & n324;
  assign n326 = n305 & n325;
  assign n327 = ~n297 & ~n301;
  assign n328 = ~n304 & n327;
  assign n329 = ~n315 & ~n320;
  assign n330 = ~n326 & n329;
  assign po01 = ~n328 | ~n330;
  assign n332 = pi039 & ~n253;
  assign n333 = pi051 & n273;
  assign n334 = n253 & n333;
  assign n335 = ~n283 & n334;
  assign n336 = pi066 & n283;
  assign n337 = n253 & n336;
  assign n338 = n273 & n337;
  assign n339 = ~n262 & n338;
  assign n340 = ~n286 & ~n332;
  assign n341 = ~n335 & ~n339;
  assign n342 = n340 & n341;
  assign n343 = n250 & ~n342;
  assign n344 = n299 & ~n342;
  assign n345 = ~n250 & n344;
  assign n346 = ~n299 & ~n342;
  assign n347 = ~n250 & n346;
  assign n348 = pi005 & n347;
  assign n349 = ~pi005 & pi091;
  assign n350 = ~n250 & n349;
  assign n351 = ~n299 & n350;
  assign n352 = n306 & n351;
  assign n353 = pi093 & ~n306;
  assign n354 = ~n299 & n353;
  assign n355 = ~n250 & n354;
  assign n356 = ~pi005 & n355;
  assign n357 = n307 & n356;
  assign n358 = pi093 & ~n307;
  assign n359 = ~pi005 & n358;
  assign n360 = ~n250 & n359;
  assign n361 = ~n299 & n360;
  assign n362 = ~n306 & n361;
  assign n363 = n305 & n362;
  assign n364 = pi096 & ~n305;
  assign n365 = ~n306 & n364;
  assign n366 = ~n299 & n365;
  assign n367 = ~n250 & n366;
  assign n368 = ~pi005 & n367;
  assign n369 = ~n307 & n368;
  assign n370 = pi095 & n369;
  assign n371 = ~pi005 & n370;
  assign n372 = ~n343 & ~n345;
  assign n373 = ~n348 & ~n352;
  assign n374 = n372 & n373;
  assign n375 = ~n357 & ~n363;
  assign n376 = ~n371 & n375;
  assign po02 = ~n374 | ~n376;
  assign n378 = ~pi006 & ~pi095;
  assign n379 = ~pi130 & n378;
  assign n380 = pi032 & ~n253;
  assign n381 = pi040 & ~n273;
  assign n382 = n253 & n381;
  assign n383 = pi044 & n273;
  assign n384 = n253 & n383;
  assign n385 = ~n283 & n384;
  assign n386 = pi059 & n283;
  assign n387 = n253 & n386;
  assign n388 = n273 & n387;
  assign n389 = ~n262 & n388;
  assign n390 = ~n380 & ~n382;
  assign n391 = ~n385 & n390;
  assign n392 = ~n286 & ~n389;
  assign n393 = n391 & n392;
  assign n394 = n379 & ~n393;
  assign n395 = pi007 & ~pi095;
  assign n396 = ~n393 & n395;
  assign n397 = ~n379 & n396;
  assign n398 = ~n393 & ~n395;
  assign n399 = ~n379 & n398;
  assign n400 = pi005 & n399;
  assign n401 = ~pi005 & pi097;
  assign n402 = ~n379 & n401;
  assign n403 = ~n395 & n402;
  assign n404 = pi095 & n403;
  assign n405 = ~pi005 & n404;
  assign n406 = ~n394 & ~n397;
  assign n407 = ~n400 & ~n405;
  assign po03 = ~n406 | ~n407;
  assign n409 = pi033 & ~n253;
  assign n410 = pi045 & n273;
  assign n411 = n253 & n410;
  assign n412 = ~n283 & n411;
  assign n413 = pi060 & n283;
  assign n414 = n253 & n413;
  assign n415 = n273 & n414;
  assign n416 = ~n262 & n415;
  assign n417 = ~n286 & ~n409;
  assign n418 = ~n412 & ~n416;
  assign n419 = n417 & n418;
  assign n420 = n379 & ~n419;
  assign n421 = n395 & ~n419;
  assign n422 = ~n379 & n421;
  assign n423 = ~n395 & ~n419;
  assign n424 = ~n379 & n423;
  assign n425 = pi005 & n424;
  assign n426 = ~pi005 & pi098;
  assign n427 = ~n379 & n426;
  assign n428 = ~n395 & n427;
  assign n429 = pi095 & n428;
  assign n430 = ~pi005 & n429;
  assign n431 = ~n420 & ~n422;
  assign n432 = ~n425 & ~n430;
  assign po04 = ~n431 | ~n432;
  assign n434 = pi034 & ~n253;
  assign n435 = pi046 & n273;
  assign n436 = n253 & n435;
  assign n437 = ~n283 & n436;
  assign n438 = pi061 & n283;
  assign n439 = n253 & n438;
  assign n440 = n273 & n439;
  assign n441 = ~n262 & n440;
  assign n442 = ~n286 & ~n434;
  assign n443 = ~n437 & ~n441;
  assign n444 = n442 & n443;
  assign n445 = n379 & ~n444;
  assign n446 = n395 & ~n444;
  assign n447 = ~n379 & n446;
  assign n448 = ~n395 & ~n444;
  assign n449 = ~n379 & n448;
  assign n450 = pi005 & n449;
  assign n451 = ~pi005 & pi099;
  assign n452 = ~n379 & n451;
  assign n453 = ~n395 & n452;
  assign n454 = pi095 & n453;
  assign n455 = ~pi005 & n454;
  assign n456 = ~n445 & ~n447;
  assign n457 = ~n450 & ~n455;
  assign po05 = ~n456 | ~n457;
  assign n459 = pi035 & ~n253;
  assign n460 = pi047 & n273;
  assign n461 = n253 & n460;
  assign n462 = ~n283 & n461;
  assign n463 = pi062 & n283;
  assign n464 = n253 & n463;
  assign n465 = n273 & n464;
  assign n466 = ~n262 & n465;
  assign n467 = ~n286 & ~n459;
  assign n468 = ~n462 & ~n466;
  assign n469 = n467 & n468;
  assign n470 = n379 & ~n469;
  assign n471 = n395 & ~n469;
  assign n472 = ~n379 & n471;
  assign n473 = ~n395 & ~n469;
  assign n474 = ~n379 & n473;
  assign n475 = pi005 & n474;
  assign n476 = ~pi005 & pi100;
  assign n477 = ~n379 & n476;
  assign n478 = ~n395 & n477;
  assign n479 = pi095 & n478;
  assign n480 = ~pi005 & n479;
  assign n481 = ~n470 & ~n472;
  assign n482 = ~n475 & ~n480;
  assign po06 = ~n481 | ~n482;
  assign n484 = pi036 & ~n253;
  assign n485 = pi048 & n273;
  assign n486 = n253 & n485;
  assign n487 = ~n283 & n486;
  assign n488 = pi063 & n283;
  assign n489 = n253 & n488;
  assign n490 = n273 & n489;
  assign n491 = ~n262 & n490;
  assign n492 = ~n286 & ~n484;
  assign n493 = ~n487 & ~n491;
  assign n494 = n492 & n493;
  assign n495 = n379 & ~n494;
  assign n496 = n395 & ~n494;
  assign n497 = ~n379 & n496;
  assign n498 = ~n395 & ~n494;
  assign n499 = ~n379 & n498;
  assign n500 = pi005 & n499;
  assign n501 = ~pi005 & pi101;
  assign n502 = ~n379 & n501;
  assign n503 = ~n395 & n502;
  assign n504 = pi095 & n503;
  assign n505 = ~pi005 & n504;
  assign n506 = ~n495 & ~n497;
  assign n507 = ~n500 & ~n505;
  assign po07 = ~n506 | ~n507;
  assign n509 = pi037 & ~n253;
  assign n510 = pi049 & n273;
  assign n511 = n253 & n510;
  assign n512 = ~n283 & n511;
  assign n513 = pi064 & n283;
  assign n514 = n253 & n513;
  assign n515 = n273 & n514;
  assign n516 = ~n262 & n515;
  assign n517 = ~n286 & ~n509;
  assign n518 = ~n512 & ~n516;
  assign n519 = n517 & n518;
  assign n520 = n379 & ~n519;
  assign n521 = n395 & ~n519;
  assign n522 = ~n379 & n521;
  assign n523 = ~n395 & ~n519;
  assign n524 = ~n379 & n523;
  assign n525 = pi005 & n524;
  assign n526 = ~pi005 & pi102;
  assign n527 = ~n379 & n526;
  assign n528 = ~n395 & n527;
  assign n529 = pi095 & n528;
  assign n530 = ~pi005 & n529;
  assign n531 = ~n520 & ~n522;
  assign n532 = ~n525 & ~n530;
  assign po08 = ~n531 | ~n532;
  assign n534 = ~pi095 & ~pi130;
  assign n535 = pi031 & ~n253;
  assign n536 = pi039 & ~n273;
  assign n537 = n253 & n536;
  assign n538 = pi043 & n273;
  assign n539 = n253 & n538;
  assign n540 = ~n283 & n539;
  assign n541 = pi058 & n283;
  assign n542 = n253 & n541;
  assign n543 = n273 & n542;
  assign n544 = ~n262 & n543;
  assign n545 = ~n535 & ~n537;
  assign n546 = ~n540 & n545;
  assign n547 = ~n286 & ~n544;
  assign n548 = n546 & n547;
  assign n549 = n534 & ~n548;
  assign n550 = n395 & ~n548;
  assign n551 = ~n534 & n550;
  assign n552 = ~n395 & ~n548;
  assign n553 = ~n534 & n552;
  assign n554 = pi005 & n553;
  assign n555 = ~pi005 & pi103;
  assign n556 = ~n534 & n555;
  assign n557 = ~n395 & n556;
  assign n558 = pi095 & n557;
  assign n559 = ~pi005 & n558;
  assign n560 = ~n549 & ~n551;
  assign n561 = ~n554 & ~n559;
  assign po09 = ~n560 | ~n561;
  assign n563 = pi029 & ~n253;
  assign n564 = pi037 & ~n273;
  assign n565 = n253 & n564;
  assign n566 = pi041 & n273;
  assign n567 = n253 & n566;
  assign n568 = ~n283 & n567;
  assign n569 = pi056 & n283;
  assign n570 = n253 & n569;
  assign n571 = n273 & n570;
  assign n572 = ~n262 & n571;
  assign n573 = ~n563 & ~n565;
  assign n574 = ~n568 & n573;
  assign n575 = ~n286 & ~n572;
  assign n576 = n574 & n575;
  assign n577 = n379 & ~n576;
  assign n578 = n395 & ~n576;
  assign n579 = ~n379 & n578;
  assign n580 = ~n395 & ~n576;
  assign n581 = ~n379 & n580;
  assign n582 = pi005 & n581;
  assign n583 = ~pi005 & pi104;
  assign n584 = ~n379 & n583;
  assign n585 = ~n395 & n584;
  assign n586 = pi095 & n585;
  assign n587 = ~pi005 & n586;
  assign n588 = ~n577 & ~n579;
  assign n589 = ~n582 & ~n587;
  assign po10 = ~n588 | ~n589;
  assign n591 = pi030 & ~n253;
  assign n592 = pi038 & ~n273;
  assign n593 = n253 & n592;
  assign n594 = pi042 & n273;
  assign n595 = n253 & n594;
  assign n596 = ~n283 & n595;
  assign n597 = pi057 & n283;
  assign n598 = n253 & n597;
  assign n599 = n273 & n598;
  assign n600 = ~n262 & n599;
  assign n601 = ~n591 & ~n593;
  assign n602 = ~n596 & n601;
  assign n603 = ~n286 & ~n600;
  assign n604 = n602 & n603;
  assign n605 = n379 & ~n604;
  assign n606 = n395 & ~n604;
  assign n607 = ~n379 & n606;
  assign n608 = ~n395 & ~n604;
  assign n609 = ~n379 & n608;
  assign n610 = pi005 & n609;
  assign n611 = ~pi005 & pi105;
  assign n612 = ~n379 & n611;
  assign n613 = ~n395 & n612;
  assign n614 = pi095 & n613;
  assign n615 = ~pi005 & n614;
  assign n616 = ~n605 & ~n607;
  assign n617 = ~n610 & ~n615;
  assign po11 = ~n616 | ~n617;
  assign n619 = ~pi001 & ~pi095;
  assign n620 = ~pi130 & n619;
  assign n621 = pi028 & ~n253;
  assign n622 = pi036 & ~n273;
  assign n623 = n253 & n622;
  assign n624 = pi039 & n273;
  assign n625 = n253 & n624;
  assign n626 = ~n283 & n625;
  assign n627 = pi055 & n283;
  assign n628 = n253 & n627;
  assign n629 = n273 & n628;
  assign n630 = ~n262 & n629;
  assign n631 = ~n621 & ~n623;
  assign n632 = ~n626 & n631;
  assign n633 = ~n286 & ~n630;
  assign n634 = n632 & n633;
  assign n635 = n620 & ~n634;
  assign n636 = ~pi002 & n378;
  assign n637 = ~pi130 & n636;
  assign n638 = ~n634 & n637;
  assign n639 = ~n620 & n638;
  assign n640 = pi000 & n534;
  assign n641 = ~n634 & ~n637;
  assign n642 = ~n620 & n641;
  assign n643 = n640 & n642;
  assign n644 = ~n634 & ~n640;
  assign n645 = ~n620 & n644;
  assign n646 = ~n637 & n645;
  assign n647 = n395 & n646;
  assign n648 = ~n395 & ~n634;
  assign n649 = ~n637 & n648;
  assign n650 = ~n620 & n649;
  assign n651 = ~n640 & n650;
  assign n652 = pi005 & n651;
  assign n653 = ~pi005 & pi106;
  assign n654 = ~n640 & n653;
  assign n655 = ~n620 & n654;
  assign n656 = ~n637 & n655;
  assign n657 = ~n395 & n656;
  assign n658 = n228 & n657;
  assign n659 = pi086 & ~n228;
  assign n660 = ~n395 & n659;
  assign n661 = ~n637 & n660;
  assign n662 = ~n620 & n661;
  assign n663 = ~n640 & n662;
  assign n664 = ~pi005 & n663;
  assign n665 = ~pi007 & n664;
  assign n666 = ~pi095 & n665;
  assign n667 = ~pi130 & n666;
  assign n668 = ~pi000 & n667;
  assign n669 = pi002 & n668;
  assign n670 = pi001 & n669;
  assign n671 = ~pi005 & n670;
  assign n672 = ~n635 & ~n639;
  assign n673 = ~n643 & ~n647;
  assign n674 = n672 & n673;
  assign n675 = ~n652 & ~n658;
  assign n676 = ~n671 & n675;
  assign po12 = ~n674 | ~n676;
  assign n678 = ~pi006 & n619;
  assign n679 = ~pi130 & n678;
  assign n680 = pi025 & ~n253;
  assign n681 = pi033 & ~n273;
  assign n682 = n253 & n681;
  assign n683 = pi036 & n273;
  assign n684 = n253 & n683;
  assign n685 = ~n283 & n684;
  assign n686 = pi052 & n283;
  assign n687 = n253 & n686;
  assign n688 = n273 & n687;
  assign n689 = ~n262 & n688;
  assign n690 = ~n680 & ~n682;
  assign n691 = ~n685 & n690;
  assign n692 = ~n286 & ~n689;
  assign n693 = n691 & n692;
  assign n694 = n679 & ~n693;
  assign n695 = n637 & ~n693;
  assign n696 = ~n679 & n695;
  assign n697 = ~n637 & ~n693;
  assign n698 = ~n679 & n697;
  assign n699 = n640 & n698;
  assign n700 = ~n640 & ~n693;
  assign n701 = ~n679 & n700;
  assign n702 = ~n637 & n701;
  assign n703 = n395 & n702;
  assign n704 = ~n395 & ~n693;
  assign n705 = ~n637 & n704;
  assign n706 = ~n679 & n705;
  assign n707 = ~n640 & n706;
  assign n708 = pi005 & n707;
  assign n709 = ~pi005 & pi107;
  assign n710 = ~n640 & n709;
  assign n711 = ~n679 & n710;
  assign n712 = ~n637 & n711;
  assign n713 = ~n395 & n712;
  assign n714 = n228 & n713;
  assign n715 = pi083 & ~n228;
  assign n716 = ~n395 & n715;
  assign n717 = ~n637 & n716;
  assign n718 = ~n679 & n717;
  assign n719 = ~n640 & n718;
  assign n720 = ~pi005 & n719;
  assign n721 = ~pi007 & n720;
  assign n722 = ~pi095 & n721;
  assign n723 = ~pi130 & n722;
  assign n724 = ~pi000 & n723;
  assign n725 = pi002 & n724;
  assign n726 = pi001 & n725;
  assign n727 = ~pi005 & n726;
  assign n728 = ~n694 & ~n696;
  assign n729 = ~n699 & ~n703;
  assign n730 = n728 & n729;
  assign n731 = ~n708 & ~n714;
  assign n732 = ~n727 & n731;
  assign po13 = ~n730 | ~n732;
  assign n734 = pi026 & ~n253;
  assign n735 = pi034 & ~n273;
  assign n736 = n253 & n735;
  assign n737 = pi037 & n273;
  assign n738 = n253 & n737;
  assign n739 = ~n283 & n738;
  assign n740 = pi053 & n283;
  assign n741 = n253 & n740;
  assign n742 = n273 & n741;
  assign n743 = ~n262 & n742;
  assign n744 = ~n734 & ~n736;
  assign n745 = ~n739 & n744;
  assign n746 = ~n286 & ~n743;
  assign n747 = n745 & n746;
  assign n748 = n679 & ~n747;
  assign n749 = n637 & ~n747;
  assign n750 = ~n679 & n749;
  assign n751 = ~n637 & ~n747;
  assign n752 = ~n679 & n751;
  assign n753 = n640 & n752;
  assign n754 = ~n640 & ~n747;
  assign n755 = ~n679 & n754;
  assign n756 = ~n637 & n755;
  assign n757 = n395 & n756;
  assign n758 = ~n395 & ~n747;
  assign n759 = ~n637 & n758;
  assign n760 = ~n679 & n759;
  assign n761 = ~n640 & n760;
  assign n762 = pi005 & n761;
  assign n763 = ~pi005 & pi108;
  assign n764 = ~n640 & n763;
  assign n765 = ~n679 & n764;
  assign n766 = ~n637 & n765;
  assign n767 = ~n395 & n766;
  assign n768 = n228 & n767;
  assign n769 = pi084 & ~n228;
  assign n770 = ~n395 & n769;
  assign n771 = ~n637 & n770;
  assign n772 = ~n679 & n771;
  assign n773 = ~n640 & n772;
  assign n774 = ~pi005 & n773;
  assign n775 = ~pi007 & n774;
  assign n776 = ~pi095 & n775;
  assign n777 = ~pi130 & n776;
  assign n778 = ~pi000 & n777;
  assign n779 = pi002 & n778;
  assign n780 = pi001 & n779;
  assign n781 = ~pi005 & n780;
  assign n782 = ~n748 & ~n750;
  assign n783 = ~n753 & ~n757;
  assign n784 = n782 & n783;
  assign n785 = ~n762 & ~n768;
  assign n786 = ~n781 & n785;
  assign po14 = ~n784 | ~n786;
  assign n788 = pi027 & ~n253;
  assign n789 = pi035 & ~n273;
  assign n790 = n253 & n789;
  assign n791 = pi038 & n273;
  assign n792 = n253 & n791;
  assign n793 = ~n283 & n792;
  assign n794 = pi054 & n283;
  assign n795 = n253 & n794;
  assign n796 = n273 & n795;
  assign n797 = ~n262 & n796;
  assign n798 = ~n788 & ~n790;
  assign n799 = ~n793 & n798;
  assign n800 = ~n286 & ~n797;
  assign n801 = n799 & n800;
  assign n802 = n679 & ~n801;
  assign n803 = n637 & ~n801;
  assign n804 = ~n679 & n803;
  assign n805 = ~n637 & ~n801;
  assign n806 = ~n679 & n805;
  assign n807 = n640 & n806;
  assign n808 = ~n640 & ~n801;
  assign n809 = ~n679 & n808;
  assign n810 = ~n637 & n809;
  assign n811 = n395 & n810;
  assign n812 = ~n395 & ~n801;
  assign n813 = ~n637 & n812;
  assign n814 = ~n679 & n813;
  assign n815 = ~n640 & n814;
  assign n816 = pi005 & n815;
  assign n817 = ~pi005 & pi109;
  assign n818 = ~n640 & n817;
  assign n819 = ~n679 & n818;
  assign n820 = ~n637 & n819;
  assign n821 = ~n395 & n820;
  assign n822 = n228 & n821;
  assign n823 = pi085 & ~n228;
  assign n824 = ~n395 & n823;
  assign n825 = ~n637 & n824;
  assign n826 = ~n679 & n825;
  assign n827 = ~n640 & n826;
  assign n828 = ~pi005 & n827;
  assign n829 = ~pi007 & n828;
  assign n830 = ~pi095 & n829;
  assign n831 = ~pi130 & n830;
  assign n832 = ~pi000 & n831;
  assign n833 = pi002 & n832;
  assign n834 = pi001 & n833;
  assign n835 = ~pi005 & n834;
  assign n836 = ~n802 & ~n804;
  assign n837 = ~n807 & ~n811;
  assign n838 = n836 & n837;
  assign n839 = ~n816 & ~n822;
  assign n840 = ~n835 & n839;
  assign po15 = ~n838 | ~n840;
  assign n842 = ~pi002 & n619;
  assign n843 = ~pi130 & n842;
  assign n844 = pi024 & ~n253;
  assign n845 = pi032 & ~n273;
  assign n846 = n253 & n845;
  assign n847 = pi035 & n273;
  assign n848 = n253 & n847;
  assign n849 = ~n283 & n848;
  assign n850 = pi039 & n283;
  assign n851 = n253 & n850;
  assign n852 = n273 & n851;
  assign n853 = ~n262 & n852;
  assign n854 = ~n844 & ~n846;
  assign n855 = ~n849 & n854;
  assign n856 = ~n286 & ~n853;
  assign n857 = n855 & n856;
  assign n858 = n843 & ~n857;
  assign n859 = n679 & ~n857;
  assign n860 = ~n843 & n859;
  assign n861 = ~n679 & ~n857;
  assign n862 = ~n843 & n861;
  assign n863 = n637 & n862;
  assign n864 = ~n637 & ~n857;
  assign n865 = ~n843 & n864;
  assign n866 = ~n679 & n865;
  assign n867 = n640 & n866;
  assign n868 = ~n640 & ~n857;
  assign n869 = ~n679 & n868;
  assign n870 = ~n843 & n869;
  assign n871 = ~n637 & n870;
  assign n872 = n395 & n871;
  assign n873 = ~n395 & ~n857;
  assign n874 = ~n637 & n873;
  assign n875 = ~n843 & n874;
  assign n876 = ~n679 & n875;
  assign n877 = ~n640 & n876;
  assign n878 = pi005 & n877;
  assign n879 = ~pi005 & pi110;
  assign n880 = ~n640 & n879;
  assign n881 = ~n679 & n880;
  assign n882 = ~n843 & n881;
  assign n883 = ~n637 & n882;
  assign n884 = ~n395 & n883;
  assign n885 = n228 & n884;
  assign n886 = pi082 & ~n228;
  assign n887 = ~n395 & n886;
  assign n888 = ~n637 & n887;
  assign n889 = ~n843 & n888;
  assign n890 = ~n679 & n889;
  assign n891 = ~n640 & n890;
  assign n892 = ~pi005 & n891;
  assign n893 = ~pi007 & n892;
  assign n894 = ~pi095 & n893;
  assign n895 = ~pi130 & n894;
  assign n896 = ~pi000 & n895;
  assign n897 = pi002 & n896;
  assign n898 = pi001 & n897;
  assign n899 = ~pi005 & n898;
  assign n900 = ~n858 & ~n860;
  assign n901 = ~n863 & ~n867;
  assign n902 = n900 & n901;
  assign n903 = ~n872 & ~n878;
  assign n904 = ~n885 & ~n899;
  assign n905 = n903 & n904;
  assign po16 = ~n902 | ~n905;
  assign n907 = pi009 & ~n253;
  assign n908 = pi017 & ~n273;
  assign n909 = n253 & n908;
  assign n910 = pi020 & n273;
  assign n911 = n253 & n910;
  assign n912 = ~n283 & n911;
  assign n913 = pi024 & n283;
  assign n914 = n253 & n913;
  assign n915 = n273 & n914;
  assign n916 = ~n262 & n915;
  assign n917 = ~n907 & ~n909;
  assign n918 = ~n912 & n917;
  assign n919 = ~n286 & ~n916;
  assign n920 = n918 & n919;
  assign n921 = n679 & ~n920;
  assign n922 = n637 & ~n920;
  assign n923 = ~n679 & n922;
  assign n924 = ~n637 & ~n920;
  assign n925 = ~n679 & n924;
  assign n926 = n640 & n925;
  assign n927 = ~n640 & ~n920;
  assign n928 = ~n679 & n927;
  assign n929 = ~n637 & n928;
  assign n930 = n395 & n929;
  assign n931 = ~n395 & ~n920;
  assign n932 = ~n637 & n931;
  assign n933 = ~n679 & n932;
  assign n934 = ~n640 & n933;
  assign n935 = pi005 & n934;
  assign n936 = ~pi005 & pi111;
  assign n937 = ~n640 & n936;
  assign n938 = ~n679 & n937;
  assign n939 = ~n637 & n938;
  assign n940 = ~n395 & n939;
  assign n941 = n228 & n940;
  assign n942 = pi067 & ~n228;
  assign n943 = ~n395 & n942;
  assign n944 = ~n637 & n943;
  assign n945 = ~n679 & n944;
  assign n946 = ~n640 & n945;
  assign n947 = ~pi005 & n946;
  assign n948 = ~pi007 & n947;
  assign n949 = ~pi095 & n948;
  assign n950 = ~pi130 & n949;
  assign n951 = ~pi000 & n950;
  assign n952 = pi002 & n951;
  assign n953 = pi001 & n952;
  assign n954 = ~pi005 & n953;
  assign n955 = ~n921 & ~n923;
  assign n956 = ~n926 & ~n930;
  assign n957 = n955 & n956;
  assign n958 = ~n935 & ~n941;
  assign n959 = ~n954 & n958;
  assign po17 = ~n957 | ~n959;
  assign n961 = pi010 & ~n253;
  assign n962 = pi018 & ~n273;
  assign n963 = n253 & n962;
  assign n964 = pi021 & n273;
  assign n965 = n253 & n964;
  assign n966 = ~n283 & n965;
  assign n967 = pi025 & n283;
  assign n968 = n253 & n967;
  assign n969 = n273 & n968;
  assign n970 = ~n262 & n969;
  assign n971 = ~n961 & ~n963;
  assign n972 = ~n966 & n971;
  assign n973 = ~n286 & ~n970;
  assign n974 = n972 & n973;
  assign n975 = n679 & ~n974;
  assign n976 = n637 & ~n974;
  assign n977 = ~n679 & n976;
  assign n978 = ~n637 & ~n974;
  assign n979 = ~n679 & n978;
  assign n980 = n640 & n979;
  assign n981 = ~n640 & ~n974;
  assign n982 = ~n679 & n981;
  assign n983 = ~n637 & n982;
  assign n984 = n395 & n983;
  assign n985 = ~n395 & ~n974;
  assign n986 = ~n637 & n985;
  assign n987 = ~n679 & n986;
  assign n988 = ~n640 & n987;
  assign n989 = pi005 & n988;
  assign n990 = ~pi005 & pi112;
  assign n991 = ~n640 & n990;
  assign n992 = ~n679 & n991;
  assign n993 = ~n637 & n992;
  assign n994 = ~n395 & n993;
  assign n995 = n228 & n994;
  assign n996 = pi068 & ~n228;
  assign n997 = ~n395 & n996;
  assign n998 = ~n637 & n997;
  assign n999 = ~n679 & n998;
  assign n1000 = ~n640 & n999;
  assign n1001 = ~pi005 & n1000;
  assign n1002 = ~pi007 & n1001;
  assign n1003 = ~pi095 & n1002;
  assign n1004 = ~pi130 & n1003;
  assign n1005 = ~pi000 & n1004;
  assign n1006 = pi002 & n1005;
  assign n1007 = pi001 & n1006;
  assign n1008 = ~pi005 & n1007;
  assign n1009 = ~n975 & ~n977;
  assign n1010 = ~n980 & ~n984;
  assign n1011 = n1009 & n1010;
  assign n1012 = ~n989 & ~n995;
  assign n1013 = ~n1008 & n1012;
  assign po18 = ~n1011 | ~n1013;
  assign n1015 = pi011 & ~n253;
  assign n1016 = pi019 & ~n273;
  assign n1017 = n253 & n1016;
  assign n1018 = pi022 & n273;
  assign n1019 = n253 & n1018;
  assign n1020 = ~n283 & n1019;
  assign n1021 = pi026 & n283;
  assign n1022 = n253 & n1021;
  assign n1023 = n273 & n1022;
  assign n1024 = ~n262 & n1023;
  assign n1025 = ~n1015 & ~n1017;
  assign n1026 = ~n1020 & n1025;
  assign n1027 = ~n286 & ~n1024;
  assign n1028 = n1026 & n1027;
  assign n1029 = n679 & ~n1028;
  assign n1030 = n637 & ~n1028;
  assign n1031 = ~n679 & n1030;
  assign n1032 = ~n637 & ~n1028;
  assign n1033 = ~n679 & n1032;
  assign n1034 = n640 & n1033;
  assign n1035 = ~n640 & ~n1028;
  assign n1036 = ~n679 & n1035;
  assign n1037 = ~n637 & n1036;
  assign n1038 = n395 & n1037;
  assign n1039 = ~n395 & ~n1028;
  assign n1040 = ~n637 & n1039;
  assign n1041 = ~n679 & n1040;
  assign n1042 = ~n640 & n1041;
  assign n1043 = pi005 & n1042;
  assign n1044 = ~pi005 & pi113;
  assign n1045 = ~n640 & n1044;
  assign n1046 = ~n679 & n1045;
  assign n1047 = ~n637 & n1046;
  assign n1048 = ~n395 & n1047;
  assign n1049 = n228 & n1048;
  assign n1050 = pi069 & ~n228;
  assign n1051 = ~n395 & n1050;
  assign n1052 = ~n637 & n1051;
  assign n1053 = ~n679 & n1052;
  assign n1054 = ~n640 & n1053;
  assign n1055 = ~pi005 & n1054;
  assign n1056 = ~pi007 & n1055;
  assign n1057 = ~pi095 & n1056;
  assign n1058 = ~pi130 & n1057;
  assign n1059 = ~pi000 & n1058;
  assign n1060 = pi002 & n1059;
  assign n1061 = pi001 & n1060;
  assign n1062 = ~pi005 & n1061;
  assign n1063 = ~n1029 & ~n1031;
  assign n1064 = ~n1034 & ~n1038;
  assign n1065 = n1063 & n1064;
  assign n1066 = ~n1043 & ~n1049;
  assign n1067 = ~n1062 & n1066;
  assign po19 = ~n1065 | ~n1067;
  assign n1069 = pi012 & ~n253;
  assign n1070 = pi020 & ~n273;
  assign n1071 = n253 & n1070;
  assign n1072 = pi023 & n273;
  assign n1073 = n253 & n1072;
  assign n1074 = ~n283 & n1073;
  assign n1075 = pi027 & n283;
  assign n1076 = n253 & n1075;
  assign n1077 = n273 & n1076;
  assign n1078 = ~n262 & n1077;
  assign n1079 = ~n1069 & ~n1071;
  assign n1080 = ~n1074 & n1079;
  assign n1081 = ~n286 & ~n1078;
  assign n1082 = n1080 & n1081;
  assign n1083 = n679 & ~n1082;
  assign n1084 = n637 & ~n1082;
  assign n1085 = ~n679 & n1084;
  assign n1086 = ~n637 & ~n1082;
  assign n1087 = ~n679 & n1086;
  assign n1088 = n640 & n1087;
  assign n1089 = ~n640 & ~n1082;
  assign n1090 = ~n679 & n1089;
  assign n1091 = ~n637 & n1090;
  assign n1092 = n395 & n1091;
  assign n1093 = ~n395 & ~n1082;
  assign n1094 = ~n637 & n1093;
  assign n1095 = ~n679 & n1094;
  assign n1096 = ~n640 & n1095;
  assign n1097 = pi005 & n1096;
  assign n1098 = ~pi005 & pi114;
  assign n1099 = ~n640 & n1098;
  assign n1100 = ~n679 & n1099;
  assign n1101 = ~n637 & n1100;
  assign n1102 = ~n395 & n1101;
  assign n1103 = n228 & n1102;
  assign n1104 = pi070 & ~n228;
  assign n1105 = ~n395 & n1104;
  assign n1106 = ~n637 & n1105;
  assign n1107 = ~n679 & n1106;
  assign n1108 = ~n640 & n1107;
  assign n1109 = ~pi005 & n1108;
  assign n1110 = ~pi007 & n1109;
  assign n1111 = ~pi095 & n1110;
  assign n1112 = ~pi130 & n1111;
  assign n1113 = ~pi000 & n1112;
  assign n1114 = pi002 & n1113;
  assign n1115 = pi001 & n1114;
  assign n1116 = ~pi005 & n1115;
  assign n1117 = ~n1083 & ~n1085;
  assign n1118 = ~n1088 & ~n1092;
  assign n1119 = n1117 & n1118;
  assign n1120 = ~n1097 & ~n1103;
  assign n1121 = ~n1116 & n1120;
  assign po20 = ~n1119 | ~n1121;
  assign n1123 = pi013 & ~n253;
  assign n1124 = pi021 & ~n273;
  assign n1125 = n253 & n1124;
  assign n1126 = pi024 & n273;
  assign n1127 = n253 & n1126;
  assign n1128 = ~n283 & n1127;
  assign n1129 = pi028 & n283;
  assign n1130 = n253 & n1129;
  assign n1131 = n273 & n1130;
  assign n1132 = ~n262 & n1131;
  assign n1133 = ~n1123 & ~n1125;
  assign n1134 = ~n1128 & n1133;
  assign n1135 = ~n286 & ~n1132;
  assign n1136 = n1134 & n1135;
  assign n1137 = n679 & ~n1136;
  assign n1138 = n637 & ~n1136;
  assign n1139 = ~n679 & n1138;
  assign n1140 = ~n637 & ~n1136;
  assign n1141 = ~n679 & n1140;
  assign n1142 = n640 & n1141;
  assign n1143 = ~n640 & ~n1136;
  assign n1144 = ~n679 & n1143;
  assign n1145 = ~n637 & n1144;
  assign n1146 = n395 & n1145;
  assign n1147 = ~n395 & ~n1136;
  assign n1148 = ~n637 & n1147;
  assign n1149 = ~n679 & n1148;
  assign n1150 = ~n640 & n1149;
  assign n1151 = pi005 & n1150;
  assign n1152 = ~pi005 & pi115;
  assign n1153 = ~n640 & n1152;
  assign n1154 = ~n679 & n1153;
  assign n1155 = ~n637 & n1154;
  assign n1156 = ~n395 & n1155;
  assign n1157 = n228 & n1156;
  assign n1158 = pi071 & ~n228;
  assign n1159 = ~n395 & n1158;
  assign n1160 = ~n637 & n1159;
  assign n1161 = ~n679 & n1160;
  assign n1162 = ~n640 & n1161;
  assign n1163 = ~pi005 & n1162;
  assign n1164 = ~pi007 & n1163;
  assign n1165 = ~pi095 & n1164;
  assign n1166 = ~pi130 & n1165;
  assign n1167 = ~pi000 & n1166;
  assign n1168 = pi002 & n1167;
  assign n1169 = pi001 & n1168;
  assign n1170 = ~pi005 & n1169;
  assign n1171 = ~n1137 & ~n1139;
  assign n1172 = ~n1142 & ~n1146;
  assign n1173 = n1171 & n1172;
  assign n1174 = ~n1151 & ~n1157;
  assign n1175 = ~n1170 & n1174;
  assign po21 = ~n1173 | ~n1175;
  assign n1177 = pi014 & ~n253;
  assign n1178 = pi022 & ~n273;
  assign n1179 = n253 & n1178;
  assign n1180 = pi025 & n273;
  assign n1181 = n253 & n1180;
  assign n1182 = ~n283 & n1181;
  assign n1183 = pi029 & n283;
  assign n1184 = n253 & n1183;
  assign n1185 = n273 & n1184;
  assign n1186 = ~n262 & n1185;
  assign n1187 = ~n1177 & ~n1179;
  assign n1188 = ~n1182 & n1187;
  assign n1189 = ~n286 & ~n1186;
  assign n1190 = n1188 & n1189;
  assign n1191 = n679 & ~n1190;
  assign n1192 = n637 & ~n1190;
  assign n1193 = ~n679 & n1192;
  assign n1194 = ~n637 & ~n1190;
  assign n1195 = ~n679 & n1194;
  assign n1196 = n640 & n1195;
  assign n1197 = ~n640 & ~n1190;
  assign n1198 = ~n679 & n1197;
  assign n1199 = ~n637 & n1198;
  assign n1200 = n395 & n1199;
  assign n1201 = ~n395 & ~n1190;
  assign n1202 = ~n637 & n1201;
  assign n1203 = ~n679 & n1202;
  assign n1204 = ~n640 & n1203;
  assign n1205 = pi005 & n1204;
  assign n1206 = ~pi005 & pi116;
  assign n1207 = ~n640 & n1206;
  assign n1208 = ~n679 & n1207;
  assign n1209 = ~n637 & n1208;
  assign n1210 = ~n395 & n1209;
  assign n1211 = n228 & n1210;
  assign n1212 = pi072 & ~n228;
  assign n1213 = ~n395 & n1212;
  assign n1214 = ~n637 & n1213;
  assign n1215 = ~n679 & n1214;
  assign n1216 = ~n640 & n1215;
  assign n1217 = ~pi005 & n1216;
  assign n1218 = ~pi007 & n1217;
  assign n1219 = ~pi095 & n1218;
  assign n1220 = ~pi130 & n1219;
  assign n1221 = ~pi000 & n1220;
  assign n1222 = pi002 & n1221;
  assign n1223 = pi001 & n1222;
  assign n1224 = ~pi005 & n1223;
  assign n1225 = ~n1191 & ~n1193;
  assign n1226 = ~n1196 & ~n1200;
  assign n1227 = n1225 & n1226;
  assign n1228 = ~n1205 & ~n1211;
  assign n1229 = ~n1224 & n1228;
  assign po22 = ~n1227 | ~n1229;
  assign n1231 = pi015 & ~n253;
  assign n1232 = pi023 & ~n273;
  assign n1233 = n253 & n1232;
  assign n1234 = pi026 & n273;
  assign n1235 = n253 & n1234;
  assign n1236 = ~n283 & n1235;
  assign n1237 = pi030 & n283;
  assign n1238 = n253 & n1237;
  assign n1239 = n273 & n1238;
  assign n1240 = ~n262 & n1239;
  assign n1241 = ~n1231 & ~n1233;
  assign n1242 = ~n1236 & n1241;
  assign n1243 = ~n286 & ~n1240;
  assign n1244 = n1242 & n1243;
  assign n1245 = n679 & ~n1244;
  assign n1246 = n637 & ~n1244;
  assign n1247 = ~n679 & n1246;
  assign n1248 = ~n637 & ~n1244;
  assign n1249 = ~n679 & n1248;
  assign n1250 = n640 & n1249;
  assign n1251 = ~n640 & ~n1244;
  assign n1252 = ~n679 & n1251;
  assign n1253 = ~n637 & n1252;
  assign n1254 = n395 & n1253;
  assign n1255 = ~n395 & ~n1244;
  assign n1256 = ~n637 & n1255;
  assign n1257 = ~n679 & n1256;
  assign n1258 = ~n640 & n1257;
  assign n1259 = pi005 & n1258;
  assign n1260 = ~pi005 & pi117;
  assign n1261 = ~n640 & n1260;
  assign n1262 = ~n679 & n1261;
  assign n1263 = ~n637 & n1262;
  assign n1264 = ~n395 & n1263;
  assign n1265 = n228 & n1264;
  assign n1266 = pi073 & ~n228;
  assign n1267 = ~n395 & n1266;
  assign n1268 = ~n637 & n1267;
  assign n1269 = ~n679 & n1268;
  assign n1270 = ~n640 & n1269;
  assign n1271 = ~pi005 & n1270;
  assign n1272 = ~pi007 & n1271;
  assign n1273 = ~pi095 & n1272;
  assign n1274 = ~pi130 & n1273;
  assign n1275 = ~pi000 & n1274;
  assign n1276 = pi002 & n1275;
  assign n1277 = pi001 & n1276;
  assign n1278 = ~pi005 & n1277;
  assign n1279 = ~n1245 & ~n1247;
  assign n1280 = ~n1250 & ~n1254;
  assign n1281 = n1279 & n1280;
  assign n1282 = ~n1259 & ~n1265;
  assign n1283 = ~n1278 & n1282;
  assign po23 = ~n1281 | ~n1283;
  assign n1285 = pi016 & ~n253;
  assign n1286 = pi024 & ~n273;
  assign n1287 = n253 & n1286;
  assign n1288 = pi027 & n273;
  assign n1289 = n253 & n1288;
  assign n1290 = ~n283 & n1289;
  assign n1291 = pi031 & n283;
  assign n1292 = n253 & n1291;
  assign n1293 = n273 & n1292;
  assign n1294 = ~n262 & n1293;
  assign n1295 = ~n1285 & ~n1287;
  assign n1296 = ~n1290 & n1295;
  assign n1297 = ~n286 & ~n1294;
  assign n1298 = n1296 & n1297;
  assign n1299 = n679 & ~n1298;
  assign n1300 = n637 & ~n1298;
  assign n1301 = ~n679 & n1300;
  assign n1302 = ~n637 & ~n1298;
  assign n1303 = ~n679 & n1302;
  assign n1304 = n640 & n1303;
  assign n1305 = ~n640 & ~n1298;
  assign n1306 = ~n679 & n1305;
  assign n1307 = ~n637 & n1306;
  assign n1308 = n395 & n1307;
  assign n1309 = ~n395 & ~n1298;
  assign n1310 = ~n637 & n1309;
  assign n1311 = ~n679 & n1310;
  assign n1312 = ~n640 & n1311;
  assign n1313 = pi005 & n1312;
  assign n1314 = ~pi005 & pi118;
  assign n1315 = ~n640 & n1314;
  assign n1316 = ~n679 & n1315;
  assign n1317 = ~n637 & n1316;
  assign n1318 = ~n395 & n1317;
  assign n1319 = n228 & n1318;
  assign n1320 = pi074 & ~n228;
  assign n1321 = ~n395 & n1320;
  assign n1322 = ~n637 & n1321;
  assign n1323 = ~n679 & n1322;
  assign n1324 = ~n640 & n1323;
  assign n1325 = ~pi005 & n1324;
  assign n1326 = ~pi007 & n1325;
  assign n1327 = ~pi095 & n1326;
  assign n1328 = ~pi130 & n1327;
  assign n1329 = ~pi000 & n1328;
  assign n1330 = pi002 & n1329;
  assign n1331 = pi001 & n1330;
  assign n1332 = ~pi005 & n1331;
  assign n1333 = ~n1299 & ~n1301;
  assign n1334 = ~n1304 & ~n1308;
  assign n1335 = n1333 & n1334;
  assign n1336 = ~n1313 & ~n1319;
  assign n1337 = ~n1332 & n1336;
  assign po24 = ~n1335 | ~n1337;
  assign n1339 = pi017 & ~n253;
  assign n1340 = pi025 & ~n273;
  assign n1341 = n253 & n1340;
  assign n1342 = pi028 & n273;
  assign n1343 = n253 & n1342;
  assign n1344 = ~n283 & n1343;
  assign n1345 = pi032 & n283;
  assign n1346 = n253 & n1345;
  assign n1347 = n273 & n1346;
  assign n1348 = ~n262 & n1347;
  assign n1349 = ~n1339 & ~n1341;
  assign n1350 = ~n1344 & n1349;
  assign n1351 = ~n286 & ~n1348;
  assign n1352 = n1350 & n1351;
  assign n1353 = n679 & ~n1352;
  assign n1354 = n637 & ~n1352;
  assign n1355 = ~n679 & n1354;
  assign n1356 = ~n637 & ~n1352;
  assign n1357 = ~n679 & n1356;
  assign n1358 = n640 & n1357;
  assign n1359 = ~n640 & ~n1352;
  assign n1360 = ~n679 & n1359;
  assign n1361 = ~n637 & n1360;
  assign n1362 = n395 & n1361;
  assign n1363 = ~n395 & ~n1352;
  assign n1364 = ~n637 & n1363;
  assign n1365 = ~n679 & n1364;
  assign n1366 = ~n640 & n1365;
  assign n1367 = pi005 & n1366;
  assign n1368 = ~pi005 & pi119;
  assign n1369 = ~n640 & n1368;
  assign n1370 = ~n679 & n1369;
  assign n1371 = ~n637 & n1370;
  assign n1372 = ~n395 & n1371;
  assign n1373 = n228 & n1372;
  assign n1374 = pi075 & ~n228;
  assign n1375 = ~n395 & n1374;
  assign n1376 = ~n637 & n1375;
  assign n1377 = ~n679 & n1376;
  assign n1378 = ~n640 & n1377;
  assign n1379 = ~pi005 & n1378;
  assign n1380 = ~pi007 & n1379;
  assign n1381 = ~pi095 & n1380;
  assign n1382 = ~pi130 & n1381;
  assign n1383 = ~pi000 & n1382;
  assign n1384 = pi002 & n1383;
  assign n1385 = pi001 & n1384;
  assign n1386 = ~pi005 & n1385;
  assign n1387 = ~n1353 & ~n1355;
  assign n1388 = ~n1358 & ~n1362;
  assign n1389 = n1387 & n1388;
  assign n1390 = ~n1367 & ~n1373;
  assign n1391 = ~n1386 & n1390;
  assign po25 = ~n1389 | ~n1391;
  assign n1393 = pi018 & ~n253;
  assign n1394 = pi026 & ~n273;
  assign n1395 = n253 & n1394;
  assign n1396 = pi029 & n273;
  assign n1397 = n253 & n1396;
  assign n1398 = ~n283 & n1397;
  assign n1399 = pi033 & n283;
  assign n1400 = n253 & n1399;
  assign n1401 = n273 & n1400;
  assign n1402 = ~n262 & n1401;
  assign n1403 = ~n1393 & ~n1395;
  assign n1404 = ~n1398 & n1403;
  assign n1405 = ~n286 & ~n1402;
  assign n1406 = n1404 & n1405;
  assign n1407 = n679 & ~n1406;
  assign n1408 = n637 & ~n1406;
  assign n1409 = ~n679 & n1408;
  assign n1410 = ~n637 & ~n1406;
  assign n1411 = ~n679 & n1410;
  assign n1412 = n640 & n1411;
  assign n1413 = ~n640 & ~n1406;
  assign n1414 = ~n679 & n1413;
  assign n1415 = ~n637 & n1414;
  assign n1416 = n395 & n1415;
  assign n1417 = ~n395 & ~n1406;
  assign n1418 = ~n637 & n1417;
  assign n1419 = ~n679 & n1418;
  assign n1420 = ~n640 & n1419;
  assign n1421 = pi005 & n1420;
  assign n1422 = ~pi005 & pi120;
  assign n1423 = ~n640 & n1422;
  assign n1424 = ~n679 & n1423;
  assign n1425 = ~n637 & n1424;
  assign n1426 = ~n395 & n1425;
  assign n1427 = n228 & n1426;
  assign n1428 = pi076 & ~n228;
  assign n1429 = ~n395 & n1428;
  assign n1430 = ~n637 & n1429;
  assign n1431 = ~n679 & n1430;
  assign n1432 = ~n640 & n1431;
  assign n1433 = ~pi005 & n1432;
  assign n1434 = ~pi007 & n1433;
  assign n1435 = ~pi095 & n1434;
  assign n1436 = ~pi130 & n1435;
  assign n1437 = ~pi000 & n1436;
  assign n1438 = pi002 & n1437;
  assign n1439 = pi001 & n1438;
  assign n1440 = ~pi005 & n1439;
  assign n1441 = ~n1407 & ~n1409;
  assign n1442 = ~n1412 & ~n1416;
  assign n1443 = n1441 & n1442;
  assign n1444 = ~n1421 & ~n1427;
  assign n1445 = ~n1440 & n1444;
  assign po26 = ~n1443 | ~n1445;
  assign n1447 = pi019 & ~n253;
  assign n1448 = pi027 & ~n273;
  assign n1449 = n253 & n1448;
  assign n1450 = pi030 & n273;
  assign n1451 = n253 & n1450;
  assign n1452 = ~n283 & n1451;
  assign n1453 = pi034 & n283;
  assign n1454 = n253 & n1453;
  assign n1455 = n273 & n1454;
  assign n1456 = ~n262 & n1455;
  assign n1457 = ~n1447 & ~n1449;
  assign n1458 = ~n1452 & n1457;
  assign n1459 = ~n286 & ~n1456;
  assign n1460 = n1458 & n1459;
  assign n1461 = n679 & ~n1460;
  assign n1462 = n637 & ~n1460;
  assign n1463 = ~n679 & n1462;
  assign n1464 = ~n637 & ~n1460;
  assign n1465 = ~n679 & n1464;
  assign n1466 = n640 & n1465;
  assign n1467 = ~n640 & ~n1460;
  assign n1468 = ~n679 & n1467;
  assign n1469 = ~n637 & n1468;
  assign n1470 = n395 & n1469;
  assign n1471 = ~n395 & ~n1460;
  assign n1472 = ~n637 & n1471;
  assign n1473 = ~n679 & n1472;
  assign n1474 = ~n640 & n1473;
  assign n1475 = pi005 & n1474;
  assign n1476 = ~pi005 & pi121;
  assign n1477 = ~n640 & n1476;
  assign n1478 = ~n679 & n1477;
  assign n1479 = ~n637 & n1478;
  assign n1480 = ~n395 & n1479;
  assign n1481 = n228 & n1480;
  assign n1482 = pi077 & ~n228;
  assign n1483 = ~n395 & n1482;
  assign n1484 = ~n637 & n1483;
  assign n1485 = ~n679 & n1484;
  assign n1486 = ~n640 & n1485;
  assign n1487 = ~pi005 & n1486;
  assign n1488 = ~pi007 & n1487;
  assign n1489 = ~pi095 & n1488;
  assign n1490 = ~pi130 & n1489;
  assign n1491 = ~pi000 & n1490;
  assign n1492 = pi002 & n1491;
  assign n1493 = pi001 & n1492;
  assign n1494 = ~pi005 & n1493;
  assign n1495 = ~n1461 & ~n1463;
  assign n1496 = ~n1466 & ~n1470;
  assign n1497 = n1495 & n1496;
  assign n1498 = ~n1475 & ~n1481;
  assign n1499 = ~n1494 & n1498;
  assign po27 = ~n1497 | ~n1499;
  assign n1501 = pi020 & ~n253;
  assign n1502 = pi028 & ~n273;
  assign n1503 = n253 & n1502;
  assign n1504 = pi031 & n273;
  assign n1505 = n253 & n1504;
  assign n1506 = ~n283 & n1505;
  assign n1507 = pi035 & n283;
  assign n1508 = n253 & n1507;
  assign n1509 = n273 & n1508;
  assign n1510 = ~n262 & n1509;
  assign n1511 = ~n1501 & ~n1503;
  assign n1512 = ~n1506 & n1511;
  assign n1513 = ~n286 & ~n1510;
  assign n1514 = n1512 & n1513;
  assign n1515 = n679 & ~n1514;
  assign n1516 = n637 & ~n1514;
  assign n1517 = ~n679 & n1516;
  assign n1518 = ~n637 & ~n1514;
  assign n1519 = ~n679 & n1518;
  assign n1520 = n640 & n1519;
  assign n1521 = ~n640 & ~n1514;
  assign n1522 = ~n679 & n1521;
  assign n1523 = ~n637 & n1522;
  assign n1524 = n395 & n1523;
  assign n1525 = ~n395 & ~n1514;
  assign n1526 = ~n637 & n1525;
  assign n1527 = ~n679 & n1526;
  assign n1528 = ~n640 & n1527;
  assign n1529 = pi005 & n1528;
  assign n1530 = ~pi005 & pi122;
  assign n1531 = ~n640 & n1530;
  assign n1532 = ~n679 & n1531;
  assign n1533 = ~n637 & n1532;
  assign n1534 = ~n395 & n1533;
  assign n1535 = n228 & n1534;
  assign n1536 = pi078 & ~n228;
  assign n1537 = ~n395 & n1536;
  assign n1538 = ~n637 & n1537;
  assign n1539 = ~n679 & n1538;
  assign n1540 = ~n640 & n1539;
  assign n1541 = ~pi005 & n1540;
  assign n1542 = ~pi007 & n1541;
  assign n1543 = ~pi095 & n1542;
  assign n1544 = ~pi130 & n1543;
  assign n1545 = ~pi000 & n1544;
  assign n1546 = pi002 & n1545;
  assign n1547 = pi001 & n1546;
  assign n1548 = ~pi005 & n1547;
  assign n1549 = ~n1515 & ~n1517;
  assign n1550 = ~n1520 & ~n1524;
  assign n1551 = n1549 & n1550;
  assign n1552 = ~n1529 & ~n1535;
  assign n1553 = ~n1548 & n1552;
  assign po28 = ~n1551 | ~n1553;
  assign n1555 = pi021 & ~n253;
  assign n1556 = pi029 & ~n273;
  assign n1557 = n253 & n1556;
  assign n1558 = pi032 & n273;
  assign n1559 = n253 & n1558;
  assign n1560 = ~n283 & n1559;
  assign n1561 = pi036 & n283;
  assign n1562 = n253 & n1561;
  assign n1563 = n273 & n1562;
  assign n1564 = ~n262 & n1563;
  assign n1565 = ~n1555 & ~n1557;
  assign n1566 = ~n1560 & n1565;
  assign n1567 = ~n286 & ~n1564;
  assign n1568 = n1566 & n1567;
  assign n1569 = n679 & ~n1568;
  assign n1570 = n637 & ~n1568;
  assign n1571 = ~n679 & n1570;
  assign n1572 = ~n637 & ~n1568;
  assign n1573 = ~n679 & n1572;
  assign n1574 = n640 & n1573;
  assign n1575 = ~n640 & ~n1568;
  assign n1576 = ~n679 & n1575;
  assign n1577 = ~n637 & n1576;
  assign n1578 = n395 & n1577;
  assign n1579 = ~n395 & ~n1568;
  assign n1580 = ~n637 & n1579;
  assign n1581 = ~n679 & n1580;
  assign n1582 = ~n640 & n1581;
  assign n1583 = pi005 & n1582;
  assign n1584 = ~pi005 & pi123;
  assign n1585 = ~n640 & n1584;
  assign n1586 = ~n679 & n1585;
  assign n1587 = ~n637 & n1586;
  assign n1588 = ~n395 & n1587;
  assign n1589 = n228 & n1588;
  assign n1590 = pi079 & ~n228;
  assign n1591 = ~n395 & n1590;
  assign n1592 = ~n637 & n1591;
  assign n1593 = ~n679 & n1592;
  assign n1594 = ~n640 & n1593;
  assign n1595 = ~pi005 & n1594;
  assign n1596 = ~pi007 & n1595;
  assign n1597 = ~pi095 & n1596;
  assign n1598 = ~pi130 & n1597;
  assign n1599 = ~pi000 & n1598;
  assign n1600 = pi002 & n1599;
  assign n1601 = pi001 & n1600;
  assign n1602 = ~pi005 & n1601;
  assign n1603 = ~n1569 & ~n1571;
  assign n1604 = ~n1574 & ~n1578;
  assign n1605 = n1603 & n1604;
  assign n1606 = ~n1583 & ~n1589;
  assign n1607 = ~n1602 & n1606;
  assign po29 = ~n1605 | ~n1607;
  assign n1609 = pi022 & ~n253;
  assign n1610 = pi030 & ~n273;
  assign n1611 = n253 & n1610;
  assign n1612 = pi033 & n273;
  assign n1613 = n253 & n1612;
  assign n1614 = ~n283 & n1613;
  assign n1615 = pi037 & n283;
  assign n1616 = n253 & n1615;
  assign n1617 = n273 & n1616;
  assign n1618 = ~n262 & n1617;
  assign n1619 = ~n1609 & ~n1611;
  assign n1620 = ~n1614 & n1619;
  assign n1621 = ~n286 & ~n1618;
  assign n1622 = n1620 & n1621;
  assign n1623 = n679 & ~n1622;
  assign n1624 = n637 & ~n1622;
  assign n1625 = ~n679 & n1624;
  assign n1626 = ~n637 & ~n1622;
  assign n1627 = ~n679 & n1626;
  assign n1628 = n640 & n1627;
  assign n1629 = ~n640 & ~n1622;
  assign n1630 = ~n679 & n1629;
  assign n1631 = ~n637 & n1630;
  assign n1632 = n395 & n1631;
  assign n1633 = ~n395 & ~n1622;
  assign n1634 = ~n637 & n1633;
  assign n1635 = ~n679 & n1634;
  assign n1636 = ~n640 & n1635;
  assign n1637 = pi005 & n1636;
  assign n1638 = ~pi005 & pi124;
  assign n1639 = ~n640 & n1638;
  assign n1640 = ~n679 & n1639;
  assign n1641 = ~n637 & n1640;
  assign n1642 = ~n395 & n1641;
  assign n1643 = n228 & n1642;
  assign n1644 = pi080 & ~n228;
  assign n1645 = ~n395 & n1644;
  assign n1646 = ~n637 & n1645;
  assign n1647 = ~n679 & n1646;
  assign n1648 = ~n640 & n1647;
  assign n1649 = ~pi005 & n1648;
  assign n1650 = ~pi007 & n1649;
  assign n1651 = ~pi095 & n1650;
  assign n1652 = ~pi130 & n1651;
  assign n1653 = ~pi000 & n1652;
  assign n1654 = pi002 & n1653;
  assign n1655 = pi001 & n1654;
  assign n1656 = ~pi005 & n1655;
  assign n1657 = ~n1623 & ~n1625;
  assign n1658 = ~n1628 & ~n1632;
  assign n1659 = n1657 & n1658;
  assign n1660 = ~n1637 & ~n1643;
  assign n1661 = ~n1656 & n1660;
  assign po30 = ~n1659 | ~n1661;
  assign n1663 = pi023 & ~n253;
  assign n1664 = pi031 & ~n273;
  assign n1665 = n253 & n1664;
  assign n1666 = pi034 & n273;
  assign n1667 = n253 & n1666;
  assign n1668 = ~n283 & n1667;
  assign n1669 = pi038 & n283;
  assign n1670 = n253 & n1669;
  assign n1671 = n273 & n1670;
  assign n1672 = ~n262 & n1671;
  assign n1673 = ~n1663 & ~n1665;
  assign n1674 = ~n1668 & n1673;
  assign n1675 = ~n286 & ~n1672;
  assign n1676 = n1674 & n1675;
  assign n1677 = n679 & ~n1676;
  assign n1678 = n637 & ~n1676;
  assign n1679 = ~n679 & n1678;
  assign n1680 = ~n637 & ~n1676;
  assign n1681 = ~n679 & n1680;
  assign n1682 = n640 & n1681;
  assign n1683 = ~n640 & ~n1676;
  assign n1684 = ~n679 & n1683;
  assign n1685 = ~n637 & n1684;
  assign n1686 = n395 & n1685;
  assign n1687 = ~n395 & ~n1676;
  assign n1688 = ~n637 & n1687;
  assign n1689 = ~n679 & n1688;
  assign n1690 = ~n640 & n1689;
  assign n1691 = pi005 & n1690;
  assign n1692 = ~pi005 & pi125;
  assign n1693 = ~n640 & n1692;
  assign n1694 = ~n679 & n1693;
  assign n1695 = ~n637 & n1694;
  assign n1696 = ~n395 & n1695;
  assign n1697 = n228 & n1696;
  assign n1698 = pi081 & ~n228;
  assign n1699 = ~n395 & n1698;
  assign n1700 = ~n637 & n1699;
  assign n1701 = ~n679 & n1700;
  assign n1702 = ~n640 & n1701;
  assign n1703 = ~pi005 & n1702;
  assign n1704 = ~pi007 & n1703;
  assign n1705 = ~pi095 & n1704;
  assign n1706 = ~pi130 & n1705;
  assign n1707 = ~pi000 & n1706;
  assign n1708 = pi002 & n1707;
  assign n1709 = pi001 & n1708;
  assign n1710 = ~pi005 & n1709;
  assign n1711 = ~n1677 & ~n1679;
  assign n1712 = ~n1682 & ~n1686;
  assign n1713 = n1711 & n1712;
  assign n1714 = ~n1691 & ~n1697;
  assign n1715 = ~n1710 & n1714;
  assign po31 = ~n1713 | ~n1715;
  assign n1717 = ~pi004 & n678;
  assign n1718 = ~pi130 & n1717;
  assign n1719 = pi067 & ~n253;
  assign n1720 = pi075 & ~n273;
  assign n1721 = n253 & n1720;
  assign n1722 = pi078 & n273;
  assign n1723 = n253 & n1722;
  assign n1724 = ~n283 & n1723;
  assign n1725 = pi082 & n283;
  assign n1726 = n253 & n1725;
  assign n1727 = n273 & n1726;
  assign n1728 = ~n262 & n1727;
  assign n1729 = ~n1719 & ~n1721;
  assign n1730 = ~n1724 & n1729;
  assign n1731 = ~n286 & ~n1728;
  assign n1732 = n1730 & n1731;
  assign n1733 = n1718 & ~n1732;
  assign n1734 = ~pi001 & pi003;
  assign n1735 = ~pi131 & n1734;
  assign n1736 = ~pi095 & n1735;
  assign n1737 = pi004 & n1736;
  assign n1738 = ~n1732 & n1737;
  assign n1739 = ~n1718 & n1738;
  assign n1740 = ~pi001 & ~pi003;
  assign n1741 = ~pi095 & n1740;
  assign n1742 = pi004 & n1741;
  assign n1743 = ~n1732 & ~n1737;
  assign n1744 = ~n1718 & n1743;
  assign n1745 = n1742 & n1744;
  assign n1746 = pi000 & n248;
  assign n1747 = ~pi130 & n1746;
  assign n1748 = ~pi006 & n1747;
  assign n1749 = ~n1732 & ~n1742;
  assign n1750 = ~n1718 & n1749;
  assign n1751 = ~n1737 & n1750;
  assign n1752 = n1748 & n1751;
  assign n1753 = pi007 & n619;
  assign n1754 = ~n1732 & ~n1748;
  assign n1755 = ~n1737 & n1754;
  assign n1756 = ~n1718 & n1755;
  assign n1757 = ~n1742 & n1756;
  assign n1758 = n1753 & n1757;
  assign n1759 = ~n1732 & ~n1753;
  assign n1760 = ~n1742 & n1759;
  assign n1761 = ~n1718 & n1760;
  assign n1762 = ~n1737 & n1761;
  assign n1763 = ~n1748 & n1762;
  assign n1764 = pi005 & n1763;
  assign n1765 = n936 & ~n1748;
  assign n1766 = ~n1737 & n1765;
  assign n1767 = ~n1718 & n1766;
  assign n1768 = ~n1742 & n1767;
  assign n1769 = ~n1753 & n1768;
  assign n1770 = pi095 & n1769;
  assign n1771 = ~pi005 & n1770;
  assign n1772 = ~n1733 & ~n1739;
  assign n1773 = ~n1745 & ~n1752;
  assign n1774 = n1772 & n1773;
  assign n1775 = ~n1758 & ~n1764;
  assign n1776 = ~n1771 & n1775;
  assign po32 = ~n1774 | ~n1776;
  assign n1778 = pi068 & ~n253;
  assign n1779 = pi076 & ~n273;
  assign n1780 = n253 & n1779;
  assign n1781 = pi079 & n273;
  assign n1782 = n253 & n1781;
  assign n1783 = ~n283 & n1782;
  assign n1784 = pi083 & n283;
  assign n1785 = n253 & n1784;
  assign n1786 = n273 & n1785;
  assign n1787 = ~n262 & n1786;
  assign n1788 = ~n1778 & ~n1780;
  assign n1789 = ~n1783 & n1788;
  assign n1790 = ~n286 & ~n1787;
  assign n1791 = n1789 & n1790;
  assign n1792 = n1718 & ~n1791;
  assign n1793 = n1737 & ~n1791;
  assign n1794 = ~n1718 & n1793;
  assign n1795 = ~n1737 & ~n1791;
  assign n1796 = ~n1718 & n1795;
  assign n1797 = n1742 & n1796;
  assign n1798 = ~n1742 & ~n1791;
  assign n1799 = ~n1718 & n1798;
  assign n1800 = ~n1737 & n1799;
  assign n1801 = n1748 & n1800;
  assign n1802 = ~n1748 & ~n1791;
  assign n1803 = ~n1737 & n1802;
  assign n1804 = ~n1718 & n1803;
  assign n1805 = ~n1742 & n1804;
  assign n1806 = n1753 & n1805;
  assign n1807 = ~n1753 & ~n1791;
  assign n1808 = ~n1742 & n1807;
  assign n1809 = ~n1718 & n1808;
  assign n1810 = ~n1737 & n1809;
  assign n1811 = ~n1748 & n1810;
  assign n1812 = pi005 & n1811;
  assign n1813 = n990 & ~n1748;
  assign n1814 = ~n1737 & n1813;
  assign n1815 = ~n1718 & n1814;
  assign n1816 = ~n1742 & n1815;
  assign n1817 = ~n1753 & n1816;
  assign n1818 = pi095 & n1817;
  assign n1819 = ~pi005 & n1818;
  assign n1820 = ~n1792 & ~n1794;
  assign n1821 = ~n1797 & ~n1801;
  assign n1822 = n1820 & n1821;
  assign n1823 = ~n1806 & ~n1812;
  assign n1824 = ~n1819 & n1823;
  assign po33 = ~n1822 | ~n1824;
  assign n1826 = pi069 & ~n253;
  assign n1827 = pi077 & ~n273;
  assign n1828 = n253 & n1827;
  assign n1829 = pi080 & n273;
  assign n1830 = n253 & n1829;
  assign n1831 = ~n283 & n1830;
  assign n1832 = pi084 & n283;
  assign n1833 = n253 & n1832;
  assign n1834 = n273 & n1833;
  assign n1835 = ~n262 & n1834;
  assign n1836 = ~n1826 & ~n1828;
  assign n1837 = ~n1831 & n1836;
  assign n1838 = ~n286 & ~n1835;
  assign n1839 = n1837 & n1838;
  assign n1840 = n1718 & ~n1839;
  assign n1841 = n1737 & ~n1839;
  assign n1842 = ~n1718 & n1841;
  assign n1843 = ~n1737 & ~n1839;
  assign n1844 = ~n1718 & n1843;
  assign n1845 = n1742 & n1844;
  assign n1846 = ~n1742 & ~n1839;
  assign n1847 = ~n1718 & n1846;
  assign n1848 = ~n1737 & n1847;
  assign n1849 = n1748 & n1848;
  assign n1850 = ~n1748 & ~n1839;
  assign n1851 = ~n1737 & n1850;
  assign n1852 = ~n1718 & n1851;
  assign n1853 = ~n1742 & n1852;
  assign n1854 = n1753 & n1853;
  assign n1855 = ~n1753 & ~n1839;
  assign n1856 = ~n1742 & n1855;
  assign n1857 = ~n1718 & n1856;
  assign n1858 = ~n1737 & n1857;
  assign n1859 = ~n1748 & n1858;
  assign n1860 = pi005 & n1859;
  assign n1861 = n1044 & ~n1748;
  assign n1862 = ~n1737 & n1861;
  assign n1863 = ~n1718 & n1862;
  assign n1864 = ~n1742 & n1863;
  assign n1865 = ~n1753 & n1864;
  assign n1866 = pi095 & n1865;
  assign n1867 = ~pi005 & n1866;
  assign n1868 = ~n1840 & ~n1842;
  assign n1869 = ~n1845 & ~n1849;
  assign n1870 = n1868 & n1869;
  assign n1871 = ~n1854 & ~n1860;
  assign n1872 = ~n1867 & n1871;
  assign po34 = ~n1870 | ~n1872;
  assign n1874 = pi070 & ~n253;
  assign n1875 = pi078 & ~n273;
  assign n1876 = n253 & n1875;
  assign n1877 = pi081 & n273;
  assign n1878 = n253 & n1877;
  assign n1879 = ~n283 & n1878;
  assign n1880 = pi085 & n283;
  assign n1881 = n253 & n1880;
  assign n1882 = n273 & n1881;
  assign n1883 = ~n262 & n1882;
  assign n1884 = ~n1874 & ~n1876;
  assign n1885 = ~n1879 & n1884;
  assign n1886 = ~n286 & ~n1883;
  assign n1887 = n1885 & n1886;
  assign n1888 = n1718 & ~n1887;
  assign n1889 = n1737 & ~n1887;
  assign n1890 = ~n1718 & n1889;
  assign n1891 = ~n1737 & ~n1887;
  assign n1892 = ~n1718 & n1891;
  assign n1893 = n1742 & n1892;
  assign n1894 = ~n1742 & ~n1887;
  assign n1895 = ~n1718 & n1894;
  assign n1896 = ~n1737 & n1895;
  assign n1897 = n1748 & n1896;
  assign n1898 = ~n1748 & ~n1887;
  assign n1899 = ~n1737 & n1898;
  assign n1900 = ~n1718 & n1899;
  assign n1901 = ~n1742 & n1900;
  assign n1902 = n1753 & n1901;
  assign n1903 = ~n1753 & ~n1887;
  assign n1904 = ~n1742 & n1903;
  assign n1905 = ~n1718 & n1904;
  assign n1906 = ~n1737 & n1905;
  assign n1907 = ~n1748 & n1906;
  assign n1908 = pi005 & n1907;
  assign n1909 = n1098 & ~n1748;
  assign n1910 = ~n1737 & n1909;
  assign n1911 = ~n1718 & n1910;
  assign n1912 = ~n1742 & n1911;
  assign n1913 = ~n1753 & n1912;
  assign n1914 = pi095 & n1913;
  assign n1915 = ~pi005 & n1914;
  assign n1916 = ~n1888 & ~n1890;
  assign n1917 = ~n1893 & ~n1897;
  assign n1918 = n1916 & n1917;
  assign n1919 = ~n1902 & ~n1908;
  assign n1920 = ~n1915 & n1919;
  assign po35 = ~n1918 | ~n1920;
  assign n1922 = pi071 & ~n253;
  assign n1923 = pi079 & ~n273;
  assign n1924 = n253 & n1923;
  assign n1925 = pi082 & n273;
  assign n1926 = n253 & n1925;
  assign n1927 = ~n283 & n1926;
  assign n1928 = pi086 & n283;
  assign n1929 = n253 & n1928;
  assign n1930 = n273 & n1929;
  assign n1931 = ~n262 & n1930;
  assign n1932 = ~n1922 & ~n1924;
  assign n1933 = ~n1927 & n1932;
  assign n1934 = ~n286 & ~n1931;
  assign n1935 = n1933 & n1934;
  assign n1936 = n1718 & ~n1935;
  assign n1937 = n1737 & ~n1935;
  assign n1938 = ~n1718 & n1937;
  assign n1939 = ~n1737 & ~n1935;
  assign n1940 = ~n1718 & n1939;
  assign n1941 = n1742 & n1940;
  assign n1942 = ~n1742 & ~n1935;
  assign n1943 = ~n1718 & n1942;
  assign n1944 = ~n1737 & n1943;
  assign n1945 = n1748 & n1944;
  assign n1946 = ~n1748 & ~n1935;
  assign n1947 = ~n1737 & n1946;
  assign n1948 = ~n1718 & n1947;
  assign n1949 = ~n1742 & n1948;
  assign n1950 = n1753 & n1949;
  assign n1951 = ~n1753 & ~n1935;
  assign n1952 = ~n1742 & n1951;
  assign n1953 = ~n1718 & n1952;
  assign n1954 = ~n1737 & n1953;
  assign n1955 = ~n1748 & n1954;
  assign n1956 = pi005 & n1955;
  assign n1957 = n1152 & ~n1748;
  assign n1958 = ~n1737 & n1957;
  assign n1959 = ~n1718 & n1958;
  assign n1960 = ~n1742 & n1959;
  assign n1961 = ~n1753 & n1960;
  assign n1962 = pi095 & n1961;
  assign n1963 = ~pi005 & n1962;
  assign n1964 = ~n1936 & ~n1938;
  assign n1965 = ~n1941 & ~n1945;
  assign n1966 = n1964 & n1965;
  assign n1967 = ~n1950 & ~n1956;
  assign n1968 = ~n1963 & n1967;
  assign po36 = ~n1966 | ~n1968;
  assign n1970 = pi072 & ~n253;
  assign n1971 = pi080 & ~n273;
  assign n1972 = n253 & n1971;
  assign n1973 = pi083 & n273;
  assign n1974 = n253 & n1973;
  assign n1975 = ~n283 & n1974;
  assign n1976 = pi041 & n283;
  assign n1977 = n253 & n1976;
  assign n1978 = n273 & n1977;
  assign n1979 = ~n262 & n1978;
  assign n1980 = ~n1970 & ~n1972;
  assign n1981 = ~n1975 & n1980;
  assign n1982 = ~n286 & ~n1979;
  assign n1983 = n1981 & n1982;
  assign n1984 = n1718 & ~n1983;
  assign n1985 = n1737 & ~n1983;
  assign n1986 = ~n1718 & n1985;
  assign n1987 = ~n1737 & ~n1983;
  assign n1988 = ~n1718 & n1987;
  assign n1989 = n1742 & n1988;
  assign n1990 = ~n1742 & ~n1983;
  assign n1991 = ~n1718 & n1990;
  assign n1992 = ~n1737 & n1991;
  assign n1993 = n1748 & n1992;
  assign n1994 = ~n1748 & ~n1983;
  assign n1995 = ~n1737 & n1994;
  assign n1996 = ~n1718 & n1995;
  assign n1997 = ~n1742 & n1996;
  assign n1998 = n1753 & n1997;
  assign n1999 = ~n1753 & ~n1983;
  assign n2000 = ~n1742 & n1999;
  assign n2001 = ~n1718 & n2000;
  assign n2002 = ~n1737 & n2001;
  assign n2003 = ~n1748 & n2002;
  assign n2004 = pi005 & n2003;
  assign n2005 = n1206 & ~n1748;
  assign n2006 = ~n1737 & n2005;
  assign n2007 = ~n1718 & n2006;
  assign n2008 = ~n1742 & n2007;
  assign n2009 = ~n1753 & n2008;
  assign n2010 = pi095 & n2009;
  assign n2011 = ~pi005 & n2010;
  assign n2012 = ~n1984 & ~n1986;
  assign n2013 = ~n1989 & ~n1993;
  assign n2014 = n2012 & n2013;
  assign n2015 = ~n1998 & ~n2004;
  assign n2016 = ~n2011 & n2015;
  assign po37 = ~n2014 | ~n2016;
  assign n2018 = pi073 & ~n253;
  assign n2019 = pi081 & ~n273;
  assign n2020 = n253 & n2019;
  assign n2021 = pi084 & n273;
  assign n2022 = n253 & n2021;
  assign n2023 = ~n283 & n2022;
  assign n2024 = pi042 & n283;
  assign n2025 = n253 & n2024;
  assign n2026 = n273 & n2025;
  assign n2027 = ~n262 & n2026;
  assign n2028 = ~n2018 & ~n2020;
  assign n2029 = ~n2023 & n2028;
  assign n2030 = ~n286 & ~n2027;
  assign n2031 = n2029 & n2030;
  assign n2032 = n1718 & ~n2031;
  assign n2033 = n1737 & ~n2031;
  assign n2034 = ~n1718 & n2033;
  assign n2035 = ~n1737 & ~n2031;
  assign n2036 = ~n1718 & n2035;
  assign n2037 = n1742 & n2036;
  assign n2038 = ~n1742 & ~n2031;
  assign n2039 = ~n1718 & n2038;
  assign n2040 = ~n1737 & n2039;
  assign n2041 = n1748 & n2040;
  assign n2042 = ~n1748 & ~n2031;
  assign n2043 = ~n1737 & n2042;
  assign n2044 = ~n1718 & n2043;
  assign n2045 = ~n1742 & n2044;
  assign n2046 = n1753 & n2045;
  assign n2047 = ~n1753 & ~n2031;
  assign n2048 = ~n1742 & n2047;
  assign n2049 = ~n1718 & n2048;
  assign n2050 = ~n1737 & n2049;
  assign n2051 = ~n1748 & n2050;
  assign n2052 = pi005 & n2051;
  assign n2053 = n1260 & ~n1748;
  assign n2054 = ~n1737 & n2053;
  assign n2055 = ~n1718 & n2054;
  assign n2056 = ~n1742 & n2055;
  assign n2057 = ~n1753 & n2056;
  assign n2058 = pi095 & n2057;
  assign n2059 = ~pi005 & n2058;
  assign n2060 = ~n2032 & ~n2034;
  assign n2061 = ~n2037 & ~n2041;
  assign n2062 = n2060 & n2061;
  assign n2063 = ~n2046 & ~n2052;
  assign n2064 = ~n2059 & n2063;
  assign po38 = ~n2062 | ~n2064;
  assign n2066 = pi074 & ~n253;
  assign n2067 = pi082 & ~n273;
  assign n2068 = n253 & n2067;
  assign n2069 = pi085 & n273;
  assign n2070 = n253 & n2069;
  assign n2071 = ~n283 & n2070;
  assign n2072 = pi043 & n283;
  assign n2073 = n253 & n2072;
  assign n2074 = n273 & n2073;
  assign n2075 = ~n262 & n2074;
  assign n2076 = ~n2066 & ~n2068;
  assign n2077 = ~n2071 & n2076;
  assign n2078 = ~n286 & ~n2075;
  assign n2079 = n2077 & n2078;
  assign n2080 = n1718 & ~n2079;
  assign n2081 = n1737 & ~n2079;
  assign n2082 = ~n1718 & n2081;
  assign n2083 = ~n1737 & ~n2079;
  assign n2084 = ~n1718 & n2083;
  assign n2085 = n1742 & n2084;
  assign n2086 = ~n1742 & ~n2079;
  assign n2087 = ~n1718 & n2086;
  assign n2088 = ~n1737 & n2087;
  assign n2089 = n1748 & n2088;
  assign n2090 = ~n1748 & ~n2079;
  assign n2091 = ~n1737 & n2090;
  assign n2092 = ~n1718 & n2091;
  assign n2093 = ~n1742 & n2092;
  assign n2094 = n1753 & n2093;
  assign n2095 = ~n1753 & ~n2079;
  assign n2096 = ~n1742 & n2095;
  assign n2097 = ~n1718 & n2096;
  assign n2098 = ~n1737 & n2097;
  assign n2099 = ~n1748 & n2098;
  assign n2100 = pi005 & n2099;
  assign n2101 = n1314 & ~n1748;
  assign n2102 = ~n1737 & n2101;
  assign n2103 = ~n1718 & n2102;
  assign n2104 = ~n1742 & n2103;
  assign n2105 = ~n1753 & n2104;
  assign n2106 = pi095 & n2105;
  assign n2107 = ~pi005 & n2106;
  assign n2108 = ~n2080 & ~n2082;
  assign n2109 = ~n2085 & ~n2089;
  assign n2110 = n2108 & n2109;
  assign n2111 = ~n2094 & ~n2100;
  assign n2112 = ~n2107 & n2111;
  assign po39 = ~n2110 | ~n2112;
  assign n2114 = pi075 & ~n253;
  assign n2115 = pi083 & ~n273;
  assign n2116 = n253 & n2115;
  assign n2117 = pi086 & n273;
  assign n2118 = n253 & n2117;
  assign n2119 = ~n283 & n2118;
  assign n2120 = pi044 & n283;
  assign n2121 = n253 & n2120;
  assign n2122 = n273 & n2121;
  assign n2123 = ~n262 & n2122;
  assign n2124 = ~n2114 & ~n2116;
  assign n2125 = ~n2119 & n2124;
  assign n2126 = ~n286 & ~n2123;
  assign n2127 = n2125 & n2126;
  assign n2128 = n1718 & ~n2127;
  assign n2129 = n1737 & ~n2127;
  assign n2130 = ~n1718 & n2129;
  assign n2131 = ~n1737 & ~n2127;
  assign n2132 = ~n1718 & n2131;
  assign n2133 = n1742 & n2132;
  assign n2134 = ~n1742 & ~n2127;
  assign n2135 = ~n1718 & n2134;
  assign n2136 = ~n1737 & n2135;
  assign n2137 = n1748 & n2136;
  assign n2138 = ~n1748 & ~n2127;
  assign n2139 = ~n1737 & n2138;
  assign n2140 = ~n1718 & n2139;
  assign n2141 = ~n1742 & n2140;
  assign n2142 = n1753 & n2141;
  assign n2143 = ~n1753 & ~n2127;
  assign n2144 = ~n1742 & n2143;
  assign n2145 = ~n1718 & n2144;
  assign n2146 = ~n1737 & n2145;
  assign n2147 = ~n1748 & n2146;
  assign n2148 = pi005 & n2147;
  assign n2149 = n1368 & ~n1748;
  assign n2150 = ~n1737 & n2149;
  assign n2151 = ~n1718 & n2150;
  assign n2152 = ~n1742 & n2151;
  assign n2153 = ~n1753 & n2152;
  assign n2154 = pi095 & n2153;
  assign n2155 = ~pi005 & n2154;
  assign n2156 = ~n2128 & ~n2130;
  assign n2157 = ~n2133 & ~n2137;
  assign n2158 = n2156 & n2157;
  assign n2159 = ~n2142 & ~n2148;
  assign n2160 = ~n2155 & n2159;
  assign po40 = ~n2158 | ~n2160;
  assign n2162 = pi076 & ~n253;
  assign n2163 = pi084 & ~n273;
  assign n2164 = n253 & n2163;
  assign n2165 = pi045 & n283;
  assign n2166 = n253 & n2165;
  assign n2167 = n273 & n2166;
  assign n2168 = ~n262 & n2167;
  assign n2169 = ~n2162 & ~n2164;
  assign n2170 = ~n568 & n2169;
  assign n2171 = ~n286 & ~n2168;
  assign n2172 = n2170 & n2171;
  assign n2173 = n1718 & ~n2172;
  assign n2174 = n1737 & ~n2172;
  assign n2175 = ~n1718 & n2174;
  assign n2176 = ~n1737 & ~n2172;
  assign n2177 = ~n1718 & n2176;
  assign n2178 = n1742 & n2177;
  assign n2179 = ~n1742 & ~n2172;
  assign n2180 = ~n1718 & n2179;
  assign n2181 = ~n1737 & n2180;
  assign n2182 = n1748 & n2181;
  assign n2183 = ~n1748 & ~n2172;
  assign n2184 = ~n1737 & n2183;
  assign n2185 = ~n1718 & n2184;
  assign n2186 = ~n1742 & n2185;
  assign n2187 = n1753 & n2186;
  assign n2188 = ~n1753 & ~n2172;
  assign n2189 = ~n1742 & n2188;
  assign n2190 = ~n1718 & n2189;
  assign n2191 = ~n1737 & n2190;
  assign n2192 = ~n1748 & n2191;
  assign n2193 = pi005 & n2192;
  assign n2194 = n1422 & ~n1748;
  assign n2195 = ~n1737 & n2194;
  assign n2196 = ~n1718 & n2195;
  assign n2197 = ~n1742 & n2196;
  assign n2198 = ~n1753 & n2197;
  assign n2199 = pi095 & n2198;
  assign n2200 = ~pi005 & n2199;
  assign n2201 = ~n2173 & ~n2175;
  assign n2202 = ~n2178 & ~n2182;
  assign n2203 = n2201 & n2202;
  assign n2204 = ~n2187 & ~n2193;
  assign n2205 = ~n2200 & n2204;
  assign po41 = ~n2203 | ~n2205;
  assign n2207 = pi077 & ~n253;
  assign n2208 = pi085 & ~n273;
  assign n2209 = n253 & n2208;
  assign n2210 = pi046 & n283;
  assign n2211 = n253 & n2210;
  assign n2212 = n273 & n2211;
  assign n2213 = ~n262 & n2212;
  assign n2214 = ~n2207 & ~n2209;
  assign n2215 = ~n596 & n2214;
  assign n2216 = ~n286 & ~n2213;
  assign n2217 = n2215 & n2216;
  assign n2218 = n1718 & ~n2217;
  assign n2219 = n1737 & ~n2217;
  assign n2220 = ~n1718 & n2219;
  assign n2221 = ~n1737 & ~n2217;
  assign n2222 = ~n1718 & n2221;
  assign n2223 = n1742 & n2222;
  assign n2224 = ~n1742 & ~n2217;
  assign n2225 = ~n1718 & n2224;
  assign n2226 = ~n1737 & n2225;
  assign n2227 = n1748 & n2226;
  assign n2228 = ~n1748 & ~n2217;
  assign n2229 = ~n1737 & n2228;
  assign n2230 = ~n1718 & n2229;
  assign n2231 = ~n1742 & n2230;
  assign n2232 = n1753 & n2231;
  assign n2233 = ~n1753 & ~n2217;
  assign n2234 = ~n1742 & n2233;
  assign n2235 = ~n1718 & n2234;
  assign n2236 = ~n1737 & n2235;
  assign n2237 = ~n1748 & n2236;
  assign n2238 = pi005 & n2237;
  assign n2239 = n1476 & ~n1748;
  assign n2240 = ~n1737 & n2239;
  assign n2241 = ~n1718 & n2240;
  assign n2242 = ~n1742 & n2241;
  assign n2243 = ~n1753 & n2242;
  assign n2244 = pi095 & n2243;
  assign n2245 = ~pi005 & n2244;
  assign n2246 = ~n2218 & ~n2220;
  assign n2247 = ~n2223 & ~n2227;
  assign n2248 = n2246 & n2247;
  assign n2249 = ~n2232 & ~n2238;
  assign n2250 = ~n2245 & n2249;
  assign po42 = ~n2248 | ~n2250;
  assign n2252 = pi078 & ~n253;
  assign n2253 = pi086 & ~n273;
  assign n2254 = n253 & n2253;
  assign n2255 = pi047 & n283;
  assign n2256 = n253 & n2255;
  assign n2257 = n273 & n2256;
  assign n2258 = ~n262 & n2257;
  assign n2259 = ~n2252 & ~n2254;
  assign n2260 = ~n540 & n2259;
  assign n2261 = ~n286 & ~n2258;
  assign n2262 = n2260 & n2261;
  assign n2263 = n1718 & ~n2262;
  assign n2264 = n1737 & ~n2262;
  assign n2265 = ~n1718 & n2264;
  assign n2266 = ~n1737 & ~n2262;
  assign n2267 = ~n1718 & n2266;
  assign n2268 = n1742 & n2267;
  assign n2269 = ~n1742 & ~n2262;
  assign n2270 = ~n1718 & n2269;
  assign n2271 = ~n1737 & n2270;
  assign n2272 = n1748 & n2271;
  assign n2273 = ~n1748 & ~n2262;
  assign n2274 = ~n1737 & n2273;
  assign n2275 = ~n1718 & n2274;
  assign n2276 = ~n1742 & n2275;
  assign n2277 = n1753 & n2276;
  assign n2278 = ~n1753 & ~n2262;
  assign n2279 = ~n1742 & n2278;
  assign n2280 = ~n1718 & n2279;
  assign n2281 = ~n1737 & n2280;
  assign n2282 = ~n1748 & n2281;
  assign n2283 = pi005 & n2282;
  assign n2284 = n1530 & ~n1748;
  assign n2285 = ~n1737 & n2284;
  assign n2286 = ~n1718 & n2285;
  assign n2287 = ~n1742 & n2286;
  assign n2288 = ~n1753 & n2287;
  assign n2289 = pi095 & n2288;
  assign n2290 = ~pi005 & n2289;
  assign n2291 = ~n2263 & ~n2265;
  assign n2292 = ~n2268 & ~n2272;
  assign n2293 = n2291 & n2292;
  assign n2294 = ~n2277 & ~n2283;
  assign n2295 = ~n2290 & n2294;
  assign po43 = ~n2293 | ~n2295;
  assign n2297 = pi079 & ~n253;
  assign n2298 = pi041 & ~n273;
  assign n2299 = n253 & n2298;
  assign n2300 = pi048 & n283;
  assign n2301 = n253 & n2300;
  assign n2302 = n273 & n2301;
  assign n2303 = ~n262 & n2302;
  assign n2304 = ~n2297 & ~n2299;
  assign n2305 = ~n385 & n2304;
  assign n2306 = ~n286 & ~n2303;
  assign n2307 = n2305 & n2306;
  assign n2308 = n1718 & ~n2307;
  assign n2309 = n1737 & ~n2307;
  assign n2310 = ~n1718 & n2309;
  assign n2311 = ~n1737 & ~n2307;
  assign n2312 = ~n1718 & n2311;
  assign n2313 = n1742 & n2312;
  assign n2314 = ~n1742 & ~n2307;
  assign n2315 = ~n1718 & n2314;
  assign n2316 = ~n1737 & n2315;
  assign n2317 = n1748 & n2316;
  assign n2318 = ~n1748 & ~n2307;
  assign n2319 = ~n1737 & n2318;
  assign n2320 = ~n1718 & n2319;
  assign n2321 = ~n1742 & n2320;
  assign n2322 = n1753 & n2321;
  assign n2323 = ~n1753 & ~n2307;
  assign n2324 = ~n1742 & n2323;
  assign n2325 = ~n1718 & n2324;
  assign n2326 = ~n1737 & n2325;
  assign n2327 = ~n1748 & n2326;
  assign n2328 = pi005 & n2327;
  assign n2329 = n1584 & ~n1748;
  assign n2330 = ~n1737 & n2329;
  assign n2331 = ~n1718 & n2330;
  assign n2332 = ~n1742 & n2331;
  assign n2333 = ~n1753 & n2332;
  assign n2334 = pi095 & n2333;
  assign n2335 = ~pi005 & n2334;
  assign n2336 = ~n2308 & ~n2310;
  assign n2337 = ~n2313 & ~n2317;
  assign n2338 = n2336 & n2337;
  assign n2339 = ~n2322 & ~n2328;
  assign n2340 = ~n2335 & n2339;
  assign po44 = ~n2338 | ~n2340;
  assign n2342 = pi080 & ~n253;
  assign n2343 = pi042 & ~n273;
  assign n2344 = n253 & n2343;
  assign n2345 = pi049 & n283;
  assign n2346 = n253 & n2345;
  assign n2347 = n273 & n2346;
  assign n2348 = ~n262 & n2347;
  assign n2349 = ~n2342 & ~n2344;
  assign n2350 = ~n412 & n2349;
  assign n2351 = ~n286 & ~n2348;
  assign n2352 = n2350 & n2351;
  assign n2353 = n1718 & ~n2352;
  assign n2354 = n1737 & ~n2352;
  assign n2355 = ~n1718 & n2354;
  assign n2356 = ~n1737 & ~n2352;
  assign n2357 = ~n1718 & n2356;
  assign n2358 = n1742 & n2357;
  assign n2359 = ~n1742 & ~n2352;
  assign n2360 = ~n1718 & n2359;
  assign n2361 = ~n1737 & n2360;
  assign n2362 = n1748 & n2361;
  assign n2363 = ~n1748 & ~n2352;
  assign n2364 = ~n1737 & n2363;
  assign n2365 = ~n1718 & n2364;
  assign n2366 = ~n1742 & n2365;
  assign n2367 = n1753 & n2366;
  assign n2368 = ~n1753 & ~n2352;
  assign n2369 = ~n1742 & n2368;
  assign n2370 = ~n1718 & n2369;
  assign n2371 = ~n1737 & n2370;
  assign n2372 = ~n1748 & n2371;
  assign n2373 = pi005 & n2372;
  assign n2374 = n1638 & ~n1748;
  assign n2375 = ~n1737 & n2374;
  assign n2376 = ~n1718 & n2375;
  assign n2377 = ~n1742 & n2376;
  assign n2378 = ~n1753 & n2377;
  assign n2379 = pi095 & n2378;
  assign n2380 = ~pi005 & n2379;
  assign n2381 = ~n2353 & ~n2355;
  assign n2382 = ~n2358 & ~n2362;
  assign n2383 = n2381 & n2382;
  assign n2384 = ~n2367 & ~n2373;
  assign n2385 = ~n2380 & n2384;
  assign po45 = ~n2383 | ~n2385;
  assign n2387 = pi081 & ~n253;
  assign n2388 = pi043 & ~n273;
  assign n2389 = n253 & n2388;
  assign n2390 = pi050 & n283;
  assign n2391 = n253 & n2390;
  assign n2392 = n273 & n2391;
  assign n2393 = ~n262 & n2392;
  assign n2394 = ~n2387 & ~n2389;
  assign n2395 = ~n437 & n2394;
  assign n2396 = ~n286 & ~n2393;
  assign n2397 = n2395 & n2396;
  assign n2398 = n1718 & ~n2397;
  assign n2399 = n1737 & ~n2397;
  assign n2400 = ~n1718 & n2399;
  assign n2401 = ~n1737 & ~n2397;
  assign n2402 = ~n1718 & n2401;
  assign n2403 = n1742 & n2402;
  assign n2404 = ~n1742 & ~n2397;
  assign n2405 = ~n1718 & n2404;
  assign n2406 = ~n1737 & n2405;
  assign n2407 = n1748 & n2406;
  assign n2408 = ~n1748 & ~n2397;
  assign n2409 = ~n1737 & n2408;
  assign n2410 = ~n1718 & n2409;
  assign n2411 = ~n1742 & n2410;
  assign n2412 = n1753 & n2411;
  assign n2413 = ~n1753 & ~n2397;
  assign n2414 = ~n1742 & n2413;
  assign n2415 = ~n1718 & n2414;
  assign n2416 = ~n1737 & n2415;
  assign n2417 = ~n1748 & n2416;
  assign n2418 = pi005 & n2417;
  assign n2419 = n1692 & ~n1748;
  assign n2420 = ~n1737 & n2419;
  assign n2421 = ~n1718 & n2420;
  assign n2422 = ~n1742 & n2421;
  assign n2423 = ~n1753 & n2422;
  assign n2424 = pi095 & n2423;
  assign n2425 = ~pi005 & n2424;
  assign n2426 = ~n2398 & ~n2400;
  assign n2427 = ~n2403 & ~n2407;
  assign n2428 = n2426 & n2427;
  assign n2429 = ~n2412 & ~n2418;
  assign n2430 = ~n2425 & n2429;
  assign po46 = ~n2428 | ~n2430;
  assign n2432 = pi082 & ~n253;
  assign n2433 = pi044 & ~n273;
  assign n2434 = n253 & n2433;
  assign n2435 = pi051 & n283;
  assign n2436 = n253 & n2435;
  assign n2437 = n273 & n2436;
  assign n2438 = ~n262 & n2437;
  assign n2439 = ~n2432 & ~n2434;
  assign n2440 = ~n462 & n2439;
  assign n2441 = ~n286 & ~n2438;
  assign n2442 = n2440 & n2441;
  assign n2443 = n1718 & ~n2442;
  assign n2444 = n1737 & ~n2442;
  assign n2445 = ~n1718 & n2444;
  assign n2446 = ~n1737 & ~n2442;
  assign n2447 = ~n1718 & n2446;
  assign n2448 = n1742 & n2447;
  assign n2449 = ~n1742 & ~n2442;
  assign n2450 = ~n1718 & n2449;
  assign n2451 = ~n1737 & n2450;
  assign n2452 = n1748 & n2451;
  assign n2453 = ~n1748 & ~n2442;
  assign n2454 = ~n1737 & n2453;
  assign n2455 = ~n1718 & n2454;
  assign n2456 = ~n1742 & n2455;
  assign n2457 = n1753 & n2456;
  assign n2458 = ~n1753 & ~n2442;
  assign n2459 = ~n1742 & n2458;
  assign n2460 = ~n1718 & n2459;
  assign n2461 = ~n1737 & n2460;
  assign n2462 = ~n1748 & n2461;
  assign n2463 = pi005 & n2462;
  assign n2464 = n879 & ~n1748;
  assign n2465 = ~n1737 & n2464;
  assign n2466 = ~n1718 & n2465;
  assign n2467 = ~n1742 & n2466;
  assign n2468 = ~n1753 & n2467;
  assign n2469 = pi095 & n2468;
  assign n2470 = ~pi005 & n2469;
  assign n2471 = ~n2443 & ~n2445;
  assign n2472 = ~n2448 & ~n2452;
  assign n2473 = n2471 & n2472;
  assign n2474 = ~n2457 & ~n2463;
  assign n2475 = ~n2470 & n2474;
  assign po47 = ~n2473 | ~n2475;
  assign n2477 = pi083 & ~n253;
  assign n2478 = pi045 & ~n273;
  assign n2479 = n253 & n2478;
  assign n2480 = pi087 & n283;
  assign n2481 = n253 & n2480;
  assign n2482 = n273 & n2481;
  assign n2483 = ~n262 & n2482;
  assign n2484 = ~n2477 & ~n2479;
  assign n2485 = ~n487 & n2484;
  assign n2486 = ~n286 & ~n2483;
  assign n2487 = n2485 & n2486;
  assign n2488 = n1718 & ~n2487;
  assign n2489 = n1737 & ~n2487;
  assign n2490 = ~n1718 & n2489;
  assign n2491 = ~n1737 & ~n2487;
  assign n2492 = ~n1718 & n2491;
  assign n2493 = n1742 & n2492;
  assign n2494 = ~n1742 & ~n2487;
  assign n2495 = ~n1718 & n2494;
  assign n2496 = ~n1737 & n2495;
  assign n2497 = n1748 & n2496;
  assign n2498 = ~n1748 & ~n2487;
  assign n2499 = ~n1737 & n2498;
  assign n2500 = ~n1718 & n2499;
  assign n2501 = ~n1742 & n2500;
  assign n2502 = n1753 & n2501;
  assign n2503 = ~n1753 & ~n2487;
  assign n2504 = ~n1742 & n2503;
  assign n2505 = ~n1718 & n2504;
  assign n2506 = ~n1737 & n2505;
  assign n2507 = ~n1748 & n2506;
  assign n2508 = pi005 & n2507;
  assign n2509 = n709 & ~n1748;
  assign n2510 = ~n1737 & n2509;
  assign n2511 = ~n1718 & n2510;
  assign n2512 = ~n1742 & n2511;
  assign n2513 = ~n1753 & n2512;
  assign n2514 = pi095 & n2513;
  assign n2515 = ~pi005 & n2514;
  assign n2516 = ~n2488 & ~n2490;
  assign n2517 = ~n2493 & ~n2497;
  assign n2518 = n2516 & n2517;
  assign n2519 = ~n2502 & ~n2508;
  assign n2520 = ~n2515 & n2519;
  assign po48 = ~n2518 | ~n2520;
  assign n2522 = pi084 & ~n253;
  assign n2523 = pi046 & ~n273;
  assign n2524 = n253 & n2523;
  assign n2525 = pi009 & n283;
  assign n2526 = n253 & n2525;
  assign n2527 = n273 & n2526;
  assign n2528 = ~n262 & n2527;
  assign n2529 = ~n2522 & ~n2524;
  assign n2530 = ~n512 & n2529;
  assign n2531 = ~n286 & ~n2528;
  assign n2532 = n2530 & n2531;
  assign n2533 = n1718 & ~n2532;
  assign n2534 = n1737 & ~n2532;
  assign n2535 = ~n1718 & n2534;
  assign n2536 = ~n1737 & ~n2532;
  assign n2537 = ~n1718 & n2536;
  assign n2538 = n1742 & n2537;
  assign n2539 = ~n1742 & ~n2532;
  assign n2540 = ~n1718 & n2539;
  assign n2541 = ~n1737 & n2540;
  assign n2542 = n1748 & n2541;
  assign n2543 = ~n1748 & ~n2532;
  assign n2544 = ~n1737 & n2543;
  assign n2545 = ~n1718 & n2544;
  assign n2546 = ~n1742 & n2545;
  assign n2547 = n1753 & n2546;
  assign n2548 = ~n1753 & ~n2532;
  assign n2549 = ~n1742 & n2548;
  assign n2550 = ~n1718 & n2549;
  assign n2551 = ~n1737 & n2550;
  assign n2552 = ~n1748 & n2551;
  assign n2553 = pi005 & n2552;
  assign n2554 = n763 & ~n1748;
  assign n2555 = ~n1737 & n2554;
  assign n2556 = ~n1718 & n2555;
  assign n2557 = ~n1742 & n2556;
  assign n2558 = ~n1753 & n2557;
  assign n2559 = pi095 & n2558;
  assign n2560 = ~pi005 & n2559;
  assign n2561 = ~n2533 & ~n2535;
  assign n2562 = ~n2538 & ~n2542;
  assign n2563 = n2561 & n2562;
  assign n2564 = ~n2547 & ~n2553;
  assign n2565 = ~n2560 & n2564;
  assign po49 = ~n2563 | ~n2565;
  assign n2567 = pi085 & ~n253;
  assign n2568 = pi047 & ~n273;
  assign n2569 = n253 & n2568;
  assign n2570 = pi010 & n283;
  assign n2571 = n253 & n2570;
  assign n2572 = n273 & n2571;
  assign n2573 = ~n262 & n2572;
  assign n2574 = ~n2567 & ~n2569;
  assign n2575 = ~n289 & n2574;
  assign n2576 = ~n286 & ~n2573;
  assign n2577 = n2575 & n2576;
  assign n2578 = n1718 & ~n2577;
  assign n2579 = n1737 & ~n2577;
  assign n2580 = ~n1718 & n2579;
  assign n2581 = ~n1737 & ~n2577;
  assign n2582 = ~n1718 & n2581;
  assign n2583 = n1742 & n2582;
  assign n2584 = ~n1742 & ~n2577;
  assign n2585 = ~n1718 & n2584;
  assign n2586 = ~n1737 & n2585;
  assign n2587 = n1748 & n2586;
  assign n2588 = ~n1748 & ~n2577;
  assign n2589 = ~n1737 & n2588;
  assign n2590 = ~n1718 & n2589;
  assign n2591 = ~n1742 & n2590;
  assign n2592 = n1753 & n2591;
  assign n2593 = ~n1753 & ~n2577;
  assign n2594 = ~n1742 & n2593;
  assign n2595 = ~n1718 & n2594;
  assign n2596 = ~n1737 & n2595;
  assign n2597 = ~n1748 & n2596;
  assign n2598 = pi005 & n2597;
  assign n2599 = n817 & ~n1748;
  assign n2600 = ~n1737 & n2599;
  assign n2601 = ~n1718 & n2600;
  assign n2602 = ~n1742 & n2601;
  assign n2603 = ~n1753 & n2602;
  assign n2604 = pi095 & n2603;
  assign n2605 = ~pi005 & n2604;
  assign n2606 = ~n2578 & ~n2580;
  assign n2607 = ~n2583 & ~n2587;
  assign n2608 = n2606 & n2607;
  assign n2609 = ~n2592 & ~n2598;
  assign n2610 = ~n2605 & n2609;
  assign po50 = ~n2608 | ~n2610;
  assign n2612 = pi086 & ~n253;
  assign n2613 = pi048 & ~n273;
  assign n2614 = n253 & n2613;
  assign n2615 = pi011 & n283;
  assign n2616 = n253 & n2615;
  assign n2617 = n273 & n2616;
  assign n2618 = ~n262 & n2617;
  assign n2619 = ~n2612 & ~n2614;
  assign n2620 = ~n335 & n2619;
  assign n2621 = ~n286 & ~n2618;
  assign n2622 = n2620 & n2621;
  assign n2623 = n1718 & ~n2622;
  assign n2624 = n1737 & ~n2622;
  assign n2625 = ~n1718 & n2624;
  assign n2626 = ~n1737 & ~n2622;
  assign n2627 = ~n1718 & n2626;
  assign n2628 = n1742 & n2627;
  assign n2629 = ~n1742 & ~n2622;
  assign n2630 = ~n1718 & n2629;
  assign n2631 = ~n1737 & n2630;
  assign n2632 = n1748 & n2631;
  assign n2633 = ~n1748 & ~n2622;
  assign n2634 = ~n1737 & n2633;
  assign n2635 = ~n1718 & n2634;
  assign n2636 = ~n1742 & n2635;
  assign n2637 = n1753 & n2636;
  assign n2638 = ~n1753 & ~n2622;
  assign n2639 = ~n1742 & n2638;
  assign n2640 = ~n1718 & n2639;
  assign n2641 = ~n1737 & n2640;
  assign n2642 = ~n1748 & n2641;
  assign n2643 = pi005 & n2642;
  assign n2644 = n653 & ~n1748;
  assign n2645 = ~n1737 & n2644;
  assign n2646 = ~n1718 & n2645;
  assign n2647 = ~n1742 & n2646;
  assign n2648 = ~n1753 & n2647;
  assign n2649 = pi095 & n2648;
  assign n2650 = ~pi005 & n2649;
  assign n2651 = ~n2623 & ~n2625;
  assign n2652 = ~n2628 & ~n2632;
  assign n2653 = n2651 & n2652;
  assign n2654 = ~n2637 & ~n2643;
  assign n2655 = ~n2650 & n2654;
  assign po51 = ~n2653 | ~n2655;
  assign n2657 = pi041 & ~n253;
  assign n2658 = pi049 & ~n273;
  assign n2659 = n253 & n2658;
  assign n2660 = pi087 & n273;
  assign n2661 = n253 & n2660;
  assign n2662 = ~n283 & n2661;
  assign n2663 = pi012 & n283;
  assign n2664 = n253 & n2663;
  assign n2665 = n273 & n2664;
  assign n2666 = ~n262 & n2665;
  assign n2667 = ~n2657 & ~n2659;
  assign n2668 = ~n2662 & n2667;
  assign n2669 = ~n286 & ~n2666;
  assign n2670 = n2668 & n2669;
  assign n2671 = n1718 & ~n2670;
  assign n2672 = n1737 & ~n2670;
  assign n2673 = ~n1718 & n2672;
  assign n2674 = ~n1737 & ~n2670;
  assign n2675 = ~n1718 & n2674;
  assign n2676 = n1742 & n2675;
  assign n2677 = ~n1742 & ~n2670;
  assign n2678 = ~n1718 & n2677;
  assign n2679 = ~n1737 & n2678;
  assign n2680 = n1748 & n2679;
  assign n2681 = ~n1748 & ~n2670;
  assign n2682 = ~n1737 & n2681;
  assign n2683 = ~n1718 & n2682;
  assign n2684 = ~n1742 & n2683;
  assign n2685 = n1753 & n2684;
  assign n2686 = ~n1753 & ~n2670;
  assign n2687 = ~n1742 & n2686;
  assign n2688 = ~n1718 & n2687;
  assign n2689 = ~n1737 & n2688;
  assign n2690 = ~n1748 & n2689;
  assign n2691 = pi005 & n2690;
  assign n2692 = n583 & ~n1748;
  assign n2693 = ~n1737 & n2692;
  assign n2694 = ~n1718 & n2693;
  assign n2695 = ~n1742 & n2694;
  assign n2696 = ~n1753 & n2695;
  assign n2697 = pi095 & n2696;
  assign n2698 = ~pi005 & n2697;
  assign n2699 = ~n2671 & ~n2673;
  assign n2700 = ~n2676 & ~n2680;
  assign n2701 = n2699 & n2700;
  assign n2702 = ~n2685 & ~n2691;
  assign n2703 = ~n2698 & n2702;
  assign po52 = ~n2701 | ~n2703;
  assign n2705 = pi042 & ~n253;
  assign n2706 = pi050 & ~n273;
  assign n2707 = n253 & n2706;
  assign n2708 = pi009 & n273;
  assign n2709 = n253 & n2708;
  assign n2710 = ~n283 & n2709;
  assign n2711 = pi013 & n283;
  assign n2712 = n253 & n2711;
  assign n2713 = n273 & n2712;
  assign n2714 = ~n262 & n2713;
  assign n2715 = ~n2705 & ~n2707;
  assign n2716 = ~n2710 & n2715;
  assign n2717 = ~n286 & ~n2714;
  assign n2718 = n2716 & n2717;
  assign n2719 = n1718 & ~n2718;
  assign n2720 = n1737 & ~n2718;
  assign n2721 = ~n1718 & n2720;
  assign n2722 = ~n1737 & ~n2718;
  assign n2723 = ~n1718 & n2722;
  assign n2724 = n1742 & n2723;
  assign n2725 = ~n1742 & ~n2718;
  assign n2726 = ~n1718 & n2725;
  assign n2727 = ~n1737 & n2726;
  assign n2728 = n1748 & n2727;
  assign n2729 = ~n1748 & ~n2718;
  assign n2730 = ~n1737 & n2729;
  assign n2731 = ~n1718 & n2730;
  assign n2732 = ~n1742 & n2731;
  assign n2733 = n1753 & n2732;
  assign n2734 = ~n1753 & ~n2718;
  assign n2735 = ~n1742 & n2734;
  assign n2736 = ~n1718 & n2735;
  assign n2737 = ~n1737 & n2736;
  assign n2738 = ~n1748 & n2737;
  assign n2739 = pi005 & n2738;
  assign n2740 = n611 & ~n1748;
  assign n2741 = ~n1737 & n2740;
  assign n2742 = ~n1718 & n2741;
  assign n2743 = ~n1742 & n2742;
  assign n2744 = ~n1753 & n2743;
  assign n2745 = pi095 & n2744;
  assign n2746 = ~pi005 & n2745;
  assign n2747 = ~n2719 & ~n2721;
  assign n2748 = ~n2724 & ~n2728;
  assign n2749 = n2747 & n2748;
  assign n2750 = ~n2733 & ~n2739;
  assign n2751 = ~n2746 & n2750;
  assign po53 = ~n2749 | ~n2751;
  assign n2753 = pi043 & ~n253;
  assign n2754 = pi051 & ~n273;
  assign n2755 = n253 & n2754;
  assign n2756 = pi010 & n273;
  assign n2757 = n253 & n2756;
  assign n2758 = ~n283 & n2757;
  assign n2759 = pi014 & n283;
  assign n2760 = n253 & n2759;
  assign n2761 = n273 & n2760;
  assign n2762 = ~n262 & n2761;
  assign n2763 = ~n2753 & ~n2755;
  assign n2764 = ~n2758 & n2763;
  assign n2765 = ~n286 & ~n2762;
  assign n2766 = n2764 & n2765;
  assign n2767 = n1718 & ~n2766;
  assign n2768 = n1737 & ~n2766;
  assign n2769 = ~n1718 & n2768;
  assign n2770 = ~n1737 & ~n2766;
  assign n2771 = ~n1718 & n2770;
  assign n2772 = n1742 & n2771;
  assign n2773 = ~n1742 & ~n2766;
  assign n2774 = ~n1718 & n2773;
  assign n2775 = ~n1737 & n2774;
  assign n2776 = n1748 & n2775;
  assign n2777 = ~n1748 & ~n2766;
  assign n2778 = ~n1737 & n2777;
  assign n2779 = ~n1718 & n2778;
  assign n2780 = ~n1742 & n2779;
  assign n2781 = n1753 & n2780;
  assign n2782 = ~n1753 & ~n2766;
  assign n2783 = ~n1742 & n2782;
  assign n2784 = ~n1718 & n2783;
  assign n2785 = ~n1737 & n2784;
  assign n2786 = ~n1748 & n2785;
  assign n2787 = pi005 & n2786;
  assign n2788 = n555 & ~n1748;
  assign n2789 = ~n1737 & n2788;
  assign n2790 = ~n1718 & n2789;
  assign n2791 = ~n1742 & n2790;
  assign n2792 = ~n1753 & n2791;
  assign n2793 = pi095 & n2792;
  assign n2794 = ~pi005 & n2793;
  assign n2795 = ~n2767 & ~n2769;
  assign n2796 = ~n2772 & ~n2776;
  assign n2797 = n2795 & n2796;
  assign n2798 = ~n2781 & ~n2787;
  assign n2799 = ~n2794 & n2798;
  assign po54 = ~n2797 | ~n2799;
  assign n2801 = pi044 & ~n253;
  assign n2802 = pi087 & ~n273;
  assign n2803 = n253 & n2802;
  assign n2804 = pi011 & n273;
  assign n2805 = n253 & n2804;
  assign n2806 = ~n283 & n2805;
  assign n2807 = pi015 & n283;
  assign n2808 = n253 & n2807;
  assign n2809 = n273 & n2808;
  assign n2810 = ~n262 & n2809;
  assign n2811 = ~n2801 & ~n2803;
  assign n2812 = ~n2806 & n2811;
  assign n2813 = ~n286 & ~n2810;
  assign n2814 = n2812 & n2813;
  assign n2815 = n1718 & ~n2814;
  assign n2816 = n1737 & ~n2814;
  assign n2817 = ~n1718 & n2816;
  assign n2818 = ~n1737 & ~n2814;
  assign n2819 = ~n1718 & n2818;
  assign n2820 = n1742 & n2819;
  assign n2821 = ~n1742 & ~n2814;
  assign n2822 = ~n1718 & n2821;
  assign n2823 = ~n1737 & n2822;
  assign n2824 = n1748 & n2823;
  assign n2825 = ~n1748 & ~n2814;
  assign n2826 = ~n1737 & n2825;
  assign n2827 = ~n1718 & n2826;
  assign n2828 = ~n1742 & n2827;
  assign n2829 = n1753 & n2828;
  assign n2830 = ~n1753 & ~n2814;
  assign n2831 = ~n1742 & n2830;
  assign n2832 = ~n1718 & n2831;
  assign n2833 = ~n1737 & n2832;
  assign n2834 = ~n1748 & n2833;
  assign n2835 = pi005 & n2834;
  assign n2836 = n401 & ~n1748;
  assign n2837 = ~n1737 & n2836;
  assign n2838 = ~n1718 & n2837;
  assign n2839 = ~n1742 & n2838;
  assign n2840 = ~n1753 & n2839;
  assign n2841 = pi095 & n2840;
  assign n2842 = ~pi005 & n2841;
  assign n2843 = ~n2815 & ~n2817;
  assign n2844 = ~n2820 & ~n2824;
  assign n2845 = n2843 & n2844;
  assign n2846 = ~n2829 & ~n2835;
  assign n2847 = ~n2842 & n2846;
  assign po55 = ~n2845 | ~n2847;
  assign n2849 = pi045 & ~n253;
  assign n2850 = pi009 & ~n273;
  assign n2851 = n253 & n2850;
  assign n2852 = pi012 & n273;
  assign n2853 = n253 & n2852;
  assign n2854 = ~n283 & n2853;
  assign n2855 = pi016 & n283;
  assign n2856 = n253 & n2855;
  assign n2857 = n273 & n2856;
  assign n2858 = ~n262 & n2857;
  assign n2859 = ~n2849 & ~n2851;
  assign n2860 = ~n2854 & n2859;
  assign n2861 = ~n286 & ~n2858;
  assign n2862 = n2860 & n2861;
  assign n2863 = n1718 & ~n2862;
  assign n2864 = n1737 & ~n2862;
  assign n2865 = ~n1718 & n2864;
  assign n2866 = ~n1737 & ~n2862;
  assign n2867 = ~n1718 & n2866;
  assign n2868 = n1742 & n2867;
  assign n2869 = ~n1742 & ~n2862;
  assign n2870 = ~n1718 & n2869;
  assign n2871 = ~n1737 & n2870;
  assign n2872 = n1748 & n2871;
  assign n2873 = ~n1748 & ~n2862;
  assign n2874 = ~n1737 & n2873;
  assign n2875 = ~n1718 & n2874;
  assign n2876 = ~n1742 & n2875;
  assign n2877 = n1753 & n2876;
  assign n2878 = ~n1753 & ~n2862;
  assign n2879 = ~n1742 & n2878;
  assign n2880 = ~n1718 & n2879;
  assign n2881 = ~n1737 & n2880;
  assign n2882 = ~n1748 & n2881;
  assign n2883 = pi005 & n2882;
  assign n2884 = n426 & ~n1748;
  assign n2885 = ~n1737 & n2884;
  assign n2886 = ~n1718 & n2885;
  assign n2887 = ~n1742 & n2886;
  assign n2888 = ~n1753 & n2887;
  assign n2889 = pi095 & n2888;
  assign n2890 = ~pi005 & n2889;
  assign n2891 = ~n2863 & ~n2865;
  assign n2892 = ~n2868 & ~n2872;
  assign n2893 = n2891 & n2892;
  assign n2894 = ~n2877 & ~n2883;
  assign n2895 = ~n2890 & n2894;
  assign po56 = ~n2893 | ~n2895;
  assign n2897 = pi046 & ~n253;
  assign n2898 = pi010 & ~n273;
  assign n2899 = n253 & n2898;
  assign n2900 = pi013 & n273;
  assign n2901 = n253 & n2900;
  assign n2902 = ~n283 & n2901;
  assign n2903 = pi017 & n283;
  assign n2904 = n253 & n2903;
  assign n2905 = n273 & n2904;
  assign n2906 = ~n262 & n2905;
  assign n2907 = ~n2897 & ~n2899;
  assign n2908 = ~n2902 & n2907;
  assign n2909 = ~n286 & ~n2906;
  assign n2910 = n2908 & n2909;
  assign n2911 = n1718 & ~n2910;
  assign n2912 = n1737 & ~n2910;
  assign n2913 = ~n1718 & n2912;
  assign n2914 = ~n1737 & ~n2910;
  assign n2915 = ~n1718 & n2914;
  assign n2916 = n1742 & n2915;
  assign n2917 = ~n1742 & ~n2910;
  assign n2918 = ~n1718 & n2917;
  assign n2919 = ~n1737 & n2918;
  assign n2920 = n1748 & n2919;
  assign n2921 = ~n1748 & ~n2910;
  assign n2922 = ~n1737 & n2921;
  assign n2923 = ~n1718 & n2922;
  assign n2924 = ~n1742 & n2923;
  assign n2925 = n1753 & n2924;
  assign n2926 = ~n1753 & ~n2910;
  assign n2927 = ~n1742 & n2926;
  assign n2928 = ~n1718 & n2927;
  assign n2929 = ~n1737 & n2928;
  assign n2930 = ~n1748 & n2929;
  assign n2931 = pi005 & n2930;
  assign n2932 = n451 & ~n1748;
  assign n2933 = ~n1737 & n2932;
  assign n2934 = ~n1718 & n2933;
  assign n2935 = ~n1742 & n2934;
  assign n2936 = ~n1753 & n2935;
  assign n2937 = pi095 & n2936;
  assign n2938 = ~pi005 & n2937;
  assign n2939 = ~n2911 & ~n2913;
  assign n2940 = ~n2916 & ~n2920;
  assign n2941 = n2939 & n2940;
  assign n2942 = ~n2925 & ~n2931;
  assign n2943 = ~n2938 & n2942;
  assign po57 = ~n2941 | ~n2943;
  assign n2945 = pi047 & ~n253;
  assign n2946 = pi011 & ~n273;
  assign n2947 = n253 & n2946;
  assign n2948 = pi014 & n273;
  assign n2949 = n253 & n2948;
  assign n2950 = ~n283 & n2949;
  assign n2951 = pi018 & n283;
  assign n2952 = n253 & n2951;
  assign n2953 = n273 & n2952;
  assign n2954 = ~n262 & n2953;
  assign n2955 = ~n2945 & ~n2947;
  assign n2956 = ~n2950 & n2955;
  assign n2957 = ~n286 & ~n2954;
  assign n2958 = n2956 & n2957;
  assign n2959 = n1718 & ~n2958;
  assign n2960 = n1737 & ~n2958;
  assign n2961 = ~n1718 & n2960;
  assign n2962 = ~n1737 & ~n2958;
  assign n2963 = ~n1718 & n2962;
  assign n2964 = n1742 & n2963;
  assign n2965 = ~n1742 & ~n2958;
  assign n2966 = ~n1718 & n2965;
  assign n2967 = ~n1737 & n2966;
  assign n2968 = n1748 & n2967;
  assign n2969 = ~n1748 & ~n2958;
  assign n2970 = ~n1737 & n2969;
  assign n2971 = ~n1718 & n2970;
  assign n2972 = ~n1742 & n2971;
  assign n2973 = n1753 & n2972;
  assign n2974 = ~n1753 & ~n2958;
  assign n2975 = ~n1742 & n2974;
  assign n2976 = ~n1718 & n2975;
  assign n2977 = ~n1737 & n2976;
  assign n2978 = ~n1748 & n2977;
  assign n2979 = pi005 & n2978;
  assign n2980 = n476 & ~n1748;
  assign n2981 = ~n1737 & n2980;
  assign n2982 = ~n1718 & n2981;
  assign n2983 = ~n1742 & n2982;
  assign n2984 = ~n1753 & n2983;
  assign n2985 = pi095 & n2984;
  assign n2986 = ~pi005 & n2985;
  assign n2987 = ~n2959 & ~n2961;
  assign n2988 = ~n2964 & ~n2968;
  assign n2989 = n2987 & n2988;
  assign n2990 = ~n2973 & ~n2979;
  assign n2991 = ~n2986 & n2990;
  assign po58 = ~n2989 | ~n2991;
  assign n2993 = pi048 & ~n253;
  assign n2994 = pi012 & ~n273;
  assign n2995 = n253 & n2994;
  assign n2996 = pi015 & n273;
  assign n2997 = n253 & n2996;
  assign n2998 = ~n283 & n2997;
  assign n2999 = pi019 & n283;
  assign n3000 = n253 & n2999;
  assign n3001 = n273 & n3000;
  assign n3002 = ~n262 & n3001;
  assign n3003 = ~n2993 & ~n2995;
  assign n3004 = ~n2998 & n3003;
  assign n3005 = ~n286 & ~n3002;
  assign n3006 = n3004 & n3005;
  assign n3007 = n1718 & ~n3006;
  assign n3008 = n1737 & ~n3006;
  assign n3009 = ~n1718 & n3008;
  assign n3010 = ~n1737 & ~n3006;
  assign n3011 = ~n1718 & n3010;
  assign n3012 = n1742 & n3011;
  assign n3013 = ~n1742 & ~n3006;
  assign n3014 = ~n1718 & n3013;
  assign n3015 = ~n1737 & n3014;
  assign n3016 = n1748 & n3015;
  assign n3017 = ~n1748 & ~n3006;
  assign n3018 = ~n1737 & n3017;
  assign n3019 = ~n1718 & n3018;
  assign n3020 = ~n1742 & n3019;
  assign n3021 = n1753 & n3020;
  assign n3022 = ~n1753 & ~n3006;
  assign n3023 = ~n1742 & n3022;
  assign n3024 = ~n1718 & n3023;
  assign n3025 = ~n1737 & n3024;
  assign n3026 = ~n1748 & n3025;
  assign n3027 = pi005 & n3026;
  assign n3028 = n501 & ~n1748;
  assign n3029 = ~n1737 & n3028;
  assign n3030 = ~n1718 & n3029;
  assign n3031 = ~n1742 & n3030;
  assign n3032 = ~n1753 & n3031;
  assign n3033 = pi095 & n3032;
  assign n3034 = ~pi005 & n3033;
  assign n3035 = ~n3007 & ~n3009;
  assign n3036 = ~n3012 & ~n3016;
  assign n3037 = n3035 & n3036;
  assign n3038 = ~n3021 & ~n3027;
  assign n3039 = ~n3034 & n3038;
  assign po59 = ~n3037 | ~n3039;
  assign n3041 = pi049 & ~n253;
  assign n3042 = pi013 & ~n273;
  assign n3043 = n253 & n3042;
  assign n3044 = pi016 & n273;
  assign n3045 = n253 & n3044;
  assign n3046 = ~n283 & n3045;
  assign n3047 = pi020 & n283;
  assign n3048 = n253 & n3047;
  assign n3049 = n273 & n3048;
  assign n3050 = ~n262 & n3049;
  assign n3051 = ~n3041 & ~n3043;
  assign n3052 = ~n3046 & n3051;
  assign n3053 = ~n286 & ~n3050;
  assign n3054 = n3052 & n3053;
  assign n3055 = n1718 & ~n3054;
  assign n3056 = n1737 & ~n3054;
  assign n3057 = ~n1718 & n3056;
  assign n3058 = ~n1737 & ~n3054;
  assign n3059 = ~n1718 & n3058;
  assign n3060 = n1742 & n3059;
  assign n3061 = ~n1742 & ~n3054;
  assign n3062 = ~n1718 & n3061;
  assign n3063 = ~n1737 & n3062;
  assign n3064 = n1748 & n3063;
  assign n3065 = ~n1748 & ~n3054;
  assign n3066 = ~n1737 & n3065;
  assign n3067 = ~n1718 & n3066;
  assign n3068 = ~n1742 & n3067;
  assign n3069 = n1753 & n3068;
  assign n3070 = ~n1753 & ~n3054;
  assign n3071 = ~n1742 & n3070;
  assign n3072 = ~n1718 & n3071;
  assign n3073 = ~n1737 & n3072;
  assign n3074 = ~n1748 & n3073;
  assign n3075 = pi005 & n3074;
  assign n3076 = n526 & ~n1748;
  assign n3077 = ~n1737 & n3076;
  assign n3078 = ~n1718 & n3077;
  assign n3079 = ~n1742 & n3078;
  assign n3080 = ~n1753 & n3079;
  assign n3081 = pi095 & n3080;
  assign n3082 = ~pi005 & n3081;
  assign n3083 = ~n3055 & ~n3057;
  assign n3084 = ~n3060 & ~n3064;
  assign n3085 = n3083 & n3084;
  assign n3086 = ~n3069 & ~n3075;
  assign n3087 = ~n3082 & n3086;
  assign po60 = ~n3085 | ~n3087;
  assign n3089 = pi050 & ~n253;
  assign n3090 = pi014 & ~n273;
  assign n3091 = n253 & n3090;
  assign n3092 = pi017 & n273;
  assign n3093 = n253 & n3092;
  assign n3094 = ~n283 & n3093;
  assign n3095 = pi021 & n283;
  assign n3096 = n253 & n3095;
  assign n3097 = n273 & n3096;
  assign n3098 = ~n262 & n3097;
  assign n3099 = ~n3089 & ~n3091;
  assign n3100 = ~n3094 & n3099;
  assign n3101 = ~n286 & ~n3098;
  assign n3102 = n3100 & n3101;
  assign n3103 = n1718 & ~n3102;
  assign n3104 = n1737 & ~n3102;
  assign n3105 = ~n1718 & n3104;
  assign n3106 = ~n1737 & ~n3102;
  assign n3107 = ~n1718 & n3106;
  assign n3108 = n1742 & n3107;
  assign n3109 = ~n1742 & ~n3102;
  assign n3110 = ~n1718 & n3109;
  assign n3111 = ~n1737 & n3110;
  assign n3112 = n1748 & n3111;
  assign n3113 = ~n1748 & ~n3102;
  assign n3114 = ~n1737 & n3113;
  assign n3115 = ~n1718 & n3114;
  assign n3116 = ~n1742 & n3115;
  assign n3117 = n1753 & n3116;
  assign n3118 = ~n1753 & ~n3102;
  assign n3119 = ~n1742 & n3118;
  assign n3120 = ~n1718 & n3119;
  assign n3121 = ~n1737 & n3120;
  assign n3122 = ~n1748 & n3121;
  assign n3123 = pi005 & n3122;
  assign n3124 = ~pi005 & pi094;
  assign n3125 = ~n1748 & n3124;
  assign n3126 = ~n1737 & n3125;
  assign n3127 = ~n1718 & n3126;
  assign n3128 = ~n1742 & n3127;
  assign n3129 = ~n1753 & n3128;
  assign n3130 = pi095 & n3129;
  assign n3131 = ~pi005 & n3130;
  assign n3132 = ~n3103 & ~n3105;
  assign n3133 = ~n3108 & ~n3112;
  assign n3134 = n3132 & n3133;
  assign n3135 = ~n3117 & ~n3123;
  assign n3136 = ~n3131 & n3135;
  assign po61 = ~n3134 | ~n3136;
  assign n3138 = pi051 & ~n253;
  assign n3139 = pi015 & ~n273;
  assign n3140 = n253 & n3139;
  assign n3141 = pi018 & n273;
  assign n3142 = n253 & n3141;
  assign n3143 = ~n283 & n3142;
  assign n3144 = pi022 & n283;
  assign n3145 = n253 & n3144;
  assign n3146 = n273 & n3145;
  assign n3147 = ~n262 & n3146;
  assign n3148 = ~n3138 & ~n3140;
  assign n3149 = ~n3143 & n3148;
  assign n3150 = ~n286 & ~n3147;
  assign n3151 = n3149 & n3150;
  assign n3152 = n1718 & ~n3151;
  assign n3153 = n1737 & ~n3151;
  assign n3154 = ~n1718 & n3153;
  assign n3155 = ~n1737 & ~n3151;
  assign n3156 = ~n1718 & n3155;
  assign n3157 = n1742 & n3156;
  assign n3158 = ~n1742 & ~n3151;
  assign n3159 = ~n1718 & n3158;
  assign n3160 = ~n1737 & n3159;
  assign n3161 = n1748 & n3160;
  assign n3162 = ~n1748 & ~n3151;
  assign n3163 = ~n1737 & n3162;
  assign n3164 = ~n1718 & n3163;
  assign n3165 = ~n1742 & n3164;
  assign n3166 = n1753 & n3165;
  assign n3167 = ~n1753 & ~n3151;
  assign n3168 = ~n1742 & n3167;
  assign n3169 = ~n1718 & n3168;
  assign n3170 = ~n1737 & n3169;
  assign n3171 = ~n1748 & n3170;
  assign n3172 = pi005 & n3171;
  assign n3173 = ~pi005 & pi096;
  assign n3174 = ~n1748 & n3173;
  assign n3175 = ~n1737 & n3174;
  assign n3176 = ~n1718 & n3175;
  assign n3177 = ~n1742 & n3176;
  assign n3178 = ~n1753 & n3177;
  assign n3179 = pi095 & n3178;
  assign n3180 = ~pi005 & n3179;
  assign n3181 = ~n3152 & ~n3154;
  assign n3182 = ~n3157 & ~n3161;
  assign n3183 = n3181 & n3182;
  assign n3184 = ~n3166 & ~n3172;
  assign n3185 = ~n3180 & n3184;
  assign po62 = ~n3183 | ~n3185;
  assign n3187 = pi087 & ~n253;
  assign n3188 = pi016 & ~n273;
  assign n3189 = n253 & n3188;
  assign n3190 = pi019 & n273;
  assign n3191 = n253 & n3190;
  assign n3192 = ~n283 & n3191;
  assign n3193 = pi023 & n283;
  assign n3194 = n253 & n3193;
  assign n3195 = n273 & n3194;
  assign n3196 = ~n262 & n3195;
  assign n3197 = ~n3187 & ~n3189;
  assign n3198 = ~n3192 & n3197;
  assign n3199 = ~n286 & ~n3196;
  assign n3200 = n3198 & n3199;
  assign n3201 = n1718 & ~n3200;
  assign n3202 = n1737 & ~n3200;
  assign n3203 = ~n1718 & n3202;
  assign n3204 = ~n1737 & ~n3200;
  assign n3205 = ~n1718 & n3204;
  assign n3206 = n1742 & n3205;
  assign n3207 = ~n1742 & ~n3200;
  assign n3208 = ~n1718 & n3207;
  assign n3209 = ~n1737 & n3208;
  assign n3210 = n1748 & n3209;
  assign n3211 = ~n1748 & ~n3200;
  assign n3212 = ~n1737 & n3211;
  assign n3213 = ~n1718 & n3212;
  assign n3214 = ~n1742 & n3213;
  assign n3215 = n1753 & n3214;
  assign n3216 = ~n1753 & ~n3200;
  assign n3217 = ~n1742 & n3216;
  assign n3218 = ~n1718 & n3217;
  assign n3219 = ~n1737 & n3218;
  assign n3220 = ~n1748 & n3219;
  assign n3221 = pi005 & n3220;
  assign n3222 = ~pi005 & pi090;
  assign n3223 = ~n1748 & n3222;
  assign n3224 = ~n1737 & n3223;
  assign n3225 = ~n1718 & n3224;
  assign n3226 = ~n1742 & n3225;
  assign n3227 = ~n1753 & n3226;
  assign n3228 = pi095 & n3227;
  assign n3229 = ~pi005 & n3228;
  assign n3230 = ~n3201 & ~n3203;
  assign n3231 = ~n3206 & ~n3210;
  assign n3232 = n3230 & n3231;
  assign n3233 = ~n3215 & ~n3221;
  assign n3234 = ~n3229 & n3233;
  assign po63 = ~n3232 | ~n3234;
  assign n3236 = ~pi006 & n842;
  assign n3237 = ~pi130 & n3236;
  assign n3238 = ~pi004 & n3237;
  assign n3239 = pi067 & n3238;
  assign n3240 = pi007 & n842;
  assign n3241 = pi067 & n3240;
  assign n3242 = ~n3238 & n3241;
  assign n3243 = pi067 & ~n3240;
  assign n3244 = ~n3238 & n3243;
  assign n3245 = pi005 & n3244;
  assign n3246 = ~pi001 & ~pi132;
  assign n3247 = ~pi002 & n3246;
  assign n3248 = ~pi131 & n3247;
  assign n3249 = ~pi005 & n3248;
  assign n3250 = pi004 & n3249;
  assign n3251 = ~pi095 & n3250;
  assign n3252 = ~pi007 & n3251;
  assign n3253 = ~n3240 & n3252;
  assign n3254 = ~n3238 & n3253;
  assign n3255 = ~pi005 & n3254;
  assign n3256 = pi108 & ~n3252;
  assign n3257 = ~n3240 & n3256;
  assign n3258 = ~n3238 & n3257;
  assign n3259 = ~pi005 & n3258;
  assign n3260 = pi095 & n3259;
  assign n3261 = ~pi005 & n3260;
  assign n3262 = ~n3239 & ~n3242;
  assign n3263 = ~n3245 & n3262;
  assign n3264 = ~n3255 & ~n3261;
  assign po64 = ~n3263 | ~n3264;
  assign n3266 = pi068 & n3238;
  assign n3267 = pi068 & n3240;
  assign n3268 = ~n3238 & n3267;
  assign n3269 = pi068 & ~n3240;
  assign n3270 = ~n3238 & n3269;
  assign n3271 = pi005 & n3270;
  assign n3272 = pi109 & ~n3252;
  assign n3273 = ~n3240 & n3272;
  assign n3274 = ~n3238 & n3273;
  assign n3275 = ~pi005 & n3274;
  assign n3276 = pi095 & n3275;
  assign n3277 = ~pi005 & n3276;
  assign n3278 = ~n3266 & ~n3268;
  assign n3279 = ~n3271 & n3278;
  assign n3280 = ~n3255 & ~n3277;
  assign po65 = ~n3279 | ~n3280;
  assign n3282 = pi069 & n3238;
  assign n3283 = pi069 & n3240;
  assign n3284 = ~n3238 & n3283;
  assign n3285 = pi069 & ~n3240;
  assign n3286 = ~n3238 & n3285;
  assign n3287 = pi005 & n3286;
  assign n3288 = pi106 & ~n3252;
  assign n3289 = ~n3240 & n3288;
  assign n3290 = ~n3238 & n3289;
  assign n3291 = ~pi005 & n3290;
  assign n3292 = pi095 & n3291;
  assign n3293 = ~pi005 & n3292;
  assign n3294 = ~n3282 & ~n3284;
  assign n3295 = ~n3287 & n3294;
  assign n3296 = ~n3255 & ~n3293;
  assign po66 = ~n3295 | ~n3296;
  assign n3298 = pi070 & n3238;
  assign n3299 = pi070 & n3240;
  assign n3300 = ~n3238 & n3299;
  assign n3301 = pi070 & ~n3240;
  assign n3302 = ~n3238 & n3301;
  assign n3303 = pi005 & n3302;
  assign n3304 = pi104 & ~n3252;
  assign n3305 = ~n3240 & n3304;
  assign n3306 = ~n3238 & n3305;
  assign n3307 = ~pi005 & n3306;
  assign n3308 = pi095 & n3307;
  assign n3309 = ~pi005 & n3308;
  assign n3310 = ~n3298 & ~n3300;
  assign n3311 = ~n3303 & n3310;
  assign n3312 = ~n3255 & ~n3309;
  assign po67 = ~n3311 | ~n3312;
  assign n3314 = pi071 & n3238;
  assign n3315 = pi071 & n3240;
  assign n3316 = ~n3238 & n3315;
  assign n3317 = pi071 & ~n3240;
  assign n3318 = ~n3238 & n3317;
  assign n3319 = pi005 & n3318;
  assign n3320 = pi105 & ~n3252;
  assign n3321 = ~n3240 & n3320;
  assign n3322 = ~n3238 & n3321;
  assign n3323 = ~pi005 & n3322;
  assign n3324 = pi095 & n3323;
  assign n3325 = ~pi005 & n3324;
  assign n3326 = ~n3314 & ~n3316;
  assign n3327 = ~n3319 & n3326;
  assign n3328 = ~n3255 & ~n3325;
  assign po68 = ~n3327 | ~n3328;
  assign n3330 = pi072 & n3238;
  assign n3331 = pi072 & n3240;
  assign n3332 = ~n3238 & n3331;
  assign n3333 = pi072 & ~n3240;
  assign n3334 = ~n3238 & n3333;
  assign n3335 = pi005 & n3334;
  assign n3336 = pi103 & ~n3252;
  assign n3337 = ~n3240 & n3336;
  assign n3338 = ~n3238 & n3337;
  assign n3339 = ~pi005 & n3338;
  assign n3340 = pi095 & n3339;
  assign n3341 = ~pi005 & n3340;
  assign n3342 = ~n3330 & ~n3332;
  assign n3343 = ~n3335 & n3342;
  assign n3344 = ~n3255 & ~n3341;
  assign po69 = ~n3343 | ~n3344;
  assign n3346 = pi073 & n3238;
  assign n3347 = pi073 & n3240;
  assign n3348 = ~n3238 & n3347;
  assign n3349 = pi073 & ~n3240;
  assign n3350 = ~n3238 & n3349;
  assign n3351 = pi005 & n3350;
  assign n3352 = pi097 & ~n3252;
  assign n3353 = ~n3240 & n3352;
  assign n3354 = ~n3238 & n3353;
  assign n3355 = ~pi005 & n3354;
  assign n3356 = pi095 & n3355;
  assign n3357 = ~pi005 & n3356;
  assign n3358 = ~n3346 & ~n3348;
  assign n3359 = ~n3351 & n3358;
  assign n3360 = ~n3255 & ~n3357;
  assign po70 = ~n3359 | ~n3360;
  assign n3362 = pi074 & n3238;
  assign n3363 = pi074 & n3240;
  assign n3364 = ~n3238 & n3363;
  assign n3365 = pi074 & ~n3240;
  assign n3366 = ~n3238 & n3365;
  assign n3367 = pi005 & n3366;
  assign n3368 = pi098 & ~n3252;
  assign n3369 = ~n3240 & n3368;
  assign n3370 = ~n3238 & n3369;
  assign n3371 = ~pi005 & n3370;
  assign n3372 = pi095 & n3371;
  assign n3373 = ~pi005 & n3372;
  assign n3374 = ~n3362 & ~n3364;
  assign n3375 = ~n3367 & n3374;
  assign n3376 = ~n3255 & ~n3373;
  assign po71 = ~n3375 | ~n3376;
  assign n3378 = pi075 & n3238;
  assign n3379 = pi075 & n3240;
  assign n3380 = ~n3238 & n3379;
  assign n3381 = pi075 & ~n3240;
  assign n3382 = ~n3238 & n3381;
  assign n3383 = pi005 & n3382;
  assign n3384 = pi099 & ~n3252;
  assign n3385 = ~n3240 & n3384;
  assign n3386 = ~n3238 & n3385;
  assign n3387 = ~pi005 & n3386;
  assign n3388 = pi095 & n3387;
  assign n3389 = ~pi005 & n3388;
  assign n3390 = ~n3378 & ~n3380;
  assign n3391 = ~n3383 & n3390;
  assign n3392 = ~n3255 & ~n3389;
  assign po72 = ~n3391 | ~n3392;
  assign n3394 = pi076 & n3238;
  assign n3395 = pi076 & n3240;
  assign n3396 = ~n3238 & n3395;
  assign n3397 = pi076 & ~n3240;
  assign n3398 = ~n3238 & n3397;
  assign n3399 = pi005 & n3398;
  assign n3400 = pi100 & ~n3252;
  assign n3401 = ~n3240 & n3400;
  assign n3402 = ~n3238 & n3401;
  assign n3403 = ~pi005 & n3402;
  assign n3404 = pi095 & n3403;
  assign n3405 = ~pi005 & n3404;
  assign n3406 = ~n3394 & ~n3396;
  assign n3407 = ~n3399 & n3406;
  assign n3408 = ~n3255 & ~n3405;
  assign po73 = ~n3407 | ~n3408;
  assign n3410 = pi077 & n3238;
  assign n3411 = pi077 & n3240;
  assign n3412 = ~n3238 & n3411;
  assign n3413 = pi077 & ~n3240;
  assign n3414 = ~n3238 & n3413;
  assign n3415 = pi005 & n3414;
  assign n3416 = pi101 & ~n3252;
  assign n3417 = ~n3240 & n3416;
  assign n3418 = ~n3238 & n3417;
  assign n3419 = ~pi005 & n3418;
  assign n3420 = pi095 & n3419;
  assign n3421 = ~pi005 & n3420;
  assign n3422 = ~n3410 & ~n3412;
  assign n3423 = ~n3415 & n3422;
  assign n3424 = ~n3255 & ~n3421;
  assign po74 = ~n3423 | ~n3424;
  assign n3426 = pi078 & n3238;
  assign n3427 = pi078 & n3240;
  assign n3428 = ~n3238 & n3427;
  assign n3429 = pi078 & ~n3240;
  assign n3430 = ~n3238 & n3429;
  assign n3431 = pi005 & n3430;
  assign n3432 = pi102 & ~n3252;
  assign n3433 = ~n3240 & n3432;
  assign n3434 = ~n3238 & n3433;
  assign n3435 = ~pi005 & n3434;
  assign n3436 = pi095 & n3435;
  assign n3437 = ~pi005 & n3436;
  assign n3438 = ~n3426 & ~n3428;
  assign n3439 = ~n3431 & n3438;
  assign n3440 = ~n3255 & ~n3437;
  assign po75 = ~n3439 | ~n3440;
  assign n3442 = pi079 & n3238;
  assign n3443 = pi079 & n3240;
  assign n3444 = ~n3238 & n3443;
  assign n3445 = pi079 & ~n3240;
  assign n3446 = ~n3238 & n3445;
  assign n3447 = pi005 & n3446;
  assign n3448 = pi094 & ~n3252;
  assign n3449 = ~n3240 & n3448;
  assign n3450 = ~n3238 & n3449;
  assign n3451 = ~pi005 & n3450;
  assign n3452 = pi095 & n3451;
  assign n3453 = ~pi005 & n3452;
  assign n3454 = ~n3442 & ~n3444;
  assign n3455 = ~n3447 & n3454;
  assign n3456 = ~n3255 & ~n3453;
  assign po76 = ~n3455 | ~n3456;
  assign n3458 = pi080 & n3238;
  assign n3459 = pi080 & n3240;
  assign n3460 = ~n3238 & n3459;
  assign n3461 = pi080 & ~n3240;
  assign n3462 = ~n3238 & n3461;
  assign n3463 = pi005 & n3462;
  assign n3464 = pi096 & ~n3252;
  assign n3465 = ~n3240 & n3464;
  assign n3466 = ~n3238 & n3465;
  assign n3467 = ~pi005 & n3466;
  assign n3468 = pi095 & n3467;
  assign n3469 = ~pi005 & n3468;
  assign n3470 = ~n3458 & ~n3460;
  assign n3471 = ~n3463 & n3470;
  assign n3472 = ~n3255 & ~n3469;
  assign po77 = ~n3471 | ~n3472;
  assign n3474 = pi081 & n3238;
  assign n3475 = pi081 & n3240;
  assign n3476 = ~n3238 & n3475;
  assign n3477 = pi081 & ~n3240;
  assign n3478 = ~n3238 & n3477;
  assign n3479 = pi005 & n3478;
  assign n3480 = pi090 & ~n3252;
  assign n3481 = ~n3240 & n3480;
  assign n3482 = ~n3238 & n3481;
  assign n3483 = ~pi005 & n3482;
  assign n3484 = pi095 & n3483;
  assign n3485 = ~pi005 & n3484;
  assign n3486 = ~n3474 & ~n3476;
  assign n3487 = ~n3479 & n3486;
  assign n3488 = ~n3255 & ~n3485;
  assign po78 = ~n3487 | ~n3488;
  assign n3490 = ~pi008 & n219;
  assign n3491 = pi007 & n3490;
  assign n3492 = pi126 & n3491;
  assign n3493 = pi002 & n263;
  assign n3494 = ~pi005 & ~n307;
  assign n3495 = ~n228 & n3494;
  assign n3496 = ~n3491 & n3495;
  assign n3497 = ~n3493 & n3496;
  assign n3498 = ~n306 & n3497;
  assign n3499 = ~pi005 & n307;
  assign n3500 = ~n228 & n3499;
  assign n3501 = ~n3491 & n3500;
  assign n3502 = ~n3493 & n3501;
  assign n3503 = ~n306 & n3502;
  assign n3504 = pi127 & ~n3493;
  assign n3505 = ~n3491 & n3504;
  assign n3506 = ~n228 & n3505;
  assign n3507 = pi005 & n3506;
  assign n3508 = n306 & ~n3493;
  assign n3509 = ~n3491 & n3508;
  assign n3510 = ~n228 & n3509;
  assign n3511 = ~pi005 & n3510;
  assign n3512 = ~n3492 & ~n3498;
  assign n3513 = ~n3503 & n3512;
  assign n3514 = ~n3507 & ~n3511;
  assign po79 = ~n3513 | ~n3514;
  assign n3516 = pi007 & n219;
  assign n3517 = pi128 & n3516;
  assign n3518 = ~pi095 & n3493;
  assign n3519 = ~n3516 & n3518;
  assign n3520 = pi129 & ~n3518;
  assign n3521 = ~n3516 & n3520;
  assign n3522 = pi005 & n3521;
  assign n3523 = ~n3517 & ~n3519;
  assign po80 = n3522 | ~n3523;
endmodule



// Benchmark "i7" written by ABC on Sun Apr 22 21:43:05 2018

module i7 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66;
  wire n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088,
    n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169;
  assign n267 = ~pi000 & pi001;
  assign n268 = pi002 & n267;
  assign n269 = ~pi000 & pi030;
  assign n270 = ~pi002 & n269;
  assign n271 = pi000 & pi058;
  assign n272 = pi002 & n271;
  assign n273 = pi000 & ~pi030;
  assign n274 = ~pi002 & n273;
  assign n275 = ~n272 & ~n274;
  assign n276 = ~n268 & ~n270;
  assign po00 = ~n275 | ~n276;
  assign n278 = ~pi000 & pi003;
  assign n279 = pi002 & n278;
  assign n280 = ~pi000 & pi031;
  assign n281 = ~pi002 & n280;
  assign n282 = pi000 & pi059;
  assign n283 = pi002 & n282;
  assign n284 = pi000 & ~pi031;
  assign n285 = ~pi002 & n284;
  assign n286 = ~n283 & ~n285;
  assign n287 = ~n279 & ~n281;
  assign po01 = ~n286 | ~n287;
  assign n289 = ~pi000 & pi004;
  assign n290 = pi002 & n289;
  assign n291 = ~pi000 & pi032;
  assign n292 = ~pi002 & n291;
  assign n293 = pi000 & pi060;
  assign n294 = pi002 & n293;
  assign n295 = pi000 & ~pi032;
  assign n296 = ~pi002 & n295;
  assign n297 = ~n294 & ~n296;
  assign n298 = ~n290 & ~n292;
  assign po02 = ~n297 | ~n298;
  assign n300 = ~pi000 & pi005;
  assign n301 = pi002 & n300;
  assign n302 = ~pi000 & pi033;
  assign n303 = ~pi002 & n302;
  assign n304 = pi000 & pi061;
  assign n305 = pi002 & n304;
  assign n306 = pi000 & ~pi033;
  assign n307 = ~pi002 & n306;
  assign n308 = ~n305 & ~n307;
  assign n309 = ~n301 & ~n303;
  assign po03 = ~n308 | ~n309;
  assign n311 = ~pi000 & pi006;
  assign n312 = pi002 & n311;
  assign n313 = ~pi000 & pi034;
  assign n314 = ~pi002 & n313;
  assign n315 = pi000 & pi062;
  assign n316 = pi002 & n315;
  assign n317 = pi000 & ~pi034;
  assign n318 = ~pi002 & n317;
  assign n319 = ~n316 & ~n318;
  assign n320 = ~n312 & ~n314;
  assign po04 = ~n319 | ~n320;
  assign n322 = ~pi000 & pi007;
  assign n323 = pi002 & n322;
  assign n324 = ~pi000 & pi035;
  assign n325 = ~pi002 & n324;
  assign n326 = pi000 & pi063;
  assign n327 = pi002 & n326;
  assign n328 = pi000 & ~pi035;
  assign n329 = ~pi002 & n328;
  assign n330 = ~n327 & ~n329;
  assign n331 = ~n323 & ~n325;
  assign po05 = ~n330 | ~n331;
  assign n333 = ~pi000 & pi008;
  assign n334 = pi002 & n333;
  assign n335 = ~pi000 & pi036;
  assign n336 = ~pi002 & n335;
  assign n337 = pi000 & pi064;
  assign n338 = pi002 & n337;
  assign n339 = pi000 & ~pi036;
  assign n340 = ~pi002 & n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = ~n334 & ~n336;
  assign po06 = ~n341 | ~n342;
  assign n344 = ~pi000 & pi009;
  assign n345 = pi002 & n344;
  assign n346 = ~pi000 & pi037;
  assign n347 = ~pi002 & n346;
  assign n348 = pi000 & pi065;
  assign n349 = pi002 & n348;
  assign n350 = pi000 & ~pi037;
  assign n351 = ~pi002 & n350;
  assign n352 = ~n349 & ~n351;
  assign n353 = ~n345 & ~n347;
  assign po07 = ~n352 | ~n353;
  assign n355 = ~pi000 & pi010;
  assign n356 = pi002 & n355;
  assign n357 = ~pi000 & pi038;
  assign n358 = ~pi002 & n357;
  assign n359 = pi000 & pi066;
  assign n360 = pi002 & n359;
  assign n361 = pi000 & ~pi038;
  assign n362 = ~pi002 & n361;
  assign n363 = ~n360 & ~n362;
  assign n364 = ~n356 & ~n358;
  assign po08 = ~n363 | ~n364;
  assign n366 = ~pi000 & pi011;
  assign n367 = pi002 & n366;
  assign n368 = ~pi000 & pi039;
  assign n369 = ~pi002 & n368;
  assign n370 = pi000 & pi067;
  assign n371 = pi002 & n370;
  assign n372 = pi000 & ~pi039;
  assign n373 = ~pi002 & n372;
  assign n374 = ~n371 & ~n373;
  assign n375 = ~n367 & ~n369;
  assign po09 = ~n374 | ~n375;
  assign n377 = ~pi000 & pi012;
  assign n378 = pi002 & n377;
  assign n379 = ~pi000 & pi040;
  assign n380 = ~pi002 & n379;
  assign n381 = pi000 & pi068;
  assign n382 = pi002 & n381;
  assign n383 = pi000 & ~pi040;
  assign n384 = ~pi002 & n383;
  assign n385 = ~n382 & ~n384;
  assign n386 = ~n378 & ~n380;
  assign po10 = ~n385 | ~n386;
  assign n388 = ~pi000 & pi013;
  assign n389 = pi002 & n388;
  assign n390 = ~pi000 & pi041;
  assign n391 = ~pi002 & n390;
  assign n392 = pi000 & pi069;
  assign n393 = pi002 & n392;
  assign n394 = pi000 & ~pi041;
  assign n395 = ~pi002 & n394;
  assign n396 = ~n393 & ~n395;
  assign n397 = ~n389 & ~n391;
  assign po11 = ~n396 | ~n397;
  assign n399 = ~pi000 & pi014;
  assign n400 = pi002 & n399;
  assign n401 = ~pi000 & pi042;
  assign n402 = ~pi002 & n401;
  assign n403 = pi000 & pi070;
  assign n404 = pi002 & n403;
  assign n405 = pi000 & ~pi042;
  assign n406 = ~pi002 & n405;
  assign n407 = ~n404 & ~n406;
  assign n408 = ~n400 & ~n402;
  assign po12 = ~n407 | ~n408;
  assign n410 = ~pi000 & pi015;
  assign n411 = pi002 & n410;
  assign n412 = ~pi000 & pi043;
  assign n413 = ~pi002 & n412;
  assign n414 = pi000 & pi071;
  assign n415 = pi002 & n414;
  assign n416 = pi000 & ~pi043;
  assign n417 = ~pi002 & n416;
  assign n418 = ~n415 & ~n417;
  assign n419 = ~n411 & ~n413;
  assign po13 = ~n418 | ~n419;
  assign n421 = ~pi000 & pi016;
  assign n422 = pi002 & n421;
  assign n423 = ~pi000 & pi044;
  assign n424 = ~pi002 & n423;
  assign n425 = pi000 & pi072;
  assign n426 = pi002 & n425;
  assign n427 = pi000 & ~pi044;
  assign n428 = ~pi002 & n427;
  assign n429 = ~n426 & ~n428;
  assign n430 = ~n422 & ~n424;
  assign po14 = ~n429 | ~n430;
  assign n432 = ~pi000 & pi017;
  assign n433 = pi002 & n432;
  assign n434 = ~pi000 & pi045;
  assign n435 = ~pi002 & n434;
  assign n436 = pi000 & pi073;
  assign n437 = pi002 & n436;
  assign n438 = pi000 & ~pi045;
  assign n439 = ~pi002 & n438;
  assign n440 = ~n437 & ~n439;
  assign n441 = ~n433 & ~n435;
  assign po15 = ~n440 | ~n441;
  assign n443 = ~pi000 & pi018;
  assign n444 = pi002 & n443;
  assign n445 = ~pi000 & pi046;
  assign n446 = ~pi002 & n445;
  assign n447 = pi000 & pi074;
  assign n448 = pi002 & n447;
  assign n449 = pi000 & ~pi046;
  assign n450 = ~pi002 & n449;
  assign n451 = ~n448 & ~n450;
  assign n452 = ~n444 & ~n446;
  assign po16 = ~n451 | ~n452;
  assign n454 = ~pi000 & pi019;
  assign n455 = pi002 & n454;
  assign n456 = ~pi000 & pi047;
  assign n457 = ~pi002 & n456;
  assign n458 = pi000 & pi075;
  assign n459 = pi002 & n458;
  assign n460 = pi000 & ~pi047;
  assign n461 = ~pi002 & n460;
  assign n462 = ~n459 & ~n461;
  assign n463 = ~n455 & ~n457;
  assign po17 = ~n462 | ~n463;
  assign n465 = ~pi000 & pi020;
  assign n466 = pi002 & n465;
  assign n467 = ~pi000 & pi048;
  assign n468 = ~pi002 & n467;
  assign n469 = pi000 & pi076;
  assign n470 = pi002 & n469;
  assign n471 = pi000 & ~pi048;
  assign n472 = ~pi002 & n471;
  assign n473 = ~n470 & ~n472;
  assign n474 = ~n466 & ~n468;
  assign po18 = ~n473 | ~n474;
  assign n476 = ~pi000 & pi021;
  assign n477 = pi002 & n476;
  assign n478 = ~pi000 & pi049;
  assign n479 = ~pi002 & n478;
  assign n480 = pi000 & pi077;
  assign n481 = pi002 & n480;
  assign n482 = pi000 & ~pi049;
  assign n483 = ~pi002 & n482;
  assign n484 = ~n481 & ~n483;
  assign n485 = ~n477 & ~n479;
  assign po19 = ~n484 | ~n485;
  assign n487 = ~pi000 & pi022;
  assign n488 = pi002 & n487;
  assign n489 = ~pi000 & pi050;
  assign n490 = ~pi002 & n489;
  assign n491 = pi000 & pi078;
  assign n492 = pi002 & n491;
  assign n493 = pi000 & ~pi050;
  assign n494 = ~pi002 & n493;
  assign n495 = ~n492 & ~n494;
  assign n496 = ~n488 & ~n490;
  assign po20 = ~n495 | ~n496;
  assign n498 = ~pi000 & pi023;
  assign n499 = pi002 & n498;
  assign n500 = ~pi000 & pi051;
  assign n501 = ~pi002 & n500;
  assign n502 = pi000 & pi079;
  assign n503 = pi002 & n502;
  assign n504 = pi000 & ~pi051;
  assign n505 = ~pi002 & n504;
  assign n506 = ~n503 & ~n505;
  assign n507 = ~n499 & ~n501;
  assign po21 = ~n506 | ~n507;
  assign n509 = ~pi000 & pi024;
  assign n510 = pi002 & n509;
  assign n511 = ~pi000 & pi052;
  assign n512 = ~pi002 & n511;
  assign n513 = pi000 & pi080;
  assign n514 = pi002 & n513;
  assign n515 = pi000 & ~pi052;
  assign n516 = ~pi002 & n515;
  assign n517 = ~n514 & ~n516;
  assign n518 = ~n510 & ~n512;
  assign po22 = ~n517 | ~n518;
  assign n520 = ~pi000 & pi025;
  assign n521 = pi002 & n520;
  assign n522 = ~pi000 & pi053;
  assign n523 = ~pi002 & n522;
  assign n524 = pi000 & pi081;
  assign n525 = pi002 & n524;
  assign n526 = pi000 & ~pi053;
  assign n527 = ~pi002 & n526;
  assign n528 = ~n525 & ~n527;
  assign n529 = ~n521 & ~n523;
  assign po23 = ~n528 | ~n529;
  assign n531 = ~pi000 & pi026;
  assign n532 = pi002 & n531;
  assign n533 = ~pi000 & pi054;
  assign n534 = ~pi002 & n533;
  assign n535 = pi000 & pi082;
  assign n536 = pi002 & n535;
  assign n537 = pi000 & ~pi054;
  assign n538 = ~pi002 & n537;
  assign n539 = ~n536 & ~n538;
  assign n540 = ~n532 & ~n534;
  assign po24 = ~n539 | ~n540;
  assign n542 = ~pi000 & pi027;
  assign n543 = pi002 & n542;
  assign n544 = ~pi000 & pi055;
  assign n545 = ~pi002 & n544;
  assign n546 = pi000 & pi083;
  assign n547 = pi002 & n546;
  assign n548 = pi000 & ~pi055;
  assign n549 = ~pi002 & n548;
  assign n550 = ~n547 & ~n549;
  assign n551 = ~n543 & ~n545;
  assign po25 = ~n550 | ~n551;
  assign n553 = ~pi000 & pi028;
  assign n554 = pi002 & n553;
  assign n555 = ~pi000 & pi056;
  assign n556 = ~pi002 & n555;
  assign n557 = pi000 & pi084;
  assign n558 = pi002 & n557;
  assign n559 = pi000 & ~pi056;
  assign n560 = ~pi002 & n559;
  assign n561 = ~n558 & ~n560;
  assign n562 = ~n554 & ~n556;
  assign po26 = ~n561 | ~n562;
  assign n564 = ~pi000 & pi029;
  assign n565 = pi002 & n564;
  assign n566 = ~pi000 & pi057;
  assign n567 = ~pi002 & n566;
  assign n568 = pi000 & pi085;
  assign n569 = pi002 & n568;
  assign n570 = pi000 & ~pi057;
  assign n571 = ~pi002 & n570;
  assign n572 = ~n569 & ~n571;
  assign n573 = ~n565 & ~n567;
  assign po27 = ~n572 | ~n573;
  assign n575 = pi002 & pi086;
  assign n576 = ~pi000 & n575;
  assign n577 = pi087 & n576;
  assign n578 = ~pi002 & pi119;
  assign n579 = ~pi000 & n578;
  assign n580 = pi087 & n579;
  assign n581 = pi002 & pi151;
  assign n582 = pi000 & n581;
  assign n583 = pi087 & n582;
  assign n584 = ~pi002 & ~pi119;
  assign n585 = pi000 & n584;
  assign n586 = pi087 & n585;
  assign n587 = pi000 & ~pi087;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~n577 & ~n580;
  assign n590 = ~n583 & n589;
  assign po28 = ~n588 | ~n590;
  assign n592 = pi002 & pi088;
  assign n593 = ~pi000 & n592;
  assign n594 = pi087 & n593;
  assign n595 = ~pi002 & pi120;
  assign n596 = ~pi000 & n595;
  assign n597 = pi087 & n596;
  assign n598 = pi002 & pi152;
  assign n599 = pi000 & n598;
  assign n600 = pi087 & n599;
  assign n601 = ~pi002 & ~pi120;
  assign n602 = pi000 & n601;
  assign n603 = pi087 & n602;
  assign n604 = ~n587 & ~n603;
  assign n605 = ~n594 & ~n597;
  assign n606 = ~n600 & n605;
  assign po29 = ~n604 | ~n606;
  assign n608 = pi002 & pi089;
  assign n609 = ~pi000 & n608;
  assign n610 = pi087 & n609;
  assign n611 = ~pi002 & pi121;
  assign n612 = ~pi000 & n611;
  assign n613 = pi087 & n612;
  assign n614 = pi002 & pi153;
  assign n615 = pi000 & n614;
  assign n616 = pi087 & n615;
  assign n617 = ~pi002 & ~pi121;
  assign n618 = pi000 & n617;
  assign n619 = pi087 & n618;
  assign n620 = ~n587 & ~n619;
  assign n621 = ~n610 & ~n613;
  assign n622 = ~n616 & n621;
  assign po30 = ~n620 | ~n622;
  assign n624 = pi002 & pi090;
  assign n625 = ~pi000 & n624;
  assign n626 = pi087 & n625;
  assign n627 = ~pi002 & pi122;
  assign n628 = ~pi000 & n627;
  assign n629 = pi087 & n628;
  assign n630 = pi002 & pi154;
  assign n631 = pi000 & n630;
  assign n632 = pi087 & n631;
  assign n633 = ~pi002 & ~pi122;
  assign n634 = pi000 & n633;
  assign n635 = pi087 & n634;
  assign n636 = ~n587 & ~n635;
  assign n637 = ~n626 & ~n629;
  assign n638 = ~n632 & n637;
  assign po31 = ~n636 | ~n638;
  assign n640 = pi002 & pi091;
  assign n641 = ~pi000 & n640;
  assign n642 = pi087 & n641;
  assign n643 = ~pi002 & pi123;
  assign n644 = ~pi000 & n643;
  assign n645 = pi087 & n644;
  assign n646 = pi002 & pi155;
  assign n647 = pi000 & n646;
  assign n648 = pi087 & n647;
  assign n649 = ~pi002 & ~pi123;
  assign n650 = pi000 & n649;
  assign n651 = pi087 & n650;
  assign n652 = ~n587 & ~n651;
  assign n653 = ~n642 & ~n645;
  assign n654 = ~n648 & n653;
  assign po32 = ~n652 | ~n654;
  assign n656 = pi002 & pi092;
  assign n657 = ~pi000 & n656;
  assign n658 = pi087 & n657;
  assign n659 = ~pi002 & pi124;
  assign n660 = ~pi000 & n659;
  assign n661 = pi087 & n660;
  assign n662 = pi002 & pi156;
  assign n663 = pi000 & n662;
  assign n664 = pi087 & n663;
  assign n665 = ~pi002 & ~pi124;
  assign n666 = pi000 & n665;
  assign n667 = pi087 & n666;
  assign n668 = ~n587 & ~n667;
  assign n669 = ~n658 & ~n661;
  assign n670 = ~n664 & n669;
  assign po33 = ~n668 | ~n670;
  assign n672 = pi002 & pi093;
  assign n673 = ~pi000 & n672;
  assign n674 = pi087 & n673;
  assign n675 = ~pi002 & pi125;
  assign n676 = ~pi000 & n675;
  assign n677 = pi087 & n676;
  assign n678 = pi002 & pi157;
  assign n679 = pi000 & n678;
  assign n680 = pi087 & n679;
  assign n681 = ~pi002 & ~pi125;
  assign n682 = pi000 & n681;
  assign n683 = pi087 & n682;
  assign n684 = ~n587 & ~n683;
  assign n685 = ~n674 & ~n677;
  assign n686 = ~n680 & n685;
  assign po34 = ~n684 | ~n686;
  assign n688 = pi002 & pi094;
  assign n689 = ~pi000 & n688;
  assign n690 = pi087 & n689;
  assign n691 = ~pi002 & pi126;
  assign n692 = ~pi000 & n691;
  assign n693 = pi087 & n692;
  assign n694 = pi002 & pi158;
  assign n695 = pi000 & n694;
  assign n696 = pi087 & n695;
  assign n697 = ~pi002 & ~pi126;
  assign n698 = pi000 & n697;
  assign n699 = pi087 & n698;
  assign n700 = ~n587 & ~n699;
  assign n701 = ~n690 & ~n693;
  assign n702 = ~n696 & n701;
  assign po35 = ~n700 | ~n702;
  assign n704 = pi002 & pi095;
  assign n705 = ~pi000 & n704;
  assign n706 = pi087 & n705;
  assign n707 = ~pi002 & pi127;
  assign n708 = ~pi000 & n707;
  assign n709 = pi087 & n708;
  assign n710 = pi002 & pi159;
  assign n711 = pi000 & n710;
  assign n712 = pi087 & n711;
  assign n713 = ~pi002 & ~pi127;
  assign n714 = pi000 & n713;
  assign n715 = pi087 & n714;
  assign n716 = ~n587 & ~n715;
  assign n717 = ~n706 & ~n709;
  assign n718 = ~n712 & n717;
  assign po36 = ~n716 | ~n718;
  assign n720 = pi002 & pi096;
  assign n721 = ~pi000 & n720;
  assign n722 = pi087 & n721;
  assign n723 = ~pi002 & pi128;
  assign n724 = ~pi000 & n723;
  assign n725 = pi087 & n724;
  assign n726 = pi002 & pi160;
  assign n727 = pi000 & n726;
  assign n728 = pi087 & n727;
  assign n729 = ~pi002 & ~pi128;
  assign n730 = pi000 & n729;
  assign n731 = pi087 & n730;
  assign n732 = ~n587 & ~n731;
  assign n733 = ~n722 & ~n725;
  assign n734 = ~n728 & n733;
  assign po37 = ~n732 | ~n734;
  assign n736 = pi002 & pi097;
  assign n737 = ~pi000 & n736;
  assign n738 = pi087 & n737;
  assign n739 = ~pi002 & pi129;
  assign n740 = ~pi000 & n739;
  assign n741 = pi087 & n740;
  assign n742 = pi002 & pi161;
  assign n743 = pi000 & n742;
  assign n744 = pi087 & n743;
  assign n745 = ~pi002 & ~pi129;
  assign n746 = pi000 & n745;
  assign n747 = pi087 & n746;
  assign n748 = ~n587 & ~n747;
  assign n749 = ~n738 & ~n741;
  assign n750 = ~n744 & n749;
  assign po38 = ~n748 | ~n750;
  assign n752 = pi002 & pi098;
  assign n753 = ~pi000 & n752;
  assign n754 = pi087 & n753;
  assign n755 = ~pi002 & pi130;
  assign n756 = ~pi000 & n755;
  assign n757 = pi087 & n756;
  assign n758 = pi002 & pi162;
  assign n759 = pi000 & n758;
  assign n760 = pi087 & n759;
  assign n761 = ~pi002 & ~pi130;
  assign n762 = pi000 & n761;
  assign n763 = pi087 & n762;
  assign n764 = ~n587 & ~n763;
  assign n765 = ~n754 & ~n757;
  assign n766 = ~n760 & n765;
  assign po39 = ~n764 | ~n766;
  assign n768 = pi002 & pi099;
  assign n769 = ~pi000 & n768;
  assign n770 = pi087 & n769;
  assign n771 = ~pi002 & pi131;
  assign n772 = ~pi000 & n771;
  assign n773 = pi087 & n772;
  assign n774 = pi002 & pi163;
  assign n775 = pi000 & n774;
  assign n776 = pi087 & n775;
  assign n777 = ~pi002 & ~pi131;
  assign n778 = pi000 & n777;
  assign n779 = pi087 & n778;
  assign n780 = ~n587 & ~n779;
  assign n781 = ~n770 & ~n773;
  assign n782 = ~n776 & n781;
  assign po40 = ~n780 | ~n782;
  assign n784 = pi002 & pi100;
  assign n785 = ~pi000 & n784;
  assign n786 = pi087 & n785;
  assign n787 = ~pi002 & pi132;
  assign n788 = ~pi000 & n787;
  assign n789 = pi087 & n788;
  assign n790 = pi002 & pi164;
  assign n791 = pi000 & n790;
  assign n792 = pi087 & n791;
  assign n793 = ~pi002 & ~pi132;
  assign n794 = pi000 & n793;
  assign n795 = pi087 & n794;
  assign n796 = ~n587 & ~n795;
  assign n797 = ~n786 & ~n789;
  assign n798 = ~n792 & n797;
  assign po41 = ~n796 | ~n798;
  assign n800 = pi002 & pi101;
  assign n801 = ~pi000 & n800;
  assign n802 = pi087 & n801;
  assign n803 = ~pi002 & pi133;
  assign n804 = ~pi000 & n803;
  assign n805 = pi087 & n804;
  assign n806 = pi002 & pi165;
  assign n807 = pi000 & n806;
  assign n808 = pi087 & n807;
  assign n809 = ~pi002 & ~pi133;
  assign n810 = pi000 & n809;
  assign n811 = pi087 & n810;
  assign n812 = ~n587 & ~n811;
  assign n813 = ~n802 & ~n805;
  assign n814 = ~n808 & n813;
  assign po42 = ~n812 | ~n814;
  assign n816 = pi002 & pi102;
  assign n817 = ~pi000 & n816;
  assign n818 = pi087 & n817;
  assign n819 = ~pi002 & pi134;
  assign n820 = ~pi000 & n819;
  assign n821 = pi087 & n820;
  assign n822 = pi002 & pi166;
  assign n823 = pi000 & n822;
  assign n824 = pi087 & n823;
  assign n825 = ~pi002 & ~pi134;
  assign n826 = pi000 & n825;
  assign n827 = pi087 & n826;
  assign n828 = ~n587 & ~n827;
  assign n829 = ~n818 & ~n821;
  assign n830 = ~n824 & n829;
  assign po43 = ~n828 | ~n830;
  assign n832 = pi002 & pi103;
  assign n833 = ~pi000 & n832;
  assign n834 = pi087 & n833;
  assign n835 = ~pi002 & pi135;
  assign n836 = ~pi000 & n835;
  assign n837 = pi087 & n836;
  assign n838 = pi002 & pi167;
  assign n839 = pi000 & n838;
  assign n840 = pi087 & n839;
  assign n841 = ~pi002 & ~pi135;
  assign n842 = pi000 & n841;
  assign n843 = pi087 & n842;
  assign n844 = ~n587 & ~n843;
  assign n845 = ~n834 & ~n837;
  assign n846 = ~n840 & n845;
  assign po44 = ~n844 | ~n846;
  assign n848 = pi002 & pi104;
  assign n849 = ~pi000 & n848;
  assign n850 = pi087 & n849;
  assign n851 = ~pi002 & pi136;
  assign n852 = ~pi000 & n851;
  assign n853 = pi087 & n852;
  assign n854 = pi002 & pi168;
  assign n855 = pi000 & n854;
  assign n856 = pi087 & n855;
  assign n857 = ~pi002 & ~pi136;
  assign n858 = pi000 & n857;
  assign n859 = pi087 & n858;
  assign n860 = ~n587 & ~n859;
  assign n861 = ~n850 & ~n853;
  assign n862 = ~n856 & n861;
  assign po45 = ~n860 | ~n862;
  assign n864 = pi002 & pi105;
  assign n865 = ~pi000 & n864;
  assign n866 = pi087 & n865;
  assign n867 = ~pi002 & pi137;
  assign n868 = ~pi000 & n867;
  assign n869 = pi087 & n868;
  assign n870 = pi002 & pi169;
  assign n871 = pi000 & n870;
  assign n872 = pi087 & n871;
  assign n873 = ~pi002 & ~pi137;
  assign n874 = pi000 & n873;
  assign n875 = pi087 & n874;
  assign n876 = ~n587 & ~n875;
  assign n877 = ~n866 & ~n869;
  assign n878 = ~n872 & n877;
  assign po46 = ~n876 | ~n878;
  assign n880 = pi002 & pi106;
  assign n881 = ~pi000 & n880;
  assign n882 = pi087 & n881;
  assign n883 = ~pi002 & pi138;
  assign n884 = ~pi000 & n883;
  assign n885 = pi087 & n884;
  assign n886 = pi002 & pi170;
  assign n887 = pi000 & n886;
  assign n888 = pi087 & n887;
  assign n889 = ~pi002 & ~pi138;
  assign n890 = pi000 & n889;
  assign n891 = pi087 & n890;
  assign n892 = ~n587 & ~n891;
  assign n893 = ~n882 & ~n885;
  assign n894 = ~n888 & n893;
  assign po47 = ~n892 | ~n894;
  assign n896 = pi002 & pi107;
  assign n897 = ~pi000 & n896;
  assign n898 = pi087 & n897;
  assign n899 = ~pi002 & pi139;
  assign n900 = ~pi000 & n899;
  assign n901 = pi087 & n900;
  assign n902 = pi002 & pi171;
  assign n903 = pi000 & n902;
  assign n904 = pi087 & n903;
  assign n905 = ~pi002 & ~pi139;
  assign n906 = pi000 & n905;
  assign n907 = pi087 & n906;
  assign n908 = ~n587 & ~n907;
  assign n909 = ~n898 & ~n901;
  assign n910 = ~n904 & n909;
  assign po48 = ~n908 | ~n910;
  assign n912 = pi002 & pi108;
  assign n913 = ~pi000 & n912;
  assign n914 = pi087 & n913;
  assign n915 = ~pi002 & pi140;
  assign n916 = ~pi000 & n915;
  assign n917 = pi087 & n916;
  assign n918 = pi002 & pi172;
  assign n919 = pi000 & n918;
  assign n920 = pi087 & n919;
  assign n921 = ~pi002 & ~pi140;
  assign n922 = pi000 & n921;
  assign n923 = pi087 & n922;
  assign n924 = ~n587 & ~n923;
  assign n925 = ~n914 & ~n917;
  assign n926 = ~n920 & n925;
  assign po49 = ~n924 | ~n926;
  assign n928 = pi002 & pi109;
  assign n929 = ~pi000 & n928;
  assign n930 = pi087 & n929;
  assign n931 = ~pi002 & pi141;
  assign n932 = ~pi000 & n931;
  assign n933 = pi087 & n932;
  assign n934 = pi002 & pi173;
  assign n935 = pi000 & n934;
  assign n936 = pi087 & n935;
  assign n937 = ~pi002 & ~pi141;
  assign n938 = pi000 & n937;
  assign n939 = pi087 & n938;
  assign n940 = ~n587 & ~n939;
  assign n941 = ~n930 & ~n933;
  assign n942 = ~n936 & n941;
  assign po50 = ~n940 | ~n942;
  assign n944 = pi002 & pi110;
  assign n945 = ~pi000 & n944;
  assign n946 = pi087 & n945;
  assign n947 = ~pi002 & pi142;
  assign n948 = ~pi000 & n947;
  assign n949 = pi087 & n948;
  assign n950 = pi002 & pi174;
  assign n951 = pi000 & n950;
  assign n952 = pi087 & n951;
  assign n953 = ~pi002 & ~pi142;
  assign n954 = pi000 & n953;
  assign n955 = pi087 & n954;
  assign n956 = ~n587 & ~n955;
  assign n957 = ~n946 & ~n949;
  assign n958 = ~n952 & n957;
  assign po51 = ~n956 | ~n958;
  assign n960 = pi002 & pi111;
  assign n961 = ~pi000 & n960;
  assign n962 = pi087 & n961;
  assign n963 = ~pi002 & pi143;
  assign n964 = ~pi000 & n963;
  assign n965 = pi087 & n964;
  assign n966 = pi002 & pi175;
  assign n967 = pi000 & n966;
  assign n968 = pi087 & n967;
  assign n969 = ~pi002 & ~pi143;
  assign n970 = pi000 & n969;
  assign n971 = pi087 & n970;
  assign n972 = ~n587 & ~n971;
  assign n973 = ~n962 & ~n965;
  assign n974 = ~n968 & n973;
  assign po52 = ~n972 | ~n974;
  assign n976 = pi002 & pi112;
  assign n977 = ~pi000 & n976;
  assign n978 = pi087 & n977;
  assign n979 = ~pi002 & pi144;
  assign n980 = ~pi000 & n979;
  assign n981 = pi087 & n980;
  assign n982 = pi002 & pi176;
  assign n983 = pi000 & n982;
  assign n984 = pi087 & n983;
  assign n985 = ~pi002 & ~pi144;
  assign n986 = pi000 & n985;
  assign n987 = pi087 & n986;
  assign n988 = ~n587 & ~n987;
  assign n989 = ~n978 & ~n981;
  assign n990 = ~n984 & n989;
  assign po53 = ~n988 | ~n990;
  assign n992 = pi002 & pi113;
  assign n993 = ~pi000 & n992;
  assign n994 = pi087 & n993;
  assign n995 = ~pi002 & pi145;
  assign n996 = ~pi000 & n995;
  assign n997 = pi087 & n996;
  assign n998 = pi002 & pi177;
  assign n999 = pi000 & n998;
  assign n1000 = pi087 & n999;
  assign n1001 = ~pi002 & ~pi145;
  assign n1002 = pi000 & n1001;
  assign n1003 = pi087 & n1002;
  assign n1004 = ~n587 & ~n1003;
  assign n1005 = ~n994 & ~n997;
  assign n1006 = ~n1000 & n1005;
  assign po54 = ~n1004 | ~n1006;
  assign n1008 = pi002 & pi114;
  assign n1009 = ~pi000 & n1008;
  assign n1010 = pi087 & n1009;
  assign n1011 = ~pi002 & pi146;
  assign n1012 = ~pi000 & n1011;
  assign n1013 = pi087 & n1012;
  assign n1014 = pi002 & pi178;
  assign n1015 = pi000 & n1014;
  assign n1016 = pi087 & n1015;
  assign n1017 = ~pi002 & ~pi146;
  assign n1018 = pi000 & n1017;
  assign n1019 = pi087 & n1018;
  assign n1020 = ~n587 & ~n1019;
  assign n1021 = ~n1010 & ~n1013;
  assign n1022 = ~n1016 & n1021;
  assign po55 = ~n1020 | ~n1022;
  assign n1024 = pi002 & pi115;
  assign n1025 = ~pi000 & n1024;
  assign n1026 = pi087 & n1025;
  assign n1027 = ~pi002 & pi147;
  assign n1028 = ~pi000 & n1027;
  assign n1029 = pi087 & n1028;
  assign n1030 = pi002 & pi179;
  assign n1031 = pi000 & n1030;
  assign n1032 = pi087 & n1031;
  assign n1033 = ~pi002 & ~pi147;
  assign n1034 = pi000 & n1033;
  assign n1035 = pi087 & n1034;
  assign n1036 = ~n587 & ~n1035;
  assign n1037 = ~n1026 & ~n1029;
  assign n1038 = ~n1032 & n1037;
  assign po56 = ~n1036 | ~n1038;
  assign n1040 = pi002 & pi116;
  assign n1041 = ~pi000 & n1040;
  assign n1042 = pi087 & n1041;
  assign n1043 = ~pi002 & pi148;
  assign n1044 = ~pi000 & n1043;
  assign n1045 = pi087 & n1044;
  assign n1046 = pi002 & pi180;
  assign n1047 = pi000 & n1046;
  assign n1048 = pi087 & n1047;
  assign n1049 = ~pi002 & ~pi148;
  assign n1050 = pi000 & n1049;
  assign n1051 = pi087 & n1050;
  assign n1052 = ~n587 & ~n1051;
  assign n1053 = ~n1042 & ~n1045;
  assign n1054 = ~n1048 & n1053;
  assign po57 = ~n1052 | ~n1054;
  assign n1056 = pi002 & pi117;
  assign n1057 = ~pi000 & n1056;
  assign n1058 = pi087 & n1057;
  assign n1059 = ~pi002 & pi149;
  assign n1060 = ~pi000 & n1059;
  assign n1061 = pi087 & n1060;
  assign n1062 = pi002 & pi181;
  assign n1063 = pi000 & n1062;
  assign n1064 = pi087 & n1063;
  assign n1065 = ~pi002 & ~pi149;
  assign n1066 = pi000 & n1065;
  assign n1067 = pi087 & n1066;
  assign n1068 = ~n587 & ~n1067;
  assign n1069 = ~n1058 & ~n1061;
  assign n1070 = ~n1064 & n1069;
  assign po58 = ~n1068 | ~n1070;
  assign n1072 = pi002 & pi118;
  assign n1073 = ~pi000 & n1072;
  assign n1074 = pi087 & n1073;
  assign n1075 = ~pi002 & pi150;
  assign n1076 = ~pi000 & n1075;
  assign n1077 = pi087 & n1076;
  assign n1078 = pi002 & pi182;
  assign n1079 = pi000 & n1078;
  assign n1080 = pi087 & n1079;
  assign n1081 = ~pi002 & ~pi150;
  assign n1082 = pi000 & n1081;
  assign n1083 = pi087 & n1082;
  assign n1084 = ~n587 & ~n1083;
  assign n1085 = ~n1074 & ~n1077;
  assign n1086 = ~n1080 & n1085;
  assign po59 = ~n1084 | ~n1086;
  assign n1088 = ~pi002 & pi188;
  assign n1089 = pi000 & n1088;
  assign n1090 = pi184 & n1089;
  assign n1091 = ~pi000 & n1088;
  assign n1092 = pi184 & n1091;
  assign po60 = n1090 | n1092;
  assign n1094 = pi000 & ~pi184;
  assign n1095 = ~pi002 & pi189;
  assign n1096 = ~pi000 & n1095;
  assign n1097 = pi184 & n1096;
  assign n1098 = pi000 & pi184;
  assign n1099 = pi002 & n1098;
  assign n1100 = ~pi002 & ~pi189;
  assign n1101 = pi000 & n1100;
  assign n1102 = pi184 & n1101;
  assign n1103 = ~n1099 & ~n1102;
  assign n1104 = ~n1094 & ~n1097;
  assign po61 = ~n1103 | ~n1104;
  assign n1106 = ~pi002 & pi190;
  assign n1107 = ~pi000 & n1106;
  assign n1108 = pi184 & n1107;
  assign n1109 = ~pi002 & ~pi190;
  assign n1110 = pi000 & n1109;
  assign n1111 = pi184 & n1110;
  assign n1112 = ~n1099 & ~n1111;
  assign n1113 = ~n1094 & ~n1108;
  assign po62 = ~n1112 | ~n1113;
  assign n1115 = pi002 & pi183;
  assign n1116 = ~pi000 & n1115;
  assign n1117 = pi184 & n1116;
  assign n1118 = ~pi002 & pi191;
  assign n1119 = ~pi000 & n1118;
  assign n1120 = pi184 & n1119;
  assign n1121 = pi195 & n1099;
  assign n1122 = ~pi002 & ~pi191;
  assign n1123 = pi000 & n1122;
  assign n1124 = pi184 & n1123;
  assign n1125 = ~n1094 & ~n1124;
  assign n1126 = ~n1117 & ~n1120;
  assign n1127 = ~n1121 & n1126;
  assign po63 = ~n1125 | ~n1127;
  assign n1129 = pi002 & pi185;
  assign n1130 = ~pi000 & n1129;
  assign n1131 = pi184 & n1130;
  assign n1132 = ~pi002 & pi192;
  assign n1133 = ~pi000 & n1132;
  assign n1134 = pi184 & n1133;
  assign n1135 = pi196 & n1099;
  assign n1136 = ~pi002 & ~pi192;
  assign n1137 = pi000 & n1136;
  assign n1138 = pi184 & n1137;
  assign n1139 = ~n1094 & ~n1138;
  assign n1140 = ~n1131 & ~n1134;
  assign n1141 = ~n1135 & n1140;
  assign po64 = ~n1139 | ~n1141;
  assign n1143 = pi002 & pi186;
  assign n1144 = ~pi000 & n1143;
  assign n1145 = pi184 & n1144;
  assign n1146 = ~pi002 & pi193;
  assign n1147 = ~pi000 & n1146;
  assign n1148 = pi184 & n1147;
  assign n1149 = pi197 & n1099;
  assign n1150 = ~pi002 & ~pi193;
  assign n1151 = pi000 & n1150;
  assign n1152 = pi184 & n1151;
  assign n1153 = ~n1094 & ~n1152;
  assign n1154 = ~n1145 & ~n1148;
  assign n1155 = ~n1149 & n1154;
  assign po65 = ~n1153 | ~n1155;
  assign n1157 = pi002 & pi187;
  assign n1158 = ~pi000 & n1157;
  assign n1159 = pi184 & n1158;
  assign n1160 = ~pi002 & pi194;
  assign n1161 = ~pi000 & n1160;
  assign n1162 = pi184 & n1161;
  assign n1163 = pi198 & n1099;
  assign n1164 = ~pi002 & ~pi194;
  assign n1165 = pi000 & n1164;
  assign n1166 = pi184 & n1165;
  assign n1167 = ~n1094 & ~n1166;
  assign n1168 = ~n1159 & ~n1162;
  assign n1169 = ~n1163 & n1168;
  assign po66 = ~n1167 | ~n1169;
endmodule



// Benchmark "alu4_cl" written by ABC on Sun Apr 22 21:42:56 2018

module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
    n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n529, n530, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756;
  assign n23 = ~pi08 & pi11;
  assign n24 = ~pi09 & pi10;
  assign n25 = ~pi10 & ~pi11;
  assign n26 = pi08 & pi09;
  assign n27 = n25 & n26;
  assign n28 = pi13 & n27;
  assign n29 = n23 & n24;
  assign n30 = ~pi13 & n29;
  assign n31 = ~n28 & ~n30;
  assign n32 = pi10 & ~pi11;
  assign n33 = ~pi08 & n32;
  assign n34 = ~pi10 & n26;
  assign n35 = pi11 & n34;
  assign n36 = pi09 & n33;
  assign n37 = ~n35 & ~n36;
  assign n38 = pi08 & ~pi09;
  assign n39 = ~pi09 & ~pi11;
  assign n40 = ~pi08 & ~pi10;
  assign n41 = pi08 & pi10;
  assign n42 = ~pi08 & pi09;
  assign n43 = n26 & n32;
  assign n44 = ~n32 & n42;
  assign n45 = pi13 & n44;
  assign n46 = ~pi09 & pi11;
  assign n47 = ~pi13 & n41;
  assign n48 = n46 & n47;
  assign n49 = ~n45 & ~n48;
  assign n50 = ~n43 & n49;
  assign n51 = ~pi08 & ~pi09;
  assign n52 = ~n26 & ~n51;
  assign n53 = pi11 & ~n52;
  assign n54 = ~pi10 & n53;
  assign n55 = pi13 & n54;
  assign n56 = ~pi09 & n33;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~pi00 & ~pi04;
  assign n59 = pi10 & pi13;
  assign n60 = ~pi13 & n25;
  assign n61 = ~n59 & ~n60;
  assign n62 = n38 & ~n61;
  assign n63 = pi09 & pi11;
  assign n64 = ~pi13 & ~n63;
  assign n65 = n40 & n64;
  assign n66 = pi00 & pi04;
  assign n67 = pi00 & ~pi04;
  assign n68 = ~pi00 & pi04;
  assign n69 = n32 & n68;
  assign n70 = ~n67 & ~n69;
  assign n71 = pi13 & ~n70;
  assign n72 = n42 & n71;
  assign n73 = ~n58 & n62;
  assign n74 = ~n57 & n66;
  assign n75 = ~n73 & ~n74;
  assign n76 = ~pi00 & n65;
  assign n77 = ~pi04 & ~n50;
  assign n78 = ~n76 & ~n77;
  assign n79 = n75 & n78;
  assign n80 = ~n72 & n79;
  assign n81 = pi13 & n32;
  assign n82 = pi09 & pi13;
  assign n83 = n23 & n82;
  assign n84 = pi00 & ~n80;
  assign n85 = ~pi00 & n80;
  assign n86 = n83 & ~n85;
  assign n87 = n51 & n80;
  assign n88 = n38 & n66;
  assign n89 = n26 & n84;
  assign n90 = ~n88 & ~n89;
  assign n91 = ~n87 & n90;
  assign n92 = n81 & ~n91;
  assign n93 = ~n86 & ~n92;
  assign n94 = pi08 & ~pi10;
  assign n95 = pi09 & n40;
  assign n96 = ~pi10 & n83;
  assign n97 = pi08 & n32;
  assign n98 = ~pi09 & pi13;
  assign n99 = n97 & n98;
  assign n100 = n66 & n96;
  assign n101 = n93 & n99;
  assign n102 = ~n100 & ~n101;
  assign n103 = ~pi10 & ~n51;
  assign n104 = pi10 & n26;
  assign n105 = ~n67 & ~n68;
  assign n106 = ~pi10 & ~n105;
  assign n107 = n38 & n106;
  assign n108 = pi10 & n39;
  assign n109 = ~pi00 & ~pi08;
  assign n110 = n108 & n109;
  assign n111 = n95 & n102;
  assign n112 = pi11 & n111;
  assign n113 = ~n110 & ~n112;
  assign n114 = ~n93 & ~n113;
  assign n115 = pi09 & ~n80;
  assign n116 = ~pi00 & ~n115;
  assign n117 = ~pi11 & ~n116;
  assign n118 = pi00 & ~pi09;
  assign n119 = n80 & n118;
  assign n120 = ~n117 & ~n119;
  assign n121 = n40 & ~n120;
  assign n122 = pi08 & n102;
  assign n123 = n108 & n122;
  assign n124 = ~pi00 & ~n103;
  assign n125 = pi11 & n124;
  assign n126 = ~n123 & ~n125;
  assign n127 = ~n80 & ~n126;
  assign n128 = pi00 & pi11;
  assign n129 = ~n26 & n128;
  assign n130 = pi08 & ~n102;
  assign n131 = n39 & n130;
  assign n132 = ~n129 & ~n131;
  assign n133 = pi10 & ~n132;
  assign n134 = n37 & ~n133;
  assign n135 = n80 & ~n134;
  assign n136 = pi04 & n94;
  assign n137 = pi00 & ~pi08;
  assign n138 = n93 & n137;
  assign n139 = ~n136 & ~n138;
  assign n140 = n39 & ~n139;
  assign n141 = n95 & ~n102;
  assign n142 = pi11 & n141;
  assign n143 = ~n43 & ~n142;
  assign n144 = n93 & ~n143;
  assign n145 = ~pi00 & n104;
  assign n146 = pi11 & n145;
  assign n147 = ~n144 & ~n146;
  assign n148 = ~n140 & n147;
  assign n149 = ~n135 & n148;
  assign n150 = ~n127 & n149;
  assign n151 = ~n121 & n150;
  assign n152 = ~n114 & n151;
  assign n153 = ~n107 & n152;
  assign n154 = pi13 & ~n153;
  assign n155 = ~pi08 & pi10;
  assign n156 = ~pi11 & ~n155;
  assign n157 = pi08 & n25;
  assign n158 = ~n155 & ~n157;
  assign n159 = pi11 & n94;
  assign n160 = pi10 & pi11;
  assign n161 = ~n40 & ~n160;
  assign n162 = pi12 & n154;
  assign n163 = ~pi12 & ~n154;
  assign n164 = ~n162 & ~n163;
  assign n165 = pi13 & ~n164;
  assign n166 = pi04 & n40;
  assign n167 = ~pi09 & ~n161;
  assign n168 = ~n166 & ~n167;
  assign n169 = ~n80 & ~n168;
  assign n170 = pi04 & n23;
  assign n171 = n33 & n58;
  assign n172 = ~n170 & ~n171;
  assign n173 = n66 & ~n156;
  assign n174 = n41 & n84;
  assign n175 = ~n173 & ~n174;
  assign n176 = n172 & n175;
  assign n177 = pi09 & ~n176;
  assign n178 = n80 & ~n158;
  assign n179 = ~pi04 & n97;
  assign n180 = ~n178 & ~n179;
  assign n181 = pi11 & n67;
  assign n182 = n68 & n159;
  assign n183 = ~n181 & ~n182;
  assign n184 = n180 & n183;
  assign n185 = ~pi09 & ~n184;
  assign n186 = ~n103 & n128;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~n177 & n187;
  assign n189 = ~n169 & n188;
  assign n190 = ~pi13 & ~n189;
  assign n191 = n31 & ~n190;
  assign po0 = n165 | ~n191;
  assign n193 = ~pi12 & n154;
  assign n194 = pi10 & ~n26;
  assign n195 = ~n51 & ~n194;
  assign n196 = pi11 & ~n195;
  assign n197 = ~pi09 & n94;
  assign n198 = pi09 & ~pi10;
  assign n199 = n23 & n198;
  assign n200 = ~pi09 & n32;
  assign n201 = pi13 & n200;
  assign n202 = n57 & ~n201;
  assign n203 = ~pi01 & ~pi05;
  assign n204 = pi01 & pi05;
  assign n205 = pi01 & ~pi05;
  assign n206 = ~pi01 & pi05;
  assign n207 = ~pi08 & pi13;
  assign n208 = n69 & n207;
  assign n209 = n202 & ~n208;
  assign n210 = n204 & ~n209;
  assign n211 = n24 & n128;
  assign n212 = n32 & n206;
  assign n213 = ~n205 & ~n212;
  assign n214 = ~n68 & ~n213;
  assign n215 = n68 & n203;
  assign n216 = ~n214 & ~n215;
  assign n217 = pi09 & ~n216;
  assign n218 = ~n211 & ~n217;
  assign n219 = ~pi08 & ~n218;
  assign n220 = pi13 & n219;
  assign n221 = n62 & ~n203;
  assign n222 = ~pi01 & n65;
  assign n223 = ~pi05 & ~n50;
  assign n224 = ~n222 & ~n223;
  assign n225 = ~n221 & n224;
  assign n226 = ~n220 & n225;
  assign n227 = ~n210 & n226;
  assign n228 = n80 & n227;
  assign n229 = ~pi01 & n227;
  assign n230 = n83 & ~n229;
  assign n231 = n51 & n227;
  assign n232 = pi09 & ~n227;
  assign n233 = pi05 & ~pi09;
  assign n234 = ~n232 & ~n233;
  assign n235 = pi08 & ~n234;
  assign n236 = pi01 & n235;
  assign n237 = ~n231 & ~n236;
  assign n238 = n81 & ~n237;
  assign n239 = ~n230 & ~n238;
  assign n240 = pi00 & ~n93;
  assign n241 = n239 & n240;
  assign n242 = ~n239 & ~n240;
  assign n243 = ~n241 & ~n242;
  assign n244 = ~n80 & ~n102;
  assign n245 = ~pi00 & ~pi01;
  assign n246 = n93 & n239;
  assign n247 = n96 & n204;
  assign n248 = n99 & n239;
  assign n249 = ~n247 & ~n248;
  assign n250 = ~n93 & ~n102;
  assign n251 = ~pi10 & n51;
  assign n252 = ~n196 & ~n251;
  assign n253 = n25 & ~n26;
  assign n254 = ~pi11 & n42;
  assign n255 = ~n35 & ~n254;
  assign n256 = n84 & n227;
  assign n257 = ~n84 & ~n227;
  assign n258 = ~n256 & ~n257;
  assign n259 = n196 & ~n258;
  assign n260 = n155 & ~n243;
  assign n261 = n39 & n260;
  assign n262 = ~n259 & ~n261;
  assign n263 = ~pi01 & ~n262;
  assign n264 = n244 & ~n249;
  assign n265 = ~n244 & n249;
  assign n266 = ~n264 & ~n265;
  assign n267 = ~n227 & ~n266;
  assign n268 = ~n244 & ~n249;
  assign n269 = n244 & n249;
  assign n270 = ~n268 & ~n269;
  assign n271 = n227 & ~n270;
  assign n272 = ~n267 & ~n271;
  assign n273 = n41 & ~n272;
  assign n274 = pi05 & n94;
  assign n275 = ~pi08 & n243;
  assign n276 = pi01 & n275;
  assign n277 = ~n274 & ~n276;
  assign n278 = ~n273 & n277;
  assign n279 = n39 & ~n278;
  assign n280 = n104 & n245;
  assign n281 = n66 & n203;
  assign n282 = n197 & n281;
  assign n283 = ~n280 & ~n282;
  assign n284 = pi11 & ~n283;
  assign n285 = ~n249 & n250;
  assign n286 = n249 & ~n250;
  assign n287 = ~n285 & ~n286;
  assign n288 = ~n239 & ~n287;
  assign n289 = n249 & n250;
  assign n290 = ~n249 & ~n250;
  assign n291 = ~n289 & ~n290;
  assign n292 = n239 & ~n291;
  assign n293 = ~n288 & ~n292;
  assign n294 = n199 & ~n293;
  assign n295 = n84 & ~n227;
  assign n296 = ~n84 & n227;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n252 & ~n297;
  assign n299 = n104 & n128;
  assign n300 = ~pi05 & ~n66;
  assign n301 = n197 & n300;
  assign n302 = ~n299 & ~n301;
  assign n303 = ~n253 & n302;
  assign n304 = ~n298 & n303;
  assign n305 = pi01 & ~n304;
  assign n306 = ~n93 & ~n239;
  assign n307 = ~n246 & ~n306;
  assign n308 = n104 & ~n307;
  assign n309 = n95 & ~n227;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~pi11 & ~n310;
  assign n312 = ~n66 & n206;
  assign n313 = n66 & n204;
  assign n314 = ~n312 & ~n313;
  assign n315 = n197 & ~n314;
  assign n316 = ~n37 & n228;
  assign n317 = ~n80 & ~n255;
  assign n318 = ~n227 & n317;
  assign n319 = ~n316 & ~n318;
  assign n320 = ~n315 & n319;
  assign n321 = ~n311 & n320;
  assign n322 = ~n305 & n321;
  assign n323 = ~n294 & n322;
  assign n324 = ~n284 & n323;
  assign n325 = ~n279 & n324;
  assign n326 = ~n263 & n325;
  assign n327 = pi13 & ~n326;
  assign n328 = ~n193 & n327;
  assign n329 = n193 & ~n327;
  assign n330 = ~n328 & ~n329;
  assign n331 = pi13 & ~n330;
  assign n332 = pi11 & ~n103;
  assign n333 = pi09 & n41;
  assign n334 = ~n227 & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = pi01 & ~n335;
  assign n337 = pi05 & n40;
  assign n338 = ~n167 & ~n337;
  assign n339 = ~n227 & ~n338;
  assign n340 = pi05 & n23;
  assign n341 = ~n156 & n204;
  assign n342 = n33 & n203;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~n340 & n343;
  assign n345 = pi09 & ~n344;
  assign n346 = pi11 & n205;
  assign n347 = n159 & n206;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n158 & n227;
  assign n350 = ~pi05 & n97;
  assign n351 = ~n349 & ~n350;
  assign n352 = n348 & n351;
  assign n353 = ~pi09 & ~n352;
  assign n354 = ~n345 & ~n353;
  assign n355 = ~n339 & n354;
  assign n356 = ~n336 & n355;
  assign n357 = ~pi13 & ~n356;
  assign n358 = n31 & ~n357;
  assign po1 = n331 | ~n358;
  assign n360 = n193 & n327;
  assign n361 = ~pi02 & ~pi06;
  assign n362 = pi02 & pi06;
  assign n363 = n68 & ~n205;
  assign n364 = ~n206 & ~n363;
  assign n365 = n32 & ~n364;
  assign n366 = pi06 & n365;
  assign n367 = pi09 & n364;
  assign n368 = ~pi06 & n367;
  assign n369 = ~n366 & ~n368;
  assign n370 = pi02 & ~n369;
  assign n371 = ~pi06 & ~n364;
  assign n372 = n32 & n364;
  assign n373 = pi06 & n372;
  assign n374 = ~n371 & ~n373;
  assign n375 = pi09 & ~n374;
  assign n376 = ~pi02 & n375;
  assign n377 = pi01 & pi11;
  assign n378 = n24 & n377;
  assign n379 = ~n376 & ~n378;
  assign n380 = ~n370 & n379;
  assign n381 = ~pi08 & ~n380;
  assign n382 = pi13 & n381;
  assign n383 = ~n202 & n362;
  assign n384 = ~pi06 & ~n50;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~pi02 & n65;
  assign n387 = n62 & ~n361;
  assign n388 = ~n386 & ~n387;
  assign n389 = n385 & n388;
  assign n390 = ~n382 & n389;
  assign n391 = n66 & ~n203;
  assign n392 = ~n204 & ~n391;
  assign n393 = n228 & n390;
  assign n394 = ~pi02 & n390;
  assign n395 = n83 & ~n394;
  assign n396 = n51 & n390;
  assign n397 = pi09 & ~n390;
  assign n398 = pi06 & ~pi09;
  assign n399 = ~n397 & ~n398;
  assign n400 = pi08 & ~n399;
  assign n401 = pi02 & n400;
  assign n402 = ~n396 & ~n401;
  assign n403 = n81 & ~n402;
  assign n404 = ~n395 & ~n403;
  assign n405 = n96 & n362;
  assign n406 = n99 & n404;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~n239 & ~n286;
  assign n409 = ~n285 & ~n408;
  assign n410 = n390 & n407;
  assign n411 = ~n390 & ~n407;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n227 & ~n265;
  assign n414 = ~n264 & ~n413;
  assign n415 = ~pi01 & ~n240;
  assign n416 = ~n239 & ~n415;
  assign n417 = pi01 & n240;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n404 & n418;
  assign n420 = n404 & ~n418;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~pi01 & ~n84;
  assign n423 = ~n227 & ~n422;
  assign n424 = pi01 & n84;
  assign n425 = ~n423 & ~n424;
  assign n426 = pi02 & pi11;
  assign n427 = ~pi02 & n245;
  assign n428 = n246 & n404;
  assign n429 = ~n252 & n425;
  assign n430 = pi02 & n429;
  assign n431 = n196 & ~n425;
  assign n432 = ~pi02 & n431;
  assign n433 = ~n430 & ~n432;
  assign n434 = n390 & ~n433;
  assign n435 = pi11 & n361;
  assign n436 = ~n362 & ~n435;
  assign n437 = ~n392 & ~n436;
  assign n438 = ~pi02 & pi06;
  assign n439 = pi02 & ~pi06;
  assign n440 = ~n438 & ~n439;
  assign n441 = n392 & ~n440;
  assign n442 = ~n437 & ~n441;
  assign n443 = n197 & ~n442;
  assign n444 = n196 & n425;
  assign n445 = ~n390 & n444;
  assign n446 = n155 & ~n421;
  assign n447 = n39 & n446;
  assign n448 = ~n445 & ~n447;
  assign n449 = ~pi02 & ~n448;
  assign n450 = ~n404 & ~n409;
  assign n451 = n404 & n409;
  assign n452 = ~n450 & ~n451;
  assign n453 = ~n407 & ~n452;
  assign n454 = ~n404 & n409;
  assign n455 = n404 & ~n409;
  assign n456 = ~n454 & ~n455;
  assign n457 = n407 & ~n456;
  assign n458 = ~n453 & ~n457;
  assign n459 = n199 & ~n458;
  assign n460 = ~n412 & ~n414;
  assign n461 = n412 & n414;
  assign n462 = ~n460 & ~n461;
  assign n463 = n41 & ~n462;
  assign n464 = pi06 & n94;
  assign n465 = ~pi08 & n421;
  assign n466 = pi02 & n465;
  assign n467 = ~n464 & ~n466;
  assign n468 = ~n463 & n467;
  assign n469 = n39 & ~n468;
  assign n470 = ~n252 & ~n425;
  assign n471 = ~n390 & n470;
  assign n472 = ~n253 & ~n471;
  assign n473 = pi02 & ~n472;
  assign n474 = ~pi11 & n95;
  assign n475 = ~n228 & ~n255;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n390 & ~n476;
  assign n478 = ~n246 & ~n404;
  assign n479 = ~n428 & ~n478;
  assign n480 = ~pi11 & ~n479;
  assign n481 = pi11 & n427;
  assign n482 = ~n245 & n426;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n480 & n483;
  assign n485 = n104 & ~n484;
  assign n486 = ~n37 & n393;
  assign n487 = ~n485 & ~n486;
  assign n488 = ~n477 & n487;
  assign n489 = ~n473 & n488;
  assign n490 = ~n469 & n489;
  assign n491 = ~n459 & n490;
  assign n492 = ~n449 & n491;
  assign n493 = ~n443 & n492;
  assign n494 = ~n434 & n493;
  assign n495 = pi13 & ~n494;
  assign n496 = ~n360 & n495;
  assign n497 = n360 & ~n495;
  assign n498 = ~n496 & ~n497;
  assign n499 = pi13 & ~n498;
  assign n500 = ~pi06 & ~pi09;
  assign n501 = n103 & ~n500;
  assign n502 = n426 & ~n501;
  assign n503 = pi06 & n40;
  assign n504 = pi02 & n41;
  assign n505 = pi09 & n504;
  assign n506 = ~n167 & ~n505;
  assign n507 = ~n503 & n506;
  assign n508 = ~n390 & ~n507;
  assign n509 = pi09 & n23;
  assign n510 = ~pi02 & n159;
  assign n511 = ~pi09 & n510;
  assign n512 = ~n509 & ~n511;
  assign n513 = pi06 & ~n512;
  assign n514 = ~n156 & n362;
  assign n515 = n33 & n361;
  assign n516 = ~n514 & ~n515;
  assign n517 = pi09 & ~n516;
  assign n518 = ~n158 & n390;
  assign n519 = ~pi06 & n97;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~pi09 & ~n520;
  assign n522 = ~n517 & ~n521;
  assign n523 = ~n513 & n522;
  assign n524 = ~n508 & n523;
  assign n525 = ~n502 & n524;
  assign n526 = ~pi13 & ~n525;
  assign n527 = n31 & ~n526;
  assign po2 = n499 | ~n527;
  assign n529 = n360 & n495;
  assign n530 = ~pi03 & ~pi07;
  assign po5 = pi03 & pi07;
  assign n532 = n364 & ~n438;
  assign n533 = ~n439 & ~n532;
  assign n534 = pi09 & ~n533;
  assign n535 = pi03 & n534;
  assign n536 = n207 & n535;
  assign n537 = n50 & ~n536;
  assign n538 = ~pi07 & ~n537;
  assign n539 = n32 & n533;
  assign n540 = pi13 & n539;
  assign n541 = ~n200 & ~n540;
  assign n542 = po5 & ~n541;
  assign n543 = ~pi10 & ~n63;
  assign n544 = ~pi13 & n543;
  assign n545 = pi07 & pi13;
  assign n546 = pi09 & n32;
  assign n547 = ~n533 & n546;
  assign n548 = n545 & n547;
  assign n549 = ~n544 & ~n548;
  assign n550 = ~pi03 & ~n549;
  assign n551 = n24 & n426;
  assign n552 = pi09 & n533;
  assign n553 = n530 & n552;
  assign n554 = ~n551 & ~n553;
  assign n555 = pi13 & ~n554;
  assign n556 = ~n550 & ~n555;
  assign n557 = ~n542 & n556;
  assign n558 = ~pi08 & ~n557;
  assign n559 = ~n54 & ~n200;
  assign n560 = pi13 & ~n559;
  assign n561 = po5 & n560;
  assign n562 = n62 & ~n530;
  assign n563 = ~n561 & ~n562;
  assign n564 = ~n558 & n563;
  assign n565 = ~n538 & n564;
  assign n566 = n393 & n565;
  assign n567 = pi03 & pi11;
  assign n568 = pi03 & ~n565;
  assign n569 = ~pi03 & n565;
  assign n570 = n83 & ~n569;
  assign n571 = n51 & n565;
  assign n572 = n26 & n568;
  assign n573 = n38 & po5;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~n571 & n574;
  assign n576 = n81 & ~n575;
  assign n577 = ~n570 & ~n576;
  assign n578 = n96 & po5;
  assign n579 = n99 & n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = n407 & n409;
  assign n582 = ~n404 & ~n581;
  assign n583 = ~n407 & ~n409;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~pi02 & n425;
  assign n586 = ~n390 & ~n585;
  assign n587 = pi02 & ~n425;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~n565 & n588;
  assign n590 = n565 & ~n588;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n361 & ~n392;
  assign n593 = ~n362 & ~n592;
  assign n594 = ~pi02 & n418;
  assign n595 = ~n404 & ~n594;
  assign n596 = pi02 & ~n418;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n565 & n580;
  assign n599 = n565 & ~n580;
  assign n600 = ~n598 & ~n599;
  assign n601 = n407 & n414;
  assign n602 = ~n390 & ~n601;
  assign n603 = ~n407 & ~n414;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~n255 & ~n393;
  assign n606 = ~n474 & ~n605;
  assign n607 = ~n565 & ~n606;
  assign n608 = n577 & ~n597;
  assign n609 = ~n577 & n597;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~pi08 & ~n610;
  assign n612 = ~pi03 & n611;
  assign n613 = n600 & ~n604;
  assign n614 = ~n600 & n604;
  assign n615 = ~n613 & ~n614;
  assign n616 = pi08 & ~n615;
  assign n617 = ~n612 & ~n616;
  assign n618 = n200 & ~n617;
  assign n619 = ~n577 & ~n584;
  assign n620 = n577 & n584;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n580 & ~n621;
  assign n623 = ~n577 & n584;
  assign n624 = n577 & ~n584;
  assign n625 = ~n623 & ~n624;
  assign n626 = n580 & ~n625;
  assign n627 = ~n622 & ~n626;
  assign n628 = n95 & ~n627;
  assign n629 = ~pi03 & n427;
  assign n630 = n104 & n629;
  assign n631 = n530 & ~n593;
  assign n632 = n197 & n631;
  assign n633 = ~n630 & ~n632;
  assign n634 = ~n628 & n633;
  assign n635 = pi11 & ~n634;
  assign n636 = n196 & ~n591;
  assign n637 = pi07 & n593;
  assign n638 = n197 & n637;
  assign n639 = ~n636 & ~n638;
  assign n640 = ~pi03 & ~n639;
  assign n641 = n428 & n577;
  assign n642 = ~n428 & ~n577;
  assign n643 = ~n641 & ~n642;
  assign n644 = n104 & ~n643;
  assign n645 = ~n577 & ~n597;
  assign n646 = n577 & n597;
  assign n647 = ~n645 & ~n646;
  assign n648 = n51 & ~n647;
  assign n649 = pi03 & n648;
  assign n650 = pi07 & n197;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n644 & n651;
  assign n653 = ~pi11 & ~n652;
  assign n654 = ~pi07 & n593;
  assign n655 = pi03 & n654;
  assign n656 = po5 & ~n593;
  assign n657 = ~n655 & ~n656;
  assign n658 = n197 & ~n657;
  assign n659 = ~n252 & n591;
  assign n660 = ~n253 & ~n659;
  assign n661 = pi03 & ~n660;
  assign n662 = ~n37 & n566;
  assign n663 = ~n427 & n567;
  assign n664 = n104 & n663;
  assign n665 = ~n662 & ~n664;
  assign n666 = ~n661 & n665;
  assign n667 = ~n658 & n666;
  assign n668 = ~n653 & n667;
  assign n669 = ~n640 & n668;
  assign n670 = ~n635 & n669;
  assign n671 = ~n618 & n670;
  assign n672 = ~n607 & n671;
  assign n673 = pi13 & ~n672;
  assign n674 = ~n529 & n673;
  assign n675 = n529 & ~n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = pi13 & ~n676;
  assign n678 = ~pi07 & ~pi09;
  assign n679 = n103 & ~n678;
  assign n680 = n567 & ~n679;
  assign n681 = pi07 & n40;
  assign n682 = ~n167 & ~n681;
  assign n683 = ~n565 & ~n682;
  assign n684 = ~pi03 & n159;
  assign n685 = ~pi09 & n684;
  assign n686 = ~n509 & ~n685;
  assign n687 = pi07 & ~n686;
  assign n688 = ~n158 & n565;
  assign n689 = ~pi07 & n97;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~pi09 & ~n690;
  assign n692 = n41 & n568;
  assign n693 = n33 & n530;
  assign n694 = ~n156 & po5;
  assign n695 = ~n693 & ~n694;
  assign n696 = ~n692 & n695;
  assign n697 = pi09 & ~n696;
  assign n698 = ~n691 & ~n697;
  assign n699 = ~n687 & n698;
  assign n700 = ~n683 & n699;
  assign n701 = ~n680 & n700;
  assign n702 = ~pi13 & ~n701;
  assign n703 = n31 & ~n702;
  assign po3 = n677 | ~n703;
  assign po4 = n530 | po5;
  assign n706 = pi10 & n42;
  assign n707 = ~pi11 & n706;
  assign n708 = ~n34 & ~n707;
  assign n709 = n566 & ~n708;
  assign n710 = n580 & n584;
  assign n711 = ~n577 & ~n710;
  assign n712 = ~n580 & ~n584;
  assign n713 = ~n711 & ~n712;
  assign n714 = n95 & ~n713;
  assign n715 = ~n530 & ~n593;
  assign n716 = ~po5 & ~n715;
  assign n717 = n197 & ~n716;
  assign n718 = ~n569 & ~n588;
  assign n719 = ~n568 & ~n718;
  assign n720 = ~n195 & ~n719;
  assign n721 = ~n630 & ~n720;
  assign n722 = ~n717 & n721;
  assign n723 = ~n714 & n722;
  assign n724 = pi11 & ~n723;
  assign n725 = ~pi03 & n597;
  assign n726 = ~n577 & ~n725;
  assign n727 = pi03 & ~n597;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~pi08 & ~n728;
  assign n730 = n565 & n604;
  assign n731 = ~n580 & ~n730;
  assign n732 = ~n565 & ~n604;
  assign n733 = ~n731 & ~n732;
  assign n734 = pi08 & ~n733;
  assign n735 = ~n729 & ~n734;
  assign n736 = n24 & ~n735;
  assign n737 = n26 & n641;
  assign n738 = ~n34 & ~n737;
  assign n739 = ~n736 & n738;
  assign n740 = ~pi11 & ~n739;
  assign n741 = n529 & n673;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~n724 & n742;
  assign n744 = ~n709 & n743;
  assign po6 = pi13 & ~n744;
  assign n746 = n245 & n362;
  assign n747 = ~pi06 & n427;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~pi05 & ~n748;
  assign n750 = ~pi04 & n749;
  assign n751 = ~n361 & ~n362;
  assign n752 = ~n58 & ~n66;
  assign n753 = n204 & ~n752;
  assign n754 = ~n281 & ~n753;
  assign n755 = ~n751 & ~n754;
  assign n756 = ~n750 & ~n755;
  assign po7 = po4 & ~n756;
endmodule



module top (
            a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63, 
            asquared_0, asquared_1, asquared_2, asquared_3, asquared_4, asquared_5, asquared_6, asquared_7, asquared_8, asquared_9, asquared_10, asquared_11, asquared_12, asquared_13, asquared_14, asquared_15, asquared_16, asquared_17, asquared_18, asquared_19, asquared_20, asquared_21, asquared_22, asquared_23, asquared_24, asquared_25, asquared_26, asquared_27, asquared_28, asquared_29, asquared_30, asquared_31, asquared_32, asquared_33, asquared_34, asquared_35, asquared_36, asquared_37, asquared_38, asquared_39, asquared_40, asquared_41, asquared_42, asquared_43, asquared_44, asquared_45, asquared_46, asquared_47, asquared_48, asquared_49, asquared_50, asquared_51, asquared_52, asquared_53, asquared_54, asquared_55, asquared_56, asquared_57, asquared_58, asquared_59, asquared_60, asquared_61, asquared_62, asquared_63, asquared_64, asquared_65, asquared_66, asquared_67, asquared_68, asquared_69, asquared_70, asquared_71, asquared_72, asquared_73, asquared_74, asquared_75, asquared_76, asquared_77, asquared_78, asquared_79, asquared_80, asquared_81, asquared_82, asquared_83, asquared_84, asquared_85, asquared_86, asquared_87, asquared_88, asquared_89, asquared_90, asquared_91, asquared_92, asquared_93, asquared_94, asquared_95, asquared_96, asquared_97, asquared_98, asquared_99, asquared_100, asquared_101, asquared_102, asquared_103, asquared_104, asquared_105, asquared_106, asquared_107, asquared_108, asquared_109, asquared_110, asquared_111, asquared_112, asquared_113, asquared_114, asquared_115, asquared_116, asquared_117, asquared_118, asquared_119, asquared_120, asquared_121, asquared_122, asquared_123, asquared_124, asquared_125, asquared_126, asquared_127);
input a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, a_16, a_17, a_18, a_19, a_20, a_21, a_22, a_23, a_24, a_25, a_26, a_27, a_28, a_29, a_30, a_31, a_32, a_33, a_34, a_35, a_36, a_37, a_38, a_39, a_40, a_41, a_42, a_43, a_44, a_45, a_46, a_47, a_48, a_49, a_50, a_51, a_52, a_53, a_54, a_55, a_56, a_57, a_58, a_59, a_60, a_61, a_62, a_63;
output asquared_0, asquared_1, asquared_2, asquared_3, asquared_4, asquared_5, asquared_6, asquared_7, asquared_8, asquared_9, asquared_10, asquared_11, asquared_12, asquared_13, asquared_14, asquared_15, asquared_16, asquared_17, asquared_18, asquared_19, asquared_20, asquared_21, asquared_22, asquared_23, asquared_24, asquared_25, asquared_26, asquared_27, asquared_28, asquared_29, asquared_30, asquared_31, asquared_32, asquared_33, asquared_34, asquared_35, asquared_36, asquared_37, asquared_38, asquared_39, asquared_40, asquared_41, asquared_42, asquared_43, asquared_44, asquared_45, asquared_46, asquared_47, asquared_48, asquared_49, asquared_50, asquared_51, asquared_52, asquared_53, asquared_54, asquared_55, asquared_56, asquared_57, asquared_58, asquared_59, asquared_60, asquared_61, asquared_62, asquared_63, asquared_64, asquared_65, asquared_66, asquared_67, asquared_68, asquared_69, asquared_70, asquared_71, asquared_72, asquared_73, asquared_74, asquared_75, asquared_76, asquared_77, asquared_78, asquared_79, asquared_80, asquared_81, asquared_82, asquared_83, asquared_84, asquared_85, asquared_86, asquared_87, asquared_88, asquared_89, asquared_90, asquared_91, asquared_92, asquared_93, asquared_94, asquared_95, asquared_96, asquared_97, asquared_98, asquared_99, asquared_100, asquared_101, asquared_102, asquared_103, asquared_104, asquared_105, asquared_106, asquared_107, asquared_108, asquared_109, asquared_110, asquared_111, asquared_112, asquared_113, asquared_114, asquared_115, asquared_116, asquared_117, asquared_118, asquared_119, asquared_120, asquared_121, asquared_122, asquared_123, asquared_124, asquared_125, asquared_126, asquared_127;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200;
assign w0 = ~w14332 & w9733;
assign w1 = a_16 & a_35;
assign w2 = (~w14263 & ~w12080) | (~w14263 & w12872) | (~w12080 & w12872);
assign w3 = a_19 & a_26;
assign w4 = ~w5186 & ~w7328;
assign w5 = ~w16252 & ~w2056;
assign w6 = ~w7756 & ~w14219;
assign w7 = a_31 & ~w13854;
assign w8 = a_22 & a_35;
assign w9 = ~w14215 & ~w2599;
assign w10 = (~w12798 & ~w15708) | (~w12798 & w3503) | (~w15708 & w3503);
assign w11 = ~w6331 & ~w11160;
assign w12 = w11789 & ~w7946;
assign w13 = ~w5010 & ~w1401;
assign w14 = ~w16795 & ~w5638;
assign w15 = w13821 & w12747;
assign w16 = (w17995 & w13082) | (w17995 & w14269) | (w13082 & w14269);
assign w17 = a_29 & a_60;
assign w18 = ~w4227 & ~w14653;
assign w19 = w2227 & ~w15499;
assign w20 = (~w3728 & ~w5219) | (~w3728 & w15773) | (~w5219 & w15773);
assign w21 = w422 & w1650;
assign w22 = w6680 & ~w19142;
assign w23 = w11991 & w16938;
assign w24 = ~w1993 & ~w6068;
assign w25 = ~w1387 & ~w828;
assign w26 = ~w6076 & w4821;
assign w27 = ~w10839 & ~w14606;
assign w28 = ~w1245 & ~w15330;
assign w29 = w8217 & w13272;
assign w30 = ~w6043 & w14593;
assign w31 = (~w6613 & ~w8367) | (~w6613 & w8593) | (~w8367 & w8593);
assign w32 = ~w3602 & w15708;
assign w33 = ~w11652 & ~w18462;
assign w34 = ~w11874 & ~w7080;
assign w35 = ~w7202 & ~w11259;
assign w36 = ~w4398 & ~w7963;
assign w37 = w8859 & w5885;
assign w38 = ~w17081 & w2865;
assign w39 = ~w9014 & ~w10222;
assign w40 = (w1596 & w7610) | (w1596 & w15671) | (w7610 & w15671);
assign w41 = (~w4589 & ~w18442) | (~w4589 & w5611) | (~w18442 & w5611);
assign w42 = ~w7248 & ~w16034;
assign w43 = ~w4065 & ~w16081;
assign w44 = w13686 & w983;
assign w45 = a_1 & a_13;
assign w46 = ~w2154 & w2093;
assign w47 = ~w15515 & ~w7603;
assign w48 = w11939 & ~w7921;
assign w49 = ~w14126 & ~w1326;
assign w50 = w11687 & w617;
assign w51 = ~w5713 & ~w6718;
assign w52 = ~w12027 & ~w9539;
assign w53 = ~w10273 & ~w1011;
assign w54 = w13082 & w1290;
assign w55 = ~w3659 & ~w3516;
assign w56 = ~w4503 & ~w17545;
assign w57 = ~w3152 & ~w7510;
assign w58 = ~w6249 & ~w14233;
assign w59 = ~w16628 & ~w17879;
assign w60 = a_35 & a_51;
assign w61 = ~w11491 & ~w9582;
assign w62 = ~w12957 & ~w5902;
assign w63 = ~w14329 & w6262;
assign w64 = w4143 & ~w16397;
assign w65 = w9027 & w7556;
assign w66 = ~w3536 & ~w10980;
assign w67 = ~w17498 & ~w12188;
assign w68 = (~w6894 & w1326) | (~w6894 & w4783) | (w1326 & w4783);
assign w69 = ~w4578 & ~w9199;
assign w70 = ~w3596 & ~w5997;
assign w71 = ~w4220 & ~w8224;
assign w72 = ~w16367 & ~w2122;
assign w73 = ~w17858 & ~w15402;
assign w74 = w7425 & ~w498;
assign w75 = w18753 & ~w2109;
assign w76 = ~w15332 & w9784;
assign w77 = ~w9713 & ~w4927;
assign w78 = ~w2946 & ~w12084;
assign w79 = ~w14965 & w12970;
assign w80 = ~w18493 & ~w19051;
assign w81 = w3672 & ~w5139;
assign w82 = w3585 & ~w18405;
assign w83 = (~w1948 & ~w12899) | (~w1948 & w15600) | (~w12899 & w15600);
assign w84 = a_25 & a_26;
assign w85 = w9926 & w8073;
assign w86 = ~w5700 & ~w5251;
assign w87 = w393 & w9760;
assign w88 = ~w9200 & ~w377;
assign w89 = ~w3082 & ~w5495;
assign w90 = ~w16576 & ~w16680;
assign w91 = a_4 & a_44;
assign w92 = ~w16612 & ~w15974;
assign w93 = ~w773 & ~w12470;
assign w94 = ~w11102 & ~w3091;
assign w95 = ~w634 & ~w6029;
assign w96 = a_11 & a_56;
assign w97 = w12229 & ~w3204;
assign w98 = ~w5058 & ~w17183;
assign w99 = a_2 & a_3;
assign w100 = ~w7365 & ~w10398;
assign w101 = w4556 & ~w12899;
assign w102 = ~w12334 & w12992;
assign w103 = w13248 & ~w16270;
assign w104 = ~w5477 & ~w3538;
assign w105 = ~w8859 & ~w5885;
assign w106 = ~w17107 & ~w12822;
assign w107 = ~w12183 & ~w5536;
assign w108 = ~w12234 & ~w8872;
assign w109 = a_17 & a_55;
assign w110 = ~w13883 & ~w6204;
assign w111 = ~w18286 & ~w9350;
assign w112 = ~w5224 & ~w12079;
assign w113 = w6896 & w4552;
assign w114 = ~w14383 & w6354;
assign w115 = a_9 & a_33;
assign w116 = ~w11353 & ~w10766;
assign w117 = w12600 & ~w8144;
assign w118 = ~w7456 & w11592;
assign w119 = a_22 & a_50;
assign w120 = ~w14129 & ~w7798;
assign w121 = (w5495 & w8661) | (w5495 & w17384) | (w8661 & w17384);
assign w122 = w15877 & w17376;
assign w123 = ~w14297 & w4303;
assign w124 = ~w16835 & ~w10715;
assign w125 = ~w6908 & ~w16142;
assign w126 = w12274 & w3658;
assign w127 = (~w13797 & ~w15808) | (~w13797 & w10380) | (~w15808 & w10380);
assign w128 = ~w14409 & ~w2470;
assign w129 = ~w17243 & ~w17090;
assign w130 = ~w6171 & w11518;
assign w131 = (w4528 & w16404) | (w4528 & w16844) | (w16404 & w16844);
assign w132 = ~w13932 & ~w6909;
assign w133 = w4993 & ~w6886;
assign w134 = a_17 & a_56;
assign w135 = w3913 & ~w19133;
assign w136 = a_14 & a_62;
assign w137 = ~w1656 & ~w12883;
assign w138 = ~w7266 & ~w3031;
assign w139 = ~w10099 & ~w3621;
assign w140 = ~w4170 & w12510;
assign w141 = w10033 & w3734;
assign w142 = ~w15838 & ~w7477;
assign w143 = (~w11004 & ~w3104) | (~w11004 & w13122) | (~w3104 & w13122);
assign w144 = ~w651 & ~w14265;
assign w145 = ~w13001 & ~w13519;
assign w146 = (w9902 & w7129) | (w9902 & w16710) | (w7129 & w16710);
assign w147 = ~w11990 & ~w17484;
assign w148 = ~w6000 & w2570;
assign w149 = a_16 & w7241;
assign w150 = ~w14085 & ~w12255;
assign w151 = (~w10883 & ~w17634) | (~w10883 & w3768) | (~w17634 & w3768);
assign w152 = ~w9799 & w7612;
assign w153 = ~w18902 & ~w2224;
assign w154 = (w3182 & w7735) | (w3182 & w2229) | (w7735 & w2229);
assign w155 = w4342 & ~w14919;
assign w156 = ~w17413 & w10500;
assign w157 = a_33 & a_35;
assign w158 = ~w18485 & w8915;
assign w159 = (w5296 & w5978) | (w5296 & w14180) | (w5978 & w14180);
assign w160 = ~w9039 & w5599;
assign w161 = ~w5203 & w1823;
assign w162 = ~w4279 & w5883;
assign w163 = ~w3043 & ~w5035;
assign w164 = ~w12880 & ~w1591;
assign w165 = ~w15982 & ~w9241;
assign w166 = ~w8193 & ~w16880;
assign w167 = ~w17389 & ~w17675;
assign w168 = w275 & ~w2991;
assign w169 = ~w12233 & ~w6170;
assign w170 = w6116 & ~w2794;
assign w171 = w3360 & ~w11533;
assign w172 = ~w8304 & w1418;
assign w173 = ~w1389 & ~w9964;
assign w174 = w6738 & ~w2014;
assign w175 = ~w15575 & ~w16072;
assign w176 = w3119 & ~w801;
assign w177 = w3915 & ~w7255;
assign w178 = ~w14833 & ~w6256;
assign w179 = w4436 & ~w11263;
assign w180 = w15048 & ~w9875;
assign w181 = w2025 & ~w18505;
assign w182 = a_0 & a_35;
assign w183 = ~w17787 & ~w10467;
assign w184 = ~w5881 & ~w17111;
assign w185 = ~w6891 & ~w3991;
assign w186 = ~w17743 & ~w5519;
assign w187 = ~w5221 & ~w4157;
assign w188 = w14993 & w1320;
assign w189 = ~w15583 & w14321;
assign w190 = a_10 & a_43;
assign w191 = ~w4373 & ~w13512;
assign w192 = ~w600 & ~w11425;
assign w193 = w13557 & w17305;
assign w194 = (~w16180 & ~w245) | (~w16180 & w9572) | (~w245 & w9572);
assign w195 = w1962 & ~w3932;
assign w196 = ~w3655 & ~w12172;
assign w197 = ~w11026 & ~w219;
assign w198 = w4339 & w11149;
assign w199 = ~w9679 & ~w11989;
assign w200 = w4770 & w2120;
assign w201 = a_12 & a_26;
assign w202 = ~w11008 & w11679;
assign w203 = a_20 & a_61;
assign w204 = ~w1700 & w17118;
assign w205 = ~w16722 & ~w12240;
assign w206 = w1753 & w2342;
assign w207 = ~w11939 & ~w18973;
assign w208 = ~w4117 & ~w2756;
assign w209 = a_15 & a_25;
assign w210 = ~w4947 & ~w16846;
assign w211 = w4478 & w5132;
assign w212 = w6669 & w16736;
assign w213 = w12430 & ~w14353;
assign w214 = ~w14336 & ~w11878;
assign w215 = ~w14341 & ~w9865;
assign w216 = w4478 & ~w12825;
assign w217 = w15899 & w11246;
assign w218 = (~w769 & ~w9635) | (~w769 & w12093) | (~w9635 & w12093);
assign w219 = w18872 & w9610;
assign w220 = ~w16551 & ~w5237;
assign w221 = ~w9381 & ~w9689;
assign w222 = w13461 & ~w12647;
assign w223 = w534 & ~w17968;
assign w224 = w13082 & ~w15163;
assign w225 = w15147 & w18617;
assign w226 = ~w14323 & w1134;
assign w227 = ~w9667 & ~w5047;
assign w228 = ~w9970 & ~w11886;
assign w229 = ~w5298 & ~w7224;
assign w230 = ~w13749 & ~w16227;
assign w231 = ~w17953 & ~w14371;
assign w232 = ~w10647 & w17279;
assign w233 = ~w1513 & ~w759;
assign w234 = ~w5420 & ~w14022;
assign w235 = ~w13198 & w6054;
assign w236 = ~w7681 & ~w3155;
assign w237 = ~w6079 & ~w6429;
assign w238 = ~w15619 & w17412;
assign w239 = w5401 & w9557;
assign w240 = (~w13938 & ~w5949) | (~w13938 & w9462) | (~w5949 & w9462);
assign w241 = w10888 & ~w14017;
assign w242 = ~w13635 & ~w8108;
assign w243 = ~w1000 & ~w1325;
assign w244 = ~w10158 & ~w17931;
assign w245 = ~w9078 & ~w16180;
assign w246 = a_17 & a_63;
assign w247 = (w4547 & w2769) | (w4547 & w7420) | (w2769 & w7420);
assign w248 = ~w11109 & ~w17631;
assign w249 = ~w13527 & ~w365;
assign w250 = a_9 & a_11;
assign w251 = ~w12171 & ~w4795;
assign w252 = (~w4006 & ~w11161) | (~w4006 & w19105) | (~w11161 & w19105);
assign w253 = a_42 & a_52;
assign w254 = w3586 & ~w3748;
assign w255 = ~a_0 & a_1;
assign w256 = w12864 & ~w5958;
assign w257 = ~w1467 & ~w14640;
assign w258 = (~w15080 & w11488) | (~w15080 & w2262) | (w11488 & w2262);
assign w259 = a_20 & a_49;
assign w260 = ~w16820 & ~w9952;
assign w261 = w935 & w6406;
assign w262 = ~w17170 & ~w6242;
assign w263 = (w1225 & w5939) | (w1225 & ~w11396) | (w5939 & ~w11396);
assign w264 = ~w10010 & w6526;
assign w265 = w2885 & w18337;
assign w266 = ~w2948 & ~w9043;
assign w267 = ~w9708 & ~w2867;
assign w268 = a_46 & a_50;
assign w269 = a_30 & a_35;
assign w270 = ~w12815 & ~w18119;
assign w271 = ~w3794 & w17385;
assign w272 = w2048 & ~w16288;
assign w273 = ~w4034 & ~w17077;
assign w274 = ~w17214 & w11091;
assign w275 = ~w6830 & ~w7164;
assign w276 = ~w7950 & ~w817;
assign w277 = ~w17129 & w16387;
assign w278 = ~w4270 & ~w14740;
assign w279 = ~w10533 & ~w15196;
assign w280 = (~w3093 & w13110) | (~w3093 & w1549) | (w13110 & w1549);
assign w281 = ~w15151 & w16388;
assign w282 = ~w10675 & ~w11850;
assign w283 = ~w15778 & ~w4912;
assign w284 = a_47 & a_54;
assign w285 = ~w9702 & ~w1943;
assign w286 = ~w11363 & ~w16365;
assign w287 = (w12263 & w12796) | (w12263 & w8405) | (w12796 & w8405);
assign w288 = ~w591 & ~w2585;
assign w289 = ~w13129 & ~w12604;
assign w290 = a_22 & a_34;
assign w291 = w18963 & w3118;
assign w292 = w14311 & ~w5952;
assign w293 = (w3020 & w6628) | (w3020 & w6472) | (w6628 & w6472);
assign w294 = w7949 & ~w18338;
assign w295 = ~w3285 & ~w16569;
assign w296 = ~w10208 & ~w15267;
assign w297 = w14135 & w901;
assign w298 = w16489 & w8063;
assign w299 = ~w14976 & w8322;
assign w300 = w13940 & ~w10833;
assign w301 = ~w15081 & ~w5109;
assign w302 = w527 & ~w1592;
assign w303 = (w6917 & w13082) | (w6917 & w10959) | (w13082 & w10959);
assign w304 = a_22 & a_38;
assign w305 = ~w15868 & ~w18278;
assign w306 = ~w14731 & ~w7651;
assign w307 = ~w5057 & ~w17587;
assign w308 = ~w1163 & ~w19062;
assign w309 = ~w16555 & ~w4498;
assign w310 = ~w15711 & ~w1174;
assign w311 = w14071 & ~w18489;
assign w312 = ~w573 & ~w3823;
assign w313 = a_34 & a_53;
assign w314 = ~w9441 & ~w14882;
assign w315 = (~w3144 & ~w5151) | (~w3144 & w12889) | (~w5151 & w12889);
assign w316 = ~w12120 & ~w15534;
assign w317 = w8502 & w6198;
assign w318 = ~w13757 & ~w13257;
assign w319 = w3718 & ~w3475;
assign w320 = ~w8337 & ~w16239;
assign w321 = ~w1525 & ~w15553;
assign w322 = w5292 & ~w3375;
assign w323 = ~w5788 & ~w1584;
assign w324 = ~w2899 & ~w2553;
assign w325 = ~w5807 & ~w11049;
assign w326 = ~w14773 & ~w2156;
assign w327 = (w901 & w13100) | (w901 & w297) | (w13100 & w297);
assign w328 = ~w9220 & ~w16871;
assign w329 = a_5 & a_51;
assign w330 = a_16 & a_39;
assign w331 = ~w14192 & ~w13471;
assign w332 = ~w14210 & w7779;
assign w333 = w15116 & ~w16983;
assign w334 = w13434 & ~w7108;
assign w335 = ~w12308 & ~w5563;
assign w336 = ~w12382 & w597;
assign w337 = a_32 & a_41;
assign w338 = ~w10705 & w10864;
assign w339 = w7709 & ~w6151;
assign w340 = w5939 & w2992;
assign w341 = ~w16012 & ~w2696;
assign w342 = ~w8956 & w10292;
assign w343 = ~w8531 & ~w16281;
assign w344 = ~w6098 & w4931;
assign w345 = w8024 & ~w18960;
assign w346 = ~w4989 & ~w12860;
assign w347 = ~w8558 & ~w14987;
assign w348 = ~w3172 & ~w16110;
assign w349 = w2580 & ~w14474;
assign w350 = ~w3331 & ~w16280;
assign w351 = ~w7451 & ~w9752;
assign w352 = a_16 & a_47;
assign w353 = a_39 & a_49;
assign w354 = w3961 & w19025;
assign w355 = w13082 & ~w18870;
assign w356 = w3596 & w5997;
assign w357 = ~w9394 & ~w6668;
assign w358 = ~w11438 & ~w4041;
assign w359 = ~w14712 & w8377;
assign w360 = w10042 & w11743;
assign w361 = ~w6447 & ~w13478;
assign w362 = a_17 & a_39;
assign w363 = ~w15234 & ~w14095;
assign w364 = (~w8636 & ~w6335) | (~w8636 & w4413) | (~w6335 & w4413);
assign w365 = w2242 & ~w13829;
assign w366 = w7242 & ~w8416;
assign w367 = ~w14408 & ~w11310;
assign w368 = a_21 & a_46;
assign w369 = (~w13493 & ~w6723) | (~w13493 & w6415) | (~w6723 & w6415);
assign w370 = ~w4588 & ~w1042;
assign w371 = a_15 & a_18;
assign w372 = w13569 & ~w17472;
assign w373 = w5327 & w7171;
assign w374 = w4996 & ~w17309;
assign w375 = w1386 & w12765;
assign w376 = ~w2591 & w15793;
assign w377 = (~w6594 & ~w7934) | (~w6594 & w6980) | (~w7934 & w6980);
assign w378 = a_13 & a_56;
assign w379 = w9515 & w18956;
assign w380 = (w11523 & w17292) | (w11523 & w18017) | (w17292 & w18017);
assign w381 = ~w17989 & ~w727;
assign w382 = w18005 & w6033;
assign w383 = ~w1273 & ~w13936;
assign w384 = w9882 & w1930;
assign w385 = a_22 & a_56;
assign w386 = ~w15676 & ~w126;
assign w387 = w10359 & ~w963;
assign w388 = ~w1081 & ~w3105;
assign w389 = ~w5325 & w13233;
assign w390 = w14625 & ~w998;
assign w391 = ~w8229 & w9429;
assign w392 = ~w11333 & w18408;
assign w393 = ~w3082 & ~w10259;
assign w394 = w9074 & ~w5268;
assign w395 = ~w11316 & w4081;
assign w396 = ~w14725 & ~w14380;
assign w397 = ~w897 & w1981;
assign w398 = ~w7308 & ~w3012;
assign w399 = ~w15607 & ~w15551;
assign w400 = w4260 & ~w11471;
assign w401 = ~w2799 & w335;
assign w402 = w6289 & ~w8696;
assign w403 = ~w12237 & ~w17173;
assign w404 = w2762 & ~w10563;
assign w405 = ~w15728 & w608;
assign w406 = ~w10881 & ~w5645;
assign w407 = (~w15233 & ~w16162) | (~w15233 & w16578) | (~w16162 & w16578);
assign w408 = (w963 & w10840) | (w963 & w6589) | (w10840 & w6589);
assign w409 = w18091 & w17170;
assign w410 = (w7038 & w8471) | (w7038 & w2958) | (w8471 & w2958);
assign w411 = w14067 & w10274;
assign w412 = ~w12764 & ~w17124;
assign w413 = ~w2161 & ~w11992;
assign w414 = w9663 & ~w879;
assign w415 = w3802 & ~w6768;
assign w416 = ~w6624 & ~w12436;
assign w417 = ~w10729 & ~w5040;
assign w418 = w4187 & ~w5396;
assign w419 = ~w4943 & ~w2334;
assign w420 = a_15 & a_61;
assign w421 = ~w10363 & w13101;
assign w422 = ~w11873 & ~w18665;
assign w423 = ~w4775 & ~w14114;
assign w424 = a_38 & w10055;
assign w425 = a_0 & a_38;
assign w426 = (w2615 & w2769) | (w2615 & w17039) | (w2769 & w17039);
assign w427 = ~w14170 & ~w9688;
assign w428 = w407 & ~w16145;
assign w429 = ~w2528 & ~w11775;
assign w430 = ~w15285 & ~w2649;
assign w431 = w3084 & w16000;
assign w432 = ~w10539 & ~w8178;
assign w433 = ~w3907 & ~w15457;
assign w434 = (~w18883 & ~w2413) | (~w18883 & w2252) | (~w2413 & w2252);
assign w435 = ~w3311 & ~w16244;
assign w436 = w17946 & ~w16275;
assign w437 = ~w11698 & ~w6967;
assign w438 = ~w15759 & ~w12980;
assign w439 = w8504 & ~w12350;
assign w440 = ~w19027 & ~w12637;
assign w441 = (~w10388 & ~w4428) | (~w10388 & w9592) | (~w4428 & w9592);
assign w442 = ~w1778 & w15429;
assign w443 = w17664 & w9613;
assign w444 = ~w18487 & w5052;
assign w445 = ~w7704 & ~w16167;
assign w446 = ~w17181 & ~w11223;
assign w447 = w5023 & ~w2571;
assign w448 = ~w9347 & w6877;
assign w449 = ~w6495 & ~w5921;
assign w450 = ~w17136 & ~w12805;
assign w451 = w2857 & ~w2275;
assign w452 = w11126 & ~w1341;
assign w453 = (~w5073 & w15845) | (~w5073 & w11294) | (w15845 & w11294);
assign w454 = ~w12933 & ~w7522;
assign w455 = ~w7465 & ~w6783;
assign w456 = ~w18598 & w12292;
assign w457 = ~w10418 & ~w16799;
assign w458 = a_46 & a_54;
assign w459 = ~w17691 & ~w3141;
assign w460 = ~w15044 & ~w10205;
assign w461 = (a_46 & w2228) | (a_46 & w9231) | (w2228 & w9231);
assign w462 = ~w3884 & ~w7675;
assign w463 = ~w6800 & ~w10106;
assign w464 = w11859 & w14069;
assign w465 = w3148 & w6016;
assign w466 = ~w2299 & ~w12574;
assign w467 = a_23 & a_26;
assign w468 = (~w15988 & w7512) | (~w15988 & w2676) | (w7512 & w2676);
assign w469 = ~w18017 & w15644;
assign w470 = w1225 & w2992;
assign w471 = ~w1153 & ~w3772;
assign w472 = ~w6301 & ~w14682;
assign w473 = ~w7503 & ~w141;
assign w474 = ~w10236 & w10806;
assign w475 = ~w4348 & ~w11200;
assign w476 = ~w2608 & ~w5502;
assign w477 = ~w16278 & ~w11453;
assign w478 = ~w16910 & ~w5821;
assign w479 = a_15 & a_22;
assign w480 = w13214 & ~w11446;
assign w481 = a_9 & a_56;
assign w482 = ~w16673 & ~w7653;
assign w483 = ~w2814 & ~w4608;
assign w484 = w18718 & ~w13979;
assign w485 = ~w14509 & w1487;
assign w486 = w18180 & w8496;
assign w487 = (~w963 & w8052) | (~w963 & w387) | (w8052 & w387);
assign w488 = ~w3508 & ~w1178;
assign w489 = ~w13198 & ~w11809;
assign w490 = a_7 & a_39;
assign w491 = w9649 & ~w3411;
assign w492 = w13940 & ~w5937;
assign w493 = ~w12613 & ~w6477;
assign w494 = w2251 & w13430;
assign w495 = w6811 & ~w17516;
assign w496 = ~w12131 & ~w17420;
assign w497 = ~w16696 & ~w277;
assign w498 = ~w13305 & ~w7986;
assign w499 = ~w8482 & w13855;
assign w500 = ~w9250 & w8636;
assign w501 = ~w17149 & w36;
assign w502 = w3972 & w2866;
assign w503 = (~w13344 & ~w10057) | (~w13344 & w7789) | (~w10057 & w7789);
assign w504 = ~w7446 & w15867;
assign w505 = (~w6917 & w4023) | (~w6917 & w5618) | (w4023 & w5618);
assign w506 = a_31 & a_37;
assign w507 = w3187 & w17743;
assign w508 = ~w13519 & ~w11462;
assign w509 = a_27 & a_43;
assign w510 = ~w2343 & w7093;
assign w511 = ~w15887 & ~w12179;
assign w512 = ~w12746 & w15145;
assign w513 = ~w15012 & ~w17394;
assign w514 = ~w18650 & w10754;
assign w515 = w19124 | w13018;
assign w516 = ~w6853 & w1007;
assign w517 = ~w2509 & ~w18605;
assign w518 = ~w16138 & ~w12461;
assign w519 = a_25 & a_34;
assign w520 = ~w8971 & ~w6928;
assign w521 = ~w11205 & w1439;
assign w522 = a_6 & a_12;
assign w523 = w318 & w3750;
assign w524 = w4459 & ~w1714;
assign w525 = ~w8942 & w17954;
assign w526 = ~w10475 & ~w10938;
assign w527 = ~w17625 & ~w9185;
assign w528 = w6926 & w13343;
assign w529 = w3805 & ~w4158;
assign w530 = a_35 & a_38;
assign w531 = (w16007 & w8645) | (w16007 & w11624) | (w8645 & w11624);
assign w532 = ~w12664 & w517;
assign w533 = ~w18186 & ~w10131;
assign w534 = a_8 & a_23;
assign w535 = ~w6688 & w14088;
assign w536 = ~w15881 & ~w6603;
assign w537 = ~w5982 & ~w19050;
assign w538 = w5977 & w68;
assign w539 = ~w2572 & w17317;
assign w540 = w927 & w9847;
assign w541 = ~w7926 & w17201;
assign w542 = w17836 & w12162;
assign w543 = ~w5974 & ~w7942;
assign w544 = w8349 & w10391;
assign w545 = ~w14429 & w3232;
assign w546 = ~w18381 & ~w8845;
assign w547 = ~w4553 & ~w10090;
assign w548 = ~w9060 & w3437;
assign w549 = ~w15858 & w8537;
assign w550 = ~w8577 & ~w6055;
assign w551 = a_11 & a_60;
assign w552 = (~w7825 & w18980) | (~w7825 & w12692) | (w18980 & w12692);
assign w553 = ~w1786 & ~w8062;
assign w554 = ~w11220 & ~w18694;
assign w555 = ~w507 & ~w213;
assign w556 = ~w9808 & ~w7135;
assign w557 = ~w15362 & ~w7665;
assign w558 = w17096 & ~w16377;
assign w559 = ~w10980 & ~w2928;
assign w560 = ~w6397 & w4316;
assign w561 = ~w7409 & w6167;
assign w562 = a_9 & a_47;
assign w563 = a_3 & a_60;
assign w564 = ~w4622 & ~w18815;
assign w565 = ~w8444 & ~w11463;
assign w566 = ~w7860 & ~w9387;
assign w567 = w16537 & ~w5316;
assign w568 = (w11351 & w10330) | (w11351 & w8566) | (w10330 & w8566);
assign w569 = ~w14533 & w1133;
assign w570 = w4940 & w909;
assign w571 = ~w11739 & ~w283;
assign w572 = ~w8467 & ~w6614;
assign w573 = w5797 & w2859;
assign w574 = ~w13077 & ~w2736;
assign w575 = ~w4233 & ~w7803;
assign w576 = a_21 & a_37;
assign w577 = (w1916 & w2769) | (w1916 & w5297) | (w2769 & w5297);
assign w578 = a_16 & a_62;
assign w579 = ~w1314 & ~w1070;
assign w580 = ~w11011 & ~w12967;
assign w581 = a_60 & a_63;
assign w582 = ~w3264 & ~w5088;
assign w583 = ~w9914 & ~w14655;
assign w584 = ~w14211 & w17448;
assign w585 = ~w2448 & w17474;
assign w586 = ~w11991 & ~w16938;
assign w587 = a_28 & a_43;
assign w588 = ~w9158 & ~w11087;
assign w589 = w4557 & ~w10897;
assign w590 = ~w17025 & ~w11378;
assign w591 = w8243 & w581;
assign w592 = ~w14745 & ~w4667;
assign w593 = ~w11115 & w2812;
assign w594 = ~w13585 & ~w12656;
assign w595 = w15288 & ~w18594;
assign w596 = a_35 & a_44;
assign w597 = ~w1102 & ~w6754;
assign w598 = w4280 & ~w4935;
assign w599 = w2880 & ~w14280;
assign w600 = a_30 & a_32;
assign w601 = w14165 & ~w6046;
assign w602 = w16440 & ~w1734;
assign w603 = w18752 & w7706;
assign w604 = ~w18861 & ~w15967;
assign w605 = ~w16403 & w12616;
assign w606 = ~w12764 & ~w14525;
assign w607 = ~w10933 & w12121;
assign w608 = ~w9988 & ~w7398;
assign w609 = ~a_10 & ~w18633;
assign w610 = w11725 & w11343;
assign w611 = ~w10744 & ~w3703;
assign w612 = a_30 & a_44;
assign w613 = ~w7965 & ~w616;
assign w614 = (~w5569 & ~w9593) | (~w5569 & w7207) | (~w9593 & w7207);
assign w615 = w13061 & ~w3001;
assign w616 = ~w7633 & ~w2472;
assign w617 = ~w8391 & ~w11298;
assign w618 = w9318 & ~w8486;
assign w619 = w14339 & w19146;
assign w620 = ~w8389 & ~w18793;
assign w621 = ~w16591 & ~w18581;
assign w622 = w9403 & ~w1522;
assign w623 = (~w16516 & ~w12901) | (~w16516 & w15885) | (~w12901 & w15885);
assign w624 = (~w15474 & ~w17272) | (~w15474 & w16511) | (~w17272 & w16511);
assign w625 = w6679 & w3555;
assign w626 = w3303 & ~w4901;
assign w627 = a_15 & a_20;
assign w628 = (~w11258 & ~w13598) | (~w11258 & w7694) | (~w13598 & w7694);
assign w629 = ~w9695 & w11667;
assign w630 = ~w7696 & ~w14763;
assign w631 = ~w4900 & w11932;
assign w632 = ~w14528 & w15522;
assign w633 = ~w14470 & ~w10552;
assign w634 = a_34 & a_51;
assign w635 = w15715 & ~w1636;
assign w636 = ~w10932 & ~w1080;
assign w637 = ~w2690 & ~w11280;
assign w638 = ~w13373 & w10442;
assign w639 = ~w867 & ~w19020;
assign w640 = ~w10190 & ~w5539;
assign w641 = w2548 & w18267;
assign w642 = ~w9762 & ~w2755;
assign w643 = ~w8665 & w15850;
assign w644 = ~w4784 & ~w1547;
assign w645 = w4372 & w17295;
assign w646 = w14356 & ~w16266;
assign w647 = ~w10349 & w1344;
assign w648 = ~w6363 & w4769;
assign w649 = w16447 & ~w14300;
assign w650 = ~w16187 & ~w60;
assign w651 = ~w3343 & ~w13477;
assign w652 = w12760 & ~w15262;
assign w653 = a_12 & a_58;
assign w654 = w1306 & ~w10549;
assign w655 = ~w5303 & ~w6947;
assign w656 = ~w7490 & ~w4238;
assign w657 = w15915 & ~w14415;
assign w658 = a_2 & a_38;
assign w659 = ~w16138 & ~w4500;
assign w660 = w4451 & ~w6069;
assign w661 = w10733 & ~w5211;
assign w662 = ~w12002 & ~w12788;
assign w663 = (w8699 & ~w1962) | (w8699 & w12943) | (~w1962 & w12943);
assign w664 = (w11667 & ~w5866) | (w11667 & w629) | (~w5866 & w629);
assign w665 = ~w14659 & ~w2668;
assign w666 = (w1566 & w515) | (w1566 & w16839) | (w515 & w16839);
assign w667 = w15901 & w17393;
assign w668 = w1320 & w44;
assign w669 = a_9 & a_17;
assign w670 = ~w11979 & ~w17965;
assign w671 = a_41 & a_53;
assign w672 = ~w6835 & ~w4437;
assign w673 = a_29 & a_37;
assign w674 = ~w10723 & ~w10695;
assign w675 = ~w14672 & ~w18568;
assign w676 = a_43 & a_60;
assign w677 = ~w12260 & ~w7264;
assign w678 = a_54 & a_58;
assign w679 = ~w10721 & ~w14687;
assign w680 = a_17 & w11297;
assign w681 = ~w16039 & w2049;
assign w682 = (w13037 & w2769) | (w13037 & w15312) | (w2769 & w15312);
assign w683 = ~w771 & ~w15981;
assign w684 = w369 & ~w1571;
assign w685 = ~w10792 & ~w7453;
assign w686 = ~w5559 & ~w13972;
assign w687 = ~w476 & ~w1539;
assign w688 = ~w14397 & ~w18280;
assign w689 = ~w4590 & ~w9050;
assign w690 = a_38 & a_49;
assign w691 = ~w1747 & ~w15724;
assign w692 = ~w207 & w7127;
assign w693 = w16493 & ~w12040;
assign w694 = a_42 & a_53;
assign w695 = ~w14377 & ~w1556;
assign w696 = ~w15732 & ~w4382;
assign w697 = a_9 & a_45;
assign w698 = w12230 & ~w11716;
assign w699 = ~w13913 & ~w4130;
assign w700 = ~w5654 & w18865;
assign w701 = ~w4527 & w13947;
assign w702 = ~w1366 & ~w16184;
assign w703 = w16287 & ~w14956;
assign w704 = ~w5418 & ~w3357;
assign w705 = a_11 & a_57;
assign w706 = ~w11430 & w3858;
assign w707 = w8588 & ~w6845;
assign w708 = ~w13752 & ~w9068;
assign w709 = ~w723 & ~w8042;
assign w710 = ~w8886 & ~w11921;
assign w711 = ~w18640 & ~w10970;
assign w712 = ~w3165 & w9950;
assign w713 = ~w5503 & ~w2845;
assign w714 = ~w9890 & ~w2945;
assign w715 = w7134 & ~w13482;
assign w716 = w7337 & w15320;
assign w717 = ~w14220 & ~w12972;
assign w718 = ~a_55 & a_56;
assign w719 = a_25 & a_61;
assign w720 = ~w2029 & ~w4256;
assign w721 = a_35 & a_53;
assign w722 = w9481 & ~w9274;
assign w723 = ~w2601 & ~w4626;
assign w724 = a_62 & a_63;
assign w725 = ~w11355 & ~w5903;
assign w726 = w6545 & ~w723;
assign w727 = ~w3069 & ~w15743;
assign w728 = ~w18052 & w7107;
assign w729 = w5697 & ~w16243;
assign w730 = ~w407 & w16145;
assign w731 = ~w19061 & ~w4452;
assign w732 = ~w13221 & ~w1885;
assign w733 = w8360 & ~w1429;
assign w734 = a_15 & a_37;
assign w735 = ~w17196 & ~w12716;
assign w736 = w17167 & w14546;
assign w737 = a_29 & a_53;
assign w738 = ~w9889 & w8137;
assign w739 = ~w12995 & ~w8852;
assign w740 = ~w10134 & ~w5722;
assign w741 = w16992 & ~w14491;
assign w742 = ~w5743 & w12887;
assign w743 = (~w12853 & ~w15918) | (~w12853 & w15977) | (~w15918 & w15977);
assign w744 = ~w963 & w1713;
assign w745 = ~w4902 & ~w7577;
assign w746 = (~w17101 & ~w927) | (~w17101 & w17705) | (~w927 & w17705);
assign w747 = ~w4030 & w4875;
assign w748 = ~w14759 & w2559;
assign w749 = ~w5022 & w18340;
assign w750 = ~w12841 & ~w10384;
assign w751 = ~w12797 & w13170;
assign w752 = (w8386 & w8345) | (w8386 & w17673) | (w8345 & w17673);
assign w753 = a_44 & a_48;
assign w754 = w2201 & ~w1640;
assign w755 = ~w6875 & ~w17979;
assign w756 = ~w13888 & w15050;
assign w757 = (w7604 & w8052) | (w7604 & w19091) | (w8052 & w19091);
assign w758 = w8286 & ~w10790;
assign w759 = w9175 & w1029;
assign w760 = (~w9710 & ~w15238) | (~w9710 & w9006) | (~w15238 & w9006);
assign w761 = w8710 & w9961;
assign w762 = w14486 & ~w7388;
assign w763 = w2881 & ~w18152;
assign w764 = ~w6000 & ~w8037;
assign w765 = ~w8788 & ~w17371;
assign w766 = w3188 & w12117;
assign w767 = ~w9682 & ~w3096;
assign w768 = w6990 & w12517;
assign w769 = w18464 & w2993;
assign w770 = ~w2969 & ~w9323;
assign w771 = w18251 & w11630;
assign w772 = ~w5448 & ~w601;
assign w773 = ~w18832 & w1388;
assign w774 = w9261 & w12869;
assign w775 = ~w369 & w18332;
assign w776 = a_7 & a_23;
assign w777 = w6550 & w3115;
assign w778 = (w6396 & w4170) | (w6396 & w14979) | (w4170 & w14979);
assign w779 = ~w6096 & w17461;
assign w780 = ~w9478 & w13396;
assign w781 = ~w8407 & ~w13636;
assign w782 = ~w5593 & w13401;
assign w783 = w15261 & ~w16629;
assign w784 = ~w15364 & ~w2066;
assign w785 = ~w3242 & ~w9683;
assign w786 = a_23 & a_53;
assign w787 = w16639 & ~w9161;
assign w788 = w7168 & w2749;
assign w789 = ~w19100 & ~w7543;
assign w790 = a_3 & a_46;
assign w791 = ~w1175 & ~w6159;
assign w792 = a_22 & a_63;
assign w793 = ~w13361 & ~w11561;
assign w794 = ~w567 & ~w1535;
assign w795 = ~w13809 & ~w2397;
assign w796 = ~w12420 & ~w17420;
assign w797 = ~w16634 & ~w18522;
assign w798 = w11822 & ~w10103;
assign w799 = ~w16426 & ~w5894;
assign w800 = w8323 & ~w10189;
assign w801 = ~w18310 & ~w14496;
assign w802 = w7298 & ~w7790;
assign w803 = ~w88 & ~w4409;
assign w804 = (w18718 & w19005) | (w18718 & w9033) | (w19005 & w9033);
assign w805 = w13086 & w4957;
assign w806 = ~w4069 & ~w19126;
assign w807 = w6770 & w4229;
assign w808 = a_8 & a_55;
assign w809 = ~w17054 & ~w15146;
assign w810 = w7388 & ~w559;
assign w811 = (~w14357 & ~w3880) | (~w14357 & w9936) | (~w3880 & w9936);
assign w812 = w10079 & ~w8003;
assign w813 = ~w13491 & ~w16777;
assign w814 = w8357 & ~w11552;
assign w815 = a_30 & a_59;
assign w816 = w7295 & ~w17951;
assign w817 = a_0 & a_42;
assign w818 = w15238 & ~w15730;
assign w819 = w205 & ~w1605;
assign w820 = ~w3818 & w9927;
assign w821 = ~w13553 & ~w18503;
assign w822 = ~w9439 & ~w7710;
assign w823 = ~w4967 & ~w8162;
assign w824 = ~w19013 & ~w1685;
assign w825 = w2868 & ~w10550;
assign w826 = ~w10222 & ~w1643;
assign w827 = ~w15794 & w7656;
assign w828 = ~w7471 & ~w15090;
assign w829 = ~w19093 & ~w17956;
assign w830 = w12688 & ~w12110;
assign w831 = w6031 & ~w12247;
assign w832 = w10615 & ~w13059;
assign w833 = ~w11818 & ~w10227;
assign w834 = a_44 & w15517;
assign w835 = w6146 & ~w197;
assign w836 = a_18 & a_46;
assign w837 = ~w14627 & ~w8882;
assign w838 = ~w5011 & ~w4473;
assign w839 = ~w17915 & ~w13514;
assign w840 = ~w9701 & ~w12595;
assign w841 = ~w14046 & ~w5848;
assign w842 = (w19099 & ~w8987) | (w19099 & w16383) | (~w8987 & w16383);
assign w843 = ~w11648 & ~w5983;
assign w844 = ~w18125 & ~w1866;
assign w845 = ~w10812 & w10803;
assign w846 = ~w182 & ~w9677;
assign w847 = w464 & ~w14949;
assign w848 = ~w84 & ~w15110;
assign w849 = ~w3880 & w13476;
assign w850 = ~w8922 & ~w11581;
assign w851 = w10234 & ~w8048;
assign w852 = ~w3587 & ~w9739;
assign w853 = a_33 & a_43;
assign w854 = ~w10025 & ~w12101;
assign w855 = ~w157 & w19002;
assign w856 = w14012 & ~w986;
assign w857 = ~w7440 & ~w10213;
assign w858 = ~w15605 & ~w18271;
assign w859 = ~w16299 & ~w8770;
assign w860 = ~w17560 & ~w17742;
assign w861 = (~w293 & ~w1836) | (~w293 & w18549) | (~w1836 & w18549);
assign w862 = ~w6903 & ~w12886;
assign w863 = (~w5610 & w19005) | (~w5610 & w15956) | (w19005 & w15956);
assign w864 = ~w16556 & ~w17708;
assign w865 = ~w3757 & ~w10037;
assign w866 = a_36 & a_58;
assign w867 = ~w12873 & ~w9939;
assign w868 = a_37 & a_39;
assign w869 = w5165 & ~w7095;
assign w870 = a_31 & a_34;
assign w871 = w4883 & ~w10490;
assign w872 = w15353 & w9217;
assign w873 = a_8 & a_46;
assign w874 = (w7102 & w10788) | (w7102 & w7811) | (w10788 & w7811);
assign w875 = ~w1135 & w12003;
assign w876 = ~w1984 & ~w5946;
assign w877 = ~w301 & ~w8823;
assign w878 = ~w920 & ~w66;
assign w879 = w4644 & w8333;
assign w880 = w15230 & ~w2309;
assign w881 = w6268 & w2488;
assign w882 = ~w12894 & ~w12133;
assign w883 = ~w13326 & w14040;
assign w884 = ~w5323 & w6542;
assign w885 = ~w12702 & ~w15278;
assign w886 = w2626 & ~w17575;
assign w887 = ~w1627 & w2459;
assign w888 = (w5781 & w5518) | (w5781 & w19147) | (w5518 & w19147);
assign w889 = ~w6853 & w7243;
assign w890 = a_6 & a_16;
assign w891 = w2834 & ~w8143;
assign w892 = a_15 & a_50;
assign w893 = ~w5973 & ~w10112;
assign w894 = ~w16496 & ~w9188;
assign w895 = w18259 & w7370;
assign w896 = ~w17268 & w18038;
assign w897 = ~w17328 & ~w3559;
assign w898 = ~w671 & ~w253;
assign w899 = w18130 & ~w4874;
assign w900 = w17395 & ~w7225;
assign w901 = ~w16345 & ~w9537;
assign w902 = ~w12521 & ~w4959;
assign w903 = w9835 & ~w12930;
assign w904 = w1577 & ~w6594;
assign w905 = ~w16232 & ~w9989;
assign w906 = w7994 & ~w4695;
assign w907 = w1811 & w18931;
assign w908 = ~w2642 & w2114;
assign w909 = ~w13445 & ~w11747;
assign w910 = ~w16285 & ~w17663;
assign w911 = w11933 & w9401;
assign w912 = w2255 & w11617;
assign w913 = ~w7589 & ~w5345;
assign w914 = ~w8956 & ~w18285;
assign w915 = ~w17050 & ~w17407;
assign w916 = ~w18704 & ~w5198;
assign w917 = ~w16327 & ~w11015;
assign w918 = ~w15041 & w4436;
assign w919 = w7276 & ~w3661;
assign w920 = w7950 & w817;
assign w921 = ~w16881 & ~w5935;
assign w922 = ~w16132 & ~w3648;
assign w923 = ~w1113 & w15659;
assign w924 = ~w8606 & w13532;
assign w925 = w10789 & w9673;
assign w926 = (~w1997 & ~w1220) | (~w1997 & w12964) | (~w1220 & w12964);
assign w927 = (~w11748 & w553) | (~w11748 & w6876) | (w553 & w6876);
assign w928 = w7868 & ~w13514;
assign w929 = a_5 & a_11;
assign w930 = a_11 & a_30;
assign w931 = ~w18886 & ~w11142;
assign w932 = ~w7815 & ~w18925;
assign w933 = a_0 & a_54;
assign w934 = w6060 & ~w3060;
assign w935 = ~w8461 & ~w13631;
assign w936 = w12946 & w16834;
assign w937 = w13067 & ~w6188;
assign w938 = ~a_12 & w6280;
assign w939 = ~w18562 & w7149;
assign w940 = ~w1465 & ~w2055;
assign w941 = a_38 & a_40;
assign w942 = ~w6259 & ~w349;
assign w943 = w15183 & ~w10182;
assign w944 = ~w16463 & w17113;
assign w945 = ~w8612 & w4721;
assign w946 = w2444 & ~w7725;
assign w947 = ~w15611 & ~w3553;
assign w948 = ~w274 & ~w9159;
assign w949 = ~w3413 & ~w11703;
assign w950 = ~w6114 & ~w15723;
assign w951 = w10264 & w13659;
assign w952 = ~w4042 & ~w9671;
assign w953 = w16384 & ~w14866;
assign w954 = w866 & ~w6020;
assign w955 = ~w13249 & ~w12085;
assign w956 = a_28 & a_35;
assign w957 = ~w10503 & ~w14540;
assign w958 = ~w5510 & ~w2997;
assign w959 = w5335 & ~w16743;
assign w960 = ~w8348 & ~w11120;
assign w961 = w10529 & ~w6136;
assign w962 = ~w12482 & ~w5275;
assign w963 = w1977 & w1621;
assign w964 = w4147 & ~w10024;
assign w965 = a_8 & a_11;
assign w966 = ~w11698 & ~w2059;
assign w967 = ~w12053 & ~w2077;
assign w968 = a_16 & a_27;
assign w969 = a_33 & a_46;
assign w970 = ~w29 & ~w6533;
assign w971 = w10629 & w8036;
assign w972 = w12805 & w17136;
assign w973 = w14012 & w7117;
assign w974 = ~w7199 & w10547;
assign w975 = ~w17759 & ~w230;
assign w976 = ~w7688 & ~w14285;
assign w977 = a_28 & a_53;
assign w978 = w267 & ~w2686;
assign w979 = w3846 & w18346;
assign w980 = w18197 & w8026;
assign w981 = ~w14407 & ~w2417;
assign w982 = w12497 & ~w1462;
assign w983 = w13979 & w18843;
assign w984 = ~w442 & ~w10695;
assign w985 = (w11173 & w2769) | (w11173 & w18254) | (w2769 & w18254);
assign w986 = ~w17006 & ~w7765;
assign w987 = ~w4389 & ~w2765;
assign w988 = ~a_15 & ~w5867;
assign w989 = ~w11936 & ~w11487;
assign w990 = ~w18656 & ~w10133;
assign w991 = ~w3180 & ~w3376;
assign w992 = ~w16433 & ~w14562;
assign w993 = a_39 & a_47;
assign w994 = w10991 & ~w10745;
assign w995 = ~w12509 & ~w12785;
assign w996 = ~w17544 & w18062;
assign w997 = ~w16878 & ~w14630;
assign w998 = w16267 & ~w18922;
assign w999 = w14398 & ~w13035;
assign w1000 = ~w2183 & w7733;
assign w1001 = ~w11905 & ~w2264;
assign w1002 = w14428 & ~w17226;
assign w1003 = w16072 & w2894;
assign w1004 = w10720 & ~w1288;
assign w1005 = ~w4734 & w13137;
assign w1006 = ~w7492 & ~w2344;
assign w1007 = (~w3175 & w10330) | (~w3175 & w14228) | (w10330 & w14228);
assign w1008 = w149 & w522;
assign w1009 = ~w4548 & w19138;
assign w1010 = a_3 & a_42;
assign w1011 = ~w14644 & ~w9985;
assign w1012 = a_36 & a_37;
assign w1013 = w15349 & w2186;
assign w1014 = ~w11501 & ~w12062;
assign w1015 = ~w5060 & ~w264;
assign w1016 = a_53 & a_62;
assign w1017 = ~w2918 & ~w2410;
assign w1018 = ~w180 & w11086;
assign w1019 = ~w10335 & ~w1739;
assign w1020 = (~w6134 & w5772) | (~w6134 & w3779) | (w5772 & w3779);
assign w1021 = ~w13698 & ~w16688;
assign w1022 = ~w15822 & ~w10743;
assign w1023 = w992 & ~w2051;
assign w1024 = w6096 & ~w17461;
assign w1025 = w7564 & ~w4964;
assign w1026 = a_28 & a_47;
assign w1027 = a_19 & a_21;
assign w1028 = w5343 & w479;
assign w1029 = ~w17063 & ~w4536;
assign w1030 = a_27 & a_50;
assign w1031 = w3076 & w13320;
assign w1032 = ~w11269 & ~w14870;
assign w1033 = w15706 & w18811;
assign w1034 = a_4 & a_31;
assign w1035 = ~w3086 & ~w6750;
assign w1036 = w10099 & ~w983;
assign w1037 = ~w6066 & ~w9356;
assign w1038 = ~w13435 & ~w3352;
assign w1039 = ~w1348 & ~w6597;
assign w1040 = ~w14793 & w564;
assign w1041 = ~w15834 & ~w4036;
assign w1042 = ~w8862 & ~w11019;
assign w1043 = w84 & w15110;
assign w1044 = w7078 & ~w14817;
assign w1045 = ~w14499 & ~w1725;
assign w1046 = ~w18846 & w989;
assign w1047 = w3308 & w12169;
assign w1048 = w6473 & ~w1227;
assign w1049 = w13732 & ~w59;
assign w1050 = (~w14184 & w16917) | (~w14184 & w7334) | (w16917 & w7334);
assign w1051 = (~w13103 & w8863) | (~w13103 & w10471) | (w8863 & w10471);
assign w1052 = ~w1806 & w8846;
assign w1053 = w17786 & w9977;
assign w1054 = a_26 & a_60;
assign w1055 = w16650 & ~w8996;
assign w1056 = ~w4106 & ~w9009;
assign w1057 = ~w1145 & ~w14234;
assign w1058 = w18510 & w4109;
assign w1059 = w8899 & ~w12931;
assign w1060 = ~w4329 & w4532;
assign w1061 = ~w17805 & ~w16156;
assign w1062 = ~w12718 & ~w1508;
assign w1063 = a_22 & a_30;
assign w1064 = w221 & ~w7047;
assign w1065 = ~w12906 & ~w15569;
assign w1066 = w16547 & w5312;
assign w1067 = w14052 & w16781;
assign w1068 = w9150 & w2956;
assign w1069 = ~w19099 & ~w17104;
assign w1070 = w3306 & w5993;
assign w1071 = ~w18406 & ~w18411;
assign w1072 = w10763 & ~w7236;
assign w1073 = a_1 & a_51;
assign w1074 = ~w15103 & w13668;
assign w1075 = ~w15768 & ~w6215;
assign w1076 = ~w12553 & ~w2423;
assign w1077 = ~w9568 & ~w2031;
assign w1078 = a_45 & a_55;
assign w1079 = ~w5805 & ~w12736;
assign w1080 = a_16 & a_44;
assign w1081 = w10810 & w3170;
assign w1082 = ~w11067 & w5025;
assign w1083 = ~w9282 & ~w18912;
assign w1084 = ~w13032 & ~w15625;
assign w1085 = ~w5651 & ~w4031;
assign w1086 = (~w7102 & w1036) | (~w7102 & w15369) | (w1036 & w15369);
assign w1087 = ~w10879 & w3355;
assign w1088 = ~w12744 & w1432;
assign w1089 = ~w15897 & ~w2324;
assign w1090 = ~w17497 & w9749;
assign w1091 = ~w580 & ~w13456;
assign w1092 = ~w220 & ~w16488;
assign w1093 = ~w8318 & w15638;
assign w1094 = ~w2433 & ~w6772;
assign w1095 = (w1898 & w5168) | (w1898 & w5933) | (w5168 & w5933);
assign w1096 = w10048 & w1766;
assign w1097 = ~w10243 & ~w10787;
assign w1098 = ~w15252 & w8721;
assign w1099 = w6089 & w6435;
assign w1100 = ~w5032 & ~w13319;
assign w1101 = w14429 & ~w9934;
assign w1102 = w16489 & w2557;
assign w1103 = ~w5255 & ~w9569;
assign w1104 = w13888 & ~w15050;
assign w1105 = a_8 & a_43;
assign w1106 = w10954 & ~w8185;
assign w1107 = w13804 & ~w3558;
assign w1108 = w8317 & ~w3718;
assign w1109 = ~w13578 & ~w8329;
assign w1110 = a_4 & a_47;
assign w1111 = ~w9986 & w18386;
assign w1112 = ~w14220 & ~w17957;
assign w1113 = w11265 & w12341;
assign w1114 = ~w16457 & ~w16588;
assign w1115 = w14722 & ~w1960;
assign w1116 = ~w15350 & w9391;
assign w1117 = w482 & w3868;
assign w1118 = ~w7760 & ~w17791;
assign w1119 = (w15755 & w18279) | (w15755 & w18772) | (w18279 & w18772);
assign w1120 = ~w8059 & ~w13511;
assign w1121 = ~w3491 & w8015;
assign w1122 = w9651 & ~w4523;
assign w1123 = ~w11435 & ~w30;
assign w1124 = ~w11898 & ~w5493;
assign w1125 = w18228 & ~w9311;
assign w1126 = ~w12565 & w11917;
assign w1127 = ~w5331 & ~w14513;
assign w1128 = w9568 & w2031;
assign w1129 = ~w1114 & ~w18876;
assign w1130 = w14758 & ~w5492;
assign w1131 = ~w9576 & ~w18283;
assign w1132 = ~w14977 & ~w8066;
assign w1133 = ~w12138 & ~w2840;
assign w1134 = ~w4270 & ~w11713;
assign w1135 = a_10 & a_32;
assign w1136 = w3525 & ~w2105;
assign w1137 = (~w15457 & ~w13652) | (~w15457 & w433) | (~w13652 & w433);
assign w1138 = a_39 & a_62;
assign w1139 = ~w9607 & ~w4520;
assign w1140 = ~w5358 & ~w14283;
assign w1141 = ~w3897 & w14968;
assign w1142 = (w18016 & w2254) | (w18016 & w18834) | (w2254 & w18834);
assign w1143 = ~w17899 & w7379;
assign w1144 = ~w6886 & ~w12328;
assign w1145 = ~w7621 & ~w772;
assign w1146 = w14667 & w14605;
assign w1147 = w4182 & w7715;
assign w1148 = w11387 & w17208;
assign w1149 = w7295 & w2976;
assign w1150 = w13082 & ~w847;
assign w1151 = ~w3439 & ~w4246;
assign w1152 = ~w7644 & ~w19092;
assign w1153 = ~w18927 & ~w13572;
assign w1154 = ~w5368 & ~w15590;
assign w1155 = ~w302 & w16683;
assign w1156 = ~w9725 & ~w6955;
assign w1157 = a_15 & a_41;
assign w1158 = a_8 & a_12;
assign w1159 = ~w7212 & ~w19125;
assign w1160 = w4494 & w2101;
assign w1161 = w791 & w822;
assign w1162 = ~w17173 & ~w13060;
assign w1163 = ~w12862 & ~w16230;
assign w1164 = ~w6988 & w11408;
assign w1165 = ~w10330 & w1986;
assign w1166 = a_23 & a_54;
assign w1167 = w10059 & ~w15124;
assign w1168 = ~w4089 & w8437;
assign w1169 = ~w17506 & w3005;
assign w1170 = ~w9036 & ~w7100;
assign w1171 = w2342 & w13290;
assign w1172 = a_21 & a_27;
assign w1173 = ~w17689 & w14524;
assign w1174 = ~w9648 & w10125;
assign w1175 = w6545 & ~w709;
assign w1176 = w13144 & w9925;
assign w1177 = ~w8718 & w15101;
assign w1178 = ~w15391 & ~w4360;
assign w1179 = ~w18330 & w8288;
assign w1180 = ~w4862 & w16387;
assign w1181 = ~w18975 & w14273;
assign w1182 = ~w12335 & ~w12742;
assign w1183 = w71 & ~w11186;
assign w1184 = w10737 & w6190;
assign w1185 = w14442 & w3043;
assign w1186 = ~w8623 & ~w951;
assign w1187 = w17128 & w837;
assign w1188 = ~w4816 & ~w1516;
assign w1189 = ~w3905 & ~w15054;
assign w1190 = w633 & ~w236;
assign w1191 = a_7 & a_16;
assign w1192 = a_22 & a_25;
assign w1193 = w8816 & w9002;
assign w1194 = a_0 & a_53;
assign w1195 = w1056 & ~w6518;
assign w1196 = ~w13542 & ~w2453;
assign w1197 = (w6279 & ~w5866) | (w6279 & w9280) | (~w5866 & w9280);
assign w1198 = w15048 & ~w13063;
assign w1199 = ~w2072 & w4712;
assign w1200 = ~w12497 & w1462;
assign w1201 = ~w6294 & w15059;
assign w1202 = ~w16552 & ~w16414;
assign w1203 = ~w15686 & w12375;
assign w1204 = ~w3272 & ~w1415;
assign w1205 = (w2746 & w7289) | (w2746 & w14091) | (w7289 & w14091);
assign w1206 = w14591 & ~w12103;
assign w1207 = ~w13458 & ~w18502;
assign w1208 = a_2 & a_37;
assign w1209 = w7526 & ~w13549;
assign w1210 = w18447 & ~w18389;
assign w1211 = w4557 & ~w14929;
assign w1212 = a_3 & a_39;
assign w1213 = ~w5711 & w16869;
assign w1214 = ~w16941 & ~w1079;
assign w1215 = a_14 & a_56;
assign w1216 = ~w17138 & w2476;
assign w1217 = ~w2422 & ~w5244;
assign w1218 = ~w4407 & ~w5570;
assign w1219 = ~w3376 & ~w13759;
assign w1220 = ~w1997 & ~w11432;
assign w1221 = ~w14084 & ~w16319;
assign w1222 = a_0 & a_24;
assign w1223 = ~w16320 & ~w5554;
assign w1224 = a_19 & a_55;
assign w1225 = ~w7863 & ~w6402;
assign w1226 = ~w12135 & ~w13025;
assign w1227 = ~w3842 & ~w12193;
assign w1228 = ~w11599 & w7719;
assign w1229 = a_2 & a_20;
assign w1230 = w7363 & w18618;
assign w1231 = ~w9297 & w17256;
assign w1232 = ~w3119 & ~w14496;
assign w1233 = ~w2834 & w8143;
assign w1234 = ~w5686 & ~w467;
assign w1235 = w1758 & w4449;
assign w1236 = w19138 & ~w13118;
assign w1237 = ~w14355 & ~w13764;
assign w1238 = w5613 & w9831;
assign w1239 = ~w2732 & w1607;
assign w1240 = a_5 & a_21;
assign w1241 = w7063 & ~w3630;
assign w1242 = ~w835 & ~w13496;
assign w1243 = ~a_45 & a_46;
assign w1244 = w9324 & w18384;
assign w1245 = w18476 & w5905;
assign w1246 = ~w16452 & ~w395;
assign w1247 = w7407 & ~w18659;
assign w1248 = w15650 & w5138;
assign w1249 = ~w1373 & ~w3518;
assign w1250 = ~w8269 & ~w5347;
assign w1251 = w15801 & w11872;
assign w1252 = ~w12108 & w16684;
assign w1253 = a_5 & a_28;
assign w1254 = a_16 & a_54;
assign w1255 = ~w18952 & ~w12233;
assign w1256 = ~w15829 & w2929;
assign w1257 = ~w353 & ~w14344;
assign w1258 = w1759 & ~w3480;
assign w1259 = ~w15126 & ~w19026;
assign w1260 = ~w14851 & ~w6287;
assign w1261 = w13061 & w17162;
assign w1262 = ~w7553 & ~w19023;
assign w1263 = w18640 & ~w10459;
assign w1264 = w4658 & ~w12164;
assign w1265 = ~w14813 & w6053;
assign w1266 = ~w10139 & ~w14652;
assign w1267 = ~w9489 & ~w14077;
assign w1268 = (~w13769 & ~w4739) | (~w13769 & w18061) | (~w4739 & w18061);
assign w1269 = w8439 & ~w3984;
assign w1270 = ~w6046 & ~w5448;
assign w1271 = ~w12122 & w9412;
assign w1272 = ~w10732 & ~w7459;
assign w1273 = ~w11870 & w15442;
assign w1274 = w3567 & w16293;
assign w1275 = ~w7358 & ~w3042;
assign w1276 = ~w6367 & ~w9440;
assign w1277 = ~w6686 & ~w502;
assign w1278 = (~w891 & ~w3189) | (~w891 & w7946) | (~w3189 & w7946);
assign w1279 = ~w3380 & ~w17607;
assign w1280 = w4749 & ~w14954;
assign w1281 = ~w12851 & ~w3430;
assign w1282 = a_56 & a_61;
assign w1283 = (~w17668 & ~w9297) | (~w17668 & w6427) | (~w9297 & w6427);
assign w1284 = a_6 & a_58;
assign w1285 = ~w6761 & ~w17873;
assign w1286 = ~w1716 & ~w4089;
assign w1287 = w5746 & ~w8005;
assign w1288 = (~w222 & ~w11323) | (~w222 & w3694) | (~w11323 & w3694);
assign w1289 = ~w2104 & w921;
assign w1290 = (w7102 & w7826) | (w7102 & w1424) | (w7826 & w1424);
assign w1291 = w8806 & ~w14059;
assign w1292 = ~w7764 & w7395;
assign w1293 = w15205 & ~w494;
assign w1294 = ~w2305 & ~w13729;
assign w1295 = ~w13082 & w5552;
assign w1296 = ~w5977 & ~w68;
assign w1297 = ~w1737 & ~w17958;
assign w1298 = ~w5399 & ~w1121;
assign w1299 = ~w11930 & ~w17238;
assign w1300 = ~w260 & ~w15186;
assign w1301 = ~w4104 & ~w8295;
assign w1302 = a_7 & a_42;
assign w1303 = w12486 & w14520;
assign w1304 = ~w8345 & w16226;
assign w1305 = ~w18258 & ~w2641;
assign w1306 = ~w16773 & ~w598;
assign w1307 = a_55 & a_58;
assign w1308 = w8836 & w12595;
assign w1309 = w18997 & w5280;
assign w1310 = w280 & w5685;
assign w1311 = ~w7193 & ~w7684;
assign w1312 = (~w14326 & ~w17749) | (~w14326 & w14058) | (~w17749 & w14058);
assign w1313 = ~w8746 & ~w16022;
assign w1314 = ~w3306 & ~w5993;
assign w1315 = a_14 & a_33;
assign w1316 = ~w13318 & ~w5936;
assign w1317 = w14798 & ~w932;
assign w1318 = ~w1551 & ~w15945;
assign w1319 = w2706 & w16758;
assign w1320 = w16918 & ~w6426;
assign w1321 = w5930 & ~w11554;
assign w1322 = w16967 & w5679;
assign w1323 = ~w8078 & ~w1033;
assign w1324 = ~w11774 & ~w15688;
assign w1325 = w2183 & ~w7733;
assign w1326 = ~w13618 & ~w18290;
assign w1327 = ~w5103 & ~w18523;
assign w1328 = ~w4650 & ~w13266;
assign w1329 = ~w3646 & ~w10466;
assign w1330 = ~w16972 & ~w417;
assign w1331 = a_21 & a_39;
assign w1332 = ~w13201 & w13934;
assign w1333 = ~w1585 & ~w5573;
assign w1334 = w4116 & w10590;
assign w1335 = ~a_52 & a_53;
assign w1336 = a_34 & a_41;
assign w1337 = w11301 & w9500;
assign w1338 = a_35 & a_54;
assign w1339 = ~w16160 & ~w15568;
assign w1340 = ~w669 & ~w2410;
assign w1341 = (~w9337 & w1792) | (~w9337 & w9623) | (w1792 & w9623);
assign w1342 = ~w15560 & w19148;
assign w1343 = ~w10733 & w4824;
assign w1344 = w4029 & ~w2448;
assign w1345 = a_0 & a_33;
assign w1346 = ~w3103 & ~w15211;
assign w1347 = w10138 & ~w7163;
assign w1348 = (~w7033 & ~w2173) | (~w7033 & w18066) | (~w2173 & w18066);
assign w1349 = ~w9917 & ~w18824;
assign w1350 = ~w7283 & w11945;
assign w1351 = (~w8097 & ~w5849) | (~w8097 & w16862) | (~w5849 & w16862);
assign w1352 = ~w3622 & ~w1211;
assign w1353 = ~w11202 & ~w12867;
assign w1354 = ~w5482 & ~w14935;
assign w1355 = w5549 & ~w13907;
assign w1356 = w3102 & w4866;
assign w1357 = ~w16097 & w2759;
assign w1358 = w10363 & ~w13101;
assign w1359 = w4585 & ~w10241;
assign w1360 = ~w2172 & ~w18221;
assign w1361 = a_28 & a_38;
assign w1362 = ~w7608 & w4195;
assign w1363 = ~w2161 & ~w8625;
assign w1364 = w18688 & ~w7503;
assign w1365 = w9525 & ~w15327;
assign w1366 = ~w15661 & ~w10480;
assign w1367 = ~w737 & ~w10317;
assign w1368 = ~w8109 & ~w4980;
assign w1369 = a_11 & a_36;
assign w1370 = ~w4896 & ~w12661;
assign w1371 = a_46 & a_51;
assign w1372 = ~w17905 & ~w12626;
assign w1373 = ~w2439 & ~w15721;
assign w1374 = ~w1336 & ~w3140;
assign w1375 = ~w7839 & ~w11285;
assign w1376 = ~w17574 & w6465;
assign w1377 = ~w1771 & ~w7075;
assign w1378 = a_8 & a_37;
assign w1379 = ~w16691 & ~w9601;
assign w1380 = (~w38 & ~w13261) | (~w38 & w12322) | (~w13261 & w12322);
assign w1381 = ~w2008 & ~w12619;
assign w1382 = ~w18293 & ~w7939;
assign w1383 = ~w17438 & w4746;
assign w1384 = w9684 & ~w13335;
assign w1385 = ~w9698 & w1120;
assign w1386 = ~w11958 & ~w14512;
assign w1387 = ~w17451 & ~w13349;
assign w1388 = ~w2341 & ~w16906;
assign w1389 = ~w12046 & ~w12937;
assign w1390 = w1705 & w7561;
assign w1391 = ~w12039 & ~w15380;
assign w1392 = ~w64 & ~w6425;
assign w1393 = a_34 & a_38;
assign w1394 = (~w3908 & w10330) | (~w3908 & w7927) | (w10330 & w7927);
assign w1395 = (w18257 & w11904) | (w18257 & w11856) | (w11904 & w11856);
assign w1396 = w5395 & ~w14905;
assign w1397 = ~w13998 & ~w1534;
assign w1398 = w14841 & w1;
assign w1399 = (w2352 & w13558) | (w2352 & w15399) | (w13558 & w15399);
assign w1400 = ~w7887 & ~w11389;
assign w1401 = (w2342 & w11496) | (w2342 & w206) | (w11496 & w206);
assign w1402 = w10183 & w4424;
assign w1403 = ~w7663 & ~w12073;
assign w1404 = ~w3373 & ~w5737;
assign w1405 = w7074 & ~w7054;
assign w1406 = ~w3319 & w15381;
assign w1407 = ~w17205 & ~w8147;
assign w1408 = a_13 & a_63;
assign w1409 = ~w6485 & ~w4517;
assign w1410 = w694 & w5816;
assign w1411 = ~w13941 & ~w11821;
assign w1412 = w10498 & ~w3094;
assign w1413 = w8612 & w15578;
assign w1414 = w16664 & w14836;
assign w1415 = ~w17152 & ~w13705;
assign w1416 = w8101 & ~w7951;
assign w1417 = w3800 & ~w2389;
assign w1418 = ~w17752 & ~w11222;
assign w1419 = ~w14530 & ~w17173;
assign w1420 = ~w17876 & ~w13890;
assign w1421 = ~w12615 & ~w18032;
assign w1422 = w8763 & ~w12473;
assign w1423 = ~w14201 & w8390;
assign w1424 = (w1320 & w16136) | (w1320 & w7826) | (w16136 & w7826);
assign w1425 = ~w10015 & ~w8363;
assign w1426 = ~w1494 & ~w15923;
assign w1427 = ~w14689 & w6517;
assign w1428 = ~w12556 & ~w1937;
assign w1429 = ~w5 & ~w6217;
assign w1430 = (w5997 & w7659) | (w5997 & w356) | (w7659 & w356);
assign w1431 = ~w12131 & w796;
assign w1432 = (a_1 & w13169) | (a_1 & w14584) | (w13169 & w14584);
assign w1433 = ~w3669 & ~w12405;
assign w1434 = ~w13212 & ~w11063;
assign w1435 = w4141 & ~w18286;
assign w1436 = a_30 & a_42;
assign w1437 = ~w17316 & ~w12563;
assign w1438 = ~w2189 & w1131;
assign w1439 = ~w5369 & ~w17676;
assign w1440 = ~w10614 & w9483;
assign w1441 = a_5 & a_42;
assign w1442 = ~w18829 & w7145;
assign w1443 = ~w5784 & ~w6337;
assign w1444 = a_37 & a_63;
assign w1445 = ~w6811 & w13796;
assign w1446 = w6395 & ~w15766;
assign w1447 = ~w755 & ~w1602;
assign w1448 = ~w730 & ~w428;
assign w1449 = ~w15647 & w4429;
assign w1450 = ~w14384 & w5725;
assign w1451 = ~w9748 & ~w3649;
assign w1452 = ~w12716 & ~w16170;
assign w1453 = w17327 & ~w5585;
assign w1454 = a_18 & a_29;
assign w1455 = ~w13461 & w12647;
assign w1456 = ~w3390 & w3749;
assign w1457 = w7377 & ~w7215;
assign w1458 = ~w4897 & ~w2101;
assign w1459 = ~w5975 & ~w6346;
assign w1460 = w10721 & w14687;
assign w1461 = w5395 & ~w18214;
assign w1462 = ~a_42 & a_43;
assign w1463 = w1299 & ~w17376;
assign w1464 = ~w3244 & ~w15802;
assign w1465 = ~w10107 & ~w11941;
assign w1466 = (w4766 & w7102) | (w4766 & w18741) | (w7102 & w18741);
assign w1467 = ~w11062 & ~w3759;
assign w1468 = ~w2689 & ~w3477;
assign w1469 = (w16423 & w11385) | (w16423 & w10283) | (w11385 & w10283);
assign w1470 = a_12 & a_20;
assign w1471 = ~w10751 & ~w8082;
assign w1472 = w7560 & ~w8272;
assign w1473 = w2243 & w7777;
assign w1474 = ~w5758 & w18252;
assign w1475 = ~w15816 & ~w4835;
assign w1476 = ~w18682 & ~w14718;
assign w1477 = w9819 & ~w8340;
assign w1478 = w19079 & w1796;
assign w1479 = w8853 & w3846;
assign w1480 = ~w15219 & w9534;
assign w1481 = ~w16640 & ~w11302;
assign w1482 = ~w1621 & ~w963;
assign w1483 = ~w11748 & ~w17053;
assign w1484 = ~w7242 & ~w14225;
assign w1485 = w8874 & ~w10690;
assign w1486 = w13125 & w5215;
assign w1487 = ~w10355 & ~w14675;
assign w1488 = ~w3023 & ~w6457;
assign w1489 = ~w4255 & ~w18211;
assign w1490 = a_12 & a_47;
assign w1491 = ~w13027 & ~w16365;
assign w1492 = a_4 & a_40;
assign w1493 = (~w2451 & ~w9904) | (~w2451 & w7332) | (~w9904 & w7332);
assign w1494 = ~w9178 & ~w6569;
assign w1495 = a_34 & a_36;
assign w1496 = ~w3878 & ~w4528;
assign w1497 = w5560 & w16685;
assign w1498 = ~w653 & ~w9063;
assign w1499 = ~w7111 & w12998;
assign w1500 = (~w15566 & ~w15288) | (~w15566 & w3959) | (~w15288 & w3959);
assign w1501 = ~w14628 & w13971;
assign w1502 = ~w7292 & ~w8381;
assign w1503 = (~w11541 & ~w13200) | (~w11541 & w2130) | (~w13200 & w2130);
assign w1504 = ~w254 & w17959;
assign w1505 = ~w12048 & w475;
assign w1506 = (~w17082 & w9963) | (~w17082 & w8210) | (w9963 & w8210);
assign w1507 = ~w8121 & w12082;
assign w1508 = ~w11321 & ~w11819;
assign w1509 = ~w5603 & ~w4402;
assign w1510 = ~w19119 & ~w17769;
assign w1511 = a_7 & a_20;
assign w1512 = ~w18443 & w18143;
assign w1513 = ~w9175 & ~w1029;
assign w1514 = ~w10044 & ~w7574;
assign w1515 = ~w5829 & ~w7173;
assign w1516 = ~w18270 & w8945;
assign w1517 = ~w17076 & ~w3393;
assign w1518 = ~w12091 & ~w4743;
assign w1519 = w18031 & w9507;
assign w1520 = ~w8411 & ~w13107;
assign w1521 = ~w15590 & ~w12384;
assign w1522 = ~w5970 & ~w3412;
assign w1523 = ~w19029 & ~w11509;
assign w1524 = (a_57 & w2227) | (a_57 & w18685) | (w2227 & w18685);
assign w1525 = ~w11549 & ~w3123;
assign w1526 = a_43 & a_55;
assign w1527 = w14668 & ~w7933;
assign w1528 = ~w4375 & w1483;
assign w1529 = ~w2123 & w5063;
assign w1530 = w10363 & w17097;
assign w1531 = ~w14659 & ~w5403;
assign w1532 = ~w7409 & w7780;
assign w1533 = ~w3057 & ~w14498;
assign w1534 = a_10 & a_22;
assign w1535 = w3304 & ~w11371;
assign w1536 = w1961 & w17024;
assign w1537 = ~w1460 & ~w15281;
assign w1538 = w18287 & ~w6773;
assign w1539 = w2608 & w5502;
assign w1540 = (~w2330 & ~w15397) | (~w2330 & w7813) | (~w15397 & w7813);
assign w1541 = w7666 & w11342;
assign w1542 = ~w8439 & w3984;
assign w1543 = ~w2583 & w4584;
assign w1544 = w12745 & ~w9469;
assign w1545 = w11067 & ~w5025;
assign w1546 = a_56 & a_58;
assign w1547 = ~w3113 & ~w6284;
assign w1548 = ~w17185 & w7657;
assign w1549 = ~w9134 & ~w3093;
assign w1550 = ~w16328 & ~w5595;
assign w1551 = ~w9547 & ~w15034;
assign w1552 = ~w15861 & w15159;
assign w1553 = ~w372 & w2960;
assign w1554 = ~w9448 & ~w18081;
assign w1555 = a_14 & a_53;
assign w1556 = w12122 & ~w15430;
assign w1557 = ~w5525 & ~w11799;
assign w1558 = w12625 & w4275;
assign w1559 = ~w3082 & w6975;
assign w1560 = a_13 & a_30;
assign w1561 = ~w5266 & ~w4167;
assign w1562 = ~w6302 & ~w12015;
assign w1563 = ~w7155 & ~w10662;
assign w1564 = ~w16209 & ~w4974;
assign w1565 = ~w2674 & w16617;
assign w1566 = ~w464 & w7338;
assign w1567 = ~w20 & ~w14075;
assign w1568 = ~w13039 & ~w17964;
assign w1569 = ~w18329 & ~w13046;
assign w1570 = ~w2697 & ~w15614;
assign w1571 = w745 & w10441;
assign w1572 = w11440 & ~w12934;
assign w1573 = (~w9354 & w8838) | (~w9354 & w6486) | (w8838 & w6486);
assign w1574 = ~w5778 & ~w16919;
assign w1575 = a_33 & a_51;
assign w1576 = ~w9810 & w19149;
assign w1577 = ~w9200 & ~w6552;
assign w1578 = w13227 & ~w15360;
assign w1579 = ~w4048 & w11740;
assign w1580 = w1137 & ~w9667;
assign w1581 = w13924 & ~w8772;
assign w1582 = w2391 & w3510;
assign w1583 = w14387 & ~w16026;
assign w1584 = ~w14223 & w6380;
assign w1585 = ~w7703 & ~w13655;
assign w1586 = (~w9392 & ~w2408) | (~w9392 & w2815) | (~w2408 & w2815);
assign w1587 = ~w9051 & ~w391;
assign w1588 = ~w13324 & ~w9333;
assign w1589 = ~w9099 & ~w16453;
assign w1590 = ~w15270 & ~w1244;
assign w1591 = ~w16201 & ~w9072;
assign w1592 = (~w8087 & ~w11103) | (~w8087 & w2839) | (~w11103 & w2839);
assign w1593 = w11645 & w19150;
assign w1594 = ~w14814 & ~w4909;
assign w1595 = (w5253 & ~w8987) | (w5253 & w12629) | (~w8987 & w12629);
assign w1596 = (~w152 & w552) | (~w152 & w15675) | (w552 & w15675);
assign w1597 = ~w7475 & ~w18105;
assign w1598 = ~w6766 & ~w1486;
assign w1599 = ~w17475 & ~w4647;
assign w1600 = ~w1194 & ~w17527;
assign w1601 = ~w4828 & ~w18844;
assign w1602 = ~w14383 & ~w7650;
assign w1603 = ~w2360 & ~w7569;
assign w1604 = ~w9307 & ~w21;
assign w1605 = ~w13694 & ~w4064;
assign w1606 = ~w13465 & ~w7167;
assign w1607 = ~w10403 & ~w11811;
assign w1608 = ~w9590 & ~w3927;
assign w1609 = ~w13246 & ~w15803;
assign w1610 = w4635 & w16504;
assign w1611 = ~w11490 & ~w4425;
assign w1612 = w3794 & ~w17385;
assign w1613 = ~w15020 & ~w5093;
assign w1614 = ~w4655 & ~w5029;
assign w1615 = ~w3921 & ~w15314;
assign w1616 = ~w279 & w3876;
assign w1617 = ~w331 & ~w10197;
assign w1618 = ~w10330 & w8691;
assign w1619 = ~w11493 & ~w234;
assign w1620 = w17851 & ~w3906;
assign w1621 = ~w17857 & ~w7070;
assign w1622 = ~w5545 & w11069;
assign w1623 = (~w11668 & ~w2579) | (~w11668 & w7094) | (~w2579 & w7094);
assign w1624 = ~w16631 & ~w16118;
assign w1625 = ~w3557 & ~w13023;
assign w1626 = w3765 & w9894;
assign w1627 = ~w8646 & ~w16993;
assign w1628 = a_0 & a_12;
assign w1629 = ~w4080 & ~w17055;
assign w1630 = ~w8282 & ~w15697;
assign w1631 = w10568 & ~w11851;
assign w1632 = ~w821 & ~w5534;
assign w1633 = a_6 & a_38;
assign w1634 = ~w4356 & ~w13547;
assign w1635 = w2107 & w9276;
assign w1636 = ~w11598 & ~w17917;
assign w1637 = ~w18112 & w10295;
assign w1638 = ~w7129 & w17207;
assign w1639 = ~w18768 & ~w3173;
assign w1640 = ~w12651 & ~w5597;
assign w1641 = ~w14520 & ~w576;
assign w1642 = ~w10470 & w4718;
assign w1643 = ~w5367 & ~w5192;
assign w1644 = w5617 & ~w574;
assign w1645 = ~w14324 & ~w9496;
assign w1646 = w10212 & ~w16689;
assign w1647 = ~w91 & w18727;
assign w1648 = (w3858 & w12973) | (w3858 & w706) | (w12973 & w706);
assign w1649 = w1448 & ~w10468;
assign w1650 = ~w8762 & ~w9307;
assign w1651 = ~w5612 & ~w6105;
assign w1652 = a_28 & a_60;
assign w1653 = w8060 & ~w11613;
assign w1654 = (~w16156 & ~w1061) | (~w16156 & w15229) | (~w1061 & w15229);
assign w1655 = a_17 & a_48;
assign w1656 = ~w12718 & w9487;
assign w1657 = w15519 & ~w2477;
assign w1658 = ~w17558 & ~w16005;
assign w1659 = w15399 & w8722;
assign w1660 = w8655 & ~w4325;
assign w1661 = (~w11877 & ~w6961) | (~w11877 & w7271) | (~w6961 & w7271);
assign w1662 = w7192 & w18589;
assign w1663 = w12492 & ~w10862;
assign w1664 = (w2769 & w3238) | (w2769 & w13810) | (w3238 & w13810);
assign w1665 = ~w5646 & ~w1392;
assign w1666 = w4652 & w5380;
assign w1667 = ~w8715 & ~w9106;
assign w1668 = ~w4696 & ~w5267;
assign w1669 = w9912 & w1830;
assign w1670 = w6701 & w18273;
assign w1671 = a_48 & a_54;
assign w1672 = w11454 & ~w4113;
assign w1673 = (~w17996 & ~w11484) | (~w17996 & w2510) | (~w11484 & w2510);
assign w1674 = ~w3592 & w1380;
assign w1675 = ~w9567 & w5406;
assign w1676 = ~w3421 & ~w11912;
assign w1677 = a_11 & a_33;
assign w1678 = a_27 & a_62;
assign w1679 = a_9 & a_63;
assign w1680 = w15389 & w16745;
assign w1681 = w6081 & ~w12836;
assign w1682 = ~w7074 & ~w16775;
assign w1683 = ~w15374 & w16286;
assign w1684 = ~w9988 & ~w12555;
assign w1685 = w15151 & ~w13737;
assign w1686 = w13373 & ~w14304;
assign w1687 = ~w142 & w10102;
assign w1688 = ~w4631 & ~w9398;
assign w1689 = ~w5641 & ~w1639;
assign w1690 = w13765 & ~w10415;
assign w1691 = ~w14161 & w10122;
assign w1692 = ~w5583 & ~w17823;
assign w1693 = ~w14720 & ~w4112;
assign w1694 = ~w11944 & ~w13798;
assign w1695 = ~w1441 & w7448;
assign w1696 = ~w16967 & ~w5679;
assign w1697 = a_11 & a_18;
assign w1698 = a_42 & a_47;
assign w1699 = ~w9609 & ~w16303;
assign w1700 = a_42 & a_61;
assign w1701 = ~w16746 & ~w10752;
assign w1702 = w3194 & ~w4657;
assign w1703 = ~w14678 & w5061;
assign w1704 = ~w1848 & ~w9109;
assign w1705 = ~w18724 & ~w14421;
assign w1706 = a_26 & a_38;
assign w1707 = w9048 & ~w10009;
assign w1708 = ~w16287 & w14956;
assign w1709 = w7449 & w13566;
assign w1710 = ~w1309 & ~w5762;
assign w1711 = ~w8664 & ~w339;
assign w1712 = w10030 & ~w14230;
assign w1713 = w13186 & w7597;
assign w1714 = ~w7178 & ~w10908;
assign w1715 = ~w11564 & ~w13410;
assign w1716 = ~w12932 & w10762;
assign w1717 = ~w17908 & w15086;
assign w1718 = w13674 & w12112;
assign w1719 = ~w4521 & ~w11869;
assign w1720 = ~w7655 & ~w18338;
assign w1721 = w11973 & ~w15022;
assign w1722 = w14550 & w17274;
assign w1723 = ~w10065 & ~w12740;
assign w1724 = ~w11528 & ~w8030;
assign w1725 = ~w2457 & w15161;
assign w1726 = (~w963 & w6968) | (~w963 & w13979) | (w6968 & w13979);
assign w1727 = ~w2388 & ~w18898;
assign w1728 = ~w3695 & ~w994;
assign w1729 = ~w4477 & w13201;
assign w1730 = ~w5523 & w2549;
assign w1731 = w17821 & ~w637;
assign w1732 = ~w3027 & ~w3013;
assign w1733 = ~w14816 & ~w5449;
assign w1734 = ~w8118 & ~w1703;
assign w1735 = w10475 & w10938;
assign w1736 = ~w15828 & ~w2484;
assign w1737 = a_7 & a_11;
assign w1738 = ~w8797 & ~w5338;
assign w1739 = ~w14308 & w4920;
assign w1740 = ~w16594 & ~w16885;
assign w1741 = ~w13375 & ~w4534;
assign w1742 = a_21 & a_55;
assign w1743 = a_7 & a_10;
assign w1744 = ~w3713 & ~w6258;
assign w1745 = w5562 & ~w11661;
assign w1746 = a_0 & a_44;
assign w1747 = ~w13429 & ~w6196;
assign w1748 = ~w3918 & ~w9737;
assign w1749 = ~w15812 & w8017;
assign w1750 = ~w9956 & ~w4708;
assign w1751 = ~w15105 & ~w7062;
assign w1752 = ~w18447 & w18389;
assign w1753 = w15218 & w14451;
assign w1754 = ~w17786 & ~w9977;
assign w1755 = a_13 & a_55;
assign w1756 = ~w208 & ~w7110;
assign w1757 = ~w3968 & ~w13200;
assign w1758 = ~w17596 & ~w17608;
assign w1759 = ~w3962 & ~w1692;
assign w1760 = w13684 & ~w7627;
assign w1761 = ~w8660 & ~w9029;
assign w1762 = ~w16489 & ~w8063;
assign w1763 = ~w11494 & ~w9445;
assign w1764 = ~w3737 & ~w4923;
assign w1765 = ~w7821 & ~w16027;
assign w1766 = ~w13355 & ~w7486;
assign w1767 = ~w9133 & ~w4861;
assign w1768 = ~w797 & ~w17459;
assign w1769 = ~w7435 & w6743;
assign w1770 = ~w2775 & w1032;
assign w1771 = ~w9943 & w4323;
assign w1772 = (~w7935 & ~w6954) | (~w7935 & w6488) | (~w6954 & w6488);
assign w1773 = ~w14260 & ~w6180;
assign w1774 = w13186 & w9799;
assign w1775 = ~w4703 & w273;
assign w1776 = ~w12671 & ~w7282;
assign w1777 = w16920 & ~w10698;
assign w1778 = ~w17813 & ~w4463;
assign w1779 = w5816 & w1935;
assign w1780 = ~w13826 & ~w5357;
assign w1781 = ~w2714 & w3354;
assign w1782 = w15316 & w12686;
assign w1783 = (~w1036 & w2607) | (~w1036 & w188) | (w2607 & w188);
assign w1784 = ~w246 & ~w8120;
assign w1785 = w5574 & ~w17621;
assign w1786 = ~w4331 & ~w7348;
assign w1787 = ~w10755 & ~w4353;
assign w1788 = ~w1244 & ~w13510;
assign w1789 = a_50 & a_61;
assign w1790 = ~w6815 & ~w10882;
assign w1791 = ~w4637 & ~w8977;
assign w1792 = w9806 & w17457;
assign w1793 = ~w7472 & ~w13613;
assign w1794 = w12719 & ~w11839;
assign w1795 = w12627 & ~w10257;
assign w1796 = ~w3453 & ~w9265;
assign w1797 = w16554 & w15734;
assign w1798 = (w16432 & w19015) | (w16432 & w5106) | (w19015 & w5106);
assign w1799 = w8753 & w15649;
assign w1800 = w15041 & ~w4436;
assign w1801 = ~w6887 & w10924;
assign w1802 = a_4 & a_32;
assign w1803 = w2405 & w9517;
assign w1804 = (~w2769 & w14542) | (~w2769 & w5470) | (w14542 & w5470);
assign w1805 = ~w14052 & ~w16781;
assign w1806 = ~w9071 & ~w3447;
assign w1807 = ~w5619 & ~w3638;
assign w1808 = w14172 & w1413;
assign w1809 = a_4 & a_11;
assign w1810 = ~w1529 & ~w16877;
assign w1811 = ~w4963 & ~w2506;
assign w1812 = ~w18068 & w16057;
assign w1813 = (w14553 & ~w12746) | (w14553 & w13358) | (~w12746 & w13358);
assign w1814 = w14572 & ~w4309;
assign w1815 = w9239 & w12217;
assign w1816 = ~w18427 & ~w8084;
assign w1817 = ~w7129 & w13374;
assign w1818 = ~w532 & ~w12181;
assign w1819 = w14078 & w4706;
assign w1820 = ~w14828 & ~w10040;
assign w1821 = ~w5043 & ~w14890;
assign w1822 = ~w16219 & ~w11847;
assign w1823 = ~w9915 & ~w6924;
assign w1824 = w518 & w4500;
assign w1825 = ~w14310 & ~w13741;
assign w1826 = (w7415 & w8989) | (w7415 & w6821) | (w8989 & w6821);
assign w1827 = ~w10455 & ~w7037;
assign w1828 = ~w13905 & ~w4925;
assign w1829 = w2799 & ~w335;
assign w1830 = ~w13637 & ~w7272;
assign w1831 = ~w107 & w5300;
assign w1832 = ~w7288 & ~w5812;
assign w1833 = w9692 & ~w16496;
assign w1834 = ~w3834 & ~w16665;
assign w1835 = w18950 & w5634;
assign w1836 = ~w293 & ~w16013;
assign w1837 = w1320 & w17036;
assign w1838 = ~w6364 & ~w15056;
assign w1839 = ~w7740 & ~w18706;
assign w1840 = ~w13818 & w3296;
assign w1841 = ~w18496 & w3624;
assign w1842 = (w14976 & w11286) | (w14976 & w11187) | (w11286 & w11187);
assign w1843 = w10464 & w11889;
assign w1844 = (~w13944 & ~w2685) | (~w13944 & w7680) | (~w2685 & w7680);
assign w1845 = ~w7019 & ~w17298;
assign w1846 = w7373 & w16779;
assign w1847 = ~w17978 & ~w11370;
assign w1848 = ~w16800 & ~w8181;
assign w1849 = a_20 & a_51;
assign w1850 = ~w2267 & ~w18586;
assign w1851 = ~w1056 & w6518;
assign w1852 = ~w10593 & ~w16589;
assign w1853 = w8165 & w9400;
assign w1854 = ~w12452 & ~w18577;
assign w1855 = ~w18970 & ~w2313;
assign w1856 = (w18365 & w9092) | (w18365 & w3870) | (w9092 & w3870);
assign w1857 = ~w18082 & ~w8184;
assign w1858 = a_36 & a_42;
assign w1859 = a_6 & a_41;
assign w1860 = ~w11976 & w16423;
assign w1861 = ~w16615 & ~w11085;
assign w1862 = (~w1665 & ~w2270) | (~w1665 & w14158) | (~w2270 & w14158);
assign w1863 = ~w15339 & ~w10013;
assign w1864 = a_16 & a_58;
assign w1865 = (~w12063 & ~w17172) | (~w12063 & w13908) | (~w17172 & w13908);
assign w1866 = w17401 & ~w18115;
assign w1867 = ~w9621 & ~w18854;
assign w1868 = ~w4145 & ~w8338;
assign w1869 = ~w7387 & ~w10117;
assign w1870 = ~w15128 & ~w7974;
assign w1871 = a_28 & a_33;
assign w1872 = ~w11280 & ~w6078;
assign w1873 = a_27 & a_47;
assign w1874 = ~w13642 & ~w14324;
assign w1875 = w4097 & w15657;
assign w1876 = (~w10382 & ~w18272) | (~w10382 & w9151) | (~w18272 & w9151);
assign w1877 = ~w16238 & ~w11442;
assign w1878 = w6381 & w13197;
assign w1879 = ~w7052 & ~w4550;
assign w1880 = ~w12627 & ~w13297;
assign w1881 = ~w8762 & w4664;
assign w1882 = ~w1120 & w18374;
assign w1883 = w14603 & w4946;
assign w1884 = w18165 & w11341;
assign w1885 = w14127 & w2858;
assign w1886 = w2068 & ~w16106;
assign w1887 = (~w5433 & ~w13083) | (~w5433 & w11216) | (~w13083 & w11216);
assign w1888 = w1983 & ~w16638;
assign w1889 = a_42 & a_59;
assign w1890 = a_28 & a_57;
assign w1891 = a_10 & a_13;
assign w1892 = w1182 & w11053;
assign w1893 = ~w7489 & ~w4171;
assign w1894 = ~w6775 & w7009;
assign w1895 = w9328 & ~w5556;
assign w1896 = ~w3135 & ~w974;
assign w1897 = ~w5734 & ~w3550;
assign w1898 = (~w18625 & ~w6399) | (~w18625 & w9108) | (~w6399 & w9108);
assign w1899 = a_23 & a_39;
assign w1900 = w8090 & w16150;
assign w1901 = a_11 & a_26;
assign w1902 = w13408 & ~w2629;
assign w1903 = (~w3376 & ~w1219) | (~w3376 & w991) | (~w1219 & w991);
assign w1904 = a_20 & a_42;
assign w1905 = w15345 & ~w6667;
assign w1906 = ~w1786 & ~w5074;
assign w1907 = w6097 & w2711;
assign w1908 = a_0 & a_30;
assign w1909 = ~w17162 & w9637;
assign w1910 = ~w6216 & ~w2463;
assign w1911 = w7161 & w11168;
assign w1912 = ~w17785 & w13370;
assign w1913 = a_3 & a_62;
assign w1914 = ~w7353 & ~w325;
assign w1915 = w1275 & w16583;
assign w1916 = (w10038 & w6653) | (w10038 & w8112) | (w6653 & w8112);
assign w1917 = ~w4539 & w2523;
assign w1918 = ~w210 & ~w5988;
assign w1919 = ~w12800 & ~w1126;
assign w1920 = ~w1803 & ~w9283;
assign w1921 = ~w2179 & ~w32;
assign w1922 = w7283 & ~w11945;
assign w1923 = ~w11497 & ~w16126;
assign w1924 = ~w11165 & ~w3372;
assign w1925 = w6177 & ~w18425;
assign w1926 = ~w11456 & ~w3896;
assign w1927 = ~w15510 & w16961;
assign w1928 = w18017 & w18216;
assign w1929 = w18486 & ~w8792;
assign w1930 = a_31 & a_39;
assign w1931 = ~w16143 & w12020;
assign w1932 = ~w1054 & w14009;
assign w1933 = w12839 & ~w4541;
assign w1934 = (w14221 & w8635) | (w14221 & w19001) | (w8635 & w19001);
assign w1935 = a_44 & a_55;
assign w1936 = w14015 & ~w5148;
assign w1937 = w8911 & ~w16261;
assign w1938 = (w13854 & w13955) | (w13854 & w3946) | (w13955 & w3946);
assign w1939 = ~w12898 & w3407;
assign w1940 = a_28 & a_50;
assign w1941 = ~w1761 & ~w9736;
assign w1942 = ~w8843 & ~w8545;
assign w1943 = ~w19101 & ~w4247;
assign w1944 = w3915 & ~w10196;
assign w1945 = ~w2089 & w483;
assign w1946 = w2684 & w5028;
assign w1947 = ~w363 & ~w3727;
assign w1948 = ~w11014 & ~w13619;
assign w1949 = ~w2299 & ~w18728;
assign w1950 = w5328 & ~w1415;
assign w1951 = ~w11061 & ~w3185;
assign w1952 = ~w14623 & w9663;
assign w1953 = ~w4833 & w6929;
assign w1954 = ~w13825 & ~w6387;
assign w1955 = ~w6060 & w3060;
assign w1956 = ~w5723 & w9246;
assign w1957 = ~w12896 & ~w1010;
assign w1958 = ~w1699 & ~w17591;
assign w1959 = ~w15915 & w14415;
assign w1960 = ~w13352 & ~w384;
assign w1961 = ~w15681 & ~w311;
assign w1962 = ~w12904 & w13254;
assign w1963 = ~w6031 & w12247;
assign w1964 = (~w477 & ~w18562) | (~w477 & w6308) | (~w18562 & w6308);
assign w1965 = w2012 & w15055;
assign w1966 = (w7243 & w2769) | (w7243 & w889) | (w2769 & w889);
assign w1967 = a_4 & a_51;
assign w1968 = ~w11883 & ~w7972;
assign w1969 = ~w8923 & ~w4525;
assign w1970 = ~w10261 & ~w4374;
assign w1971 = (w18923 & w11686) | (w18923 & w7539) | (w11686 & w7539);
assign w1972 = w11776 & ~w2444;
assign w1973 = w11760 & ~w1000;
assign w1974 = (w7102 & w4341) | (w7102 & w10785) | (w4341 & w10785);
assign w1975 = w14349 & w10328;
assign w1976 = w5558 & w9904;
assign w1977 = w4002 & ~w4337;
assign w1978 = ~w5424 & ~w2320;
assign w1979 = w5179 & w1755;
assign w1980 = a_26 & a_39;
assign w1981 = ~w6986 & ~w15529;
assign w1982 = ~w3645 & w15103;
assign w1983 = a_35 & a_37;
assign w1984 = ~w493 & w8937;
assign w1985 = ~w16954 & w789;
assign w1986 = ~w13082 & w3845;
assign w1987 = w8947 & ~w6865;
assign w1988 = w2202 & w10205;
assign w1989 = ~w13781 & ~w10306;
assign w1990 = (w10122 & w9764) | (w10122 & w3908) | (w9764 & w3908);
assign w1991 = ~w2154 & ~w13966;
assign w1992 = w14014 & w8650;
assign w1993 = ~w411 & ~w9645;
assign w1994 = a_8 & a_25;
assign w1995 = ~w4277 & ~w17567;
assign w1996 = ~w11036 & ~w17559;
assign w1997 = w10981 & w11808;
assign w1998 = ~w18905 & ~w15689;
assign w1999 = (~w16858 & ~w8947) | (~w16858 & w2129) | (~w8947 & w2129);
assign w2000 = ~w7025 & ~w9073;
assign w2001 = ~w4259 & ~w7730;
assign w2002 = (w14255 & w11909) | (w14255 & w16995) | (w11909 & w16995);
assign w2003 = w14620 & w9870;
assign w2004 = ~w6169 & ~w10665;
assign w2005 = a_16 & a_48;
assign w2006 = a_2 & a_53;
assign w2007 = w2189 & ~w1131;
assign w2008 = w269 & ~w10952;
assign w2009 = w13805 & ~w11135;
assign w2010 = a_39 & a_43;
assign w2011 = ~w3141 & ~w18796;
assign w2012 = ~w7514 & ~w2138;
assign w2013 = ~w15247 & w15256;
assign w2014 = ~w7032 & ~w19104;
assign w2015 = w10325 & ~w3620;
assign w2016 = ~w18871 & ~w13614;
assign w2017 = ~w11197 & ~w2509;
assign w2018 = ~w4674 & ~w4271;
assign w2019 = w14216 & ~w10960;
assign w2020 = w12958 & ~w16702;
assign w2021 = ~w3857 & ~w1663;
assign w2022 = ~w6960 & w14685;
assign w2023 = a_29 & a_33;
assign w2024 = w17543 & w2478;
assign w2025 = a_10 & a_31;
assign w2026 = ~w2769 & w8726;
assign w2027 = w15982 & w15832;
assign w2028 = w10503 & w14540;
assign w2029 = a_8 & a_31;
assign w2030 = ~w1753 & ~w2342;
assign w2031 = ~w15207 & ~w4690;
assign w2032 = ~w15694 & w7546;
assign w2033 = a_37 & a_40;
assign w2034 = (~w12290 & ~w6702) | (~w12290 & w9314) | (~w6702 & w9314);
assign w2035 = a_11 & a_25;
assign w2036 = ~w15083 & ~w18320;
assign w2037 = ~w15486 & ~w18406;
assign w2038 = w3341 & ~w13599;
assign w2039 = w9713 & w4927;
assign w2040 = ~w8641 & w143;
assign w2041 = a_18 & a_51;
assign w2042 = ~w11489 & ~w4972;
assign w2043 = ~w10033 & ~w7801;
assign w2044 = ~w15911 & w8347;
assign w2045 = ~w3765 & ~w895;
assign w2046 = w8479 & ~w13194;
assign w2047 = ~w18980 & w17225;
assign w2048 = (~w6977 & ~w12680) | (~w6977 & w3707) | (~w12680 & w3707);
assign w2049 = ~w14503 & ~w1952;
assign w2050 = ~w275 & w2991;
assign w2051 = w1995 & ~w16692;
assign w2052 = (~w9594 & ~w2240) | (~w9594 & w12598) | (~w2240 & w12598);
assign w2053 = (~w16400 & ~w8356) | (~w16400 & w5377) | (~w8356 & w5377);
assign w2054 = w11161 & ~w12640;
assign w2055 = w10107 & w11941;
assign w2056 = a_26 & a_30;
assign w2057 = w5452 & ~w17904;
assign w2058 = ~w10179 & ~w630;
assign w2059 = w17259 & w2971;
assign w2060 = ~w4224 & ~w2528;
assign w2061 = w676 & ~w18563;
assign w2062 = w10518 & w16889;
assign w2063 = ~w859 & ~w12843;
assign w2064 = ~w17765 & w628;
assign w2065 = ~w1257 & ~w10990;
assign w2066 = ~w17840 & w6510;
assign w2067 = (~w13113 & w14329) | (~w13113 & w10982) | (w14329 & w10982);
assign w2068 = a_43 & a_49;
assign w2069 = (w15329 & w1974) | (w15329 & w10099) | (w1974 & w10099);
assign w2070 = ~w5042 & ~w13234;
assign w2071 = ~w18781 & ~w13832;
assign w2072 = ~w12738 & w14791;
assign w2073 = ~w5173 & w9519;
assign w2074 = w290 & w13869;
assign w2075 = a_34 & a_50;
assign w2076 = w4598 & w12758;
assign w2077 = w18996 & ~w16953;
assign w2078 = ~w10320 & ~w2223;
assign w2079 = a_15 & a_30;
assign w2080 = ~w14419 & ~w594;
assign w2081 = ~w18429 & ~w14821;
assign w2082 = ~w16828 & ~w475;
assign w2083 = a_17 & a_60;
assign w2084 = ~w18802 & ~w8321;
assign w2085 = ~w10183 & ~w4424;
assign w2086 = ~w14667 & ~w14605;
assign w2087 = (~w7610 & w6857) | (~w7610 & w16567) | (w6857 & w16567);
assign w2088 = w18407 & w11208;
assign w2089 = ~w15505 & ~w9156;
assign w2090 = w1935 & w8547;
assign w2091 = ~w702 & ~w11751;
assign w2092 = ~w3855 & ~w838;
assign w2093 = ~w11422 & ~w15735;
assign w2094 = a_22 & a_26;
assign w2095 = w7365 & w18104;
assign w2096 = ~w16306 & ~w13185;
assign w2097 = ~w10954 & w8185;
assign w2098 = ~w10683 & ~w16350;
assign w2099 = ~w5015 & ~w18201;
assign w2100 = ~w8778 & ~w14391;
assign w2101 = ~w3821 & ~w11950;
assign w2102 = ~w14074 & ~w12483;
assign w2103 = w4068 & ~w18851;
assign w2104 = (~w1245 & ~w28) | (~w1245 & w13038) | (~w28 & w13038);
assign w2105 = ~w11301 & ~w9500;
assign w2106 = ~w14492 & w16385;
assign w2107 = ~w16499 & ~w19061;
assign w2108 = ~w2002 & ~w2168;
assign w2109 = ~w13637 & ~w4333;
assign w2110 = w3418 & ~w386;
assign w2111 = w8875 & w5586;
assign w2112 = ~w10176 & ~w6775;
assign w2113 = ~w2384 & w536;
assign w2114 = ~w4301 & ~w9664;
assign w2115 = ~w3567 & ~w16293;
assign w2116 = ~w903 & ~w8518;
assign w2117 = w5102 & w8710;
assign w2118 = ~w9016 & w8095;
assign w2119 = w4304 & w3529;
assign w2120 = ~w5703 & ~w17313;
assign w2121 = ~w4312 & w10795;
assign w2122 = ~w8793 & w12444;
assign w2123 = ~w8404 & ~w13616;
assign w2124 = ~w13761 & ~w3214;
assign w2125 = ~w7377 & w7215;
assign w2126 = ~w14546 & ~w3781;
assign w2127 = w15941 & w10193;
assign w2128 = ~w15829 & w8340;
assign w2129 = w6865 & ~w16858;
assign w2130 = ~w3968 & ~w11541;
assign w2131 = ~w15376 & ~w17176;
assign w2132 = w10591 & ~w3672;
assign w2133 = (~w7006 & w11450) | (~w7006 & w5750) | (w11450 & w5750);
assign w2134 = ~w12850 & ~w13954;
assign w2135 = w10315 & w18103;
assign w2136 = ~w9001 & w4275;
assign w2137 = ~w7298 & w16776;
assign w2138 = ~w6423 & ~w5600;
assign w2139 = (~w3292 & ~w5089) | (~w3292 & w5827) | (~w5089 & w5827);
assign w2140 = ~w4084 & ~w13059;
assign w2141 = w15060 & ~w5811;
assign w2142 = ~w5417 & ~w10515;
assign w2143 = ~w11266 & ~w16370;
assign w2144 = ~w10942 & ~w3366;
assign w2145 = ~w3636 & ~w5989;
assign w2146 = ~w9466 & w546;
assign w2147 = ~w7977 & ~w10273;
assign w2148 = ~w1330 & w16349;
assign w2149 = ~w5386 & ~w3657;
assign w2150 = ~w14375 & ~w7518;
assign w2151 = a_1 & a_56;
assign w2152 = ~w13338 & ~w8682;
assign w2153 = ~w752 & ~w12067;
assign w2154 = ~w4383 & ~w12031;
assign w2155 = w8134 & ~w6113;
assign w2156 = ~w17908 & ~w15046;
assign w2157 = w2431 & ~w12360;
assign w2158 = ~w16224 & ~w13485;
assign w2159 = ~w5837 & ~w12733;
assign w2160 = w13016 & ~w5222;
assign w2161 = ~w16144 & w8308;
assign w2162 = ~w15458 & ~w12058;
assign w2163 = a_2 & a_47;
assign w2164 = ~w5682 & ~w5926;
assign w2165 = ~w15389 & ~w16745;
assign w2166 = (~w1805 & ~w10896) | (~w1805 & w19094) | (~w10896 & w19094);
assign w2167 = ~w1963 & ~w16408;
assign w2168 = ~w11388 & w6321;
assign w2169 = a_31 & a_59;
assign w2170 = ~w8500 & ~w2685;
assign w2171 = w12769 & ~w178;
assign w2172 = a_27 & a_55;
assign w2173 = ~w2781 & ~w7033;
assign w2174 = ~w17721 & ~w11784;
assign w2175 = (w7341 & w8154) | (w7341 & w364) | (w8154 & w364);
assign w2176 = ~w15470 & ~w9359;
assign w2177 = ~w9230 & ~w359;
assign w2178 = w4219 & ~w11527;
assign w2179 = w3602 & ~w15708;
assign w2180 = w7830 & ~w15427;
assign w2181 = ~w15204 & ~w15271;
assign w2182 = a_7 & a_47;
assign w2183 = ~w16810 & ~w14923;
assign w2184 = ~w14597 & ~w14155;
assign w2185 = ~w300 & ~w3184;
assign w2186 = ~w18019 & ~w9804;
assign w2187 = w6641 & ~w15033;
assign w2188 = ~w15717 & ~w5537;
assign w2189 = a_12 & a_21;
assign w2190 = ~w15594 & ~w15313;
assign w2191 = ~w8380 & ~w14788;
assign w2192 = ~w18270 & ~w4816;
assign w2193 = a_0 & a_58;
assign w2194 = w15415 & ~w17686;
assign w2195 = ~w5656 & w10652;
assign w2196 = ~w5087 & w4747;
assign w2197 = ~w11548 & ~w7151;
assign w2198 = ~w7307 & ~w8900;
assign w2199 = w5378 & ~w17143;
assign w2200 = ~w15931 & ~w15255;
assign w2201 = ~w8966 & ~w8881;
assign w2202 = ~w15044 & ~w2073;
assign w2203 = ~w2426 & ~w3079;
assign w2204 = ~w16308 & ~w18110;
assign w2205 = w12839 & ~w11320;
assign w2206 = ~w9560 & ~w1189;
assign w2207 = w4184 & w4666;
assign w2208 = ~w18131 & w18178;
assign w2209 = (~w18818 & ~w16018) | (~w18818 & w18506) | (~w16018 & w18506);
assign w2210 = ~w8517 & ~w8002;
assign w2211 = w14087 & ~w2663;
assign w2212 = w13491 & w16777;
assign w2213 = w11105 & w8576;
assign w2214 = ~w6310 & ~w5869;
assign w2215 = ~w4886 & ~w15089;
assign w2216 = w5832 & w7716;
assign w2217 = ~w922 & ~w12174;
assign w2218 = (w19005 & w7366) | (w19005 & w15163) | (w7366 & w15163);
assign w2219 = w1951 & ~w4791;
assign w2220 = a_43 & a_63;
assign w2221 = ~w17648 & ~w6801;
assign w2222 = ~w2530 & ~w207;
assign w2223 = ~w14741 & ~w2375;
assign w2224 = w12987 & ~w2428;
assign w2225 = a_33 & a_37;
assign w2226 = ~w3143 & w8006;
assign w2227 = a_51 & a_62;
assign w2228 = a_29 & a_62;
assign w2229 = ~w6919 & w9065;
assign w2230 = w12334 & ~w296;
assign w2231 = a_8 & a_18;
assign w2232 = ~w2922 & ~w7647;
assign w2233 = w1874 & w17105;
assign w2234 = ~w10490 & ~w15847;
assign w2235 = w14602 & ~w18716;
assign w2236 = ~w8384 & ~w3625;
assign w2237 = a_11 & a_46;
assign w2238 = ~w3560 & w231;
assign w2239 = ~w11748 & w17101;
assign w2240 = ~w9594 & ~w7275;
assign w2241 = ~w2141 & ~w17262;
assign w2242 = ~w17276 & ~w6813;
assign w2243 = ~w10165 & ~w12408;
assign w2244 = (~w4580 & ~w5311) | (~w4580 & w7540) | (~w5311 & w7540);
assign w2245 = ~w8611 & ~w9725;
assign w2246 = a_35 & a_41;
assign w2247 = w13851 & ~w18117;
assign w2248 = ~w3641 & ~w1524;
assign w2249 = a_1 & a_30;
assign w2250 = w10053 & ~w5608;
assign w2251 = ~w16853 & ~w17609;
assign w2252 = w1127 & ~w18883;
assign w2253 = ~w11678 & ~w15171;
assign w2254 = (w9821 & ~w10803) | (w9821 & w7466) | (~w10803 & w7466);
assign w2255 = ~w4869 & ~w18635;
assign w2256 = ~w14201 & ~w3509;
assign w2257 = w15584 & ~w14284;
assign w2258 = w11177 & ~w19064;
assign w2259 = ~w15629 & w8128;
assign w2260 = ~w11060 & ~w4720;
assign w2261 = w9604 & ~w7162;
assign w2262 = w14465 & w1320;
assign w2263 = ~w3920 & w15522;
assign w2264 = ~w1819 & ~w333;
assign w2265 = ~w6961 & ~w13470;
assign w2266 = ~w5214 & ~w3408;
assign w2267 = w14447 & w1318;
assign w2268 = ~w11413 & w18444;
assign w2269 = ~w5850 & ~w16079;
assign w2270 = ~w1665 & ~w14774;
assign w2271 = w9482 & ~w14580;
assign w2272 = ~w15387 & ~w14772;
assign w2273 = ~w7175 & ~w7342;
assign w2274 = (~w8353 & ~w15501) | (~w8353 & w13703) | (~w15501 & w13703);
assign w2275 = (~w18545 & ~w3805) | (~w18545 & w3890) | (~w3805 & w3890);
assign w2276 = w13807 & w5393;
assign w2277 = ~w18065 & ~w14116;
assign w2278 = ~w10552 & ~w6143;
assign w2279 = ~w2836 & w127;
assign w2280 = ~w16690 & ~w15907;
assign w2281 = ~w15913 & ~w14963;
assign w2282 = ~w14727 & ~w12070;
assign w2283 = ~w18289 & ~w15555;
assign w2284 = ~w12022 & ~w11759;
assign w2285 = ~w12501 & w12402;
assign w2286 = ~w18190 & ~w8023;
assign w2287 = a_28 & a_40;
assign w2288 = ~w350 & ~w8926;
assign w2289 = ~w14668 & w7933;
assign w2290 = ~w8701 & w5626;
assign w2291 = ~w11324 & ~w9944;
assign w2292 = w565 & ~w7461;
assign w2293 = w11362 & w5119;
assign w2294 = ~w5788 & ~w19075;
assign w2295 = a_11 & a_19;
assign w2296 = ~w15785 & ~w15943;
assign w2297 = w7915 & ~w5143;
assign w2298 = w10724 & w17862;
assign w2299 = ~w2764 & ~w15177;
assign w2300 = ~w15268 & ~w1161;
assign w2301 = ~w16359 & ~w12754;
assign w2302 = a_33 & a_39;
assign w2303 = ~w18963 & ~w3118;
assign w2304 = a_7 & a_36;
assign w2305 = w6216 & w3418;
assign w2306 = ~w13352 & ~w11052;
assign w2307 = ~w7853 & ~w18196;
assign w2308 = a_45 & a_60;
assign w2309 = ~w12209 & ~w10565;
assign w2310 = w11582 & w8189;
assign w2311 = w107 & ~w5300;
assign w2312 = ~w2349 & ~w16770;
assign w2313 = w250 & w9421;
assign w2314 = ~w11997 & ~w19126;
assign w2315 = w12343 & ~w14417;
assign w2316 = ~w7389 & ~w8773;
assign w2317 = ~w16448 & w8864;
assign w2318 = ~w17360 & w7075;
assign w2319 = a_15 & a_21;
assign w2320 = a_30 & a_34;
assign w2321 = ~w7050 & ~w15869;
assign w2322 = ~w12865 & ~w4253;
assign w2323 = ~w2271 & ~w2567;
assign w2324 = ~w17578 & ~w18836;
assign w2325 = ~w15782 & w1324;
assign w2326 = w18246 & w11289;
assign w2327 = w16741 & ~w10650;
assign w2328 = a_4 & a_33;
assign w2329 = ~w7178 & ~w8775;
assign w2330 = ~w7513 & ~w17436;
assign w2331 = w15245 & ~w9735;
assign w2332 = w2949 & ~w12299;
assign w2333 = ~w10225 & ~w5573;
assign w2334 = w11577 & ~w16500;
assign w2335 = ~w17471 & ~w14276;
assign w2336 = w5874 & w7227;
assign w2337 = w9616 & w14664;
assign w2338 = w13971 & w4966;
assign w2339 = ~w10899 & ~w9460;
assign w2340 = ~w15048 & w13063;
assign w2341 = (~w11651 & w10072) | (~w11651 & w2634) | (w10072 & w2634);
assign w2342 = a_30 & a_61;
assign w2343 = ~w3409 & ~w8617;
assign w2344 = w2401 & w1157;
assign w2345 = ~w1988 & ~w2511;
assign w2346 = ~w3396 & ~w12575;
assign w2347 = ~w18587 & ~w1985;
assign w2348 = ~w11710 & ~w9382;
assign w2349 = w330 & ~w12092;
assign w2350 = w9579 & w19046;
assign w2351 = ~w2834 & ~w15150;
assign w2352 = w18170 & w8135;
assign w2353 = a_19 & a_38;
assign w2354 = ~w8848 & w16212;
assign w2355 = ~w8106 & ~w17415;
assign w2356 = ~w15715 & w1636;
assign w2357 = ~w830 & ~w5282;
assign w2358 = ~w12077 & ~w18711;
assign w2359 = a_32 & a_50;
assign w2360 = w1629 & w14481;
assign w2361 = ~w9695 & w2615;
assign w2362 = w18899 & w5169;
assign w2363 = ~w6906 & ~w820;
assign w2364 = ~w15182 & w13235;
assign w2365 = w306 & w15085;
assign w2366 = ~w5352 & ~w6897;
assign w2367 = ~w16704 & ~w12493;
assign w2368 = ~w14407 & ~w819;
assign w2369 = ~w7201 & ~w4189;
assign w2370 = ~w10632 & ~w12580;
assign w2371 = w17521 & ~w922;
assign w2372 = ~w8343 & ~w8108;
assign w2373 = ~w19103 & ~w18452;
assign w2374 = ~w1883 & ~w11618;
assign w2375 = ~w11503 & w18414;
assign w2376 = w16912 & ~w12638;
assign w2377 = ~w7877 & w3394;
assign w2378 = (~w12335 & ~w1182) | (~w12335 & w2412) | (~w1182 & w2412);
assign w2379 = a_19 & a_20;
assign w2380 = ~w12796 & w12926;
assign w2381 = ~w15912 & ~w1695;
assign w2382 = w7754 & ~w16913;
assign w2383 = ~w11574 & w1242;
assign w2384 = ~w15758 & ~w14489;
assign w2385 = ~w14599 & ~w230;
assign w2386 = w12739 & w15322;
assign w2387 = a_6 & a_24;
assign w2388 = a_14 & a_40;
assign w2389 = ~w14913 & ~w15476;
assign w2390 = w10340 & w11708;
assign w2391 = ~w192 & ~w10672;
assign w2392 = ~w12164 & ~w3058;
assign w2393 = ~w2378 & w6637;
assign w2394 = w10285 & ~w8573;
assign w2395 = w4074 & w3722;
assign w2396 = ~w11447 & ~w11420;
assign w2397 = ~w17248 & ~w14203;
assign w2398 = ~w15349 & ~w2186;
assign w2399 = ~w11742 & w1576;
assign w2400 = ~w464 & ~w12682;
assign w2401 = a_8 & a_48;
assign w2402 = w142 & ~w10102;
assign w2403 = ~w8685 & ~w14107;
assign w2404 = w19018 & w13196;
assign w2405 = (~w3781 & ~w17167) | (~w3781 & w2126) | (~w17167 & w2126);
assign w2406 = ~w11858 & ~w17798;
assign w2407 = ~w17340 & ~w8894;
assign w2408 = ~w9392 & ~w18515;
assign w2409 = w5544 & ~w12028;
assign w2410 = w16703 & w18037;
assign w2411 = ~w6245 & ~w18875;
assign w2412 = ~w11053 & ~w12335;
assign w2413 = ~w18883 & ~w18415;
assign w2414 = ~w15830 & ~w5872;
assign w2415 = ~w18362 & ~w10341;
assign w2416 = w18985 & ~w14932;
assign w2417 = ~w12163 & ~w819;
assign w2418 = a_33 & a_40;
assign w2419 = a_25 & a_38;
assign w2420 = a_5 & a_60;
assign w2421 = (w18650 & w15787) | (w18650 & w3740) | (w15787 & w3740);
assign w2422 = ~w16485 & ~w15266;
assign w2423 = ~w9389 & ~w9436;
assign w2424 = ~w15227 & w4777;
assign w2425 = w9513 & ~w5261;
assign w2426 = ~w3409 & ~w14454;
assign w2427 = ~w7614 & ~w12220;
assign w2428 = ~w4028 & ~w5868;
assign w2429 = ~w117 & w6790;
assign w2430 = w7435 & ~w6743;
assign w2431 = a_4 & a_19;
assign w2432 = ~w280 & ~w5685;
assign w2433 = w2905 & ~w10815;
assign w2434 = ~w14387 & w16026;
assign w2435 = ~w7169 & ~w16314;
assign w2436 = w12262 & w3683;
assign w2437 = w6820 & w15797;
assign w2438 = ~w7701 & w16606;
assign w2439 = a_47 & a_51;
assign w2440 = ~w6609 & ~w1380;
assign w2441 = ~w3487 & ~w14663;
assign w2442 = ~w12859 & ~w3767;
assign w2443 = w12622 & w16172;
assign w2444 = ~w5635 & ~w8248;
assign w2445 = (~w4917 & ~w8252) | (~w4917 & w11968) | (~w8252 & w11968);
assign w2446 = ~w7815 & ~w9647;
assign w2447 = ~w6844 & ~w2203;
assign w2448 = ~w11093 & ~w1113;
assign w2449 = a_42 & a_44;
assign w2450 = ~w941 & ~w15347;
assign w2451 = w4650 & w13266;
assign w2452 = ~w4262 & ~w14807;
assign w2453 = ~w15149 & w4785;
assign w2454 = (w1566 & w13904) | (w1566 & w13872) | (w13904 & w13872);
assign w2455 = w557 & ~w4489;
assign w2456 = w12485 & ~w5394;
assign w2457 = a_13 & a_48;
assign w2458 = ~w14082 & ~w17477;
assign w2459 = ~w13454 & ~w8490;
assign w2460 = (~w10735 & w10875) | (~w10735 & w9541) | (w10875 & w9541);
assign w2461 = w2221 & ~w13828;
assign w2462 = ~w3777 & w14656;
assign w2463 = a_27 & a_42;
assign w2464 = ~w14521 & ~w5113;
assign w2465 = ~w1709 & ~w9138;
assign w2466 = ~w15293 & ~w5843;
assign w2467 = ~w3585 & ~w7474;
assign w2468 = ~w7181 & ~w17808;
assign w2469 = a_16 & a_19;
assign w2470 = ~w225 & ~w5457;
assign w2471 = w13072 & w1339;
assign w2472 = w420 & ~w16778;
assign w2473 = ~w7305 & w13577;
assign w2474 = w7114 & ~w7842;
assign w2475 = ~w2916 & w1838;
assign w2476 = ~w10606 & ~w6991;
assign w2477 = ~w16990 & ~w12145;
assign w2478 = (~w15461 & ~w5808) | (~w15461 & w9377) | (~w5808 & w9377);
assign w2479 = a_8 & a_41;
assign w2480 = w17031 & w13253;
assign w2481 = ~w5412 & ~w16806;
assign w2482 = ~w2394 & ~w10864;
assign w2483 = (w9902 & w10330) | (w9902 & w11697) | (w10330 & w11697);
assign w2484 = ~w13164 & w17535;
assign w2485 = ~w15821 & ~w9456;
assign w2486 = w9631 & w11217;
assign w2487 = w13559 & w4910;
assign w2488 = ~w10902 & ~w1720;
assign w2489 = w9625 & w7084;
assign w2490 = ~w7689 & w2347;
assign w2491 = ~w5422 & ~w6804;
assign w2492 = ~w10663 & w13523;
assign w2493 = ~w18975 & ~w11396;
assign w2494 = a_12 & a_30;
assign w2495 = w5683 & w12762;
assign w2496 = w2154 & w13966;
assign w2497 = w1845 & ~w5745;
assign w2498 = w9580 & ~w824;
assign w2499 = (~w5714 & w12041) | (~w5714 & w15436) | (w12041 & w15436);
assign w2500 = w17052 & ~w10450;
assign w2501 = w17452 & w11293;
assign w2502 = ~w16165 & ~w11566;
assign w2503 = w2968 & ~w2435;
assign w2504 = a_11 & a_49;
assign w2505 = ~w562 & ~w18652;
assign w2506 = w8878 & ~w8393;
assign w2507 = ~w11933 & ~w9401;
assign w2508 = w10699 & w8294;
assign w2509 = ~w13404 & ~w6223;
assign w2510 = w10 & ~w17996;
assign w2511 = ~w2202 & ~w10205;
assign w2512 = a_32 & a_57;
assign w2513 = a_11 & a_43;
assign w2514 = ~w11313 & w12728;
assign w2515 = ~w5530 & w3784;
assign w2516 = a_2 & a_14;
assign w2517 = ~w12973 & w11430;
assign w2518 = w6458 & w5009;
assign w2519 = ~w4702 & w15158;
assign w2520 = (w7253 & w2769) | (w7253 & w12327) | (w2769 & w12327);
assign w2521 = ~w11616 & ~w16374;
assign w2522 = w16998 & ~w1711;
assign w2523 = ~w17937 & ~w7672;
assign w2524 = ~w11660 & ~w520;
assign w2525 = ~w6633 & ~w10303;
assign w2526 = (w8780 & w5527) | (w8780 & w12383) | (w5527 & w12383);
assign w2527 = w1890 & w792;
assign w2528 = w1301 & ~w4217;
assign w2529 = ~w9028 & ~w15939;
assign w2530 = ~a_34 & ~w18850;
assign w2531 = a_6 & a_32;
assign w2532 = a_17 & a_54;
assign w2533 = a_3 & a_14;
assign w2534 = w7899 & ~w2065;
assign w2535 = w2450 & ~w18200;
assign w2536 = ~w7961 & ~w1260;
assign w2537 = ~w5909 & ~w12890;
assign w2538 = w4535 & ~w17399;
assign w2539 = ~w10693 & w4111;
assign w2540 = ~w12876 & ~w138;
assign w2541 = ~w19097 & ~w19001;
assign w2542 = ~w14145 & ~w1634;
assign w2543 = ~w5125 & ~w15608;
assign w2544 = w8417 & ~w16823;
assign w2545 = w14383 & ~w6354;
assign w2546 = ~w16070 & ~w7683;
assign w2547 = a_34 & a_48;
assign w2548 = ~w12428 & ~w11998;
assign w2549 = ~w9930 & ~w4263;
assign w2550 = w8324 & w16845;
assign w2551 = w9691 & ~w7072;
assign w2552 = ~w4558 & w7479;
assign w2553 = ~w1563 & ~w215;
assign w2554 = w8552 & ~w4361;
assign w2555 = w7106 & w14197;
assign w2556 = ~w5955 & ~w13363;
assign w2557 = a_25 & a_52;
assign w2558 = ~w13803 & ~w15298;
assign w2559 = ~w17933 & ~w9083;
assign w2560 = w11141 & ~w3999;
assign w2561 = w2838 & ~w3339;
assign w2562 = ~w17679 & ~w615;
assign w2563 = a_42 & a_63;
assign w2564 = ~w13594 & ~w18035;
assign w2565 = w12100 & ~w5967;
assign w2566 = ~w10114 & ~w8452;
assign w2567 = ~w9482 & w14580;
assign w2568 = w6363 & ~w4769;
assign w2569 = ~w1710 & ~w4806;
assign w2570 = ~w5670 & ~w8037;
assign w2571 = ~w17819 & ~w16712;
assign w2572 = ~w3610 & ~w14089;
assign w2573 = a_37 & a_41;
assign w2574 = ~w10289 & ~w554;
assign w2575 = ~w4194 & ~w9756;
assign w2576 = ~w13147 & ~w5414;
assign w2577 = ~w15237 & ~w3283;
assign w2578 = w11601 & ~w6626;
assign w2579 = ~w11668 & ~w14673;
assign w2580 = ~w12676 & ~w5730;
assign w2581 = w5871 & w13438;
assign w2582 = ~w2684 & ~w5028;
assign w2583 = a_45 & a_54;
assign w2584 = ~w8839 & ~w17916;
assign w2585 = ~w16465 & w9798;
assign w2586 = w2689 & w3477;
assign w2587 = w5226 & ~w426;
assign w2588 = ~w1369 & ~w7372;
assign w2589 = ~w17418 & w14957;
assign w2590 = ~w17160 & ~w6746;
assign w2591 = ~w4052 & ~w12185;
assign w2592 = ~w15854 & ~w4403;
assign w2593 = ~w7498 & ~w8542;
assign w2594 = w321 & ~w6622;
assign w2595 = (~w16896 & w18006) | (~w16896 & w4312) | (w18006 & w4312);
assign w2596 = w4228 & w16346;
assign w2597 = w4871 & ~w12210;
assign w2598 = ~w17173 & ~w12625;
assign w2599 = w7148 & ~w13695;
assign w2600 = ~w5984 & ~w17911;
assign w2601 = a_53 & a_61;
assign w2602 = w350 & w8926;
assign w2603 = ~w8213 & ~w2597;
assign w2604 = ~w16051 & ~w3497;
assign w2605 = ~w10421 & ~w13431;
assign w2606 = ~w12715 & ~w2462;
assign w2607 = (w14993 & w7610) | (w14993 & w14707) | (w7610 & w14707);
assign w2608 = (~w15766 & ~w11536) | (~w15766 & w1446) | (~w11536 & w1446);
assign w2609 = ~w2046 & ~w13731;
assign w2610 = ~w7527 & ~w13517;
assign w2611 = ~w14277 & ~w3020;
assign w2612 = w8886 & w11921;
assign w2613 = ~w2359 & w4851;
assign w2614 = ~w7788 & ~w6467;
assign w2615 = w16072 & w15575;
assign w2616 = a_0 & a_26;
assign w2617 = ~w6996 & ~w3434;
assign w2618 = ~w4968 & ~w15354;
assign w2619 = w11606 & w11155;
assign w2620 = ~w113 & ~w18730;
assign w2621 = ~w2593 & w17367;
assign w2622 = ~w12372 & ~w8575;
assign w2623 = ~w7209 & ~w2869;
assign w2624 = ~w18344 & ~w6015;
assign w2625 = a_8 & a_27;
assign w2626 = ~w1068 & ~w14889;
assign w2627 = ~w11127 & ~w10592;
assign w2628 = w1294 & ~w12541;
assign w2629 = ~w14851 & ~w9862;
assign w2630 = ~w523 & ~w435;
assign w2631 = ~w6289 & w8696;
assign w2632 = ~w7836 & ~w4899;
assign w2633 = ~w10888 & w14017;
assign w2634 = w5360 & ~w11651;
assign w2635 = ~w3006 & ~w13893;
assign w2636 = ~w11736 & ~w10506;
assign w2637 = ~w13742 & ~w5947;
assign w2638 = w4027 & w18289;
assign w2639 = w4750 & ~w13439;
assign w2640 = ~w5105 & w16869;
assign w2641 = ~w10083 & ~w18897;
assign w2642 = ~w17356 & ~w2071;
assign w2643 = ~w6483 & ~w3270;
assign w2644 = w15035 & w6320;
assign w2645 = w6214 & w13981;
assign w2646 = a_12 & a_52;
assign w2647 = w16071 & w11133;
assign w2648 = ~w2193 & ~w13587;
assign w2649 = ~w3950 & ~w6838;
assign w2650 = w4369 & w885;
assign w2651 = ~w10712 & ~w18673;
assign w2652 = ~w7851 & ~w8172;
assign w2653 = w7929 & ~w13171;
assign w2654 = ~w9419 & ~w1854;
assign w2655 = ~w10052 & ~w6560;
assign w2656 = ~w3075 & w2852;
assign w2657 = ~w4627 & ~w11257;
assign w2658 = w11601 & ~w18770;
assign w2659 = ~a_61 & a_62;
assign w2660 = ~w7047 & ~w9080;
assign w2661 = ~w9430 & w13934;
assign w2662 = a_3 & a_18;
assign w2663 = ~w8936 & ~w18383;
assign w2664 = ~w3016 & ~w17002;
assign w2665 = ~w14372 & ~w2662;
assign w2666 = ~w9779 & ~w5521;
assign w2667 = ~w15396 & ~w17677;
assign w2668 = w14239 & w3092;
assign w2669 = w5216 & ~w7976;
assign w2670 = ~w14453 & ~w13171;
assign w2671 = ~w10639 & ~w5923;
assign w2672 = w10542 & ~w1311;
assign w2673 = ~w8786 & w7814;
assign w2674 = ~w8885 & ~w18951;
assign w2675 = ~w6904 & ~w10928;
assign w2676 = (w6359 & ~w5464) | (w6359 & w3828) | (~w5464 & w3828);
assign w2677 = ~w5592 & w642;
assign w2678 = ~w13607 & ~w8266;
assign w2679 = w17963 & ~w18435;
assign w2680 = (w6323 & w10653) | (w6323 & w17517) | (w10653 & w17517);
assign w2681 = ~w7485 & ~w2276;
assign w2682 = ~w18528 & ~w5207;
assign w2683 = w17034 & ~w7196;
assign w2684 = (~w11575 & ~w9526) | (~w11575 & w4007) | (~w9526 & w4007);
assign w2685 = ~w13944 & ~w18881;
assign w2686 = ~w16515 & ~w6292;
assign w2687 = ~w6905 & ~w17247;
assign w2688 = w1661 & ~w17674;
assign w2689 = (~w9667 & ~w227) | (~w9667 & w1580) | (~w227 & w1580);
assign w2690 = ~w6128 & ~w14690;
assign w2691 = a_16 & ~w2249;
assign w2692 = ~w3169 & ~w8563;
assign w2693 = w18236 & w6792;
assign w2694 = ~w18601 & w6524;
assign w2695 = w3650 & w6508;
assign w2696 = w6523 & w17391;
assign w2697 = ~w16475 & ~w5133;
assign w2698 = ~w209 & w11911;
assign w2699 = ~w8530 & ~w1606;
assign w2700 = ~w2190 & ~w14219;
assign w2701 = w15182 & ~w13235;
assign w2702 = ~w425 & ~w13721;
assign w2703 = a_12 & a_44;
assign w2704 = w1574 & ~w315;
assign w2705 = ~w12739 & ~w584;
assign w2706 = (~w13784 & ~w5661) | (~w13784 & w14855) | (~w5661 & w14855);
assign w2707 = ~w18974 & ~w3395;
assign w2708 = ~w18924 & ~w164;
assign w2709 = (~w5527 & w18006) | (~w5527 & w7772) | (w18006 & w7772);
assign w2710 = a_19 & a_33;
assign w2711 = a_24 & a_56;
assign w2712 = ~w4029 & w2448;
assign w2713 = ~w12463 & ~w18241;
assign w2714 = a_28 & a_54;
assign w2715 = w6200 & ~w6353;
assign w2716 = (~w2165 & ~w10623) | (~w2165 & w10637) | (~w10623 & w10637);
assign w2717 = ~w16948 & w6953;
assign w2718 = w12678 & ~w18539;
assign w2719 = ~w9110 & ~w4785;
assign w2720 = w17634 & w10404;
assign w2721 = w11935 & w2792;
assign w2722 = w11154 & ~w1471;
assign w2723 = ~w216 & ~w11633;
assign w2724 = ~w5832 & ~w7716;
assign w2725 = a_2 & a_46;
assign w2726 = w10049 & ~w3131;
assign w2727 = ~w14034 & ~w6981;
assign w2728 = ~w17282 & w10347;
assign w2729 = ~w11996 & ~w9214;
assign w2730 = (w7341 & w11245) | (w7341 & w12280) | (w11245 & w12280);
assign w2731 = w8668 & ~w5864;
assign w2732 = ~w15265 & ~w16672;
assign w2733 = ~w18602 & ~w1498;
assign w2734 = (w14519 & w2769) | (w14519 & w4958) | (w2769 & w4958);
assign w2735 = ~w13075 & ~w8561;
assign w2736 = ~w14724 & ~w11473;
assign w2737 = w9913 & ~w4730;
assign w2738 = ~w14150 & ~w12580;
assign w2739 = w11483 & ~w16203;
assign w2740 = w7361 & ~w13392;
assign w2741 = ~w3080 & ~w8020;
assign w2742 = ~w18522 & ~w11611;
assign w2743 = ~w12203 & ~w18519;
assign w2744 = ~w12781 & w9984;
assign w2745 = w187 & ~w17980;
assign w2746 = a_40 & a_63;
assign w2747 = ~w3610 & ~w13387;
assign w2748 = w4944 & ~w8151;
assign w2749 = ~w5722 & ~w14808;
assign w2750 = ~w9515 & ~w18956;
assign w2751 = w11973 & ~w6819;
assign w2752 = ~w7195 & ~w3177;
assign w2753 = ~w14622 & w9526;
assign w2754 = w3405 & ~w1611;
assign w2755 = ~w11781 & ~w3332;
assign w2756 = ~w8319 & w9281;
assign w2757 = a_7 & a_48;
assign w2758 = ~w1261 & ~w10156;
assign w2759 = ~w15900 & ~w7573;
assign w2760 = ~w8889 & ~w14952;
assign w2761 = ~w11514 & w2357;
assign w2762 = ~w17047 & ~w9426;
assign w2763 = w15030 & ~w14287;
assign w2764 = a_4 & a_43;
assign w2765 = w13347 & w7818;
assign w2766 = (~w11945 & w6325) | (~w11945 & w1922) | (w6325 & w1922);
assign w2767 = a_34 & a_54;
assign w2768 = w17757 & ~w12245;
assign w2769 = ~w2896 & w2994;
assign w2770 = ~w3544 & ~w6210;
assign w2771 = ~w11867 & ~w14643;
assign w2772 = (~w11263 & ~w15041) | (~w11263 & w179) | (~w15041 & w179);
assign w2773 = ~w11080 & w5344;
assign w2774 = ~w4891 & ~w14065;
assign w2775 = a_3 & a_24;
assign w2776 = ~w6548 & ~w6478;
assign w2777 = ~w10909 & w3138;
assign w2778 = ~w12874 & ~w8522;
assign w2779 = ~w13248 & w16270;
assign w2780 = ~w13695 & ~w14215;
assign w2781 = ~w5631 & w13211;
assign w2782 = w8054 & ~w4395;
assign w2783 = ~w11562 & ~w7993;
assign w2784 = ~w19102 & w11243;
assign w2785 = ~w8323 & w10189;
assign w2786 = ~w8453 & w11507;
assign w2787 = ~w551 & w9210;
assign w2788 = w2201 & ~w5597;
assign w2789 = ~w16074 & ~w5959;
assign w2790 = ~w3847 & ~w232;
assign w2791 = ~w16988 & ~w3299;
assign w2792 = a_25 & a_35;
assign w2793 = (~w11227 & ~w12411) | (~w11227 & w14991) | (~w12411 & w14991);
assign w2794 = ~w8985 & ~w11994;
assign w2795 = ~w11134 & ~w5759;
assign w2796 = ~w15528 & ~w9123;
assign w2797 = ~w3083 & ~w8396;
assign w2798 = ~w2073 & ~w460;
assign w2799 = a_13 & a_46;
assign w2800 = w12861 & w7297;
assign w2801 = ~w19073 & ~w7611;
assign w2802 = a_11 & a_41;
assign w2803 = w13082 & w10961;
assign w2804 = w8069 & w16098;
assign w2805 = w8937 & ~w6477;
assign w2806 = ~w4346 & ~w12246;
assign w2807 = a_13 & a_20;
assign w2808 = w91 & w9607;
assign w2809 = w2048 & ~w18370;
assign w2810 = ~w5551 & ~w14078;
assign w2811 = ~w9142 & ~w11302;
assign w2812 = ~w291 & ~w2303;
assign w2813 = ~w982 & ~w1200;
assign w2814 = w1019 & ~w16772;
assign w2815 = ~w7816 & ~w9392;
assign w2816 = ~w7688 & ~w17417;
assign w2817 = ~w17173 & w8442;
assign w2818 = w18203 & w1088;
assign w2819 = ~w12594 & w731;
assign w2820 = w6777 & ~w15253;
assign w2821 = ~w10386 & ~w17194;
assign w2822 = ~w7161 & ~w11168;
assign w2823 = ~w6855 & w13456;
assign w2824 = w1906 & ~w7341;
assign w2825 = w4753 & ~w4570;
assign w2826 = ~w7732 & w18664;
assign w2827 = ~w11158 & ~w18532;
assign w2828 = w3658 & ~w1382;
assign w2829 = ~w8306 & w6644;
assign w2830 = a_7 & a_12;
assign w2831 = ~w2217 & w17521;
assign w2832 = (w15415 & w12741) | (w15415 & w4447) | (w12741 & w4447);
assign w2833 = ~w18 & ~w13535;
assign w2834 = ~w10731 & ~w6810;
assign w2835 = ~w8060 & ~w872;
assign w2836 = ~w17045 & ~w3764;
assign w2837 = a_9 & a_49;
assign w2838 = a_52 & a_59;
assign w2839 = w2312 & ~w8087;
assign w2840 = ~w17017 & w17617;
assign w2841 = w11683 & ~w13462;
assign w2842 = ~w6189 & ~w5030;
assign w2843 = a_10 & a_34;
assign w2844 = ~w14739 & ~w9153;
assign w2845 = ~w8125 & ~w9227;
assign w2846 = ~w13861 & ~w18813;
assign w2847 = (~w12833 & ~w12134) | (~w12833 & w6270) | (~w12134 & w6270);
assign w2848 = ~w13362 & ~w18126;
assign w2849 = ~w5548 & w12733;
assign w2850 = ~w2842 & ~w13727;
assign w2851 = w17685 & w16250;
assign w2852 = ~w6062 & ~w8105;
assign w2853 = w2420 & ~w1557;
assign w2854 = w12459 & w18782;
assign w2855 = ~w12808 & ~w25;
assign w2856 = ~w12150 & w9326;
assign w2857 = ~w18020 & ~w12051;
assign w2858 = a_2 & a_4;
assign w2859 = a_45 & a_61;
assign w2860 = (~w14600 & ~w15204) | (~w14600 & w3623) | (~w15204 & w3623);
assign w2861 = a_37 & a_58;
assign w2862 = ~w15104 & ~w8355;
assign w2863 = ~w11088 & ~w2250;
assign w2864 = ~w9656 & w15240;
assign w2865 = ~w16009 & ~w1374;
assign w2866 = ~w18284 & ~w1427;
assign w2867 = ~w10773 & w13098;
assign w2868 = a_12 & a_34;
assign w2869 = ~w7249 & w1316;
assign w2870 = ~w8052 & ~w7673;
assign w2871 = ~w12946 & ~w16834;
assign w2872 = ~w10393 & ~w4648;
assign w2873 = ~w18981 & ~w14476;
assign w2874 = w18245 & ~w4742;
assign w2875 = ~w12001 & ~w588;
assign w2876 = a_19 & a_58;
assign w2877 = ~w13064 & ~w4142;
assign w2878 = a_45 & a_62;
assign w2879 = ~w4122 & ~w2208;
assign w2880 = (~w3987 & ~w17947) | (~w3987 & w12225) | (~w17947 & w12225);
assign w2881 = (~w3282 & w8986) | (~w3282 & w13222) | (w8986 & w13222);
assign w2882 = ~w7795 & ~w11308;
assign w2883 = a_51 & a_55;
assign w2884 = ~w3120 & ~w13121;
assign w2885 = a_7 & a_25;
assign w2886 = w15025 & ~w7834;
assign w2887 = ~w11336 & ~w1070;
assign w2888 = ~w1881 & ~w15272;
assign w2889 = w8302 & ~w6724;
assign w2890 = w13564 & ~w15213;
assign w2891 = (~w2100 & w12255) | (~w2100 & w10884) | (w12255 & w10884);
assign w2892 = w6462 & ~w8809;
assign w2893 = ~w16669 & ~w7417;
assign w2894 = ~w6249 & ~w16137;
assign w2895 = ~w9867 & ~w4407;
assign w2896 = ~w18747 & w12950;
assign w2897 = ~w15235 & ~w7767;
assign w2898 = ~w5956 & ~w11797;
assign w2899 = w7155 & w10662;
assign w2900 = ~w13303 & ~w17227;
assign w2901 = w5525 & w18891;
assign w2902 = ~w13082 & w1817;
assign w2903 = ~w14976 & w11733;
assign w2904 = ~w8201 & w1323;
assign w2905 = (~w11881 & ~w15823) | (~w11881 & w12605) | (~w15823 & w12605);
assign w2906 = ~w8358 & ~w8435;
assign w2907 = w16292 & w16434;
assign w2908 = ~w12824 & ~w780;
assign w2909 = ~w7856 & w12011;
assign w2910 = w14724 & w9555;
assign w2911 = ~w15343 & ~w6577;
assign w2912 = w5066 & w15494;
assign w2913 = ~w16135 & ~w4775;
assign w2914 = (~w13979 & w10840) | (~w13979 & w408) | (w10840 & w408);
assign w2915 = w11889 & ~w17848;
assign w2916 = ~w13263 & ~w10245;
assign w2917 = ~w10305 & ~w3956;
assign w2918 = ~w16703 & ~w18037;
assign w2919 = ~w667 & ~w3422;
assign w2920 = ~w4598 & w3350;
assign w2921 = a_22 & a_60;
assign w2922 = w17116 & ~w17023;
assign w2923 = ~w10111 & ~w8049;
assign w2924 = w2714 & ~w3354;
assign w2925 = ~w11649 & ~w4042;
assign w2926 = w17150 & w352;
assign w2927 = ~w18023 & ~w2314;
assign w2928 = ~w8685 & ~w15835;
assign w2929 = ~w2452 & ~w6983;
assign w2930 = (~w5115 & ~w17611) | (~w5115 & w15282) | (~w17611 & w15282);
assign w2931 = ~w18471 & ~w12903;
assign w2932 = ~w2189 & ~w18283;
assign w2933 = ~w1588 & ~w14571;
assign w2934 = w18959 & w17582;
assign w2935 = w8923 & w4525;
assign w2936 = w10873 & ~w9549;
assign w2937 = ~w424 & ~w16276;
assign w2938 = w4539 & ~w2523;
assign w2939 = ~w14165 & w1270;
assign w2940 = w5161 & w17541;
assign w2941 = w10852 & w1864;
assign w2942 = w1109 & w18305;
assign w2943 = w13281 & ~w2446;
assign w2944 = w3260 & w3297;
assign w2945 = ~w1138 & w14825;
assign w2946 = w1490 & w2457;
assign w2947 = w14533 & ~w1133;
assign w2948 = ~w16886 & ~w16140;
assign w2949 = ~w18707 & ~w13980;
assign w2950 = a_28 & w18620;
assign w2951 = a_32 & a_51;
assign w2952 = ~w5884 & ~w5320;
assign w2953 = ~w8885 & w16617;
assign w2954 = ~w9596 & ~w13119;
assign w2955 = ~w6200 & w6353;
assign w2956 = a_0 & a_27;
assign w2957 = ~w3606 & w4365;
assign w2958 = ~w4357 & w7038;
assign w2959 = w16189 & w828;
assign w2960 = ~w13569 & w17472;
assign w2961 = a_29 & a_35;
assign w2962 = ~w1441 & ~w11361;
assign w2963 = a_18 & a_27;
assign w2964 = ~w5074 & ~w17101;
assign w2965 = (~w1244 & ~w1788) | (~w1244 & w1590) | (~w1788 & w1590);
assign w2966 = a_12 & a_57;
assign w2967 = w1202 & ~w9091;
assign w2968 = a_14 & a_54;
assign w2969 = a_25 & a_30;
assign w2970 = ~w18155 & ~w17446;
assign w2971 = ~w15178 & ~w11525;
assign w2972 = (~w17433 & w5028) | (~w17433 & w9892) | (w5028 & w9892);
assign w2973 = ~w15584 & w14284;
assign w2974 = a_33 & a_55;
assign w2975 = ~w37 & ~w105;
assign w2976 = a_24 & a_39;
assign w2977 = ~w6101 & w11981;
assign w2978 = (~w6697 & ~w16669) | (~w6697 & w8383) | (~w16669 & w8383);
assign w2979 = ~w14011 & ~w13475;
assign w2980 = ~w3405 & w1611;
assign w2981 = w13078 & w16945;
assign w2982 = ~w10596 & ~w8385;
assign w2983 = w669 & ~w1017;
assign w2984 = ~w15941 & ~w10193;
assign w2985 = a_49 & a_51;
assign w2986 = ~w16662 & w4733;
assign w2987 = a_26 & a_44;
assign w2988 = a_36 & a_44;
assign w2989 = a_12 & a_55;
assign w2990 = ~w12779 & ~w2941;
assign w2991 = ~w5473 & ~w11783;
assign w2992 = w16918 & w6426;
assign w2993 = ~w733 & ~w3406;
assign w2994 = w9420 & w12243;
assign w2995 = w7177 & w19151;
assign w2996 = ~w11051 & ~w18923;
assign w2997 = ~w18627 & ~w9166;
assign w2998 = w1861 & ~w13687;
assign w2999 = w7565 & ~w9982;
assign w3000 = w621 & ~w17091;
assign w3001 = ~w8000 & ~w18306;
assign w3002 = w8426 & ~w14282;
assign w3003 = ~w9913 & w4730;
assign w3004 = w2817 & ~w15416;
assign w3005 = ~w16404 & w1496;
assign w3006 = ~w17812 & ~w11781;
assign w3007 = w18277 & ~w16928;
assign w3008 = ~w16177 & ~w5858;
assign w3009 = ~w1911 & ~w2822;
assign w3010 = ~w12481 & ~w4819;
assign w3011 = (~w3700 & w13082) | (~w3700 & w13575) | (w13082 & w13575);
assign w3012 = a_11 & a_59;
assign w3013 = a_2 & a_30;
assign w3014 = ~w1513 & ~w13645;
assign w3015 = ~w845 & ~w12655;
assign w3016 = ~w620 & ~w16066;
assign w3017 = ~w4908 & ~w18454;
assign w3018 = ~w17670 & ~w9334;
assign w3019 = w6853 & w3985;
assign w3020 = ~w16337 & ~w2159;
assign w3021 = (~w9987 & w5258) | (~w9987 & w4324) | (w5258 & w4324);
assign w3022 = ~w17842 & w14634;
assign w3023 = w16420 & w19111;
assign w3024 = ~w13600 & ~w8494;
assign w3025 = ~w4140 & ~w13720;
assign w3026 = ~w12037 & w4597;
assign w3027 = a_0 & a_32;
assign w3028 = ~w5046 & ~w18392;
assign w3029 = ~w10514 & ~w17624;
assign w3030 = a_23 & a_31;
assign w3031 = ~w18194 & ~w8698;
assign w3032 = ~w9502 & ~w13629;
assign w3033 = w461 & ~w13395;
assign w3034 = a_31 & a_43;
assign w3035 = ~w5365 & w7829;
assign w3036 = ~w14809 & ~w15606;
assign w3037 = ~w6964 & ~w16653;
assign w3038 = w11936 & w11487;
assign w3039 = w13294 & ~w17037;
assign w3040 = w6006 & w13815;
assign w3041 = w2975 & w1701;
assign w3042 = w5677 & w16421;
assign w3043 = ~w6501 & ~w4306;
assign w3044 = ~w8969 & ~w18565;
assign w3045 = (~w2396 & w15538) | (~w2396 & w18757) | (w15538 & w18757);
assign w3046 = ~w11561 & ~w12953;
assign w3047 = ~w4381 & ~w5606;
assign w3048 = ~w1587 & ~w4432;
assign w3049 = w4939 & w8657;
assign w3050 = w18147 & ~w1588;
assign w3051 = a_14 & a_47;
assign w3052 = w2723 & w784;
assign w3053 = ~w5765 & w11687;
assign w3054 = a_3 & a_51;
assign w3055 = w15335 & ~w11054;
assign w3056 = w15418 & ~w9528;
assign w3057 = ~w13311 & ~w786;
assign w3058 = w4502 & w12617;
assign w3059 = ~w14892 & ~w4709;
assign w3060 = ~w9813 & ~w10630;
assign w3061 = (w5464 & w17784) | (w5464 & w8336) | (w17784 & w8336);
assign w3062 = a_17 & a_32;
assign w3063 = w8083 & ~w14275;
assign w3064 = ~w17005 & ~w2346;
assign w3065 = w10697 & w17294;
assign w3066 = ~w9129 & w15351;
assign w3067 = ~w11079 & w13693;
assign w3068 = ~w3824 & ~w10798;
assign w3069 = w11106 & ~w7142;
assign w3070 = w2217 & ~w17521;
assign w3071 = (~w37 & ~w2975) | (~w37 & w9086) | (~w2975 & w9086);
assign w3072 = w2716 & w13626;
assign w3073 = w15734 & ~w16223;
assign w3074 = a_9 & a_25;
assign w3075 = ~w10097 & ~w4003;
assign w3076 = a_23 & a_25;
assign w3077 = a_44 & a_57;
assign w3078 = a_16 & a_49;
assign w3079 = ~w6124 & ~w2490;
assign w3080 = a_20 & a_35;
assign w3081 = a_8 & a_53;
assign w3082 = w10811 & w4209;
assign w3083 = ~w2035 & ~w1802;
assign w3084 = (~w10332 & ~w12656) | (~w10332 & w14626) | (~w12656 & w14626);
assign w3085 = (w14993 & ~w10099) | (w14993 & w4751) | (~w10099 & w4751);
assign w3086 = w10180 & ~w14093;
assign w3087 = ~w14757 & ~w18288;
assign w3088 = ~w13557 & ~w17305;
assign w3089 = a_20 & a_22;
assign w3090 = a_3 & a_34;
assign w3091 = ~w18089 & w3632;
assign w3092 = a_0 & a_59;
assign w3093 = w1652 & w16628;
assign w3094 = ~w17522 & ~w15615;
assign w3095 = w2502 & ~w11201;
assign w3096 = w3877 & ~w11913;
assign w3097 = w10861 & ~w13845;
assign w3098 = ~w14387 & ~w12054;
assign w3099 = a_6 & a_17;
assign w3100 = ~w19108 & ~w3900;
assign w3101 = ~w8546 & ~w14679;
assign w3102 = (~w17801 & ~w8392) | (~w17801 & w17871) | (~w8392 & w17871);
assign w3103 = (w2769 & w16759) | (w2769 & w18108) | (w16759 & w18108);
assign w3104 = ~w11004 & ~w1430;
assign w3105 = ~w17985 & w2363;
assign w3106 = ~w17733 & w15141;
assign w3107 = (w15988 & w16666) | (w15988 & w3760) | (w16666 & w3760);
assign w3108 = w15902 & w12236;
assign w3109 = ~w10827 & ~w15008;
assign w3110 = ~w4967 & w8783;
assign w3111 = w14608 & ~w11802;
assign w3112 = ~w318 & ~w3750;
assign w3113 = w17422 & ~w13483;
assign w3114 = (~w1962 & w486) | (~w1962 & w10622) | (w486 & w10622);
assign w3115 = a_36 & a_39;
assign w3116 = a_26 & a_57;
assign w3117 = ~w15980 & ~w8075;
assign w3118 = ~w18835 & ~w15658;
assign w3119 = a_18 & a_34;
assign w3120 = w6564 & ~w13360;
assign w3121 = a_5 & a_59;
assign w3122 = w16095 & ~w14916;
assign w3123 = ~w9105 & ~w436;
assign w3124 = w10261 & w3171;
assign w3125 = a_22 & a_59;
assign w3126 = w3378 & w10316;
assign w3127 = a_18 & a_25;
assign w3128 = ~w2540 & w10373;
assign w3129 = (~w5928 & ~w8017) | (~w5928 & w17839) | (~w8017 & w17839);
assign w3130 = a_17 & a_28;
assign w3131 = ~w17330 & ~w12475;
assign w3132 = ~w13608 & ~w4078;
assign w3133 = ~w8162 & ~w3110;
assign w3134 = ~w7089 & ~w6908;
assign w3135 = w7199 & ~w10547;
assign w3136 = w13005 & w4811;
assign w3137 = ~w11845 & ~w11308;
assign w3138 = ~w18049 & ~w7766;
assign w3139 = ~w18070 & ~w8768;
assign w3140 = w14333 & w5614;
assign w3141 = (~w1536 & ~w10475) | (~w1536 & w4191) | (~w10475 & w4191);
assign w3142 = ~w12134 & ~w8111;
assign w3143 = ~w10026 & ~w16336;
assign w3144 = ~w11537 & ~w3202;
assign w3145 = ~w4462 & ~w13427;
assign w3146 = ~w5890 & ~w18507;
assign w3147 = ~w14253 & w14347;
assign w3148 = ~w9088 & ~w18325;
assign w3149 = (~w2330 & w1540) | (~w2330 & w18128) | (w1540 & w18128);
assign w3150 = (~w12620 & ~w16882) | (~w12620 & w4707) | (~w16882 & w4707);
assign w3151 = w1857 & w7835;
assign w3152 = a_53 & a_57;
assign w3153 = ~w16327 & ~w610;
assign w3154 = ~w2772 & ~w3479;
assign w3155 = ~w16439 & w120;
assign w3156 = a_17 & a_21;
assign w3157 = w18422 & ~w1599;
assign w3158 = ~w17534 & w18281;
assign w3159 = ~w4268 & ~w14066;
assign w3160 = w3721 & w6842;
assign w3161 = ~w2455 & ~w13503;
assign w3162 = w2104 & ~w921;
assign w3163 = ~w8232 & ~w6909;
assign w3164 = w14001 & ~w14439;
assign w3165 = (w5673 & w2769) | (w5673 & w5826) | (w2769 & w5826);
assign w3166 = w14569 & ~w7276;
assign w3167 = ~w3246 & ~w11441;
assign w3168 = w1154 & ~w12384;
assign w3169 = ~w13049 & w13092;
assign w3170 = ~w2568 & ~w648;
assign w3171 = ~w4374 & ~w9101;
assign w3172 = a_3 & a_56;
assign w3173 = ~w14414 & w17974;
assign w3174 = ~w5670 & ~w764;
assign w3175 = (~w7102 & w14068) | (~w7102 & w6142) | (w14068 & w6142);
assign w3176 = ~w2078 & ~w18416;
assign w3177 = w10842 & ~w12526;
assign w3178 = w1434 & w17904;
assign w3179 = (~w18980 & w13945) | (~w18980 & w6791) | (w13945 & w6791);
assign w3180 = ~w18229 & ~w10906;
assign w3181 = ~w14624 & ~w16568;
assign w3182 = (w17620 & w12095) | (w17620 & w3600) | (w12095 & w3600);
assign w3183 = a_16 & a_29;
assign w3184 = ~w13940 & w10833;
assign w3185 = ~w8447 & ~w6213;
assign w3186 = ~w3188 & ~w12117;
assign w3187 = a_47 & a_56;
assign w3188 = a_0 & a_18;
assign w3189 = ~w1233 & ~w891;
assign w3190 = ~w1499 & ~w4754;
assign w3191 = ~w15810 & ~w1841;
assign w3192 = ~w10117 & ~w17085;
assign w3193 = w5123 & ~w4380;
assign w3194 = a_54 & a_63;
assign w3195 = a_12 & a_24;
assign w3196 = ~w17536 & ~w8546;
assign w3197 = w10029 & ~w17744;
assign w3198 = w6733 & w7386;
assign w3199 = w12501 & w12376;
assign w3200 = ~w9630 & ~w18739;
assign w3201 = ~w6858 & ~w2335;
assign w3202 = ~w17100 & ~w17086;
assign w3203 = w8943 & ~w5068;
assign w3204 = ~w4461 & ~w17019;
assign w3205 = w12324 & w15121;
assign w3206 = ~w15976 & w9451;
assign w3207 = w2185 & w12650;
assign w3208 = (~w16652 & ~w11683) | (~w16652 & w17439) | (~w11683 & w17439);
assign w3209 = ~w14765 & ~w8425;
assign w3210 = w10909 & ~w3138;
assign w3211 = ~w16595 & w2466;
assign w3212 = ~w14418 & w7913;
assign w3213 = ~w14930 & w6321;
assign w3214 = w6531 & w18889;
assign w3215 = ~w16778 & ~w7633;
assign w3216 = w9390 & ~w6317;
assign w3217 = w5523 & ~w2549;
assign w3218 = w10889 & ~w14809;
assign w3219 = ~w10198 & w9143;
assign w3220 = w10879 & ~w3355;
assign w3221 = a_14 & a_55;
assign w3222 = ~w1727 & ~w18935;
assign w3223 = w18116 & w17286;
assign w3224 = ~w4813 & ~w1470;
assign w3225 = a_10 & a_46;
assign w3226 = w19004 & ~w4364;
assign w3227 = a_43 & a_62;
assign w3228 = w11551 & ~w5594;
assign w3229 = ~w5255 & ~w9832;
assign w3230 = ~w3426 & ~w14350;
assign w3231 = ~w7032 & ~w5873;
assign w3232 = ~w12595 & ~w17581;
assign w3233 = ~w1829 & ~w401;
assign w3234 = ~w10580 & w11380;
assign w3235 = (w15380 & w8780) | (w15380 & w12205) | (w8780 & w12205);
assign w3236 = a_16 & a_61;
assign w3237 = ~w11578 & ~w10365;
assign w3238 = ~w9337 & w17049;
assign w3239 = a_5 & a_52;
assign w3240 = w8507 & ~w4949;
assign w3241 = w6476 & w2281;
assign w3242 = w17284 & w10356;
assign w3243 = w17588 & w509;
assign w3244 = w11040 & ~w12125;
assign w3245 = ~w3463 & ~w1697;
assign w3246 = w16498 & ~w13299;
assign w3247 = ~w7409 & w18490;
assign w3248 = ~w156 & ~w18204;
assign w3249 = w5323 & ~w6542;
assign w3250 = a_47 & a_57;
assign w3251 = w4968 & w15354;
assign w3252 = ~w1758 & ~w4449;
assign w3253 = ~w12852 & ~w13179;
assign w3254 = ~w1824 & ~w6195;
assign w3255 = (w2526 & w2769) | (w2526 & w15720) | (w2769 & w15720);
assign w3256 = w8687 & w11241;
assign w3257 = ~w14121 & w16994;
assign w3258 = w4603 & w328;
assign w3259 = ~w7714 & ~w8209;
assign w3260 = ~w10941 & ~w12355;
assign w3261 = ~w2864 & w16270;
assign w3262 = ~w10676 & ~w12144;
assign w3263 = a_57 & a_59;
assign w3264 = ~w14881 & ~w981;
assign w3265 = ~w9708 & ~w14949;
assign w3266 = w2042 & ~w4623;
assign w3267 = ~w6297 & ~w18824;
assign w3268 = ~w8408 & ~w1528;
assign w3269 = ~w9351 & ~w7157;
assign w3270 = ~w3444 & ~w14081;
assign w3271 = ~w15632 & ~w939;
assign w3272 = w3533 & ~w13974;
assign w3273 = ~w14994 & ~w18665;
assign w3274 = (w16842 & w10330) | (w16842 & w8273) | (w10330 & w8273);
assign w3275 = ~w3260 & ~w3297;
assign w3276 = a_40 & a_50;
assign w3277 = (~w5778 & ~w1574) | (~w5778 & w11427) | (~w1574 & w11427);
assign w3278 = ~w799 & ~w14672;
assign w3279 = w139 & w19152;
assign w3280 = w8352 & w15414;
assign w3281 = (w16174 & w4170) | (w16174 & w8981) | (w4170 & w8981);
assign w3282 = ~w1865 & w9223;
assign w3283 = w5475 & w18470;
assign w3284 = (~w998 & ~w17454) | (~w998 & w390) | (~w17454 & w390);
assign w3285 = a_41 & a_46;
assign w3286 = ~w1035 & ~w17172;
assign w3287 = ~a_41 & a_42;
assign w3288 = w3616 & w18424;
assign w3289 = a_4 & a_49;
assign w3290 = ~w2478 & ~w7432;
assign w3291 = ~w2655 & ~w17012;
assign w3292 = w11701 & w2021;
assign w3293 = ~w18383 & w2541;
assign w3294 = ~w14302 & w6675;
assign w3295 = w11189 & ~w17969;
assign w3296 = ~w14805 & ~w4745;
assign w3297 = ~w9797 & ~w10605;
assign w3298 = w5434 & w8649;
assign w3299 = a_1 & a_25;
assign w3300 = ~w6275 & ~w153;
assign w3301 = w12048 & ~w475;
assign w3302 = ~w16599 & ~w17215;
assign w3303 = (~w4586 & ~w13666) | (~w4586 & w15164) | (~w13666 & w15164);
assign w3304 = ~w15126 & ~w14859;
assign w3305 = w4299 & w14878;
assign w3306 = a_27 & a_57;
assign w3307 = w9807 & ~w14449;
assign w3308 = ~w8738 & ~w5094;
assign w3309 = ~w16753 & ~w17525;
assign w3310 = a_43 & a_53;
assign w3311 = w3770 & ~w1570;
assign w3312 = w11455 & ~w16929;
assign w3313 = ~w5262 & ~w13053;
assign w3314 = a_2 & a_58;
assign w3315 = w6304 & w2228;
assign w3316 = a_23 & a_33;
assign w3317 = ~w19076 & ~w900;
assign w3318 = ~w6538 & ~w3923;
assign w3319 = ~w256 & ~w10211;
assign w3320 = w12812 & w16213;
assign w3321 = w12331 & ~w8004;
assign w3322 = ~w17772 & ~w2338;
assign w3323 = ~w2724 & ~w14946;
assign w3324 = w18175 & ~w10504;
assign w3325 = ~w8016 & ~w10530;
assign w3326 = ~w5311 & ~w13982;
assign w3327 = ~w11547 & w11075;
assign w3328 = ~w1390 & ~w12767;
assign w3329 = ~w4449 & ~w17596;
assign w3330 = ~w16833 & ~w12783;
assign w3331 = ~a_24 & ~w17912;
assign w3332 = a_10 & a_23;
assign w3333 = ~w7711 & w13997;
assign w3334 = ~w18604 & ~w3869;
assign w3335 = ~w14615 & w1140;
assign w3336 = ~w12812 & ~w16213;
assign w3337 = ~w10484 & ~w14373;
assign w3338 = (~w6834 & w6291) | (~w6834 & w1596) | (w6291 & w1596);
assign w3339 = ~w5793 & ~w17566;
assign w3340 = w1366 & w16184;
assign w3341 = a_23 & a_41;
assign w3342 = ~w7567 & ~w3049;
assign w3343 = ~w9597 & w14769;
assign w3344 = ~w3765 & ~w9894;
assign w3345 = (w2615 & w2361) | (w2615 & w10231) | (w2361 & w10231);
assign w3346 = ~w5213 & w18960;
assign w3347 = ~w9134 & w13110;
assign w3348 = ~w3937 & ~w16056;
assign w3349 = ~w15823 & ~w7139;
assign w3350 = ~w848 & ~w1043;
assign w3351 = ~w12939 & ~w2851;
assign w3352 = w7090 & ~w14915;
assign w3353 = ~w1304 & ~w752;
assign w3354 = ~w1360 & ~w9659;
assign w3355 = ~w2339 & ~w3733;
assign w3356 = ~w13304 & ~w8095;
assign w3357 = (w4559 & w3232) | (w4559 & w9730) | (w3232 & w9730);
assign w3358 = ~w9870 & ~w14997;
assign w3359 = w17258 & w3068;
assign w3360 = ~w16103 & ~w2191;
assign w3361 = (w9893 & w2769) | (w9893 & w12329) | (w2769 & w12329);
assign w3362 = ~w3223 & ~w8110;
assign w3363 = ~w1300 & ~w18071;
assign w3364 = w10733 & ~w4824;
assign w3365 = ~w2588 & ~w12115;
assign w3366 = ~w2901 & ~w6561;
assign w3367 = w12789 & ~w14906;
assign w3368 = ~w13105 & ~w8850;
assign w3369 = w5695 & ~w16764;
assign w3370 = w9096 & w15733;
assign w3371 = w2142 & ~w17874;
assign w3372 = a_40 & a_45;
assign w3373 = a_2 & a_23;
assign w3374 = w9060 & ~w3437;
assign w3375 = ~w12572 & ~w11032;
assign w3376 = (w11176 & w2235) | (w11176 & w8420) | (w2235 & w8420);
assign w3377 = a_22 & a_46;
assign w3378 = a_21 & a_32;
assign w3379 = ~w1674 & ~w16258;
assign w3380 = ~w8034 & ~w6847;
assign w3381 = ~w18341 & ~w1965;
assign w3382 = w16135 & w4775;
assign w3383 = w2035 & w1802;
assign w3384 = w9612 & w8745;
assign w3385 = ~w14327 & ~w3484;
assign w3386 = ~w17471 & w4292;
assign w3387 = ~w7349 & ~w5467;
assign w3388 = (~w4541 & w1648) | (~w4541 & w1933) | (w1648 & w1933);
assign w3389 = w4048 & ~w11740;
assign w3390 = ~w7984 & ~w9205;
assign w3391 = a_1 & a_48;
assign w3392 = ~w16446 & ~w2070;
assign w3393 = ~w12137 & w5821;
assign w3394 = ~w3445 & ~w11763;
assign w3395 = ~w2861 & ~w9510;
assign w3396 = ~w12784 & ~w1292;
assign w3397 = w10228 & ~w16977;
assign w3398 = a_27 & a_38;
assign w3399 = ~w7465 & w15865;
assign w3400 = ~w12922 & ~w14703;
assign w3401 = ~w7911 & w1500;
assign w3402 = ~w8736 & w6471;
assign w3403 = a_41 & a_42;
assign w3404 = ~w18882 & ~w5160;
assign w3405 = (~w741 & ~w3777) | (~w741 & w6822) | (~w3777 & w6822);
assign w3406 = ~w8360 & w1429;
assign w3407 = ~w17872 & ~w1458;
assign w3408 = w13998 & w1534;
assign w3409 = w15004 & w17106;
assign w3410 = w17515 & w45;
assign w3411 = ~w13187 & ~w17263;
assign w3412 = w776 & w2387;
assign w3413 = ~w17549 & ~w4152;
assign w3414 = ~w13186 & w6834;
assign w3415 = ~w13282 & ~w6539;
assign w3416 = w15918 & ~w17169;
assign w3417 = ~w4420 & w10231;
assign w3418 = a_27 & a_44;
assign w3419 = (w2769 & w13007) | (w2769 & w13554) | (w13007 & w13554);
assign w3420 = ~w10955 & ~w6394;
assign w3421 = w7004 & ~w7736;
assign w3422 = ~w15901 & ~w17393;
assign w3423 = w18828 & ~w5342;
assign w3424 = ~w7754 & w5578;
assign w3425 = ~w5059 & ~w7287;
assign w3426 = ~w4998 & w1999;
assign w3427 = ~w6304 & ~w17;
assign w3428 = ~w5270 & w18929;
assign w3429 = w8904 & ~w3689;
assign w3430 = ~w21 & ~w16624;
assign w3431 = a_49 & a_52;
assign w3432 = ~w5438 & w1923;
assign w3433 = ~w6888 & ~w7239;
assign w3434 = ~w6595 & ~w11042;
assign w3435 = ~w468 & ~w13341;
assign w3436 = w15126 & w19026;
assign w3437 = ~w9125 & ~w2718;
assign w3438 = w13036 & ~w2210;
assign w3439 = w12477 & ~w10517;
assign w3440 = w11332 & w15601;
assign w3441 = w15858 & ~w8537;
assign w3442 = ~w5852 & ~w2052;
assign w3443 = (~w6547 & w10937) | (~w6547 & w17289) | (w10937 & w17289);
assign w3444 = w2313 & w6030;
assign w3445 = w734 & ~w915;
assign w3446 = ~w7129 & w12218;
assign w3447 = w17600 & ~w6935;
assign w3448 = w5194 & w13083;
assign w3449 = w5482 & w14935;
assign w3450 = ~w851 & ~w14178;
assign w3451 = w10010 & ~w15978;
assign w3452 = ~w8344 & ~w1825;
assign w3453 = w18838 & ~w5134;
assign w3454 = (~w14747 & ~w13135) | (~w14747 & w8483) | (~w13135 & w8483);
assign w3455 = ~w5480 & ~w1558;
assign w3456 = ~w12701 & ~w15197;
assign w3457 = ~w882 & ~w11646;
assign w3458 = w10679 & w5752;
assign w3459 = ~w8568 & ~w9715;
assign w3460 = w6829 & ~w6734;
assign w3461 = w4257 & ~w17837;
assign w3462 = w5506 & ~w17197;
assign w3463 = a_10 & a_19;
assign w3464 = ~w8806 & w14059;
assign w3465 = w2844 & w19153;
assign w3466 = a_37 & a_55;
assign w3467 = ~w16890 & ~w18804;
assign w3468 = a_12 & a_25;
assign w3469 = ~w6551 & ~w11666;
assign w3470 = ~w6649 & ~w12577;
assign w3471 = ~w11644 & w13923;
assign w3472 = w1191 & ~w16838;
assign w3473 = w3176 & w17009;
assign w3474 = ~w7786 & w6358;
assign w3475 = w17526 & w3385;
assign w3476 = w14361 & ~w6699;
assign w3477 = (~w18844 & ~w1601) | (~w18844 & w3940) | (~w1601 & w3940);
assign w3478 = w13306 & ~w13670;
assign w3479 = ~w7131 & ~w14638;
assign w3480 = ~w18591 & ~w7141;
assign w3481 = w17471 & ~w4292;
assign w3482 = ~w8508 & ~w15502;
assign w3483 = w6274 & ~w564;
assign w3484 = w15726 & ~w17156;
assign w3485 = w3549 & w5256;
assign w3486 = ~w6163 & w10917;
assign w3487 = a_0 & a_61;
assign w3488 = w9079 & ~w10061;
assign w3489 = a_29 & a_38;
assign w3490 = w13820 & w5790;
assign w3491 = a_40 & a_47;
assign w3492 = (~w3088 & ~w17497) | (~w3088 & w10101) | (~w17497 & w10101);
assign w3493 = ~w6349 & w5001;
assign w3494 = ~a_33 & ~w1913;
assign w3495 = w3591 & ~w15093;
assign w3496 = w2590 & w8249;
assign w3497 = w7293 & w11033;
assign w3498 = ~w5340 & ~w14563;
assign w3499 = ~w6443 & ~w18749;
assign w3500 = ~w5541 & w9922;
assign w3501 = ~w10261 & ~w3171;
assign w3502 = a_15 & a_43;
assign w3503 = w3602 & ~w12798;
assign w3504 = a_6 & a_46;
assign w3505 = w12703 & w10336;
assign w3506 = a_20 & a_27;
assign w3507 = ~w8234 & ~w620;
assign w3508 = ~w18672 & w18954;
assign w3509 = w4976 & w7216;
assign w3510 = ~w4984 & ~w10949;
assign w3511 = w14759 & ~w2559;
assign w3512 = ~w2079 & w12126;
assign w3513 = w3952 & ~w112;
assign w3514 = a_7 & a_44;
assign w3515 = ~w15367 & ~w9826;
assign w3516 = w18432 & w3231;
assign w3517 = ~w14204 & w3675;
assign w3518 = w8782 & w4585;
assign w3519 = (w9337 & w12353) | (w9337 & w17165) | (w12353 & w17165);
assign w3520 = ~w929 & w8309;
assign w3521 = ~w6326 & ~w17212;
assign w3522 = ~w9301 & ~w3126;
assign w3523 = w5465 & ~w2624;
assign w3524 = w13210 & ~w13992;
assign w3525 = ~w17199 & ~w18526;
assign w3526 = ~w7418 & ~w18154;
assign w3527 = w9741 & w2790;
assign w3528 = ~w8909 & w5644;
assign w3529 = ~w7076 & ~w5800;
assign w3530 = ~w17571 & ~w12852;
assign w3531 = (w16892 & w18980) | (w16892 & w12366) | (w18980 & w12366);
assign w3532 = ~w4435 & ~w2816;
assign w3533 = ~w18227 & ~w736;
assign w3534 = a_6 & a_52;
assign w3535 = w12971 & ~w13237;
assign w3536 = ~w3089 & ~w8589;
assign w3537 = ~w14909 & ~w12445;
assign w3538 = ~w11273 & w8594;
assign w3539 = ~w13922 & ~w4720;
assign w3540 = ~w2682 & ~w3780;
assign w3541 = ~w5108 & w16437;
assign w3542 = a_11 & a_63;
assign w3543 = ~w6860 & ~w15021;
assign w3544 = w14183 & w2010;
assign w3545 = ~w14167 & w16729;
assign w3546 = w12761 & w385;
assign w3547 = a_20 & a_63;
assign w3548 = ~w11551 & ~w1398;
assign w3549 = a_7 & a_15;
assign w3550 = ~w8791 & ~w1015;
assign w3551 = w11136 & ~w1625;
assign w3552 = ~w7408 & ~w2556;
assign w3553 = w1267 & w3302;
assign w3554 = ~w9586 & w8865;
assign w3555 = ~w18551 & ~w12370;
assign w3556 = ~w18937 & ~w2436;
assign w3557 = w5397 & ~w18126;
assign w3558 = ~w16382 & ~w18377;
assign w3559 = w4872 & ~w14422;
assign w3560 = ~w8830 & ~w10673;
assign w3561 = ~w18753 & w2109;
assign w3562 = a_51 & a_53;
assign w3563 = w5019 & ~w485;
assign w3564 = ~w1995 & w16692;
assign w3565 = ~w7242 & w8416;
assign w3566 = w17680 & w3284;
assign w3567 = ~w1149 & ~w8980;
assign w3568 = w3337 & w1807;
assign w3569 = ~w1845 & ~w9543;
assign w3570 = (~w12344 & ~w6278) | (~w12344 & w1813) | (~w6278 & w1813);
assign w3571 = ~w19070 & ~w2895;
assign w3572 = (w1920 & ~w6575) | (w1920 & w4417) | (~w6575 & w4417);
assign w3573 = a_1 & a_29;
assign w3574 = a_0 & a_6;
assign w3575 = ~w4611 & w4166;
assign w3576 = ~w5360 & w11651;
assign w3577 = ~w17821 & w637;
assign w3578 = ~a_21 & ~w4744;
assign w3579 = ~w7454 & ~w3977;
assign w3580 = ~w625 & ~w8140;
assign w3581 = w17123 & w8962;
assign w3582 = a_15 & a_16;
assign w3583 = a_7 & a_17;
assign w3584 = w16532 & w2232;
assign w3585 = ~w834 & ~w14794;
assign w3586 = ~w11320 & ~w10805;
assign w3587 = ~w8197 & ~w2552;
assign w3588 = w13522 & ~w5315;
assign w3589 = ~w11357 & w15241;
assign w3590 = w7751 & w12078;
assign w3591 = a_47 & a_59;
assign w3592 = ~w1125 & ~w6609;
assign w3593 = w8637 & ~w2875;
assign w3594 = ~w6673 & ~w4136;
assign w3595 = ~w4266 & ~w2256;
assign w3596 = w5453 & w12319;
assign w3597 = ~w621 & w17091;
assign w3598 = w11350 & ~w16417;
assign w3599 = w10455 & w14896;
assign w3600 = ~w7360 & w17620;
assign w3601 = (w63 & w5389) | (w63 & w8472) | (w5389 & w8472);
assign w3602 = (~w6944 & ~w5090) | (~w6944 & w13314) | (~w5090 & w13314);
assign w3603 = ~w9711 & ~w4504;
assign w3604 = ~w2133 & w781;
assign w3605 = ~w14990 & ~w7041;
assign w3606 = a_3 & a_21;
assign w3607 = a_20 & a_41;
assign w3608 = w18017 & w14161;
assign w3609 = ~w2140 & w10068;
assign w3610 = ~w1298 & ~w1989;
assign w3611 = ~w1730 & w6542;
assign w3612 = w91 & ~w18727;
assign w3613 = w17466 & ~w12597;
assign w3614 = a_10 & a_28;
assign w3615 = a_24 & a_28;
assign w3616 = ~w18914 & ~w8688;
assign w3617 = ~w11570 & w11364;
assign w3618 = w15025 & w11395;
assign w3619 = ~w12690 & ~w214;
assign w3620 = ~w9766 & ~w2124;
assign w3621 = (~w2541 & w7610) | (~w2541 & w12198) | (w7610 & w12198);
assign w3622 = ~w4557 & w14929;
assign w3623 = ~w15271 & ~w14600;
assign w3624 = ~w1146 & ~w2086;
assign w3625 = ~w1564 & ~w3941;
assign w3626 = ~w10621 & ~w9507;
assign w3627 = w1576 & w1320;
assign w3628 = ~w440 & ~w6634;
assign w3629 = a_21 & a_22;
assign w3630 = w86 & ~w18078;
assign w3631 = w5904 & w17701;
assign w3632 = ~w1978 & ~w17397;
assign w3633 = a_24 & a_58;
assign w3634 = w9586 & ~w8865;
assign w3635 = w10109 & w2863;
assign w3636 = ~w10456 & ~w5450;
assign w3637 = ~w4419 & ~w10247;
assign w3638 = ~w7756 & w2700;
assign w3639 = ~w1109 & ~w18305;
assign w3640 = ~w8001 & ~w1606;
assign w3641 = w678 & w11340;
assign w3642 = ~w4770 & ~w2120;
assign w3643 = ~w209 & ~w8888;
assign w3644 = w17272 & ~w833;
assign w3645 = ~w11390 & w12734;
assign w3646 = ~w2592 & ~w9271;
assign w3647 = ~w15873 & ~w6778;
assign w3648 = ~w13359 & ~w9602;
assign w3649 = a_58 & a_63;
assign w3650 = ~w17070 & ~w5487;
assign w3651 = ~w15822 & ~w4926;
assign w3652 = a_55 & a_63;
assign w3653 = ~w24 & ~w13543;
assign w3654 = ~w11551 & w5594;
assign w3655 = ~w5204 & ~w9428;
assign w3656 = w10419 & ~w4021;
assign w3657 = w8334 & ~w11318;
assign w3658 = a_29 & a_43;
assign w3659 = ~w18432 & ~w3231;
assign w3660 = w18690 & w16760;
assign w3661 = ~w9825 & w2783;
assign w3662 = ~w6984 & ~w1842;
assign w3663 = ~w13312 & w13134;
assign w3664 = ~w17580 & w8072;
assign w3665 = w9172 & ~w2363;
assign w3666 = a_18 & a_30;
assign w3667 = ~w9959 & ~w18982;
assign w3668 = ~w14581 & ~w8712;
assign w3669 = ~w17768 & ~w2741;
assign w3670 = ~w4108 & ~w10084;
assign w3671 = w18942 & ~w2678;
assign w3672 = (~w10066 & ~w12296) | (~w10066 & w10994) | (~w12296 & w10994);
assign w3673 = w5604 & w14094;
assign w3674 = w10495 & ~w14342;
assign w3675 = ~w15053 & ~w10281;
assign w3676 = w7754 & ~w5578;
assign w3677 = ~w14771 & ~w9652;
assign w3678 = ~w19115 & ~w17012;
assign w3679 = w8012 & ~w4415;
assign w3680 = ~w2176 & w5756;
assign w3681 = ~w18236 & ~w6792;
assign w3682 = ~w4880 & w655;
assign w3683 = a_33 & a_45;
assign w3684 = ~w5401 & ~w9557;
assign w3685 = ~w11399 & ~w17187;
assign w3686 = w8469 & ~w8560;
assign w3687 = ~w9650 & ~w14128;
assign w3688 = ~w15713 & ~w18161;
assign w3689 = ~w15587 & ~w14490;
assign w3690 = (w19005 & w2069) | (w19005 & w12708) | (w2069 & w12708);
assign w3691 = w13884 & w12820;
assign w3692 = ~w16513 & w1959;
assign w3693 = w11079 & ~w13693;
assign w3694 = ~w10631 & ~w222;
assign w3695 = ~w9778 & ~w994;
assign w3696 = w1839 & ~w15884;
assign w3697 = ~w2978 & ~w10964;
assign w3698 = w7564 & ~w5938;
assign w3699 = a_25 & a_45;
assign w3700 = ~w9668 & ~w10603;
assign w3701 = ~w5019 & w15172;
assign w3702 = ~w1629 & ~w14481;
assign w3703 = ~w12274 & ~w11461;
assign w3704 = w6855 & ~w13456;
assign w3705 = ~w18942 & w2678;
assign w3706 = ~w691 & w15106;
assign w3707 = w1673 & ~w6977;
assign w3708 = w8950 & ~w11771;
assign w3709 = ~w7701 & w7441;
assign w3710 = (w17890 & w729) | (w17890 & w9935) | (w729 & w9935);
assign w3711 = ~w17794 & ~w1676;
assign w3712 = w15833 & ~w18967;
assign w3713 = a_20 & a_62;
assign w3714 = ~w9817 & ~w11632;
assign w3715 = ~w4481 & w5871;
assign w3716 = ~w19087 & ~w5999;
assign w3717 = ~w7856 & ~w6263;
assign w3718 = ~w14548 & ~w11046;
assign w3719 = ~w4346 & w16358;
assign w3720 = w12781 & ~w18253;
assign w3721 = (~w2432 & ~w13818) | (~w2432 & w6219) | (~w13818 & w6219);
assign w3722 = ~w5602 & w11887;
assign w3723 = w10469 & w5810;
assign w3724 = ~w14904 & w14267;
assign w3725 = ~w5829 & ~w4601;
assign w3726 = ~w11440 & w12934;
assign w3727 = w15234 & w14095;
assign w3728 = ~w10449 & w18219;
assign w3729 = ~w18723 & ~w1105;
assign w3730 = ~w4009 & ~w19076;
assign w3731 = ~w13017 & ~w2072;
assign w3732 = ~w13238 & ~w3399;
assign w3733 = w13827 & w2163;
assign w3734 = a_43 & a_47;
assign w3735 = w13486 & w2860;
assign w3736 = ~w16382 & ~w9240;
assign w3737 = a_3 & a_5;
assign w3738 = (w961 & w4889) | (w961 & ~w5108) | (w4889 & ~w5108);
assign w3739 = ~w963 & w16863;
assign w3740 = w7086 & w17139;
assign w3741 = w1671 & ~w13389;
assign w3742 = w4138 & ~w5041;
assign w3743 = w11786 & w18661;
assign w3744 = a_0 & a_15;
assign w3745 = ~w6109 & ~w14176;
assign w3746 = ~w13158 & w10854;
assign w3747 = w16830 & ~w14260;
assign w3748 = ~w12839 & ~w14780;
assign w3749 = ~w2336 & ~w7056;
assign w3750 = ~w7092 & ~w8395;
assign w3751 = ~w5927 & ~w11185;
assign w3752 = ~w3104 & ~w194;
assign w3753 = ~w17374 & ~w15479;
assign w3754 = ~w15519 & w2477;
assign w3755 = ~w9627 & ~w13239;
assign w3756 = a_2 & a_35;
assign w3757 = a_16 & a_56;
assign w3758 = a_4 & a_52;
assign w3759 = ~w18157 & ~w6147;
assign w3760 = w8974 & w16661;
assign w3761 = ~w10509 & ~w3581;
assign w3762 = w10495 & w8574;
assign w3763 = (~w559 & ~w14486) | (~w559 & w810) | (~w14486 & w810);
assign w3764 = w16494 & w9299;
assign w3765 = ~w18259 & ~w7370;
assign w3766 = ~w18017 & w11852;
assign w3767 = w3668 & ~w9193;
assign w3768 = ~w10404 & ~w10883;
assign w3769 = ~w7059 & ~w6629;
assign w3770 = a_11 & a_28;
assign w3771 = w9914 & ~w13920;
assign w3772 = w17829 & w12114;
assign w3773 = a_16 & a_43;
assign w3774 = ~w11146 & w4960;
assign w3775 = ~w10171 & ~w7687;
assign w3776 = w208 & w7110;
assign w3777 = ~w6556 & ~w741;
assign w3778 = ~w4206 & ~w10953;
assign w3779 = ~w5438 & w12449;
assign w3780 = w3574 & w6534;
assign w3781 = w7390 & w15425;
assign w3782 = ~w4996 & w17309;
assign w3783 = ~w14926 & ~w7742;
assign w3784 = ~w16321 & ~w15924;
assign w3785 = w10393 & w5182;
assign w3786 = w12919 & ~w5712;
assign w3787 = ~w6920 & ~w15908;
assign w3788 = ~w3309 & w9666;
assign w3789 = a_46 & a_57;
assign w3790 = ~w6313 & ~w16685;
assign w3791 = ~w4405 & w1531;
assign w3792 = w10616 & ~w9933;
assign w3793 = w13466 & ~w1924;
assign w3794 = w6372 & ~w10218;
assign w3795 = a_3 & a_54;
assign w3796 = ~w8203 & ~w14861;
assign w3797 = ~w5643 & ~w281;
assign w3798 = w8939 & ~w9195;
assign w3799 = ~w14110 & ~w17944;
assign w3800 = a_32 & a_46;
assign w3801 = w9476 & w6097;
assign w3802 = ~w12123 & ~w8815;
assign w3803 = w98 & w4978;
assign w3804 = ~w5896 & ~w3416;
assign w3805 = ~w18545 & ~w16616;
assign w3806 = w14980 & w19154;
assign w3807 = (w6567 & ~w12288) | (w6567 & ~w999) | (~w12288 & ~w999);
assign w3808 = w511 & ~w12533;
assign w3809 = ~w1448 & w10468;
assign w3810 = (~w11436 & ~w16761) | (~w11436 & w8102) | (~w16761 & w8102);
assign w3811 = ~w18916 & ~w8057;
assign w3812 = ~w16536 & ~w11326;
assign w3813 = w1575 & ~w10634;
assign w3814 = w13054 & ~w14466;
assign w3815 = w3542 & ~w10324;
assign w3816 = ~w17034 & w7196;
assign w3817 = ~w10617 & ~w6449;
assign w3818 = a_22 & a_39;
assign w3819 = ~w15128 & w10808;
assign w3820 = ~w6578 & ~w5830;
assign w3821 = w7099 & ~w6309;
assign w3822 = ~w10381 & ~w11937;
assign w3823 = w2563 & ~w14328;
assign w3824 = w4946 & w7919;
assign w3825 = ~a_58 & a_59;
assign w3826 = ~w15170 & ~w18861;
assign w3827 = ~w7034 & w8740;
assign w3828 = ~w6660 & w6359;
assign w3829 = ~w4856 & ~w10229;
assign w3830 = ~w18595 & ~w15518;
assign w3831 = ~w3111 & ~w17042;
assign w3832 = a_14 & a_19;
assign w3833 = a_21 & a_38;
assign w3834 = w3194 & ~w7699;
assign w3835 = ~w2401 & ~w1157;
assign w3836 = ~w5961 & ~w8921;
assign w3837 = ~w17553 & ~w7220;
assign w3838 = w3277 & ~w7796;
assign w3839 = a_32 & a_43;
assign w3840 = ~w9512 & w5376;
assign w3841 = ~w14112 & ~w17486;
assign w3842 = w9896 & ~w13473;
assign w3843 = ~w7280 & ~w7400;
assign w3844 = ~w7430 & w4580;
assign w3845 = w15763 & ~w4979;
assign w3846 = a_51 & a_54;
assign w3847 = w10647 & ~w17279;
assign w3848 = ~w7407 & w18659;
assign w3849 = w17585 & ~w4748;
assign w3850 = ~w14379 & ~w9769;
assign w3851 = w8574 & ~w5291;
assign w3852 = ~w763 & ~w18825;
assign w3853 = (w14650 & w5142) | (w14650 & ~w11689) | (w5142 & ~w11689);
assign w3854 = w14598 & w4338;
assign w3855 = ~w18648 & w3271;
assign w3856 = ~w11538 & ~w632;
assign w3857 = ~w12492 & w10862;
assign w3858 = ~w13457 & w14990;
assign w3859 = ~w17274 & ~w15340;
assign w3860 = w8525 & w12666;
assign w3861 = ~w6528 & ~w3432;
assign w3862 = (~w13076 & ~w13294) | (~w13076 & w12709) | (~w13294 & w12709);
assign w3863 = ~w12226 & ~w9218;
assign w3864 = ~w16448 & ~w13806;
assign w3865 = ~w3605 & ~w1648;
assign w3866 = ~w4831 & ~w9160;
assign w3867 = a_38 & a_55;
assign w3868 = ~w1223 & ~w11028;
assign w3869 = w6996 & w3434;
assign w3870 = ~w10447 & ~w2143;
assign w3871 = w2010 & w10302;
assign w3872 = w11118 & ~w13270;
assign w3873 = w17374 & w15479;
assign w3874 = a_5 & a_37;
assign w3875 = w6098 & ~w4931;
assign w3876 = (~w5400 & ~w15252) | (~w5400 & w12607) | (~w15252 & w12607);
assign w3877 = ~w18324 & ~w10062;
assign w3878 = ~w15353 & ~w9217;
assign w3879 = ~w609 & ~w13198;
assign w3880 = ~w14357 & ~w17213;
assign w3881 = ~w13425 & ~w4614;
assign w3882 = ~w18943 & w17462;
assign w3883 = a_22 & a_61;
assign w3884 = ~w13806 & ~w2317;
assign w3885 = ~w13286 & ~w12942;
assign w3886 = w18598 & ~w12292;
assign w3887 = ~w17634 & ~w10404;
assign w3888 = a_25 & a_44;
assign w3889 = w15937 & ~w9280;
assign w3890 = w4158 & ~w18545;
assign w3891 = ~w865 & ~w13056;
assign w3892 = w4268 & w14066;
assign w3893 = ~w16189 & ~w828;
assign w3894 = w914 & ~w10292;
assign w3895 = w18025 & ~w3918;
assign w3896 = ~w18765 & w13517;
assign w3897 = ~w16591 & ~w14686;
assign w3898 = ~w16364 & ~w7288;
assign w3899 = ~w3219 & ~w8046;
assign w3900 = w2557 & ~w14209;
assign w3901 = w8339 & ~w18309;
assign w3902 = ~w2892 & ~w15302;
assign w3903 = w10932 & w1080;
assign w3904 = ~w18030 & ~w16176;
assign w3905 = ~w15999 & ~w17878;
assign w3906 = ~w6751 & ~w18072;
assign w3907 = ~w1443 & ~w15457;
assign w3908 = (w10122 & w1691) | (w10122 & w18733) | (w1691 & w18733);
assign w3909 = ~w1597 & ~w13236;
assign w3910 = w13979 & w3739;
assign w3911 = ~w10546 & ~w13568;
assign w3912 = w2322 & w17251;
assign w3913 = ~w1082 & ~w1545;
assign w3914 = ~w2620 & ~w17346;
assign w3915 = ~w5026 & ~w4685;
assign w3916 = ~w6853 & w17797;
assign w3917 = (~w8203 & ~w3796) | (~w8203 & w11159) | (~w3796 & w11159);
assign w3918 = ~w3276 & ~w18615;
assign w3919 = w14637 & w362;
assign w3920 = ~w19079 & ~w1796;
assign w3921 = a_6 & a_47;
assign w3922 = w16386 & w2373;
assign w3923 = ~w17809 & w9877;
assign w3924 = a_16 & a_60;
assign w3925 = ~w5510 & ~w9135;
assign w3926 = ~w4808 & w12724;
assign w3927 = ~w16055 & w1632;
assign w3928 = w11401 & w11165;
assign w3929 = ~w1057 & w9705;
assign w3930 = w16597 & ~w2919;
assign w3931 = ~w6923 & ~w5642;
assign w3932 = ~w16375 & ~w14172;
assign w3933 = ~w19080 & ~w8707;
assign w3934 = ~w15544 & ~w4349;
assign w3935 = w7877 & ~w3394;
assign w3936 = ~w18532 & ~w7103;
assign w3937 = ~w6059 & ~w8418;
assign w3938 = ~w15989 & ~w15859;
assign w3939 = (w9894 & w15585) | (w9894 & w1626) | (w15585 & w1626);
assign w3940 = w17859 & ~w18844;
assign w3941 = w17065 & ~w6140;
assign w3942 = ~w13369 & ~w12895;
assign w3943 = ~w15915 & ~w11723;
assign w3944 = ~w13851 & w18117;
assign w3945 = w866 & ~w13537;
assign w3946 = ~a_31 & w13854;
assign w3947 = ~w3542 & w4723;
assign w3948 = ~w424 & ~w16876;
assign w3949 = a_4 & a_62;
assign w3950 = ~w3629 & ~w9728;
assign w3951 = ~w11701 & ~w2021;
assign w3952 = (~w1571 & ~w18332) | (~w1571 & w684) | (~w18332 & w684);
assign w3953 = ~w6442 & ~w17080;
assign w3954 = w16637 & ~w554;
assign w3955 = ~w6466 & ~w5310;
assign w3956 = ~w8540 & ~w13378;
assign w3957 = ~w6534 & w8208;
assign w3958 = ~w7180 & ~w1066;
assign w3959 = w18594 & ~w15566;
assign w3960 = (~w10992 & ~w8148) | (~w10992 & w5489) | (~w8148 & w5489);
assign w3961 = (~w5851 & ~w11417) | (~w5851 & w10221) | (~w11417 & w10221);
assign w3962 = w5583 & w17823;
assign w3963 = ~w7204 & ~w4538;
assign w3964 = ~w6233 & ~w5704;
assign w3965 = (~w5495 & w13159) | (~w5495 & w18042) | (w13159 & w18042);
assign w3966 = a_35 & a_55;
assign w3967 = (w7102 & w3085) | (w7102 & w1783) | (w3085 & w1783);
assign w3968 = ~w4063 & ~w13128;
assign w3969 = ~w3715 & ~w8567;
assign w3970 = w3666 & w8634;
assign w3971 = ~w7910 & ~w368;
assign w3972 = ~w10511 & ~w15745;
assign w3973 = w5463 & ~w14207;
assign w3974 = ~w18426 & ~w5294;
assign w3975 = ~w3309 & ~w13743;
assign w3976 = w17224 & ~w6598;
assign w3977 = w11812 & w1338;
assign w3978 = ~w4961 & ~w13383;
assign w3979 = w15806 & w14010;
assign w3980 = w6112 & ~w18063;
assign w3981 = w14678 & ~w7743;
assign w3982 = w18701 & w1022;
assign w3983 = ~w18450 & ~w10163;
assign w3984 = ~w15599 & ~w15254;
assign w3985 = ~w7129 & w1184;
assign w3986 = ~w18918 & ~w10973;
assign w3987 = ~w10664 & ~w1379;
assign w3988 = ~w16392 & ~w17443;
assign w3989 = w16726 & ~w17113;
assign w3990 = w16245 & w10866;
assign w3991 = ~w12536 & ~w14464;
assign w3992 = a_7 & a_59;
assign w3993 = ~w18255 & ~w2265;
assign w3994 = ~w4459 & w1714;
assign w3995 = w5530 & ~w3784;
assign w3996 = a_38 & a_46;
assign w3997 = ~w17416 & ~w3710;
assign w3998 = ~w7071 & ~w7602;
assign w3999 = w4674 & w4271;
assign w4000 = ~w17175 & ~w5801;
assign w4001 = ~w17747 & ~w4443;
assign w4002 = ~w7998 & ~w7394;
assign w4003 = ~w11065 & ~w6895;
assign w4004 = w6745 & w11356;
assign w4005 = ~w5987 & ~w3711;
assign w4006 = w16631 & w16118;
assign w4007 = w14622 & ~w11575;
assign w4008 = ~w12904 & w10382;
assign w4009 = ~w8115 & ~w900;
assign w4010 = ~w9750 & w7847;
assign w4011 = ~w13301 & ~w12349;
assign w4012 = w2359 & ~w10646;
assign w4013 = w10584 & w11993;
assign w4014 = w15219 & ~w9534;
assign w4015 = ~w3915 & w7255;
assign w4016 = w4511 & ~w14350;
assign w4017 = w7156 & ~w2602;
assign w4018 = w331 & w10197;
assign w4019 = w10053 & ~w6570;
assign w4020 = ~w10278 & ~w725;
assign w4021 = ~w351 & w1684;
assign w4022 = ~w13034 & ~w9968;
assign w4023 = ~w2769 & w7128;
assign w4024 = ~w16866 & ~w15127;
assign w4025 = (w7768 & w7864) | (w7768 & w9790) | (w7864 & w9790);
assign w4026 = ~w10651 & w7739;
assign w4027 = a_39 & a_60;
assign w4028 = a_44 & a_49;
assign w4029 = (~w11099 & ~w12625) | (~w11099 & w4416) | (~w12625 & w4416);
assign w4030 = ~w1412 & ~w6498;
assign w4031 = ~w4453 & w13905;
assign w4032 = ~w9508 & ~w9262;
assign w4033 = a_25 & a_47;
assign w4034 = w13086 & w6568;
assign w4035 = ~w8121 & w1168;
assign w4036 = w18096 & w13385;
assign w4037 = ~w11616 & ~w8344;
assign w4038 = ~w8870 & ~w5498;
assign w4039 = ~w534 & ~w3660;
assign w4040 = (w5866 & w12413) | (w5866 & w3889) | (w12413 & w3889);
assign w4041 = w13734 & ~w15851;
assign w4042 = ~w12624 & ~w14033;
assign w4043 = (w794 & w5882) | (w794 & w17616) | (w5882 & w17616);
assign w4044 = ~w11606 & ~w11155;
assign w4045 = a_28 & a_51;
assign w4046 = w5775 & ~w17922;
assign w4047 = w134 & ~w17345;
assign w4048 = ~w3854 & ~w11643;
assign w4049 = w16232 & w9989;
assign w4050 = a_9 & a_15;
assign w4051 = ~w11566 & w11201;
assign w4052 = ~w11761 & w12333;
assign w4053 = ~w18721 & ~w14056;
assign w4054 = ~w6034 & w11175;
assign w4055 = w9170 & w4705;
assign w4056 = w5339 & ~w3515;
assign w4057 = w2593 & ~w17367;
assign w4058 = ~w3230 & w4511;
assign w4059 = w3871 & w9208;
assign w4060 = w17150 & w7160;
assign w4061 = ~w7566 & w13452;
assign w4062 = w9560 & ~w9543;
assign w4063 = ~w2468 & w15634;
assign w4064 = ~w17359 & w10496;
assign w4065 = ~w6519 & ~w15422;
assign w4066 = w5074 & w17101;
assign w4067 = w13186 & w1596;
assign w4068 = ~w1274 & ~w2115;
assign w4069 = w1761 & w9736;
assign w4070 = ~w1852 & ~w5655;
assign w4071 = (~w6477 & ~w493) | (~w6477 & w2805) | (~w493 & w2805);
assign w4072 = w10806 & ~w2569;
assign w4073 = ~w17097 & ~w2169;
assign w4074 = ~w3199 & ~w2285;
assign w4075 = ~w15295 & ~w13755;
assign w4076 = ~w8493 & ~w5460;
assign w4077 = ~w3167 & ~w2813;
assign w4078 = ~w6660 & w19155;
assign w4079 = w6171 & ~w11518;
assign w4080 = w4535 & ~w5018;
assign w4081 = ~w11637 & ~w217;
assign w4082 = (w7341 & w13126) | (w7341 & w746) | (w13126 & w746);
assign w4083 = ~w7524 & ~w9874;
assign w4084 = w12583 & w4571;
assign w4085 = ~w12693 & w18864;
assign w4086 = ~w11532 & w12821;
assign w4087 = w4188 & w5727;
assign w4088 = ~w18307 & ~w18213;
assign w4089 = w12932 & ~w10762;
assign w4090 = ~w3938 & w1822;
assign w4091 = ~w9764 & w10961;
assign w4092 = ~w1942 & ~w15206;
assign w4093 = w853 & ~w14537;
assign w4094 = w9430 & ~w13934;
assign w4095 = ~w13009 & ~w11710;
assign w4096 = ~w16186 & ~w2237;
assign w4097 = a_11 & a_39;
assign w4098 = ~w4516 & ~w13856;
assign w4099 = w10140 & w15726;
assign w4100 = w18014 & w8601;
assign w4101 = ~w16541 & ~w17640;
assign w4102 = ~w3204 & ~w9475;
assign w4103 = ~w17772 & ~w9622;
assign w4104 = ~w14692 & w10771;
assign w4105 = ~w18555 & ~w3258;
assign w4106 = ~w10287 & w10934;
assign w4107 = ~w9238 & ~w2717;
assign w4108 = (~w11308 & ~w2882) | (~w11308 & w3137) | (~w2882 & w3137);
assign w4109 = ~w14571 & ~w3050;
assign w4110 = ~w348 & ~w6657;
assign w4111 = ~w17453 & w15026;
assign w4112 = ~w8382 & w1123;
assign w4113 = ~w9891 & ~w5092;
assign w4114 = a_11 & a_23;
assign w4115 = (w11864 & w2475) | (w11864 & w8361) | (w2475 & w8361);
assign w4116 = a_6 & a_48;
assign w4117 = w8319 & ~w9281;
assign w4118 = w9300 & ~w12542;
assign w4119 = w16639 & ~w4725;
assign w4120 = ~w15665 & ~w5175;
assign w4121 = a_47 & a_60;
assign w4122 = w18131 & ~w18178;
assign w4123 = (w18733 & w17698) | (w18733 & w11068) | (w17698 & w11068);
assign w4124 = ~w16465 & ~w591;
assign w4125 = ~w6658 & ~w12242;
assign w4126 = ~w14885 & ~w13582;
assign w4127 = w7657 & ~w9472;
assign w4128 = w17827 & ~w15678;
assign w4129 = ~w14135 & ~w901;
assign w4130 = ~w8019 & ~w10524;
assign w4131 = ~w10666 & w9213;
assign w4132 = w17438 & ~w4746;
assign w4133 = a_26 & a_48;
assign w4134 = w17184 & ~w17410;
assign w4135 = a_23 & a_34;
assign w4136 = ~w15602 & w10032;
assign w4137 = ~w10805 & ~w7067;
assign w4138 = a_36 & a_63;
assign w4139 = ~w19007 & ~w12523;
assign w4140 = ~w1628 & ~w11094;
assign w4141 = ~w7194 & ~w10429;
assign w4142 = ~w7523 & ~w3150;
assign w4143 = a_38 & a_63;
assign w4144 = ~w15738 & ~w5305;
assign w4145 = ~w6521 & ~w8100;
assign w4146 = ~w8056 & ~w18677;
assign w4147 = ~w18469 & ~w2727;
assign w4148 = ~w5381 & ~w15836;
assign w4149 = w107 & ~w13283;
assign w4150 = w11979 & w17965;
assign w4151 = w18823 & ~w14937;
assign w4152 = a_9 & a_60;
assign w4153 = a_15 & a_46;
assign w4154 = w11536 & ~w6395;
assign w4155 = w12030 & w7350;
assign w4156 = ~w12385 & ~w6636;
assign w4157 = ~w9983 & w11288;
assign w4158 = ~w181 & ~w5776;
assign w4159 = a_17 & a_19;
assign w4160 = ~w14500 & ~w4676;
assign w4161 = (~w9797 & ~w3297) | (~w9797 & w13839) | (~w3297 & w13839);
assign w4162 = ~w11143 & ~w970;
assign w4163 = ~w9204 & ~w17849;
assign w4164 = a_2 & w14127;
assign w4165 = ~w4054 & ~w11082;
assign w4166 = ~w18983 & ~w10756;
assign w4167 = w15167 & w11920;
assign w4168 = ~w8733 & ~w9364;
assign w4169 = ~w14092 & ~w11573;
assign w4170 = (~w2960 & w5978) | (~w2960 & w17597) | (w5978 & w17597);
assign w4171 = ~w4385 & ~w7852;
assign w4172 = ~w15854 & ~w14649;
assign w4173 = ~w6490 & ~w8666;
assign w4174 = w9091 & ~w16552;
assign w4175 = w5216 & ~w14247;
assign w4176 = ~w14015 & w5148;
assign w4177 = w8230 & w399;
assign w4178 = w16236 & ~w9611;
assign w4179 = ~w1100 & w4212;
assign w4180 = a_6 & a_50;
assign w4181 = w2861 & ~w9820;
assign w4182 = ~w1228 & ~w4206;
assign w4183 = w9750 & ~w7847;
assign w4184 = ~w5466 & ~w2575;
assign w4185 = w941 & w15347;
assign w4186 = ~w17068 & w11029;
assign w4187 = ~w813 & ~w2212;
assign w4188 = a_3 & a_25;
assign w4189 = ~w14018 & ~w4956;
assign w4190 = ~w10056 & ~w12224;
assign w4191 = ~w10938 & ~w1536;
assign w4192 = ~w11193 & w14589;
assign w4193 = w18351 & ~w16416;
assign w4194 = ~w16283 & w7559;
assign w4195 = ~w18303 & ~w4230;
assign w4196 = w8625 & w18363;
assign w4197 = ~w5544 & w12028;
assign w4198 = ~w9119 & ~w4600;
assign w4199 = ~w17428 & w12958;
assign w4200 = w19070 & w2895;
assign w4201 = ~w2300 & ~w15268;
assign w4202 = a_25 & a_27;
assign w4203 = ~w2950 & ~w1908;
assign w4204 = ~w5202 & ~w15702;
assign w4205 = w672 & w13871;
assign w4206 = w11599 & ~w7719;
assign w4207 = ~w12977 & ~w11383;
assign w4208 = a_5 & a_53;
assign w4209 = ~w10259 & ~w603;
assign w4210 = ~w19010 & w3580;
assign w4211 = a_11 & a_48;
assign w4212 = ~w16253 & ~w12596;
assign w4213 = ~w1208 & w10300;
assign w4214 = w4733 & ~w1092;
assign w4215 = w12411 & ~w14185;
assign w4216 = ~w11749 & ~w5878;
assign w4217 = ~w18011 & ~w7346;
assign w4218 = ~w1773 & w16830;
assign w4219 = (~w15864 & ~w6148) | (~w15864 & w14693) | (~w6148 & w14693);
assign w4220 = ~w10681 & ~w10972;
assign w4221 = w18723 & w1105;
assign w4222 = ~w2633 & ~w241;
assign w4223 = w15128 & ~w10808;
assign w4224 = ~w1301 & w4217;
assign w4225 = w5095 & ~w12441;
assign w4226 = w15622 & ~w16361;
assign w4227 = a_20 & a_57;
assign w4228 = ~w18554 & ~w5533;
assign w4229 = ~w12722 & ~w8811;
assign w4230 = (w16432 & w13400) | (w16432 & w16401) | (w13400 & w16401);
assign w4231 = a_1 & a_3;
assign w4232 = ~w9718 & w3279;
assign w4233 = (~w14549 & w17825) | (~w14549 & w8529) | (w17825 & w8529);
assign w4234 = w13785 & ~w7339;
assign w4235 = w558 & ~w9113;
assign w4236 = ~w4492 & ~w3072;
assign w4237 = ~w5190 & ~w3233;
assign w4238 = w12301 & w4907;
assign w4239 = ~w16471 & w14730;
assign w4240 = w4889 | w961;
assign w4241 = ~w8060 & ~w11613;
assign w4242 = a_41 & a_57;
assign w4243 = ~w13524 & ~w16260;
assign w4244 = ~w12207 & ~w6083;
assign w4245 = ~w18321 & ~w16573;
assign w4246 = ~w12477 & w10517;
assign w4247 = ~w11970 & ~w17011;
assign w4248 = w13646 & w1411;
assign w4249 = ~w5157 & ~w1169;
assign w4250 = ~w1047 & ~w12763;
assign w4251 = ~w11629 & ~w8022;
assign w4252 = ~w14629 & ~w1425;
assign w4253 = ~w7411 & w8616;
assign w4254 = ~w6168 & ~w3512;
assign w4255 = w11755 & w18040;
assign w4256 = w2379 & w14618;
assign w4257 = a_2 & a_7;
assign w4258 = w13082 & w9025;
assign w4259 = w3489 & ~w6753;
assign w4260 = (w5175 & w6080) | (w5175 & w14257) | (w6080 & w14257);
assign w4261 = w4405 & ~w1531;
assign w4262 = ~w248 & ~w1437;
assign w4263 = ~w17365 & ~w36;
assign w4264 = ~w13267 & w8448;
assign w4265 = ~w4318 & ~w9449;
assign w4266 = ~w4976 & ~w7216;
assign w4267 = a_30 & a_50;
assign w4268 = ~w3724 & ~w19131;
assign w4269 = ~w18101 & ~w12087;
assign w4270 = ~w11211 & ~w7254;
assign w4271 = ~w13635 & ~w2372;
assign w4272 = ~w9690 & ~w2904;
assign w4273 = ~w7117 & ~w9035;
assign w4274 = a_35 & a_63;
assign w4275 = ~w1956 & ~w12237;
assign w4276 = ~w13756 & ~w16342;
assign w4277 = w14910 & w18131;
assign w4278 = ~w4192 & ~w5345;
assign w4279 = (~w10202 & ~w15219) | (~w10202 & w8449) | (~w15219 & w8449);
assign w4280 = ~w11180 & ~w1843;
assign w4281 = ~w17038 & ~w1445;
assign w4282 = ~w16113 & w3274;
assign w4283 = a_44 & a_61;
assign w4284 = ~w11157 & ~w4499;
assign w4285 = ~w17526 & ~w3385;
assign w4286 = w5808 & w9738;
assign w4287 = ~w1466 & ~w18713;
assign w4288 = ~w4467 & ~w3814;
assign w4289 = w7590 & ~w14734;
assign w4290 = w17606 & ~w877;
assign w4291 = ~w12611 & ~w7861;
assign w4292 = ~w6858 & ~w14276;
assign w4293 = ~w13928 & ~w2445;
assign w4294 = a_15 & a_60;
assign w4295 = ~w10597 & ~w14162;
assign w4296 = a_18 & a_63;
assign w4297 = w14660 & ~w17349;
assign w4298 = ~w12108 & ~w1853;
assign w4299 = ~w5818 & ~w6377;
assign w4300 = ~w11330 & ~w5082;
assign w4301 = w6759 & ~w8328;
assign w4302 = ~w10844 & ~w16939;
assign w4303 = ~w12187 & ~w11860;
assign w4304 = ~w7101 & ~w8491;
assign w4305 = ~w9362 & ~w14290;
assign w4306 = ~w10356 & ~w2090;
assign w4307 = ~w13477 & ~w16007;
assign w4308 = a_13 & a_29;
assign w4309 = ~w18012 & ~w1660;
assign w4310 = ~w16864 & ~w11490;
assign w4311 = w16389 & ~w8171;
assign w4312 = w3235 & ~w16269;
assign w4313 = ~w7115 & ~w8058;
assign w4314 = w12893 & ~w9259;
assign w4315 = a_49 & a_50;
assign w4316 = ~w8850 & ~w14576;
assign w4317 = w9774 & w6964;
assign w4318 = w5005 & w18401;
assign w4319 = ~w9836 & ~w13976;
assign w4320 = ~w7784 & ~w10559;
assign w4321 = w7303 & ~w17983;
assign w4322 = ~w2318 & ~w10248;
assign w4323 = ~w10848 & ~w1775;
assign w4324 = w11539 & ~w9987;
assign w4325 = ~w16848 & ~w18541;
assign w4326 = (w4979 & w13082) | (w4979 & w17191) | (w13082 & w17191);
assign w4327 = ~w10260 & ~w12730;
assign w4328 = (~w4570 & ~w9258) | (~w4570 & w2825) | (~w9258 & w2825);
assign w4329 = ~w15756 & w16953;
assign w4330 = ~w3866 & ~w18208;
assign w4331 = ~w575 & ~w4937;
assign w4332 = ~w2380 & ~w287;
assign w4333 = w7941 & w8300;
assign w4334 = ~w1894 & w4542;
assign w4335 = ~w6825 & ~w583;
assign w4336 = w14170 & w9688;
assign w4337 = (~w3154 & ~w13871) | (~w3154 & w15112) | (~w13871 & w15112);
assign w4338 = ~w15138 & ~w4975;
assign w4339 = ~w7674 & ~w2424;
assign w4340 = w14765 & w8425;
assign w4341 = (w1576 & ~w15399) | (w1576 & w10654) | (~w15399 & w10654);
assign w4342 = (~w3500 & ~w14145) | (~w3500 & w14586) | (~w14145 & w14586);
assign w4343 = ~w8362 & w5048;
assign w4344 = ~w17285 & ~w18497;
assign w4345 = ~w12706 & ~w10740;
assign w4346 = w15542 & ~w16973;
assign w4347 = ~w18892 & ~w3793;
assign w4348 = ~w4159 & ~w14251;
assign w4349 = (~w8733 & ~w4168) | (~w8733 & w8795) | (~w4168 & w8795);
assign w4350 = ~w10022 & ~w14258;
assign w4351 = w4846 & w10518;
assign w4352 = (w8965 & w6940) | (w8965 & ~w5108) | (w6940 & ~w5108);
assign w4353 = ~w16611 & w1816;
assign w4354 = ~w16755 & w13261;
assign w4355 = ~w12627 & w10257;
assign w4356 = ~w16564 & w17947;
assign w4357 = ~w5924 & ~w16004;
assign w4358 = w7404 & ~w3761;
assign w4359 = w8468 & w8982;
assign w4360 = ~w345 & ~w7318;
assign w4361 = ~w898 & ~w9381;
assign w4362 = ~w3289 & ~w18081;
assign w4363 = ~w17955 & ~w13096;
assign w4364 = ~w12152 & ~w1875;
assign w4365 = ~w15185 & ~w13628;
assign w4366 = ~w18868 & w15645;
assign w4367 = (w4043 & w9221) | (w4043 & w7943) | (w9221 & w7943);
assign w4368 = ~w8703 & ~w9942;
assign w4369 = ~w14367 & w1787;
assign w4370 = w9768 & w5382;
assign w4371 = ~w7643 & ~w12025;
assign w4372 = ~w3551 & ~w17217;
assign w4373 = a_33 & a_59;
assign w4374 = w15190 & w10344;
assign w4375 = ~w18917 & ~w18550;
assign w4376 = ~w10195 & ~w5080;
assign w4377 = ~w17259 & w11875;
assign w4378 = ~w8054 & w4395;
assign w4379 = a_0 & a_41;
assign w4380 = ~w17613 & ~w12339;
assign w4381 = ~w18373 & ~w11512;
assign w4382 = w10896 & ~w16681;
assign w4383 = w15166 & w16050;
assign w4384 = ~w12911 & ~w8158;
assign w4385 = ~w12632 & ~w5979;
assign w4386 = w11532 & ~w12821;
assign w4387 = ~w6643 & w9951;
assign w4388 = ~w5136 & ~w10288;
assign w4389 = a_17 & a_22;
assign w4390 = ~w6430 & ~w135;
assign w4391 = ~w6839 & w16754;
assign w4392 = ~w4820 & w11450;
assign w4393 = w9654 & ~w10142;
assign w4394 = (~w8530 & ~w10615) | (~w8530 & w5370) | (~w10615 & w5370);
assign w4395 = ~w15930 & ~w9255;
assign w4396 = ~w1678 & w5630;
assign w4397 = w12547 & w5006;
assign w4398 = ~w4188 & ~w5727;
assign w4399 = w2908 & w12630;
assign w4400 = ~w503 & w8978;
assign w4401 = ~w11457 & ~w9665;
assign w4402 = ~w14182 & ~w12929;
assign w4403 = ~w12170 & ~w14649;
assign w4404 = w10357 & ~w17776;
assign w4405 = ~w6657 & ~w15070;
assign w4406 = w12421 & w12996;
assign w4407 = w11291 & ~w1509;
assign w4408 = ~w10693 & ~w2998;
assign w4409 = ~w8723 & ~w11458;
assign w4410 = w11707 & ~w2758;
assign w4411 = ~w538 & ~w1296;
assign w4412 = ~w9573 & ~w10585;
assign w4413 = w8612 & w10728;
assign w4414 = ~w11103 & w2312;
assign w4415 = (w6475 & w3460) | (w6475 & w11038) | (w3460 & w11038);
assign w4416 = ~w17173 & ~w11099;
assign w4417 = ~w14642 & w1920;
assign w4418 = w3285 & w1698;
assign w4419 = w17058 & w13760;
assign w4420 = ~w16284 & ~w11656;
assign w4421 = ~w3443 & ~w12310;
assign w4422 = w1587 & w4432;
assign w4423 = a_34 & a_35;
assign w4424 = ~w15409 & ~w3528;
assign w4425 = ~w16864 & w624;
assign w4426 = ~w18206 & w4597;
assign w4427 = w12296 & ~w4216;
assign w4428 = ~w10388 & ~w8223;
assign w4429 = ~w11709 & ~w26;
assign w4430 = w12558 & ~w3318;
assign w4431 = w290 & w3316;
assign w4432 = ~w5813 & ~w17723;
assign w4433 = ~w13155 & w2770;
assign w4434 = w17282 & ~w10347;
assign w4435 = w7688 & w17417;
assign w4436 = ~w16757 & ~w14317;
assign w4437 = ~w16601 & w1834;
assign w4438 = a_11 & a_22;
assign w4439 = ~w2502 & w11201;
assign w4440 = w11910 & ~w278;
assign w4441 = ~w11786 & ~w18661;
assign w4442 = w15833 & ~w5724;
assign w4443 = ~w7488 & w19129;
assign w4444 = ~w12769 & w178;
assign w4445 = ~w191 & ~w5891;
assign w4446 = ~w1247 & ~w3848;
assign w4447 = w17375 & ~w5678;
assign w4448 = w67 & ~w16102;
assign w4449 = ~w3226 & ~w16202;
assign w4450 = w10236 & ~w10806;
assign w4451 = ~w13426 & ~w883;
assign w4452 = ~w16499 & ~w9276;
assign w4453 = ~w13022 & ~w13916;
assign w4454 = ~w4559 & w6288;
assign w4455 = (w6567 & ~w12288) | (w6567 & w4123) | (~w12288 & w4123);
assign w4456 = w12781 & ~w9984;
assign w4457 = ~w17491 & w4350;
assign w4458 = ~w1641 & ~w18905;
assign w4459 = ~w7535 & ~w639;
assign w4460 = w2956 & w9267;
assign w4461 = a_17 & a_49;
assign w4462 = ~w17755 & ~w144;
assign w4463 = ~w6702 & w4882;
assign w4464 = ~w1128 & ~w11367;
assign w4465 = w8685 & ~w11612;
assign w4466 = ~w9999 & w16491;
assign w4467 = ~w13054 & w14466;
assign w4468 = w11266 & w18365;
assign w4469 = w13095 & w17998;
assign w4470 = ~w14535 & ~w9484;
assign w4471 = ~w10185 & ~w9128;
assign w4472 = ~w14741 & ~w11503;
assign w4473 = w1964 & ~w12881;
assign w4474 = (~w3772 & ~w13661) | (~w3772 & w471) | (~w13661 & w471);
assign w4475 = w10912 & ~w18281;
assign w4476 = ~w8768 & w6993;
assign w4477 = ~w12876 & ~w18039;
assign w4478 = a_3 & a_47;
assign w4479 = ~w17302 & ~w17153;
assign w4480 = ~w481 & w10962;
assign w4481 = ~w15921 & ~w7349;
assign w4482 = ~w17133 & ~w5609;
assign w4483 = a_4 & a_27;
assign w4484 = w8675 & w8142;
assign w4485 = ~w11439 & w3904;
assign w4486 = ~w177 & ~w4015;
assign w4487 = w2579 & ~w15527;
assign w4488 = w17138 & ~w2476;
assign w4489 = ~w8398 & ~w7125;
assign w4490 = ~w14428 & ~w7121;
assign w4491 = ~w2724 & ~w2216;
assign w4492 = ~w2716 & ~w13626;
assign w4493 = w5499 & ~w17846;
assign w4494 = ~w4897 & ~w17872;
assign w4495 = ~w10321 & ~w12132;
assign w4496 = a_24 & a_60;
assign w4497 = ~w11366 & w15039;
assign w4498 = ~w18124 & ~w11635;
assign w4499 = ~w15411 & ~w12584;
assign w4500 = ~w10395 & ~w6480;
assign w4501 = w10382 & ~w4367;
assign w4502 = a_35 & a_42;
assign w4503 = ~w12285 & w17503;
assign w4504 = w16478 & w14090;
assign w4505 = w14132 & ~w9995;
assign w4506 = ~w9464 & ~w6173;
assign w4507 = (~w7768 & w2338) | (~w7768 & w9622) | (w2338 & w9622);
assign w4508 = ~w16883 & ~w1644;
assign w4509 = ~w16987 & ~w8040;
assign w4510 = ~w2097 & ~w11734;
assign w4511 = ~w7097 & ~w13968;
assign w4512 = a_3 & a_22;
assign w4513 = ~w6154 & ~w777;
assign w4514 = ~w18203 & ~w1088;
assign w4515 = ~w3289 & w1554;
assign w4516 = w10865 & ~w15341;
assign w4517 = (w6553 & w11366) | (w6553 & w15412) | (w11366 & w15412);
assign w4518 = w2583 & ~w4584;
assign w4519 = ~w10974 & ~w1096;
assign w4520 = a_15 & a_35;
assign w4521 = w15042 & ~w606;
assign w4522 = (w15337 & w2769) | (w15337 & w12454) | (w2769 & w12454);
assign w4523 = ~w19038 & ~w1248;
assign w4524 = ~w6422 & ~w9652;
assign w4525 = ~w18906 & ~w9046;
assign w4526 = w11464 & w15525;
assign w4527 = ~w17607 & ~w14869;
assign w4528 = ~w6679 & ~w11792;
assign w4529 = ~w4312 & w8780;
assign w4530 = (w2769 & w2824) | (w2769 & w14146) | (w2824 & w14146);
assign w4531 = ~w14231 & ~w2213;
assign w4532 = ~w11387 & ~w17208;
assign w4533 = ~w10873 & w8747;
assign w4534 = ~w9139 & ~w682;
assign w4535 = a_20 & a_39;
assign w4536 = ~w13736 & ~w10407;
assign w4537 = ~w8732 & ~w17601;
assign w4538 = (~w4287 & w12089) | (~w4287 & w12773) | (w12089 & w12773);
assign w4539 = a_11 & a_20;
assign w4540 = w3988 & ~w13789;
assign w4541 = ~w14780 & ~w11320;
assign w4542 = ~w9291 & w5949;
assign w4543 = ~w3993 & ~w11900;
assign w4544 = w6529 & ~w14559;
assign w4545 = ~w16067 & ~w11207;
assign w4546 = ~w7385 & ~w10573;
assign w4547 = (w8008 & w10330) | (w8008 & w18726) | (w10330 & w18726);
assign w4548 = ~w13118 & ~w12241;
assign w4549 = a_40 & a_62;
assign w4550 = ~w14725 & w15815;
assign w4551 = w143 & ~w16751;
assign w4552 = ~w11684 & ~w12951;
assign w4553 = ~w6605 & ~w8608;
assign w4554 = ~w17938 & ~w6551;
assign w4555 = w15629 & ~w8128;
assign w4556 = (~w10167 & ~w11492) | (~w10167 & w7112) | (~w11492 & w7112);
assign w4557 = ~w17168 & ~w7626;
assign w4558 = ~w1116 & ~w14573;
assign w4559 = ~w15988 & w7878;
assign w4560 = ~w4575 & ~w3420;
assign w4561 = w17721 & w11784;
assign w4562 = ~w12456 & w6794;
assign w4563 = ~w13853 & w17354;
assign w4564 = w2906 & w14518;
assign w4565 = ~w13259 & ~w6939;
assign w4566 = ~w1563 & ~w2899;
assign w4567 = ~w18989 & ~w14187;
assign w4568 = w17201 & ~w14064;
assign w4569 = ~w2533 & ~w9218;
assign w4570 = ~w7973 & ~w12847;
assign w4571 = (~w359 & w8458) | (~w359 & w8755) | (w8458 & w8755);
assign w4572 = w5402 & ~w3150;
assign w4573 = a_8 & a_22;
assign w4574 = ~w7462 & w9077;
assign w4575 = ~w18966 & ~w17614;
assign w4576 = w4281 & w13896;
assign w4577 = ~w12370 & ~w3878;
assign w4578 = w13371 & w5948;
assign w4579 = ~w6487 & ~w15297;
assign w4580 = ~w9404 & ~w529;
assign w4581 = ~w15684 & ~w8206;
assign w4582 = ~w2846 & ~w15703;
assign w4583 = ~w12509 & w11421;
assign w4584 = ~w2414 & ~w13885;
assign w4585 = a_48 & a_51;
assign w4586 = (~w4791 & w10601) | (~w4791 & w2219) | (w10601 & w2219);
assign w4587 = w5982 & w19050;
assign w4588 = w8862 & w11019;
assign w4589 = ~w3964 & ~w10730;
assign w4590 = a_13 & a_34;
assign w4591 = w1575 & ~w16668;
assign w4592 = ~w1998 & ~w7537;
assign w4593 = w7493 & w3032;
assign w4594 = ~w16022 & ~w8618;
assign w4595 = ~w11779 & w15559;
assign w4596 = w1862 & ~w18519;
assign w4597 = ~w3295 & ~w8948;
assign w4598 = a_11 & a_40;
assign w4599 = ~w16372 & ~w930;
assign w4600 = a_20 & a_50;
assign w4601 = w1515 & ~w571;
assign w4602 = ~w11429 & w14027;
assign w4603 = ~w9884 & ~w15331;
assign w4604 = (~w14064 & ~w7926) | (~w14064 & w4568) | (~w7926 & w4568);
assign w4605 = (~w8530 & ~w7544) | (~w8530 & w10562) | (~w7544 & w10562);
assign w4606 = ~w17955 & ~w14148;
assign w4607 = ~w14217 & w3328;
assign w4608 = ~w1019 & w16772;
assign w4609 = ~w3183 & ~w3130;
assign w4610 = a_12 & a_39;
assign w4611 = ~w14131 & ~w6443;
assign w4612 = ~w8116 & w4938;
assign w4613 = ~w9417 & ~w5070;
assign w4614 = w330 & ~w19084;
assign w4615 = w4772 & ~w11772;
assign w4616 = ~w9576 & ~w2932;
assign w4617 = w4009 & w19076;
assign w4618 = w10873 & w3624;
assign w4619 = ~w4419 & ~w6888;
assign w4620 = ~w986 & ~w12979;
assign w4621 = a_26 & a_51;
assign w4622 = w4872 & ~w9164;
assign w4623 = ~w5941 & ~w14477;
assign w4624 = ~w15291 & ~w4121;
assign w4625 = w16022 & w8618;
assign w4626 = a_52 & a_62;
assign w4627 = w10626 & ~w7996;
assign w4628 = w13354 & ~w251;
assign w4629 = ~w5056 & ~w855;
assign w4630 = ~w10581 & w18153;
assign w4631 = ~w6148 & w2776;
assign w4632 = ~w15789 & w8067;
assign w4633 = a_19 & a_34;
assign w4634 = ~w322 & ~w3131;
assign w4635 = ~w13447 & ~w3206;
assign w4636 = ~w19042 & ~w5184;
assign w4637 = ~w3195 & ~w10411;
assign w4638 = ~w13513 & w5257;
assign w4639 = ~w13388 & ~w12749;
assign w4640 = (~w1597 & ~w3909) | (~w1597 & w15811) | (~w3909 & w15811);
assign w4641 = ~w18264 & ~w6436;
assign w4642 = w9286 & ~w35;
assign w4643 = ~w2153 & ~w9998;
assign w4644 = ~w1764 & ~w18197;
assign w4645 = ~w8176 & w16237;
assign w4646 = w3936 & w11158;
assign w4647 = w3582 & w5907;
assign w4648 = w6447 & w13478;
assign w4649 = ~w5691 & ~w18597;
assign w4650 = a_15 & a_47;
assign w4651 = w8474 & w10299;
assign w4652 = ~w2791 & ~w9150;
assign w4653 = ~w17046 & ~w8963;
assign w4654 = w17785 & ~w13370;
assign w4655 = w7120 & w16408;
assign w4656 = ~w17762 & w1547;
assign w4657 = ~w18451 & ~w1282;
assign w4658 = a_23 & a_55;
assign w4659 = w18034 & w5034;
assign w4660 = w10376 & w10697;
assign w4661 = w16788 & ~w15805;
assign w4662 = a_26 & a_56;
assign w4663 = w1220 & w950;
assign w4664 = ~w11085 & ~w9545;
assign w4665 = ~w2602 & ~w2288;
assign w4666 = ~w11125 & ~w10814;
assign w4667 = ~w1488 & ~w13455;
assign w4668 = ~w1737 & ~w766;
assign w4669 = ~w853 & w14537;
assign w4670 = ~w7871 & w16117;
assign w4671 = ~w7478 & w14466;
assign w4672 = ~w17656 & w8676;
assign w4673 = a_19 & a_41;
assign w4674 = ~w18380 & ~w7838;
assign w4675 = ~w2966 & ~w378;
assign w4676 = ~w17836 & ~w12162;
assign w4677 = a_7 & a_46;
assign w4678 = ~w12854 & ~w4115;
assign w4679 = ~w3148 & ~w6016;
assign w4680 = w10392 & ~w18638;
assign w4681 = ~w3607 & ~w9325;
assign w4682 = ~w3198 & ~w14275;
assign w4683 = ~w15806 & ~w14010;
assign w4684 = w5100 & w11796;
assign w4685 = ~w16084 & ~w16393;
assign w4686 = ~w2860 & ~w14557;
assign w4687 = a_1 & a_36;
assign w4688 = w6756 & ~w13250;
assign w4689 = ~w7916 & ~w10748;
assign w4690 = ~w1208 & ~w10159;
assign w4691 = ~w18100 & ~w13991;
assign w4692 = a_20 & a_44;
assign w4693 = w17491 & ~w4350;
assign w4694 = ~w1722 & ~w5118;
assign w4695 = ~w10751 & ~w13620;
assign w4696 = w9740 & w11593;
assign w4697 = w9943 & ~w4323;
assign w4698 = w11230 & ~w15277;
assign w4699 = w12221 & w8847;
assign w4700 = (~w4501 & w2769) | (~w4501 & w12287) | (w2769 & w12287);
assign w4701 = ~w14235 & w18425;
assign w4702 = ~w2769 & w14268;
assign w4703 = ~w16766 & ~w17766;
assign w4704 = (w5866 & w17854) | (w5866 & w10966) | (w17854 & w10966);
assign w4705 = a_14 & a_24;
assign w4706 = a_22 & a_44;
assign w4707 = w2729 & ~w12620;
assign w4708 = ~w1452 & w3415;
assign w4709 = ~w14144 & ~w6663;
assign w4710 = w16357 & ~w15063;
assign w4711 = ~w9727 & ~w5098;
assign w4712 = ~w6914 & ~w17427;
assign w4713 = w9540 & w6222;
assign w4714 = a_24 & a_48;
assign w4715 = ~w1453 & ~w4729;
assign w4716 = ~w13795 & w9951;
assign w4717 = ~w4847 & ~w10555;
assign w4718 = ~w10078 & ~w17724;
assign w4719 = ~w1154 & w12384;
assign w4720 = w3273 & ~w9552;
assign w4721 = ~w8756 & ~w12347;
assign w4722 = ~w8574 & ~w14159;
assign w4723 = ~w10324 & ~w15672;
assign w4724 = ~a_18 & w13356;
assign w4725 = ~w7981 & ~w4294;
assign w4726 = ~w6588 & ~w2804;
assign w4727 = ~w420 & w3215;
assign w4728 = w4322 & ~w3264;
assign w4729 = ~w17327 & w5585;
assign w4730 = ~w18466 & ~w16024;
assign w4731 = w7020 & ~w16714;
assign w4732 = w5298 & w7224;
assign w4733 = ~w17288 & ~w18080;
assign w4734 = ~w9600 & ~w3939;
assign w4735 = ~w1354 & ~w3449;
assign w4736 = ~w6302 & ~w4340;
assign w4737 = ~w16678 & ~w10761;
assign w4738 = ~w7900 & ~w12399;
assign w4739 = ~w13769 & ~w19121;
assign w4740 = ~w1250 & w10816;
assign w4741 = w9937 & ~w11043;
assign w4742 = ~w10667 & ~w11801;
assign w4743 = (~w18824 & ~w3267) | (~w18824 & w1349) | (~w3267 & w1349);
assign w4744 = a_1 & a_40;
assign w4745 = ~w13732 & w5076;
assign w4746 = ~w4398 & ~w4087;
assign w4747 = (~w14483 & ~w7119) | (~w14483 & w7619) | (~w7119 & w7619);
assign w4748 = ~w11849 & ~w13676;
assign w4749 = a_24 & a_47;
assign w4750 = a_6 & a_23;
assign w4751 = w13979 & w12878;
assign w4752 = w1737 & w17958;
assign w4753 = ~w11938 & ~w9168;
assign w4754 = w7111 & ~w12998;
assign w4755 = ~w12124 & ~w15082;
assign w4756 = ~w15398 & ~w15866;
assign w4757 = w14126 & w1326;
assign w4758 = ~w12157 & ~w17092;
assign w4759 = w18814 & w16565;
assign w4760 = w15976 & w14428;
assign w4761 = ~w5592 & ~w9762;
assign w4762 = ~w1147 & ~w14694;
assign w4763 = ~w3315 & ~w1049;
assign w4764 = (~w16660 & ~w4812) | (~w16660 & w11830) | (~w4812 & w11830);
assign w4765 = ~w14797 & ~w8863;
assign w4766 = ~w12782 & ~w722;
assign w4767 = ~w15336 & w10687;
assign w4768 = ~w11003 & w11231;
assign w4769 = ~w4681 & ~w9779;
assign w4770 = ~w12631 & ~w14647;
assign w4771 = ~a_5 & ~w12021;
assign w4772 = a_22 & a_57;
assign w4773 = ~w14910 & w1791;
assign w4774 = (~w10856 & ~w6546) | (~w10856 & w6744) | (~w6546 & w6744);
assign w4775 = (~w3671 & ~w6923) | (~w3671 & w10526) | (~w6923 & w10526);
assign w4776 = ~w2841 & ~w15142;
assign w4777 = ~w14139 & ~w12068;
assign w4778 = w9700 & ~w9081;
assign w4779 = w12258 | w1540;
assign w4780 = ~w4583 & w4355;
assign w4781 = ~w12704 & ~w9639;
assign w4782 = w15005 & w10113;
assign w4783 = w9678 & ~w6894;
assign w4784 = ~w13161 & w16908;
assign w4785 = ~w17195 & ~w9459;
assign w4786 = ~w16247 & ~w9734;
assign w4787 = ~w10587 & ~w17174;
assign w4788 = ~w18777 & ~w136;
assign w4789 = ~w8196 & ~w14437;
assign w4790 = ~w13913 & ~w10071;
assign w4791 = (~w10880 & ~w7361) | (~w10880 & w9242) | (~w7361 & w9242);
assign w4792 = ~w3327 & ~w16425;
assign w4793 = a_27 & a_29;
assign w4794 = ~w8833 & ~w14545;
assign w4795 = ~w341 & w765;
assign w4796 = ~w4886 & ~w7126;
assign w4797 = ~w17178 & ~w8342;
assign w4798 = ~w8669 & ~w17514;
assign w4799 = ~w10410 & ~w3919;
assign w4800 = a_28 & a_30;
assign w4801 = w9712 & w128;
assign w4802 = w11080 & ~w3028;
assign w4803 = w8819 & ~w16850;
assign w4804 = a_47 & a_62;
assign w4805 = w5011 & ~w15016;
assign w4806 = ~w13582 & ~w15670;
assign w4807 = ~w3962 & w3480;
assign w4808 = ~w2221 & w13828;
assign w4809 = w16636 & w6989;
assign w4810 = ~w11504 & w17713;
assign w4811 = ~w12965 & ~w7634;
assign w4812 = ~w16660 & ~w13145;
assign w4813 = a_13 & a_19;
assign w4814 = w16882 & ~w2729;
assign w4815 = ~w8243 & w9269;
assign w4816 = w14244 & w14856;
assign w4817 = ~w11230 & w15277;
assign w4818 = ~w3533 & w13974;
assign w4819 = w1677 & w8810;
assign w4820 = ~w2283 & ~w7006;
assign w4821 = ~w17362 & w13577;
assign w4822 = ~w4314 & ~w18901;
assign w4823 = ~w5303 & ~w5650;
assign w4824 = ~w5211 & ~w16644;
assign w4825 = ~w10357 & w17776;
assign w4826 = ~w9172 & w2363;
assign w4827 = w2385 & w17759;
assign w4828 = ~w2080 & w4636;
assign w4829 = ~w1712 & ~w13682;
assign w4830 = a_12 & a_63;
assign w4831 = ~w5915 & ~w14032;
assign w4832 = ~w14548 & ~w2527;
assign w4833 = (~w879 & ~w14623) | (~w879 & w414) | (~w14623 & w414);
assign w4834 = ~w13617 & ~w3831;
assign w4835 = w15593 & ~w7841;
assign w4836 = w9079 & ~w2795;
assign w4837 = ~w3795 & w556;
assign w4838 = a_1 & a_55;
assign w4839 = w11178 & ~w80;
assign w4840 = w11798 & w6827;
assign w4841 = ~w15524 & ~w7079;
assign w4842 = ~w7907 & ~w9059;
assign w4843 = w9995 & ~w6152;
assign w4844 = (~w14829 & ~w14539) | (~w14829 & w13817) | (~w14539 & w13817);
assign w4845 = ~w9909 & ~w10427;
assign w4846 = ~w11859 & ~w14069;
assign w4847 = ~w14872 & ~w9848;
assign w4848 = w3227 & ~w1335;
assign w4849 = a_18 & a_31;
assign w4850 = ~w11879 & ~w360;
assign w4851 = ~w10646 & ~w10154;
assign w4852 = ~w11372 & ~w13050;
assign w4853 = ~w2197 & ~w8159;
assign w4854 = w6248 & ~w7077;
assign w4855 = ~w5204 & ~w12172;
assign w4856 = a_37 & a_45;
assign w4857 = ~w11556 & ~w16939;
assign w4858 = w10356 & ~w11980;
assign w4859 = ~w11385 & ~w12266;
assign w4860 = ~w3337 & ~w1807;
assign w4861 = ~w16379 & w11738;
assign w4862 = ~w17129 & ~w16696;
assign w4863 = w4616 & w10310;
assign w4864 = ~w13813 & ~w2802;
assign w4865 = w7284 & ~w17455;
assign w4866 = ~w12628 & ~w2893;
assign w4867 = a_14 & a_16;
assign w4868 = w15567 & ~w3365;
assign w4869 = w10294 & w18475;
assign w4870 = ~w14658 & ~w5392;
assign w4871 = ~w15382 & ~w14190;
assign w4872 = a_10 & a_56;
assign w4873 = (~w18555 & ~w4105) | (~w18555 & w13019) | (~w4105 & w13019);
assign w4874 = ~w2845 & ~w13048;
assign w4875 = ~w4593 & ~w4426;
assign w4876 = w4310 & ~w624;
assign w4877 = (~w16751 & ~w8641) | (~w16751 & w4551) | (~w8641 & w4551);
assign w4878 = ~w4190 & ~w15094;
assign w4879 = ~w1874 & ~w17105;
assign w4880 = a_34 & a_43;
assign w4881 = ~w9571 & ~w14193;
assign w4882 = ~w15191 & ~w10184;
assign w4883 = (~w13364 & ~w7830) | (~w13364 & w14445) | (~w7830 & w14445);
assign w4884 = ~w13484 & w4236;
assign w4885 = w9806 & w1553;
assign w4886 = ~w459 & ~w18107;
assign w4887 = w4316 & ~w1971;
assign w4888 = w929 & ~w8309;
assign w4889 = (w15755 & w6221) | (w15755 & w17353) | (w6221 & w17353);
assign w4890 = ~w11825 & ~w76;
assign w4891 = a_21 & a_48;
assign w4892 = w1575 & w16187;
assign w4893 = ~w10327 & ~w17603;
assign w4894 = a_8 & a_34;
assign w4895 = ~w639 & ~w10521;
assign w4896 = a_22 & a_31;
assign w4897 = w6181 & w15809;
assign w4898 = ~w1667 & ~w9675;
assign w4899 = ~w2734 & w5901;
assign w4900 = ~w17518 & w2140;
assign w4901 = ~w4205 & ~w6788;
assign w4902 = ~w9371 & w16525;
assign w4903 = ~w18351 & w16416;
assign w4904 = ~w7490 & ~w11543;
assign w4905 = ~w1669 & ~w8364;
assign w4906 = ~w7101 & ~w11443;
assign w4907 = a_5 & a_24;
assign w4908 = w7485 & ~w10438;
assign w4909 = w11023 & ~w4870;
assign w4910 = (~w7725 & ~w11776) | (~w7725 & w946) | (~w11776 & w946);
assign w4911 = w16565 & ~w5154;
assign w4912 = ~w2619 & ~w4044;
assign w4913 = w7180 & w14457;
assign w4914 = w4747 & ~w16832;
assign w4915 = ~w14313 & w16117;
assign w4916 = a_49 & a_54;
assign w4917 = w6153 & w9228;
assign w4918 = ~w8192 & ~w18840;
assign w4919 = w7617 & ~w8170;
assign w4920 = ~w18342 & ~w12351;
assign w4921 = a_11 & a_24;
assign w4922 = (w4900 & w63) | (w4900 & w18619) | (w63 & w18619);
assign w4923 = a_1 & a_7;
assign w4924 = w2642 & ~w2114;
assign w4925 = ~w16123 & ~w13193;
assign w4926 = w16246 & w14138;
assign w4927 = ~w3494 & ~w5149;
assign w4928 = w9835 & ~w1456;
assign w4929 = a_9 & a_18;
assign w4930 = ~w18580 & w5600;
assign w4931 = ~w15125 & ~w12437;
assign w4932 = w13459 & ~w687;
assign w4933 = w8640 & w6666;
assign w4934 = ~w11262 & w7682;
assign w4935 = (a_49 & w16565) | (a_49 & w10627) | (w16565 & w10627);
assign w4936 = ~w7958 & ~w1193;
assign w4937 = w17062 & w3191;
assign w4938 = ~w8484 & ~w1021;
assign w4939 = a_7 & a_29;
assign w4940 = ~w6026 & ~w5277;
assign w4941 = ~w7692 & ~w15468;
assign w4942 = (w11687 & ~w14279) | (w11687 & w3053) | (~w14279 & w3053);
assign w4943 = (w16374 & w3452) | (w16374 & w8365) | (w3452 & w8365);
assign w4944 = ~w8679 & ~w8867;
assign w4945 = ~w11609 & ~w7277;
assign w4946 = a_51 & a_60;
assign w4947 = w6934 & ~w2654;
assign w4948 = ~w18059 & ~w18978;
assign w4949 = ~w7692 & ~w5286;
assign w4950 = a_27 & a_41;
assign w4951 = ~w4046 & ~w10697;
assign w4952 = ~w16900 & ~w2023;
assign w4953 = (~w9571 & w14130) | (~w9571 & w7036) | (w14130 & w7036);
assign w4954 = w17638 & ~w6972;
assign w4955 = w16186 & w2237;
assign w4956 = ~w5188 & ~w18785;
assign w4957 = a_25 & a_39;
assign w4958 = ~w8665 & w14519;
assign w4959 = w3874 & w2494;
assign w4960 = (w9221 & w4240) | (w9221 & w3738) | (w4240 & w3738);
assign w4961 = w18437 & ~w14332;
assign w4962 = w834 & w6283;
assign w4963 = w10995 & w18451;
assign w4964 = ~w5938 & ~w5385;
assign w4965 = (~w2105 & ~w12561) | (~w2105 & w1136) | (~w12561 & w1136);
assign w4966 = w8341 & ~w16711;
assign w4967 = ~w18990 & w12699;
assign w4968 = w15777 & ~w12148;
assign w4969 = ~w14662 & ~w16472;
assign w4970 = ~w3939 & ~w5319;
assign w4971 = w2045 & ~w5227;
assign w4972 = ~w10138 & w8758;
assign w4973 = ~w18789 & w1823;
assign w4974 = ~w2481 & ~w12837;
assign w4975 = ~w4045 & w18274;
assign w4976 = a_3 & a_31;
assign w4977 = (w2448 & w10349) | (w2448 & w2712) | (w10349 & w2712);
assign w4978 = ~w11047 & ~w1512;
assign w4979 = ~w9369 & ~w16700;
assign w4980 = ~w2119 & w15393;
assign w4981 = ~w16384 & w14866;
assign w4982 = w6056 & w10935;
assign w4983 = ~w527 & w1592;
assign w4984 = ~w13505 & ~w10047;
assign w4985 = a_62 & w15910;
assign w4986 = ~w7015 & w11948;
assign w4987 = ~w12461 & ~w659;
assign w4988 = ~w14940 & ~w7175;
assign w4989 = a_41 & a_45;
assign w4990 = ~w12009 & ~w5421;
assign w4991 = ~w16822 & ~w10309;
assign w4992 = ~w10377 & ~w3948;
assign w4993 = ~w12094 & ~w18269;
assign w4994 = ~w16468 & ~w1187;
assign w4995 = w13343 & w18182;
assign w4996 = a_23 & a_46;
assign w4997 = a_22 & a_55;
assign w4998 = ~w12844 & ~w13548;
assign w4999 = ~w15015 & ~w9855;
assign w5000 = w14608 & ~w15751;
assign w5001 = (a_43 & w12497) | (a_43 & w18896) | (w12497 & w18896);
assign w5002 = ~w15577 & w12250;
assign w5003 = ~w17450 & ~w17924;
assign w5004 = ~w11161 & w12640;
assign w5005 = ~w4013 & ~w5208;
assign w5006 = ~w2647 & ~w5210;
assign w5007 = ~w13933 & ~w14072;
assign w5008 = ~w17766 & w273;
assign w5009 = a_21 & a_53;
assign w5010 = ~w11496 & w2030;
assign w5011 = ~w1964 & w12881;
assign w5012 = (w8058 & w1062) | (w8058 & w11325) | (w1062 & w11325);
assign w5013 = ~w17096 & w16377;
assign w5014 = a_4 & a_34;
assign w5015 = w12157 & w17092;
assign w5016 = ~w9768 & ~w5382;
assign w5017 = a_35 & a_52;
assign w5018 = ~w17399 & ~w13247;
assign w5019 = ~w18933 & ~w11234;
assign w5020 = ~w8424 & ~w17911;
assign w5021 = ~w9476 & ~w3546;
assign w5022 = ~w10080 & ~w9184;
assign w5023 = a_39 & a_41;
assign w5024 = ~w13678 & w19112;
assign w5025 = ~w1779 & ~w13865;
assign w5026 = ~w2796 & ~w4300;
assign w5027 = ~w13919 & ~w16771;
assign w5028 = ~w13017 & ~w1199;
assign w5029 = ~w7120 & ~w16408;
assign w5030 = a_7 & a_30;
assign w5031 = ~w2648 & ~w17644;
assign w5032 = ~w15358 & ~w8627;
assign w5033 = ~w18762 & ~w1330;
assign w5034 = a_29 & a_50;
assign w5035 = ~w16198 & ~w15498;
assign w5036 = ~w1633 & ~w4819;
assign w5037 = ~w8687 & ~w11241;
assign w5038 = a_4 & a_16;
assign w5039 = w17121 & ~w15995;
assign w5040 = ~w4502 & w4990;
assign w5041 = ~w12633 & ~w3108;
assign w5042 = w11374 & ~w10123;
assign w5043 = ~w8681 & ~w2181;
assign w5044 = ~w1831 & ~w2311;
assign w5045 = (~w1465 & ~w940) | (~w1465 & w7697) | (~w940 & w7697);
assign w5046 = a_49 & a_59;
assign w5047 = ~w2707 & ~w13167;
assign w5048 = ~w62 & ~w6045;
assign w5049 = w5893 & ~w11894;
assign w5050 = w15812 & ~w8017;
assign w5051 = (~w18388 & ~w15198) | (~w18388 & w10160) | (~w15198 & w10160);
assign w5052 = ~w5266 & ~w6704;
assign w5053 = ~w15814 & ~w5079;
assign w5054 = ~w10230 & w18204;
assign w5055 = (~w4925 & w4453) | (~w4925 & w1828) | (w4453 & w1828);
assign w5056 = w157 & ~w19002;
assign w5057 = w419 & ~w8187;
assign w5058 = w16085 & w2584;
assign w5059 = ~w14105 & ~w8808;
assign w5060 = w10010 & ~w6526;
assign w5061 = ~w7743 & ~w12448;
assign w5062 = ~w5715 & w3342;
assign w5063 = ~w11307 & ~w15775;
assign w5064 = ~w18323 & ~w13458;
assign w5065 = w14928 & ~w3017;
assign w5066 = (~w5163 & ~w13195) | (~w5163 & w5766) | (~w13195 & w5766);
assign w5067 = ~w18959 & ~w7670;
assign w5068 = ~w9118 & ~w10656;
assign w5069 = ~w8852 & ~w18047;
assign w5070 = ~w10885 & w14743;
assign w5071 = ~w19053 & ~w9641;
assign w5072 = ~w13269 & ~w9837;
assign w5073 = ~w10337 & w9993;
assign w5074 = w4331 & w7348;
assign w5075 = a_10 & a_30;
assign w5076 = ~w59 & ~w3315;
assign w5077 = (~w10222 & ~w826) | (~w10222 & w39) | (~w826 & w39);
assign w5078 = a_29 & a_46;
assign w5079 = w15114 & w17435;
assign w5080 = ~w14940 & ~w2273;
assign w5081 = a_13 & a_60;
assign w5082 = ~w17702 & ~w16454;
assign w5083 = ~w2025 & ~w1815;
assign w5084 = ~w14506 & ~w4020;
assign w5085 = w2878 & ~w10141;
assign w5086 = ~w6511 & ~w10742;
assign w5087 = ~w1538 & ~w16832;
assign w5088 = w14881 & w981;
assign w5089 = ~w3292 & ~w3951;
assign w5090 = ~w4982 & ~w6944;
assign w5091 = (~w14148 & ~w13096) | (~w14148 & w4606) | (~w13096 & w4606);
assign w5092 = ~w6187 & w14960;
assign w5093 = a_35 & a_48;
assign w5094 = ~w2182 & w10800;
assign w5095 = a_50 & a_63;
assign w5096 = ~w9520 & ~w17561;
assign w5097 = ~w17652 & ~w69;
assign w5098 = ~w7058 & ~w2241;
assign w5099 = w1428 & w6240;
assign w5100 = ~w9551 & ~w12195;
assign w5101 = ~w2331 & ~w8227;
assign w5102 = a_18 & a_45;
assign w5103 = ~w10082 & ~w4207;
assign w5104 = (w4960 & w2769) | (w4960 & w3774) | (w2769 & w3774);
assign w5105 = ~w5711 & ~w4576;
assign w5106 = w3009 & ~w8556;
assign w5107 = w4776 & ~w12440;
assign w5108 = ~w3932 & w7211;
assign w5109 = a_4 & a_7;
assign w5110 = ~w6360 & ~w8719;
assign w5111 = ~w7570 & ~w2855;
assign w5112 = a_1 & a_27;
assign w5113 = ~w10978 & ~w6384;
assign w5114 = w7305 & ~w13577;
assign w5115 = ~w695 & w4445;
assign w5116 = ~w12587 & ~w9739;
assign w5117 = w15867 & ~w8195;
assign w5118 = ~w14550 & ~w17274;
assign w5119 = ~w12809 & ~w2610;
assign w5120 = w581 & ~w2659;
assign w5121 = w351 & ~w1684;
assign w5122 = ~w13805 & w11135;
assign w5123 = a_10 & a_50;
assign w5124 = w14360 & w15401;
assign w5125 = ~w14361 & w6699;
assign w5126 = ~w13975 & ~w12658;
assign w5127 = w14983 & w15997;
assign w5128 = w15151 & w11134;
assign w5129 = ~w5879 & ~w12623;
assign w5130 = w952 & w3133;
assign w5131 = ~w15549 & ~w1440;
assign w5132 = a_4 & a_48;
assign w5133 = a_5 & a_34;
assign w5134 = ~w7259 & ~w13967;
assign w5135 = ~w18094 & ~w3804;
assign w5136 = w8029 & ~w19136;
assign w5137 = w420 & ~w3215;
assign w5138 = ~w3710 & ~w18509;
assign w5139 = ~w8127 & w18198;
assign w5140 = w13970 & ~w17301;
assign w5141 = w11932 & w9252;
assign w5142 = (~w724 & ~w7825) | (~w724 & w14650) | (~w7825 & w14650);
assign w5143 = ~w10308 & ~w13990;
assign w5144 = ~w13708 & ~w4369;
assign w5145 = ~w4179 & ~w9941;
assign w5146 = (~w5566 & w15771) | (~w5566 & w12016) | (w15771 & w12016);
assign w5147 = ~w7824 & ~w14089;
assign w5148 = ~w10199 & ~w13783;
assign w5149 = ~w1655 & ~w9147;
assign w5150 = ~w239 & ~w3684;
assign w5151 = ~w3144 & ~w17265;
assign w5152 = w17955 & w13096;
assign w5153 = ~w7751 & ~w12078;
assign w5154 = ~a_48 & a_49;
assign w5155 = ~w2799 & ~w5563;
assign w5156 = ~w4420 & ~w994;
assign w5157 = (w4528 & w17506) | (w4528 & w131) | (w17506 & w131);
assign w5158 = w10038 & ~w7513;
assign w5159 = ~w3468 & ~w2328;
assign w5160 = a_8 & a_32;
assign w5161 = a_9 & a_30;
assign w5162 = ~w9958 & ~w16484;
assign w5163 = ~w10277 & ~w13857;
assign w5164 = w1998 & w7537;
assign w5165 = a_4 & a_36;
assign w5166 = ~w10145 & ~w16657;
assign w5167 = w17671 & ~w15174;
assign w5168 = ~w12095 & w7360;
assign w5169 = ~w14056 & ~w2325;
assign w5170 = ~w1479 & ~w4954;
assign w5171 = ~w11607 & ~w13992;
assign w5172 = ~w306 & ~w15085;
assign w5173 = ~w4505 & ~w17299;
assign w5174 = w1594 & ~w15287;
assign w5175 = ~w6451 & ~w17709;
assign w5176 = a_20 & a_56;
assign w5177 = w15098 & ~w17717;
assign w5178 = w2616 & w2231;
assign w5179 = a_12 & a_54;
assign w5180 = (~w18423 & ~w11067) | (~w18423 & w15130) | (~w11067 & w15130);
assign w5181 = ~w4136 & ~w14558;
assign w5182 = ~w361 & ~w4648;
assign w5183 = ~w10572 & ~w18722;
assign w5184 = ~w13061 & w18798;
assign w5185 = w14441 & w16032;
assign w5186 = w17772 & w4507;
assign w5187 = ~w10850 & ~w11803;
assign w5188 = (w5640 & w4298) | (w5640 & w18445) | (w4298 & w18445);
assign w5189 = ~w1627 & ~w14845;
assign w5190 = ~w16956 & ~w11467;
assign w5191 = ~w13852 & ~w18087;
assign w5192 = ~w12952 & ~w7410;
assign w5193 = ~w16695 & ~w155;
assign w5194 = ~w14358 & ~w11769;
assign w5195 = ~w11615 & w14972;
assign w5196 = a_13 & a_50;
assign w5197 = w10456 & w5450;
assign w5198 = w316 & w677;
assign w5199 = a_11 & a_29;
assign w5200 = (~w6186 & ~w12232) | (~w6186 & w9136) | (~w12232 & w9136);
assign w5201 = ~w1404 & ~w16944;
assign w5202 = ~w2844 & w19197;
assign w5203 = ~w1905 & ~w18789;
assign w5204 = w850 & ~w13995;
assign w5205 = w8080 & ~w8836;
assign w5206 = ~w14895 & ~w3498;
assign w5207 = a_0 & a_8;
assign w5208 = ~w10584 & ~w11993;
assign w5209 = w2240 & ~w13070;
assign w5210 = ~w16071 & ~w11133;
assign w5211 = ~w3377 & ~w18600;
assign w5212 = a_32 & a_56;
assign w5213 = w14202 & w7997;
assign w5214 = a_14 & a_18;
assign w5215 = a_23 & a_28;
assign w5216 = ~w7374 & ~w2471;
assign w5217 = ~w9801 & ~w762;
assign w5218 = ~w2048 & w16288;
assign w5219 = ~w3728 & ~w18360;
assign w5220 = ~w14127 & w19065;
assign w5221 = w9983 & ~w11288;
assign w5222 = ~w9431 & ~w14002;
assign w5223 = ~w11982 & w1500;
assign w5224 = w11995 & ~w1893;
assign w5225 = ~w2203 & ~w16619;
assign w5226 = ~w16934 & ~w16580;
assign w5227 = ~w18761 & ~w16963;
assign w5228 = ~w3221 & w10830;
assign w5229 = ~w3125 & ~w11741;
assign w5230 = w1596 & w1320;
assign w5231 = ~w6365 & ~w10224;
assign w5232 = ~w2693 & ~w3681;
assign w5233 = ~w16826 & ~w7857;
assign w5234 = ~w9419 & ~w18577;
assign w5235 = w4279 & ~w5883;
assign w5236 = ~w8904 & w3689;
assign w5237 = ~w7732 & ~w2550;
assign w5238 = w13761 & ~w15088;
assign w5239 = a_6 & a_42;
assign w5240 = ~w3639 & ~w11916;
assign w5241 = ~w8113 & ~w12660;
assign w5242 = w18172 & ~w11814;
assign w5243 = w12406 & ~w2652;
assign w5244 = w16485 & w15266;
assign w5245 = w6481 & ~w2682;
assign w5246 = ~w8224 & ~w11186;
assign w5247 = a_43 & a_51;
assign w5248 = ~w18147 & w2933;
assign w5249 = a_12 & a_46;
assign w5250 = ~w17005 & ~w16029;
assign w5251 = ~w1329 & w17358;
assign w5252 = ~w14939 & ~w12959;
assign w5253 = w12295 & w4241;
assign w5254 = ~w10315 & ~w18103;
assign w5255 = ~w17307 & w4844;
assign w5256 = a_8 & a_14;
assign w5257 = ~w18159 & ~w11012;
assign w5258 = ~w6499 & w8003;
assign w5259 = a_16 & a_37;
assign w5260 = (~w13355 & ~w1766) | (~w13355 & w7532) | (~w1766 & w7532);
assign w5261 = ~w6515 & ~w7914;
assign w5262 = w5943 & ~w6994;
assign w5263 = w17544 & ~w18062;
assign w5264 = ~w2974 & ~w2767;
assign w5265 = w5884 & w5320;
assign w5266 = ~w15167 & ~w11920;
assign w5267 = ~w9740 & ~w11593;
assign w5268 = ~w11111 & ~w3142;
assign w5269 = ~w614 & ~w537;
assign w5270 = ~w7069 & ~w8865;
assign w5271 = ~w10601 & w9899;
assign w5272 = ~w12104 & w7597;
assign w5273 = a_50 & a_54;
assign w5274 = w4308 & ~w902;
assign w5275 = ~w13827 & w9198;
assign w5276 = ~w5023 & w13591;
assign w5277 = w18200 & w7435;
assign w5278 = ~w6021 & w7035;
assign w5279 = w10823 & w14472;
assign w5280 = a_44 & a_59;
assign w5281 = ~w3404 & ~w18642;
assign w5282 = ~w12688 & w12110;
assign w5283 = a_6 & a_13;
assign w5284 = ~w16196 & ~w13565;
assign w5285 = ~w4202 & ~w1073;
assign w5286 = w16859 & w17283;
assign w5287 = w3594 & ~w14558;
assign w5288 = ~w10967 & ~w11239;
assign w5289 = ~w13698 & ~w8484;
assign w5290 = ~w2374 & ~w12052;
assign w5291 = ~w1234 & ~w14159;
assign w5292 = ~w13154 & ~w235;
assign w5293 = ~w4308 & ~w4959;
assign w5294 = (~w2039 & ~w5761) | (~w2039 & w18022) | (~w5761 & w18022);
assign w5295 = ~w13736 & w7662;
assign w5296 = ~w372 & ~w2960;
assign w5297 = ~w16480 & w1916;
assign w5298 = ~w13372 & ~w15513;
assign w5299 = ~w8708 & ~w18634;
assign w5300 = ~w3827 & ~w13283;
assign w5301 = ~w10918 & ~w5908;
assign w5302 = (~w18674 & w17718) | (~w18674 & w15466) | (w17718 & w15466);
assign w5303 = ~w4997 & ~w4621;
assign w5304 = ~w7390 & ~w15425;
assign w5305 = ~w18702 & w14578;
assign w5306 = w4024 & ~w11242;
assign w5307 = ~w16646 & ~w7741;
assign w5308 = w5077 & w10069;
assign w5309 = ~w17829 & ~w12114;
assign w5310 = w13094 & ~w7333;
assign w5311 = ~w16647 & ~w3346;
assign w5312 = (~w16047 & ~w7737) | (~w16047 & w6627) | (~w7737 & w6627);
assign w5313 = a_24 & a_62;
assign w5314 = w18829 & ~w16304;
assign w5315 = ~w15064 & ~w211;
assign w5316 = (~w10136 & ~w6063) | (~w10136 & w16396) | (~w6063 & w16396);
assign w5317 = w1773 & ~w16830;
assign w5318 = ~w8419 & w4345;
assign w5319 = w4734 & ~w13137;
assign w5320 = ~w12039 & ~w12642;
assign w5321 = w1623 & ~w10048;
assign w5322 = ~w12630 & ~w780;
assign w5323 = ~w1730 & ~w3217;
assign w5324 = a_11 & a_47;
assign w5325 = ~w7606 & ~w16720;
assign w5326 = ~w4164 & w16424;
assign w5327 = ~w4760 & ~w13726;
assign w5328 = ~w4818 & ~w3272;
assign w5329 = ~w2961 & ~w9331;
assign w5330 = ~w11235 & ~w16883;
assign w5331 = w6943 & ~w15769;
assign w5332 = w13621 & ~w18629;
assign w5333 = (~w6971 & ~w14931) | (~w6971 & w13836) | (~w14931 & w13836);
assign w5334 = w11570 & ~w11364;
assign w5335 = ~w13546 & ~w16980;
assign w5336 = ~w4537 & w4715;
assign w5337 = a_31 & a_44;
assign w5338 = w10137 & ~w12253;
assign w5339 = a_15 & a_23;
assign w5340 = w13724 & ~w8509;
assign w5341 = (w7341 & w17539) | (w7341 & w5071) | (w17539 & w5071);
assign w5342 = ~w2152 & ~w17398;
assign w5343 = a_14 & a_23;
assign w5344 = ~w3028 & ~w16540;
assign w5345 = w11193 & ~w14589;
assign w5346 = w15579 & ~w9969;
assign w5347 = ~w3024 & w3222;
assign w5348 = ~w2667 & ~w14902;
assign w5349 = ~w11073 & ~w16306;
assign w5350 = ~w16506 & ~w9887;
assign w5351 = a_16 & a_42;
assign w5352 = ~w4624 & ~w6897;
assign w5353 = ~w18578 & w11794;
assign w5354 = ~w8853 & ~w4916;
assign w5355 = ~w8098 & w19156;
assign w5356 = ~w18145 & ~w4760;
assign w5357 = ~w508 & w17308;
assign w5358 = ~w17976 & ~w18649;
assign w5359 = a_1 & a_5;
assign w5360 = ~w10720 & w1288;
assign w5361 = w12600 & w5141;
assign w5362 = w18904 & ~w4372;
assign w5363 = ~w10851 & w12512;
assign w5364 = ~w16028 & w7575;
assign w5365 = (~w1037 & ~w18702) | (~w1037 & w5687) | (~w18702 & w5687);
assign w5366 = w18067 & ~w14522;
assign w5367 = ~w14612 & ~w7799;
assign w5368 = ~w13291 & w4173;
assign w5369 = ~w15098 & w17717;
assign w5370 = w13059 & ~w8530;
assign w5371 = ~w6535 & w2862;
assign w5372 = w4428 & w10641;
assign w5373 = w14153 & w9495;
assign w5374 = ~w10201 & ~w13331;
assign w5375 = ~w13182 & ~w4446;
assign w5376 = ~w10598 & ~w9588;
assign w5377 = ~w13384 & ~w16400;
assign w5378 = a_24 & a_44;
assign w5379 = ~w15488 & ~w13814;
assign w5380 = ~w18169 & ~w9222;
assign w5381 = a_27 & a_46;
assign w5382 = a_27 & a_30;
assign w5383 = w6441 & ~w926;
assign w5384 = a_15 & a_36;
assign w5385 = w3236 & w14868;
assign w5386 = w7548 & ~w13199;
assign w5387 = a_14 & a_25;
assign w5388 = ~w17369 & w12848;
assign w5389 = w4605 | w4394;
assign w5390 = w11905 & w2264;
assign w5391 = ~w3224 & ~w11989;
assign w5392 = ~w5770 & w11595;
assign w5393 = a_25 & a_28;
assign w5394 = ~w17843 & ~w11426;
assign w5395 = a_28 & a_63;
assign w5396 = ~w11505 & ~w17602;
assign w5397 = ~w14229 & ~w13362;
assign w5398 = w15134 & ~w17889;
assign w5399 = w3491 & ~w8015;
assign w5400 = ~w12910 & ~w3181;
assign w5401 = ~w18660 & ~w5039;
assign w5402 = ~w13064 & ~w7523;
assign w5403 = ~w6500 & ~w2668;
assign w5404 = ~w14035 & ~w4682;
assign w5405 = (w8699 & w2769) | (w8699 & w663) | (w2769 & w663);
assign w5406 = ~w18564 & ~w14320;
assign w5407 = (w7969 & w13082) | (w7969 & w13733) | (w13082 & w13733);
assign w5408 = w14910 & ~w1791;
assign w5409 = (w14650 & w5142) | (w14650 & ~w19001) | (w5142 & ~w19001);
assign w5410 = (~w1391 & w5527) | (~w1391 & w15027) | (w5527 & w15027);
assign w5411 = ~w15883 & ~w5876;
assign w5412 = a_4 & a_13;
assign w5413 = ~w2304 & ~w17769;
assign w5414 = ~w9898 & ~w6137;
assign w5415 = (~w8158 & ~w6513) | (~w8158 & w4384) | (~w6513 & w4384);
assign w5416 = ~w18471 & ~w16719;
assign w5417 = ~w9115 & w1896;
assign w5418 = (~w4559 & w17531) | (~w4559 & w17716) | (w17531 & w17716);
assign w5419 = ~w1957 & ~w2467;
assign w5420 = w6002 & ~w4451;
assign w5421 = w10635 & w2573;
assign w5422 = ~w13794 & ~w5045;
assign w5423 = a_32 & a_48;
assign w5424 = a_31 & a_33;
assign w5425 = ~w10670 & ~w13876;
assign w5426 = ~w18891 & ~w10801;
assign w5427 = w8288 & ~w8727;
assign w5428 = ~w357 & w876;
assign w5429 = ~w5963 & ~w14343;
assign w5430 = ~w6571 & w948;
assign w5431 = ~w16886 & ~w9043;
assign w5432 = ~w4372 & ~w17295;
assign w5433 = (w13603 & w17529) | (w13603 & w13081) | (w17529 & w13081);
assign w5434 = ~w3875 & ~w344;
assign w5435 = ~w9746 & ~w8858;
assign w5436 = a_44 & a_54;
assign w5437 = ~w16260 & w6747;
assign w5438 = ~w16073 & ~w4058;
assign w5439 = ~w5172 & ~w7810;
assign w5440 = ~w1085 & w4925;
assign w5441 = (~w12463 & ~w2713) | (~w12463 & w16010) | (~w2713 & w16010);
assign w5442 = a_7 & a_19;
assign w5443 = w17413 & ~w10500;
assign w5444 = ~w13515 & ~w7109;
assign w5445 = ~w11660 & ~w12206;
assign w5446 = w16587 & w12503;
assign w5447 = ~w11459 & ~w13152;
assign w5448 = w596 & w18537;
assign w5449 = w17337 & ~w4024;
assign w5450 = a_18 & a_41;
assign w5451 = w9629 & ~w15032;
assign w5452 = ~w6371 & ~w17230;
assign w5453 = ~w12794 & ~w10280;
assign w5454 = ~w15861 & w8481;
assign w5455 = ~w13774 & ~w6898;
assign w5456 = w15010 & ~w9562;
assign w5457 = ~w12300 & ~w12923;
assign w5458 = ~w2935 & ~w11209;
assign w5459 = a_50 & a_55;
assign w5460 = w4137 & w19157;
assign w5461 = w6326 & w17212;
assign w5462 = a_17 & a_45;
assign w5463 = (~w7126 & ~w15089) | (~w7126 & w4796) | (~w15089 & w4796);
assign w5464 = (~w2433 & w11390) | (~w2433 & w6721) | (w11390 & w6721);
assign w5465 = ~w13074 & ~w1485;
assign w5466 = w16283 & ~w7559;
assign w5467 = ~w15921 & w5871;
assign w5468 = a_2 & a_9;
assign w5469 = ~w3569 & ~w4062;
assign w5470 = (~w17101 & w4082) | (~w17101 & w13381) | (w4082 & w13381);
assign w5471 = ~w17040 & ~w3532;
assign w5472 = ~w10057 & w10400;
assign w5473 = ~w4649 & ~w8776;
assign w5474 = w9396 | w840;
assign w5475 = (~w4340 & ~w12015) | (~w4340 & w4736) | (~w12015 & w4736);
assign w5476 = ~w2644 & ~w11661;
assign w5477 = w11273 & ~w8594;
assign w5478 = a_14 & a_30;
assign w5479 = ~w2076 & ~w17135;
assign w5480 = w17173 & w12625;
assign w5481 = w9634 & ~w4041;
assign w5482 = a_5 & a_15;
assign w5483 = w4549 & ~w18566;
assign w5484 = ~w8711 & ~w12289;
assign w5485 = ~w18397 & w14169;
assign w5486 = (w17797 & w2769) | (w17797 & w3916) | (w2769 & w3916);
assign w5487 = ~w10907 & ~w1608;
assign w5488 = ~w11983 & ~w2419;
assign w5489 = w18548 & ~w10992;
assign w5490 = ~w5095 & w12441;
assign w5491 = a_7 & a_61;
assign w5492 = ~w1198 & ~w2340;
assign w5493 = a_42 & a_58;
assign w5494 = a_16 & a_57;
assign w5495 = (w15103 & w15988) | (w15103 & w1982) | (w15988 & w1982);
assign w5496 = ~w14340 & ~w15973;
assign w5497 = w8806 & ~w7185;
assign w5498 = ~w2672 & ~w16075;
assign w5499 = ~w10387 & ~w5941;
assign w5500 = (w9337 & w16205) | (w9337 & w3281) | (w16205 & w3281);
assign w5501 = w7844 & ~w14607;
assign w5502 = ~w1690 & ~w14588;
assign w5503 = w8125 & w9227;
assign w5504 = ~w15567 & ~w12115;
assign w5505 = w6655 & ~w466;
assign w5506 = w3459 & ~w17694;
assign w5507 = a_6 & a_54;
assign w5508 = w5183 & ~w17584;
assign w5509 = ~w5426 & ~w17133;
assign w5510 = w18627 & w9166;
assign w5511 = a_34 & a_56;
assign w5512 = ~w14405 & ~w7558;
assign w5513 = ~w16076 & ~w10085;
assign w5514 = w14895 & w3498;
assign w5515 = w5513 & ~w3254;
assign w5516 = ~w6751 & ~w5130;
assign w5517 = w5415 & ~w3745;
assign w5518 = ~w8974 & w5781;
assign w5519 = a_47 & a_58;
assign w5520 = (~w17197 & w691) | (~w17197 & w3462) | (w691 & w3462);
assign w5521 = w6363 & ~w4681;
assign w5522 = w10083 & ~w9955;
assign w5523 = ~w928 & ~w16922;
assign w5524 = ~w228 & ~w16441;
assign w5525 = a_7 & a_58;
assign w5526 = ~w396 & w15299;
assign w5527 = (w16025 & w9221) | (w16025 & w6432) | (w9221 & w6432);
assign w5528 = ~w4700 & w10595;
assign w5529 = ~w7303 & w14604;
assign w5530 = a_28 & a_56;
assign w5531 = ~w8946 & w4604;
assign w5532 = a_15 & a_40;
assign w5533 = w16344 & w5774;
assign w5534 = w13553 & w18503;
assign w5535 = ~w8700 & w1990;
assign w5536 = w1654 & ~w14579;
assign w5537 = ~w1489 & w9947;
assign w5538 = w3810 & ~w10684;
assign w5539 = w10538 & ~w6938;
assign w5540 = w17496 & ~w1920;
assign w5541 = (~w16969 & ~w12423) | (~w16969 & w17343) | (~w12423 & w17343);
assign w5542 = (w17294 & w2026) | (w17294 & w9266) | (w2026 & w9266);
assign w5543 = w14069 & ~w16515;
assign w5544 = a_2 & a_52;
assign w5545 = a_52 & a_58;
assign w5546 = ~w14118 & ~w13112;
assign w5547 = ~w16691 & ~w14761;
assign w5548 = ~w7639 & w8292;
assign w5549 = ~w7658 & ~w13623;
assign w5550 = w16206 & ~w6115;
assign w5551 = a_22 & a_42;
assign w5552 = w9372 & ~w6917;
assign w5553 = w18182 & ~w2358;
assign w5554 = a_4 & a_18;
assign w5555 = w7273 & ~w13500;
assign w5556 = ~w18169 & ~w13183;
assign w5557 = ~w15507 & ~w10867;
assign w5558 = a_16 & a_46;
assign w5559 = w11597 & ~w15652;
assign w5560 = ~w16713 & ~w13892;
assign w5561 = ~w8262 & ~w3906;
assign w5562 = ~w2644 & ~w5889;
assign w5563 = w5735 & w15228;
assign w5564 = ~w9608 & ~w10633;
assign w5565 = ~w3363 & ~w12524;
assign w5566 = ~w1209 & ~w12498;
assign w5567 = ~w6782 & ~w7427;
assign w5568 = ~w11131 & ~w4359;
assign w5569 = ~w5077 & ~w10069;
assign w5570 = w19070 & ~w9867;
assign w5571 = a_24 & a_53;
assign w5572 = ~w11079 & ~w16339;
assign w5573 = w7703 & w13655;
assign w5574 = a_11 & a_17;
assign w5575 = ~w15882 & w12142;
assign w5576 = ~w2923 & w8351;
assign w5577 = ~w11409 & ~w7602;
assign w5578 = ~w16913 & ~w9030;
assign w5579 = w6610 & w8550;
assign w5580 = w18750 & w1071;
assign w5581 = ~w2228 & w1243;
assign w5582 = w8905 & w1305;
assign w5583 = ~w14100 & ~w10188;
assign w5584 = w13155 & ~w2770;
assign w5585 = ~w5744 & ~w9087;
assign w5586 = ~w7931 & ~w2082;
assign w5587 = ~w9026 & ~w14999;
assign w5588 = ~w2532 & ~w18140;
assign w5589 = ~w16163 & w3783;
assign w5590 = ~w528 & ~w17913;
assign w5591 = ~w16370 & ~w5555;
assign w5592 = ~w680 & ~w8280;
assign w5593 = ~w12356 & ~w3223;
assign w5594 = ~w15452 & ~w1398;
assign w5595 = ~w4186 & ~w5840;
assign w5596 = ~w3083 & ~w3383;
assign w5597 = w4474 & w3841;
assign w5598 = ~w5002 & ~w5916;
assign w5599 = ~w4198 & ~w9464;
assign w5600 = ~w17304 & ~w13419;
assign w5601 = ~w6853 & w6052;
assign w5602 = (~w5967 & w15904) | (~w5967 & w2565) | (w15904 & w2565);
assign w5603 = ~w15139 & ~w17552;
assign w5604 = ~w13571 & ~w14818;
assign w5605 = w15701 & ~w11319;
assign w5606 = ~w16450 & ~w17738;
assign w5607 = ~w13960 & ~w7300;
assign w5608 = ~w4706 & ~w9344;
assign w5609 = w16562 & ~w5426;
assign w5610 = ~w17604 & ~w7969;
assign w5611 = w18109 & ~w4589;
assign w5612 = w92 & w6070;
assign w5613 = ~w5456 & ~w18174;
assign w5614 = a_25 & a_50;
assign w5615 = w1887 & ~w5150;
assign w5616 = ~w11455 & w8459;
assign w5617 = ~w18603 & ~w338;
assign w5618 = ~w10330 & w1295;
assign w5619 = w7756 & ~w2700;
assign w5620 = w18893 & w1537;
assign w5621 = a_18 & a_28;
assign w5622 = a_8 & a_63;
assign w5623 = ~w5844 & ~w809;
assign w5624 = ~w11939 & w7921;
assign w5625 = ~w2307 & w15165;
assign w5626 = ~w10321 & ~w10219;
assign w5627 = w2295 & w18731;
assign w5628 = ~w3494 & ~w9147;
assign w5629 = ~w10286 & ~w9353;
assign w5630 = ~a_44 & a_45;
assign w5631 = ~w15154 & ~w10168;
assign w5632 = ~w14792 & w7136;
assign w5633 = w4265 & ~w5767;
assign w5634 = a_14 & a_37;
assign w5635 = w458 & ~w15965;
assign w5636 = ~w15511 & w15378;
assign w5637 = w3390 & ~w3749;
assign w5638 = ~w12612 & w16380;
assign w5639 = ~w13210 & w13992;
assign w5640 = ~w15813 & ~w9918;
assign w5641 = ~w13903 & ~w17152;
assign w5642 = ~w14434 & ~w17966;
assign w5643 = w15151 & ~w16388;
assign w5644 = ~w13276 & ~w7783;
assign w5645 = ~w12170 & w4172;
assign w5646 = ~w6615 & ~w18628;
assign w5647 = ~w15660 & ~w14061;
assign w5648 = ~w10050 & ~w14609;
assign w5649 = ~w4491 & w16152;
assign w5650 = ~w4880 & ~w6947;
assign w5651 = w4453 & ~w13905;
assign w5652 = ~w5199 & ~w7183;
assign w5653 = w4545 & ~w16641;
assign w5654 = a_15 & a_62;
assign w5655 = ~w6966 & ~w7234;
assign w5656 = a_7 & a_28;
assign w5657 = w10397 | w13037;
assign w5658 = ~w11797 & ~w17341;
assign w5659 = w10596 & w8385;
assign w5660 = (~w3604 & ~w9045) | (~w3604 & w10463) | (~w9045 & w10463);
assign w5661 = ~w9864 & ~w13784;
assign w5662 = ~w5932 & w2525;
assign w5663 = w12302 & w5003;
assign w5664 = ~w1013 & ~w3017;
assign w5665 = ~w13804 & w3558;
assign w5666 = ~w1706 & w15122;
assign w5667 = a_5 & a_48;
assign w5668 = w5415 & ~w18222;
assign w5669 = ~w14810 & ~w15580;
assign w5670 = ~w3547 & ~w3883;
assign w5671 = w16362 & ~w5857;
assign w5672 = ~w7572 & ~w4256;
assign w5673 = (~w12288 & w10330) | (~w12288 & w10923) | (w10330 & w10923);
assign w5674 = w815 & ~w8757;
assign w5675 = w6426 & w11523;
assign w5676 = (w18187 & ~w14095) | (w18187 & w17952) | (~w14095 & w17952);
assign w5677 = ~w12906 & ~w11311;
assign w5678 = w18640 & w10970;
assign w5679 = ~w3210 & ~w2777;
assign w5680 = ~w8946 & ~w12711;
assign w5681 = ~w18887 & ~w13102;
assign w5682 = ~w18934 & ~w19120;
assign w5683 = (~w569 & ~w13158) | (~w569 & w8027) | (~w13158 & w8027);
assign w5684 = (~w4195 & w12278) | (~w4195 & w18856) | (w12278 & w18856);
assign w5685 = ~w15244 & ~w12474;
assign w5686 = a_24 & a_25;
assign w5687 = w14578 & ~w1037;
assign w5688 = ~w12234 & ~w12984;
assign w5689 = ~w4320 & w6468;
assign w5690 = ~w8134 & w6113;
assign w5691 = w3514 & ~w18630;
assign w5692 = ~w11971 & ~w14639;
assign w5693 = w13353 & w9721;
assign w5694 = ~w13301 & ~w12815;
assign w5695 = ~w3384 & ~w18367;
assign w5696 = a_16 & a_22;
assign w5697 = a_39 & a_45;
assign w5698 = ~w16308 & ~w13563;
assign w5699 = ~w2376 & ~w15241;
assign w5700 = w1329 & ~w17358;
assign w5701 = w17773 & ~w16895;
assign w5702 = ~w15276 & w12216;
assign w5703 = ~w10823 & ~w14472;
assign w5704 = ~w10269 & w5096;
assign w5705 = ~w14893 & ~w17700;
assign w5706 = w8240 & w1566;
assign w5707 = ~w11923 & ~w17864;
assign w5708 = ~w12529 & w8328;
assign w5709 = w2465 & ~w10669;
assign w5710 = w7074 & w15753;
assign w5711 = ~w4281 & ~w13896;
assign w5712 = ~w9477 & ~w6036;
assign w5713 = (w4471 & w3219) | (w4471 & w18708) | (w3219 & w18708);
assign w5714 = ~w13968 & ~w14543;
assign w5715 = a_6 & a_30;
assign w5716 = w1353 & ~w16614;
assign w5717 = ~w14742 & w1368;
assign w5718 = w7926 & ~w17201;
assign w5719 = w10861 & ~w10412;
assign w5720 = ~w1559 & ~w17910;
assign w5721 = w13161 & ~w16908;
assign w5722 = w5093 & w16498;
assign w5723 = ~w1402 & ~w2085;
assign w5724 = ~w18907 & ~w18967;
assign w5725 = (~w16012 & ~w341) | (~w16012 & w12425) | (~w341 & w12425);
assign w5726 = ~w7841 & ~w15816;
assign w5727 = a_4 & a_24;
assign w5728 = ~w16638 & ~w16063;
assign w5729 = w1962 & w7592;
assign w5730 = ~w8917 & w9684;
assign w5731 = ~w5754 & w8215;
assign w5732 = w8233 & ~w14262;
assign w5733 = ~w7872 & ~w2099;
assign w5734 = w8791 & w1015;
assign w5735 = a_29 & a_30;
assign w5736 = w7786 & ~w846;
assign w5737 = a_0 & a_25;
assign w5738 = a_29 & a_52;
assign w5739 = ~w13567 & ~w12361;
assign w5740 = w15415 & w7294;
assign w5741 = ~w1196 & ~w4479;
assign w5742 = ~w6097 & ~w2711;
assign w5743 = w17914 & w12178;
assign w5744 = w8799 & ~w5792;
assign w5745 = ~w7019 & ~w2206;
assign w5746 = (~w17033 & ~w15401) | (~w17033 & w12223) | (~w15401 & w12223);
assign w5747 = ~w9328 & w5556;
assign w5748 = w14294 & ~w11609;
assign w5749 = w1363 & ~w16428;
assign w5750 = ~w4820 & ~w7006;
assign w5751 = ~w5416 & ~w1949;
assign w5752 = ~w12823 & ~w18877;
assign w5753 = ~w3208 & w2300;
assign w5754 = ~w10462 & ~w17853;
assign w5755 = w2 & ~w17707;
assign w5756 = ~w10677 & ~w1717;
assign w5757 = w17419 & w10719;
assign w5758 = ~w9204 & ~w17939;
assign w5759 = a_31 & a_50;
assign w5760 = a_5 & a_30;
assign w5761 = ~w2039 & ~w77;
assign w5762 = w4549 & ~w11940;
assign w5763 = ~w8165 & ~w9400;
assign w5764 = ~w15942 & ~w8835;
assign w5765 = (~w18576 & ~w6096) | (~w18576 & w18712) | (~w6096 & w18712);
assign w5766 = w14435 & ~w5163;
assign w5767 = ~w3441 & ~w549;
assign w5768 = ~w11970 & ~w15435;
assign w5769 = ~w14042 & ~w9352;
assign w5770 = w15970 & ~w11737;
assign w5771 = (~w13342 & ~w17491) | (~w13342 & w12462) | (~w17491 & w12462);
assign w5772 = ~w6528 & ~w11398;
assign w5773 = ~w7517 & ~w6163;
assign w5774 = ~w15073 & ~w17166;
assign w5775 = (~w17277 & ~w9896) | (~w17277 & w5785) | (~w9896 & w5785);
assign w5776 = ~w2025 & w18505;
assign w5777 = ~w13761 & w15088;
assign w5778 = ~w18375 & w388;
assign w5779 = w1655 & ~w5628;
assign w5780 = ~w4676 & ~w542;
assign w5781 = ~w10811 & ~w4209;
assign w5782 = w6228 & ~w1276;
assign w5783 = (~w9077 & w14792) | (~w9077 & w11805) | (w14792 & w11805);
assign w5784 = a_35 & a_60;
assign w5785 = w13473 & ~w17277;
assign w5786 = ~w14944 & w12072;
assign w5787 = ~w3873 & ~w3753;
assign w5788 = (w15832 & w14223) | (w15832 & w2027) | (w14223 & w2027);
assign w5789 = w15897 & w2324;
assign w5790 = ~w15752 & ~w10461;
assign w5791 = ~w6948 & w2396;
assign w5792 = ~w13933 & ~w8796;
assign w5793 = a_54 & a_57;
assign w5794 = w14167 & ~w11486;
assign w5795 = ~w6673 & ~w5181;
assign w5796 = ~w3771 & ~w9811;
assign w5797 = a_44 & a_60;
assign w5798 = w12667 & ~w15987;
assign w5799 = w948 & ~w17322;
assign w5800 = ~w16357 & ~w16378;
assign w5801 = ~w19055 & w4126;
assign w5802 = w16211 & ~w11419;
assign w5803 = w11577 & ~w6391;
assign w5804 = w18234 & ~w16670;
assign w5805 = ~w18407 & ~w11208;
assign w5806 = a_10 & a_54;
assign w5807 = w13151 & ~w9309;
assign w5808 = ~w15461 & ~w4077;
assign w5809 = ~w11215 & ~w4689;
assign w5810 = ~w10177 & ~w12116;
assign w5811 = ~w16605 & ~w12177;
assign w5812 = ~w13433 & ~w8394;
assign w5813 = w11822 & ~w16728;
assign w5814 = (~w10266 & w11644) | (~w10266 & w16715) | (w11644 & w16715);
assign w5815 = w14915 & ~w4834;
assign w5816 = a_43 & a_54;
assign w5817 = ~w10018 & ~w18684;
assign w5818 = ~w17945 & ~w9305;
assign w5819 = w15663 & w7756;
assign w5820 = ~w13343 & ~w13413;
assign w5821 = ~w4888 & ~w3520;
assign w5822 = ~w301 & ~w14459;
assign w5823 = w16427 & ~w9471;
assign w5824 = ~w17528 & ~w13541;
assign w5825 = (~w16966 & ~w12559) | (~w16966 & w14799) | (~w12559 & w14799);
assign w5826 = ~w6853 & w5673;
assign w5827 = ~w3433 & ~w3292;
assign w5828 = ~w7717 & ~w13506;
assign w5829 = ~w13398 & ~w15944;
assign w5830 = ~w12459 & ~w18782;
assign w5831 = w6974 & ~w3714;
assign w5832 = ~w12981 & ~w12367;
assign w5833 = w6409 & ~w8183;
assign w5834 = w8080 & ~w8122;
assign w5835 = ~w16807 & w16234;
assign w5836 = (~w12791 & ~w6503) | (~w12791 & w18569) | (~w6503 & w18569);
assign w5837 = ~w16822 & ~w5548;
assign w5838 = w3606 & ~w4365;
assign w5839 = ~w7551 & ~w968;
assign w5840 = w17068 & ~w11029;
assign w5841 = ~w15562 & w6769;
assign w5842 = a_1 & a_53;
assign w5843 = ~w7529 & w17948;
assign w5844 = ~w16731 & ~w5038;
assign w5845 = ~w12324 & ~w15121;
assign w5846 = w1237 & ~w56;
assign w5847 = a_4 & a_21;
assign w5848 = ~w6600 & ~w14750;
assign w5849 = ~w8887 & ~w8097;
assign w5850 = ~w12846 & w2248;
assign w5851 = ~w3084 & ~w16000;
assign w5852 = ~w3953 & ~w11236;
assign w5853 = w3930 & ~w2161;
assign w5854 = w8918 & ~w5084;
assign w5855 = (~w9760 & w5495) | (~w9760 & w15926) | (w5495 & w15926);
assign w5856 = w7248 & w16034;
assign w5857 = ~w604 & ~w7238;
assign w5858 = ~w8504 & w10599;
assign w5859 = a_13 & a_15;
assign w5860 = ~w6158 & w3911;
assign w5861 = ~w676 & w18563;
assign w5862 = w6951 & ~w15637;
assign w5863 = ~w1951 & ~w16011;
assign w5864 = ~w4060 & ~w13047;
assign w5865 = a_15 & a_55;
assign w5866 = ~w12904 & ~w10231;
assign w5867 = a_1 & a_28;
assign w5868 = a_43 & a_50;
assign w5869 = (~w7768 & w585) | (~w7768 & w647) | (w585 & w647);
assign w5870 = a_0 & a_48;
assign w5871 = a_20 & a_60;
assign w5872 = a_46 & a_53;
assign w5873 = ~w6738 & ~w19104;
assign w5874 = (~w7675 & ~w6912) | (~w7675 & w462) | (~w6912 & w462);
assign w5875 = a_3 & a_8;
assign w5876 = ~w5803 & ~w8521;
assign w5877 = a_19 & a_56;
assign w5878 = ~w7148 & w2780;
assign w5879 = ~w17803 & ~w1770;
assign w5880 = ~w6655 & w466;
assign w5881 = ~w6494 & ~w3855;
assign w5882 = (w11659 & w553) | (w11659 & w18546) | (w553 & w18546);
assign w5883 = ~w6937 & ~w16219;
assign w5884 = w14217 & ~w3328;
assign w5885 = ~w7206 & ~w7088;
assign w5886 = ~w5987 & ~w12311;
assign w5887 = ~w3594 & w14558;
assign w5888 = w9258 & ~w4753;
assign w5889 = ~w15035 & ~w6320;
assign w5890 = a_36 & w9421;
assign w5891 = ~w18647 & ~w15232;
assign w5892 = w4833 & ~w6929;
assign w5893 = (a_52 & w10851) | (a_52 & w7956) | (w10851 & w7956);
assign w5894 = (~w9696 & ~w4184) | (~w9696 & w18482) | (~w4184 & w18482);
assign w5895 = a_5 & a_12;
assign w5896 = ~w15918 & w17169;
assign w5897 = ~w8920 & ~w18058;
assign w5898 = ~w10223 & ~w5806;
assign w5899 = ~w2847 & w572;
assign w5900 = w6541 & ~w1132;
assign w5901 = ~w1259 & ~w3436;
assign w5902 = a_32 & a_52;
assign w5903 = ~w18295 & ~w10643;
assign w5904 = w1621 & ~w2663;
assign w5905 = ~w14833 & ~w10126;
assign w5906 = ~w11717 & ~w10422;
assign w5907 = a_14 & a_17;
assign w5908 = ~w8160 & w5001;
assign w5909 = ~w5660 & ~w15408;
assign w5910 = ~w1109 & w12679;
assign w5911 = w9254 & w11558;
assign w5912 = ~w15047 & w1266;
assign w5913 = ~w15753 & w9114;
assign w5914 = a_1 & a_38;
assign w5915 = a_6 & a_51;
assign w5916 = w15577 & ~w12250;
assign w5917 = a_36 & a_41;
assign w5918 = w5622 & w13333;
assign w5919 = a_7 & a_41;
assign w5920 = ~w2937 & w7159;
assign w5921 = ~w4683 & ~w3979;
assign w5922 = ~w2653 & ~w16257;
assign w5923 = w14372 & w2662;
assign w5924 = w12232 & w10474;
assign w5925 = ~w8603 & ~w6654;
assign w5926 = ~w13206 & ~w2907;
assign w5927 = w2847 & ~w572;
assign w5928 = ~w7029 & ~w9781;
assign w5929 = (~w537 & ~w19114) | (~w537 & w5269) | (~w19114 & w5269);
assign w5930 = ~w16207 & ~w3370;
assign w5931 = w17573 & ~w7978;
assign w5932 = ~w18806 & ~w3596;
assign w5933 = ~w18093 & w1898;
assign w5934 = ~w14903 & ~w4162;
assign w5935 = ~w3763 & ~w8150;
assign w5936 = ~w17956 & w4139;
assign w5937 = w10058 & w10947;
assign w5938 = ~w578 & ~w16422;
assign w5939 = ~w18975 & w1225;
assign w5940 = ~w11194 & w14931;
assign w5941 = ~w16280 & ~w5870;
assign w5942 = w6433 & w16371;
assign w5943 = a_27 & a_54;
assign w5944 = (~w8901 & ~w7464) | (~w8901 & w14529) | (~w7464 & w14529);
assign w5945 = a_43 & a_52;
assign w5946 = w493 & ~w8937;
assign w5947 = w13021 & ~w17368;
assign w5948 = ~w8964 & ~w11903;
assign w5949 = ~w4642 & ~w13938;
assign w5950 = a_2 & a_54;
assign w5951 = a_59 & a_61;
assign w5952 = ~w9842 & ~w8985;
assign w5953 = ~w4924 & ~w908;
assign w5954 = w4895 & w4842;
assign w5955 = ~w17115 & w2001;
assign w5956 = ~w17341 & ~w9112;
assign w5957 = w8414 & ~w16341;
assign w5958 = ~w18429 & ~w16099;
assign w5959 = ~w15294 & ~w6013;
assign w5960 = w15728 & ~w608;
assign w5961 = ~w9807 & w14449;
assign w5962 = w582 & ~w4322;
assign w5963 = ~w310 & w688;
assign w5964 = a_60 & a_61;
assign w5965 = w1710 & w4806;
assign w5966 = ~w565 & w7461;
assign w5967 = ~w4488 & ~w1216;
assign w5968 = w675 & w799;
assign w5969 = ~w10231 & w9695;
assign w5970 = ~w776 & ~w2387;
assign w5971 = ~w19035 & w7604;
assign w5972 = ~w15808 & w11057;
assign w5973 = w3998 & w5447;
assign w5974 = ~w6926 & ~w14790;
assign w5975 = w5289 & ~w16688;
assign w5976 = ~w1859 & ~w1315;
assign w5977 = ~w7030 & ~w14096;
assign w5978 = w2977 & ~w14959;
assign w5979 = ~w16061 & ~w7024;
assign w5980 = w9405 & ~w12840;
assign w5981 = ~w8228 & ~w12389;
assign w5982 = ~w12154 & ~w10478;
assign w5983 = ~w1706 & ~w17281;
assign w5984 = w13495 & w17565;
assign w5985 = ~w17450 & ~w18257;
assign w5986 = ~a_9 & ~w13123;
assign w5987 = w17794 & w1676;
assign w5988 = ~w2436 & ~w14565;
assign w5989 = ~w16706 & ~w5197;
assign w5990 = ~w6212 & ~w7381;
assign w5991 = ~w13459 & w687;
assign w5992 = w5261 & ~w18913;
assign w5993 = a_30 & a_54;
assign w5994 = ~w14428 & w17226;
assign w5995 = ~w2075 & w740;
assign w5996 = ~w18924 & ~w12880;
assign w5997 = ~w17815 & ~w14733;
assign w5998 = ~w4633 & w3522;
assign w5999 = ~w11331 & ~w5707;
assign w6000 = a_27 & a_56;
assign w6001 = ~w2514 & ~w13917;
assign w6002 = ~w6069 & ~w2326;
assign w6003 = a_4 & a_6;
assign w6004 = ~w16371 & ~w14005;
assign w6005 = w11504 & ~w17445;
assign w6006 = ~w5408 & ~w4773;
assign w6007 = w14218 & ~w5069;
assign w6008 = ~w2391 & ~w3510;
assign w6009 = a_6 & a_40;
assign w6010 = ~w9474 & w7186;
assign w6011 = ~w18118 & ~w2855;
assign w6012 = ~w2093 & w13241;
assign w6013 = ~w10626 & ~w10696;
assign w6014 = (w1320 & w487) | (w1320 & w1726) | (w487 & w1726);
assign w6015 = w245 & ~w367;
assign w6016 = ~w16369 & ~w3545;
assign w6017 = a_5 & a_61;
assign w6018 = ~w403 & w19158;
assign w6019 = ~w12935 & w16093;
assign w6020 = ~w13537 & ~w15586;
assign w6021 = ~w8913 & ~w10088;
assign w6022 = w12782 & ~w19035;
assign w6023 = ~w2769 & w7188;
assign w6024 = w14636 & ~w6823;
assign w6025 = w4105 & ~w4546;
assign w6026 = ~w13399 & ~w10545;
assign w6027 = a_24 & a_33;
assign w6028 = w10350 & ~w1373;
assign w6029 = a_33 & a_52;
assign w6030 = a_0 & a_21;
assign w6031 = ~w2272 & ~w6918;
assign w6032 = w2533 & ~w3863;
assign w6033 = ~w14085 & w5663;
assign w6034 = ~w16817 & ~w2137;
assign w6035 = w13249 & w12085;
assign w6036 = w13504 & w12790;
assign w6037 = ~w2810 & ~w6687;
assign w6038 = w12326 & ~w13551;
assign w6039 = ~w13820 & ~w5790;
assign w6040 = ~w7807 & ~w7768;
assign w6041 = ~w2606 & ~w15484;
assign w6042 = w12810 & ~w13983;
assign w6043 = a_5 & a_58;
assign w6044 = (w9957 & w14332) | (w9957 & w13688) | (w14332 & w13688);
assign w6045 = w17028 & w9700;
assign w6046 = ~w7691 & ~w2988;
assign w6047 = w2979 & w16111;
assign w6048 = w5214 & ~w14259;
assign w6049 = ~w9410 & ~w19083;
assign w6050 = ~w8793 & ~w2940;
assign w6051 = ~w2107 & ~w9276;
assign w6052 = (~w847 & w10330) | (~w847 & w1150) | (w10330 & w1150);
assign w6053 = ~w15996 & ~w9070;
assign w6054 = ~w15767 & ~w11809;
assign w6055 = ~w8417 & ~w17430;
assign w6056 = ~w7862 & ~w4740;
assign w6057 = ~w7698 & ~w14345;
assign w6058 = ~w2079 & ~w6099;
assign w6059 = ~w2918 & ~w1340;
assign w6060 = a_13 & a_40;
assign w6061 = (~w11406 & w9395) | (~w11406 & w17540) | (w9395 & w17540);
assign w6062 = ~w15068 & ~w11196;
assign w6063 = ~w3022 & ~w10136;
assign w6064 = a_8 & a_58;
assign w6065 = ~w9012 & ~w14368;
assign w6066 = ~w19125 & ~w16780;
assign w6067 = w15235 & w7767;
assign w6068 = ~w7392 & ~w15719;
assign w6069 = ~w18246 & ~w11289;
assign w6070 = ~w12308 & ~w5155;
assign w6071 = ~a_57 & a_58;
assign w6072 = ~w7061 & ~w3752;
assign w6073 = w2270 & ~w1879;
assign w6074 = (w1540 & w12258) | (w1540 & ~w5108) | (w12258 & ~w5108);
assign w6075 = ~w4135 & ~w8;
assign w6076 = ~w7305 & ~w16916;
assign w6077 = ~w7401 & w17942;
assign w6078 = w17821 & ~w2690;
assign w6079 = ~w17537 & ~w13443;
assign w6080 = ~w10000 & w17669;
assign w6081 = ~w376 & ~w18146;
assign w6082 = ~w15418 & w9528;
assign w6083 = a_1 & a_43;
assign w6084 = ~w14617 & w8194;
assign w6085 = ~w13677 & ~w2433;
assign w6086 = ~w1671 & w13389;
assign w6087 = w12404 & ~w6136;
assign w6088 = ~w17109 & ~w17623;
assign w6089 = ~w9098 & ~w652;
assign w6090 = w1034 & ~w2063;
assign w6091 = w9475 & w17252;
assign w6092 = w18575 & w4936;
assign w6093 = ~w2111 & w14730;
assign w6094 = ~w2131 & ~w314;
assign w6095 = (~w11815 & ~w18028) | (~w11815 & w15348) | (~w18028 & w15348);
assign w6096 = ~w18576 & ~w19037;
assign w6097 = a_26 & a_54;
assign w6098 = ~w18643 & ~w13310;
assign w6099 = w3183 & w3130;
assign w6100 = a_16 & a_24;
assign w6101 = ~w538 & ~w10368;
assign w6102 = ~w7823 & ~w449;
assign w6103 = w7479 & ~w14573;
assign w6104 = ~w13962 & w8553;
assign w6105 = ~w92 & ~w6070;
assign w6106 = ~w10609 & ~w10173;
assign w6107 = ~w10645 & w18697;
assign w6108 = ~w18521 & ~w7471;
assign w6109 = ~w12685 & ~w17130;
assign w6110 = ~w5287 & ~w5887;
assign w6111 = ~w17921 & ~w8278;
assign w6112 = ~w2518 & ~w2578;
assign w6113 = ~w7840 & ~w12200;
assign w6114 = w17576 & ~w1242;
assign w6115 = ~w6770 & ~w4229;
assign w6116 = w10305 & w3956;
assign w6117 = ~w13277 & ~w7202;
assign w6118 = ~w6912 & ~w3884;
assign w6119 = ~w1857 & ~w17934;
assign w6120 = ~w6411 & ~w505;
assign w6121 = ~w9979 & w12483;
assign w6122 = ~w4792 & ~w11681;
assign w6123 = ~w13005 & ~w4811;
assign w6124 = w7689 & ~w2347;
assign w6125 = ~w19001 & w9799;
assign w6126 = (w5081 & w1888) | (w5081 & w14098) | (w1888 & w14098);
assign w6127 = w10617 & w6449;
assign w6128 = a_29 & a_44;
assign w6129 = w17367 & ~w8542;
assign w6130 = ~w16533 & ~w12443;
assign w6131 = w12753 & ~w12005;
assign w6132 = ~w1662 & ~w9066;
assign w6133 = w2858 & w5359;
assign w6134 = ~w16531 & ~w8131;
assign w6135 = ~w18097 & ~w18585;
assign w6136 = w15397 & w5158;
assign w6137 = ~w14020 & ~w14469;
assign w6138 = w5199 & ~w6400;
assign w6139 = ~w541 & ~w5718;
assign w6140 = w16209 & w4974;
assign w6141 = a_1 & a_50;
assign w6142 = (w15080 & w1399) | (w15080 & w14063) | (w1399 & w14063);
assign w6143 = ~w14470 & w236;
assign w6144 = ~w11586 & ~w3902;
assign w6145 = ~w10878 & ~w14764;
assign w6146 = a_21 & a_47;
assign w6147 = ~w1897 & w2200;
assign w6148 = ~w15864 & ~w3976;
assign w6149 = w9039 & ~w5599;
assign w6150 = w15823 & w7139;
assign w6151 = ~w16114 & ~w2561;
assign w6152 = w2197 & w8159;
assign w6153 = ~w4858 & ~w11843;
assign w6154 = ~w6550 & ~w3115;
assign w6155 = a_13 & a_61;
assign w6156 = ~w5339 & w3515;
assign w6157 = w13713 & w1030;
assign w6158 = ~w10676 & ~w5135;
assign w6159 = ~w6545 & w709;
assign w6160 = ~w2450 & ~w4185;
assign w6161 = (~w18200 & w17737) | (~w18200 & w2535) | (w17737 & w2535);
assign w6162 = ~w5951 & ~w19054;
assign w6163 = ~w7669 & ~w8009;
assign w6164 = w4420 & w994;
assign w6165 = ~w12589 & ~w11544;
assign w6166 = ~w7518 & ~w13888;
assign w6167 = ~w4312 & w15061;
assign w6168 = w2079 & ~w12126;
assign w6169 = ~w12622 & ~w16172;
assign w6170 = w1980 & ~w18952;
assign w6171 = ~w7305 & ~w9177;
assign w6172 = ~w3330 & w16479;
assign w6173 = w653 & w14071;
assign w6174 = ~w9435 & ~w17627;
assign w6175 = ~w11083 & ~w931;
assign w6176 = ~w11620 & ~w9121;
assign w6177 = ~w14235 & ~w1877;
assign w6178 = ~w13633 & ~w6871;
assign w6179 = w14130 & ~w15481;
assign w6180 = ~w6438 & ~w4284;
assign w6181 = ~w176 & ~w10128;
assign w6182 = ~w14305 & ~w16503;
assign w6183 = w8320 & ~w3454;
assign w6184 = a_10 & a_58;
assign w6185 = ~w15644 & w13777;
assign w6186 = ~w4328 & w3071;
assign w6187 = ~w1117 & ~w15627;
assign w6188 = ~w13702 & ~w8764;
assign w6189 = a_6 & a_31;
assign w6190 = ~w18017 & w15243;
assign w6191 = ~w8498 & ~w8031;
assign w6192 = ~w12068 & ~w12557;
assign w6193 = ~w16657 & ~w13509;
assign w6194 = ~w4809 & ~w16670;
assign w6195 = ~w518 & ~w4500;
assign w6196 = ~w17087 & ~w7618;
assign w6197 = ~w16147 & w2352;
assign w6198 = ~w5174 & ~w16451;
assign w6199 = ~w6728 & w15393;
assign w6200 = ~w8587 & ~w1321;
assign w6201 = (~w17101 & w17665) | (~w17101 & w16522) | (w17665 & w16522);
assign w6202 = ~w6278 & w14553;
assign w6203 = ~w14699 & w12740;
assign w6204 = ~w370 & w12057;
assign w6205 = ~w8230 & ~w1866;
assign w6206 = a_53 & a_60;
assign w6207 = w10651 & ~w7739;
assign w6208 = w8156 & w15517;
assign w6209 = ~w11106 & ~w4370;
assign w6210 = w5943 & ~w4273;
assign w6211 = a_15 & a_48;
assign w6212 = ~w10988 & w6952;
assign w6213 = ~w1016 & w6071;
assign w6214 = w18346 & w16036;
assign w6215 = (w13215 & w18660) | (w13215 & w6976) | (w18660 & w6976);
assign w6216 = a_26 & a_43;
assign w6217 = w16252 & w2056;
assign w6218 = w12439 & w5131;
assign w6219 = w3296 & ~w2432;
assign w6220 = (~w980 & ~w12312) | (~w980 & w15633) | (~w12312 & w15633);
assign w6221 = (w10529 & w961) | (w10529 & w18128) | (w961 & w18128);
assign w6222 = ~w4061 & ~w10215;
assign w6223 = ~w11452 & ~w1918;
assign w6224 = ~w13237 & ~w16879;
assign w6225 = ~w7122 & ~w13136;
assign w6226 = ~w12100 & ~w15426;
assign w6227 = ~w18769 & w2812;
assign w6228 = ~w4406 & ~w7907;
assign w6229 = ~w9525 & w15327;
assign w6230 = ~w12917 & w6295;
assign w6231 = ~w2563 & w11206;
assign w6232 = ~w15459 & ~w18667;
assign w6233 = w10269 & ~w5096;
assign w6234 = ~w9258 & w4753;
assign w6235 = ~w11154 & w1471;
assign w6236 = (~w18816 & ~w11394) | (~w18816 & w9397) | (~w11394 & w9397);
assign w6237 = ~w10246 & ~w17876;
assign w6238 = ~w12696 & ~w360;
assign w6239 = ~w6090 & ~w9057;
assign w6240 = ~w539 & ~w15221;
assign w6241 = ~w1953 & ~w5892;
assign w6242 = (w11700 & w10414) | (w11700 & w9709) | (w10414 & w9709);
assign w6243 = ~w17951 & ~w15639;
assign w6244 = w1836 & w11888;
assign w6245 = w8089 & ~w2651;
assign w6246 = (w8169 & w19005) | (w8169 & w13481) | (w19005 & w13481);
assign w6247 = ~w9928 & ~w2826;
assign w6248 = a_3 & a_52;
assign w6249 = w3492 & ~w18561;
assign w6250 = ~w15360 & ~w3762;
assign w6251 = (~w19005 & w757) | (~w19005 & w13704) | (w757 & w13704);
assign w6252 = a_9 & a_36;
assign w6253 = ~w8022 & ~w15731;
assign w6254 = w9748 & w3649;
assign w6255 = ~w18257 & w11868;
assign w6256 = w13390 & w8211;
assign w6257 = w18329 & w13046;
assign w6258 = w13438 & w8614;
assign w6259 = ~w2580 & w14474;
assign w6260 = w1172 & w2094;
assign w6261 = ~w9841 & ~w13848;
assign w6262 = w1846 & ~w8286;
assign w6263 = ~w8065 & ~w15597;
assign w6264 = w2348 & w13009;
assign w6265 = ~w6818 & ~w5920;
assign w6266 = ~w16860 & ~w11548;
assign w6267 = ~w18725 & ~w6901;
assign w6268 = ~w13640 & ~w11167;
assign w6269 = ~w16512 & ~w3888;
assign w6270 = ~w8111 & ~w12833;
assign w6271 = ~w3404 & ~w6630;
assign w6272 = ~w17228 & ~w15680;
assign w6273 = (w8250 & ~w13082) | (w8250 & w17693) | (~w13082 & w17693);
assign w6274 = ~w7483 & ~w14793;
assign w6275 = ~w15589 & ~w10797;
assign w6276 = ~w3717 & w12011;
assign w6277 = a_48 & a_55;
assign w6278 = ~w512 & ~w12344;
assign w6279 = w13037 & w9139;
assign w6280 = w11494 & w9445;
assign w6281 = ~w5535 & ~w10768;
assign w6282 = a_29 & a_42;
assign w6283 = ~w2427 & ~w10879;
assign w6284 = ~w17422 & w13483;
assign w6285 = ~w17495 & w18862;
assign w6286 = ~w19069 & w949;
assign w6287 = ~w13408 & ~w9862;
assign w6288 = ~w1074 & w14429;
assign w6289 = ~w8391 & ~w4942;
assign w6290 = ~w15610 & w9793;
assign w6291 = (w152 & w15862) | (w152 & w1934) | (w15862 & w1934);
assign w6292 = ~w14531 & w18622;
assign w6293 = (~w4683 & ~w5921) | (~w4683 & w11571) | (~w5921 & w11571);
assign w6294 = (~w6115 & ~w11089) | (~w6115 & w5550) | (~w11089 & w5550);
assign w6295 = ~w3806 & ~w12578;
assign w6296 = ~w18830 & ~w13766;
assign w6297 = ~w11226 & ~w5950;
assign w6298 = ~w14424 & w10822;
assign w6299 = w5593 & ~w13401;
assign w6300 = (w18980 & w6334) | (w18980 & w3853) | (w6334 & w3853);
assign w6301 = w16915 & ~w12724;
assign w6302 = ~w9662 & ~w8798;
assign w6303 = ~w14874 & ~w6497;
assign w6304 = a_28 & a_61;
assign w6305 = ~w1557 & ~w15290;
assign w6306 = a_17 & a_23;
assign w6307 = (w16917 & w470) | (w16917 & w340) | (w470 & w340);
assign w6308 = w7149 & ~w477;
assign w6309 = ~w12022 & ~w1799;
assign w6310 = (w7768 & w16197) | (w7768 & w4977) | (w16197 & w4977);
assign w6311 = ~w10416 & ~w8938;
assign w6312 = w4772 & ~w13190;
assign w6313 = ~w11415 & ~w9614;
assign w6314 = ~w16366 & ~w6208;
assign w6315 = (~w4374 & ~w3171) | (~w4374 & w1970) | (~w3171 & w1970);
assign w6316 = ~w5495 & w87;
assign w6317 = ~w17223 & ~w4995;
assign w6318 = ~w17728 & ~w18671;
assign w6319 = (w7102 & w2350) | (w7102 & w14611) | (w2350 & w14611);
assign w6320 = ~w10758 & ~w5572;
assign w6321 = ~w13468 & ~w18135;
assign w6322 = ~w17314 & ~w17108;
assign w6323 = ~w11373 & ~w13218;
assign w6324 = w16695 & w17788;
assign w6325 = ~w8960 & ~w8537;
assign w6326 = (a_56 & w15289) | (a_56 & w9313) | (w15289 & w9313);
assign w6327 = w10230 & ~w18204;
assign w6328 = ~w491 & w1818;
assign w6329 = ~w15500 & ~w15914;
assign w6330 = a_42 & a_56;
assign w6331 = w14435 & ~w13195;
assign w6332 = ~w6388 & w8671;
assign w6333 = ~w4904 & ~w52;
assign w6334 = w5142 | w14650;
assign w6335 = ~w9250 & ~w11391;
assign w6336 = ~w14508 & w16603;
assign w6337 = a_36 & a_59;
assign w6338 = ~w13022 & ~w17806;
assign w6339 = ~w18964 & w19085;
assign w6340 = w3431 & w8853;
assign w6341 = ~w3549 & ~w5256;
assign w6342 = ~w9621 & ~w72;
assign w6343 = ~w5429 & ~w16884;
assign w6344 = ~w16928 & ~w10162;
assign w6345 = ~w11645 & w3640;
assign w6346 = ~w5289 & w16688;
assign w6347 = ~w7610 & ~w11204;
assign w6348 = ~w3583 & ~w1718;
assign w6349 = ~w8160 & ~w10918;
assign w6350 = ~w10114 & w6516;
assign w6351 = ~w9442 & ~w17186;
assign w6352 = ~w10083 & w9955;
assign w6353 = ~w9856 & ~w11775;
assign w6354 = ~w755 & ~w7650;
assign w6355 = ~w18132 & ~w14828;
assign w6356 = (~w4834 & ~w7090) | (~w4834 & w5815) | (~w7090 & w5815);
assign w6357 = (~w18538 & ~w9923) | (~w18538 & w12119) | (~w9923 & w12119);
assign w6358 = ~w846 & ~w9485;
assign w6359 = ~w12030 & ~w7350;
assign w6360 = ~w13912 & w4429;
assign w6361 = (~w14436 & w14974) | (~w14436 & w15844) | (w14974 & w15844);
assign w6362 = w9016 & ~w8095;
assign w6363 = a_6 & a_55;
assign w6364 = (~w7887 & ~w1400) | (~w7887 & w12525) | (~w1400 & w12525);
assign w6365 = w13633 & w6871;
assign w6366 = ~w14087 & w18843;
assign w6367 = ~w1172 & ~w2094;
assign w6368 = ~w4517 & ~w4497;
assign w6369 = ~w13265 & ~w12603;
assign w6370 = ~w592 & w18311;
assign w6371 = ~w3925 & w1434;
assign w6372 = ~w2766 & ~w13778;
assign w6373 = ~w7393 & ~w3367;
assign w6374 = ~a_25 & ~w3391;
assign w6375 = ~w9308 & ~w17178;
assign w6376 = ~w15582 & ~w17923;
assign w6377 = w17945 & w9305;
assign w6378 = ~w10352 & ~w16461;
assign w6379 = w10969 & ~w11122;
assign w6380 = ~w15982 & ~w15832;
assign w6381 = ~w3618 & ~w6131;
assign w6382 = a_29 & a_34;
assign w6383 = ~w16856 & ~w3572;
assign w6384 = w4124 & ~w9798;
assign w6385 = ~w17107 & ~w2536;
assign w6386 = ~w12601 & ~w6155;
assign w6387 = a_50 & a_52;
assign w6388 = ~w9028 & ~w16159;
assign w6389 = ~w14971 & ~w18054;
assign w6390 = w15992 & w11138;
assign w6391 = ~w16500 & ~w4943;
assign w6392 = w15692 & ~w15612;
assign w6393 = ~w3036 & w10889;
assign w6394 = w17218 & ~w8412;
assign w6395 = ~w5823 & ~w9272;
assign w6396 = ~w15264 & ~w17326;
assign w6397 = ~w14884 & ~w1971;
assign w6398 = a_17 & a_24;
assign w6399 = ~w18967 & ~w9924;
assign w6400 = ~w11764 & ~w7183;
assign w6401 = ~w3699 & w11722;
assign w6402 = ~w14398 & w13035;
assign w6403 = ~w13883 & ~w6369;
assign w6404 = ~w13067 & w6188;
assign w6405 = ~w3664 & ~w4471;
assign w6406 = ~w8257 & ~w3483;
assign w6407 = (~w1798 & w10330) | (~w1798 & w18955) | (w10330 & w18955);
assign w6408 = ~w9729 & w3025;
assign w6409 = a_4 & a_14;
assign w6410 = ~w3040 & ~w11921;
assign w6411 = ~w4023 & w16904;
assign w6412 = ~w10339 & w16645;
assign w6413 = a_37 & a_43;
assign w6414 = w8151 & ~w8679;
assign w6415 = w2760 & ~w13493;
assign w6416 = (w804 & w18821) | (w804 & w11244) | (w18821 & w11244);
assign w6417 = ~w13707 & ~w6122;
assign w6418 = ~w6476 & ~w2281;
assign w6419 = ~w15524 & ~w15783;
assign w6420 = a_39 & a_56;
assign w6421 = a_40 & a_58;
assign w6422 = ~w3062 & ~w4849;
assign w6423 = ~w18580 & ~w61;
assign w6424 = w10786 & ~w767;
assign w6425 = ~w4143 & w16397;
assign w6426 = ~w999 & w2411;
assign w6427 = (w17256 & ~w6294) | (w17256 & w19058) | (~w6294 & w19058);
assign w6428 = w9841 & w13848;
assign w6429 = ~w18484 & ~w448;
assign w6430 = ~w3913 & w19133;
assign w6431 = ~w1756 & ~w9427;
assign w6432 = ~w5108 & w16025;
assign w6433 = ~w14005 & ~w5299;
assign w6434 = w9999 & ~w16491;
assign w6435 = ~w9559 & ~w3626;
assign w6436 = w28 & w550;
assign w6437 = a_38 & a_54;
assign w6438 = ~w11132 & ~w14942;
assign w6439 = w17967 & w6191;
assign w6440 = w141 & w10727;
assign w6441 = ~w16125 & ~w8398;
assign w6442 = ~w10207 & ~w18046;
assign w6443 = ~w4250 & ~w14292;
assign w6444 = w6761 & w17873;
assign w6445 = w4749 & ~w18784;
assign w6446 = ~w2038 & ~w14526;
assign w6447 = a_13 & a_42;
assign w6448 = w1048 & ~w4951;
assign w6449 = ~w18368 & ~w18530;
assign w6450 = ~w11417 & w17099;
assign w6451 = w1867 & w72;
assign w6452 = w3078 & ~w4969;
assign w6453 = (~w2095 & ~w10734) | (~w2095 & w18122) | (~w10734 & w18122);
assign w6454 = ~w7849 & ~w9015;
assign w6455 = w897 & ~w1981;
assign w6456 = ~w11148 & ~w15014;
assign w6457 = ~w16420 & ~w19111;
assign w6458 = a_20 & a_52;
assign w6459 = w4133 & ~w145;
assign w6460 = a_54 & a_59;
assign w6461 = ~w3999 & ~w2018;
assign w6462 = ~w11471 & ~w4260;
assign w6463 = ~w4692 & w6037;
assign w6464 = ~w13175 & w14386;
assign w6465 = ~w13296 & ~w14291;
assign w6466 = ~w13094 & w7333;
assign w6467 = ~w13028 & w4360;
assign w6468 = (~w17442 & ~w12985) | (~w17442 & w16774) | (~w12985 & w16774);
assign w6469 = (~w120 & w15526) | (~w120 & w12403) | (w15526 & w12403);
assign w6470 = ~w18578 & ~w15129;
assign w6471 = ~w4200 & ~w3571;
assign w6472 = w14277 & w3020;
assign w6473 = (~w16689 & ~w18127) | (~w16689 & w1646) | (~w18127 & w1646);
assign w6474 = a_1 & a_62;
assign w6475 = ~w1468 & ~w2586;
assign w6476 = ~w1582 & ~w6008;
assign w6477 = ~w9247 & ~w324;
assign w6478 = ~w15888 & w19052;
assign w6479 = ~w9312 & ~w18939;
assign w6480 = ~w1194 & w11892;
assign w6481 = a_4 & w15464;
assign w6482 = w18911 & ~w1520;
assign w6483 = ~w2313 & ~w6030;
assign w6484 = ~w13429 & ~w9263;
assign w6485 = ~w3002 & ~w15543;
assign w6486 = w11108 & ~w9354;
assign w6487 = ~w14423 & ~w13671;
assign w6488 = ~w5922 & ~w7935;
assign w6489 = ~w8143 & w8315;
assign w6490 = w2307 & ~w15165;
assign w6491 = (~w1433 & ~w14920) | (~w1433 & w16455) | (~w14920 & w16455);
assign w6492 = w8603 & w6654;
assign w6493 = ~w7701 & w5939;
assign w6494 = w18648 & ~w3271;
assign w6495 = ~w9931 & ~w10963;
assign w6496 = ~w15395 & ~w371;
assign w6497 = (~w2769 & w6164) | (~w2769 & w12109) | (w6164 & w12109);
assign w6498 = ~w10498 & w3094;
assign w6499 = w3101 & ~w5648;
assign w6500 = a_26 & a_33;
assign w6501 = ~w1935 & ~w8547;
assign w6502 = ~w16402 & ~w18988;
assign w6503 = ~w12791 & ~w17465;
assign w6504 = ~w7494 & w16259;
assign w6505 = ~w16447 & w14300;
assign w6506 = w5078 & w12452;
assign w6507 = ~w3207 & ~w14866;
assign w6508 = ~w2160 & ~w10741;
assign w6509 = ~w5796 & ~w9548;
assign w6510 = ~w16971 & ~w16354;
assign w6511 = a_31 & a_56;
assign w6512 = w13036 & ~w8517;
assign w6513 = ~w8158 & ~w6580;
assign w6514 = ~w1800 & ~w918;
assign w6515 = w3833 & w3818;
assign w6516 = ~w8452 & w16724;
assign w6517 = ~w18763 & ~w4985;
assign w6518 = ~w16255 & ~w6410;
assign w6519 = a_3 & a_45;
assign w6520 = ~w13602 & ~w1203;
assign w6521 = a_3 & a_15;
assign w6522 = w9506 & ~w7296;
assign w6523 = ~w8476 & ~w6005;
assign w6524 = (~w10490 & ~w2234) | (~w10490 & w871) | (~w2234 & w871);
assign w6525 = w4856 & w3996;
assign w6526 = ~w15978 & ~w12634;
assign w6527 = ~w6041 & ~w8792;
assign w6528 = w5438 & ~w1923;
assign w6529 = a_51 & a_57;
assign w6530 = ~w5651 & ~w3663;
assign w6531 = a_8 & a_17;
assign w6532 = w4320 & ~w6468;
assign w6533 = ~w8217 & ~w13272;
assign w6534 = a_2 & a_8;
assign w6535 = ~w18754 & ~w2199;
assign w6536 = w13617 & w3831;
assign w6537 = ~w15988 & w14815;
assign w6538 = w17809 & ~w9877;
assign w6539 = w6315 & w6617;
assign w6540 = ~w3239 & w9940;
assign w6541 = a_10 & a_48;
assign w6542 = (~w12947 & ~w14364) | (~w12947 & w17683) | (~w14364 & w17683);
assign w6543 = a_35 & a_56;
assign w6544 = w17161 & w18997;
assign w6545 = a_51 & a_63;
assign w6546 = ~w10856 & ~w2487;
assign w6547 = ~w11384 & ~w47;
assign w6548 = ~w13700 & ~w1715;
assign w6549 = ~w10296 & ~w17035;
assign w6550 = a_35 & a_40;
assign w6551 = w12477 & w5378;
assign w6552 = w252 & w7934;
assign w6553 = ~w10414 & ~w10443;
assign w6554 = ~w11412 & w12151;
assign w6555 = w10851 & w2563;
assign w6556 = ~w16992 & w14491;
assign w6557 = w1054 & ~w14009;
assign w6558 = w797 & w17459;
assign w6559 = ~w5564 & w2091;
assign w6560 = a_17 & a_44;
assign w6561 = w15622 & ~w10036;
assign w6562 = w13825 & w5273;
assign w6563 = (~w5786 & ~w9743) | (~w5786 & w12392) | (~w9743 & w12392);
assign w6564 = ~w8629 & ~w8596;
assign w6565 = ~w11650 & ~w3680;
assign w6566 = a_54 & a_60;
assign w6567 = (w13150 & w666) | (w13150 & w18282) | (w666 & w18282);
assign w6568 = a_25 & a_41;
assign w6569 = ~w12050 & ~w8833;
assign w6570 = ~w5608 & ~w11088;
assign w6571 = ~w17322 & ~w16149;
assign w6572 = ~w14982 & w8164;
assign w6573 = w9340 & ~w2222;
assign w6574 = w6856 & ~w5357;
assign w6575 = ~w4818 & ~w1204;
assign w6576 = ~w16640 & w2811;
assign w6577 = ~w17950 & w13156;
assign w6578 = ~w11005 & ~w13641;
assign w6579 = ~w5990 & w18358;
assign w6580 = w18276 & w4893;
assign w6581 = w9707 & w10366;
assign w6582 = ~w15346 & ~w16835;
assign w6583 = w1839 & ~w14322;
assign w6584 = ~w16165 & ~w4051;
assign w6585 = a_13 & a_24;
assign w6586 = w11469 & ~w2733;
assign w6587 = ~w14745 & w18068;
assign w6588 = a_0 & a_7;
assign w6589 = (w2352 & w13558) | (w2352 & ~w13186) | (w13558 & ~w13186);
assign w6590 = ~w15134 & w17889;
assign w6591 = w14996 & w7991;
assign w6592 = ~w16644 & ~w661;
assign w6593 = a_13 & ~w17557;
assign w6594 = ~w15446 & ~w17570;
assign w6595 = ~w7985 & ~w12494;
assign w6596 = ~w1577 & w6594;
assign w6597 = ~w13460 & ~w17364;
assign w6598 = ~w50 & ~w15588;
assign w6599 = ~w11546 & ~w18810;
assign w6600 = w5516 & ~w8281;
assign w6601 = w11107 & w16322;
assign w6602 = ~w13177 & ~w18857;
assign w6603 = ~w15495 & ~w8949;
assign w6604 = ~w15100 & ~w519;
assign w6605 = w12252 & ~w8856;
assign w6606 = w18001 & w12515;
assign w6607 = w3016 & w17002;
assign w6608 = ~w5532 & ~w10213;
assign w6609 = ~w18228 & w9311;
assign w6610 = ~w16185 & ~w6470;
assign w6611 = ~w11316 & ~w217;
assign w6612 = ~w3139 & w6993;
assign w6613 = w15616 & w14;
assign w6614 = ~w11104 & ~w17749;
assign w6615 = w1889 & ~w7549;
assign w6616 = ~w15861 & w16045;
assign w6617 = (~w14350 & ~w3230) | (~w14350 & w4016) | (~w3230 & w4016);
assign w6618 = ~w11922 & ~w12545;
assign w6619 = ~w2019 & ~w7123;
assign w6620 = w16296 & w14482;
assign w6621 = ~w9267 & ~w10973;
assign w6622 = ~w16756 & ~w4810;
assign w6623 = ~w14385 & ~w11679;
assign w6624 = w16560 & w13405;
assign w6625 = ~w3499 & ~w9546;
assign w6626 = ~w14149 & ~w10425;
assign w6627 = ~w18176 & ~w16047;
assign w6628 = ~w8907 & ~w1520;
assign w6629 = ~w4839 & ~w11746;
assign w6630 = ~w14595 & ~w18642;
assign w6631 = ~w6146 & ~w219;
assign w6632 = w17544 & ~w11931;
assign w6633 = ~w5622 & ~w13333;
assign w6634 = ~w11273 & ~w10948;
assign w6635 = ~w14803 & ~w17287;
assign w6636 = ~w102 & ~w18319;
assign w6637 = ~w16819 & ~w9511;
assign w6638 = ~w1041 & w6446;
assign w6639 = w15407 & ~w13658;
assign w6640 = ~w3994 & ~w524;
assign w6641 = ~w16805 & ~w9886;
assign w6642 = ~w10761 & w7310;
assign w6643 = ~w13795 & ~w12500;
assign w6644 = ~w16390 & ~w16407;
assign w6645 = w16659 & ~w18359;
assign w6646 = ~w8101 & w7951;
assign w6647 = a_0 & a_62;
assign w6648 = w491 & ~w1818;
assign w6649 = w18304 & ~w3430;
assign w6650 = (~w4041 & ~w358) | (~w4041 & w5481) | (~w358 & w5481);
assign w6651 = w17580 & ~w8072;
assign w6652 = w12098 & ~w1475;
assign w6653 = (w16437 & w9221) | (w16437 & w3541) | (w9221 & w3541);
assign w6654 = ~w8779 & ~w12662;
assign w6655 = a_3 & a_44;
assign w6656 = ~w4161 & w15210;
assign w6657 = w14418 & w8034;
assign w6658 = w6677 & ~w18026;
assign w6659 = w4890 & w13819;
assign w6660 = ~w6772 & ~w12030;
assign w6661 = ~w12731 & ~w13245;
assign w6662 = w17571 & w12852;
assign w6663 = ~w3157 & ~w9191;
assign w6664 = ~w16060 & ~w7778;
assign w6665 = w13227 & ~w6250;
assign w6666 = a_9 & a_14;
assign w6667 = ~w9428 & ~w4855;
assign w6668 = ~w5538 & ~w13057;
assign w6669 = ~w14446 & ~w3857;
assign w6670 = ~w2743 & w1862;
assign w6671 = w16554 & w6618;
assign w6672 = ~w7915 & w5143;
assign w6673 = w15602 & ~w10032;
assign w6674 = w6001 & ~w2562;
assign w6675 = ~w15197 & ~w9306;
assign w6676 = ~w12739 & ~w15322;
assign w6677 = ~w8117 & ~w8769;
assign w6678 = ~w3686 & ~w3974;
assign w6679 = w10794 & w6710;
assign w6680 = ~w8327 & ~w16415;
assign w6681 = ~w16824 & ~w11220;
assign w6682 = (~w2769 & w2730) | (~w2769 & w15062) | (w2730 & w15062);
assign w6683 = w1983 & w15552;
assign w6684 = ~w15289 & w718;
assign w6685 = w3180 & w1219;
assign w6686 = ~w2658 & ~w9823;
assign w6687 = w16825 & w16873;
assign w6688 = ~w16502 & ~w463;
assign w6689 = w18458 & ~w12034;
assign w6690 = w7399 & ~w10764;
assign w6691 = ~w5935 & ~w8180;
assign w6692 = w3997 & ~w14676;
assign w6693 = ~w2663 & w19159;
assign w6694 = ~w6777 & w15253;
assign w6695 = w11092 & w4781;
assign w6696 = ~w11346 & ~w10661;
assign w6697 = w18240 & ~w3174;
assign w6698 = ~w7726 & ~w18981;
assign w6699 = ~w4592 & ~w18371;
assign w6700 = ~w1361 & ~w673;
assign w6701 = a_10 & a_55;
assign w6702 = ~w12290 & ~w8621;
assign w6703 = ~w9531 & ~w7179;
assign w6704 = ~w6027 & ~w4167;
assign w6705 = a_16 & a_20;
assign w6706 = w9630 & w18739;
assign w6707 = w2359 & ~w4851;
assign w6708 = ~w1235 & ~w3252;
assign w6709 = ~w15338 & ~w18941;
assign w6710 = ~w287 & ~w11007;
assign w6711 = w4462 & w13427;
assign w6712 = w5723 & ~w9246;
assign w6713 = w16318 & ~w15283;
assign w6714 = ~w11644 & w16802;
assign w6715 = ~w16540 & ~w4802;
assign w6716 = w8519 & ~w6402;
assign w6717 = ~w1058 & ~w15546;
assign w6718 = ~w3219 & w6405;
assign w6719 = ~w7925 & ~w17015;
assign w6720 = ~w5128 & ~w17847;
assign w6721 = ~w6085 & ~w2433;
assign w6722 = ~w15596 & ~w9783;
assign w6723 = ~w13493 & ~w17487;
assign w6724 = ~w15480 & ~w12088;
assign w6725 = ~w7492 & w17891;
assign w6726 = w14820 & ~w18593;
assign w6727 = ~w9053 & ~w15314;
assign w6728 = ~w8109 & ~w2119;
assign w6729 = w10942 & w3366;
assign w6730 = ~w9654 & w10142;
assign w6731 = ~w630 & ~w4884;
assign w6732 = w11333 & ~w18408;
assign w6733 = ~w14848 & ~w692;
assign w6734 = (~w16818 & w3477) | (~w16818 & w18839) | (w3477 & w18839);
assign w6735 = ~w8930 & w27;
assign w6736 = a_45 & a_59;
assign w6737 = w6982 & w16440;
assign w6738 = a_12 & a_17;
assign w6739 = a_28 & a_44;
assign w6740 = (w7350 & w4155) | (w7350 & w7023) | (w4155 & w7023);
assign w6741 = ~w8466 & ~w8524;
assign w6742 = ~w6990 & ~w12517;
assign w6743 = ~a_40 & a_41;
assign w6744 = ~w696 & ~w10856;
assign w6745 = ~w12949 & ~w8924;
assign w6746 = w11623 & ~w8761;
assign w6747 = ~w18788 & ~w11880;
assign w6748 = w6661 & w16611;
assign w6749 = a_43 & a_48;
assign w6750 = ~w10180 & w14093;
assign w6751 = ~w952 & ~w3133;
assign w6752 = ~w13388 & ~w5336;
assign w6753 = ~w8401 & ~w1979;
assign w6754 = w868 & ~w9919;
assign w6755 = ~w15935 & w17102;
assign w6756 = ~w6729 & ~w2144;
assign w6757 = ~w5574 & w17621;
assign w6758 = ~w257 & ~w11284;
assign w6759 = ~w12529 & ~w6361;
assign w6760 = ~w13837 & w12099;
assign w6761 = ~w19131 & ~w3892;
assign w6762 = (w7102 & w1726) | (w7102 & w6014) | (w1726 & w6014);
assign w6763 = w14165 & ~w1270;
assign w6764 = w3075 & ~w2852;
assign w6765 = ~w5486 & w863;
assign w6766 = ~w13125 & ~w5215;
assign w6767 = ~w6215 & ~w11720;
assign w6768 = ~w2316 & ~w1370;
assign w6769 = ~w14173 & ~w9163;
assign w6770 = (~w13570 & ~w8911) | (~w13570 & w16804) | (~w8911 & w16804);
assign w6771 = ~w13216 & ~w7623;
assign w6772 = w18156 & ~w129;
assign w6773 = ~w8033 & ~w4490;
assign w6774 = ~w16718 & ~w19044;
assign w6775 = w6241 & w15581;
assign w6776 = ~w15861 & w5410;
assign w6777 = a_10 & a_20;
assign w6778 = ~w14535 & ~w12417;
assign w6779 = w5780 & w14500;
assign w6780 = ~w12983 & w14109;
assign w6781 = ~w16128 & ~w8642;
assign w6782 = ~w17357 & ~w2856;
assign w6783 = w7551 & w968;
assign w6784 = w5273 & w2883;
assign w6785 = w3800 & ~w14913;
assign w6786 = ~w17627 & ~w18540;
assign w6787 = w17976 & w18649;
assign w6788 = ~w672 & ~w13871;
assign w6789 = w14492 & ~w16385;
assign w6790 = w4196 & w4471;
assign w6791 = (w2352 & w13945) | (w2352 & w11689) | (w13945 & w11689);
assign w6792 = ~w12045 & ~w7124;
assign w6793 = w12678 & ~w12283;
assign w6794 = ~w14051 & w8474;
assign w6795 = w2541 & w2047;
assign w6796 = ~w12008 & w10239;
assign w6797 = w3334 & w16705;
assign w6798 = ~w951 & ~w17865;
assign w6799 = w11148 & w15014;
assign w6800 = w17444 & ~w11367;
assign w6801 = ~w16808 & w8392;
assign w6802 = w13186 & w14993;
assign w6803 = ~a_36 & ~w8906;
assign w6804 = w16151 & ~w8583;
assign w6805 = w6728 & ~w15393;
assign w6806 = ~w6211 & w15863;
assign w6807 = w5190 & w3233;
assign w6808 = ~w1502 & w6351;
assign w6809 = ~w6513 & ~w12911;
assign w6810 = w18433 & ~w6715;
assign w6811 = a_23 & a_63;
assign w6812 = w11960 & ~w16648;
assign w6813 = w9868 & w7995;
assign w6814 = a_19 & a_59;
assign w6815 = ~w6841 & ~w14898;
assign w6816 = w6960 & ~w14685;
assign w6817 = w8229 & ~w398;
assign w6818 = w2937 & ~w7159;
assign w6819 = ~w2513 & ~w12426;
assign w6820 = ~w11181 & ~w10868;
assign w6821 = w2627 & w7415;
assign w6822 = w14656 & ~w741;
assign w6823 = ~w13863 & ~w15444;
assign w6824 = w8998 & ~w13977;
assign w6825 = ~w17551 & ~w6814;
assign w6826 = ~w4556 & w12899;
assign w6827 = ~w2196 & ~w18803;
assign w6828 = w10812 & ~w15952;
assign w6829 = ~w13316 & ~w18391;
assign w6830 = w14431 & w3457;
assign w6831 = w1312 & ~w7654;
assign w6832 = w13089 & ~w12347;
assign w6833 = w4905 & w12819;
assign w6834 = (~w152 & w3531) | (~w152 & w8713) | (w3531 & w8713);
assign w6835 = w16601 & ~w1834;
assign w6836 = ~w18926 & ~w1231;
assign w6837 = ~w2979 & ~w16111;
assign w6838 = ~w15663 & ~w16181;
assign w6839 = ~w15308 & ~w18223;
assign w6840 = ~w4312 & ~w1391;
assign w6841 = a_5 & a_31;
assign w6842 = (~w14439 & ~w6987) | (~w14439 & w3164) | (~w6987 & w3164);
assign w6843 = ~w7517 & w10965;
assign w6844 = w2426 & w3079;
assign w6845 = ~w13524 & ~w5437;
assign w6846 = a_31 & a_63;
assign w6847 = a_4 & a_56;
assign w6848 = ~w18750 & ~w1071;
assign w6849 = ~w4290 & ~w9343;
assign w6850 = ~w4454 & ~w3965;
assign w6851 = w11273 & w5551;
assign w6852 = w10879 & ~w2339;
assign w6853 = w7594 & w10869;
assign w6854 = w9990 & ~w8754;
assign w6855 = ~w17344 & ~w580;
assign w6856 = ~w16872 & ~w5719;
assign w6857 = ~w9799 & w19001;
assign w6858 = ~w18364 & ~w1560;
assign w6859 = w183 & w18999;
assign w6860 = a_50 & a_60;
assign w6861 = w3051 & w12286;
assign w6862 = ~w6745 & ~w11356;
assign w6863 = ~w17389 & ~w1230;
assign w6864 = ~w14329 & w1846;
assign w6865 = (~w17627 & ~w6786) | (~w17627 & w6174) | (~w6786 & w6174);
assign w6866 = ~w15623 & ~w15799;
assign w6867 = ~w1088 & ~w12744;
assign w6868 = w1196 & w4479;
assign w6869 = w11829 & w15363;
assign w6870 = ~w10804 & ~w5185;
assign w6871 = ~w4186 & ~w11153;
assign w6872 = w12679 & ~w13870;
assign w6873 = a_21 & a_60;
assign w6874 = ~w8053 & ~w6012;
assign w6875 = a_0 & a_43;
assign w6876 = ~w13830 & ~w11748;
assign w6877 = ~w4952 & ~w10671;
assign w6878 = w17753 & ~w8265;
assign w6879 = w15248 & w8290;
assign w6880 = w721 & ~w543;
assign w6881 = ~w2304 & w1510;
assign w6882 = ~w3189 & ~w15150;
assign w6883 = ~w3070 & ~w2831;
assign w6884 = w13361 & w11561;
assign w6885 = ~w11657 & ~w13747;
assign w6886 = ~w17119 & ~w12567;
assign w6887 = a_33 & a_50;
assign w6888 = w3637 & ~w16231;
assign w6889 = ~w2045 & w5227;
assign w6890 = ~w12347 & w11659;
assign w6891 = w12536 & w14464;
assign w6892 = w13082 & ~w11001;
assign w6893 = w1780 & ~w6856;
assign w6894 = ~w10100 & ~w12476;
assign w6895 = ~w14574 & ~w12817;
assign w6896 = ~w17929 & ~w18807;
assign w6897 = w10008 & w8332;
assign w6898 = ~w15744 & w10595;
assign w6899 = ~w1707 & ~w8114;
assign w6900 = ~w17054 & w8465;
assign w6901 = ~w16249 & w16023;
assign w6902 = w12552 & ~w137;
assign w6903 = ~w11658 & ~w5666;
assign w6904 = w6376 & ~w686;
assign w6905 = w286 & w13027;
assign w6906 = w3818 & ~w9927;
assign w6907 = ~w1527 & ~w2289;
assign w6908 = ~w5699 & w8456;
assign w6909 = w11465 & w3313;
assign w6910 = (~w15437 & ~w7472) | (~w15437 & w15371) | (~w7472 & w15371);
assign w6911 = ~w9399 & ~w1753;
assign w6912 = ~w7675 & ~w1681;
assign w6913 = ~w15861 & w16033;
assign w6914 = ~w13961 & w14880;
assign w6915 = (~w11835 & ~w8264) | (~w11835 & w16553) | (~w8264 & w16553);
assign w6916 = w16413 & w10857;
assign w6917 = ~w8477 & ~w7279;
assign w6918 = w15387 & w14772;
assign w6919 = ~w9924 & ~w18625;
assign w6920 = w2192 & ~w8945;
assign w6921 = w14396 & w7749;
assign w6922 = ~w8225 & ~w10322;
assign w6923 = ~w3671 & ~w3705;
assign w6924 = w12465 & ~w13598;
assign w6925 = ~w800 & ~w2785;
assign w6926 = a_37 & a_51;
assign w6927 = ~w15025 & w7834;
assign w6928 = (~w14839 & ~w17204) | (~w14839 & w17637) | (~w17204 & w17637);
assign w6929 = ~w12538 & ~w15208;
assign w6930 = ~w9926 & ~w14970;
assign w6931 = ~w2435 & ~w7257;
assign w6932 = a_27 & a_60;
assign w6933 = ~w12939 & ~w11915;
assign w6934 = ~w12399 & ~w12348;
assign w6935 = ~w1039 & ~w7954;
assign w6936 = ~w6228 & w1276;
assign w6937 = w16251 & w6771;
assign w6938 = ~w3166 & ~w7600;
assign w6939 = ~w15934 & ~w12490;
assign w6940 = (w15755 & w10668) | (w15755 & w12102) | (w10668 & w12102);
assign w6941 = w13859 & w5294;
assign w6942 = ~w14426 & ~w4639;
assign w6943 = a_35 & a_47;
assign w6944 = ~w6056 & ~w10935;
assign w6945 = w13135 & ~w5681;
assign w6946 = w1320 & w8485;
assign w6947 = w4997 & w4621;
assign w6948 = w12456 & w6794;
assign w6949 = w10893 & ~w18230;
assign w6950 = w13801 & w13138;
assign w6951 = a_18 & a_40;
assign w6952 = (~w4521 & w2278) | (~w4521 & w8237) | (w2278 & w8237);
assign w6953 = ~w10606 & ~w13937;
assign w6954 = ~w7935 & ~w10717;
assign w6955 = ~w2 & w17707;
assign w6956 = ~w10155 & w16711;
assign w6957 = w7608 & ~w4195;
assign w6958 = w17638 & ~w13000;
assign w6959 = w7201 & w4189;
assign w6960 = ~w15242 & ~w4543;
assign w6961 = ~w11877 & ~w1238;
assign w6962 = ~w5833 & ~w12645;
assign w6963 = a_26 & a_29;
assign w6964 = ~w19059 & ~w886;
assign w6965 = a_18 & a_44;
assign w6966 = w10969 & ~w15275;
assign w6967 = ~w2927 & w7718;
assign w6968 = (~w963 & w8052) | (~w963 & w10359) | (w8052 & w10359);
assign w6969 = (~w14817 & ~w8765) | (~w14817 & w1044) | (~w8765 & w1044);
assign w6970 = w9129 & ~w15351;
assign w6971 = ~w4339 & ~w11149;
assign w6972 = ~w5273 & ~w3562;
assign w6973 = w18737 & ~w10564;
assign w6974 = ~w17520 & ~w8378;
assign w6975 = ~w10259 & ~w10440;
assign w6976 = w14309 & w13215;
assign w6977 = w9805 & ~w11807;
assign w6978 = a_52 & a_54;
assign w6979 = ~w1857 & ~w7835;
assign w6980 = ~w252 & ~w6594;
assign w6981 = ~w12814 & ~w15610;
assign w6982 = ~w18759 & ~w13640;
assign w6983 = ~w7008 & w9693;
assign w6984 = ~w11286 & w12689;
assign w6985 = ~w5741 & ~w9156;
assign w6986 = ~w8247 & ~w12358;
assign w6987 = ~w14439 & ~w8129;
assign w6988 = ~w8717 & ~w10939;
assign w6989 = ~w15292 & ~w226;
assign w6990 = a_6 & a_22;
assign w6991 = ~w16948 & ~w13937;
assign w6992 = (w16045 & w2769) | (w16045 & w6616) | (w2769 & w6616);
assign w6993 = ~w17429 & ~w10841;
assign w6994 = ~w4273 & ~w3544;
assign w6995 = ~w7700 & ~w7463;
assign w6996 = ~w18604 & ~w4845;
assign w6997 = ~w7601 & w17666;
assign w6998 = ~w11368 & w18518;
assign w6999 = ~w16318 & w15283;
assign w7000 = w6935 & ~w18263;
assign w7001 = ~w12719 & w17568;
assign w7002 = ~w16483 & w497;
assign w7003 = a_36 & a_55;
assign w7004 = a_14 & a_46;
assign w7005 = ~w4852 & w167;
assign w7006 = w15872 & w12447;
assign w7007 = ~w8532 & w18421;
assign w7008 = w4262 & w14807;
assign w7009 = ~w1953 & w11017;
assign w7010 = ~w7316 & ~w5031;
assign w7011 = w9824 & ~w6075;
assign w7012 = ~w16386 & ~w2373;
assign w7013 = ~w1967 & ~w2006;
assign w7014 = ~w10079 & w8003;
assign w7015 = ~w14085 & w12302;
assign w7016 = ~w4869 & w9698;
assign w7017 = ~w5013 & w8789;
assign w7018 = w14211 & ~w17448;
assign w7019 = ~w10172 & ~w16622;
assign w7020 = a_32 & a_55;
assign w7021 = ~w7533 & ~w8113;
assign w7022 = ~w6712 & ~w1956;
assign w7023 = w6660 & ~w2433;
assign w7024 = ~w4096 & ~w15643;
assign w7025 = ~w10657 & ~w16277;
assign w7026 = w8001 & ~w3601;
assign w7027 = ~w3481 & ~w3386;
assign w7028 = w14530 & ~w7022;
assign w7029 = ~w7515 & ~w11172;
assign w7030 = w14458 & ~w453;
assign w7031 = a_50 & a_51;
assign w7032 = ~w17856 & ~w15051;
assign w7033 = w5631 & ~w13211;
assign w7034 = ~w13708 & ~w1051;
assign w7035 = ~w2115 & ~w16195;
assign w7036 = ~w15481 & ~w9571;
assign w7037 = a_38 & a_51;
assign w7038 = ~w10217 & ~w123;
assign w7039 = (~w3300 & ~w10602) | (~w3300 & w17695) | (~w10602 & w17695);
assign w7040 = w9480 & w2359;
assign w7041 = (~w13457 & w12973) | (~w13457 & w11078) | (w12973 & w11078);
assign w7042 = ~w10298 & w6375;
assign w7043 = ~w890 & ~w1229;
assign w7044 = ~w7314 & w14820;
assign w7045 = w16650 & ~w74;
assign w7046 = ~w8763 & w12473;
assign w7047 = w2004 & w7065;
assign w7048 = a_1 & a_44;
assign w7049 = ~w955 & ~w6035;
assign w7050 = w6500 & ~w665;
assign w7051 = ~w2665 & ~w2671;
assign w7052 = w14725 & ~w15815;
assign w7053 = ~w10241 & ~w8241;
assign w7054 = ~w10329 & ~w16775;
assign w7055 = w6853 & w19102;
assign w7056 = ~w5874 & ~w7227;
assign w7057 = (w12578 & w12917) | (w12578 & w17636) | (w12917 & w17636);
assign w7058 = ~w8055 & ~w8528;
assign w7059 = ~w5841 & ~w8155;
assign w7060 = ~w15888 & ~w6548;
assign w7061 = w3104 & w194;
assign w7062 = w7020 & ~w295;
assign w7063 = ~w18529 & ~w14857;
assign w7064 = ~w7806 & ~w5348;
assign w7065 = ~w10749 & ~w15454;
assign w7066 = ~w2135 & ~w5254;
assign w7067 = w14381 & ~w9209;
assign w7068 = w4169 & w11837;
assign w7069 = w83 & ~w12118;
assign w7070 = w16112 & ~w18215;
assign w7071 = w9538 & ~w17380;
assign w7072 = ~w13914 & ~w12499;
assign w7073 = ~w14894 & ~w9013;
assign w7074 = a_10 & a_57;
assign w7075 = (~w11641 & ~w17967) | (~w11641 & w8291) | (~w17967 & w8291);
assign w7076 = ~w6398 & ~w14852;
assign w7077 = ~w14351 & ~w2501;
assign w7078 = ~w16799 & ~w17615;
assign w7079 = ~w4764 & ~w15783;
assign w7080 = ~w566 & ~w15455;
assign w7081 = w3208 & ~w2300;
assign w7082 = ~w4801 & ~w3783;
assign w7083 = ~w514 & ~w16732;
assign w7084 = ~w4223 & ~w3819;
assign w7085 = w3361 & w3268;
assign w7086 = ~w1838 & ~w7581;
assign w7087 = w16941 & w1079;
assign w7088 = ~w8371 & w15224;
assign w7089 = (~w5952 & w5699) | (~w5952 & w292) | (w5699 & w292);
assign w7090 = ~w4834 & ~w6536;
assign w7091 = ~w8051 & ~w332;
assign w7092 = w2029 & ~w5672;
assign w7093 = ~w2635 & ~w2102;
assign w7094 = w15527 & ~w11668;
assign w7095 = ~w1754 & ~w1053;
assign w7096 = ~w9008 & ~w1486;
assign w7097 = ~w3117 & w10020;
assign w7098 = a_1 & a_10;
assign w7099 = a_14 & a_38;
assign w7100 = w10110 & w7781;
assign w7101 = ~w17361 & ~w12435;
assign w7102 = (w1566 & w14303) | (w1566 & w380) | (w14303 & w380);
assign w7103 = ~w15871 & w17748;
assign w7104 = a_32 & a_33;
assign w7105 = w16675 & ~w12546;
assign w7106 = a_6 & a_57;
assign w7107 = ~w2636 & ~w13955;
assign w7108 = (~w9998 & ~w9809) | (~w9998 & w4643) | (~w9809 & w4643);
assign w7109 = ~w9216 & ~w1418;
assign w7110 = (~w17341 & ~w5956) | (~w17341 & w5658) | (~w5956 & w5658);
assign w7111 = ~w11924 & ~w3513;
assign w7112 = w11140 & ~w10167;
assign w7113 = w13168 & ~w2204;
assign w7114 = ~w11107 & ~w16322;
assign w7115 = (w11515 & w15826) | (w11515 & w972) | (w15826 & w972);
assign w7116 = ~w3461 & ~w8274;
assign w7117 = a_38 & a_43;
assign w7118 = ~w14597 & ~w18776;
assign w7119 = ~w18763 & ~w17291;
assign w7120 = ~w1963 & ~w831;
assign w7121 = w7219 & w11329;
assign w7122 = w14134 & ~w15482;
assign w7123 = ~w14216 & w10960;
assign w7124 = w4830 & w5877;
assign w7125 = ~w16125 & w926;
assign w7126 = w3787 & w3843;
assign w7127 = ~w2530 & ~w17189;
assign w7128 = w6853 & w9372;
assign w7129 = ~w10697 & ~w2254;
assign w7130 = ~w12214 & ~w12801;
assign w7131 = w18558 & ~w3825;
assign w7132 = w9556 & ~w18361;
assign w7133 = ~w994 & w19160;
assign w7134 = a_31 & a_36;
assign w7135 = w7948 & w10674;
assign w7136 = ~w14959 & w7903;
assign w7137 = w9394 & w6668;
assign w7138 = a_2 & a_42;
assign w7139 = ~w12775 & ~w6144;
assign w7140 = ~w9453 & ~w13831;
assign w7141 = ~w15193 & ~w931;
assign w7142 = ~w5016 & ~w4370;
assign w7143 = ~w16430 & ~w9755;
assign w7144 = (w18654 & w11853) | (w18654 & w16403) | (w11853 & w16403);
assign w7145 = ~w16304 & ~w6784;
assign w7146 = ~w3112 & ~w2630;
assign w7147 = (w6938 & w13138) | (w6938 & w13256) | (w13138 & w13256);
assign w7148 = a_30 & a_56;
assign w7149 = ~w9374 & ~w16964;
assign w7150 = ~w7191 & ~w10782;
assign w7151 = ~w16860 & ~w3100;
assign w7152 = ~w171 & ~w12321;
assign w7153 = w11719 & ~w7682;
assign w7154 = a_34 & a_44;
assign w7155 = ~w15305 & ~w8064;
assign w7156 = ~w14981 & ~w18477;
assign w7157 = ~w9067 & w13860;
assign w7158 = ~w7229 & ~w4440;
assign w7159 = ~w3256 & ~w5037;
assign w7160 = a_12 & a_53;
assign w7161 = w10968 & ~w6774;
assign w7162 = ~w12963 & ~w265;
assign w7163 = ~w12514 & ~w9834;
assign w7164 = ~w14431 & ~w3457;
assign w7165 = w17259 & w7340;
assign w7166 = w5011 & ~w10459;
assign w7167 = ~w1572 & ~w8684;
assign w7168 = ~w10322 & ~w14561;
assign w7169 = a_16 & a_52;
assign w7170 = ~w15744 & ~w15677;
assign w7171 = ~w6683 & ~w13939;
assign w7172 = w15610 & ~w9793;
assign w7173 = w13398 & w15944;
assign w7174 = ~w15538 & w17234;
assign w7175 = w16658 & w7859;
assign w7176 = ~w4019 & ~w18390;
assign w7177 = ~w12909 & ~w9906;
assign w7178 = ~w13844 & ~w17112;
assign w7179 = ~w14671 & ~w5375;
assign w7180 = ~w16547 & ~w5312;
assign w7181 = w16923 & w1444;
assign w7182 = w13373 & ~w10442;
assign w7183 = w15099 & w5075;
assign w7184 = ~w4465 & ~w8119;
assign w7185 = ~w2859 & ~w10008;
assign w7186 = ~w9584 & ~w11956;
assign w7187 = w1320 & w9579;
assign w7188 = ~w12904 & w11787;
assign w7189 = ~w16603 & w457;
assign w7190 = ~w17245 & ~w4515;
assign w7191 = w10602 & ~w13029;
assign w7192 = ~w17300 & ~w7988;
assign w7193 = ~w9789 & ~w14867;
assign w7194 = w10844 & ~w4857;
assign w7195 = ~w10842 & w12526;
assign w7196 = ~w1223 & ~w12106;
assign w7197 = ~w1030 & w4738;
assign w7198 = ~w15324 & ~w15173;
assign w7199 = ~w17008 & ~w19109;
assign w7200 = w5915 & w14032;
assign w7201 = ~w10314 & ~w599;
assign w7202 = w2623 & w13657;
assign w7203 = ~w5144 & ~w1051;
assign w7204 = ~w12089 & w12066;
assign w7205 = a_29 & a_49;
assign w7206 = w8371 & ~w15224;
assign w7207 = w10086 & ~w5569;
assign w7208 = w17453 & ~w15026;
assign w7209 = w7249 & ~w1316;
assign w7210 = w14298 & ~w11827;
assign w7211 = w8612 & w18272;
assign w7212 = ~w6330 & ~w4242;
assign w7213 = ~w6889 & ~w4971;
assign w7214 = (~w14557 & ~w13486) | (~w14557 & w4686) | (~w13486 & w4686);
assign w7215 = ~w9493 & ~w12213;
assign w7216 = a_4 & a_30;
assign w7217 = ~w14108 & w12882;
assign w7218 = ~w9403 & w1522;
assign w7219 = a_18 & a_56;
assign w7220 = ~w16429 & ~w14937;
assign w7221 = w5895 & w16311;
assign w7222 = ~w9840 & w4495;
assign w7223 = w11336 & w7355;
assign w7224 = ~w9966 & ~w6684;
assign w7225 = ~w9566 & ~w15257;
assign w7226 = ~w13999 & ~w9288;
assign w7227 = ~w5520 & ~w3706;
assign w7228 = ~w5402 & w3150;
assign w7229 = ~w11910 & w278;
assign w7230 = ~w15242 & ~w6816;
assign w7231 = ~w5814 & w15469;
assign w7232 = ~w1317 & ~w12294;
assign w7233 = (~w11242 & ~w17337) | (~w11242 & w5306) | (~w17337 & w5306);
assign w7234 = ~w10969 & w15275;
assign w7235 = ~w18017 & w14547;
assign w7236 = ~w18434 & ~w17595;
assign w7237 = w3018 & w3192;
assign w7238 = ~w1675 & ~w14029;
assign w7239 = ~w3637 & w16231;
assign w7240 = a_10 & a_12;
assign w7241 = a_1 & a_9;
assign w7242 = a_23 & a_32;
assign w7243 = (~w13481 & w10330) | (~w13481 & w10828) | (w10330 & w10828);
assign w7244 = w2384 & ~w536;
assign w7245 = ~w12641 & w1514;
assign w7246 = w15563 & w17029;
assign w7247 = ~w15604 & ~w7761;
assign w7248 = ~w3458 & ~w16373;
assign w7249 = ~w7087 & ~w1214;
assign w7250 = ~w494 & ~w17869;
assign w7251 = ~w5292 & w3375;
assign w7252 = w11 & ~w15198;
assign w7253 = (w13160 & w10330) | (w13160 & w16334) | (w10330 & w16334);
assign w7254 = a_0 & a_13;
assign w7255 = ~w3021 & ~w10196;
assign w7256 = ~w11619 & ~w18217;
assign w7257 = w11570 & w16131;
assign w7258 = (~w17983 & ~w14604) | (~w17983 & w4321) | (~w14604 & w4321);
assign w7259 = ~w16867 & ~w3081;
assign w7260 = w6392 & w6139;
assign w7261 = w4212 & ~w5032;
assign w7262 = w18417 & w5661;
assign w7263 = ~w16392 & w13789;
assign w7264 = ~w5797 & ~w17293;
assign w7265 = ~w9181 & ~w16986;
assign w7266 = ~w5789 & ~w1089;
assign w7267 = a_17 & a_33;
assign w7268 = ~w9188 & ~w1833;
assign w7269 = ~w2465 & w10669;
assign w7270 = ~w9256 & ~w118;
assign w7271 = ~w13470 & ~w11877;
assign w7272 = ~w18753 & ~w4333;
assign w7273 = (~w11284 & ~w8503) | (~w11284 & w6758) | (~w8503 & w6758);
assign w7274 = w16576 & w16680;
assign w7275 = w14314 & ~w860;
assign w7276 = ~w3193 & ~w12902;
assign w7277 = w519 & w9348;
assign w7278 = w8343 & ~w242;
assign w7279 = w2454 & w11128;
assign w7280 = w5064 & ~w1421;
assign w7281 = ~w2541 & w6125;
assign w7282 = ~w15317 & ~w5794;
assign w7283 = w17480 & ~w14331;
assign w7284 = ~w7044 & ~w15284;
assign w7285 = ~w285 & w12757;
assign w7286 = ~w18417 & ~w5661;
assign w7287 = w14105 & w8808;
assign w7288 = ~w429 & w13580;
assign w7289 = w1671 & ~w1954;
assign w7290 = ~w5387 & w15855;
assign w7291 = (w6087 & w14488) | (w6087 & ~w5108) | (w14488 & ~w5108);
assign w7292 = ~w2108 & w16146;
assign w7293 = a_5 & a_32;
assign w7294 = ~w5011 & w15016;
assign w7295 = a_23 & a_38;
assign w7296 = ~w2694 & ~w14135;
assign w7297 = ~w15485 & ~w4396;
assign w7298 = w1027 & w10483;
assign w7299 = ~w14054 & ~w10913;
assign w7300 = ~w15443 & w10608;
assign w7301 = w16128 & w8642;
assign w7302 = ~w3197 & ~w19071;
assign w7303 = ~w10853 & ~w7487;
assign w7304 = ~w1655 & w5628;
assign w7305 = ~w1118 & w17432;
assign w7306 = a_10 & a_14;
assign w7307 = ~w8900 & ~w9795;
assign w7308 = a_10 & a_60;
assign w7309 = ~w5860 & ~w12915;
assign w7310 = ~w2618 & ~w3251;
assign w7311 = w4992 & ~w14527;
assign w7312 = a_13 & a_43;
assign w7313 = ~w745 & ~w10441;
assign w7314 = ~w10569 & ~w18593;
assign w7315 = (w1225 & w5939) | (w1225 & w14273) | (w5939 & w14273);
assign w7316 = ~w8672 & ~w7343;
assign w7317 = ~w13718 & ~w2353;
assign w7318 = ~w8024 & w18960;
assign w7319 = w14316 & w17333;
assign w7320 = w7066 & w18318;
assign w7321 = ~w14928 & w3017;
assign w7322 = (~w14732 & ~w15760) | (~w14732 & w18298) | (~w15760 & w18298);
assign w7323 = ~w17031 & ~w13253;
assign w7324 = w11009 & ~w12041;
assign w7325 = ~w10225 & w1333;
assign w7326 = w6302 & w12015;
assign w7327 = w4877 & ~w343;
assign w7328 = (w7768 & w4103) | (w7768 & w3322) | (w4103 & w3322);
assign w7329 = ~w11942 & ~w11419;
assign w7330 = w5990 & ~w18358;
assign w7331 = w6640 & w13722;
assign w7332 = ~w5558 & ~w2451;
assign w7333 = ~w8599 & ~w11071;
assign w7334 = ~w18975 & ~w14184;
assign w7335 = ~w9206 & w8422;
assign w7336 = w8166 & ~w18785;
assign w7337 = a_31 & a_55;
assign w7338 = w267 & w9085;
assign w7339 = ~w6689 & ~w8513;
assign w7340 = w4022 & ~w2971;
assign w7341 = (~w3932 & w9337) | (~w3932 & w10582) | (w9337 & w10582);
assign w7342 = ~w16658 & ~w7859;
assign w7343 = ~w8702 & ~w15853;
assign w7344 = w14201 & ~w8390;
assign w7345 = w9651 & ~w1248;
assign w7346 = ~w110 & ~w6369;
assign w7347 = w12667 & ~w14860;
assign w7348 = ~w7509 & ~w9370;
assign w7349 = w11428 & w3125;
assign w7350 = ~w16003 & ~w15295;
assign w7351 = ~w13014 & ~w12103;
assign w7352 = ~w12259 & ~w9992;
assign w7353 = ~w2015 & ~w8510;
assign w7354 = ~w19086 & w7150;
assign w7355 = a_38 & a_48;
assign w7356 = w923 & ~w9001;
assign w7357 = w13513 & ~w5257;
assign w7358 = ~w5677 & ~w16421;
assign w7359 = ~w6820 & ~w15797;
assign w7360 = ~w10245 & w7700;
assign w7361 = ~w6998 & ~w10880;
assign w7362 = ~w3200 & ~w6706;
assign w7363 = ~w14373 & ~w17688;
assign w7364 = ~w19066 & ~w6135;
assign w7365 = a_29 & w2151;
assign w7366 = ~w7610 & w9687;
assign w7367 = (~w539 & ~w6240) | (~w539 & w9319) | (~w6240 & w9319);
assign w7368 = w16498 & ~w16340;
assign w7369 = ~w12393 & ~w2740;
assign w7370 = ~w831 & ~w2167;
assign w7371 = ~w4539 & ~w7672;
assign w7372 = a_9 & a_38;
assign w7373 = ~w13113 & ~w18885;
assign w7374 = ~w13072 & ~w1339;
assign w7375 = w9598 & ~w8305;
assign w7376 = w10450 & ~w3047;
assign w7377 = a_8 & a_33;
assign w7378 = w17211 & w6933;
assign w7379 = ~w8686 & ~w212;
assign w7380 = ~w3871 & ~w9208;
assign w7381 = w10988 & ~w6952;
assign w7382 = w3969 & w8138;
assign w7383 = ~w8704 & ~w8879;
assign w7384 = w17593 & ~w5557;
assign w7385 = w11516 & ~w739;
assign w7386 = ~w8061 & ~w5913;
assign w7387 = ~w3839 & ~w13166;
assign w7388 = ~w13634 & ~w17507;
assign w7389 = a_24 & a_29;
assign w7390 = ~w8953 & ~w15954;
assign w7391 = w15764 & ~w2369;
assign w7392 = ~w17826 & ~w6635;
assign w7393 = ~w12789 & w14906;
assign w7394 = w19082 & w13748;
assign w7395 = ~w16950 & ~w15419;
assign w7396 = ~w1253 & ~w7649;
assign w7397 = w6660 & w5464;
assign w7398 = w12442 & w7003;
assign w7399 = (~w13956 & ~w8249) | (~w13956 & w16094) | (~w8249 & w16094);
assign w7400 = ~w5064 & w1421;
assign w7401 = w17454 & ~w14625;
assign w7402 = ~w15079 & ~w18848;
assign w7403 = w15541 & ~w18205;
assign w7404 = a_9 & a_29;
assign w7405 = ~w17300 & ~w18589;
assign w7406 = ~w18701 & ~w1022;
assign w7407 = ~w6709 & ~w10255;
assign w7408 = ~w18817 & ~w924;
assign w7409 = w6136 & w3235;
assign w7410 = ~w13648 & w2070;
assign w7411 = a_0 & a_37;
assign w7412 = ~w14351 & ~w13525;
assign w7413 = (w17294 & w2254) | (w17294 & w3065) | (w2254 & w3065);
assign w7414 = ~w7897 & ~w7741;
assign w7415 = ~w14113 & ~w10736;
assign w7416 = ~w14026 & ~w3785;
assign w7417 = ~w16936 & ~w4343;
assign w7418 = ~w16199 & ~w18606;
assign w7419 = ~w15297 & ~w12362;
assign w7420 = ~w6853 & w4547;
assign w7421 = w8277 & ~w18500;
assign w7422 = (~w1092 & ~w16662) | (~w1092 & w4214) | (~w16662 & w4214);
assign w7423 = ~w6992 & ~w11386;
assign w7424 = ~w9634 & w358;
assign w7425 = ~w10510 & ~w9124;
assign w7426 = w2710 & ~w7668;
assign w7427 = ~w4311 & ~w10031;
assign w7428 = w5143 & ~w707;
assign w7429 = ~w15450 & ~w9542;
assign w7430 = ~w3326 & ~w18302;
assign w7431 = ~w14591 & w12103;
assign w7432 = ~w15357 & w6910;
assign w7433 = ~w12877 & ~w7578;
assign w7434 = ~w17737 & w18946;
assign w7435 = a_19 & a_62;
assign w7436 = (w9221 & w4779) | (w9221 & w6074) | (w4779 & w6074);
assign w7437 = ~w8350 & ~w9199;
assign w7438 = ~w5072 & ~w11199;
assign w7439 = ~w18197 & ~w8026;
assign w7440 = ~w13224 & ~w13346;
assign w7441 = w16918 & w5939;
assign w7442 = ~w3099 & ~w774;
assign w7443 = a_14 & a_15;
assign w7444 = w7485 & w8343;
assign w7445 = ~w10890 & ~w16137;
assign w7446 = ~w8195 & ~w7552;
assign w7447 = ~w14698 & ~w15037;
assign w7448 = ~w5976 & ~w11361;
assign w7449 = ~w6851 & ~w9055;
assign w7450 = ~w18828 & w5342;
assign w7451 = w3734 & w753;
assign w7452 = ~w5845 & ~w17179;
assign w7453 = w14786 & ~w2395;
assign w7454 = ~w11812 & ~w1338;
assign w7455 = ~w9770 & w1014;
assign w7456 = a_26 & a_63;
assign w7457 = ~w7671 & w17069;
assign w7458 = ~w2174 & ~w12202;
assign w7459 = ~w48 & ~w5624;
assign w7460 = ~w3795 & ~w7135;
assign w7461 = ~w7433 & ~w10831;
assign w7462 = ~w15144 & ~w8628;
assign w7463 = (~w10245 & w16740) | (~w10245 & w15117) | (w16740 & w15117);
assign w7464 = ~w4599 & ~w8901;
assign w7465 = a_14 & a_29;
assign w7466 = w10812 & w9821;
assign w7467 = ~w10804 & w17003;
assign w7468 = w9300 & ~w1642;
assign w7469 = ~w16302 & ~w2315;
assign w7470 = w17629 & ~w8636;
assign w7471 = ~w12683 & ~w6271;
assign w7472 = ~w15437 & ~w17250;
assign w7473 = w6834 & ~w1320;
assign w7474 = w12896 & w1010;
assign w7475 = ~w11947 & ~w14236;
assign w7476 = ~w9405 & w12840;
assign w7477 = w8643 & ~w8854;
assign w7478 = w6095 & w2692;
assign w7479 = ~w8970 & ~w148;
assign w7480 = w2388 & w18898;
assign w7481 = ~w8417 & w16823;
assign w7482 = ~w1839 & w14322;
assign w7483 = w1151 & w7176;
assign w7484 = ~w1273 & ~w10846;
assign w7485 = a_11 & a_42;
assign w7486 = w17145 & w1623;
assign w7487 = w13552 & w1218;
assign w7488 = a_13 & a_62;
assign w7489 = w4385 & w7852;
assign w7490 = ~w12301 & ~w4907;
assign w7491 = w3964 & w10730;
assign w7492 = a_16 & a_40;
assign w7493 = ~w5238 & ~w5777;
assign w7494 = ~w7406 & ~w3982;
assign w7495 = w17204 & ~w18354;
assign w7496 = ~w3775 & w9570;
assign w7497 = (~w17294 & w13082) | (~w17294 & w7584) | (w13082 & w7584);
assign w7498 = w16412 & ~w3628;
assign w7499 = ~w2428 & ~w18902;
assign w7500 = ~w13674 & ~w12112;
assign w7501 = a_9 & a_42;
assign w7502 = ~w6452 & ~w7536;
assign w7503 = ~w1698 & ~w15218;
assign w7504 = ~w3969 & ~w8138;
assign w7505 = ~w320 & w12727;
assign w7506 = ~w18690 & ~w16760;
assign w7507 = w1806 & ~w8846;
assign w7508 = (w9869 & w2769) | (w9869 & w13583) | (w2769 & w13583);
assign w7509 = w7307 & ~w3850;
assign w7510 = a_54 & a_56;
assign w7511 = ~w15303 & ~w6675;
assign w7512 = w6359 & ~w7023;
assign w7513 = w3259 & ~w93;
assign w7514 = w6423 & w5600;
assign w7515 = w8655 & ~w17542;
assign w7516 = ~w8807 & ~w14795;
assign w7517 = ~w3159 & ~w3892;
assign w7518 = w1207 & w1188;
assign w7519 = ~w7381 & w18358;
assign w7520 = w15753 & ~w4675;
assign w7521 = ~w7086 & ~w11864;
assign w7522 = ~w4053 & ~w15964;
assign w7523 = w5217 & w1645;
assign w7524 = ~w18176 & ~w7737;
assign w7525 = ~w3802 & w6768;
assign w7526 = ~w6123 & ~w3136;
assign w7527 = ~w15520 & w446;
assign w7528 = w14617 & ~w8194;
assign w7529 = a_4 & a_55;
assign w7530 = w12509 & ~w11421;
assign w7531 = w17963 & w16782;
assign w7532 = (~w10048 & w17145) | (~w10048 & w5321) | (w17145 & w5321);
assign w7533 = ~w13808 & ~w4289;
assign w7534 = ~w7707 & w13811;
assign w7535 = w867 & w19020;
assign w7536 = ~w3078 & w4969;
assign w7537 = ~w8188 & ~w18791;
assign w7538 = ~w11814 & ~w8492;
assign w7539 = w11051 & w18923;
assign w7540 = ~w13982 & ~w4580;
assign w7541 = w17656 & ~w8676;
assign w7542 = (~w5417 & ~w2142) | (~w5417 & w7975) | (~w2142 & w7975);
assign w7543 = w4114 & w9454;
assign w7544 = (~w13059 & ~w2140) | (~w13059 & w8242) | (~w2140 & w8242);
assign w7545 = a_5 & a_36;
assign w7546 = (w15850 & w2769) | (w15850 & w643) | (w2769 & w643);
assign w7547 = ~w12553 & ~w9436;
assign w7548 = ~w7483 & ~w1040;
assign w7549 = ~w8407 & ~w6544;
assign w7550 = a_32 & a_63;
assign w7551 = a_15 & a_28;
assign w7552 = w3537 & w10448;
assign w7553 = a_46 & a_49;
assign w7554 = (~w1818 & w944) | (~w1818 & w6648) | (w944 & w6648);
assign w7555 = w11934 & w10903;
assign w7556 = a_16 & a_41;
assign w7557 = ~w12918 & ~w17832;
assign w7558 = w16727 & w7119;
assign w7559 = ~w1943 & ~w8785;
assign w7560 = ~w19081 & ~w18149;
assign w7561 = ~w6428 & ~w6261;
assign w7562 = (~w16679 & ~w14218) | (~w16679 & w9107) | (~w14218 & w9107);
assign w7563 = ~w17419 & ~w10719;
assign w7564 = a_15 & a_63;
assign w7565 = ~w11321 & ~w3901;
assign w7566 = ~w3792 & ~w10035;
assign w7567 = ~w4939 & ~w8657;
assign w7568 = ~w12029 & ~w11018;
assign w7569 = ~w3702 & w2321;
assign w7570 = ~w18118 & ~w12921;
assign w7571 = ~w13220 & w7268;
assign w7572 = ~w2379 & ~w14618;
assign w7573 = ~w10984 & w10454;
assign w7574 = w18579 & w5442;
assign w7575 = ~w8807 & ~w10284;
assign w7576 = ~w14959 & ~w6988;
assign w7577 = w9371 & ~w16525;
assign w7578 = a_3 & a_6;
assign w7579 = a_32 & a_36;
assign w7580 = w3099 & ~w11163;
assign w7581 = w6364 & w15056;
assign w7582 = w9873 & ~w17626;
assign w7583 = ~w14949 & ~w15710;
assign w7584 = ~w2254 & w13773;
assign w7585 = w7844 & ~w6604;
assign w7586 = (~w18315 & ~w10336) | (~w18315 & w15413) | (~w10336 & w15413);
assign w7587 = ~w1826 & ~w7677;
assign w7588 = ~w9261 & ~w12869;
assign w7589 = ~w9670 & ~w570;
assign w7590 = ~w13964 & ~w5751;
assign w7591 = ~w15764 & w11495;
assign w7592 = (w1906 & w16375) | (w1906 & w11908) | (w16375 & w11908);
assign w7593 = a_3 & a_28;
assign w7594 = w13254 & w5108;
assign w7595 = ~w10174 & ~w14630;
assign w7596 = (w10961 & w10330) | (w10961 & w2803) | (w10330 & w2803);
assign w7597 = (~w152 & w6300) | (~w152 & w5409) | (w6300 & w5409);
assign w7598 = ~w6987 & w14001;
assign w7599 = ~w18327 & w6565;
assign w7600 = ~w14569 & w7276;
assign w7601 = a_20 & a_28;
assign w7602 = ~w9538 & w17380;
assign w7603 = ~w8815 & ~w13412;
assign w7604 = ~w1977 & ~w1621;
assign w7605 = ~w10058 & ~w10947;
assign w7606 = ~w12419 & w9025;
assign w7607 = ~w16061 & ~w12632;
assign w7608 = w12456 & w4651;
assign w7609 = w4633 & ~w3522;
assign w7610 = (w18843 & w8052) | (w18843 & w6366) | (w8052 & w6366);
assign w7611 = w8957 & w5101;
assign w7612 = ~w18980 & w11689;
assign w7613 = ~w9501 & ~w7762;
assign w7614 = a_22 & a_24;
assign w7615 = w2206 & w2835;
assign w7616 = w16761 & w13625;
assign w7617 = (~w11471 & w8809) | (~w11471 & w400) | (w8809 & w400);
assign w7618 = w2543 & ~w15628;
assign w7619 = ~w16727 & ~w14483;
assign w7620 = ~w184 & ~w17192;
assign w7621 = (~w5277 & ~w909) | (~w5277 & w15222) | (~w909 & w15222);
assign w7622 = ~w10311 & ~w2804;
assign w7623 = ~w2577 & w990;
assign w7624 = ~w1063 & ~w18691;
assign w7625 = ~w18737 & w10564;
assign w7626 = ~a_30 & w12128;
assign w7627 = ~w18596 & ~w1652;
assign w7628 = ~w9303 & ~w15071;
assign w7629 = ~w844 & w18331;
assign w7630 = ~w9034 & ~w15604;
assign w7631 = ~w9027 & ~w7556;
assign w7632 = ~w8174 & ~w7429;
assign w7633 = w7981 & w2083;
assign w7634 = ~w10604 & ~w16031;
assign w7635 = ~w13970 & w17301;
assign w7636 = w12037 & ~w4597;
assign w7637 = w1144 & ~w4993;
assign w7638 = ~w1976 & ~w16449;
assign w7639 = ~w1946 & ~w2972;
assign w7640 = ~w4147 & w10024;
assign w7641 = ~w13384 & ~w8356;
assign w7642 = w5424 & w2320;
assign w7643 = w12180 & ~w13091;
assign w7644 = w8041 & w1734;
assign w7645 = w4088 & w6192;
assign w7646 = w15510 & ~w16961;
assign w7647 = ~w17116 & w17023;
assign w7648 = w18629 & ~w3160;
assign w7649 = w1994 & w13714;
assign w7650 = w6875 & w17979;
assign w7651 = ~w12274 & w8585;
assign w7652 = ~w15749 & w14456;
assign w7653 = ~a_12 & ~w15843;
assign w7654 = ~w6685 & ~w17312;
assign w7655 = w9292 & ~w16395;
assign w7656 = (~w381 & ~w15674) | (~w381 & w16294) | (~w15674 & w16294);
assign w7657 = (~w3875 & ~w5434) | (~w3875 & w12364) | (~w5434 & w12364);
assign w7658 = ~w12038 & ~w1589;
assign w7659 = ~w18806 & ~w2525;
assign w7660 = w53 & w7977;
assign w7661 = a_36 & a_50;
assign w7662 = ~w17063 & ~w10407;
assign w7663 = a_26 & a_50;
assign w7664 = ~w15057 & ~w5472;
assign w7665 = w13604 & ~w6132;
assign w7666 = ~w17470 & ~w9011;
assign w7667 = ~w5398 & w6547;
assign w7668 = ~w11957 & ~w9757;
assign w7669 = ~w4412 & ~w9486;
assign w7670 = w12654 & ~w13436;
assign w7671 = ~w4441 & ~w3743;
assign w7672 = w10522 & w10835;
assign w7673 = ~w4002 & w4337;
assign w7674 = w15227 & ~w4777;
assign w7675 = ~w6081 & w12836;
assign w7676 = w10577 & w1533;
assign w7677 = ~w4079 & ~w130;
assign w7678 = w11119 & w4254;
assign w7679 = w15276 & ~w12216;
assign w7680 = ~w8500 & ~w13944;
assign w7681 = w16439 & ~w120;
assign w7682 = ~w3849 & ~w10054;
assign w7683 = ~w2554 & ~w11261;
assign w7684 = w12122 & w12622;
assign w7685 = w5102 & ~w10362;
assign w7686 = ~w7129 & w12400;
assign w7687 = (w3649 & w8580) | (w3649 & w6254) | (w8580 & w6254);
assign w7688 = (~w14997 & ~w14620) | (~w14997 & w3358) | (~w14620 & w3358);
assign w7689 = ~w4863 & ~w10435;
assign w7690 = w6969 & ~w19123;
assign w7691 = a_35 & a_45;
assign w7692 = ~w16859 & ~w17283;
assign w7693 = ~w6853 & w14256;
assign w7694 = w12465 & ~w11258;
assign w7695 = ~w13763 & ~w11919;
assign w7696 = ~w3277 & w7796;
assign w7697 = w11275 & ~w1465;
assign w7698 = w1747 & w17013;
assign w7699 = ~w4657 & ~w13782;
assign w7700 = ~w8436 & ~w17134;
assign w7701 = w17396 & w17103;
assign w7702 = ~w627 & ~w14754;
assign w7703 = a_13 & a_32;
assign w7704 = (~w7434 & ~w9889) | (~w7434 & w11375) | (~w9889 & w11375);
assign w7705 = a_15 & a_58;
assign w7706 = ~w1968 & ~w5411;
assign w7707 = ~w2322 & ~w17251;
assign w7708 = ~w10873 & ~w3624;
assign w7709 = ~w5461 & ~w3521;
assign w7710 = ~w6566 & w18986;
assign w7711 = (w11174 & w2769) | (w11174 & w15736) | (w2769 & w15736);
assign w7712 = w15116 & ~w12189;
assign w7713 = ~w14980 & w11585;
assign w7714 = (w15569 & w3042) | (w15569 & w15536) | (w3042 & w15536);
assign w7715 = ~w18812 & ~w5731;
assign w7716 = ~w7766 & ~w14137;
assign w7717 = w3250 & w13142;
assign w7718 = ~w3872 & ~w6623;
assign w7719 = ~w9146 & ~w2708;
assign w7720 = ~w10901 & ~w1760;
assign w7721 = ~w7278 & ~w10746;
assign w7722 = ~w11437 & ~w13032;
assign w7723 = w12971 & ~w6224;
assign w7724 = w15768 & w6767;
assign w7725 = ~w3029 & ~w8814;
assign w7726 = ~w12863 & ~w18233;
assign w7727 = (~w3695 & w12904) | (~w3695 & w14163) | (w12904 & w14163);
assign w7728 = w9729 & ~w3025;
assign w7729 = w3641 & w1524;
assign w7730 = ~w3489 & w6753;
assign w7731 = w5180 & w14674;
assign w7732 = a_8 & a_42;
assign w7733 = ~w849 & ~w19024;
assign w7734 = ~w13909 & w4554;
assign w7735 = ~w6919 & ~w18967;
assign w7736 = ~w2735 & ~w2946;
assign w7737 = ~w16047 & ~w354;
assign w7738 = ~w8326 & ~w9041;
assign w7739 = ~w10749 & ~w6879;
assign w7740 = w6356 & ~w2537;
assign w7741 = ~w8269 & ~w12811;
assign w7742 = ~w2954 & w3595;
assign w7743 = w15704 & ~w14666;
assign w7744 = ~w5378 & w10576;
assign w7745 = ~w7251 & ~w4634;
assign w7746 = a_17 & a_57;
assign w7747 = a_9 & a_50;
assign w7748 = ~w10340 & ~w11708;
assign w7749 = ~w15718 & ~w5649;
assign w7750 = ~w8039 & w18719;
assign w7751 = ~w10660 & ~w8431;
assign w7752 = ~w5542 & ~w12373;
assign w7753 = ~w14168 & ~w6357;
assign w7754 = (~w4237 & ~w14875) | (~w4237 & w10760) | (~w14875 & w10760);
assign w7755 = ~w18437 & ~w16476;
assign w7756 = a_10 & a_35;
assign w7757 = w13919 & w16771;
assign w7758 = ~w10504 & ~w6024;
assign w7759 = (~w8436 & ~w7700) | (~w8436 & w8354) | (~w7700 & w8354);
assign w7760 = ~w15183 & w10182;
assign w7761 = ~w8592 & ~w1431;
assign w7762 = ~w6707 & ~w2613;
assign w7763 = w19063 & w664;
assign w7764 = a_14 & a_34;
assign w7765 = a_38 & a_41;
assign w7766 = w6550 & w5917;
assign w7767 = a_4 & a_41;
assign w7768 = ~w18747 & w8860;
assign w7769 = ~w5371 & ~w15652;
assign w7770 = ~w8899 & w12931;
assign w7771 = w9692 & ~w894;
assign w7772 = (w7409 & ~w16896) | (w7409 & w2595) | (~w16896 & w2595);
assign w7773 = ~w920 & ~w276;
assign w7774 = ~w2337 & ~w15779;
assign w7775 = ~w7322 & ~w10993;
assign w7776 = (~w5724 & w3182) | (~w5724 & w4442) | (w3182 & w4442);
assign w7777 = ~w957 & ~w2028;
assign w7778 = (w16322 & w6601) | (w16322 & w13280) | (w6601 & w13280);
assign w7779 = ~w17692 & ~w5471;
assign w7780 = ~w4312 & w1386;
assign w7781 = ~w10711 & ~w1637;
assign w7782 = ~w9165 & ~w15387;
assign w7783 = ~w6057 & w8613;
assign w7784 = w6373 & w5145;
assign w7785 = w4548 & ~w19138;
assign w7786 = w12271 & w14473;
assign w7787 = ~w13003 & w18979;
assign w7788 = w13028 & ~w4360;
assign w7789 = w10400 & ~w13344;
assign w7790 = ~w4379 & ~w8653;
assign w7791 = ~w16675 & w12546;
assign w7792 = ~w1923 & w6134;
assign w7793 = ~w16248 & w17696;
assign w7794 = w11150 & ~w15181;
assign w7795 = ~w10108 & ~w15102;
assign w7796 = (~w282 & ~w15793) | (~w282 & w8932) | (~w15793 & w8932);
assign w7797 = ~w586 & ~w14013;
assign w7798 = ~w13332 & w2321;
assign w7799 = w7538 & ~w18172;
assign w7800 = ~w18232 & ~w12061;
assign w7801 = a_41 & a_47;
assign w7802 = w14069 & w15762;
assign w7803 = ~w11800 & ~w17350;
assign w7804 = ~w15629 & ~w17319;
assign w7805 = ~w8052 & w17833;
assign w7806 = ~w12284 & ~w11828;
assign w7807 = ~w16358 & ~w9285;
assign w7808 = w13689 & w3;
assign w7809 = ~w7019 & w17381;
assign w7810 = w11205 & ~w1439;
assign w7811 = w8485 & w13479;
assign w7812 = ~w6417 & ~w12768;
assign w7813 = ~w5158 & ~w2330;
assign w7814 = ~w12826 & ~w18004;
assign w7815 = ~w16254 & ~w313;
assign w7816 = ~w11393 & ~w6276;
assign w7817 = a_10 & a_38;
assign w7818 = a_12 & a_27;
assign w7819 = ~w16767 & w3797;
assign w7820 = ~w13306 & w13670;
assign w7821 = w12935 & ~w16093;
assign w7822 = ~w12885 & ~w16608;
assign w7823 = w6495 & w5921;
assign w7824 = ~w2747 & ~w14224;
assign w7825 = ~w18170 & ~w288;
assign w7826 = (w7604 & ~w2870) | (w7604 & w9636) | (~w2870 & w9636);
assign w7827 = ~w1313 & w19139;
assign w7828 = ~w16637 & w554;
assign w7829 = ~w8307 & ~w7731;
assign w7830 = ~w13364 & ~w1251;
assign w7831 = w7550 & w18814;
assign w7832 = w16405 & w18467;
assign w7833 = w2911 & ~w3837;
assign w7834 = ~w16621 & ~w17662;
assign w7835 = ~w7895 & ~w17934;
assign w7836 = w2734 & ~w19026;
assign w7837 = ~w15622 & w16361;
assign w7838 = w4793 & w4838;
assign w7839 = w3921 & ~w6727;
assign w7840 = w8648 & ~w13192;
assign w7841 = ~w18537 & ~w9341;
assign w7842 = w16493 & ~w832;
assign w7843 = w10220 & ~w16286;
assign w7844 = a_23 & a_36;
assign w7845 = ~w14360 & ~w15401;
assign w7846 = ~w14452 & w19161;
assign w7847 = ~w17095 & ~w10143;
assign w7848 = w9799 & ~w11689;
assign w7849 = ~w10983 & ~w3633;
assign w7850 = ~w3341 & ~w805;
assign w7851 = ~w8012 & w8207;
assign w7852 = ~w4330 & ~w2574;
assign w7853 = w4590 & ~w8554;
assign w7854 = ~w12406 & w2652;
assign w7855 = ~w10147 & ~w2713;
assign w7856 = w8065 & w15597;
assign w7857 = ~w10333 & ~w6870;
assign w7858 = a_1 & a_37;
assign w7859 = ~w16355 & ~w3844;
assign w7860 = a_21 & a_33;
assign w7861 = ~w18682 & w9974;
assign w7862 = w1250 & ~w10816;
assign w7863 = ~w1903 & w11449;
assign w7864 = w403 & ~w1956;
assign w7865 = ~w422 & ~w16821;
assign w7866 = (~w7102 & w8497) | (~w7102 & w15795) | (w8497 & w15795);
assign w7867 = ~w12365 & ~w6714;
assign w7868 = ~w17915 & ~w4203;
assign w7869 = a_5 & a_57;
assign w7870 = ~w4867 & ~w3573;
assign w7871 = ~w16625 & ~w14313;
assign w7872 = ~w3882 & ~w16092;
assign w7873 = ~w8286 & w10790;
assign w7874 = ~w3048 & w2477;
assign w7875 = a_41 & a_54;
assign w7876 = (w8169 & ~w1320) | (w8169 & w14021) | (~w1320 & w14021);
assign w7877 = ~w6862 & ~w4004;
assign w7878 = w13668 & w3645;
assign w7879 = ~w12278 & w11605;
assign w7880 = w5283 & w2830;
assign w7881 = ~w6781 & ~w10076;
assign w7882 = w9824 & ~w10279;
assign w7883 = ~w717 & w7213;
assign w7884 = ~w3448 & ~w13516;
assign w7885 = (w7341 & w15133) | (w7341 & w5071) | (w15133 & w5071);
assign w7886 = ~w4312 & w5882;
assign w7887 = ~w7158 & ~w8091;
assign w7888 = ~w13494 & ~w12535;
assign w7889 = w18551 & ~w12370;
assign w7890 = ~w1449 & w18374;
assign w7891 = a_0 & a_36;
assign w7892 = w15270 & w1788;
assign w7893 = ~w16406 & w15097;
assign w7894 = w18442 & ~w18109;
assign w7895 = ~w947 & w12023;
assign w7896 = ~w9420 & w2206;
assign w7897 = ~w16523 & w6602;
assign w7898 = ~w15116 & w12189;
assign w7899 = a_29 & a_59;
assign w7900 = ~w18034 & ~w17408;
assign w7901 = w12390 & ~w15623;
assign w7902 = ~w14182 & ~w5603;
assign w7903 = ~w7462 & ~w19118;
assign w7904 = w15510 & ~w16350;
assign w7905 = ~w13082 & w3446;
assign w7906 = a_17 & a_42;
assign w7907 = ~w12421 & ~w12996;
assign w7908 = ~w14353 & ~w507;
assign w7909 = w13921 & w16530;
assign w7910 = a_26 & a_41;
assign w7911 = w13889 & w10360;
assign w7912 = ~w18372 & ~w15258;
assign w7913 = ~w2648 & ~w17275;
assign w7914 = w17116 & ~w17270;
assign w7915 = ~w12677 & ~w707;
assign w7916 = w2177 & w8458;
assign w7917 = ~w18212 & w18683;
assign w7918 = w10298 & ~w6375;
assign w7919 = a_52 & a_61;
assign w7920 = w18128 & w19162;
assign w7921 = ~w2530 & ~w18973;
assign w7922 = ~w4168 & ~w7367;
assign w7923 = w320 & ~w12727;
assign w7924 = ~w6491 & w10558;
assign w7925 = a_7 & a_51;
assign w7926 = ~w14064 & ~w11219;
assign w7927 = w13082 & ~w3908;
assign w7928 = ~w18129 & ~w6202;
assign w7929 = ~w8826 & ~w14453;
assign w7930 = ~w16505 & w14776;
assign w7931 = ~w14299 & ~w7891;
assign w7932 = a_23 & a_60;
assign w7933 = ~w17767 & ~w9852;
assign w7934 = ~w16240 & ~w17220;
assign w7935 = ~w7774 & ~w16965;
assign w7936 = ~w6316 & ~w5855;
assign w7937 = w5014 & w18859;
assign w7938 = ~w16357 & w15063;
assign w7939 = w14617 & w16546;
assign w7940 = w14286 & ~w4906;
assign w7941 = a_0 & a_31;
assign w7942 = w16250 & w10455;
assign w7943 = ~w5108 & w4043;
assign w7944 = ~w3907 & ~w13652;
assign w7945 = ~w12864 & w5958;
assign w7946 = (~w15150 & w8143) | (~w15150 & w2351) | (w8143 & w2351);
assign w7947 = ~w15714 & ~w17458;
assign w7948 = a_4 & a_53;
assign w7949 = ~w10902 & ~w7655;
assign w7950 = a_40 & w13653;
assign w7951 = ~w6793 & ~w12323;
assign w7952 = ~w5507 & ~w4673;
assign w7953 = ~w16809 & ~w6507;
assign w7954 = ~w11499 & w6357;
assign w7955 = ~w8877 & w15097;
assign w7956 = a_51 & a_52;
assign w7957 = ~w18944 & ~w8730;
assign w7958 = ~w8816 & ~w9002;
assign w7959 = ~w10085 & ~w3254;
assign w7960 = w16406 & ~w15097;
assign w7961 = ~w7500 & ~w6348;
assign w7962 = ~w16579 & ~w14635;
assign w7963 = ~w17438 & ~w4087;
assign w7964 = ~w17418 & ~w3903;
assign w7965 = ~w6157 & ~w14370;
assign w7966 = w10675 & w11850;
assign w7967 = w11515 & w11406;
assign w7968 = w16070 & w7683;
assign w7969 = (w7102 & w8485) | (w7102 & w6946) | (w8485 & w6946);
assign w7970 = ~w16006 & ~w8652;
assign w7971 = ~w1826 & ~w17463;
assign w7972 = ~w10618 & ~w5733;
assign w7973 = ~w4181 & ~w16049;
assign w7974 = w3463 & w1697;
assign w7975 = w17874 & ~w5417;
assign w7976 = ~w14247 & ~w5954;
assign w7977 = (~w14114 & ~w16135) | (~w14114 & w423) | (~w16135 & w423);
assign w7978 = ~w13717 & ~w3402;
assign w7979 = ~w6610 & ~w747;
assign w7980 = (~w16896 & w2709) | (~w16896 & w15861) | (w2709 & w15861);
assign w7981 = a_16 & a_59;
assign w7982 = a_17 & a_30;
assign w7983 = ~w5007 & ~w12502;
assign w7984 = w18910 & w12549;
assign w7985 = ~w13453 & ~w12197;
assign w7986 = w16769 & ~w12422;
assign w7987 = w18127 & ~w10212;
assign w7988 = ~w13879 & w10784;
assign w7989 = w15677 & ~w10149;
assign w7990 = w2968 & ~w6931;
assign w7991 = a_25 & a_29;
assign w7992 = (~w8792 & ~w6527) | (~w8792 & w1929) | (~w6527 & w1929);
assign w7993 = ~w4211 & ~w18880;
assign w7994 = ~w10943 & ~w18643;
assign w7995 = ~w5385 & ~w3698;
assign w7996 = ~w15294 & ~w10696;
assign w7997 = ~w1969 & ~w5458;
assign w7998 = ~w19082 & ~w13748;
assign w7999 = ~w17593 & w13593;
assign w8000 = a_39 & a_57;
assign w8001 = ~w14998 & ~w1606;
assign w8002 = w1054 & w18596;
assign w8003 = ~w7833 & ~w12592;
assign w8004 = ~w1403 & ~w6157;
assign w8005 = ~w15761 & ~w17075;
assign w8006 = (~w2875 & ~w17546) | (~w2875 & w3593) | (~w17546 & w3593);
assign w8007 = ~w10049 & w3131;
assign w8008 = (w7102 & w11050) | (w7102 & w13244) | (w11050 & w13244);
assign w8009 = ~w16654 & ~w15181;
assign w8010 = ~w16737 & ~w451;
assign w8011 = w551 & ~w9210;
assign w8012 = (~w6645 & ~w8299) | (~w6645 & w14399) | (~w8299 & w14399);
assign w8013 = ~w8443 & ~w12160;
assign w8014 = ~w6878 & ~w17229;
assign w8015 = ~w5086 & ~w15700;
assign w8016 = w562 & ~w17562;
assign w8017 = ~w5928 & ~w15493;
assign w8018 = w5425 & ~w6296;
assign w8019 = w8343 & w16186;
assign w8020 = w11726 & w15898;
assign w8021 = a_9 & a_10;
assign w8022 = w13333 & w11203;
assign w8023 = ~w9530 & ~w9523;
assign w8024 = ~w5213 & ~w16647;
assign w8025 = w17643 & ~w8251;
assign w8026 = a_0 & a_9;
assign w8027 = w10854 & ~w569;
assign w8028 = w2666 & ~w17329;
assign w8029 = a_40 & a_42;
assign w8030 = ~w2110 & ~w18799;
assign w8031 = ~w1980 & w1255;
assign w8032 = w19114 & w614;
assign w8033 = ~w7219 & ~w11329;
assign w8034 = a_3 & a_57;
assign w8035 = ~w13227 & w6250;
assign w8036 = a_28 & a_39;
assign w8037 = w3547 & w3883;
assign w8038 = ~w16120 & ~w13594;
assign w8039 = a_7 & a_53;
assign w8040 = w612 & w7746;
assign w8041 = ~w18504 & ~w6737;
assign w8042 = w7919 & w1016;
assign w8043 = ~w859 & ~w18822;
assign w8044 = a_25 & a_54;
assign w8045 = (~w7341 & w18441) | (~w7341 & w15922) | (w18441 & w15922);
assign w8046 = (~w13280 & w5749) | (~w13280 & w12770) | (w5749 & w12770);
assign w8047 = w12994 & w7720;
assign w8048 = ~w13957 & ~w9527;
assign w8049 = (~w16234 & w7329) | (~w16234 & w13862) | (w7329 & w13862);
assign w8050 = a_26 & w6141;
assign w8051 = w14210 & ~w7779;
assign w8052 = (~w19035 & ~w9703) | (~w19035 & w6022) | (~w9703 & w6022);
assign w8053 = w2093 & ~w13241;
assign w8054 = (~w16663 & ~w15199) | (~w16663 & w9997) | (~w15199 & w9997);
assign w8055 = ~w7152 & w16271;
assign w8056 = ~w9843 & ~w19060;
assign w8057 = w14755 & ~w1693;
assign w8058 = ~w18457 & ~w9360;
assign w8059 = w15384 & ~w2291;
assign w8060 = w12008 & ~w10239;
assign w8061 = w15753 & ~w9114;
assign w8062 = w18917 & w18550;
assign w8063 = a_22 & a_53;
assign w8064 = w2976 & ~w5488;
assign w8065 = ~w12309 & ~w10505;
assign w8066 = w3502 & w5324;
assign w8067 = ~w11522 & ~w18097;
assign w8068 = ~w3339 & ~w16114;
assign w8069 = a_2 & a_5;
assign w8070 = w12776 & w12007;
assign w8071 = ~w4053 & w17961;
assign w8072 = ~w18376 & ~w8557;
assign w8073 = ~w8958 & ~w14970;
assign w8074 = ~w3514 & ~w4221;
assign w8075 = ~w16162 & ~w14450;
assign w8076 = ~w17248 & w16739;
assign w8077 = (~w2769 & w14412) | (~w2769 & w18961) | (w14412 & w18961);
assign w8078 = ~w15706 & ~w18811;
assign w8079 = w13158 & ~w10854;
assign w8080 = w18666 & w11530;
assign w8081 = a_24 & a_52;
assign w8082 = w9704 & w3127;
assign w8083 = ~w14035 & ~w3198;
assign w8084 = w7230 & ~w6661;
assign w8085 = w14140 & w6686;
assign w8086 = ~w17231 & w16683;
assign w8087 = w7416 & ~w7721;
assign w8088 = ~w1542 & ~w1269;
assign w8089 = (~w12953 & ~w13361) | (~w12953 & w3046) | (~w13361 & w3046);
assign w8090 = ~w14582 & ~w10497;
assign w8091 = ~w16274 & ~w6194;
assign w8092 = ~w16316 & ~w15539;
assign w8093 = ~w16554 & ~w6618;
assign w8094 = w4472 & w18414;
assign w8095 = ~w276 & ~w878;
assign w8096 = ~w17336 & ~w10018;
assign w8097 = ~w14705 & w4941;
assign w8098 = ~w1687 & ~w2402;
assign w8099 = ~w18841 & ~w18698;
assign w8100 = a_2 & a_16;
assign w8101 = ~w4560 & ~w17490;
assign w8102 = ~w13625 & ~w11436;
assign w8103 = ~w14871 & ~w1689;
assign w8104 = ~w11924 & w12998;
assign w8105 = ~w10568 & ~w18557;
assign w8106 = w11434 & w165;
assign w8107 = w14365 & ~w13811;
assign w8108 = w15095 & w6963;
assign w8109 = ~w4304 & ~w3529;
assign w8110 = ~w12356 & w13401;
assign w8111 = ~w16216 & ~w6882;
assign w8112 = ~w15397 & w10038;
assign w8113 = ~w18209 & w15342;
assign w8114 = ~w9048 & w10009;
assign w8115 = ~w17395 & w7225;
assign w8116 = ~w15373 & ~w7068;
assign w8117 = w6520 & w9450;
assign w8118 = w14678 & ~w5061;
assign w8119 = ~w8685 & w11612;
assign w8120 = a_29 & a_51;
assign w8121 = ~w5591 & w18666;
assign w8122 = (w12595 & w14429) | (w12595 & w8836) | (w14429 & w8836);
assign w8123 = (w9549 & w8747) | (w9549 & w18410) | (w8747 & w18410);
assign w8124 = ~w2849 & w4991;
assign w8125 = ~w15452 & ~w3548;
assign w8126 = ~w4137 & ~w11320;
assign w8127 = (~w16082 & ~w10137) | (~w16082 & w13409) | (~w10137 & w13409);
assign w8128 = ~w11587 & ~w17319;
assign w8129 = w15152 & w14846;
assign w8130 = w18578 & ~w11794;
assign w8131 = ~w3433 & ~w5089;
assign w8132 = w563 & w9422;
assign w8133 = ~w534 & w17968;
assign w8134 = ~w15664 & ~w17051;
assign w8135 = a_62 & ~w10389;
assign w8136 = ~w712 & ~w16548;
assign w8137 = ~w3058 & ~w1264;
assign w8138 = ~w12979 & ~w856;
assign w8139 = w14041 & ~w19122;
assign w8140 = w11792 & ~w3555;
assign w8141 = ~w5452 & w17904;
assign w8142 = ~w5484 & ~w5546;
assign w8143 = (~w296 & ~w12992) | (~w296 & w2230) | (~w12992 & w2230);
assign w8144 = w16493 & ~w631;
assign w8145 = w16640 & ~w2811;
assign w8146 = a_29 & a_47;
assign w8147 = w8176 & ~w16237;
assign w8148 = ~w10992 & ~w11627;
assign w8149 = w2970 & ~w13226;
assign w8150 = ~w14250 & ~w3356;
assign w8151 = ~w17605 & ~w14307;
assign w8152 = ~w11782 & w12488;
assign w8153 = w4328 & ~w3071;
assign w8154 = (~w8636 & w11391) | (~w8636 & w17629) | (w11391 & w17629);
assign w8155 = w15562 & ~w6769;
assign w8156 = a_11 & a_13;
assign w8157 = ~w6777 & ~w5627;
assign w8158 = ~w18276 & ~w4893;
assign w8159 = ~w16846 & ~w11724;
assign w8160 = ~w5313 & ~w719;
assign w8161 = ~w2255 & ~w11617;
assign w8162 = w18990 & ~w12699;
assign w8163 = ~w12940 & w18903;
assign w8164 = ~w186 & ~w7717;
assign w8165 = (~w16323 & ~w9901) | (~w16323 & w9881) | (~w9901 & w9881);
assign w8166 = ~w14018 & ~w5188;
assign w8167 = w12987 & ~w7499;
assign w8168 = ~w14365 & w13811;
assign w8169 = ~w17690 & ~w8992;
assign w8170 = ~w8302 & w6724;
assign w8171 = ~w10436 & ~w4060;
assign w8172 = w8012 & ~w8207;
assign w8173 = a_44 & a_45;
assign w8174 = ~w4854 & ~w18676;
assign w8175 = a_16 & a_21;
assign w8176 = ~w17205 & ~w10726;
assign w8177 = ~w7355 & ~w716;
assign w8178 = ~w412 & w12801;
assign w8179 = ~w9986 & ~w15432;
assign w8180 = w2104 & ~w16881;
assign w8181 = ~w3674 & ~w8931;
assign w8182 = ~w3257 & ~w17450;
assign w8183 = ~w4145 & ~w15916;
assign w8184 = w5849 & ~w5897;
assign w8185 = ~w1583 & ~w2434;
assign w8186 = w16313 & ~w12211;
assign w8187 = ~w16221 & ~w4118;
assign w8188 = w4135 & w15100;
assign w8189 = ~w17441 & ~w17569;
assign w8190 = a_6 & a_37;
assign w8191 = w14862 & w910;
assign w8192 = (w2249 & w12128) | (w2249 & w11563) | (w12128 & w11563);
assign w8193 = (w12255 & w11948) | (w12255 & w4986) | (w11948 & w4986);
assign w8194 = ~w14408 & ~w6581;
assign w8195 = ~w3537 & ~w10448;
assign w8196 = w8375 & w2821;
assign w8197 = w4558 & ~w7479;
assign w8198 = (~w15195 & ~w10254) | (~w15195 & w11358) | (~w10254 & w11358);
assign w8199 = ~w9746 & ~w6378;
assign w8200 = ~w3176 & ~w17009;
assign w8201 = a_14 & a_49;
assign w8202 = ~w11874 & ~w15455;
assign w8203 = w9 & ~w10186;
assign w8204 = w10150 & w2469;
assign w8205 = ~w9235 & ~w9653;
assign w8206 = w5796 & w9548;
assign w8207 = ~w4415 & ~w11861;
assign w8208 = ~w5805 & ~w2088;
assign w8209 = w15786 & ~w5647;
assign w8210 = w17046 & ~w17082;
assign w8211 = a_11 & a_31;
assign w8212 = ~w16430 & ~w14983;
assign w8213 = ~w4871 & w12210;
assign w8214 = ~w5927 & ~w5899;
assign w8215 = ~w7728 & ~w6408;
assign w8216 = ~w1358 & ~w421;
assign w8217 = ~w13993 & ~w6392;
assign w8218 = w3330 & ~w16479;
assign w8219 = ~w5033 & w16349;
assign w8220 = w3239 & ~w7317;
assign w8221 = w6919 & w19163;
assign w8222 = w5541 & ~w9922;
assign w8223 = ~w680 & ~w13526;
assign w8224 = w10681 & w10972;
assign w8225 = ~w11664 & ~w8268;
assign w8226 = w7369 & ~w18314;
assign w8227 = ~w15245 & w9735;
assign w8228 = ~w15837 & w9318;
assign w8229 = a_9 & a_61;
assign w8230 = ~w17401 & w18115;
assign w8231 = ~w15288 & w18594;
assign w8232 = (~w1776 & ~w18701) | (~w1776 & w11016) | (~w18701 & w11016);
assign w8233 = ~w13184 & ~w15920;
assign w8234 = w8389 & w18793;
assign w8235 = a_0 & a_4;
assign w8236 = ~w9434 & ~w12855;
assign w8237 = w11869 & ~w4521;
assign w8238 = ~w17046 & w17082;
assign w8239 = a_17 & a_59;
assign w8240 = ~w978 & ~w18017;
assign w8241 = w6330 & w17466;
assign w8242 = w17518 & ~w13059;
assign w8243 = a_59 & a_62;
assign w8244 = w2625 & w17893;
assign w8245 = w5055 & ~w14073;
assign w8246 = ~w7222 & w2466;
assign w8247 = a_9 & a_57;
assign w8248 = ~w458 & w15965;
assign w8249 = ~w1616 & ~w13956;
assign w8250 = (w139 & w19005) | (w139 & w16748) | (w19005 & w16748);
assign w8251 = ~w6869 & ~w5553;
assign w8252 = ~w4917 & ~w16204;
assign w8253 = (w14652 & w15047) | (w14652 & w17240) | (w15047 & w17240);
assign w8254 = (~w15340 & ~w14550) | (~w15340 & w3859) | (~w14550 & w3859);
assign w8255 = w6940 | w8965;
assign w8256 = ~w16805 & ~w15033;
assign w8257 = ~w6274 & w564;
assign w8258 = w1638 & w11249;
assign w8259 = ~w8429 & ~w426;
assign w8260 = ~w15663 & w9916;
assign w8261 = ~w13189 & ~w2268;
assign w8262 = w6417 & w12768;
assign w8263 = w243 & ~w11760;
assign w8264 = ~w11835 & ~w1020;
assign w8265 = ~w1910 & ~w3243;
assign w8266 = ~w13805 & ~w3440;
assign w8267 = w10587 & w17174;
assign w8268 = a_23 & a_61;
assign w8269 = w3024 & ~w3222;
assign w8270 = ~w4439 & ~w3095;
assign w8271 = ~w13901 & ~w6652;
assign w8272 = ~w8191 & ~w7351;
assign w8273 = (w16842 & w13082) | (w16842 & w9747) | (w13082 & w9747);
assign w8274 = ~w4257 & w17837;
assign w8275 = ~w464 & ~w5543;
assign w8276 = w2680 & ~w17779;
assign w8277 = ~w5480 & w19164;
assign w8278 = w11170 & ~w10043;
assign w8279 = w10701 & w873;
assign w8280 = ~a_17 & ~w11297;
assign w8281 = ~w15991 & ~w4661;
assign w8282 = ~w1966 & w6246;
assign w8283 = ~w3696 & w16264;
assign w8284 = ~w11739 & ~w15778;
assign w8285 = ~w4004 & ~w15137;
assign w8286 = ~w3830 & ~w18141;
assign w8287 = w16001 & w9017;
assign w8288 = ~w17894 & ~w3701;
assign w8289 = ~w11314 & ~w4659;
assign w8290 = a_39 & a_55;
assign w8291 = ~w6191 & ~w11641;
assign w8292 = ~w6872 & ~w10371;
assign w8293 = w10663 & ~w13523;
assign w8294 = a_56 & a_63;
assign w8295 = ~w4684 & w15571;
assign w8296 = w7786 & ~w6358;
assign w8297 = ~w10568 & w11851;
assign w8298 = a_52 & a_53;
assign w8299 = ~w15007 & ~w6645;
assign w8300 = a_9 & a_22;
assign w8301 = ~w4310 & w624;
assign w8302 = ~w2078 & ~w10950;
assign w8303 = ~w5280 & ~w14683;
assign w8304 = ~w9216 & ~w13515;
assign w8305 = ~w3773 & ~w7906;
assign w8306 = a_11 & a_55;
assign w8307 = ~w5180 & ~w14674;
assign w8308 = ~w13469 & ~w5430;
assign w8309 = ~w5703 & ~w5279;
assign w8310 = ~w15370 & ~w7734;
assign w8311 = w9461 & w6242;
assign w8312 = ~w443 & ~w12588;
assign w8313 = ~w15310 & w1868;
assign w8314 = w8127 & ~w18198;
assign w8315 = w2834 & w11789;
assign w8316 = ~w18678 & w9693;
assign w8317 = ~w4285 & ~w3475;
assign w8318 = ~w349 & ~w10378;
assign w8319 = ~w4070 & ~w17678;
assign w8320 = ~w9310 & ~w7676;
assign w8321 = a_14 & a_48;
assign w8322 = w8214 & w19165;
assign w8323 = a_17 & a_41;
assign w8324 = a_13 & a_37;
assign w8325 = ~w9700 & w9081;
assign w8326 = ~w13713 & ~w17264;
assign w8327 = (w17252 & w97) | (w17252 & w6091) | (w97 & w6091);
assign w8328 = ~w15249 & ~w2761;
assign w8329 = ~w10206 & ~w16831;
assign w8330 = w7214 & ~w14393;
assign w8331 = ~w15115 & w14943;
assign w8332 = a_47 & a_61;
assign w8333 = ~w10311 & ~w4726;
assign w8334 = (~w14005 & ~w6433) | (~w14005 & w6004) | (~w6433 & w6004);
assign w8335 = ~w14724 & ~w9555;
assign w8336 = (w7350 & w4155) | (w7350 & w6660) | (w4155 & w6660);
assign w8337 = w4812 & w6925;
assign w8338 = ~w6409 & ~w15916;
assign w8339 = (~w15613 & ~w13380) | (~w15613 & w14443) | (~w13380 & w14443);
assign w8340 = ~w8828 & ~w4814;
assign w8341 = ~w14628 & ~w3794;
assign w8342 = w10298 & ~w9308;
assign w8343 = a_12 & a_43;
assign w8344 = ~w8010 & ~w14849;
assign w8345 = ~w16612 & ~w6070;
assign w8346 = w3688 & w12049;
assign w8347 = ~w11476 & ~w17520;
assign w8348 = w15003 & w13120;
assign w8349 = ~w10353 & ~w8687;
assign w8350 = ~w4578 & ~w17652;
assign w8351 = ~w6579 & ~w7330;
assign w8352 = ~w2701 & ~w2364;
assign w8353 = ~w12861 & ~w7297;
assign w8354 = w10245 & ~w8436;
assign w8355 = ~w17963 & ~w11274;
assign w8356 = ~w5110 & ~w5024;
assign w8357 = ~w10003 & ~w1541;
assign w8358 = w16363 & ~w4582;
assign w8359 = a_10 & a_41;
assign w8360 = a_24 & a_32;
assign w8361 = ~w2916 & ~w16256;
assign w8362 = a_26 & a_58;
assign w8363 = ~w1284 & ~w16043;
assign w8364 = ~w9912 & ~w1830;
assign w8365 = w11616 & w16374;
assign w8366 = w2743 & ~w1862;
assign w8367 = ~w6613 & ~w12832;
assign w8368 = ~w17960 & w2067;
assign w8369 = ~w10508 & ~w9554;
assign w8370 = w17826 & w6635;
assign w8371 = a_33 & a_62;
assign w8372 = ~w17061 & ~w967;
assign w8373 = ~w15824 & w8986;
assign w8374 = w4243 & w6747;
assign w8375 = ~w101 & ~w6826;
assign w8376 = w16318 & ~w16020;
assign w8377 = ~w15711 & w18007;
assign w8378 = w15911 & ~w11476;
assign w8379 = ~w5051 & ~w3943;
assign w8380 = ~w7262 & ~w7286;
assign w8381 = w2108 & ~w16146;
assign w8382 = ~w15953 & ~w12418;
assign w8383 = ~w7417 & ~w6697;
assign w8384 = ~w11190 & ~w3527;
assign w8385 = ~w17997 & ~w803;
assign w8386 = ~w16297 & ~w12352;
assign w8387 = w14622 & ~w9526;
assign w8388 = ~w7423 & w11969;
assign w8389 = ~w14389 & ~w6881;
assign w8390 = ~w4266 & ~w3509;
assign w8391 = ~w14279 & ~w5765;
assign w8392 = ~w10272 & ~w17801;
assign w8393 = ~w14985 & ~w3263;
assign w8394 = ~w881 & ~w1226;
assign w8395 = ~w2029 & w5672;
assign w8396 = ~w14181 & ~w3383;
assign w8397 = ~w3125 & w16335;
assign w8398 = w6985 & ~w2675;
assign w8399 = ~w17515 & ~w45;
assign w8400 = ~w14660 & w17349;
assign w8401 = ~w2989 & ~w13699;
assign w8402 = ~w16103 & ~w17480;
assign w8403 = a_22 & a_58;
assign w8404 = ~w7638 & w9468;
assign w8405 = w13762 & w12263;
assign w8406 = ~w14442 & ~w3043;
assign w8407 = ~w17161 & ~w18997;
assign w8408 = w4375 & ~w1483;
assign w8409 = w5023 & ~w13591;
assign w8410 = ~w3486 & ~w12989;
assign w8411 = ~w944 & w6328;
assign w8412 = ~w4946 & ~w1789;
assign w8413 = a_7 & a_40;
assign w8414 = ~w13129 & ~w547;
assign w8415 = ~w3688 & ~w12049;
assign w8416 = ~w770 & ~w14225;
assign w8417 = a_17 & a_25;
assign w8418 = ~w13914 & ~w9463;
assign w8419 = ~w5620 & ~w8752;
assign w8420 = w16794 & w11176;
assign w8421 = w13684 & ~w17142;
assign w8422 = ~w15938 & ~w9786;
assign w8423 = a_7 & a_45;
assign w8424 = ~w5984 & ~w12248;
assign w8425 = ~w9378 & ~w18018;
assign w8426 = (~w18593 & ~w7314) | (~w18593 & w6726) | (~w7314 & w6726);
assign w8427 = ~w15948 & w662;
assign w8428 = ~w11568 & ~w15750;
assign w8429 = (~w2769 & w175) | (~w2769 & w10146) | (w175 & w10146);
assign w8430 = (w19096 & w2769) | (w19096 & w12155) | (w2769 & w12155);
assign w8431 = w8410 & w10370;
assign w8432 = w9593 & ~w10086;
assign w8433 = ~w3431 & ~w3077;
assign w8434 = ~w161 & ~w12780;
assign w8435 = ~w16363 & w4582;
assign w8436 = ~w9120 & w16723;
assign w8437 = ~w14079 & ~w12509;
assign w8438 = w15575 & w18292;
assign w8439 = ~w10258 & ~w10401;
assign w8440 = ~w6340 & ~w2746;
assign w8441 = ~w16664 & ~w14836;
assign w8442 = ~w11099 & ~w11093;
assign w8443 = ~w2139 & w18653;
assign w8444 = w16331 & w829;
assign w8445 = w4841 & w16168;
assign w8446 = ~w5549 & w13907;
assign w8447 = w1016 & ~w6071;
assign w8448 = ~w12415 & ~w18614;
assign w8449 = w9534 & ~w10202;
assign w8450 = w3469 & ~w17888;
assign w8451 = ~w14249 & w9339;
assign w8452 = w3855 & w838;
assign w8453 = ~w2354 & ~w12706;
assign w8454 = ~w9830 & ~w13586;
assign w8455 = ~w5108 & w7920;
assign w8456 = ~w14311 & w5952;
assign w8457 = ~w5165 & w7095;
assign w8458 = ~w10129 & ~w19056;
assign w8459 = ~w16929 & ~w6506;
assign w8460 = w18385 & ~w1459;
assign w8461 = ~w19134 & w8951;
assign w8462 = ~w8450 & ~w14340;
assign w8463 = ~w4883 & w2234;
assign w8464 = ~w4702 & w16765;
assign w8465 = ~w5844 & ~w15146;
assign w8466 = w11990 & ~w18349;
assign w8467 = w11104 & w17749;
assign w8468 = a_32 & a_37;
assign w8469 = ~w16766 & ~w5008;
assign w8470 = ~w4308 & w902;
assign w8471 = (~w2597 & ~w2603) | (~w2597 & w18527) | (~w2603 & w18527);
assign w8472 = (w4394 & w4605) | (w4394 & ~w9252) | (w4605 & ~w9252);
assign w8473 = w14783 & ~w4146;
assign w8474 = ~w464 & ~w3265;
assign w8475 = ~w5949 & w19166;
assign w8476 = w9044 & w3152;
assign w8477 = (w17004 & ~w2454) | (w17004 & w18890) | (~w2454 & w18890);
assign w8478 = ~w16834 & ~w788;
assign w8479 = ~w4612 & ~w10871;
assign w8480 = ~w8737 & w8454;
assign w8481 = (w10795 & w5527) | (w10795 & w8973) | (w5527 & w8973);
assign w8482 = ~w4503 & ~w14133;
assign w8483 = w5681 & ~w14747;
assign w8484 = ~w16054 & ~w13910;
assign w8485 = w10099 & w983;
assign w8486 = w10158 & w17931;
assign w8487 = w8909 & ~w7783;
assign w8488 = ~w5319 & ~w1005;
assign w8489 = ~w17211 & ~w6933;
assign w8490 = ~w16529 & w9179;
assign w8491 = ~w14286 & ~w11443;
assign w8492 = w3400 & ~w14779;
assign w8493 = (w1648 & w8126) | (w1648 & w13588) | (w8126 & w13588);
assign w8494 = w5544 & ~w9900;
assign w8495 = ~w19008 & ~w3361;
assign w8496 = ~w16709 & ~w16175;
assign w8497 = ~w9579 & ~w19046;
assign w8498 = w1980 & ~w1255;
assign w8499 = w15504 & ~w2949;
assign w8500 = ~w14577 & ~w4487;
assign w8501 = ~w7501 & w3942;
assign w8502 = ~w1060 & ~w10540;
assign w8503 = ~w6038 & ~w11284;
assign w8504 = w4202 & w1073;
assign w8505 = ~w10271 & ~w373;
assign w8506 = ~w4764 & ~w6419;
assign w8507 = a_35 & a_58;
assign w8508 = w13221 & w3826;
assign w8509 = ~w2612 & ~w710;
assign w8510 = ~w10325 & w3620;
assign w8511 = w461 & ~w2458;
assign w8512 = ~w17851 & w3906;
assign w8513 = ~w18458 & w12034;
assign w8514 = w19032 & ~w430;
assign w8515 = ~w10965 & ~w11702;
assign w8516 = w14024 & ~w12264;
assign w8517 = ~w6932 & ~w14147;
assign w8518 = ~w9835 & w12930;
assign w8519 = w1903 & ~w11449;
assign w8520 = ~w4116 & ~w10590;
assign w8521 = ~w11577 & w6391;
assign w8522 = w7992 & ~w9174;
assign w8523 = w13303 & w17227;
assign w8524 = ~w11990 & w18349;
assign w8525 = (~w3999 & ~w6461) | (~w3999 & w2560) | (~w6461 & w2560);
assign w8526 = ~w6766 & ~w7096;
assign w8527 = w9729 & ~w4140;
assign w8528 = w7152 & ~w16271;
assign w8529 = w8868 & ~w14549;
assign w8530 = ~w13024 & w14762;
assign w8531 = (w15788 & w10532) | (w15788 & w10977) | (w10532 & w10977);
assign w8532 = ~w18520 & ~w15548;
assign w8533 = w13647 & ~w18087;
assign w8534 = ~w4411 & w15140;
assign w8535 = ~w490 & ~w17423;
assign w8536 = (~w12526 & ~w14300) | (~w12526 & w15038) | (~w14300 & w15038);
assign w8537 = ~w9505 & ~w7455;
assign w8538 = ~w6338 & w13963;
assign w8539 = ~w11934 & ~w10903;
assign w8540 = w5337 & ~w1869;
assign w8541 = ~w18908 & w14404;
assign w8542 = ~w16412 & w3628;
assign w8543 = ~w6089 & ~w6435;
assign w8544 = a_3 & a_48;
assign w8545 = (~w5357 & ~w1780) | (~w5357 & w6574) | (~w1780 & w6574);
assign w8546 = w1733 & ~w17884;
assign w8547 = a_41 & a_58;
assign w8548 = ~w7704 & w16613;
assign w8549 = (w6347 & w19005) | (w6347 & w18870) | (w19005 & w18870);
assign w8550 = ~w747 & ~w13564;
assign w8551 = ~w6737 & ~w9638;
assign w8552 = a_40 & a_54;
assign w8553 = ~w8196 & ~w11252;
assign w8554 = ~w11254 & ~w9050;
assign w8555 = ~w12464 & ~w9959;
assign w8556 = (w8896 & w9058) | (w8896 & w15662) | (w9058 & w15662);
assign w8557 = ~w7469 & ~w14270;
assign w8558 = w9320 & w13701;
assign w8559 = w10648 & ~w18995;
assign w8560 = ~w1001 & ~w18378;
assign w8561 = a_13 & a_47;
assign w8562 = ~w11582 & ~w8189;
assign w8563 = ~w14619 & ~w13192;
assign w8564 = (~w1426 & ~w10183) | (~w1426 & w10895) | (~w10183 & w10895);
assign w8565 = w5378 & ~w10576;
assign w8566 = (w11351 & w13082) | (w11351 & w9863) | (w13082 & w9863);
assign w8567 = w4481 & ~w5871;
assign w8568 = w9809 & w2153;
assign w8569 = ~w4154 & ~w8804;
assign w8570 = a_48 & a_52;
assign w8571 = w9117 & w12735;
assign w8572 = ~w9192 & ~w17810;
assign w8573 = ~w12984 & ~w108;
assign w8574 = a_11 & a_38;
assign w8575 = w16143 & ~w12020;
assign w8576 = a_17 & a_20;
assign w8577 = ~w10793 & ~w16347;
assign w8578 = ~w1780 & w6856;
assign w8579 = a_2 & a_51;
assign w8580 = w17476 & ~w6162;
assign w8581 = w2253 & w4071;
assign w8582 = w4296 & ~w17198;
assign w8583 = w13794 & w5045;
assign w8584 = ~w10242 & w6033;
assign w8585 = ~w10744 & ~w11461;
assign w8586 = w4233 & w7803;
assign w8587 = ~w5930 & w11554;
assign w8588 = ~w9981 & ~w1672;
assign w8589 = a_1 & a_41;
assign w8590 = ~w15209 & ~w13472;
assign w8591 = ~w3606 & ~w13628;
assign w8592 = w12131 & ~w796;
assign w8593 = ~w9744 & ~w6613;
assign w8594 = ~w440 & ~w10948;
assign w8595 = ~w357 & ~w7137;
assign w8596 = w1921 & w10457;
assign w8597 = a_6 & a_11;
assign w8598 = ~w17638 & w13000;
assign w8599 = w2068 & ~w17556;
assign w8600 = ~w2695 & ~w13691;
assign w8601 = ~w783 & ~w11101;
assign w8602 = ~w506 & ~w7579;
assign w8603 = ~w12871 & ~w9497;
assign w8604 = w4798 & w10105;
assign w8605 = w6356 & ~w5909;
assign w8606 = ~w11045 & ~w18160;
assign w8607 = w15596 & w9783;
assign w8608 = ~w12252 & w8856;
assign w8609 = w11399 & w17187;
assign w8610 = ~w15237 & w990;
assign w8611 = ~w6955 & ~w5755;
assign w8612 = ~w5074 & w13830;
assign w8613 = ~w10346 & ~w18055;
assign w8614 = a_31 & a_51;
assign w8615 = ~w16063 & ~w5081;
assign w8616 = ~w5159 & ~w9660;
assign w8617 = ~w15004 & ~w17106;
assign w8618 = ~w1895 & ~w5747;
assign w8619 = ~w13720 & ~w8527;
assign w8620 = w1336 & ~w16508;
assign w8621 = w9581 & w7502;
assign w8622 = ~w16076 & ~w7959;
assign w8623 = ~w10264 & ~w13659;
assign w8624 = w16095 & w1873;
assign w8625 = ~w3664 & ~w6651;
assign w8626 = a_23 & a_29;
assign w8627 = ~w8167 & ~w8766;
assign w8628 = (~w16702 & ~w17428) | (~w16702 & w2020) | (~w17428 & w2020);
assign w8629 = ~w1921 & ~w10457;
assign w8630 = w12586 & w1614;
assign w8631 = ~w4305 & ~w10343;
assign w8632 = ~w7958 & ~w6092;
assign w8633 = ~w3995 & ~w2515;
assign w8634 = a_19 & a_29;
assign w8635 = w7825 & w14221;
assign w8636 = ~w15126 & ~w5846;
assign w8637 = (~w2569 & ~w10236) | (~w2569 & w4072) | (~w10236 & w4072);
assign w8638 = ~w11 & w15198;
assign w8639 = ~w4312 & ~w7409;
assign w8640 = a_8 & a_15;
assign w8641 = ~w16751 & ~w4898;
assign w8642 = ~w14534 & ~w11130;
assign w8643 = ~w2064 & ~w12254;
assign w8644 = w14642 & w6575;
assign w8645 = ~w3343 & ~w14265;
assign w8646 = ~w2247 & ~w3944;
assign w8647 = w3713 & ~w14111;
assign w8648 = ~w3169 & ~w14619;
assign w8649 = (~w430 & ~w14770) | (~w430 & w8514) | (~w14770 & w8514);
assign w8650 = ~w6711 & ~w3145;
assign w8651 = ~w17993 & ~w7375;
assign w8652 = a_10 & a_39;
assign w8653 = a_2 & a_39;
assign w8654 = w5956 & w11797;
assign w8655 = (a_55 & w4804) | (a_55 & w14936) | (w4804 & w14936);
assign w8656 = a_19 & a_52;
assign w8657 = a_8 & a_28;
assign w8658 = w16626 & ~w6911;
assign w8659 = w7073 & w10944;
assign w8660 = w11559 & ~w9257;
assign w8661 = w8098 & ~w17910;
assign w8662 = w3221 & ~w10830;
assign w8663 = ~w6853 & w6407;
assign w8664 = ~w7709 & w6151;
assign w8665 = w1962 & w11604;
assign w8666 = ~w5625 & ~w6137;
assign w8667 = ~w17834 & ~w18650;
assign w8668 = ~w18657 & ~w17775;
assign w8669 = ~w11123 & ~w5200;
assign w8670 = (w3601 & w10405) | (w3601 & w6345) | (w10405 & w6345);
assign w8671 = ~w4688 & ~w14048;
assign w8672 = ~w17855 & ~w3534;
assign w8673 = ~w1724 & ~w13402;
assign w8674 = ~w4068 & w18851;
assign w8675 = ~w14299 & ~w15189;
assign w8676 = ~w1457 & ~w2125;
assign w8677 = ~w18070 & ~w4476;
assign w8678 = ~w12297 & w394;
assign w8679 = ~w18099 & w18139;
assign w8680 = w18640 & w19167;
assign w8681 = w15204 & w15271;
assign w8682 = a_20 & a_29;
assign w8683 = ~w15595 & w1306;
assign w8684 = w11546 & w18810;
assign w8685 = a_42 & w15843;
assign w8686 = ~w6669 & ~w16736;
assign w8687 = w14199 & w7858;
assign w8688 = ~w18820 & ~w6389;
assign w8689 = ~w6899 & ~w14953;
assign w8690 = a_31 & a_54;
assign w8691 = ~w13082 & w7686;
assign w8692 = a_16 & a_26;
assign w8693 = ~w5285 & ~w8504;
assign w8694 = ~w721 & w543;
assign w8695 = ~w17272 & w833;
assign w8696 = ~w7327 & ~w10997;
assign w8697 = w16161 & w11076;
assign w8698 = ~w14539 & ~w16220;
assign w8699 = (~w9337 & w13595) | (~w9337 & w140) | (w13595 & w140);
assign w8700 = (w1394 & w2769) | (w1394 & w13929) | (w2769 & w13929);
assign w8701 = a_25 & a_33;
assign w8702 = a_3 & a_55;
assign w8703 = w8803 & ~w5240;
assign w8704 = (w2769 & w15825) | (w2769 & w7763) | (w15825 & w7763);
assign w8705 = w16486 & w7051;
assign w8706 = w6535 & ~w2862;
assign w8707 = ~w16510 & w18382;
assign w8708 = ~w2456 & ~w16598;
assign w8709 = ~w11798 & ~w6827;
assign w8710 = a_19 & a_46;
assign w8711 = a_8 & a_26;
assign w8712 = ~w4948 & ~w4001;
assign w8713 = w16892 & ~w19001;
assign w8714 = ~w10763 & w7236;
assign w8715 = w8505 & ~w11147;
assign w8716 = ~w1586 & w10192;
assign w8717 = ~w16942 & ~w9973;
assign w8718 = a_33 & a_53;
assign w8719 = ~w17463 & ~w7587;
assign w8720 = ~w11045 & w13532;
assign w8721 = ~w15960 & ~w5363;
assign w8722 = (w6834 & ~w13979) | (w6834 & w10820) | (~w13979 & w10820);
assign w8723 = w3898 & ~w5812;
assign w8724 = ~w8842 & ~w11700;
assign w8725 = ~w13088 & ~w3720;
assign w8726 = ~w7129 & w6853;
assign w8727 = w5587 & w14455;
assign w8728 = w6527 & ~w18486;
assign w8729 = ~w6204 & ~w6403;
assign w8730 = ~w5636 & w17509;
assign w8731 = w12423 & ~w9141;
assign w8732 = ~w9625 & ~w7084;
assign w8733 = ~w11305 & w7947;
assign w8734 = ~w7074 & w7054;
assign w8735 = w12430 & ~w7908;
assign w8736 = ~w6781 & ~w7301;
assign w8737 = w18033 & w3379;
assign w8738 = w2182 & ~w10800;
assign w8739 = w5739 & w308;
assign w8740 = ~w4369 & ~w885;
assign w8741 = w7270 & ~w11591;
assign w8742 = a_24 & a_38;
assign w8743 = w17982 & ~w2931;
assign w8744 = w2970 & w8509;
assign w8745 = a_32 & a_59;
assign w8746 = w2016 & w19068;
assign w8747 = (~w332 & ~w7091) | (~w332 & w15748) | (~w7091 & w15748);
assign w8748 = ~w9390 & w6317;
assign w8749 = a_36 & a_48;
assign w8750 = ~w1666 & ~w3094;
assign w8751 = ~w12874 & ~w17041;
assign w8752 = ~w18893 & ~w1537;
assign w8753 = a_9 & a_43;
assign w8754 = ~w9464 & ~w17060;
assign w8755 = w9230 & ~w359;
assign w8756 = ~w11192 & w3470;
assign w8757 = ~w2512 & ~w9612;
assign w8758 = ~w7163 & ~w2808;
assign w8759 = a_41 & a_43;
assign w8760 = ~w1321 & w6353;
assign w8761 = ~w6958 & ~w8598;
assign w8762 = w16474 & w17334;
assign w8763 = a_34 & a_39;
assign w8764 = ~w6754 & w9342;
assign w8765 = ~w14817 & ~w18003;
assign w8766 = ~w12987 & w7499;
assign w8767 = ~w5780 & ~w14500;
assign w8768 = w6253 & w17261;
assign w8769 = ~w6520 & ~w9450;
assign w8770 = a_10 & a_25;
assign w8771 = a_40 & a_55;
assign w8772 = ~w4937 & ~w17687;
assign w8773 = a_23 & a_30;
assign w8774 = ~w12657 & ~w2765;
assign w8775 = w13844 & w17112;
assign w8776 = ~w18438 & ~w8501;
assign w8777 = ~w15420 & ~w15024;
assign w8778 = w17681 & w3362;
assign w8779 = w8555 & ~w2614;
assign w8780 = ~w5884 & ~w12642;
assign w8781 = ~w3869 & ~w2617;
assign w8782 = a_47 & a_50;
assign w8783 = ~w2103 & ~w8674;
assign w8784 = w9634 & ~w358;
assign w8785 = ~w9702 & w12757;
assign w8786 = ~w7504 & ~w7382;
assign w8787 = ~w4658 & w2392;
assign w8788 = w11897 & ~w16017;
assign w8789 = ~w4297 & ~w12610;
assign w8790 = w4108 & w10084;
assign w8791 = ~w13498 & ~w7002;
assign w8792 = w2606 & w15484;
assign w8793 = a_6 & a_33;
assign w8794 = w4694 & w15340;
assign w8795 = ~w7367 & ~w8733;
assign w8796 = w17280 & w10915;
assign w8797 = ~w10137 & w12253;
assign w8798 = ~w4278 & ~w7589;
assign w8799 = a_13 & a_17;
assign w8800 = ~w7505 & ~w8155;
assign w8801 = w329 & w13058;
assign w8802 = ~w3496 & ~w17860;
assign w8803 = ~w2310 & ~w8562;
assign w8804 = ~w11536 & w6395;
assign w8805 = ~w1739 & ~w16772;
assign w8806 = a_44 & a_62;
assign w8807 = ~w9803 & ~w1871;
assign w8808 = ~w3363 & ~w16932;
assign w8809 = ~w1285 & ~w16134;
assign w8810 = a_7 & a_37;
assign w8811 = w11907 & ~w1751;
assign w8812 = ~w18647 & w9674;
assign w8813 = w695 & ~w4445;
assign w8814 = ~w14402 & ~w12143;
assign w8815 = ~w14306 & ~w14596;
assign w8816 = (~w1000 & ~w243) | (~w1000 & w1973) | (~w243 & w1973);
assign w8817 = w16039 & ~w2049;
assign w8818 = ~w4684 & ~w15571;
assign w8819 = ~w4261 & ~w3791;
assign w8820 = w12042 & w7568;
assign w8821 = w17282 & w16389;
assign w8822 = ~w17295 & w17267;
assign w8823 = w15081 & w5109;
assign w8824 = ~w5263 & ~w996;
assign w8825 = w15764 & ~w11495;
assign w8826 = ~w12468 & w8851;
assign w8827 = w6643 & ~w9951;
assign w8828 = ~w16882 & w2729;
assign w8829 = a_33 & a_34;
assign w8830 = ~w18249 & w14621;
assign w8831 = ~w5617 & w574;
assign w8832 = ~w7702 & ~w15943;
assign w8833 = (~w6624 & w14831) | (~w6624 & w14806) | (w14831 & w14806);
assign w8834 = w15948 & ~w662;
assign w8835 = ~w16188 & w17378;
assign w8836 = w12595 & w17581;
assign w8837 = ~w8060 & w11613;
assign w8838 = w18508 & w14438;
assign w8839 = w10817 & ~w17163;
assign w8840 = ~w12807 & w18662;
assign w8841 = w3655 & w12172;
assign w8842 = ~w3960 & ~w1407;
assign w8843 = (~w16832 & ~w5087) | (~w16832 & w4914) | (~w5087 & w4914);
assign w8844 = ~w187 & w17980;
assign w8845 = w9996 & w15045;
assign w8846 = ~w2661 & ~w4094;
assign w8847 = ~w4724 & ~w12573;
assign w8848 = ~w17363 & ~w5589;
assign w8849 = ~w18113 & ~w4837;
assign w8850 = w5247 & w13061;
assign w8851 = ~w15107 & ~w14164;
assign w8852 = w17819 & w737;
assign w8853 = a_50 & a_53;
assign w8854 = ~w1905 & ~w4973;
assign w8855 = ~w11894 & ~w6555;
assign w8856 = ~w14574 & ~w9575;
assign w8857 = w18188 & ~w16121;
assign w8858 = ~w1810 & w10718;
assign w8859 = ~w18972 & ~w15666;
assign w8860 = ~w8584 & w14713;
assign w8861 = ~w8819 & w16850;
assign w8862 = ~w5177 & ~w5369;
assign w8863 = ~w15362 & ~w2455;
assign w8864 = (~w16913 & ~w5578) | (~w16913 & w2382) | (~w5578 & w2382);
assign w8865 = (~w135 & ~w4390) | (~w135 & w18120) | (~w4390 & w18120);
assign w8866 = ~w18938 & ~w2505;
assign w8867 = w18099 & ~w18139;
assign w8868 = ~w16785 & w472;
assign w8869 = w16462 & w2355;
assign w8870 = ~w3240 & ~w16829;
assign w8871 = w1586 & ~w10192;
assign w8872 = ~w15767 & ~w489;
assign w8873 = ~w2051 & ~w3564;
assign w8874 = ~w4150 & ~w670;
assign w8875 = ~w6815 & ~w12318;
assign w8876 = w15115 & ~w14943;
assign w8877 = w15749 & ~w14456;
assign w8878 = a_55 & a_61;
assign w8879 = (~w2769 & w17854) | (~w2769 & w4704) | (w17854 & w4704);
assign w8880 = w16229 & w2516;
assign w8881 = ~w4665 & w7156;
assign w8882 = ~w15411 & w18780;
assign w8883 = ~w13858 & ~w15788;
assign w8884 = ~w14920 & w7412;
assign w8885 = w10824 & ~w640;
assign w8886 = ~w3040 & ~w16255;
assign w8887 = w14705 & ~w4941;
assign w8888 = w6100 & w6306;
assign w8889 = w6027 & ~w1561;
assign w8890 = ~w13030 & w14081;
assign w8891 = w12893 & ~w13902;
assign w8892 = ~w2603 & w6193;
assign w8893 = ~w13821 & ~w12747;
assign w8894 = ~w1478 & ~w2263;
assign w8895 = ~w5530 & ~w15924;
assign w8896 = ~w7161 & ~w10224;
assign w8897 = ~w10604 & ~w12965;
assign w8898 = w7951 & ~w4560;
assign w8899 = w12807 & ~w18662;
assign w8900 = ~w18977 & w17339;
assign w8901 = w16372 & w930;
assign w8902 = ~w12163 & ~w2368;
assign w8903 = a_30 & a_58;
assign w8904 = ~w5164 & ~w4592;
assign w8905 = ~w17331 & ~w2403;
assign w8906 = a_9 & a_62;
assign w8907 = w2752 & w19048;
assign w8908 = ~w9626 & w2442;
assign w8909 = ~w3458 & ~w5856;
assign w8910 = ~w4003 & ~w17763;
assign w8911 = ~w2943 & ~w13570;
assign w8912 = ~w5189 & w2459;
assign w8913 = ~w9880 & ~w10945;
assign w8914 = w9705 & ~w1145;
assign w8915 = ~a_34 & a_35;
assign w8916 = w12627 & ~w896;
assign w8917 = ~w13335 & ~w7678;
assign w8918 = ~w9279 & ~w202;
assign w8919 = ~w15563 & ~w17029;
assign w8920 = w18711 & w671;
assign w8921 = ~w6473 & w1227;
assign w8922 = w17830 & w2877;
assign w8923 = ~w10509 & ~w16089;
assign w8924 = ~w12010 & w12969;
assign w8925 = w10350 & ~w1249;
assign w8926 = ~w821 & ~w14174;
assign w8927 = w10557 & ~w4832;
assign w8928 = a_32 & a_45;
assign w8929 = w3907 & w13652;
assign w8930 = (~w9957 & ~w2771) | (~w9957 & w0) | (~w2771 & w0);
assign w8931 = ~w10495 & w14342;
assign w8932 = w2591 & ~w282;
assign w8933 = w6853 & w15763;
assign w8934 = ~w5732 & ~w2719;
assign w8935 = ~w16160 & ~w8571;
assign w8936 = ~w10473 & w11955;
assign w8937 = (~w1709 & ~w2465) | (~w1709 & w14143) | (~w2465 & w14143);
assign w8938 = ~w16818 & ~w6475;
assign w8939 = ~w6444 & ~w1285;
assign w8940 = ~w11745 & w2879;
assign w8941 = w11287 & w3348;
assign w8942 = ~w16240 & ~w11460;
assign w8943 = a_48 & a_61;
assign w8944 = w2361 | w2615;
assign w8945 = ~w6459 & ~w10870;
assign w8946 = w13744 & ~w3323;
assign w8947 = ~w16858 & ~w1356;
assign w8948 = ~w11189 & w17969;
assign w8949 = ~w9211 & ~w14700;
assign w8950 = ~w10153 & ~w7833;
assign w8951 = ~w16279 & ~w19137;
assign w8952 = w157 & ~w4269;
assign w8953 = ~w14316 & ~w17333;
assign w8954 = ~w17963 & w18435;
assign w8955 = (~w766 & ~w17958) | (~w766 & w4668) | (~w17958 & w4668);
assign w8956 = ~w17599 & w6584;
assign w8957 = ~w19073 & ~w8630;
assign w8958 = w6798 & ~w5404;
assign w8959 = w5257 & ~w18069;
assign w8960 = ~w171 & w8402;
assign w8961 = w17753 & ~w1910;
assign w8962 = a_8 & a_30;
assign w8963 = w5091 & w6720;
assign w8964 = w18051 & ~w7362;
assign w8965 = ~w18654 & w11949;
assign w8966 = w4665 & ~w7156;
assign w8967 = (w13981 & w18868) | (w13981 & w2645) | (w18868 & w2645);
assign w8968 = w7607 & w7024;
assign w8969 = w14595 & ~w5281;
assign w8970 = w6000 & ~w2570;
assign w8971 = ~w2596 & ~w18534;
assign w8972 = (w63 & w16041) | (w63 & w17203) | (w16041 & w17203);
assign w8973 = ~w7409 & w2121;
assign w8974 = ~w10811 & ~w10767;
assign w8975 = w13979 & w15011;
assign w8976 = w9405 & ~w5820;
assign w8977 = w3195 & w10411;
assign w8978 = ~w10406 & ~w5330;
assign w8979 = a_55 & a_57;
assign w8980 = w12060 & ~w12755;
assign w8981 = ~w19116 & w16174;
assign w8982 = a_33 & a_36;
assign w8983 = w8214 & w8678;
assign w8984 = w8786 & ~w7814;
assign w8985 = w12391 & w9031;
assign w8986 = ~w8686 & ~w14681;
assign w8987 = (w2206 & w2896) | (w2206 & w7896) | (w2896 & w7896);
assign w8988 = (~w3695 & w2769) | (~w3695 & w7727) | (w2769 & w7727);
assign w8989 = ~w12369 & w731;
assign w8990 = w15619 & ~w17412;
assign w8991 = ~w16462 & ~w2355;
assign w8992 = w12782 & ~w9703;
assign w8993 = w3830 & w18141;
assign w8994 = ~w2324 & ~w1610;
assign w8995 = ~w11692 & ~w2381;
assign w8996 = ~w74 & ~w13739;
assign w8997 = w14012 & ~w4620;
assign w8998 = ~w12710 & ~w1076;
assign w8999 = ~w10792 & ~w2395;
assign w9000 = ~w4351 & w2519;
assign w9001 = w11610 & ~w11093;
assign w9002 = (~w5139 & ~w10591) | (~w5139 & w81) | (~w10591 & w81);
assign w9003 = ~w9475 & ~w17252;
assign w9004 = ~w16425 & ~w16154;
assign w9005 = ~w5244 & ~w10326;
assign w9006 = w15730 & ~w9710;
assign w9007 = w6853 & w8258;
assign w9008 = a_21 & a_30;
assign w9009 = w10287 & ~w10934;
assign w9010 = a_1 & a_54;
assign w9011 = ~w4180 & w4799;
assign w9012 = ~w10624 & ~w3653;
assign w9013 = ~w7902 & w12929;
assign w9014 = ~w6638 & ~w16535;
assign w9015 = w16503 & w10140;
assign w9016 = ~w13304 & ~w14250;
assign w9017 = ~w1397 & ~w2266;
assign w9018 = w12797 & ~w13170;
assign w9019 = ~w18786 & ~w3744;
assign w9020 = ~w17397 & ~w11102;
assign w9021 = ~w11862 & w3755;
assign w9022 = w6446 & ~w15834;
assign w9023 = w16131 & w2532;
assign w9024 = ~w1679 & w4251;
assign w9025 = w2454 & ~w17589;
assign w9026 = w11977 & ~w3933;
assign w9027 = a_8 & a_49;
assign w9028 = ~w9980 & ~w15848;
assign w9029 = ~w11559 & w9257;
assign w9030 = ~w1603 & ~w1651;
assign w9031 = ~w6154 & ~w9672;
assign w9032 = w2531 & w3614;
assign w9033 = (~w7102 & w484) | (~w7102 & w16716) | (w484 & w16716);
assign w9034 = ~w4107 & w13225;
assign w9035 = a_39 & a_42;
assign w9036 = ~w10110 & ~w7781;
assign w9037 = ~w15332 & ~w16490;
assign w9038 = ~w12060 & w16052;
assign w9039 = a_21 & a_49;
assign w9040 = ~w904 & ~w6596;
assign w9041 = ~w13851 & ~w10561;
assign w9042 = ~w16784 & ~w12845;
assign w9043 = ~w1950 & ~w15212;
assign w9044 = a_52 & a_56;
assign w9045 = ~w3604 & ~w9676;
assign w9046 = ~w201 & ~w7937;
assign w9047 = w12108 & ~w16684;
assign w9048 = ~w3336 & ~w3320;
assign w9049 = ~a_2 & a_3;
assign w9050 = w15428 & w8413;
assign w9051 = w8229 & ~w9429;
assign w9052 = ~w16744 & ~w1108;
assign w9053 = ~w14714 & ~w4677;
assign w9054 = a_30 & a_49;
assign w9055 = w6043 & ~w14243;
assign w9056 = ~w10596 & ~w803;
assign w9057 = ~w1034 & w2063;
assign w9058 = ~w6178 & ~w6365;
assign w9059 = ~w4406 & ~w1276;
assign w9060 = ~w13174 & ~w10375;
assign w9061 = ~w15508 & ~w12368;
assign w9062 = ~w18185 & w2879;
assign w9063 = w16782 & w12675;
assign w9064 = a_29 & a_45;
assign w9065 = (~w18967 & ~w5724) | (~w18967 & w3712) | (~w5724 & w3712);
assign w9066 = ~w7192 & ~w18589;
assign w9067 = w2367 & w5444;
assign w9068 = (~w17276 & ~w2242) | (~w17276 & w16059) | (~w2242 & w16059);
assign w9069 = ~w17101 & w746;
assign w9070 = ~w14106 & ~w13205;
assign w9071 = ~w17600 & w6935;
assign w9072 = a_4 & a_8;
assign w9073 = w10657 & w16277;
assign w9074 = ~w9945 & ~w18065;
assign w9075 = a_42 & a_62;
assign w9076 = a_21 & a_35;
assign w9077 = ~w2977 & ~w19118;
assign w9078 = ~w13153 & ~w17650;
assign w9079 = a_30 & a_51;
assign w9080 = ~w2004 & ~w7065;
assign w9081 = ~w95 & ~w4892;
assign w9082 = ~w10557 & w4832;
assign w9083 = w808 & w13926;
assign w9084 = ~w7747 & ~w2981;
assign w9085 = (~w17700 & w5231) | (~w17700 & w5705) | (w5231 & w5705);
assign w9086 = ~w1701 & ~w37;
assign w9087 = ~w8799 & w5792;
assign w9088 = w12617 & ~w3651;
assign w9089 = ~w6385 & w12822;
assign w9090 = ~w13090 & ~w10535;
assign w9091 = ~w10722 & ~w2786;
assign w9092 = ~w10447 & w16370;
assign w9093 = ~w645 & ~w5432;
assign w9094 = w14813 & ~w6053;
assign w9095 = (~w6834 & w6291) | (~w6834 & w18199) | (w6291 & w18199);
assign w9096 = ~w1945 & ~w16207;
assign w9097 = ~w6654 & ~w9497;
assign w9098 = ~w12760 & w15262;
assign w9099 = ~w1061 & w6650;
assign w9100 = ~w16761 & ~w13625;
assign w9101 = ~w15190 & ~w10344;
assign w9102 = (w9337 & w18894) | (w9337 & w17532) | (w18894 & w17532);
assign w9103 = ~w11859 & w16515;
assign w9104 = ~w18240 & w3174;
assign w9105 = w15291 & w4804;
assign w9106 = ~w8505 & w11147;
assign w9107 = w5069 & ~w16679;
assign w9108 = w18560 & ~w18625;
assign w9109 = ~w18734 & ~w2381;
assign w9110 = ~w8233 & w14262;
assign w9111 = (~w19082 & w15009) | (~w19082 & w9215) | (w15009 & w9215);
assign w9112 = ~w104 & ~w5288;
assign w9113 = ~w1519 & ~w9197;
assign w9114 = ~w4675 & ~w7531;
assign w9115 = ~w13843 & ~w2215;
assign w9116 = ~w2449 & ~w9883;
assign w9117 = a_6 & a_43;
assign w9118 = ~w14603 & ~w18296;
assign w9119 = a_19 & a_51;
assign w9120 = ~w10572 & ~w5508;
assign w9121 = ~w1275 & ~w17547;
assign w9122 = ~w247 & ~w10096;
assign w9123 = ~w4421 & ~w14047;
assign w9124 = ~w15621 & w17669;
assign w9125 = w5793 & w1307;
assign w9126 = a_30 & a_36;
assign w9127 = ~w13207 & ~w12907;
assign w9128 = ~w11117 & w18092;
assign w9129 = ~w14843 & ~w1008;
assign w9130 = ~w9250 & ~w1413;
assign w9131 = ~w7326 & ~w1562;
assign w9132 = (~w18975 & ~w17396) | (~w18975 & w13953) | (~w17396 & w13953);
assign w9133 = w16379 & ~w11738;
assign w9134 = ~w3427 & ~w3093;
assign w9135 = w958 & ~w8729;
assign w9136 = ~w10474 & ~w6186;
assign w9137 = w18095 & ~w9910;
assign w9138 = ~w7449 & ~w13566;
assign w9139 = ~w15936 & ~w10892;
assign w9140 = ~w2706 & ~w16758;
assign w9141 = ~w9355 & ~w12579;
assign w9142 = ~w2225 & ~w1495;
assign w9143 = ~w117 & w4196;
assign w9144 = w7355 & w353;
assign w9145 = w13522 & ~w15064;
assign w9146 = w18924 & w164;
assign w9147 = a_33 & w1913;
assign w9148 = ~w2723 & ~w784;
assign w9149 = w4700 & ~w3419;
assign w9150 = w16988 & w3299;
assign w9151 = ~w8612 & ~w10382;
assign w9152 = ~w11742 & w14465;
assign w9153 = w1772 & ~w9853;
assign w9154 = ~w5073 & ~w13894;
assign w9155 = a_6 & a_15;
assign w9156 = w18773 & ~w6678;
assign w9157 = ~w1915 & ~w12466;
assign w9158 = w5893 & ~w8855;
assign w9159 = w17214 & ~w11091;
assign w9160 = ~w12268 & ~w7200;
assign w9161 = ~w4725 & ~w11773;
assign w9162 = ~w1139 & ~w10713;
assign w9163 = ~w3860 & w218;
assign w9164 = ~w14422 & ~w17328;
assign w9165 = ~w15894 & ~w18620;
assign w9166 = ~w16940 & ~w7894;
assign w9167 = ~w6325 & w1350;
assign w9168 = ~w7875 & w15831;
assign w9169 = w19069 & ~w3413;
assign w9170 = a_13 & a_25;
assign w9171 = ~w5760 & ~w8244;
assign w9172 = ~w1081 & ~w17985;
assign w9173 = w4880 & ~w655;
assign w9174 = ~w13675 & ~w14938;
assign w9175 = ~w3971 & ~w13711;
assign w9176 = ~w523 & ~w3112;
assign w9177 = w1118 & ~w17432;
assign w9178 = w12050 & w8833;
assign w9179 = ~w16935 & ~w11806;
assign w9180 = ~w16050 & ~w10738;
assign w9181 = ~w17611 & w12534;
assign w9182 = ~w17740 & ~w10115;
assign w9183 = a_13 & a_33;
assign w9184 = w13534 & w17255;
assign w9185 = w11141 & ~w6461;
assign w9186 = ~w18189 & ~w19045;
assign w9187 = w209 & ~w11911;
assign w9188 = w18451 & w10699;
assign w9189 = ~w4989 & w16343;
assign w9190 = ~w9298 & w41;
assign w9191 = ~w18422 & w1599;
assign w9192 = w18715 & ~w3736;
assign w9193 = ~w14467 & ~w8912;
assign w9194 = ~w6263 & ~w2909;
assign w9195 = ~w3288 & ~w16129;
assign w9196 = ~w4585 & w7053;
assign w9197 = ~w18031 & ~w9507;
assign w9198 = ~w2897 & ~w6067;
assign w9199 = ~w14847 & ~w13984;
assign w9200 = ~w252 & ~w7934;
assign w9201 = ~w8822 & ~w14873;
assign w9202 = ~w18112 & ~w11963;
assign w9203 = ~w13745 & ~w6578;
assign w9204 = w3044 & w3822;
assign w9205 = ~w18910 & ~w12549;
assign w9206 = ~w13468 & ~w17010;
assign w9207 = a_21 & a_25;
assign w9208 = (a_42 & w17379) | (a_42 & w3403) | (w17379 & w3403);
assign w9209 = ~w1992 & ~w16730;
assign w9210 = ~w6633 & ~w5918;
assign w9211 = w5564 & ~w2091;
assign w9212 = ~w13664 & ~w4371;
assign w9213 = ~w17288 & ~w925;
assign w9214 = ~w14701 & w14723;
assign w9215 = w12267 & ~w19082;
assign w9216 = w10243 & w933;
assign w9217 = ~w16002 & ~w16721;
assign w9218 = w1743 & w11039;
assign w9219 = w3314 & ~w1279;
assign w9220 = w15593 & ~w5726;
assign w9221 = ~w9337 & w13052;
assign w9222 = ~w9328 & ~w13183;
assign w9223 = ~w10204 & ~w3234;
assign w9224 = ~w5151 & w1045;
assign w9225 = w2921 & ~w7849;
assign w9226 = ~w1097 & w5479;
assign w9227 = ~w3729 & ~w8074;
assign w9228 = ~w4518 & ~w1543;
assign w9229 = ~w18699 & ~w3388;
assign w9230 = (~w18007 & w14712) | (~w18007 & w15119) | (w14712 & w15119);
assign w9231 = a_45 & a_46;
assign w9232 = w369 & ~w18332;
assign w9233 = ~w6455 & ~w2863;
assign w9234 = ~w7342 & ~w4988;
assign w9235 = ~w3551 & ~w14768;
assign w9236 = w6034 & ~w11175;
assign w9237 = ~w4338 & ~w2486;
assign w9238 = w16948 & ~w6953;
assign w9239 = a_9 & a_32;
assign w9240 = w12337 & w12539;
assign w9241 = ~w1850 & w7258;
assign w9242 = w13392 & ~w10880;
assign w9243 = (~w3485 & ~w16771) | (~w3485 & w15849) | (~w16771 & w15849);
assign w9244 = w2732 & ~w1607;
assign w9245 = ~w13082 & w10860;
assign w9246 = ~w10111 & ~w18379;
assign w9247 = ~w16360 & ~w11780;
assign w9248 = ~w1938 & ~w15269;
assign w9249 = ~w2348 & ~w13009;
assign w9250 = w8482 & ~w13855;
assign w9251 = ~w16267 & w18922;
assign w9252 = (~w5809 & w10770) | (~w5809 & w17641) | (w10770 & w17641);
assign w9253 = ~w2955 & ~w2715;
assign w9254 = ~w5862 & ~w13391;
assign w9255 = w13080 & w17110;
assign w9256 = w7456 & ~w11592;
assign w9257 = ~w15400 & ~w18347;
assign w9258 = ~w4570 & ~w11376;
assign w9259 = ~w13902 & ~w17538;
assign w9260 = ~w19072 & ~w959;
assign w9261 = a_5 & a_18;
assign w9262 = ~w11834 & w15111;
assign w9263 = ~w15423 & ~w2543;
assign w9264 = w10690 & ~w4150;
assign w9265 = ~w18838 & w5134;
assign w9266 = ~w10330 & w17895;
assign w9267 = a_2 & a_29;
assign w9268 = w3591 & ~w10420;
assign w9269 = ~a_60 & a_61;
assign w9270 = (w10232 & w17132) | (w10232 & w1596) | (w17132 & w1596);
assign w9271 = ~w7702 & ~w2296;
assign w9272 = ~w16427 & w9471;
assign w9273 = ~w5667 & ~w5259;
assign w9274 = (~w8226 & ~w16655) | (~w8226 & w17348) | (~w16655 & w17348);
assign w9275 = ~w6169 & ~w2443;
assign w9276 = ~w15627 & ~w12713;
assign w9277 = ~w12761 & ~w385;
assign w9278 = a_27 & a_37;
assign w9279 = w11008 & ~w11679;
assign w9280 = ~w9695 & w6279;
assign w9281 = ~w404 & ~w10832;
assign w9282 = w11711 & w13130;
assign w9283 = ~w2405 & ~w9517;
assign w9284 = (w12151 & w17506) | (w12151 & w6554) | (w17506 & w6554);
assign w9285 = ~w18747 & w13612;
assign w9286 = ~w11731 & ~w1777;
assign w9287 = ~w10639 & w10238;
assign w9288 = w15552 & ~w12968;
assign w9289 = w10541 & ~w5863;
assign w9290 = ~w4098 & ~w4272;
assign w9291 = w15882 & ~w12142;
assign w9292 = ~w12639 & ~w13556;
assign w9293 = (~w2769 & w11853) | (~w2769 & w7144) | (w11853 & w7144);
assign w9294 = w17109 & ~w18144;
assign w9295 = ~w4299 & ~w14878;
assign w9296 = (w10232 & w17132) | (w10232 & w18199) | (w17132 & w18199);
assign w9297 = ~w1201 & ~w17668;
assign w9298 = ~w14024 & w12264;
assign w9299 = ~w2846 & ~w14030;
assign w9300 = (~w230 & ~w2385) | (~w230 & w975) | (~w2385 & w975);
assign w9301 = ~w3378 & ~w10316;
assign w9302 = w8196 & w11252;
assign w9303 = ~w5260 & w309;
assign w9304 = w8341 & w13971;
assign w9305 = ~w10118 & ~w6573;
assign w9306 = w4662 & ~w12701;
assign w9307 = ~w16474 & ~w17334;
assign w9308 = ~w13895 & ~w8690;
assign w9309 = ~w12990 & ~w5178;
assign w9310 = ~w10577 & ~w1533;
assign w9311 = ~w9334 & ~w19021;
assign w9312 = ~w6974 & w3714;
assign w9313 = a_55 & a_56;
assign w9314 = w4882 & ~w12290;
assign w9315 = ~w4194 & ~w5466;
assign w9316 = w2870 & w13420;
assign w9317 = w18182 & ~w11714;
assign w9318 = ~w16879 & ~w3535;
assign w9319 = (~w1428 & w2572) | (~w1428 & w12191) | (w2572 & w12191);
assign w9320 = ~w1018 & ~w10430;
assign w9321 = w8611 & w9725;
assign w9322 = (w11949 & w1119) | (w11949 & ~w5108) | (w1119 & ~w5108);
assign w9323 = a_24 & a_31;
assign w9324 = ~w11569 & ~w10971;
assign w9325 = a_21 & a_40;
assign w9326 = ~w5898 & ~w18613;
assign w9327 = ~w15125 & ~w2789;
assign w9328 = a_5 & a_20;
assign w9329 = ~w10361 & ~w16632;
assign w9330 = ~w3283 & ~w8610;
assign w9331 = a_28 & a_36;
assign w9332 = w15547 & ~w4291;
assign w9333 = a_2 & a_21;
assign w9334 = ~w18775 & w7738;
assign w9335 = w8006 & ~w16336;
assign w9336 = ~w7922 & ~w18535;
assign w9337 = ~w8438 & w5632;
assign w9338 = w1135 & ~w12003;
assign w9339 = ~w10481 & ~w5957;
assign w9340 = ~w17189 & ~w14848;
assign w9341 = a_37 & a_44;
assign w9342 = ~w1102 & ~w13499;
assign w9343 = ~w17606 & w877;
assign w9344 = a_21 & a_45;
assign w9345 = ~w13106 & ~w3977;
assign w9346 = w134 & ~w4148;
assign w9347 = a_27 & a_35;
assign w9348 = a_26 & a_35;
assign w9349 = ~w6692 & ~w11264;
assign w9350 = w3450 & w12884;
assign w9351 = ~w2367 & ~w5444;
assign w9352 = ~w4662 & w3456;
assign w9353 = ~w14921 & ~w2884;
assign w9354 = ~w16130 & ~w3213;
assign w9355 = w5547 & ~w12916;
assign w9356 = ~w1843 & ~w14274;
assign w9357 = ~w12971 & w6224;
assign w9358 = w11405 & w13380;
assign w9359 = w8955 & ~w11096;
assign w9360 = w18175 & ~w7758;
assign w9361 = ~w8988 & ~w6023;
assign w9362 = a_34 & a_63;
assign w9363 = w458 & w14566;
assign w9364 = w11305 & ~w7947;
assign w9365 = w12910 & w3181;
assign w9366 = ~w6514 & ~w13666;
assign w9367 = ~w18899 & ~w5169;
assign w9368 = ~w7273 & w13500;
assign w9369 = ~w1566 & w18419;
assign w9370 = ~w7307 & w3850;
assign w9371 = ~w18333 & ~w444;
assign w9372 = w12419 & w10210;
assign w9373 = w13384 & w8356;
assign w9374 = w17311 & w18655;
assign w9375 = ~w11304 & ~w4190;
assign w9376 = ~w14854 & ~w14775;
assign w9377 = ~w9738 & ~w15461;
assign w9378 = ~w940 & w11275;
assign w9379 = ~w9053 & ~w1615;
assign w9380 = w11656 & ~w16284;
assign w9381 = w15363 & w694;
assign w9382 = w12273 & ~w12714;
assign w9383 = w16028 & ~w7575;
assign w9384 = w12898 & ~w3407;
assign w9385 = w150 & ~w5676;
assign w9386 = w8636 & w15957;
assign w9387 = a_22 & a_32;
assign w9388 = (w6139 & w9656) | (w6139 & w7260) | (w9656 & w7260);
assign w9389 = ~w14487 & ~w16495;
assign w9390 = a_37 & a_54;
assign w9391 = ~w17903 & ~w10064;
assign w9392 = ~w18418 & w5953;
assign w9393 = ~w6658 & w12892;
assign w9394 = (~w11839 & ~w17568) | (~w11839 & w1794) | (~w17568 & w1794);
assign w9395 = ~w15508 & ~w18100;
assign w9396 = (~w9701 & ~w12595) | (~w9701 & w10385) | (~w12595 & w10385);
assign w9397 = w611 & ~w18816;
assign w9398 = w6148 & ~w2776;
assign w9399 = ~w3734 & ~w14362;
assign w9400 = ~w17619 & ~w14995;
assign w9401 = (~w11678 & ~w2253) | (~w11678 & w13026) | (~w2253 & w13026);
assign w9402 = ~w3603 & w16481;
assign w9403 = a_5 & a_25;
assign w9404 = ~w3805 & w4158;
assign w9405 = a_36 & a_54;
assign w9406 = ~w12783 & w16479;
assign w9407 = ~w12332 & ~w10489;
assign w9408 = ~w8430 & ~w1804;
assign w9409 = ~w4164 & ~w3482;
assign w9410 = w432 & ~w11844;
assign w9411 = w8362 & ~w62;
assign w9412 = ~w15430 & ~w14377;
assign w9413 = w1901 & w2604;
assign w9414 = w7353 & w325;
assign w9415 = ~w18860 & ~w1793;
assign w9416 = ~w18911 & w1520;
assign w9417 = w10885 & ~w14743;
assign w9418 = ~w372 & w9806;
assign w9419 = ~w13489 & ~w11400;
assign w9420 = ~w9137 & w18873;
assign w9421 = a_1 & a_19;
assign w9422 = a_4 & a_61;
assign w9423 = ~w14286 & w4906;
assign w9424 = ~w4772 & w11772;
assign w9425 = (w3624 & ~w8747) | (w3624 & w4618) | (~w8747 & w4618);
assign w9426 = ~a_32 & ~w6474;
assign w9427 = ~w3776 & ~w8949;
assign w9428 = ~w850 & w13995;
assign w9429 = ~w398 & ~w14242;
assign w9430 = ~w14803 & ~w1729;
assign w9431 = ~w16836 & ~w9207;
assign w9432 = (w4287 & w13082) | (w4287 & w17988) | (w13082 & w17988);
assign w9433 = (w12255 & w1395) | (w12255 & w14945) | (w1395 & w14945);
assign w9434 = w10472 & w9379;
assign w9435 = (~w10738 & ~w15166) | (~w10738 & w9180) | (~w15166 & w9180);
assign w9436 = w14487 & w16495;
assign w9437 = ~w15846 & ~w15372;
assign w9438 = w10355 & w14675;
assign w9439 = w6566 & ~w18986;
assign w9440 = ~w7601 & ~w6260;
assign w9441 = w18024 & ~w12745;
assign w9442 = w16643 & w16353;
assign w9443 = ~w8090 & ~w16150;
assign w9444 = (w15734 & w6618) | (w15734 & w1797) | (w6618 & w1797);
assign w9445 = a_1 & a_11;
assign w9446 = ~w9173 & ~w3682;
assign w9447 = ~w1314 & ~w2887;
assign w9448 = ~w15554 & ~w17485;
assign w9449 = ~w5005 & ~w18401;
assign w9450 = ~w13114 & ~w9857;
assign w9451 = ~w865 & ~w18778;
assign w9452 = a_16 & a_36;
assign w9453 = ~w18308 & ~w11691;
assign w9454 = a_12 & a_22;
assign w9455 = w12690 & w214;
assign w9456 = a_19 & a_32;
assign w9457 = a_27 & a_45;
assign w9458 = ~w13086 & ~w4957;
assign w9459 = ~w11570 & ~w15157;
assign w9460 = a_2 & a_45;
assign w9461 = ~w14538 & ~w16763;
assign w9462 = w9291 & ~w13938;
assign w9463 = ~w9691 & ~w12499;
assign w9464 = w15911 & w1849;
assign w9465 = ~w14086 & w10874;
assign w9466 = a_5 & a_22;
assign w9467 = ~w3636 & ~w5197;
assign w9468 = ~w4434 & ~w2728;
assign w9469 = ~w19018 & ~w13196;
assign w9470 = w11862 & ~w3755;
assign w9471 = ~w9019 & ~w10476;
assign w9472 = w14086 & ~w10874;
assign w9473 = w10208 & w15267;
assign w9474 = ~w17373 & ~w12192;
assign w9475 = w3078 & w14744;
assign w9476 = a_25 & a_53;
assign w9477 = ~w13504 & ~w12790;
assign w9478 = ~w18248 & ~w8940;
assign w9479 = w12719 & ~w17568;
assign w9480 = a_31 & a_49;
assign w9481 = ~w14544 & ~w9366;
assign w9482 = ~w1939 & ~w9384;
assign w9483 = ~w16236 & ~w14850;
assign w9484 = w4153 & w16273;
assign w9485 = w1345 & w3756;
assign w9486 = ~w13119 & ~w10275;
assign w9487 = ~w7115 & ~w1508;
assign w9488 = w15256 & ~w5526;
assign w9489 = w6846 & w10014;
assign w9490 = ~w9348 & w7516;
assign w9491 = w16328 & w5595;
assign w9492 = a_37 & a_49;
assign w9493 = ~w18592 & ~w16909;
assign w9494 = w11290 & ~w13204;
assign w9495 = ~w8231 & ~w595;
assign w9496 = ~w13642 & ~w17105;
assign w9497 = w1996 & w13127;
assign w9498 = ~w2481 & ~w13867;
assign w9499 = ~w4598 & ~w1043;
assign w9500 = ~w6562 & ~w11025;
assign w9501 = ~w8647 & ~w15023;
assign w9502 = w13771 & ~w5201;
assign w9503 = ~w8590 & ~w3824;
assign w9504 = ~w12331 & w8004;
assign w9505 = w9770 & ~w1014;
assign w9506 = ~w7784 & ~w6532;
assign w9507 = ~w1474 & ~w17325;
assign w9508 = w11834 & ~w15111;
assign w9509 = ~w1961 & ~w17024;
assign w9510 = w15251 & w8771;
assign w9511 = ~w16607 & w19112;
assign w9512 = ~w14392 & ~w10843;
assign w9513 = ~w13946 & ~w18913;
assign w9514 = ~w5972 & ~w14378;
assign w9515 = ~w4646 & ~w16538;
assign w9516 = ~w13827 & ~w6067;
assign w9517 = ~w18493 & ~w7924;
assign w9518 = w14145 & w1634;
assign w9519 = ~w12711 & ~w5531;
assign w9520 = ~w5865 & ~w1215;
assign w9521 = w6853 & w14721;
assign w9522 = w13753 & ~w17014;
assign w9523 = ~w5574 & ~w1782;
assign w9524 = ~w15659 & w8442;
assign w9525 = ~w17303 & ~w16487;
assign w9526 = ~w11575 & ~w14706;
assign w9527 = w9119 & w6458;
assign w9528 = (~w14903 & ~w5934) | (~w14903 & w19074) | (~w5934 & w19074);
assign w9529 = w1085 & ~w4925;
assign w9530 = ~w15316 & ~w12686;
assign w9531 = ~w10364 & ~w1477;
assign w9532 = w7190 & w3008;
assign w9533 = ~w2295 & ~w18731;
assign w9534 = ~w11930 & ~w13574;
assign w9535 = w3418 & w17821;
assign w9536 = ~w18575 & ~w4936;
assign w9537 = ~w6487 & ~w7419;
assign w9538 = (~w12120 & ~w316) | (~w12120 & w13930) | (~w316 & w13930);
assign w9539 = ~w4750 & ~w10809;
assign w9540 = ~w16317 & ~w14911;
assign w9541 = w18211 & ~w10735;
assign w9542 = ~w5532 & w857;
assign w9543 = ~w8060 & ~w6796;
assign w9544 = a_10 & a_17;
assign w9545 = w8632 & ~w13031;
assign w9546 = ~w9816 & ~w5307;
assign w9547 = ~w12167 & ~w5020;
assign w9548 = ~w17209 & ~w18962;
assign w9549 = ~w3124 & ~w3501;
assign w9550 = w6402 & ~w999;
assign w9551 = w14395 & w17941;
assign w9552 = ~w13282 & ~w9796;
assign w9553 = ~w1575 & w16668;
assign w9554 = ~w1812 & w3498;
assign w9555 = ~w11473 & ~w13077;
assign w9556 = ~w2842 & ~w11477;
assign w9557 = ~w7854 & ~w5243;
assign w9558 = w11059 & ~w5419;
assign w9559 = (w15997 & w7143) | (w15997 & w5127) | (w7143 & w5127);
assign w9560 = w3905 & w15054;
assign w9561 = w13178 & ~w9234;
assign w9562 = ~w9127 & ~w12794;
assign w9563 = ~w1924 & ~w18892;
assign w9564 = ~w13973 & ~w5079;
assign w9565 = ~w4101 & w13776;
assign w9566 = ~w5934 & w15273;
assign w9567 = ~w18412 & ~w6133;
assign w9568 = ~w2697 & ~w18994;
assign w9569 = w17307 & ~w4844;
assign w9570 = ~w15537 & ~w4815;
assign w9571 = w1352 & w8270;
assign w9572 = w367 & ~w16180;
assign w9573 = ~w8675 & ~w8142;
assign w9574 = (~w18361 & ~w9585) | (~w18361 & w7132) | (~w9585 & w7132);
assign w9575 = w1492 & w5478;
assign w9576 = ~w2807 & ~w3832;
assign w9577 = ~w10215 & ~w9872;
assign w9578 = w6211 & ~w18623;
assign w9579 = w4766 & w9703;
assign w9580 = ~w13673 & ~w1878;
assign w9581 = ~w18010 & ~w18703;
assign w9582 = ~w2157 & ~w9731;
assign w9583 = w9767 & w8261;
assign w9584 = w9327 & ~w7184;
assign w9585 = ~w544 & ~w18361;
assign w9586 = ~w13768 & ~w7069;
assign w9587 = w17989 & w727;
assign w9588 = ~w10282 & ~w15684;
assign w9589 = w15433 & w590;
assign w9590 = w16055 & ~w1632;
assign w9591 = ~w12276 & ~w447;
assign w9592 = ~w10641 & ~w10388;
assign w9593 = ~w5569 & ~w5308;
assign w9594 = ~w14314 & w860;
assign w9595 = a_0 & ~w16542;
assign w9596 = w12888 & w917;
assign w9597 = ~w12500 & ~w4716;
assign w9598 = a_8 & a_51;
assign w9599 = ~w10220 & w16286;
assign w9600 = ~w15585 & w3344;
assign w9601 = ~w14761 & w12916;
assign w9602 = ~w17379 & w3287;
assign w9603 = ~w17561 & ~w11414;
assign w9604 = a_8 & a_24;
assign w9605 = w10761 & ~w15354;
assign w9606 = ~w18245 & w4742;
assign w9607 = a_5 & a_45;
assign w9608 = ~w9248 & ~w78;
assign w9609 = ~w13541 & ~w17838;
assign w9610 = a_6 & a_62;
assign w9611 = ~w12527 & ~w16575;
assign w9612 = a_31 & a_58;
assign w9613 = ~w12591 & ~w2195;
assign w9614 = (w5560 & w9184) | (w5560 & w18511) | (w9184 & w18511);
assign w9615 = ~w14907 & ~w5931;
assign w9616 = (~w10504 & ~w7758) | (~w10504 & w3324) | (~w7758 & w3324);
assign w9617 = (w1286 & w18212) | (w1286 & w16592) | (w18212 & w16592);
assign w9618 = w6954 & w5922;
assign w9619 = w7594 & w4008;
assign w9620 = (~w2794 & w15113) | (~w2794 & w170) | (w15113 & w170);
assign w9621 = w14016 & w13772;
assign w9622 = w9304 & ~w6956;
assign w9623 = w2960 & w9932;
assign w9624 = ~w19016 & w2081;
assign w9625 = ~w174 & ~w10039;
assign w9626 = (~w14709 & ~w17422) | (~w14709 & w10836) | (~w17422 & w10836);
assign w9627 = ~w2319 & ~w6705;
assign w9628 = w18821 & w804;
assign w9629 = ~w18343 & ~w2669;
assign w9630 = a_19 & a_25;
assign w9631 = ~w14468 & ~w14883;
assign w9632 = ~w16726 & w17113;
assign w9633 = w10796 & ~w14298;
assign w9634 = (~w14672 & ~w675) | (~w14672 & w3278) | (~w675 & w3278);
assign w9635 = ~w769 & ~w11098;
assign w9636 = w4766 & w5971;
assign w9637 = ~w17962 & ~w3242;
assign w9638 = (~w1734 & w6982) | (~w1734 & w602) | (w6982 & w602);
assign w9639 = w13217 & ~w1268;
assign w9640 = ~w18125 & ~w6205;
assign w9641 = w5074 & ~w1786;
assign w9642 = w18027 & ~w2000;
assign w9643 = ~w16398 & w14288;
assign w9644 = ~w7722 & w15625;
assign w9645 = ~w14067 & ~w10274;
assign w9646 = w15663 & ~w9916;
assign w9647 = ~w14798 & ~w18925;
assign w9648 = (~w5084 & ~w18488) | (~w5084 & w5854) | (~w18488 & w5854);
assign w9649 = ~w6183 & ~w12504;
assign w9650 = ~w15496 & ~w9287;
assign w9651 = (~w788 & ~w12946) | (~w788 & w8478) | (~w12946 & w8478);
assign w9652 = w3062 & w4849;
assign w9653 = ~w2664 & ~w11836;
assign w9654 = ~w8085 & ~w18479;
assign w9655 = ~w3045 & ~w7174;
assign w9656 = ~w13993 & ~w13272;
assign w9657 = a_11 & a_32;
assign w9658 = ~w13353 & ~w9721;
assign w9659 = w2172 & w18221;
assign w9660 = w3468 & w2328;
assign w9661 = (~w3670 & ~w17643) | (~w3670 & w18123) | (~w17643 & w18123);
assign w9662 = w4278 & w7589;
assign w9663 = ~w15155 & ~w11238;
assign w9664 = ~w6759 & w8328;
assign w9665 = (~w13118 & ~w4548) | (~w13118 & w1236) | (~w4548 & w1236);
assign w9666 = (a_58 & w1016) | (a_58 & w10527) | (w1016 & w10527);
assign w9667 = w2707 & w13167;
assign w9668 = (w1566 & w2903) | (w1566 & w299) | (w2903 & w299);
assign w9669 = ~w3487 & w11020;
assign w9670 = ~w4940 & ~w909;
assign w9671 = ~w11649 & ~w16333;
assign w9672 = ~w11506 & ~w777;
assign w9673 = a_23 & a_27;
assign w9674 = ~w191 & ~w15232;
assign w9675 = (~w502 & ~w14140) | (~w502 & w1277) | (~w14140 & w1277);
assign w9676 = w2133 & ~w781;
assign w9677 = a_2 & a_33;
assign w9678 = w10100 & w12476;
assign w9679 = a_11 & a_21;
assign w9680 = ~w9096 & ~w15733;
assign w9681 = w16843 & ~w4823;
assign w9682 = ~w3877 & w11913;
assign w9683 = w17162 & ~w17962;
assign w9684 = ~w82 & ~w11508;
assign w9685 = ~w3570 & ~w3190;
assign w9686 = ~w243 & w11760;
assign w9687 = w11742 & w6834;
assign w9688 = a_7 & a_8;
assign w9689 = w8552 & ~w898;
assign w9690 = w8201 & ~w1323;
assign w9691 = a_4 & a_22;
assign w9692 = a_56 & a_62;
assign w9693 = ~w6824 & ~w16208;
assign w9694 = ~w11108 & w9354;
assign w9695 = w3695 & ~w11656;
assign w9696 = ~w3063 & ~w15323;
assign w9697 = ~w16518 & ~w2425;
assign w9698 = (~w16653 & ~w9774) | (~w16653 & w3037) | (~w9774 & w3037);
assign w9699 = ~w1719 & w2278;
assign w9700 = a_32 & a_53;
assign w9701 = ~w5694 & ~w12147;
assign w9702 = w19101 & w4247;
assign w9703 = ~w626 & ~w19035;
assign w9704 = a_19 & a_24;
assign w9705 = ~w3488 & ~w16431;
assign w9706 = w2844 & w19168;
assign w9707 = a_31 & a_40;
assign w9708 = w14531 & ~w18622;
assign w9709 = w8842 & w11700;
assign w9710 = ~w19130 & ~w13918;
assign w9711 = ~w16478 & ~w14090;
assign w9712 = ~w15673 & ~w16649;
assign w9713 = ~w10452 & ~w15136;
assign w9714 = w11323 & w10631;
assign w9715 = ~w9809 & ~w2153;
assign w9716 = ~w7097 & ~w13488;
assign w9717 = ~w9824 & w10279;
assign w9718 = (w7102 & w3910) | (w7102 & w13663) | (w3910 & w13663);
assign w9719 = ~w12390 & w6866;
assign w9720 = ~w9922 & ~w1634;
assign w9721 = ~w3990 & ~w18434;
assign w9722 = ~w14759 & ~w9083;
assign w9723 = w2562 & ~w13917;
assign w9724 = ~w13731 & ~w14888;
assign w9725 = ~w12161 & ~w13414;
assign w9726 = ~w5919 & w2329;
assign w9727 = w7058 & w2241;
assign w9728 = a_20 & a_23;
assign w9729 = a_3 & a_9;
assign w9730 = (w3232 & w545) | (w3232 & w1074) | (w545 & w1074);
assign w9731 = ~w2431 & w12360;
assign w9732 = ~w2666 & w17329;
assign w9733 = w18437 & ~w9957;
assign w9734 = ~w6082 & ~w3056;
assign w9735 = ~w12081 & ~w478;
assign w9736 = ~w622 & ~w7218;
assign w9737 = w17706 & w13487;
assign w9738 = ~w7918 & ~w7042;
assign w9739 = w6883 & ~w15707;
assign w9740 = ~w11698 & w18492;
assign w9741 = ~w18717 & ~w12543;
assign w9742 = a_29 & a_54;
assign w9743 = ~w5786 & ~w12581;
assign w9744 = ~w10957 & ~w11521;
assign w9745 = w11385 & w12266;
assign w9746 = w1810 & ~w10718;
assign w9747 = ~w3985 & w16842;
assign w9748 = w10699 & w8243;
assign w9749 = ~w4617 & ~w3730;
assign w9750 = ~w7181 & ~w13128;
assign w9751 = ~w8166 & w18785;
assign w9752 = w6543 & ~w10216;
assign w9753 = ~w1994 & ~w13714;
assign w9754 = ~w15760 & ~w2284;
assign w9755 = (~w2051 & ~w8873) | (~w2051 & w1023) | (~w8873 & w1023);
assign w9756 = ~w18160 & ~w8720;
assign w9757 = w13522 & w10121;
assign w9758 = ~w3080 & w18687;
assign w9759 = ~w4607 & ~w5884;
assign w9760 = ~w10440 & ~w17910;
assign w9761 = ~w8360 & ~w6217;
assign w9762 = w11781 & w3332;
assign w9763 = ~w4962 & ~w9933;
assign w9764 = (w8240 & w2254) | (w8240 & w16164) | (w2254 & w16164);
assign w9765 = w4035 & ~w5205;
assign w9766 = ~w6531 & ~w18889;
assign w9767 = ~w11816 & ~w13560;
assign w9768 = a_28 & a_29;
assign w9769 = ~w3861 & ~w11398;
assign w9770 = ~w1319 & ~w9140;
assign w9771 = ~w18051 & ~w6706;
assign w9772 = w15052 & w5621;
assign w9773 = ~w18339 & ~w16157;
assign w9774 = ~w16653 & ~w5129;
assign w9775 = w14920 & ~w7412;
assign w9776 = w8471 & ~w4357;
assign w9777 = w9742 & ~w10659;
assign w9778 = ~w10991 & w10745;
assign w9779 = w17116 & w11273;
assign w9780 = w8532 & ~w18421;
assign w9781 = ~w15449 & ~w1622;
assign w9782 = ~w15674 & w4567;
assign w9783 = ~w10710 & ~w7624;
assign w9784 = ~w2485 & ~w16490;
assign w9785 = ~w14614 & ~w14400;
assign w9786 = ~w15123 & w14013;
assign w9787 = w4512 & w5847;
assign w9788 = ~w14151 & w12216;
assign w9789 = a_32 & a_61;
assign w9790 = w403 & w15928;
assign w9791 = w1313 & ~w19139;
assign w9792 = ~w5355 & ~w121;
assign w9793 = ~w18624 & ~w4460;
assign w9794 = ~w1939 & ~w14255;
assign w9795 = ~w9425 & w8123;
assign w9796 = (w1452 & ~w6617) | (w1452 & w18987) | (~w6617 & w18987);
assign w9797 = (w10390 & w5107) | (w10390 & w17140) | (w5107 & w17140);
assign w9798 = (a_61 & w8243) | (a_61 & w5964) | (w8243 & w5964);
assign w9799 = ~w18980 & ~w2464;
assign w9800 = ~w16161 & ~w17699;
assign w9801 = ~w14486 & w7388;
assign w9802 = ~w1303 & ~w8220;
assign w9803 = a_27 & a_34;
assign w9804 = ~w4896 & w14654;
assign w9805 = ~w953 & ~w4981;
assign w9806 = w2524 & w6396;
assign w9807 = (~w6215 & ~w6767) | (~w6215 & w1075) | (~w6767 & w1075);
assign w9808 = ~w7948 & ~w10674;
assign w9809 = ~w9998 & ~w2407;
assign w9810 = w18980 & ~w11689;
assign w9811 = ~w9914 & w13920;
assign w9812 = ~w13689 & ~w3;
assign w9813 = ~w12758 & ~w190;
assign w9814 = ~w7794 & ~w15462;
assign w9815 = ~w567 & w7170;
assign w9816 = w16646 & w7741;
assign w9817 = ~w16131 & ~w259;
assign w9818 = w6853 & w19005;
assign w9819 = ~w1256 & ~w14099;
assign w9820 = ~w18974 & ~w9510;
assign w9821 = ~w1048 & w4951;
assign w9822 = ~w3978 & w16476;
assign w9823 = ~w11601 & w18770;
assign w9824 = a_21 & a_36;
assign w9825 = ~w13875 & ~w2589;
assign w9826 = w5696 & w3156;
assign w9827 = w4749 & w16363;
assign w9828 = ~w2868 & w10550;
assign w9829 = ~w5874 & ~w3706;
assign w9830 = w13116 & w14778;
assign w9831 = ~w1280 & ~w16962;
assign w9832 = (~w14011 & ~w2979) | (~w14011 & w19127) | (~w2979 & w19127);
assign w9833 = ~w5488 & ~w15305;
assign w9834 = a_5 & a_44;
assign w9835 = (~w14545 & ~w12050) | (~w14545 & w4794) | (~w12050 & w4794);
assign w9836 = ~w3334 & w12856;
assign w9837 = a_7 & a_14;
assign w9838 = ~w98 & ~w4978;
assign w9839 = ~w12819 & ~w1669;
assign w9840 = ~w18491 & ~w17266;
assign w9841 = ~w19031 & ~w14338;
assign w9842 = w18777 & w136;
assign w9843 = a_6 & a_7;
assign w9844 = ~w12537 & ~w15725;
assign w9845 = ~w1173 & w10144;
assign w9846 = w3036 & ~w10889;
assign w9847 = (w17101 & ~w13830) | (w17101 & w4066) | (~w13830 & w4066);
assign w9848 = a_5 & a_41;
assign w9849 = w13450 & w995;
assign w9850 = ~w3599 & ~w8976;
assign w9851 = ~w6241 & ~w1953;
assign w9852 = w13480 & w11164;
assign w9853 = ~w5124 & ~w7845;
assign w9854 = a_46 & a_56;
assign w9855 = ~w11277 & w5824;
assign w9856 = ~w2060 & w454;
assign w9857 = ~w5384 & ~w1835;
assign w9858 = a_46 & a_47;
assign w9859 = ~w899 & ~w14108;
assign w9860 = w6021 & ~w7035;
assign w9861 = w1018 & ~w10430;
assign w9862 = w4050 & w7306;
assign w9863 = ~w3985 & w11351;
assign w9864 = ~w6431 & w11603;
assign w9865 = ~w16287 & ~w2926;
assign w9866 = ~w9627 & ~w12838;
assign w9867 = ~w11291 & w1509;
assign w9868 = ~w17662 & ~w10226;
assign w9869 = (w1290 & w10330) | (w1290 & w54) | (w10330 & w54);
assign w9870 = ~w5742 & ~w17746;
assign w9871 = ~w11789 & w7946;
assign w9872 = ~w9540 & ~w4061;
assign w9873 = ~w13165 & ~w10638;
assign w9874 = w18176 & w7737;
assign w9875 = ~w15188 & w10600;
assign w9876 = ~w1106 & ~w4510;
assign w9877 = ~w5264 & ~w11480;
assign w9878 = w16793 & ~w15526;
assign w9879 = w11281 & ~w5906;
assign w9880 = ~w18466 & ~w14760;
assign w9881 = ~w2406 & ~w16323;
assign w9882 = a_30 & a_40;
assign w9883 = a_32 & a_54;
assign w9884 = w4296 & ~w18720;
assign w9885 = a_23 & a_47;
assign w9886 = w8198 & ~w11218;
assign w9887 = ~w2808 & ~w1347;
assign w9888 = ~w1979 & ~w12778;
assign w9889 = ~w7434 & ~w6161;
assign w9890 = w1138 & ~w14825;
assign w9891 = w6187 & ~w14960;
assign w9892 = w2684 & ~w17433;
assign w9893 = w19053 & w19169;
assign w9894 = ~w17918 & ~w2236;
assign w9895 = ~w13323 & ~w16217;
assign w9896 = ~w17277 & ~w2238;
assign w9897 = a_52 & a_57;
assign w9898 = ~w5625 & ~w6490;
assign w9899 = ~w1951 & w4791;
assign w9900 = ~w3054 & ~w14410;
assign w9901 = ~w16323 & ~w8047;
assign w9902 = (w1566 & w11733) | (w1566 & w8322) | (w11733 & w8322);
assign w9903 = ~w8510 & ~w15143;
assign w9904 = ~w1328 & ~w2451;
assign w9905 = (~w2769 & w11636) | (~w2769 & w17881) | (w11636 & w17881);
assign w9906 = ~w6117 & w4762;
assign w9907 = w5545 & ~w57;
assign w9908 = w14248 & w4163;
assign w9909 = ~w17411 & ~w12434;
assign w9910 = w7022 & w1419;
assign w9911 = ~w8974 & w19147;
assign w9912 = ~w17937 & ~w7371;
assign w9913 = a_9 & a_53;
assign w9914 = a_18 & a_60;
assign w9915 = ~w12465 & w13598;
assign w9916 = ~w3950 & ~w16181;
assign w9917 = a_54 & w5867;
assign w9918 = w12751 & ~w5695;
assign w9919 = ~w17618 & ~w8081;
assign w9920 = ~w19114 & ~w614;
assign w9921 = ~w12452 & w5234;
assign w9922 = ~w17745 & ~w17059;
assign w9923 = ~w18538 & ~w6949;
assign w9924 = ~w4970 & w1919;
assign w9925 = ~w15799 & ~w7901;
assign w9926 = (~w3336 & ~w9048) | (~w3336 & w14782) | (~w9048 & w14782);
assign w9927 = ~w15759 & ~w6916;
assign w9928 = w7732 & ~w18664;
assign w9929 = w4800 & w18517;
assign w9930 = ~w13115 & ~w15028;
assign w9931 = w5193 & ~w6885;
assign w9932 = ~w4170 & w9418;
assign w9933 = ~w2190 & ~w6;
assign w9934 = w5694 & w12147;
assign w9935 = w3928 & w17890;
assign w9936 = w13476 & ~w14357;
assign w9937 = a_31 & w13854;
assign w9938 = a_17 & a_51;
assign w9939 = ~w15261 & ~w3970;
assign w9940 = ~w7317 & ~w1303;
assign w9941 = w1100 & ~w4212;
assign w9942 = ~w18895 & ~w11341;
assign w9943 = (~w3619 & ~w10496) | (~w3619 & w15565) | (~w10496 & w15565);
assign w9944 = ~w17483 & w19113;
assign w9945 = (w6636 & w15543) | (w6636 & w10537) | (w15543 & w10537);
assign w9946 = w15669 & ~w5607;
assign w9947 = ~w16786 & ~w13899;
assign w9948 = (~w16418 & ~w10180) | (~w16418 & w10780) | (~w10180 & w10780);
assign w9949 = w11628 & w17447;
assign w9950 = (w14339 & w1638) | (w14339 & w16742) | (w1638 & w16742);
assign w9951 = ~w3472 & ~w13891;
assign w9952 = ~w3217 & ~w3611;
assign w9953 = ~w10349 & w14886;
assign w9954 = a_20 & a_59;
assign w9955 = ~w18258 & ~w18897;
assign w9956 = w1452 & ~w3415;
assign w9957 = ~w8538 & ~w13916;
assign w9958 = w4804 & ~w13287;
assign w9959 = (~w9113 & w7017) | (~w9113 & w4235) | (w7017 & w4235);
assign w9960 = w18671 & w10838;
assign w9961 = a_11 & a_54;
assign w9962 = ~a_46 & a_47;
assign w9963 = ~w8963 & ~w3387;
assign w9964 = ~w79 & ~w14554;
assign w9965 = w824 & ~w13673;
assign w9966 = w15289 & ~w718;
assign w9967 = ~w8619 & ~w10929;
assign w9968 = w14364 & ~w15352;
assign w9969 = ~w13240 & ~w2098;
assign w9970 = ~w19110 & w10556;
assign w9971 = w1553 & w15975;
assign w9972 = w9336 & ~w17249;
assign w9973 = w14646 & w15691;
assign w9974 = ~w14718 & ~w9685;
assign w9975 = ~w2963 & w17533;
assign w9976 = w1673 & ~w12680;
assign w9977 = a_5 & a_35;
assign w9978 = ~w14055 & ~w701;
assign w9979 = ~w14074 & ~w2635;
assign w9980 = ~w22 & ~w11171;
assign w9981 = ~w11454 & w4113;
assign w9982 = ~w3598 & ~w11974;
assign w9983 = ~w6859 & ~w18771;
assign w9984 = ~w18253 & ~w13088;
assign w9985 = ~w10702 & ~w5662;
assign w9986 = a_5 & a_47;
assign w9987 = ~w18736 & ~w266;
assign w9988 = ~w12442 & ~w7003;
assign w9989 = a_28 & a_55;
assign w9990 = ~w9844 & ~w6173;
assign w9991 = w10339 & ~w16645;
assign w9992 = ~w16550 & ~w10451;
assign w9993 = ~w16236 & w9611;
assign w9994 = w9008 & ~w1598;
assign w9995 = (~w8206 & ~w10282) | (~w8206 & w4581) | (~w10282 & w4581);
assign w9996 = a_12 & a_15;
assign w9997 = w13163 & ~w16663;
assign w9998 = w17340 & w8894;
assign w9999 = a_3 & a_53;
assign w10000 = w16200 & w15983;
assign w10001 = w481 & ~w10962;
assign w10002 = ~w16472 & ~w18057;
assign w10003 = ~w7666 & ~w11342;
assign w10004 = ~w2402 & ~w13590;
assign w10005 = ~w3269 & ~w15747;
assign w10006 = w14530 & ~w1956;
assign w10007 = w3669 & w12405;
assign w10008 = a_46 & a_60;
assign w10009 = ~w5605 & ~w13162;
assign w10010 = (~w13964 & ~w7590) | (~w13964 & w15690) | (~w7590 & w15690);
assign w10011 = w18845 & ~w18940;
assign w10012 = w18688 & ~w473;
assign w10013 = ~w17347 & ~w185;
assign w10014 = (a_47 & w13290) | (a_47 & w9858) | (w13290 & w9858);
assign w10015 = ~w16699 & ~w16596;
assign w10016 = (~w2769 & w12413) | (~w2769 & w4040) | (w12413 & w4040);
assign w10017 = w5715 & ~w3342;
assign w10018 = w11812 & w12442;
assign w10019 = ~w9045 & w4000;
assign w10020 = ~w504 & ~w16893;
assign w10021 = (w8802 & w3696) | (w8802 & w12484) | (w3696 & w12484);
assign w10022 = w14771 & ~w4524;
assign w10023 = ~w13008 & w13770;
assign w10024 = ~w18381 & ~w10063;
assign w10025 = ~w329 & ~w13058;
assign w10026 = ~w916 & w17241;
assign w10027 = (~w10375 & w3437) | (~w10375 & w12866) | (w3437 & w12866);
assign w10028 = w3068 & w13462;
assign w10029 = ~w13377 & ~w15880;
assign w10030 = a_37 & a_50;
assign w10031 = ~w16389 & w8171;
assign w10032 = ~w11565 & ~w1744;
assign w10033 = a_42 & a_46;
assign w10034 = w11336 & ~w579;
assign w10035 = ~w10616 & w9933;
assign w10036 = ~w3992 & ~w6064;
assign w10037 = a_23 & a_49;
assign w10038 = ~w13214 & ~w11446;
assign w10039 = ~w6738 & w2014;
assign w10040 = w7494 & ~w16259;
assign w10041 = w9854 & w3250;
assign w10042 = a_9 & a_19;
assign w10043 = ~w3935 & ~w2377;
assign w10044 = ~w18579 & ~w5442;
assign w10045 = w14613 & w15903;
assign w10046 = ~w17665 & w2239;
assign w10047 = a_29 & a_32;
assign w10048 = ~w12165 & ~w14119;
assign w10049 = ~w7251 & ~w322;
assign w10050 = ~w17994 & w7233;
assign w10051 = (~w17294 & w10330) | (~w17294 & w7497) | (w10330 & w7497);
assign w10052 = a_9 & a_52;
assign w10053 = a_20 & a_46;
assign w10054 = ~w17585 & w4748;
assign w10055 = a_1 & a_20;
assign w10056 = ~w2356 & ~w635;
assign w10057 = ~w13344 & ~w1472;
assign w10058 = ~w10607 & ~w1518;
assign w10059 = a_8 & a_36;
assign w10060 = w13484 & ~w4236;
assign w10061 = ~w2795 & ~w7040;
assign w10062 = ~w14715 & w5374;
assign w10063 = ~w9466 & ~w8845;
assign w10064 = ~w18495 & w18474;
assign w10065 = ~w18033 & ~w3379;
assign w10066 = ~w17943 & ~w15932;
assign w10067 = w4113 & ~w10170;
assign w10068 = ~w5809 & ~w10790;
assign w10069 = (~w10334 & ~w16741) | (~w10334 & w13996) | (~w16741 & w13996);
assign w10070 = w1286 & ~w11855;
assign w10071 = w8866 & w854;
assign w10072 = ~w1004 & ~w18827;
assign w10073 = ~w16998 & ~w11070;
assign w10074 = ~w17409 & ~w7082;
assign w10075 = w7517 & w6163;
assign w10076 = ~w7301 & ~w6471;
assign w10077 = ~w5463 & w14207;
assign w10078 = w14789 & ~w14802;
assign w10079 = ~w11539 & ~w6499;
assign w10080 = ~w7214 & w14393;
assign w10081 = w13246 & w15803;
assign w10082 = ~w11254 & ~w689;
assign w10083 = a_3 & a_41;
assign w10084 = ~w14564 & ~w1886;
assign w10085 = ~w17335 & ~w4222;
assign w10086 = ~w5223 & ~w13260;
assign w10087 = ~w17767 & ~w11929;
assign w10088 = ~w16840 & ~w6053;
assign w10089 = ~w16639 & w9161;
assign w10090 = ~w1167 & ~w17414;
assign w10091 = ~w1062 & w4313;
assign w10092 = ~w10724 & ~w17862;
assign w10093 = ~w17967 & ~w6191;
assign w10094 = w815 & ~w15765;
assign w10095 = a_43 & a_61;
assign w10096 = (~w19005 & w487) | (~w19005 & w6762) | (w487 & w6762);
assign w10097 = w11065 & w6895;
assign w10098 = ~w5715 & ~w3049;
assign w10099 = ~w7610 & w3293;
assign w10100 = ~w14004 & ~w6203;
assign w10101 = w9749 & ~w3088;
assign w10102 = ~w11891 & ~w6227;
assign w10103 = ~w12925 & ~w1254;
assign w10104 = a_52 & a_63;
assign w10105 = (~w12187 & ~w4303) | (~w12187 & w12379) | (~w4303 & w12379);
assign w10106 = ~w17444 & w11367;
assign w10107 = ~w6973 & ~w7625;
assign w10108 = a_42 & a_50;
assign w10109 = ~w6455 & ~w397;
assign w10110 = ~w10987 & ~w7467;
assign w10111 = ~w7329 & w5835;
assign w10112 = ~w3998 & ~w5447;
assign w10113 = ~w8826 & ~w2670;
assign w10114 = w838 & w1504;
assign w10115 = w13268 & w10930;
assign w10116 = ~w13621 & w18629;
assign w10117 = w13589 & w853;
assign w10118 = ~w9340 & w2222;
assign w10119 = ~w13571 & ~w3673;
assign w10120 = w9449 & ~w4318;
assign w10121 = a_3 & a_50;
assign w10122 = ~w394 & ~w8214;
assign w10123 = ~w1978 & ~w7642;
assign w10124 = ~w7289 & w8440;
assign w10125 = ~w884 & ~w3249;
assign w10126 = ~w12769 & ~w6256;
assign w10127 = w10179 & w630;
assign w10128 = ~w3119 & w801;
assign w10129 = w7962 & ~w5565;
assign w10130 = ~w14511 & ~w8092;
assign w10131 = ~w18884 & w17861;
assign w10132 = ~w9945 & ~w13415;
assign w10133 = ~w16151 & w16265;
assign w10134 = ~w12090 & ~w8749;
assign w10135 = w8641 & ~w143;
assign w10136 = w17842 & ~w14634;
assign w10137 = ~w16082 & ~w15521;
assign w10138 = a_0 & a_49;
assign w10139 = ~w15573 & ~w10087;
assign w10140 = a_24 & a_59;
assign w10141 = ~a_53 & a_54;
assign w10142 = ~w8499 & ~w16897;
assign w10143 = w12508 & ~w714;
assign w10144 = ~w2520 & ~w14485;
assign w10145 = w19086 & w7586;
assign w10146 = (~w12904 & w175) | (~w12904 & w18074) | (w175 & w18074);
assign w10147 = ~w7507 & ~w12183;
assign w10148 = w10193 & w17593;
assign w10149 = w6293 & ~w9157;
assign w10150 = a_17 & a_18;
assign w10151 = ~w1220 & ~w950;
assign w10152 = ~w9708 & w9058;
assign w10153 = ~w2911 & w3837;
assign w10154 = w18356 & w15020;
assign w10155 = ~w14530 & w7022;
assign w10156 = w5816 & ~w6322;
assign w10157 = w5688 & ~w8872;
assign w10158 = ~w2152 & ~w11237;
assign w10159 = w16868 & w18921;
assign w10160 = w11 & ~w18388;
assign w10161 = w15396 & w17677;
assign w10162 = w14978 & w6043;
assign w10163 = w12317 & ~w17184;
assign w10164 = w18564 & ~w14320;
assign w10165 = ~w5352 & w17141;
assign w10166 = ~w11416 & w17433;
assign w10167 = ~w4088 & ~w6192;
assign w10168 = w18636 & ~w1294;
assign w10169 = ~w16793 & w15526;
assign w10170 = w5825 & ~w9876;
assign w10171 = ~w8580 & w1451;
assign w10172 = ~w2460 & ~w16435;
assign w10173 = ~w4344 & ~w12901;
assign w10174 = w16087 & ~w4335;
assign w10175 = w6585 & ~w12270;
assign w10176 = ~w6241 & ~w15581;
assign w10177 = w1408 & ~w4276;
assign w10178 = ~w10197 & ~w13471;
assign w10179 = ~w4884 & ~w10060;
assign w10180 = ~w16418 & ~w12432;
assign w10181 = ~w16042 & ~w15955;
assign w10182 = ~w15185 & ~w8591;
assign w10183 = ~w1426 & ~w17730;
assign w10184 = w9020 & ~w16999;
assign w10185 = w11117 & ~w18092;
assign w10186 = ~w9116 & ~w346;
assign w10187 = a_0 & a_5;
assign w10188 = ~w18764 & w2357;
assign w10189 = ~w15605 & ~w13952;
assign w10190 = ~w10538 & w6938;
assign w10191 = ~w14218 & w5069;
assign w10192 = ~w15072 & ~w2967;
assign w10193 = a_0 & a_60;
assign w10194 = ~w2834 & ~w11789;
assign w10195 = w14940 & w2273;
assign w10196 = ~w5258 & w11715;
assign w10197 = ~w15739 & ~w2498;
assign w10198 = ~w63 & w5361;
assign w10199 = ~w8710 & ~w9961;
assign w10200 = (~w3047 & ~w17052) | (~w3047 & w7376) | (~w17052 & w7376);
assign w10201 = ~w12726 & w218;
assign w10202 = w9131 & ~w2798;
assign w10203 = a_31 & a_45;
assign w10204 = w10580 & ~w11380;
assign w10205 = ~w2046 & ~w9724;
assign w10206 = ~w7555 & ~w8539;
assign w10207 = w12648 & ~w2184;
assign w10208 = (~w6069 & ~w6002) | (~w6069 & w660) | (~w6002 & w660);
assign w10209 = (~w8437 & w17734) | (~w8437 & w19170) | (w17734 & w19170);
assign w10210 = ~w7863 & w2454;
assign w10211 = ~w7945 & ~w9783;
assign w10212 = ~w18689 & ~w17269;
assign w10213 = w13224 & w13346;
assign w10214 = a_33 & a_57;
assign w10215 = w7566 & ~w13452;
assign w10216 = ~w14451 & ~w6749;
assign w10217 = w14297 & ~w4303;
assign w10218 = ~w16435 & ~w8372;
assign w10219 = w13350 & w15325;
assign w10220 = ~w15374 & ~w3552;
assign w10221 = w17099 & ~w5851;
assign w10222 = w5367 & w5192;
assign w10223 = a_15 & a_49;
assign w10224 = ~w10968 & w6774;
assign w10225 = a_14 & a_31;
assign w10226 = w15025 & ~w16621;
assign w10227 = ~w14294 & w4945;
assign w10228 = ~w5366 & ~w18352;
assign w10229 = a_36 & a_46;
assign w10230 = ~w156 & ~w5443;
assign w10231 = (~w12370 & w6679) | (~w12370 & w7889) | (w6679 & w7889);
assign w10232 = a_63 & ~w2659;
assign w10233 = w1475 & ~w16667;
assign w10234 = a_21 & a_50;
assign w10235 = ~w7252 & ~w8638;
assign w10236 = ~w2569 & ~w5965;
assign w10237 = (w8340 & w2929) | (w8340 & w2128) | (w2929 & w2128);
assign w10238 = ~w2665 & ~w5923;
assign w10239 = ~w5659 & ~w2982;
assign w10240 = ~w1103 & w9832;
assign w10241 = ~w11600 & ~w16104;
assign w10242 = w17513 & w15386;
assign w10243 = a_52 & w5112;
assign w10244 = ~w1170 & ~w13417;
assign w10245 = ~w11826 & ~w14504;
assign w10246 = w1855 & w326;
assign w10247 = ~w17058 & ~w13760;
assign w10248 = w17360 & ~w7075;
assign w10249 = w3125 & ~w16335;
assign w10250 = ~w3353 & ~w14427;
assign w10251 = w10581 & ~w18153;
assign w10252 = w11309 & w15501;
assign w10253 = (~w10003 & ~w8357) | (~w10003 & w16524) | (~w8357 & w16524);
assign w10254 = ~w15195 & ~w12176;
assign w10255 = w15338 & w18941;
assign w10256 = ~w15698 & w9773;
assign w10257 = ~w896 & ~w13297;
assign w10258 = ~w10140 & ~w7932;
assign w10259 = ~w18752 & ~w7706;
assign w10260 = ~w4691 & w3262;
assign w10261 = ~w13644 & ~w3673;
assign w10262 = a_18 & a_55;
assign w10263 = w11779 & ~w15559;
assign w10264 = ~w14900 & ~w6286;
assign w10265 = ~w13381 & w8045;
assign w10266 = (w1576 & w7610) | (w1576 & w2399) | (w7610 & w2399);
assign w10267 = ~w2258 & ~w17083;
assign w10268 = ~w12839 & w4541;
assign w10269 = a_22 & a_48;
assign w10270 = ~w5016 & ~w6209;
assign w10271 = ~w5327 & ~w7171;
assign w10272 = ~w8088 & w14984;
assign w10273 = w14644 & w9985;
assign w10274 = ~w698 & ~w17882;
assign w10275 = ~w9596 & ~w3595;
assign w10276 = a_43 & a_59;
assign w10277 = ~w12397 & ~w17789;
assign w10278 = w11355 & w5903;
assign w10279 = ~w6075 & ~w2074;
assign w10280 = w15010 & ~w9127;
assign w10281 = ~w2838 & w8068;
assign w10282 = ~w8206 & ~w6509;
assign w10283 = w12266 & w16423;
assign w10284 = ~w9348 & ~w14795;
assign w10285 = ~w1107 & ~w5665;
assign w10286 = w14921 & w2884;
assign w10287 = ~w5716 & ~w13386;
assign w10288 = ~w8029 & w19136;
assign w10289 = w3866 & w18208;
assign w10290 = a_15 & a_45;
assign w10291 = a_24 & a_26;
assign w10292 = (~w10897 & ~w14929) | (~w10897 & w589) | (~w14929 & w589);
assign w10293 = w8258 & ~w4287;
assign w10294 = ~w964 & ~w7640;
assign w10295 = ~w12835 & ~w11963;
assign w10296 = w10704 & w11734;
assign w10297 = a_17 & a_27;
assign w10298 = a_29 & a_56;
assign w10299 = (w9058 & ~w14949) | (w9058 & w10152) | (~w14949 & w10152);
assign w10300 = ~w15207 & ~w10159;
assign w10301 = ~w9049 & ~w10187;
assign w10302 = a_40 & a_44;
assign w10303 = ~w551 & ~w5918;
assign w10304 = ~w16191 & w15781;
assign w10305 = ~w8620 & ~w16443;
assign w10306 = ~w11965 & w10958;
assign w10307 = ~w13294 & w17037;
assign w10308 = w3381 & w12184;
assign w10309 = ~w12113 & ~w13411;
assign w10310 = ~w2755 & ~w4761;
assign w10311 = ~w8069 & ~w16098;
assign w10312 = a_34 & a_47;
assign w10313 = w7316 & w5031;
assign w10314 = ~w2880 & w14280;
assign w10315 = a_8 & a_62;
assign w10316 = a_20 & a_33;
assign w10317 = a_30 & a_52;
assign w10318 = ~w11365 & ~w14854;
assign w10319 = ~w14889 & ~w10989;
assign w10320 = ~w16609 & ~w17219;
assign w10321 = ~w13350 & ~w15325;
assign w10322 = w3883 & w12497;
assign w10323 = ~w8212 & ~w9755;
assign w10324 = ~w13589 & ~w3034;
assign w10325 = ~w16944 & ~w17731;
assign w10326 = ~w4670 & ~w10872;
assign w10327 = ~w4005 & w11842;
assign w10328 = ~w7970 & ~w6088;
assign w10329 = ~w96 & ~w16315;
assign w10330 = (w7920 & w9221) | (w7920 & w8455) | (w9221 & w8455);
assign w10331 = ~w2297 & ~w6672;
assign w10332 = w12332 & w10489;
assign w10333 = ~w14441 & ~w16032;
assign w10334 = ~w14153 & ~w9495;
assign w10335 = w14308 & ~w4920;
assign w10336 = ~w18315 & ~w7832;
assign w10337 = w10614 & ~w14850;
assign w10338 = ~w2766 & ~w9167;
assign w10339 = ~w10139 & ~w11221;
assign w10340 = ~w8743 & ~w15465;
assign w10341 = ~w19011 & ~w6907;
assign w10342 = ~w1759 & w3480;
assign w10343 = w9362 & w14290;
assign w10344 = ~w3809 & ~w1649;
assign w10345 = (~w2178 & ~w10624) | (~w2178 & w12044) | (~w10624 & w12044);
assign w10346 = w2778 & w17041;
assign w10347 = ~w2084 & ~w15471;
assign w10348 = w10666 & ~w9213;
assign w10349 = ~w10155 & w1558;
assign w10350 = a_46 & a_52;
assign w10351 = w15456 & ~w12563;
assign w10352 = w13597 & ~w12626;
assign w10353 = ~w14199 & ~w7858;
assign w10354 = ~w8957 & ~w5101;
assign w10355 = ~w7881 & ~w7309;
assign w10356 = a_40 & a_59;
assign w10357 = ~w17355 & ~w19106;
assign w10358 = ~w13367 & ~w13866;
assign w10359 = ~w14087 & ~w963;
assign w10360 = ~w11642 & ~w18632;
assign w10361 = ~w1601 & w17859;
assign w10362 = ~w1163 & ~w18043;
assign w10363 = a_31 & a_57;
assign w10364 = ~w9819 & w8340;
assign w10365 = ~w2557 & w14115;
assign w10366 = a_32 & a_39;
assign w10367 = ~w4635 & ~w16504;
assign w10368 = w4411 & ~w15140;
assign w10369 = ~w18127 & w10212;
assign w10370 = ~w10075 & w18243;
assign w10371 = ~w12679 & w13870;
assign w10372 = ~w1299 & w17376;
assign w10373 = ~w8516 & ~w9190;
assign w10374 = a_7 & a_63;
assign w10375 = w13472 & w2601;
assign w10376 = ~w12487 & ~w6178;
assign w10377 = w424 & w16876;
assign w10378 = ~w6259 & w6691;
assign w10379 = ~w7949 & w18338;
assign w10380 = w11057 & ~w13797;
assign w10381 = w15541 & ~w13994;
assign w10382 = ~w16101 & ~w15744;
assign w10383 = a_15 & a_59;
assign w10384 = (~w10753 & ~w14349) | (~w10753 & w15049) | (~w14349 & w15049);
assign w10385 = ~w17581 & ~w9701;
assign w10386 = w4390 & w4144;
assign w10387 = w16280 & w5870;
assign w10388 = w680 & w13526;
assign w10389 = a_61 & a_63;
assign w10390 = ~w10073 & ~w14933;
assign w10391 = ~w17555 & ~w4531;
assign w10392 = ~w13367 & ~w6424;
assign w10393 = a_10 & a_45;
assign w10394 = ~w16338 & w6135;
assign w10395 = w1194 & ~w11892;
assign w10396 = w6912 & w3884;
assign w10397 = ~w9695 & w13037;
assign w10398 = ~a_29 & ~w2151;
assign w10399 = w17899 & ~w7379;
assign w10400 = ~w2910 & ~w8335;
assign w10401 = w10983 & w4496;
assign w10402 = w8718 & ~w650;
assign w10403 = ~w6723 & w2760;
assign w10404 = ~w17351 & ~w13823;
assign w10405 = ~w11645 & ~w1606;
assign w10406 = w11235 & w16883;
assign w10407 = w14744 & w1555;
assign w10408 = ~w19102 & w17667;
assign w10409 = ~w5165 & ~w1053;
assign w10410 = ~w14637 & ~w362;
assign w10411 = a_13 & a_23;
assign w10412 = ~w1864 & ~w10383;
assign w10413 = ~w6532 & ~w5689;
assign w10414 = ~w5577 & w12743;
assign w10415 = ~w16536 & ~w8880;
assign w10416 = w16818 & w6475;
assign w10417 = ~w18422 & ~w4647;
assign w10418 = w14508 & w5836;
assign w10419 = ~w10887 & ~w1271;
assign w10420 = ~w13142 & ~w12306;
assign w10421 = ~w6285 & w18969;
assign w10422 = ~w2886 & ~w6927;
assign w10423 = ~w7564 & w4964;
assign w10424 = (w6125 & w18383) | (w6125 & w7281) | (w18383 & w7281);
assign w10425 = a_21 & a_52;
assign w10426 = a_38 & a_44;
assign w10427 = ~w3211 & ~w12458;
assign w10428 = a_49 & a_58;
assign w10429 = ~w10844 & w4857;
assign w10430 = (w5006 & w180) | (w5006 & w4397) | (w180 & w4397);
assign w10431 = w4658 & ~w2392;
assign w10432 = ~w394 & w18975;
assign w10433 = ~w6641 & w15033;
assign w10434 = ~w15387 & ~w7221;
assign w10435 = ~w4616 & ~w10310;
assign w10436 = ~w18235 & ~w2646;
assign w10437 = ~w8001 & w3601;
assign w10438 = ~w14189 & ~w2276;
assign w10439 = ~w17393 & ~w10834;
assign w10440 = w307 & ~w8434;
assign w10441 = ~w8968 & ~w11121;
assign w10442 = ~w14463 & ~w14304;
assign w10443 = w5577 & ~w12743;
assign w10444 = ~w2134 & ~w17500;
assign w10445 = ~w7866 & ~w6319;
assign w10446 = w14742 & ~w1368;
assign w10447 = ~w5555 & ~w9368;
assign w10448 = ~w4591 & ~w9553;
assign w10449 = (~w10143 & ~w7847) | (~w10143 & w17919) | (~w7847 & w17919);
assign w10450 = ~w10094 & ~w15156;
assign w10451 = ~w2722 & ~w6235;
assign w10452 = ~w870 & ~w7104;
assign w10453 = w5947 & ~w3856;
assign w10454 = ~a_59 & a_60;
assign w10455 = a_37 & a_52;
assign w10456 = a_7 & a_52;
assign w10457 = ~w11437 & ~w1084;
assign w10458 = ~w8428 & ~w14892;
assign w10459 = w2378 & ~w6637;
assign w10460 = (~w15416 & ~w7356) | (~w15416 & w3004) | (~w7356 & w3004);
assign w10461 = ~w9014 & ~w826;
assign w10462 = w12371 & w5822;
assign w10463 = w4000 & ~w3604;
assign w10464 = a_36 & a_61;
assign w10465 = ~w16053 & ~w8025;
assign w10466 = w2592 & w9271;
assign w10467 = (w7749 & ~w4092) | (w7749 & w6921) | (~w4092 & w6921);
assign w10468 = ~w2871 & ~w936;
assign w10469 = ~w4093 & ~w4669;
assign w10470 = ~w17498 & ~w4448;
assign w10471 = w13518 & ~w13103;
assign w10472 = ~w9273 & ~w1600;
assign w10473 = (~w15876 & ~w17091) | (~w15876 & w11229) | (~w17091 & w11229);
assign w10474 = ~w560 & ~w17647;
assign w10475 = ~w1536 & ~w9509;
assign w10476 = w18786 & w3744;
assign w10477 = ~w1008 & ~w15351;
assign w10478 = w16178 & ~w13632;
assign w10479 = ~w6229 & w14436;
assign w10480 = ~w8039 & ~w16458;
assign w10481 = ~w8414 & w16341;
assign w10482 = ~w17137 & w1790;
assign w10483 = a_1 & a_39;
assign w10484 = w1736 & w962;
assign w10485 = ~w9076 & w11162;
assign w10486 = ~w8762 & ~w4664;
assign w10487 = ~w10826 & ~w9332;
assign w10488 = ~w1738 & w9052;
assign w10489 = a_40 & a_56;
assign w10490 = w10465 & w7265;
assign w10491 = ~w1012 & ~w530;
assign w10492 = ~w12820 & ~w750;
assign w10493 = ~w3787 & ~w3843;
assign w10494 = ~w16415 & w19142;
assign w10495 = a_10 & a_37;
assign w10496 = ~w3619 & ~w9455;
assign w10497 = ~w12753 & w10680;
assign w10498 = ~w1666 & ~w11680;
assign w10499 = w16603 & ~w457;
assign w10500 = ~w13247 & ~w2538;
assign w10501 = w1389 & w9964;
assign w10502 = w9474 & ~w7186;
assign w10503 = ~w17048 & ~w9643;
assign w10504 = ~w14636 & w6823;
assign w10505 = ~w2447 & w16619;
assign w10506 = a_1 & a_59;
assign w10507 = ~w10262 & ~w5446;
assign w10508 = (w19014 & w18068) | (w19014 & w15040) | (w18068 & w15040);
assign w10509 = ~w17123 & ~w8962;
assign w10510 = w15621 & ~w17669;
assign w10511 = w10262 & ~w13651;
assign w10512 = ~w3566 & ~w14494;
assign w10513 = ~w10116 & ~w5332;
assign w10514 = w17773 & ~w16979;
assign w10515 = w9115 & ~w1896;
assign w10516 = (~w13335 & ~w8917) | (~w13335 & w1384) | (~w8917 & w1384);
assign w10517 = ~w6986 & ~w12388;
assign w10518 = (~w11244 & w2769) | (~w11244 & w14887) | (w2769 & w14887);
assign w10519 = ~w6730 & ~w4393;
assign w10520 = a_38 & a_59;
assign w10521 = ~w7535 & ~w1714;
assign w10522 = a_12 & a_19;
assign w10523 = ~w10062 & w11913;
assign w10524 = w14356 & ~w11292;
assign w10525 = ~w1217 & w10326;
assign w10526 = ~w5642 & ~w3671;
assign w10527 = a_57 & a_58;
assign w10528 = ~w14189 & ~w2681;
assign w10529 = ~w2330 & ~w4607;
assign w10530 = ~w562 & w17562;
assign w10531 = ~w8829 & ~w12966;
assign w10532 = w7199 & ~w2279;
assign w10533 = ~w12561 & w3525;
assign w10534 = (~w4038 & ~w12789) | (~w4038 & w12813) | (~w12789 & w12813);
assign w10535 = ~w16562 & w5509;
assign w10536 = w5116 & w3587;
assign w10537 = w12385 & w6636;
assign w10538 = ~w6950 & ~w12336;
assign w10539 = w412 & ~w12801;
assign w10540 = (w17208 & w4329) | (w17208 & w1148) | (w4329 & w1148);
assign w10541 = ~w16079 & ~w18531;
assign w10542 = a_30 & a_63;
assign w10543 = ~w17469 & ~w10209;
assign w10544 = ~w11906 & ~w16322;
assign w10545 = a_19 & a_61;
assign w10546 = w11674 & ~w4295;
assign w10547 = ~w13858 & ~w2279;
assign w10548 = w15205 & ~w7250;
assign w10549 = ~w17481 & ~w16391;
assign w10550 = ~w8535 & ~w14981;
assign w10551 = ~w12974 & ~w1069;
assign w10552 = ~w8781 & w7953;
assign w10553 = ~w18640 & w10459;
assign w10554 = w1568 & ~w12941;
assign w10555 = w14872 & w9848;
assign w10556 = ~w17424 & ~w15013;
assign w10557 = a_35 & a_50;
assign w10558 = ~w11000 & ~w10891;
assign w10559 = ~w6373 & ~w5145;
assign w10560 = a_31 & a_41;
assign w10561 = w13713 & w17264;
assign w10562 = ~w10615 & ~w8530;
assign w10563 = ~w13317 & ~w14019;
assign w10564 = ~w5742 & ~w1907;
assign w10565 = w7553 & w8782;
assign w10566 = ~w2873 & ~w7226;
assign w10567 = w685 & w1668;
assign w10568 = a_5 & a_39;
assign w10569 = ~w13328 & w12024;
assign w10570 = ~w8175 & w18670;
assign w10571 = (w11243 & w10330) | (w11243 & w13950) | (w10330 & w13950);
assign w10572 = ~w16604 & w1517;
assign w10573 = ~w11516 & w739;
assign w10574 = w5944 & ~w15321;
assign w10575 = ~w413 & w1363;
assign w10576 = ~w17143 & ~w18754;
assign w10577 = ~w613 & ~w15905;
assign w10578 = ~w14758 & w5492;
assign w10579 = ~w5401 & ~w7854;
assign w10580 = (~w17410 & ~w12317) | (~w17410 & w4134) | (~w12317 & w4134);
assign w10581 = a_37 & a_56;
assign w10582 = ~w13052 & ~w3932;
assign w10583 = ~w13927 & ~w3106;
assign w10584 = ~w12238 & ~w16786;
assign w10585 = ~w4484 & ~w5698;
assign w10586 = ~a_42 & w10980;
assign w10587 = ~w10286 & ~w10849;
assign w10588 = ~w18610 & ~w4865;
assign w10589 = ~w6713 & ~w6999;
assign w10590 = a_16 & a_38;
assign w10591 = ~w5139 & ~w8314;
assign w10592 = ~w13840 & ~w6717;
assign w10593 = w2976 & ~w9833;
assign w10594 = w8878 & ~w17866;
assign w10595 = ~w15677 & ~w10149;
assign w10596 = ~w16141 & ~w12796;
assign w10597 = w14194 & ~w8935;
assign w10598 = w10282 & w15684;
assign w10599 = ~w12350 & ~w18224;
assign w10600 = ~w2973 & w4774;
assign w10601 = ~w10541 & w5863;
assign w10602 = ~w3300 & ~w16528;
assign w10603 = w14976 & w19198;
assign w10604 = w10940 & w16801;
assign w10605 = ~w4776 & w19171;
assign w10606 = ~w17622 & ~w1511;
assign w10607 = w11268 & w13943;
assign w10608 = ~w1762 & ~w298;
assign w10609 = w4344 & w12901;
assign w10610 = w15935 & ~w17102;
assign w10611 = ~w7793 & ~w10691;
assign w10612 = (w8509 & ~w13226) | (w8509 & w8744) | (~w13226 & w8744);
assign w10613 = (~w2769 & w15503) | (~w2769 & w17377) | (w15503 & w17377);
assign w10614 = (~w4840 & ~w13370) | (~w4840 & w18158) | (~w13370 & w18158);
assign w10615 = ~w8530 & ~w14688;
assign w10616 = ~w4962 & ~w18449;
assign w10617 = ~w13369 & ~w13842;
assign w10618 = w7872 & w2099;
assign w10619 = ~w2970 & w13226;
assign w10620 = ~w19077 & ~w16957;
assign w10621 = ~w7143 & w18766;
assign w10622 = w18180 & ~w16175;
assign w10623 = ~w2165 & ~w1680;
assign w10624 = ~w16096 & ~w2178;
assign w10625 = ~w13172 & ~w6824;
assign w10626 = a_12 & a_31;
assign w10627 = a_48 & a_49;
assign w10628 = w2564 & w17725;
assign w10629 = a_27 & a_40;
assign w10630 = w12758 & w190;
assign w10631 = ~w8463 & ~w12944;
assign w10632 = ~w11669 & ~w9126;
assign w10633 = ~a_60 & w13955;
assign w10634 = ~w4496 & ~w12566;
assign w10635 = a_36 & a_40;
assign w10636 = (w16611 & ~w7230) | (w16611 & w6748) | (~w7230 & w6748);
assign w10637 = w18394 & ~w2165;
assign w10638 = ~w696 & ~w6546;
assign w10639 = a_5 & a_16;
assign w10640 = a_5 & a_27;
assign w10641 = ~w6496 & ~w15741;
assign w10642 = ~w18341 & ~w12184;
assign w10643 = ~w18543 & w656;
assign w10644 = ~w1090 & ~w18758;
assign w10645 = ~w5012 & ~w10091;
assign w10646 = ~w2547 & ~w16790;
assign w10647 = a_5 & a_14;
assign w10648 = ~w6859 & ~w11169;
assign w10649 = ~w18350 & w13723;
assign w10650 = ~w7418 & ~w15933;
assign w10651 = a_37 & a_57;
assign w10652 = ~w15985 & ~w8204;
assign w10653 = w9873 & ~w3428;
assign w10654 = w13979 & w16272;
assign w10655 = ~w3042 & w1065;
assign w10656 = w5046 & w6860;
assign w10657 = a_11 & a_34;
assign w10658 = ~w4992 & w14527;
assign w10659 = ~w15754 & ~w3871;
assign w10660 = (~w18243 & ~w8410) | (~w18243 & w17896) | (~w8410 & w17896);
assign w10661 = w10611 & ~w17592;
assign w10662 = ~w8821 & ~w9578;
assign w10663 = a_3 & a_30;
assign w10664 = ~w5960 & ~w405;
assign w10665 = ~w13169 & ~w2443;
assign w10666 = a_22 & a_28;
assign w10667 = w2725 & ~w43;
assign w10668 = ~w18654 & w18279;
assign w10669 = ~w17933 & ~w9722;
assign w10670 = w13011 & w8631;
assign w10671 = w16900 & w2023;
assign w10672 = w600 & w11425;
assign w10673 = ~w12097 & ~w12599;
assign w10674 = a_2 & a_55;
assign w10675 = ~w18611 & ~w18326;
assign w10676 = w18094 & w3804;
assign w10677 = w17908 & ~w15086;
assign w10678 = ~w13753 & w17014;
assign w10679 = ~w19043 & ~w8728;
assign w10680 = ~w12005 & ~w3618;
assign w10681 = ~w2702 & ~w3146;
assign w10682 = (~w63 & w3609) | (~w63 & w6639) | (w3609 & w6639);
assign w10683 = ~w1927 & ~w7646;
assign w10684 = ~w14413 & ~w14752;
assign w10685 = ~w11515 & ~w11406;
assign w10686 = ~w4994 & ~w8910;
assign w10687 = ~w7025 & ~w16933;
assign w10688 = ~w3518 & ~w6028;
assign w10689 = ~w7404 & w3761;
assign w10690 = ~w9527 & ~w16169;
assign w10691 = w16248 & ~w17696;
assign w10692 = ~w9604 & w7162;
assign w10693 = ~w1861 & w13687;
assign w10694 = w8174 & w7429;
assign w10695 = ~w9860 & ~w13149;
assign w10696 = w9657 & w8190;
assign w10697 = ~w5775 & w17922;
assign w10698 = ~w2292 & ~w5966;
assign w10699 = a_58 & a_61;
assign w10700 = ~w12908 & ~w14515;
assign w10701 = a_15 & a_39;
assign w10702 = w5932 & ~w2525;
assign w10703 = ~w633 & w236;
assign w10704 = ~w2097 & ~w1106;
assign w10705 = ~w18584 & ~w2394;
assign w10706 = (~w16353 & w8448) | (~w16353 & w18193) | (w8448 & w18193);
assign w10707 = w16850 & ~w4261;
assign w10708 = w17777 & w7542;
assign w10709 = w15458 & w12058;
assign w10710 = ~w8626 & ~w3615;
assign w10711 = w18112 & ~w10295;
assign w10712 = w14585 & w16655;
assign w10713 = w9607 & w4520;
assign w10714 = ~w16206 & w11089;
assign w10715 = ~w15215 & ~w1381;
assign w10716 = a_43 & a_44;
assign w10717 = w7774 & w16965;
assign w10718 = ~w8654 & ~w2898;
assign w10719 = a_19 & a_40;
assign w10720 = ~w3151 & ~w6979;
assign w10721 = ~w6361 & ~w5708;
assign w10722 = w8453 & ~w11507;
assign w10723 = ~w442 & ~w15523;
assign w10724 = ~w3835 & ~w1006;
assign w10725 = ~w15785 & w8832;
assign w10726 = ~w2220 & ~w18404;
assign w10727 = (a_45 & w1678) | (a_45 & w8173) | (w1678 & w8173);
assign w10728 = w15578 & ~w8636;
assign w10729 = w4502 & ~w4990;
assign w10730 = ~w12018 & ~w6401;
assign w10731 = ~w18433 & w6715;
assign w10732 = ~w715 & ~w12026;
assign w10733 = a_20 & a_48;
assign w10734 = ~w2095 & ~w14708;
assign w10735 = ~w10433 & ~w2187;
assign w10736 = ~w7049 & w17816;
assign w10737 = ~w978 & w7701;
assign w10738 = w9501 & w7762;
assign w10739 = w19016 & ~w2081;
assign w10740 = ~w2354 & w11507;
assign w10741 = ~w13016 & w5222;
assign w10742 = a_33 & a_54;
assign w10743 = ~w12617 & ~w4926;
assign w10744 = ~w9885 & ~w10374;
assign w10745 = ~w14212 & ~w7855;
assign w10746 = ~w8343 & w242;
assign w10747 = (~w14304 & ~w10442) | (~w14304 & w1686) | (~w10442 & w1686);
assign w10748 = ~w2177 & ~w8458;
assign w10749 = ~w15248 & ~w8290;
assign w10750 = ~w91 & ~w8523;
assign w10751 = ~w9704 & ~w3127;
assign w10752 = ~w694 & w3368;
assign w10753 = w1114 & w18876;
assign w10754 = ~w13647 & w5191;
assign w10755 = w16611 & ~w1816;
assign w10756 = ~w7484 & ~w13936;
assign w10757 = ~w18091 & ~w17170;
assign w10758 = ~w12256 & ~w3506;
assign w10759 = w10277 & w13857;
assign w10760 = w6329 & ~w4237;
assign w10761 = (w8481 & w2769) | (w8481 & w5454) | (w2769 & w5454);
assign w10762 = ~w5346 & ~w14388;
assign w10763 = ~w1752 & ~w1210;
assign w10764 = ~w17392 & ~w6094;
assign w10765 = ~w13502 & ~w14950;
assign w10766 = ~w5090 & ~w16749;
assign w10767 = w13788 & w11195;
assign w10768 = ~w11286 & w2483;
assign w10769 = ~w10091 & ~w18697;
assign w10770 = ~w13113 & ~w8993;
assign w10771 = ~w5818 & ~w14767;
assign w10772 = w8212 & w9755;
assign w10773 = (~w10021 & ~w15903) | (~w10021 & w13530) | (~w15903 & w13530);
assign w10774 = (~w3189 & w9871) | (~w3189 & w15776) | (w9871 & w15776);
assign w10775 = ~w15344 & ~w18166;
assign w10776 = ~w16161 & ~w11076;
assign w10777 = ~w461 & w13395;
assign w10778 = ~w2421 & ~w7521;
assign w10779 = ~w15335 & w11054;
assign w10780 = w14093 & ~w16418;
assign w10781 = (~w16350 & ~w16961) | (~w16350 & w7904) | (~w16961 & w7904);
assign w10782 = ~w10602 & w13029;
assign w10783 = a_14 & a_58;
assign w10784 = ~w1657 & ~w3754;
assign w10785 = (~w15080 & w10266) | (~w15080 & w3627) | (w10266 & w3627);
assign w10786 = ~w11832 & ~w13440;
assign w10787 = ~a_27 & ~w13816;
assign w10788 = w10099 & w11634;
assign w10789 = a_18 & a_32;
assign w10790 = ~w5809 & ~w17518;
assign w10791 = w8677 & w13654;
assign w10792 = (~w11887 & ~w4074) | (~w11887 & w11369) | (~w4074 & w11369);
assign w10793 = a_18 & a_24;
assign w10794 = ~w1355 & ~w8446;
assign w10795 = ~w11958 & w18353;
assign w10796 = ~w11827 & ~w11100;
assign w10797 = ~w13169 & w9275;
assign w10798 = w11271 & ~w8590;
assign w10799 = ~w14778 & ~w3840;
assign w10800 = ~w16704 & ~w8279;
assign w10801 = a_9 & a_58;
assign w10802 = ~w17957 & ~w7883;
assign w10803 = ~w5961 & w15952;
assign w10804 = a_0 & a_14;
assign w10805 = ~w14381 & w9209;
assign w10806 = ~w11959 & ~w204;
assign w10807 = ~w1319 & w1014;
assign w10808 = ~w3245 & ~w7974;
assign w10809 = w7443 & w11354;
assign w10810 = ~w12912 & ~w9669;
assign w10811 = ~w13788 & ~w11195;
assign w10812 = ~w4968 & ~w3307;
assign w10813 = ~w1352 & ~w8270;
assign w10814 = ~w1186 & w8014;
assign w10815 = ~w6492 & ~w5925;
assign w10816 = ~w9477 & ~w17790;
assign w10817 = a_25 & a_42;
assign w10818 = ~a_14 & ~w14403;
assign w10819 = w9626 & ~w12859;
assign w10820 = (w6834 & w963) | (w6834 & w3414) | (w963 & w3414);
assign w10821 = ~w9970 & ~w16441;
assign w10822 = ~w6992 & w3015;
assign w10823 = a_6 & a_10;
assign w10824 = ~w3513 & ~w8104;
assign w10825 = (w1962 & w5500) | (w1962 & w9102) | (w5500 & w9102);
assign w10826 = ~w15547 & w4291;
assign w10827 = ~w1958 & w12532;
assign w10828 = w13082 & ~w13481;
assign w10829 = ~w3862 & w12985;
assign w10830 = ~w2774 & ~w12094;
assign w10831 = ~w4257 & ~w14560;
assign w10832 = ~w2762 & w10563;
assign w10833 = ~w5937 & ~w7605;
assign w10834 = w8419 & ~w4345;
assign w10835 = a_13 & a_18;
assign w10836 = w13483 & ~w14709;
assign w10837 = w12691 & ~w7749;
assign w10838 = ~w33 & ~w13647;
assign w10839 = w9260 & ~w17632;
assign w10840 = w13558 | w2352;
assign w10841 = ~w109 & ~w12438;
assign w10842 = ~w6505 & ~w649;
assign w10843 = w16693 & ~w11281;
assign w10844 = a_33 & a_38;
assign w10845 = ~w11680 & ~w8750;
assign w10846 = w11870 & ~w15442;
assign w10847 = ~w12260 & ~w17293;
assign w10848 = w4703 & ~w273;
assign w10849 = ~w9353 & w4486;
assign w10850 = w9064 & ~w4509;
assign w10851 = a_41 & a_62;
assign w10852 = a_15 & a_57;
assign w10853 = ~w6640 & ~w13722;
assign w10854 = (~w12859 & ~w2442) | (~w12859 & w10819) | (~w2442 & w10819);
assign w10855 = a_39 & a_50;
assign w10856 = ~w13559 & ~w4910;
assign w10857 = a_25 & a_36;
assign w10858 = ~w67 & w16102;
assign w10859 = ~w5249 & ~w12069;
assign w10860 = w6948 & ~w2396;
assign w10861 = a_14 & a_60;
assign w10862 = ~w10488 & ~w14446;
assign w10863 = ~a_2 & ~w14127;
assign w10864 = ~w3687 & ~w11152;
assign w10865 = a_23 & a_40;
assign w10866 = ~w6333 & ~w14964;
assign w10867 = a_3 & a_61;
assign w10868 = ~w8050 & ~w8693;
assign w10869 = ~w12904 & ~w13082;
assign w10870 = ~w4133 & w145;
assign w10871 = w8116 & ~w4938;
assign w10872 = w7871 & ~w16117;
assign w10873 = (~w6939 & ~w16520) | (~w6939 & w4565) | (~w16520 & w4565);
assign w10874 = ~w17714 & ~w4767;
assign w10875 = ~w4255 & ~w9947;
assign w10876 = ~w5528 & ~w18709;
assign w10877 = ~w5576 & ~w18379;
assign w10878 = ~w8858 & ~w8199;
assign w10879 = w7614 & w12220;
assign w10880 = (w10104 & w11368) | (w10104 & w17925) | (w11368 & w17925);
assign w10881 = w12170 & ~w4172;
assign w10882 = w6841 & w14898;
assign w10883 = (w11487 & w18846) | (w11487 & w3038) | (w18846 & w3038);
assign w10884 = ~w12491 & ~w2100;
assign w10885 = a_2 & a_13;
assign w10886 = ~w4841 & ~w16168;
assign w10887 = w12122 & ~w9412;
assign w10888 = ~w9532 & ~w13767;
assign w10889 = ~w5721 & ~w644;
assign w10890 = ~w10345 & w10644;
assign w10891 = w6681 & ~w100;
assign w10892 = (~w17352 & w7445) | (~w17352 & w14801) | (w7445 & w14801);
assign w10893 = ~w18133 & ~w12621;
assign w10894 = ~w10077 & ~w11716;
assign w10895 = ~w4424 & ~w1426;
assign w10896 = ~w1805 & ~w1067;
assign w10897 = ~w15984 & ~w18748;
assign w10898 = ~w3756 & ~w3090;
assign w10899 = a_0 & a_47;
assign w10900 = w16471 & ~w14730;
assign w10901 = w6932 & w6304;
assign w10902 = ~w9292 & w16395;
assign w10903 = ~w2430 & ~w1769;
assign w10904 = ~w9533 & ~w8157;
assign w10905 = w10447 & w19172;
assign w10906 = w12080 & ~w3129;
assign w10907 = ~w12955 & ~w18008;
assign w10908 = ~w5919 & ~w8775;
assign w10909 = a_34 & a_42;
assign w10910 = ~w12124 & w12357;
assign w10911 = w11255 & w16982;
assign w10912 = ~w13750 & ~w17534;
assign w10913 = w3731 & ~w4712;
assign w10914 = ~w8947 & w6865;
assign w10915 = a_9 & a_21;
assign w10916 = ~w13050 & ~w167;
assign w10917 = w7517 & w10965;
assign w10918 = w17890 & w11965;
assign w10919 = w6839 & ~w16754;
assign w10920 = a_51 & a_56;
assign w10921 = w4862 & ~w16387;
assign w10922 = ~w14853 & ~w18242;
assign w10923 = w13082 & ~w12288;
assign w10924 = ~w1613 & ~w12397;
assign w10925 = w3699 & w16095;
assign w10926 = ~w10964 & ~w2912;
assign w10927 = ~w18028 & ~w10904;
assign w10928 = ~w6376 & w686;
assign w10929 = ~w6280 & ~w18920;
assign w10930 = a_38 & a_56;
assign w10931 = ~w3109 & ~w16444;
assign w10932 = a_9 & a_51;
assign w10933 = a_47 & a_53;
assign w10934 = ~w15946 & ~w9042;
assign w10935 = ~w11886 & ~w10821;
assign w10936 = w1449 & ~w18374;
assign w10937 = ~w6590 & ~w13156;
assign w10938 = ~w7939 & ~w14366;
assign w10939 = ~w6172 & ~w8218;
assign w10940 = ~w9470 & ~w9021;
assign w10941 = ~w5067 & w13012;
assign w10942 = ~w11426 & ~w14124;
assign w10943 = w3201 & w1447;
assign w10944 = ~w5487 & ~w13133;
assign w10945 = ~w4952 & ~w14967;
assign w10946 = ~w6832 & ~w1413;
assign w10947 = ~w10071 & ~w699;
assign w10948 = w19027 & w12637;
assign w10949 = ~w2457 & ~w14811;
assign w10950 = ~w18416 & ~w17009;
assign w10951 = w11390 & ~w6085;
assign w10952 = ~w10452 & ~w19088;
assign w10953 = ~w1228 & ~w7715;
assign w10954 = ~w7757 & ~w5027;
assign w10955 = w6860 & w15209;
assign w10956 = w5890 & ~w10996;
assign w10957 = w8702 & ~w12293;
assign w10958 = ~a_43 & a_44;
assign w10959 = ~w9372 & w6917;
assign w10960 = ~w18399 & ~w4759;
assign w10961 = (w18216 & w1566) | (w18216 & w1928) | (w1566 & w1928);
assign w10962 = ~w18366 & ~w1670;
assign w10963 = ~w5193 & w6885;
assign w10964 = ~w5066 & ~w15494;
assign w10965 = ~w8168 & ~w8107;
assign w10966 = ~w19063 & ~w629;
assign w10967 = w9937 & ~w13203;
assign w10968 = (~w4865 & ~w15160) | (~w4865 & w10588) | (~w15160 & w10588);
assign w10969 = a_27 & a_36;
assign w10970 = (~w10459 & ~w15016) | (~w10459 & w7166) | (~w15016 & w7166);
assign w10971 = w9901 & w2406;
assign w10972 = ~w11210 & ~w18355;
assign w10973 = w7593 & w4483;
assign w10974 = ~w10048 & ~w1766;
assign w10975 = w18495 & ~w8099;
assign w10976 = w7246 & ~w2657;
assign w10977 = w13858 & w15788;
assign w10978 = ~w4124 & w9798;
assign w10979 = w1502 & ~w6351;
assign w10980 = w3089 & w8589;
assign w10981 = ~w16064 & ~w17672;
assign w10982 = ~w1846 & ~w13113;
assign w10983 = a_23 & a_59;
assign w10984 = a_57 & a_62;
assign w10985 = ~w16296 & ~w14482;
assign w10986 = a_14 & a_36;
assign w10987 = w10804 & ~w17003;
assign w10988 = ~w14737 & ~w5668;
assign w10989 = ~w1068 & ~w17575;
assign w10990 = w690 & w10855;
assign w10991 = (~w13283 & ~w5300) | (~w13283 & w4149) | (~w5300 & w4149);
assign w10992 = ~w5828 & ~w312;
assign w10993 = ~w12415 & ~w1406;
assign w10994 = w4216 & ~w10066;
assign w10995 = a_56 & a_59;
assign w10996 = ~w2702 & ~w18507;
assign w10997 = ~w4877 & w343;
assign w10998 = ~w13949 & ~w15451;
assign w10999 = (w6134 & w5438) | (w6134 & w7792) | (w5438 & w7792);
assign w11000 = ~w6681 & w100;
assign w11001 = w1974 & ~w3967;
assign w11002 = w6426 & w19046;
assign w11003 = a_41 & a_55;
assign w11004 = ~w7659 & w70;
assign w11005 = ~w14786 & w8999;
assign w11006 = (w7768 & w18797) | (w7768 & w14232) | (w18797 & w14232);
assign w11007 = ~w2380 & ~w16218;
assign w11008 = ~w3872 & ~w14385;
assign w11009 = ~w10914 & ~w1987;
assign w11010 = ~w17682 & w5566;
assign w11011 = ~w12921 & ~w6011;
assign w11012 = ~w18277 & w6344;
assign w11013 = ~w15162 & w4743;
assign w11014 = (~w6848 & ~w11707) | (~w6848 & w16173) | (~w11707 & w16173);
assign w11015 = ~w13545 & ~w610;
assign w11016 = ~w1022 & ~w1776;
assign w11017 = ~w9291 & ~w5575;
assign w11018 = ~w18397 & ~w17007;
assign w11019 = ~w7257 & ~w2503;
assign w11020 = ~w12249 & ~w14663;
assign w11021 = (~w3523 & ~w17674) | (~w3523 & w15561) | (~w17674 & w15561);
assign w11022 = ~w14922 & w4717;
assign w11023 = ~w2054 & ~w5004;
assign w11024 = ~w2973 & ~w2257;
assign w11025 = w6277 & ~w5354;
assign w11026 = ~w18872 & ~w9610;
assign w11027 = w9281 & ~w4070;
assign w11028 = ~w17034 & ~w12106;
assign w11029 = (~w13206 & ~w5926) | (~w13206 & w14346) | (~w5926 & w14346);
assign w11030 = w6543 & ~w18693;
assign w11031 = ~w1568 & w12941;
assign w11032 = ~w10647 & ~w7880;
assign w11033 = a_10 & a_27;
assign w11034 = w15794 & ~w7656;
assign w11035 = w13533 & ~w2277;
assign w11036 = ~w12495 & w7617;
assign w11037 = ~w14583 & ~w8316;
assign w11038 = w6829 & w1468;
assign w11039 = a_8 & a_9;
assign w11040 = a_40 & a_48;
assign w11041 = ~w16884 & ~w10567;
assign w11042 = ~w14696 & w7656;
assign w11043 = ~w6647 & ~w15434;
assign w11044 = a_18 & a_48;
assign w11045 = ~w9090 & ~w8310;
assign w11046 = ~w10557 & ~w2527;
assign w11047 = w18443 & ~w18143;
assign w11048 = ~w18488 & w8918;
assign w11049 = ~w13151 & w9309;
assign w11050 = (~w963 & w1482) | (~w963 & ~w16291) | (w1482 & ~w16291);
assign w11051 = w12433 & w268;
assign w11052 = ~w14722 & ~w384;
assign w11053 = ~w18909 & ~w17456;
assign w11054 = ~w12793 & ~w10725;
assign w11055 = w18831 & ~w7063;
assign w11056 = ~w11519 & ~w16090;
assign w11057 = ~w1422 & ~w7046;
assign w11058 = w9979 & ~w12483;
assign w11059 = ~w14728 & ~w16974;
assign w11060 = ~w3273 & w9552;
assign w11061 = ~w14736 & ~w9719;
assign w11062 = (~w14073 & ~w6530) | (~w14073 & w8245) | (~w6530 & w8245);
assign w11063 = w11943 & ~w41;
assign w11064 = ~w12042 & ~w7568;
assign w11065 = ~w12481 & ~w5036;
assign w11066 = w7059 & w6629;
assign w11067 = ~w18423 & ~w14070;
assign w11068 = (~w16917 & w16062) | (~w16917 & w18171) | (w16062 & w18171);
assign w11069 = ~w57 & ~w17807;
assign w11070 = (~w229 & ~w14204) | (~w229 & w12816) | (~w14204 & w12816);
assign w11071 = ~w2068 & w17556;
assign w11072 = w12983 & ~w14109;
assign w11073 = w11021 & ~w6072;
assign w11074 = ~w13833 & w14325;
assign w11075 = ~w862 & ~w3392;
assign w11076 = ~w17699 & ~w10304;
assign w11077 = ~w3099 & w11163;
assign w11078 = ~w11430 & ~w13457;
assign w11079 = a_19 & a_28;
assign w11080 = a_48 & a_60;
assign w11081 = a_7 & a_26;
assign w11082 = ~w9236 & ~w15479;
assign w11083 = w14511 & w8092;
assign w11084 = ~w9457 & ~w6739;
assign w11085 = ~w8632 & w13031;
assign w11086 = ~w12547 & ~w5006;
assign w11087 = ~w5893 & w8855;
assign w11088 = w14330 & w13909;
assign w11089 = ~w6115 & ~w807;
assign w11090 = w9889 & ~w8137;
assign w11091 = ~w5146 & ~w12320;
assign w11092 = ~w10396 & ~w6118;
assign w11093 = ~w11265 & ~w12341;
assign w11094 = a_2 & a_10;
assign w11095 = ~w1515 & w571;
assign w11096 = ~w14843 & ~w10477;
assign w11097 = w55 & ~w17342;
assign w11098 = ~w18464 & ~w2993;
assign w11099 = w4711 & ~w2209;
assign w11100 = w2793 & ~w4032;
assign w11101 = ~w15261 & w16629;
assign w11102 = w9422 & w15841;
assign w11103 = ~w17795 & ~w8087;
assign w11104 = ~w17387 & ~w2235;
assign w11105 = a_18 & a_19;
assign w11106 = a_12 & a_45;
assign w11107 = ~w8871 & ~w13043;
assign w11108 = w11893 & w2323;
assign w11109 = ~w13630 & ~w12550;
assign w11110 = a_28 & a_58;
assign w11111 = w12134 & w8111;
assign w11112 = ~w5436 & ~w1526;
assign w11113 = ~w7355 & w17867;
assign w11114 = ~w6208 & w6593;
assign w11115 = w2771 & w6044;
assign w11116 = ~w12752 & ~w16307;
assign w11117 = ~w6150 & ~w3349;
assign w11118 = ~w2639 & ~w18064;
assign w11119 = ~w9642 & ~w13799;
assign w11120 = ~w15003 & ~w13120;
assign w11121 = ~w7607 & ~w7024;
assign w11122 = ~w6382 & ~w956;
assign w11123 = ~w18583 & ~w17273;
assign w11124 = ~w12667 & w15987;
assign w11125 = w1186 & ~w8014;
assign w11126 = ~w13449 & ~w17440;
assign w11127 = ~w15223 & ~w9089;
assign w11128 = ~w7863 & ~w17004;
assign w11129 = w10187 & w9049;
assign w11130 = ~w12803 & ~w8659;
assign w11131 = ~w8468 & ~w8982;
assign w11132 = ~w15052 & ~w5621;
assign w11133 = ~w15300 & ~w2558;
assign w11134 = a_32 & a_49;
assign w11135 = ~w13607 & ~w3440;
assign w11136 = ~w3568 & ~w4860;
assign w11137 = a_0 & a_20;
assign w11138 = (~w14573 & ~w4558) | (~w14573 & w6103) | (~w4558 & w6103);
assign w11139 = ~w13889 & ~w10360;
assign w11140 = ~w12732 & ~w12014;
assign w11141 = (~w4648 & ~w5182) | (~w4648 & w2872) | (~w5182 & w2872);
assign w11142 = ~w11081 & w17820;
assign w11143 = ~w12182 & ~w12107;
assign w11144 = ~w5890 & ~w11918;
assign w11145 = ~w1284 & w13441;
assign w11146 = w7594 & w14296;
assign w11147 = ~w3097 & ~w13010;
assign w11148 = ~w7968 & ~w2546;
assign w11149 = ~w4911 & ~w12936;
assign w11150 = ~w16654 & ~w7669;
assign w11151 = ~w11266 & ~w18365;
assign w11152 = ~w11317 & ~w8572;
assign w11153 = (~w16328 & w11029) | (~w16328 & w17799) | (w11029 & w17799);
assign w11154 = a_17 & a_26;
assign w11155 = (~w17775 & ~w8668) | (~w17775 & w12196) | (~w8668 & w12196);
assign w11156 = ~w17429 & ~w12438;
assign w11157 = ~w6009 & ~w9183;
assign w11158 = ~w7018 & ~w2705;
assign w11159 = w16419 & ~w8203;
assign w11160 = ~w14435 & w13195;
assign w11161 = ~w4006 & ~w1624;
assign w11162 = ~w10025 & ~w8801;
assign w11163 = ~w7588 & ~w774;
assign w11164 = a_20 & a_30;
assign w11165 = a_41 & a_44;
assign w11166 = ~w15968 & ~w16492;
assign w11167 = ~w15655 & ~w14266;
assign w11168 = ~w17700 & ~w11035;
assign w11169 = ~w183 & ~w18999;
assign w11170 = ~w1160 & ~w11967;
assign w11171 = ~w6680 & w19142;
assign w11172 = ~w8655 & w17542;
assign w11173 = (~w15163 & w10330) | (~w15163 & w224) | (w10330 & w224);
assign w11174 = (w9221 & w11397) | (w9221 & w7291) | (w11397 & w7291);
assign w11175 = ~w1754 & ~w10409;
assign w11176 = ~w3517 & ~w14334;
assign w11177 = a_6 & a_44;
assign w11178 = ~w17633 & ~w641;
assign w11179 = (w4355 & w16015) | (w4355 & w4780) | (w16015 & w4780);
assign w11180 = ~w11224 & ~w17237;
assign w11181 = w8050 & w8693;
assign w11182 = ~w5857 & ~w17210;
assign w11183 = w233 & ~w9888;
assign w11184 = w9248 & w78;
assign w11185 = ~w11396 & ~w6831;
assign w11186 = ~w15367 & ~w11952;
assign w11187 = ~w10330 & w2902;
assign w11188 = w15443 & w4997;
assign w11189 = a_6 & a_19;
assign w11190 = ~w9741 & ~w2790;
assign w11191 = a_40 & a_41;
assign w11192 = (~w4720 & ~w2260) | (~w4720 & w3539) | (~w2260 & w3539);
assign w11193 = ~w5152 & ~w4363;
assign w11194 = (~w1971 & ~w6397) | (~w1971 & w4887) | (~w6397 & w4887);
assign w11195 = ~w12127 & ~w12540;
assign w11196 = a_13 & a_31;
assign w11197 = w13404 & w6223;
assign w11198 = w1035 & w17172;
assign w11199 = w13269 & w9837;
assign w11200 = w4159 & w14251;
assign w11201 = ~w6048 & ~w16543;
assign w11202 = ~a_36 & w11200;
assign w11203 = a_11 & a_62;
assign w11204 = (~w2663 & w963) | (~w2663 & w18402) | (w963 & w18402);
assign w11205 = ~w5172 & ~w2365;
assign w11206 = ~w14328 & ~w573;
assign w11207 = ~w15726 & w16708;
assign w11208 = a_0 & a_10;
assign w11209 = ~w15076 & ~w12868;
assign w11210 = ~w9170 & ~w4705;
assign w11211 = a_4 & a_9;
assign w11212 = ~w284 & ~w16792;
assign w11213 = ~w6682 & ~w2734;
assign w11214 = w15824 & ~w8986;
assign w11215 = (~w16884 & ~w11041) | (~w16884 & w6343) | (~w11041 & w6343);
assign w11216 = ~w5194 & ~w5433;
assign w11217 = ~w8997 & ~w12636;
assign w11218 = ~w11095 & ~w4601;
assign w11219 = w9446 & w3237;
assign w11220 = ~w7838 & ~w16514;
assign w11221 = w15573 & w10087;
assign w11222 = w11987 & w5842;
assign w11223 = ~w4128 & ~w15506;
assign w11224 = a_36 & a_62;
assign w11225 = ~w14631 & ~w12075;
assign w11226 = a_0 & a_56;
assign w11227 = ~w4890 & ~w13819;
assign w11228 = ~w5587 & ~w14455;
assign w11229 = w621 & ~w15876;
assign w11230 = ~w3663 & ~w14073;
assign w11231 = ~w18181 & ~w1410;
assign w11232 = w12885 & w16608;
assign w11233 = ~w2968 & w6931;
assign w11234 = ~w4327 & w15890;
assign w11235 = ~w8831 & ~w1644;
assign w11236 = w6442 & w17080;
assign w11237 = ~w18828 & ~w17398;
assign w11238 = ~w6481 & w3540;
assign w11239 = ~w9937 & w13203;
assign w11240 = ~w15230 & w2309;
assign w11241 = a_0 & a_39;
assign w11242 = ~w18567 & ~w4987;
assign w11243 = (w13777 & w666) | (w13777 & w6185) | (w666 & w6185);
assign w11244 = ~w13082 & ~w10330;
assign w11245 = (~w8636 & w11391) | (~w8636 & w7470) | (w11391 & w7470);
assign w11246 = a_12 & a_29;
assign w11247 = ~w10660 & w18674;
assign w11248 = ~w55 & w17342;
assign w11249 = (~w18733 & w5675) | (~w18733 & w6307) | (w5675 & w6307);
assign w11250 = ~w3988 & w13789;
assign w11251 = w3353 & w14427;
assign w11252 = ~w3554 & ~w3634;
assign w11253 = ~w2609 & w14888;
assign w11254 = ~w15428 & ~w8413;
assign w11255 = ~w3423 & ~w7450;
assign w11256 = ~w15058 & ~w3957;
assign w11257 = ~w10626 & w7996;
assign w11258 = ~w18001 & ~w12515;
assign w11259 = ~w2623 & ~w13657;
assign w11260 = ~w3507 & ~w7027;
assign w11261 = ~w8552 & w4361;
assign w11262 = ~w8849 & ~w11824;
assign w11263 = ~w13144 & ~w9925;
assign w11264 = ~w3997 & w14676;
assign w11265 = ~w8528 & ~w9727;
assign w11266 = ~w16370 & ~w4248;
assign w11267 = ~w13864 & w5568;
assign w11268 = ~w14973 & ~w17338;
assign w11269 = ~w17524 & ~w12489;
assign w11270 = w15061 & ~w4951;
assign w11271 = a_49 & a_63;
assign w11272 = a_9 & a_48;
assign w11273 = a_21 & a_41;
assign w11274 = w1755 & w9938;
assign w11275 = ~w8409 & ~w5276;
assign w11276 = ~w2995 & ~w12071;
assign w11277 = a_31 & a_60;
assign w11278 = ~w225 & ~w14409;
assign w11279 = w15890 & ~w12730;
assign w11280 = w3658 & w612;
assign w11281 = ~w11557 & ~w15790;
assign w11282 = ~w11278 & ~w5457;
assign w11283 = w14181 & ~w5596;
assign w11284 = ~w12326 & w13551;
assign w11285 = ~w3921 & w6727;
assign w11286 = ~w2769 & w9521;
assign w11287 = ~w7012 & ~w3922;
assign w11288 = ~w10372 & ~w1463;
assign w11289 = ~w16048 & ~w5497;
assign w11290 = a_5 & a_50;
assign w11291 = ~w13397 & ~w4493;
assign w11292 = ~w7312 & ~w2703;
assign w11293 = a_17 & a_38;
assign w11294 = w13894 & ~w5073;
assign w11295 = (w3279 & w19005) | (w3279 & w4232) | (w19005 & w4232);
assign w11296 = a_35 & a_61;
assign w11297 = a_1 & a_32;
assign w11298 = w14279 & w5765;
assign w11299 = ~w15669 & w5607;
assign w11300 = ~w2984 & ~w16324;
assign w11301 = ~w10041 & ~w15699;
assign w11302 = w2225 & w1495;
assign w11303 = a_24 & a_50;
assign w11304 = ~w15930 & ~w15696;
assign w11305 = ~w15667 & ~w10714;
assign w11306 = a_14 & a_45;
assign w11307 = w1904 & ~w18639;
assign w11308 = w10108 & w15102;
assign w11309 = ~w3347 & ~w16783;
assign w11310 = ~w14617 & ~w6581;
assign w11311 = w18571 & ~w10413;
assign w11312 = ~w4607 & ~w12039;
assign w11313 = w15230 & ~w12209;
assign w11314 = ~w7205 & ~w1940;
assign w11315 = w7704 & ~w16613;
assign w11316 = a_14 & a_27;
assign w11317 = w9650 & w14128;
assign w11318 = ~w7548 & w13199;
assign w11319 = ~w9817 & ~w15840;
assign w11320 = ~w15796 & w10331;
assign w11321 = ~w8339 & w18309;
assign w11322 = (~w3953 & ~w5852) | (~w3953 & w13421) | (~w5852 & w13421);
assign w11323 = ~w1455 & ~w222;
assign w11324 = w17483 & ~w19113;
assign w11325 = w7115 & w8058;
assign w11326 = ~w13765 & ~w8880;
assign w11327 = w17402 & w9033;
assign w11328 = ~w1727 & ~w7480;
assign w11329 = a_25 & a_49;
assign w11330 = w17702 & w16454;
assign w11331 = (~w10462 & ~w5754) | (~w10462 & w17739) | (~w5754 & w17739);
assign w11332 = a_29 & a_40;
assign w11333 = a_23 & a_42;
assign w11334 = ~w12277 & ~w8313;
assign w11335 = w14684 & w4829;
assign w11336 = a_37 & a_47;
assign w11337 = ~w13356 & ~w3879;
assign w11338 = a_62 & w6252;
assign w11339 = w17898 & ~w843;
assign w11340 = a_55 & a_59;
assign w11341 = ~w7893 & ~w7960;
assign w11342 = ~w646 & ~w17523;
assign w11343 = a_15 & a_19;
assign w11344 = ~w12271 & ~w14473;
assign w11345 = w17425 & w14055;
assign w11346 = ~w10611 & w17592;
assign w11347 = w2881 & ~w11639;
assign w11348 = ~w6585 & w12270;
assign w11349 = w9825 & ~w2783;
assign w11350 = ~w8876 & ~w8331;
assign w11351 = (w7102 & w17822) | (w7102 & w9095) | (w17822 & w9095);
assign w11352 = w4037 & ~w1825;
assign w11353 = w5090 & w16749;
assign w11354 = a_13 & a_16;
assign w11355 = ~w2489 & ~w8732;
assign w11356 = ~w11890 & ~w1111;
assign w11357 = ~w14311 & ~w2376;
assign w11358 = ~w15036 & ~w15195;
assign w11359 = ~w2408 & ~w7816;
assign w11360 = ~w8574 & w5291;
assign w11361 = w1859 & w1315;
assign w11362 = ~w15705 & ~w10355;
assign w11363 = ~w12960 & w5333;
assign w11364 = ~w17195 & ~w15157;
assign w11365 = ~w427 & ~w14252;
assign w11366 = ~w12795 & w893;
assign w11367 = ~w12657 & ~w987;
assign w11368 = w6566 & ~w17991;
assign w11369 = w5602 & ~w11887;
assign w11370 = a_7 & a_55;
assign w11371 = ~w9250 & ~w5846;
assign w11372 = w2576 & w9577;
assign w11373 = w5219 & w1038;
assign w11374 = a_14 & a_50;
assign w11375 = w8137 & ~w7434;
assign w11376 = w7973 & w12847;
assign w11377 = ~w3018 & ~w3192;
assign w11378 = ~w16814 & ~w8789;
assign w11379 = ~w12380 & ~w11560;
assign w11380 = ~w15714 & ~w14025;
assign w11381 = ~w6311 & ~w864;
assign w11382 = w7899 & ~w1257;
assign w11383 = ~w10495 & ~w14925;
assign w11384 = w15515 & w7603;
assign w11385 = (~w10040 & ~w18132) | (~w10040 & w1820) | (~w18132 & w1820);
assign w11386 = ~w2254 & ~w6448;
assign w11387 = ~w5929 & w1765;
assign w11388 = ~w11909 & w9794;
assign w11389 = w7158 & w8091;
assign w11390 = ~w9128 & ~w18668;
assign w11391 = (w15578 & w17665) | (w15578 & w14835) | (w17665 & w14835);
assign w11392 = ~w6370 & ~w6587;
assign w11393 = w3717 & ~w12011;
assign w11394 = ~w18816 & ~w17324;
assign w11395 = a_21 & a_59;
assign w11396 = ~w1312 & w7654;
assign w11397 = w14488 | w6087;
assign w11398 = ~w14281 & ~w2499;
assign w11399 = ~w5831 & ~w9312;
assign w11400 = a_31 & a_46;
assign w11401 = a_40 & a_43;
assign w11402 = w11241 & w17471;
assign w11403 = ~w10313 & ~w7010;
assign w11404 = ~w8875 & ~w5586;
assign w11405 = ~w3735 & ~w18790;
assign w11406 = ~w3691 & ~w15979;
assign w11407 = w12333 & ~w9732;
assign w11408 = ~w372 & ~w17326;
assign w11409 = ~w16959 & ~w16109;
assign w11410 = ~w14949 & ~w8275;
assign w11411 = ~w2710 & w7668;
assign w11412 = ~w3878 & ~w16404;
assign w11413 = a_9 & a_59;
assign w11414 = w10269 & ~w9520;
assign w11415 = ~w9184 & w14394;
assign w11416 = ~w1946 & ~w2582;
assign w11417 = ~w5851 & ~w431;
assign w11418 = ~w8182 & w14391;
assign w11419 = ~w9685 & ~w1476;
assign w11420 = w16432 & ~w9058;
assign w11421 = ~w12785 & ~w12627;
assign w11422 = ~w2413 & w1127;
assign w11423 = ~w13351 & ~w4768;
assign w11424 = ~w582 & w4322;
assign w11425 = a_1 & a_61;
assign w11426 = w9422 & w18850;
assign w11427 = w315 & ~w5778;
assign w11428 = a_21 & a_58;
assign w11429 = ~w18714 & ~w3937;
assign w11430 = w15472 & w1898;
assign w11431 = w3775 & ~w9570;
assign w11432 = ~w10981 & ~w11808;
assign w11433 = ~w13253 & ~w19034;
assign w11434 = (~w12730 & ~w4327) | (~w12730 & w11279) | (~w4327 & w11279);
assign w11435 = w6043 & ~w14593;
assign w11436 = w4098 & w4272;
assign w11437 = ~w116 & ~w8103;
assign w11438 = ~w13734 & w15851;
assign w11439 = ~w19028 & ~w17492;
assign w11440 = ~w11250 & ~w4540;
assign w11441 = ~w16498 & w13299;
assign w11442 = ~w79 & ~w11718;
assign w11443 = w17361 & w12435;
assign w11444 = ~w16650 & w8996;
assign w11445 = w8442 & w1162;
assign w11446 = w11752 & w6176;
assign w11447 = ~w16432 & w9058;
assign w11448 = w16505 & ~w14776;
assign w11449 = ~w9321 & ~w2245;
assign w11450 = ~w13709 & ~w14195;
assign w11451 = ~w6543 & w18693;
assign w11452 = w210 & w5988;
assign w11453 = ~w17131 & ~w2819;
assign w11454 = ~w14834 & ~w10170;
assign w11455 = a_28 & a_48;
assign w11456 = w18765 & ~w13517;
assign w11457 = ~w7695 & w4074;
assign w11458 = ~w3898 & w5812;
assign w11459 = w8148 & ~w18548;
assign w11460 = w3725 & w17760;
assign w11461 = w9885 & w10374;
assign w11462 = w4133 & ~w13001;
assign w11463 = ~w16331 & ~w829;
assign w11464 = a_15 & a_24;
assign w11465 = (~w13673 & ~w9580) | (~w13673 & w9965) | (~w9580 & w9965);
assign w11466 = ~w15768 & ~w6767;
assign w11467 = ~w4211 & w13528;
assign w11468 = ~w6830 & w2991;
assign w11469 = ~w14242 & ~w6817;
assign w11470 = ~w12997 & ~w16228;
assign w11471 = ~w6080 & w4120;
assign w11472 = ~w8412 & ~w10955;
assign w11473 = w3799 & w12945;
assign w11474 = w3960 & w1407;
assign w11475 = w10519 & w7957;
assign w11476 = ~w2041 & ~w18428;
assign w11477 = ~w13581 & ~w13727;
assign w11478 = w12427 & ~w4470;
assign w11479 = ~w2253 & ~w4071;
assign w11480 = w10742 & w18688;
assign w11481 = (w13508 & w18316) | (w13508 & w14430) | (w18316 & w14430);
assign w11482 = ~w12737 & ~w10358;
assign w11483 = a_50 & a_56;
assign w11484 = ~w7457 & ~w17996;
assign w11485 = ~w14080 & ~w16641;
assign w11486 = ~w16674 & ~w596;
assign w11487 = (a_54 & w2878) | (a_54 & w14335) | (w2878 & w14335);
assign w11488 = (w14465 & w7610) | (w14465 & w9152) | (w7610 & w9152);
assign w11489 = w10138 & ~w8758;
assign w11490 = ~w9697 & ~w18266;
assign w11491 = ~w7580 & ~w11077;
assign w11492 = ~w10167 & ~w7645;
assign w11493 = ~w1473 & ~w13791;
assign w11494 = a_5 & a_7;
assign w11495 = ~w6959 & ~w2369;
assign w11496 = w16626 & ~w9399;
assign w11497 = ~w12776 & ~w12007;
assign w11498 = ~w15959 & ~w6323;
assign w11499 = w1348 & w6597;
assign w11500 = ~w17028 & ~w4049;
assign w11501 = w8595 & ~w876;
assign w11502 = ~w10912 & w18281;
assign w11503 = w11116 & w14988;
assign w11504 = a_51 & a_58;
assign w11505 = ~w11334 & ~w2742;
assign w11506 = a_23 & a_52;
assign w11507 = ~w2071 & ~w19019;
assign w11508 = ~w3585 & w18405;
assign w11509 = w6943 & ~w3829;
assign w11510 = ~w8991 & ~w5346;
assign w11511 = ~w14719 & ~w17732;
assign w11512 = ~w13106 & w3579;
assign w11513 = ~w16847 & ~w6466;
assign w11514 = w15990 & w15491;
assign w11515 = ~w17136 & ~w12033;
assign w11516 = a_26 & a_55;
assign w11517 = ~w7565 & w9982;
assign w11518 = ~w9414 & ~w1914;
assign w11519 = ~w3116 & ~w2951;
assign w11520 = w16533 & w12443;
assign w11521 = ~w8702 & w12293;
assign w11522 = ~w2302 & ~w1393;
assign w11523 = (w16917 & w2438) | (w16917 & w3709) | (w2438 & w3709);
assign w11524 = ~w11362 & ~w5119;
assign w11525 = ~w16701 & ~w2291;
assign w11526 = ~w7994 & w4695;
assign w11527 = ~w10708 & ~w18483;
assign w11528 = ~w7528 & ~w6084;
assign w11529 = ~w8232 & ~w132;
assign w11530 = ~w9701 & ~w4248;
assign w11531 = ~w5354 & ~w6562;
assign w11532 = (~w14352 & ~w12673) | (~w14352 & w15259) | (~w12673 & w15259);
assign w11533 = ~w5520 & ~w9829;
assign w11534 = ~w4694 & ~w15340;
assign w11535 = w10565 & w10464;
assign w11536 = ~w15766 & ~w5233;
assign w11537 = ~w11478 & ~w15286;
assign w11538 = w14528 & ~w15522;
assign w11539 = ~w3101 & w5648;
assign w11540 = a_57 & a_61;
assign w11541 = w13928 & w2445;
assign w11542 = w4527 & ~w13947;
assign w11543 = ~w18543 & ~w4238;
assign w11544 = w19012 & w13835;
assign w11545 = (~w18913 & ~w9513) | (~w18913 & w5992) | (~w9513 & w5992);
assign w11546 = ~w3726 & ~w1572;
assign w11547 = ~w18083 & ~w2731;
assign w11548 = (w16582 & w15737) | (w16582 & w14587) | (w15737 & w14587);
assign w11549 = ~w3203 & ~w11688;
assign w11550 = w8080 & ~w13639;
assign w11551 = a_18 & a_33;
assign w11552 = ~w15417 & ~w6725;
assign w11553 = ~w2062 & w12231;
assign w11554 = ~w16803 & ~w5383;
assign w11555 = ~w14932 & ~w3801;
assign w11556 = ~w19098 & ~w15473;
assign w11557 = w9476 & ~w17157;
assign w11558 = ~w8990 & ~w238;
assign w11559 = a_3 & a_27;
assign w11560 = (~w4318 & w5767) | (~w4318 & w10120) | (w5767 & w10120);
assign w11561 = ~w7081 & ~w5753;
assign w11562 = ~w11306 & ~w1490;
assign w11563 = ~a_16 & w2249;
assign w11564 = ~w5349 & w13185;
assign w11565 = ~w13438 & ~w8614;
assign w11566 = ~w7912 & ~w1767;
assign w11567 = ~w12703 & ~w10336;
assign w11568 = w9267 & ~w3986;
assign w11569 = ~w9901 & ~w2406;
assign w11570 = a_15 & a_52;
assign w11571 = ~w6495 & ~w4683;
assign w11572 = ~w12821 & ~w5811;
assign w11573 = ~w2573 & w6160;
assign w11574 = ~w9767 & ~w8261;
assign w11575 = w12652 & w249;
assign w11576 = ~w8636 & w1413;
assign w11577 = ~w4827 & ~w17992;
assign w11578 = w2557 & ~w14115;
assign w11579 = w1063 & ~w16460;
assign w11580 = ~w12804 & w16642;
assign w11581 = ~w17830 & ~w2877;
assign w11582 = ~w10191 & ~w6007;
assign w11583 = ~w13742 & w4640;
assign w11584 = w2772 & w3479;
assign w11585 = w16155 & ~w2508;
assign w11586 = ~w5302 & ~w16235;
assign w11587 = ~w11696 & ~w10640;
assign w11588 = ~w18906 & ~w7937;
assign w11589 = ~w16332 & ~w7928;
assign w11590 = ~w12346 & ~w11188;
assign w11591 = ~w16482 & ~w13868;
assign w11592 = ~w12363 & ~w18030;
assign w11593 = ~w6967 & ~w16579;
assign w11594 = ~w14440 & ~w13679;
assign w11595 = ~w1925 & ~w13274;
assign w11596 = w8701 & ~w5626;
assign w11597 = ~w8706 & ~w5371;
assign w11598 = w868 & ~w17907;
assign w11599 = (~w7087 & ~w7249) | (~w7087 & w13728) | (~w7249 & w13728);
assign w11600 = a_42 & a_57;
assign w11601 = a_22 & a_51;
assign w11602 = w13949 & w15451;
assign w11603 = ~w18916 & ~w17026;
assign w11604 = (w1413 & w16375) | (w1413 & w1808) | (w16375 & w1808);
assign w11605 = (w4195 & w10330) | (w4195 & w16618) | (w10330 & w16618);
assign w11606 = ~w3335 & ~w11774;
assign w11607 = w7806 & w5348;
assign w11608 = w10428 & w18953;
assign w11609 = ~w2792 & ~w17885;
assign w11610 = ~w4711 & w2209;
assign w11611 = ~w16634 & ~w17459;
assign w11612 = ~w17331 & ~w14107;
assign w11613 = ~w872 & ~w3878;
assign w11614 = w16402 & w18988;
assign w11615 = ~w14830 & ~w4319;
assign w11616 = w8010 & w14849;
assign w11617 = ~w14567 & ~w1385;
assign w11618 = w11897 & ~w3543;
assign w11619 = ~w6106 & w4613;
assign w11620 = ~w9931 & w17177;
assign w11621 = ~w4710 & ~w7938;
assign w11622 = ~w15786 & w5647;
assign w11623 = ~w13667 & ~w18547;
assign w11624 = w13477 & w16007;
assign w11625 = ~w5434 & ~w8649;
assign w11626 = w12275 & ~w17825;
assign w11627 = w5828 & w312;
assign w11628 = ~w1396 & ~w12511;
assign w11629 = ~w14401 & ~w18858;
assign w11630 = ~w7723 & ~w9357;
assign w11631 = w8232 & w132;
assign w11632 = ~w15701 & ~w15840;
assign w11633 = ~w4478 & w12825;
assign w11634 = w13979 & w13985;
assign w11635 = ~w9047 & ~w1252;
assign w11636 = (~w10330 & w15201) | (~w10330 & w6273) | (w15201 & w6273);
assign w11637 = ~w15899 & ~w11246;
assign w11638 = a_5 & a_56;
assign w11639 = ~w9336 & w17249;
assign w11640 = ~w5011 & ~w2393;
assign w11641 = w14614 & w14400;
assign w11642 = w18582 & ~w1425;
assign w11643 = ~w14598 & ~w4338;
assign w11644 = ~w2769 & w9818;
assign w11645 = ~w8871 & ~w8716;
assign w11646 = ~w13330 & w14109;
assign w11647 = ~w15492 & w9162;
assign w11648 = ~w2005 & ~w12282;
assign w11649 = w12624 & w14033;
assign w11650 = w2176 & ~w5756;
assign w11651 = ~w13897 & ~w8892;
assign w11652 = ~w11840 & ~w13279;
assign w11653 = (~w15668 & ~w13046) | (~w15668 & w12802) | (~w13046 & w12802);
assign w11654 = ~w3182 & w14238;
assign w11655 = a_14 & a_51;
assign w11656 = w6065 & ~w5441;
assign w11657 = w1283 & ~w10513;
assign w11658 = w1706 & ~w15122;
assign w11659 = ~w11748 & ~w8756;
assign w11660 = w8971 & w6928;
assign w11661 = ~w5976 & ~w2962;
assign w11662 = a_36 & a_53;
assign w11663 = ~w12150 & ~w18613;
assign w11664 = a_22 & a_62;
assign w11665 = w4619 & ~w18745;
assign w11666 = w13909 & ~w17938;
assign w11667 = w17473 & w8438;
assign w11668 = ~w14123 & ~w8216;
assign w11669 = a_31 & a_35;
assign w11670 = ~w17774 & w11054;
assign w11671 = ~w15404 & ~w13309;
assign w11672 = w12433 & ~w9182;
assign w11673 = ~w8596 & ~w13360;
assign w11674 = ~w17793 & ~w771;
assign w11675 = ~w17550 & ~w8244;
assign w11676 = w9410 & w19083;
assign w11677 = ~w15 & ~w8601;
assign w11678 = ~w2034 & ~w18705;
assign w11679 = ~w17278 & ~w13040;
assign w11680 = ~w4652 & ~w5380;
assign w11681 = (~w15834 & ~w1041) | (~w15834 & w9022) | (~w1041 & w9022);
assign w11682 = ~w12810 & ~w1334;
assign w11683 = ~w16652 & ~w3359;
assign w11684 = w14150 & ~w2370;
assign w11685 = ~w1182 & ~w11053;
assign w11686 = w6420 & ~w1262;
assign w11687 = ~w2040 & ~w10135;
assign w11688 = ~w8943 & w5068;
assign w11689 = ~w7825 & ~w13986;
assign w11690 = w17999 & ~w11595;
assign w11691 = ~w5816 & w17548;
assign w11692 = ~w18734 & ~w1848;
assign w11693 = ~w8597 & w9498;
assign w11694 = a_9 & a_35;
assign w11695 = ~w14698 & ~w11778;
assign w11696 = a_4 & a_28;
assign w11697 = (w9902 & w13082) | (w9902 & w146) | (w13082 & w146);
assign w11698 = ~w17259 & ~w2971;
assign w11699 = w4877 & ~w8531;
assign w11700 = ~w3887 & ~w2720;
assign w11701 = ~w17778 & ~w2024;
assign w11702 = ~w5773 & ~w10075;
assign w11703 = w11413 & w7308;
assign w11704 = ~w10414 & w8724;
assign w11705 = a_15 & a_17;
assign w11706 = (w13979 & w17016) | (w13979 & w18842) | (w17016 & w18842);
assign w11707 = ~w6848 & ~w5580;
assign w11708 = ~w3220 & ~w1087;
assign w11709 = w6076 & w17468;
assign w11710 = ~w12273 & w12714;
assign w11711 = ~w379 & ~w2750;
assign w11712 = ~w3932 & ~w15109;
assign w11713 = w11211 & w7254;
assign w11714 = ~w2358 & ~w6869;
assign w11715 = ~w11539 & w9987;
assign w11716 = ~w1912 & ~w4654;
assign w11717 = ~w1417 & ~w13437;
assign w11718 = ~w1389 & ~w14554;
assign w11719 = ~w11262 & ~w12111;
assign w11720 = ~w18660 & w15889;
assign w11721 = ~w11511 & ~w3933;
assign w11722 = ~w12064 & ~w2305;
assign w11723 = ~w3087 & w9349;
assign w11724 = ~w4947 & ~w5988;
assign w11725 = a_14 & a_20;
assign w11726 = a_22 & a_33;
assign w11727 = ~w14922 & ~w10555;
assign w11728 = (~w5221 & ~w187) | (~w5221 & w13337) | (~w187 & w13337);
assign w11729 = ~w5513 & w3254;
assign w11730 = ~w15875 & ~w11110;
assign w11731 = ~w6220 & ~w11256;
assign w11732 = w17162 & ~w9637;
assign w11733 = w8214 & w19175;
assign w11734 = ~w2683 & ~w3816;
assign w11735 = (w6794 & w13082) | (w6794 & w4562) | (w13082 & w4562);
assign w11736 = a_29 & a_31;
assign w11737 = ~w7843 & ~w9599;
assign w11738 = ~w1732 & ~w17303;
assign w11739 = ~w19057 & ~w9004;
assign w11740 = ~w7819 & ~w12257;
assign w11741 = w14305 & w16503;
assign w11742 = ~w18383 & w17564;
assign w11743 = a_10 & a_18;
assign w11744 = w16338 & ~w6135;
assign w11745 = ~w16651 & ~w15078;
assign w11746 = ~w11178 & w80;
assign w11747 = ~w4045 & ~w15798;
assign w11748 = ~w6915 & w1221;
assign w11749 = w7148 & ~w2780;
assign w11750 = ~w9450 & ~w1203;
assign w11751 = ~w3340 & ~w11300;
assign w11752 = ~w11622 & ~w8209;
assign w11753 = ~w18005 & w10242;
assign w11754 = ~w13880 & ~w3397;
assign w11755 = ~w8032 & ~w9920;
assign w11756 = w6226 & ~w14800;
assign w11757 = ~w7764 & ~w15419;
assign w11758 = ~w3410 & ~w1809;
assign w11759 = ~w7099 & ~w1799;
assign w11760 = ~w19038 & ~w7345;
assign w11761 = ~w8028 & ~w9732;
assign w11762 = (~w7658 & ~w5549) | (~w7658 & w11768) | (~w5549 & w11768);
assign w11763 = ~w734 & w915;
assign w11764 = ~w15099 & ~w5075;
assign w11765 = a_39 & a_48;
assign w11766 = w7303 & ~w14604;
assign w11767 = ~w11336 & w579;
assign w11768 = w13907 & ~w7658;
assign w11769 = ~w6969 & w19047;
assign w11770 = ~w18489 & ~w15681;
assign w11771 = ~w8794 & ~w11534;
assign w11772 = ~w13190 & ~w16326;
assign w11773 = w10383 & w3924;
assign w11774 = w14615 & ~w1140;
assign w11775 = w2060 & ~w454;
assign w11776 = ~w7725 & ~w17863;
assign w11777 = ~w13562 & ~w11260;
assign w11778 = (~w4859 & ~w11976) | (~w4859 & w1469) | (~w11976 & w1469);
assign w11779 = ~w2390 & ~w7748;
assign w11780 = ~w8739 & w17378;
assign w11781 = w11705 & w13223;
assign w11782 = ~w8714 & ~w1072;
assign w11783 = ~w11833 & ~w15803;
assign w11784 = a_2 & a_17;
assign w11785 = a_30 & a_48;
assign w11786 = ~w1414 & ~w8441;
assign w11787 = ~w10231 & w3695;
assign w11788 = ~w4752 & ~w1297;
assign w11789 = ~w5050 & ~w1749;
assign w11790 = w6853 & w6948;
assign w11791 = a_7 & a_13;
assign w11792 = ~w10794 & ~w6710;
assign w11793 = w5063 & ~w13616;
assign w11794 = ~w16185 & ~w15129;
assign w11795 = w458 & ~w1124;
assign w11796 = ~w13750 & ~w3158;
assign w11797 = ~w2737 & ~w3003;
assign w11798 = ~w11064 & ~w8820;
assign w11799 = a_6 & a_59;
assign w11800 = w11972 & ~w5714;
assign w11801 = ~w2725 & w43;
assign w11802 = ~w15751 & ~w13988;
assign w11803 = ~w9064 & w4509;
assign w11804 = w11413 & ~w15722;
assign w11805 = w7462 & ~w9077;
assign w11806 = w13790 & w8146;
assign w11807 = ~w18324 & ~w10523;
assign w11808 = ~w11502 & ~w4475;
assign w11809 = w11791 & w11137;
assign w11810 = w18458 & ~w13339;
assign w11811 = w6723 & ~w2760;
assign w11812 = a_33 & a_56;
assign w11813 = a_23 & a_24;
assign w11814 = ~w3400 & w14779;
assign w11815 = w5007 & w12502;
assign w11816 = w4950 & ~w4245;
assign w11817 = w17421 & ~w17757;
assign w11818 = w14294 & ~w4945;
assign w11819 = ~w3901 & w9982;
assign w11820 = w6220 & w11256;
assign w11821 = w18740 & ~w16630;
assign w11822 = a_18 & a_52;
assign w11823 = (~w6085 & w15988) | (~w6085 & w10951) | (w15988 & w10951);
assign w11824 = ~w18626 & ~w6540;
assign w11825 = w15332 & ~w9784;
assign w11826 = ~w18928 & ~w5508;
assign w11827 = ~w2793 & w4032;
assign w11828 = ~w12688 & ~w18220;
assign w11829 = a_40 & a_51;
assign w11830 = ~w6925 & ~w16660;
assign w11831 = (~w16175 & ~w1962) | (~w16175 & w8496) | (~w1962 & w8496);
assign w11832 = ~w10 & w11484;
assign w11833 = w4649 & w8776;
assign w11834 = ~w6127 & ~w3817;
assign w11835 = ~w5772 & w10999;
assign w11836 = ~w6607 & ~w14802;
assign w11837 = ~w10431 & ~w8787;
assign w11838 = w1284 & ~w13441;
assign w11839 = ~w13834 & w5764;
assign w11840 = w19087 & w3778;
assign w11841 = w15591 & w9591;
assign w11842 = ~w18448 & ~w10910;
assign w11843 = ~w10356 & w11980;
assign w11844 = ~w1190 & ~w10703;
assign w11845 = a_34 & a_58;
assign w11846 = w10487 & w18874;
assign w11847 = w4279 & ~w6937;
assign w11848 = w14922 & ~w4717;
assign w11849 = ~w11272 & ~w19128;
assign w11850 = ~w3241 & ~w6418;
assign w11851 = ~w6062 & ~w18557;
assign w11852 = ~w978 & w14184;
assign w11853 = ~w18218 & w18654;
assign w11854 = w18459 & w7267;
assign w11855 = ~w9368 & ~w5591;
assign w11856 = w17450 & w18257;
assign w11857 = w13008 & ~w13770;
assign w11858 = ~w8903 & ~w5212;
assign w11859 = ~w347 & w16445;
assign w11860 = w2280 & ~w6563;
assign w11861 = ~w6829 & w19176;
assign w11862 = a_14 & a_22;
assign w11863 = (~w8454 & w1723) | (~w8454 & w13877) | (w1723 & w13877);
assign w11864 = (~w18087 & w18650) | (~w18087 & w17139) | (w18650 & w17139);
assign w11865 = a_1 & a_58;
assign w11866 = (~w4415 & ~w8207) | (~w4415 & w3679) | (~w8207 & w3679);
assign w11867 = w14332 & w12467;
assign w11868 = (~w17450 & w7015) | (~w17450 & w18608) | (w7015 & w18608);
assign w11869 = ~w15042 & w606;
assign w11870 = (~w15455 & ~w7080) | (~w15455 & w8202) | (~w7080 & w8202);
assign w11871 = ~w13273 & w12453;
assign w11872 = ~w9317 & ~w15375;
assign w11873 = ~w4619 & w18745;
assign w11874 = a_19 & a_35;
assign w11875 = w4022 & w2971;
assign w11876 = ~w9585 & w9556;
assign w11877 = ~w5613 & ~w9831;
assign w11878 = ~w2420 & w6305;
assign w11879 = a_2 & a_26;
assign w11880 = ~w13683 & w7745;
assign w11881 = ~w15433 & ~w590;
assign w11882 = ~w1901 & ~w2604;
assign w11883 = (~w6703 & ~w12536) | (~w6703 & w16841) | (~w12536 & w16841);
assign w11884 = w10737 & w15043;
assign w11885 = w6165 & ~w5496;
assign w11886 = w19110 & ~w10556;
assign w11887 = ~w18635 & ~w7016;
assign w11888 = ~w5235 & ~w162;
assign w11889 = a_37 & a_62;
assign w11890 = w9986 & ~w18386;
assign w11891 = w18769 & ~w2812;
assign w11892 = ~w9273 & ~w17527;
assign w11893 = ~w7335 & ~w12544;
assign w11894 = ~w12396 & ~w9075;
assign w11895 = w18052 & ~w7107;
assign w11896 = ~w9681 & w6188;
assign w11897 = a_49 & a_61;
assign w11898 = a_41 & a_59;
assign w11899 = ~w12296 & w4216;
assign w11900 = ~w15962 & ~w15216;
assign w11901 = ~w11907 & w1751;
assign w11902 = ~w14041 & w19122;
assign w11903 = ~w18051 & w7362;
assign w11904 = ~w14391 & ~w3257;
assign w11905 = ~w15290 & ~w2853;
assign w11906 = ~w16597 & w2919;
assign w11907 = ~w12722 & ~w13800;
assign w11908 = w14172 & w1906;
assign w11909 = ~w9384 & ~w14580;
assign w11910 = ~w11614 & ~w6502;
assign w11911 = ~w15592 & ~w8888;
assign w11912 = ~w7004 & w7736;
assign w11913 = ~w11988 & ~w13228;
assign w11914 = w7673 & w7604;
assign w11915 = ~w5017 & ~w2851;
assign w11916 = (w12679 & ~w18305) | (w12679 & w5910) | (~w18305 & w5910);
assign w11917 = ~w1206 & ~w7431;
assign w11918 = ~a_19 & ~w4687;
assign w11919 = ~w14478 & ~w5602;
assign w11920 = a_25 & a_32;
assign w11921 = ~w10017 & ~w5062;
assign w11922 = w18867 & w12712;
assign w11923 = w16016 & w8619;
assign w11924 = ~w3952 & w112;
assign w11925 = ~w14701 & ~w13446;
assign w11926 = w5927 & w11185;
assign w11927 = ~w16784 & ~w15946;
assign w11928 = w11417 & ~w17099;
assign w11929 = ~w14668 & ~w9852;
assign w11930 = w15877 & ~w7299;
assign w11931 = w3269 & w15747;
assign w11932 = ~w13059 & ~w14688;
assign w11933 = (~w261 & ~w13632) | (~w261 & w14610) | (~w13632 & w14610);
assign w11934 = ~w10249 & ~w8397;
assign w11935 = a_24 & a_34;
assign w11936 = w2883 & w9044;
assign w11937 = ~w15541 & w13994;
assign w11938 = w7875 & ~w15831;
assign w11939 = a_18 & a_49;
assign w11940 = ~w12725 & ~w10276;
assign w11941 = ~w5798 & ~w11124;
assign w11942 = w5195 & w12771;
assign w11943 = ~w9298 & ~w8516;
assign w11944 = a_8 & a_10;
assign w11945 = ~w10256 & ~w18641;
assign w11946 = ~w11391 & w500;
assign w11947 = w16706 & ~w9467;
assign w11948 = w8182 & ~w14391;
assign w11949 = (~w11446 & ~w15397) | (~w11446 & w480) | (~w15397 & w480);
assign w11950 = ~w7099 & w6309;
assign w11951 = ~w10109 & ~w2863;
assign w11952 = ~w5339 & ~w9826;
assign w11953 = ~w15084 & w3526;
assign w11954 = (~w15016 & ~w15415) | (~w15016 & w4805) | (~w15415 & w4805);
assign w11955 = ~w6230 & ~w7057;
assign w11956 = ~w9327 & w7184;
assign w11957 = ~w13202 & ~w18992;
assign w11958 = ~w1887 & w5150;
assign w11959 = w1700 & ~w17118;
assign w11960 = ~w2581 & ~w8582;
assign w11961 = a_23 & a_37;
assign w11962 = w7256 & w16571;
assign w11963 = w16738 & w15685;
assign w11964 = ~w19005 & w17711;
assign w11965 = a_25 & a_62;
assign w11966 = ~w12423 & w9141;
assign w11967 = ~w4494 & ~w2101;
assign w11968 = ~w12891 & ~w4917;
assign w11969 = (~w2769 & w12479) | (~w2769 & w7980) | (w12479 & w7980);
assign w11970 = ~w17886 & ~w12649;
assign w11971 = ~w12559 & w2643;
assign w11972 = ~w14281 & ~w7324;
assign w11973 = a_13 & a_41;
assign w11974 = ~w11350 & w16417;
assign w11975 = w10873 & ~w8747;
assign w11976 = ~w4859 & ~w9745;
assign w11977 = ~w11511 & ~w14702;
assign w11978 = w11147 & ~w10271;
assign w11979 = ~w6803 & ~w15572;
assign w11980 = ~w6501 & ~w2090;
assign w11981 = ~w9973 & ~w19145;
assign w11982 = ~w11139 & ~w7911;
assign w11983 = a_26 & a_37;
assign w11984 = ~w12160 & ~w18076;
assign w11985 = ~w11904 & w5985;
assign w11986 = w10030 & ~w15653;
assign w11987 = a_26 & a_28;
assign w11988 = ~w11754 & w10253;
assign w11989 = w4813 & w1470;
assign w11990 = a_30 & a_38;
assign w11991 = ~w12340 & ~w8179;
assign w11992 = w16144 & ~w8308;
assign w11993 = ~w17239 & ~w841;
assign w11994 = ~w12391 & ~w9031;
assign w11995 = (~w444 & ~w9371) | (~w444 & w18162) | (~w9371 & w18162);
assign w11996 = w14701 & ~w14723;
assign w11997 = ~w4069 & ~w1941;
assign w11998 = ~w8367 & ~w9744;
assign w11999 = (w17904 & ~w3925) | (w17904 & w3178) | (~w3925 & w3178);
assign w12000 = ~w13864 & ~w4359;
assign w12001 = (~w1205 & ~w14041) | (~w1205 & w14497) | (~w14041 & w14497);
assign w12002 = w9635 & w3325;
assign w12003 = ~w13634 & ~w13719;
assign w12004 = ~w16119 & ~w8680;
assign w12005 = ~w11428 & ~w9954;
assign w12006 = ~w14910 & ~w8977;
assign w12007 = ~w10919 & ~w4391;
assign w12008 = ~w15420 & ~w15999;
assign w12009 = ~w5917 & ~w2033;
assign w12010 = a_10 & a_42;
assign w12011 = ~w17443 & ~w7263;
assign w12012 = w13273 & ~w12453;
assign w12013 = ~w6272 & ~w12227;
assign w12014 = ~w15902 & w1159;
assign w12015 = ~w4340 & ~w3209;
assign w12016 = w17682 & ~w5566;
assign w12017 = ~w9409 & ~w1885;
assign w12018 = w3699 & ~w11722;
assign w12019 = ~w10937 & w7667;
assign w12020 = ~w5802 & ~w14125;
assign w12021 = a_1 & a_8;
assign w12022 = ~w8753 & ~w15649;
assign w12023 = (~w5032 & ~w1100) | (~w5032 & w7261) | (~w1100 & w7261);
assign w12024 = (~w9469 & ~w18024) | (~w9469 & w1544) | (~w18024 & w1544);
assign w12025 = ~w12180 & w13091;
assign w12026 = ~w7134 & w13482;
assign w12027 = ~w7443 & ~w11354;
assign w12028 = ~w9900 & ~w13600;
assign w12029 = ~w5009 & ~w1224;
assign w12030 = ~w18156 & w129;
assign w12031 = ~w15166 & ~w16050;
assign w12032 = w9176 & w435;
assign w12033 = w9395 & w8725;
assign w12034 = ~w13339 & ~w9827;
assign w12035 = (~w15301 & ~w17311) | (~w15301 & w18609) | (~w17311 & w18609);
assign w12036 = ~w1339 & ~w5350;
assign w12037 = ~w18206 & ~w4593;
assign w12038 = ~w16541 & ~w13751;
assign w12039 = ~w15909 & w7884;
assign w12040 = w10615 & w7544;
assign w12041 = ~w2461 & ~w3926;
assign w12042 = ~w10566 & ~w14003;
assign w12043 = ~w669 & w1017;
assign w12044 = ~w3653 & ~w2178;
assign w12045 = ~w4830 & ~w5877;
assign w12046 = ~w5761 & w10002;
assign w12047 = ~w5688 & w8872;
assign w12048 = ~w16828 & ~w7931;
assign w12049 = ~w6010 & ~w10502;
assign w12050 = ~w14545 & ~w6695;
assign w12051 = w10747 & w4165;
assign w12052 = ~w17807 & ~w9907;
assign w12053 = ~w18996 & w16953;
assign w12054 = w890 & w1229;
assign w12055 = ~w18959 & ~w17582;
assign w12056 = w7533 & w5241;
assign w12057 = ~w9583 & ~w2383;
assign w12058 = (~w14809 & ~w3036) | (~w14809 & w3218) | (~w3036 & w3218);
assign w12059 = w15975 & w1341;
assign w12060 = a_22 & a_40;
assign w12061 = w16673 & w1222;
assign w12062 = ~w8595 & w876;
assign w12063 = w5147 & w3983;
assign w12064 = ~w509 & ~w2987;
assign w12065 = ~w11287 & ~w3348;
assign w12066 = (w4287 & w10330) | (w4287 & w9432) | (w10330 & w9432);
assign w12067 = ~w1304 & ~w14427;
assign w12068 = w268 & w2439;
assign w12069 = a_13 & a_45;
assign w12070 = w151 & w5162;
assign w12071 = (w1894 & w13609) | (w1894 & w16356) | (w13609 & w16356);
assign w12072 = ~w7944 & ~w8929;
assign w12073 = a_27 & a_49;
assign w12074 = w7116 & w15656;
assign w12075 = (~w10257 & w1795) | (~w10257 & w742) | (w1795 & w742);
assign w12076 = ~w14697 & ~w10402;
assign w12077 = a_41 & a_51;
assign w12078 = ~w3798 & ~w18036;
assign w12079 = ~w11995 & w1893;
assign w12080 = ~w1450 & ~w14263;
assign w12081 = ~w623 & w16409;
assign w12082 = ~w4089 & ~w14079;
assign w12083 = a_1 & a_42;
assign w12084 = w7004 & ~w2735;
assign w12085 = ~w2983 & ~w12043;
assign w12086 = (w8250 & w11295) | (w8250 & w11244) | (w11295 & w11244);
assign w12087 = a_19 & a_49;
assign w12088 = ~w14028 & w463;
assign w12089 = ~w2769 & w9007;
assign w12090 = a_35 & a_49;
assign w12091 = ~w11268 & ~w13943;
assign w12092 = ~w19084 & ~w13425;
assign w12093 = ~w3325 & ~w769;
assign w12094 = w6146 & w10269;
assign w12095 = ~w16740 & w16768;
assign w12096 = ~w8624 & ~w9346;
assign w12097 = (w14457 & w18249) | (w14457 & w4913) | (w18249 & w4913);
assign w12098 = ~w6812 & ~w16667;
assign w12099 = (w19005 & w1399) | (w19005 & w18480) | (w1399 & w18480);
assign w12100 = w10845 & ~w9903;
assign w12101 = ~w9076 & ~w8801;
assign w12102 = ~w18654 & w18772;
assign w12103 = ~w2726 & ~w8007;
assign w12104 = ~w18383 & w6795;
assign w12105 = a_5 & a_29;
assign w12106 = w16320 & w5554;
assign w12107 = ~w4878 & ~w11304;
assign w12108 = (~w11591 & ~w13365) | (~w11591 & w8741) | (~w13365 & w8741);
assign w12109 = w4420 & w19199;
assign w12110 = ~w12284 & ~w18220;
assign w12111 = w8849 & w11824;
assign w12112 = a_6 & a_18;
assign w12113 = w12156 & ~w3532;
assign w12114 = ~w1585 & ~w2333;
assign w12115 = w1369 & w7372;
assign w12116 = ~w1408 & w4276;
assign w12117 = a_5 & a_13;
assign w12118 = ~w15421 & ~w1972;
assign w12119 = w14827 & ~w18538;
assign w12120 = ~w555 & ~w5170;
assign w12121 = ~w12136 & ~w13709;
assign w12122 = a_32 & a_60;
assign w12123 = w14306 & w14596;
assign w12124 = a_5 & a_55;
assign w12125 = ~w11858 & ~w14616;
assign w12126 = ~w4609 & ~w6099;
assign w12127 = w12834 & w5876;
assign w12128 = w4867 & w3573;
assign w12129 = ~w8444 & ~w7461;
assign w12130 = ~w15509 & ~w2117;
assign w12131 = a_8 & a_19;
assign w12132 = ~w8701 & ~w10219;
assign w12133 = ~w1139 & ~w12269;
assign w12134 = ~w15774 & ~w12833;
assign w12135 = w12235 & w9696;
assign w12136 = ~w8570 & ~w2985;
assign w12137 = ~w12081 & ~w16910;
assign w12138 = w17017 & ~w17617;
assign w12139 = ~w9908 & w15262;
assign w12140 = ~w154 & ~w8221;
assign w12141 = ~w2775 & ~w14870;
assign w12142 = ~w1777 & ~w15448;
assign w12143 = ~w17466 & w15187;
assign w12144 = ~w5135 & w3911;
assign w12145 = ~w653 & w18965;
assign w12146 = (~w19053 & w5341) | (~w19053 & w5729) | (w5341 & w5729);
assign w12147 = ~w16991 & ~w11821;
assign w12148 = ~w7724 & ~w11466;
assign w12149 = ~w15270 & ~w1788;
assign w12150 = a_9 & a_55;
assign w12151 = w4528 & ~w3555;
assign w12152 = ~w4097 & ~w15657;
assign w12153 = ~w5421 & ~w16582;
assign w12154 = ~w16178 & w13632;
assign w12155 = ~w13381 & w19096;
assign w12156 = ~w17692 & ~w17040;
assign w12157 = ~w17366 & ~w12139;
assign w12158 = w10059 & ~w13850;
assign w12159 = ~w8098 & w10004;
assign w12160 = w2139 & ~w18653;
assign w12161 = w1711 & w10390;
assign w12162 = ~w15617 & ~w9644;
assign w12163 = ~w6439 & ~w10093;
assign w12164 = ~w18393 & ~w1858;
assign w12165 = w13365 & ~w7270;
assign w12166 = w645 & w10181;
assign w12167 = w8424 & w17911;
assign w12168 = (w12404 & w6087) | (w12404 & w18128) | (w6087 & w18128);
assign w12169 = ~w2409 & ~w4197;
assign w12170 = a_3 & a_32;
assign w12171 = w341 & ~w765;
assign w12172 = (~w3882 & w2099) | (~w3882 & w14804) | (w2099 & w14804);
assign w12173 = ~w18874 & ~w9332;
assign w12174 = w16132 & w3648;
assign w12175 = w11455 & ~w8459;
assign w12176 = ~w14924 & ~w18574;
assign w12177 = ~w12219 & ~w5848;
assign w12178 = w1507 & w1101;
assign w12179 = w12673 & ~w18993;
assign w12180 = ~w5540 & ~w17704;
assign w12181 = w12664 & ~w517;
assign w12182 = w4878 & w11304;
assign w12183 = ~w1654 & w14579;
assign w12184 = ~w18584 & ~w2482;
assign w12185 = w11761 & ~w12333;
assign w12186 = w6839 & ~w6390;
assign w12187 = ~w2280 & w6563;
assign w12188 = w7352 & w11777;
assign w12189 = ~w16983 & ~w1819;
assign w12190 = ~w11405 & ~w13380;
assign w12191 = ~w17317 & ~w1428;
assign w12192 = w14770 & ~w19032;
assign w12193 = ~w9896 & w13473;
assign w12194 = w5760 & ~w11675;
assign w12195 = ~w14864 & w17383;
assign w12196 = w5864 & ~w17775;
assign w12197 = w10734 & w10270;
assign w12198 = w18383 & ~w2541;
assign w12199 = w15760 & w2284;
assign w12200 = ~w8648 & w13192;
assign w12201 = ~w7129 & w17661;
assign w12202 = ~w15630 & ~w4561;
assign w12203 = ~w15135 & w2166;
assign w12204 = w13423 & ~w270;
assign w12205 = w12039 & w15380;
assign w12206 = ~w13924 & w8772;
assign w12207 = a_21 & a_23;
assign w12208 = w6211 & ~w15863;
assign w12209 = ~w268 & ~w15366;
assign w12210 = (~w17934 & ~w7835) | (~w17934 & w6119) | (~w7835 & w6119);
assign w12211 = ~w8050 & ~w14007;
assign w12212 = w13450 & ~w1880;
assign w12213 = w18592 & w16909;
assign w12214 = ~w18787 & ~w2748;
assign w12215 = ~w5199 & w6400;
assign w12216 = ~w14505 & ~w3929;
assign w12217 = a_7 & a_34;
assign w12218 = w10737 & w15202;
assign w12219 = ~w14046 & ~w17239;
assign w12220 = a_1 & a_45;
assign w12221 = ~w14315 & ~w6900;
assign w12222 = a_20 & a_54;
assign w12223 = ~w14360 & ~w17033;
assign w12224 = ~w18833 & ~w3589;
assign w12225 = w16564 & ~w3987;
assign w12226 = ~w1743 & ~w11039;
assign w12227 = ~w7116 & ~w15656;
assign w12228 = w1983 & ~w5728;
assign w12229 = a_32 & a_34;
assign w12230 = ~w3973 & ~w10077;
assign w12231 = ~w19036 & w18499;
assign w12232 = ~w6186 & ~w8153;
assign w12233 = w9278 & w1361;
assign w12234 = w5623 & w16870;
assign w12235 = ~w2207 & ~w16426;
assign w12236 = a_39 & a_61;
assign w12237 = w8564 & ~w1658;
assign w12238 = ~w13887 & ~w17887;
assign w12239 = ~w12030 & ~w16003;
assign w12240 = ~w124 & ~w15346;
assign w12241 = ~w7979 & w18300;
assign w12242 = ~w6677 & w18026;
assign w12243 = ~w16404 & w15969;
assign w12244 = ~w12411 & w14185;
assign w12245 = ~w9254 & ~w11558;
assign w12246 = ~w11904 & w5003;
assign w12247 = ~w6032 & ~w14969;
assign w12248 = ~w13495 & ~w17565;
assign w12249 = ~w12697 & ~w11638;
assign w12250 = ~w14710 & ~w16509;
assign w12251 = ~w17660 & ~w7753;
assign w12252 = a_16 & a_28;
assign w12253 = ~w7223 & ~w7368;
assign w12254 = w17765 & ~w628;
assign w12255 = (w10242 & w5743) | (w10242 & w11753) | (w5743 & w11753);
assign w12256 = a_21 & a_26;
assign w12257 = w16767 & ~w3797;
assign w12258 = (w15755 & w3149) | (w15755 & w15239) | (w3149 & w15239);
assign w12259 = w16550 & w10451;
assign w12260 = ~w6736 & ~w10095;
assign w12261 = (w2254 & w11410) | (w2254 & w7583) | (w11410 & w7583);
assign w12262 = a_32 & a_44;
assign w12263 = ~w17188 & ~w4765;
assign w12264 = ~w4422 & ~w7874;
assign w12265 = w18837 & ~w10419;
assign w12266 = (~w13471 & ~w331) | (~w13471 & w10178) | (~w331 & w10178);
assign w12267 = ~w7771 & ~w16194;
assign w12268 = a_18 & a_39;
assign w12269 = ~w15492 & ~w10713;
assign w12270 = ~w16433 & ~w1028;
assign w12271 = a_16 & a_18;
assign w12272 = ~w71 & w11186;
assign w12273 = ~w14691 & ~w6612;
assign w12274 = a_28 & a_42;
assign w12275 = ~w8868 & ~w14549;
assign w12276 = w14138 & w977;
assign w12277 = w15310 & ~w1868;
assign w12278 = ~w2769 & w18002;
assign w12279 = ~w8587 & ~w8760;
assign w12280 = (~w8636 & ~w6335) | (~w8636 & w11576) | (~w6335 & w11576);
assign w12281 = w18975 & ~w16917;
assign w12282 = a_8 & a_56;
assign w12283 = ~w18539 & ~w9125;
assign w12284 = ~w1345 & ~w4438;
assign w12285 = ~w15029 & ~w7865;
assign w12286 = a_12 & a_49;
assign w12287 = ~w9619 & ~w4501;
assign w12288 = ~w666 & w15644;
assign w12289 = a_7 & a_27;
assign w12290 = ~w9581 & ~w7502;
assign w12291 = ~w3076 & ~w13320;
assign w12292 = ~w17977 & ~w19041;
assign w12293 = ~w8672 & ~w15853;
assign w12294 = ~w14798 & w932;
assign w12295 = ~w9560 & ~w6796;
assign w12296 = ~w10066 & ~w13951;
assign w12297 = ~w9074 & w5268;
assign w12298 = w16662 & ~w4733;
assign w12299 = ~w12305 & w3891;
assign w12300 = w14118 & ~w15712;
assign w12301 = a_7 & a_22;
assign w12302 = ~w8267 & w2100;
assign w12303 = w3418 & ~w15676;
assign w12304 = ~w4264 & ~w10706;
assign w12305 = ~w4047 & ~w12342;
assign w12306 = a_49 & a_57;
assign w12307 = w3064 & w16029;
assign w12308 = ~w5735 & ~w15228;
assign w12309 = w2447 & ~w16619;
assign w12310 = ~w12019 & w7233;
assign w12311 = ~w3711 & w11842;
assign w12312 = ~w980 & ~w7439;
assign w12313 = w9466 & ~w546;
assign w12314 = w8433 & ~w14986;
assign w12315 = ~w9753 & ~w7649;
assign w12316 = ~w17204 & w18354;
assign w12317 = ~w17410 & ~w11335;
assign w12318 = ~w17137 & ~w10882;
assign w12319 = ~w10925 & ~w6445;
assign w12320 = ~w15771 & w11010;
assign w12321 = ~w3360 & w11533;
assign w12322 = w16755 & ~w38;
assign w12323 = ~w12678 & w12283;
assign w12324 = a_13 & a_52;
assign w12325 = w11080 & ~w5344;
assign w12326 = ~w14907 & ~w12961;
assign w12327 = ~w6853 & w7253;
assign w12328 = w17119 & w12567;
assign w12329 = ~w5729 & w9893;
assign w12330 = w12452 & ~w5234;
assign w12331 = a_18 & a_58;
assign w12332 = a_37 & a_59;
assign w12333 = ~w13967 & ~w13779;
assign w12334 = (~w957 & ~w7777) | (~w957 & w15791) | (~w7777 & w15791);
assign w12335 = w12035 & w17512;
assign w12336 = ~w13801 & ~w13138;
assign w12337 = a_10 & a_11;
assign w12338 = w6708 & w2415;
assign w12339 = w10290 & w2504;
assign w12340 = ~w9452 & ~w3504;
assign w12341 = ~w5633 & ~w13340;
assign w12342 = ~w134 & w17345;
assign w12343 = ~w3590 & ~w5153;
assign w12344 = w12746 & ~w15145;
assign w12345 = ~w8331 & ~w16417;
assign w12346 = ~w1742 & ~w13793;
assign w12347 = ~w9250 & ~w499;
assign w12348 = w1030 & ~w7900;
assign w12349 = ~w593 & w6735;
assign w12350 = ~w10121 & ~w8579;
assign w12351 = ~w1272 & w2001;
assign w12352 = ~w7295 & w6243;
assign w12353 = w11126 & ~w4885;
assign w12354 = ~w8320 & w3454;
assign w12355 = w5067 & ~w13012;
assign w12356 = ~w18116 & ~w17286;
assign w12357 = ~w7952 & ~w15082;
assign w12358 = a_24 & a_42;
assign w12359 = ~w15992 & ~w11138;
assign w12360 = ~w18871 & ~w17159;
assign w12361 = ~w10865 & ~w2555;
assign w12362 = w7039 & ~w18446;
assign w12363 = ~w10855 & ~w17706;
assign w12364 = ~w8649 & ~w3875;
assign w12365 = (w7597 & w7610) | (w7597 & w5272) | (w7610 & w5272);
assign w12366 = ~w11689 & w16892;
assign w12367 = ~w2876 & w2833;
assign w12368 = ~w5981 & ~w683;
assign w12369 = w11127 & w10592;
assign w12370 = w11762 & ~w5044;
assign w12371 = ~w19007 & ~w18760;
assign w12372 = ~w2809 & w6049;
assign w12373 = ~w2026 & w10051;
assign w12374 = ~w14996 & ~w7991;
assign w12375 = ~w2485 & ~w9037;
assign w12376 = w13763 & ~w5967;
assign w12377 = ~w558 & w9113;
assign w12378 = ~a_62 & w10389;
assign w12379 = w14297 & ~w12187;
assign w12380 = ~w13778 & ~w16572;
assign w12381 = w9531 & w7179;
assign w12382 = ~w13702 & ~w13499;
assign w12383 = ~w7409 & w4529;
assign w12384 = ~w4100 & ~w14914;
assign w12385 = w11493 & w234;
assign w12386 = ~w17109 & w18144;
assign w12387 = w12532 & ~w1699;
assign w12388 = w8247 & w12358;
assign w12389 = w15837 & ~w9318;
assign w12390 = a_54 & a_61;
assign w12391 = ~w9842 & ~w4788;
assign w12392 = w1351 & ~w5786;
assign w12393 = ~w7361 & w13392;
assign w12394 = w13186 & w1576;
assign w12395 = ~w14722 & w1960;
assign w12396 = a_41 & a_63;
assign w12397 = w2547 & w12090;
assign w12398 = ~w2517 & w15583;
assign w12399 = w11455 & w7205;
assign w12400 = w11884 & ~w17604;
assign w12401 = ~w233 & w9888;
assign w12402 = w13763 & w5967;
assign w12403 = ~w16793 & ~w120;
assign w12404 = ~w2330 & w9759;
assign w12405 = ~w770 & ~w1484;
assign w12406 = (~w19123 & ~w19047) | (~w19123 & w7690) | (~w19047 & w7690);
assign w12407 = ~w11901 & ~w8811;
assign w12408 = w5352 & ~w17141;
assign w12409 = ~w6995 & ~w5168;
assign w12410 = ~w1723 & w8480;
assign w12411 = ~w11227 & ~w6659;
assign w12412 = w425 & w17248;
assign w12413 = w15937 & ~w6279;
assign w12414 = ~w13417 & ~w9036;
assign w12415 = w3319 & ~w15381;
assign w12416 = a_19 & a_45;
assign w12417 = ~w12427 & ~w9484;
assign w12418 = w1493 & w4822;
assign w12419 = ~w7129 & w3766;
assign w12420 = ~w9544 & ~w4929;
assign w12421 = ~w4065 & ~w14507;
assign w12422 = ~w8094 & ~w16527;
assign w12423 = ~w16969 & ~w17583;
assign w12424 = ~w8464 & ~w13900;
assign w12425 = w765 & ~w16012;
assign w12426 = a_12 & a_42;
assign w12427 = a_16 & a_45;
assign w12428 = w8367 & w9744;
assign w12429 = w4994 & w8910;
assign w12430 = a_46 & a_58;
assign w12431 = ~w3425 & w15574;
assign w12432 = w7232 & w5301;
assign w12433 = a_45 & a_49;
assign w12434 = w14875 & ~w6329;
assign w12435 = a_15 & a_26;
assign w12436 = ~w16560 & ~w13405;
assign w12437 = ~w2789 & ~w7184;
assign w12438 = w13284 & w6458;
assign w12439 = ~w3973 & ~w10894;
assign w12440 = (~w1711 & w11070) | (~w1711 & w2522) | (w11070 & w2522);
assign w12441 = ~w16192 & ~w3641;
assign w12442 = a_34 & a_57;
assign w12443 = a_9 & a_44;
assign w12444 = ~w15558 & ~w2940;
assign w12445 = ~w16849 & w6922;
assign w12446 = ~w6145 & ~w13235;
assign w12447 = a_41 & a_61;
assign w12448 = ~w15704 & w14666;
assign w12449 = w1923 & ~w6134;
assign w12450 = ~w15647 & ~w15986;
assign w12451 = ~w3361 & ~w3268;
assign w12452 = a_30 & a_47;
assign w12453 = ~w18692 & ~w4431;
assign w12454 = ~w6853 & w15337;
assign w12455 = ~w5010 & ~w5817;
assign w12456 = (w2254 & w5543) | (w2254 & w7802) | (w5543 & w7802);
assign w12457 = w5598 & w15447;
assign w12458 = w16595 & ~w2466;
assign w12459 = ~w12665 & ~w11048;
assign w12460 = ~w6896 & ~w4552;
assign w12461 = ~w16891 & ~w1375;
assign w12462 = w4350 & ~w13342;
assign w12463 = ~w1688 & w18679;
assign w12464 = ~w7017 & w12377;
assign w12465 = (~w1642 & ~w12542) | (~w1642 & w7468) | (~w12542 & w7468);
assign w12466 = ~w1275 & ~w16583;
assign w12467 = w18437 & ~w16476;
assign w12468 = (~w18532 & ~w3936) | (~w18532 & w2827) | (~w3936 & w2827);
assign w12469 = ~w14181 & w5596;
assign w12470 = w18832 & ~w1388;
assign w12471 = ~w866 & w6020;
assign w12472 = ~w19143 & ~w7541;
assign w12473 = ~w10491 & ~w6683;
assign w12474 = w17804 & ~w18226;
assign w12475 = ~w1158 & w4735;
assign w12476 = ~w16620 & ~w15641;
assign w12477 = a_23 & a_43;
assign w12478 = ~w3227 & w1335;
assign w12479 = ~w16896 & w19178;
assign w12480 = a_21 & a_51;
assign w12481 = ~w1677 & ~w8810;
assign w12482 = w13827 & ~w9198;
assign w12483 = ~w7506 & ~w4039;
assign w12484 = w1567 & w8802;
assign w12485 = a_3 & a_63;
assign w12486 = a_19 & a_37;
assign w12487 = w10773 & ~w13098;
assign w12488 = ~w14912 & ~w14319;
assign w12489 = a_4 & a_23;
assign w12490 = ~w1991 & ~w18919;
assign w12491 = (~w8267 & ~w18559) | (~w8267 & w14753) | (~w18559 & w14753);
assign w12492 = (~w10964 & ~w10926) | (~w10964 & w3697) | (~w10926 & w3697);
assign w12493 = ~w2182 & ~w8279;
assign w12494 = ~w12111 & ~w4934;
assign w12495 = ~w2889 & ~w8170;
assign w12496 = ~w5808 & ~w9738;
assign w12497 = a_23 & a_62;
assign w12498 = ~w7526 & w13549;
assign w12499 = w19141 & w1240;
assign w12500 = w9243 & w15804;
assign w12501 = ~w12100 & ~w15904;
assign w12502 = ~w15400 & ~w18250;
assign w12503 = a_19 & a_54;
assign w12504 = ~w12354 & w1459;
assign w12505 = ~w6656 & ~w12991;
assign w12506 = ~w1821 & w13670;
assign w12507 = ~w2891 & ~w15879;
assign w12508 = ~w4392 & ~w18570;
assign w12509 = ~w11510 & w12614;
assign w12510 = ~w372 & ~w6396;
assign w12511 = ~w5395 & w14905;
assign w12512 = ~a_51 & a_52;
assign w12513 = (~w2977 & ~w9077) | (~w2977 & w16694) | (~w9077 & w16694);
assign w12514 = a_4 & a_45;
assign w12515 = ~w15031 & ~w10525;
assign w12516 = a_8 & a_47;
assign w12517 = a_5 & a_23;
assign w12518 = w14517 & ~w6383;
assign w12519 = w7150 & w5166;
assign w12520 = ~w19022 & ~w1523;
assign w12521 = ~w3874 & ~w2494;
assign w12522 = w3966 & ~w8096;
assign w12523 = w5468 & w5875;
assign w12524 = w1300 & w18071;
assign w12525 = ~w14444 & ~w7887;
assign w12526 = ~w4018 & ~w1617;
assign w12527 = ~w3134 & w16142;
assign w12528 = ~w713 & w8526;
assign w12529 = ~w14974 & w10479;
assign w12530 = ~w7576 & w12513;
assign w12531 = w8306 & ~w6644;
assign w12532 = ~w15359 & ~w1461;
assign w12533 = ~w13276 & ~w8487;
assign w12534 = ~w1171 & ~w8511;
assign w12535 = ~w4226 & ~w7837;
assign w12536 = ~w6703 & ~w12381;
assign w12537 = a_12 & a_59;
assign w12538 = w6272 & w18645;
assign w12539 = a_9 & a_12;
assign w12540 = ~w12834 & ~w5876;
assign w12541 = ~w11469 & w2733;
assign w12542 = ~w1642 & ~w16851;
assign w12543 = ~w15630 & w16854;
assign w12544 = w9206 & ~w8422;
assign w12545 = ~w16975 & ~w16436;
assign w12546 = ~w14461 & ~w8920;
assign w12547 = (~w4774 & w15188) | (~w4774 & w12646) | (w15188 & w12646);
assign w12548 = w1967 & w2006;
assign w12549 = ~w2754 & ~w14657;
assign w12550 = ~w5387 & ~w4526;
assign w12551 = ~w5656 & ~w8204;
assign w12552 = ~w7646 & ~w10781;
assign w12553 = a_3 & a_37;
assign w12554 = ~w17671 & w15174;
assign w12555 = ~w15728 & ~w7398;
assign w12556 = ~w8911 & w16261;
assign w12557 = w15227 & ~w14139;
assign w12558 = ~w7378 & ~w8489;
assign w12559 = ~w16966 & ~w8705;
assign w12560 = ~w14864 & ~w9551;
assign w12561 = ~w2105 & ~w1337;
assign w12562 = a_16 & a_30;
assign w12563 = ~w5037 & ~w14941;
assign w12564 = w2880 & ~w16282;
assign w12565 = ~w15431 & ~w418;
assign w12566 = a_25 & a_59;
assign w12567 = ~w7531 & ~w7520;
assign w12568 = ~w14039 & ~w13942;
assign w12569 = w721 & ~w5974;
assign w12570 = ~w16888 & ~w10016;
assign w12571 = ~w14134 & ~w65;
assign w12572 = ~w5283 & ~w2830;
assign w12573 = ~w11337 & w1868;
assign w12574 = w2764 & w15177;
assign w12575 = ~w15695 & ~w9726;
assign w12576 = ~w18366 & ~w18743;
assign w12577 = ~w18304 & w3430;
assign w12578 = ~w14318 & ~w17032;
assign w12579 = ~w5547 & w12916;
assign w12580 = w11669 & w9126;
assign w12581 = w14944 & ~w12072;
assign w12582 = ~w11764 & ~w5652;
assign w12583 = ~w17390 & ~w12431;
assign w12584 = w6009 & w9183;
assign w12585 = w8942 & ~w17954;
assign w12586 = ~w476 & ~w17844;
assign w12587 = ~w6883 & w15707;
assign w12588 = ~w17664 & ~w9613;
assign w12589 = ~w19012 & ~w13835;
assign w12590 = ~w15470 & w5756;
assign w12591 = w5656 & ~w10652;
assign w12592 = ~w10153 & ~w11771;
assign w12593 = ~w17550 & ~w9171;
assign w12594 = ~w12369 & ~w2627;
assign w12595 = ~w9934 & ~w9701;
assign w12596 = ~w13290 & w9962;
assign w12597 = ~w1078 & ~w15279;
assign w12598 = w13070 & ~w9594;
assign w12599 = ~w18137 & ~w1757;
assign w12600 = ~w11107 & w17479;
assign w12601 = a_12 & a_62;
assign w12602 = w10737 & w469;
assign w12603 = ~w533 & ~w6592;
assign w12604 = ~w547 & w16341;
assign w12605 = ~w7139 & ~w11881;
assign w12606 = a_37 & a_60;
assign w12607 = w8721 & ~w5400;
assign w12608 = ~w7747 & w19006;
assign w12609 = ~w8640 & ~w6666;
assign w12610 = ~w8400 & w12422;
assign w12611 = w18682 & ~w9974;
assign w12612 = a_14 & a_44;
assign w12613 = w9247 & w324;
assign w12614 = ~w8857 & ~w14175;
assign w12615 = w15552 & ~w15192;
assign w12616 = (w9221 & w8255) | (w9221 & w4352) | (w8255 & w4352);
assign w12617 = a_36 & a_43;
assign w12618 = w17248 & ~w16739;
assign w12619 = ~w269 & w10952;
assign w12620 = ~w13298 & ~w12756;
assign w12621 = w111 & ~w4141;
assign w12622 = a_33 & a_61;
assign w12623 = ~w12313 & ~w2146;
assign w12624 = ~w9094 & ~w1265;
assign w12625 = ~w11610 & ~w11099;
assign w12626 = ~w18826 & ~w9038;
assign w12627 = w18732 & ~w1083;
assign w12628 = w16669 & w7417;
assign w12629 = w1845 & w5253;
assign w12630 = ~w1183 & ~w12272;
assign w12631 = w16558 & w3812;
assign w12632 = w9802 & ~w14819;
assign w12633 = ~w4027 & ~w15564;
assign w12634 = ~w15598 & ~w1327;
assign w12635 = w13745 & w6578;
assign w12636 = ~w14012 & w4620;
assign w12637 = a_26 & a_36;
assign w12638 = ~w1762 & ~w18400;
assign w12639 = w9315 & w9756;
assign w12640 = (~w2507 & ~w18899) | (~w2507 & w12858) | (~w18899 & w12858);
assign w12641 = a_2 & a_24;
assign w12642 = w15909 & ~w7884;
assign w12643 = w18028 & w10904;
assign w12644 = ~w19115 & w3291;
assign w12645 = ~w6409 & w8183;
assign w12646 = w2973 & ~w4774;
assign w12647 = (~w16282 & ~w14280) | (~w16282 & w12564) | (~w14280 & w12564);
assign w12648 = a_27 & a_33;
assign w12649 = a_13 & a_53;
assign w12650 = ~w13880 & ~w17057;
assign w12651 = ~w4474 & ~w3841;
assign w12652 = ~w738 & ~w11090;
assign w12653 = ~w10875 & w18268;
assign w12654 = ~w5461 & ~w339;
assign w12655 = w5961 & ~w15952;
assign w12656 = ~w9407 & ~w10332;
assign w12657 = ~w13347 & ~w7818;
assign w12658 = ~w5697 & w14495;
assign w12659 = w3161 & ~w1152;
assign w12660 = w18209 & ~w15342;
assign w12661 = w7389 & w8773;
assign w12662 = ~w8555 & w2614;
assign w12663 = ~w11146 & w7436;
assign w12664 = ~w1579 & ~w3389;
assign w12665 = w18488 & ~w8918;
assign w12666 = ~w17355 & ~w17437;
assign w12667 = a_25 & a_55;
assign w12668 = w1953 & ~w9291;
assign w12669 = w7114 & ~w693;
assign w12670 = w14231 & ~w15993;
assign w12671 = ~w3801 & ~w2416;
assign w12672 = ~w5912 & ~w7422;
assign w12673 = ~w14352 & ~w3280;
assign w12674 = w12925 & w13284;
assign w12675 = a_24 & a_46;
assign w12676 = w8917 & ~w9684;
assign w12677 = ~w8588 & w6845;
assign w12678 = a_53 & a_59;
assign w12679 = ~w16534 & ~w6025;
assign w12680 = ~w14992 & ~w6977;
assign w12681 = ~w13036 & w2210;
assign w12682 = w4846 & ~w15762;
assign w12683 = ~w7950 & ~w3578;
assign w12684 = w12917 & ~w3806;
assign w12685 = ~w4739 & w11322;
assign w12686 = a_12 & a_16;
assign w12687 = w15789 & ~w8067;
assign w12688 = a_2 & a_31;
assign w12689 = (~w3700 & w10330) | (~w3700 & w3011) | (w10330 & w3011);
assign w12690 = ~w7712 & ~w7898;
assign w12691 = ~w17787 & ~w14198;
assign w12692 = ~w11689 & ~w7825;
assign w12693 = a_27 & a_39;
assign w12694 = w10225 & ~w1333;
assign w12695 = ~w12558 & w3318;
assign w12696 = ~w10042 & ~w11743;
assign w12697 = a_2 & a_59;
assign w12698 = a_29 & a_39;
assign w12699 = (~w9732 & ~w11761) | (~w9732 & w11407) | (~w11761 & w11407);
assign w12700 = ~w9420 & w16857;
assign w12701 = ~w2010 & ~w10426;
assign w12702 = w7060 & ~w19052;
assign w12703 = (~w6466 & ~w3955) | (~w6466 & w11513) | (~w3955 & w11513);
assign w12704 = ~w13217 & w1268;
assign w12705 = w4585 & ~w7053;
assign w12706 = w8848 & ~w16212;
assign w12707 = ~w18671 & ~w10838;
assign w12708 = (w15329 & w1974) | (w15329 & w1086) | (w1974 & w1086);
assign w12709 = w17037 & ~w13076;
assign w12710 = w12553 & w2423;
assign w12711 = ~w13744 & w3323;
assign w12712 = ~w12448 & ~w3981;
assign w12713 = ~w1117 & ~w14960;
assign w12714 = ~w11744 & ~w10394;
assign w12715 = w3777 & ~w14656;
assign w12716 = ~w10119 & w13959;
assign w12717 = ~w17499 & ~w16943;
assign w12718 = ~w7967 & w450;
assign w12719 = (~w4070 & ~w8319) | (~w4070 & w11027) | (~w8319 & w11027);
assign w12720 = ~w4022 & ~w966;
assign w12721 = ~w15456 & w12563;
assign w12722 = w15168 & w15682;
assign w12723 = ~w11707 & w2758;
assign w12724 = ~w13055 & ~w16108;
assign w12725 = a_44 & a_58;
assign w12726 = ~w14173 & ~w3860;
assign w12727 = ~w13329 & ~w11817;
assign w12728 = ~w10565 & ~w10464;
assign w12729 = w80 & ~w17633;
assign w12730 = w4691 & ~w3262;
assign w12731 = ~w14822 & w17509;
assign w12732 = w15902 & ~w1159;
assign w12733 = ~w649 & ~w8536;
assign w12734 = w6085 & w12239;
assign w12735 = a_14 & a_35;
assign w12736 = ~w6534 & ~w2088;
assign w12737 = ~w17579 & ~w9976;
assign w12738 = ~w16914 & ~w13334;
assign w12739 = ~w17628 & ~w9633;
assign w12740 = ~w8460 & ~w18317;
assign w12741 = w17375 & ~w1263;
assign w12742 = ~w12035 & ~w17512;
assign w12743 = ~w8842 & ~w11474;
assign w12744 = w6474 & w7550;
assign w12745 = ~w13685 & ~w6572;
assign w12746 = ~w1414 & ~w3743;
assign w12747 = ~w16952 & ~w6997;
assign w12748 = ~w2113 & ~w12549;
assign w12749 = ~w5336 & ~w17235;
assign w12750 = w18330 & ~w8288;
assign w12751 = ~w16764 & ~w14411;
assign w12752 = w201 & ~w11588;
assign w12753 = a_19 & a_60;
assign w12754 = (w18365 & w17323) | (w18365 & w7917) | (w17323 & w7917);
assign w12755 = ~w1899 & ~w8742;
assign w12756 = ~w2544 & ~w7481;
assign w12757 = ~w1405 & ~w8734;
assign w12758 = a_12 & a_41;
assign w12759 = w6656 & w13232;
assign w12760 = ~w17366 & ~w9908;
assign w12761 = a_24 & a_54;
assign w12762 = ~w2779 & ~w103;
assign w12763 = ~w15532 & w17084;
assign w12764 = w8800 & ~w12214;
assign w12765 = ~w10697 & w3836;
assign w12766 = (w16033 & w2769) | (w16033 & w6913) | (w2769 & w6913);
assign w12767 = ~w1705 & ~w7561;
assign w12768 = ~w17155 & ~w674;
assign w12769 = a_6 & a_36;
assign w12770 = (w1363 & w17770) | (w1363 & w10575) | (w17770 & w10575);
assign w12771 = ~w16899 & ~w1565;
assign w12772 = ~w8873 & w992;
assign w12773 = ~w10330 & w16989;
assign w12774 = w16482 & w13868;
assign w12775 = w11586 & w3902;
assign w12776 = (~w9739 & ~w5116) | (~w9739 & w852) | (~w5116 & w852);
assign w12777 = w8547 & w1889;
assign w12778 = w3489 & ~w8401;
assign w12779 = ~w7705 & ~w5494;
assign w12780 = w5203 & ~w1823;
assign w12781 = ~w1975 & ~w14632;
assign w12782 = ~w9481 & w9274;
assign w12783 = w11728 & ~w16635;
assign w12784 = w7764 & ~w7395;
assign w12785 = ~w18732 & w1083;
assign w12786 = w2609 & ~w14888;
assign w12787 = ~w6108 & w12582;
assign w12788 = ~w9635 & ~w3325;
assign w12789 = ~w4038 & ~w13416;
assign w12790 = a_5 & a_49;
assign w12791 = ~w2930 & ~w9661;
assign w12792 = ~w3236 & w3556;
assign w12793 = w15785 & ~w8832;
assign w12794 = w5865 & w3757;
assign w12795 = (~w16336 & ~w3143) | (~w16336 & w9335) | (~w3143 & w9335);
assign w12796 = w16590 & ~w12279;
assign w12797 = a_23 & a_48;
assign w12798 = w3499 & w9546;
assign w12799 = ~w12061 & ~w6314;
assign w12800 = w12565 & ~w11917;
assign w12801 = ~w17078 & ~w8506;
assign w12802 = ~w18329 & ~w15668;
assign w12803 = ~w16468 & ~w12429;
assign w12804 = ~w7890 & ~w10936;
assign w12805 = ~w13180 & ~w16158;
assign w12806 = w6715 & ~w8967;
assign w12807 = ~w200 & ~w3642;
assign w12808 = w17451 & w13349;
assign w12809 = w15520 & ~w446;
assign w12810 = a_17 & a_37;
assign w12811 = ~w5347 & ~w10816;
assign w12812 = ~w16707 & ~w11267;
assign w12813 = w14906 & ~w4038;
assign w12814 = ~w5859 & ~w5112;
assign w12815 = w4011 & ~w7302;
assign w12816 = w3675 & ~w229;
assign w12817 = ~w12252 & ~w9575;
assign w12818 = (~w12245 & ~w17421) | (~w12245 & w2768) | (~w17421 & w2768);
assign w12819 = ~w18918 & ~w6621;
assign w12820 = (~w3052 & ~w19011) | (~w3052 & w14735) | (~w19011 & w14735);
assign w12821 = ~w10127 & ~w2058;
assign w12822 = ~w18232 & ~w12799;
assign w12823 = ~w3864 & w8864;
assign w12824 = w9478 & ~w13396;
assign w12825 = ~w17654 & ~w11854;
assign w12826 = w4267 & ~w16083;
assign w12827 = ~w15238 & w15730;
assign w12828 = ~w6162 & ~w9748;
assign w12829 = w1904 & ~w1847;
assign w12830 = (w7436 & w2769) | (w7436 & w12663) | (w2769 & w12663);
assign w12831 = w14101 & ~w18616;
assign w12832 = ~w15616 & ~w14;
assign w12833 = (w18091 & w16133) | (w18091 & w8311) | (w16133 & w8311);
assign w12834 = ~w15883 & ~w1968;
assign w12835 = ~w16738 & ~w15685;
assign w12836 = ~w2704 & ~w19000;
assign w12837 = ~w8597 & ~w13867;
assign w12838 = ~w11862 & ~w13239;
assign w12839 = w503 & ~w8978;
assign w12840 = ~w5820 & ~w3599;
assign w12841 = (~w5350 & ~w13072) | (~w5350 & w12036) | (~w13072 & w12036);
assign w12842 = ~w13135 & w5681;
assign w12843 = w16299 & w8770;
assign w12844 = ~w10926 & ~w2978;
assign w12845 = ~w15985 & ~w12551;
assign w12846 = w5095 & ~w16192;
assign w12847 = ~w15586 & ~w3945;
assign w12848 = ~w18121 & ~w18658;
assign w12849 = ~w2269 & w10027;
assign w12850 = ~w14157 & ~w1442;
assign w12851 = ~w16951 & w18573;
assign w12852 = ~w10499 & ~w7189;
assign w12853 = ~w11255 & ~w16982;
assign w12854 = w2916 & w19179;
assign w12855 = ~w10472 & ~w9379;
assign w12856 = ~w13987 & ~w13507;
assign w12857 = a_58 & a_60;
assign w12858 = ~w5169 & ~w2507;
assign w12859 = ~w3668 & w9193;
assign w12860 = w2449 & w9883;
assign w12861 = ~w10012 & ~w14781;
assign w12862 = a_17 & a_46;
assign w12863 = a_34 & a_40;
assign w12864 = ~w9757 & ~w17460;
assign w12865 = w7411 & ~w8616;
assign w12866 = ~w9060 & ~w10375;
assign w12867 = ~w11200 & ~w11144;
assign w12868 = ~w18369 & ~w9032;
assign w12869 = a_3 & a_20;
assign w12870 = w11439 & ~w3904;
assign w12871 = ~w1996 & ~w13127;
assign w12872 = w3129 & ~w14263;
assign w12873 = ~w3666 & ~w8634;
assign w12874 = ~w7992 & w9174;
assign w12875 = ~w6541 & ~w8066;
assign w12876 = w7266 & w3031;
assign w12877 = a_4 & a_5;
assign w12878 = ~w963 & w6802;
assign w12879 = ~w14130 & w15481;
assign w12880 = w16201 & w9072;
assign w12881 = ~w1892 & ~w11685;
assign w12882 = (~w1203 & ~w6520) | (~w1203 & w11750) | (~w6520 & w11750);
assign w12883 = (w1508 & w12718) | (w1508 & w14823) | (w12718 & w14823);
assign w12884 = ~w11448 & ~w7930;
assign w12885 = ~w7392 & ~w8370;
assign w12886 = ~w18779 & ~w15406;
assign w12887 = ~w16015 & w4583;
assign w12888 = ~w19100 & ~w16623;
assign w12889 = w1045 & ~w3144;
assign w12890 = w5660 & w15408;
assign w12891 = ~w12705 & ~w9196;
assign w12892 = ~w15296 & ~w12528;
assign w12893 = a_2 & a_61;
assign w12894 = ~w12152 & ~w18312;
assign w12895 = w4610 & w8359;
assign w12896 = w12207 & w6083;
assign w12897 = (w7356 & w16593) | (w7356 & w14777) | (w16593 & w14777);
assign w12898 = ~w3817 & ~w16549;
assign w12899 = ~w1948 & ~w15852;
assign w12900 = a_37 & a_48;
assign w12901 = ~w16516 & ~w11758;
assign w12902 = ~w5123 & w4380;
assign w12903 = w1454 & w7982;
assign w12904 = ~w16857 & w12243;
assign w12905 = ~w9239 & ~w12217;
assign w12906 = ~w18571 & w10413;
assign w12907 = a_16 & a_55;
assign w12908 = ~w16362 & w11182;
assign w12909 = w6117 & ~w4762;
assign w12910 = ~w2061 & ~w5861;
assign w12911 = (~w8679 & ~w4944) | (~w8679 & w6414) | (~w4944 & w6414);
assign w12912 = w3487 & ~w11020;
assign w12913 = w14216 & ~w18399;
assign w12914 = ~w10105 & ~w8669;
assign w12915 = w6158 & ~w3911;
assign w12916 = ~w7454 & ~w9345;
assign w12917 = (w7268 & w18852) | (w7268 & w7713) | (w18852 & w7713);
assign w12918 = w14444 & w1400;
assign w12919 = a_20 & a_34;
assign w12920 = ~w8643 & ~w12254;
assign w12921 = ~w4641 & w15940;
assign w12922 = w3121 & ~w12130;
assign w12923 = ~w14118 & w15712;
assign w12924 = ~w1969 & ~w2935;
assign w12925 = a_17 & a_53;
assign w12926 = ~w13762 & ~w12263;
assign w12927 = w14827 & ~w9923;
assign w12928 = ~w10607 & w1518;
assign w12929 = ~w15814 & ~w9564;
assign w12930 = ~w5637 & ~w1456;
assign w12931 = ~w6558 & ~w1768;
assign w12932 = (~w8727 & ~w18330) | (~w8727 & w5427) | (~w18330 & w5427);
assign w12933 = ~w2529 & ~w2149;
assign w12934 = ~w14912 & ~w19090;
assign w12935 = ~w5962 & ~w11424;
assign w12936 = ~w16565 & w5154;
assign w12937 = w5761 & ~w10002;
assign w12938 = ~w6060 & ~w10630;
assign w12939 = ~w17685 & ~w16250;
assign w12940 = ~w10927 & ~w12643;
assign w12941 = (~w14320 & ~w9567) | (~w14320 & w10164) | (~w9567 & w10164);
assign w12942 = ~w16113 & w568;
assign w12943 = w13595 & w19180;
assign w12944 = w4883 & ~w2234;
assign w12945 = ~w10157 & ~w12047;
assign w12946 = ~w788 & ~w14726;
assign w12947 = w18190 & w8023;
assign w12948 = ~w7846 & ~w3182;
assign w12949 = w12010 & ~w12969;
assign w12950 = ~w8584 & w16088;
assign w12951 = ~w14150 & w2370;
assign w12952 = w13648 & ~w2070;
assign w12953 = (w17582 & w12355) | (w17582 & w2934) | (w12355 & w2934);
assign w12954 = (w14256 & w2769) | (w14256 & w7693) | (w2769 & w7693);
assign w12955 = w13973 & ~w5053;
assign w12956 = ~w5763 & ~w5640;
assign w12957 = a_31 & a_53;
assign w12958 = ~w4757 & ~w49;
assign w12959 = (~w7022 & w7768) | (~w7022 & w7028) | (w7768 & w7028);
assign w12960 = ~w12723 & ~w4410;
assign w12961 = ~w5931 & ~w1926;
assign w12962 = ~w16442 & ~w3333;
assign w12963 = ~w2885 & ~w18337;
assign w12964 = ~w950 & ~w1997;
assign w12965 = ~w10940 & ~w16801;
assign w12966 = a_32 & a_35;
assign w12967 = ~w3162 & ~w1289;
assign w12968 = ~w13148 & ~w11303;
assign w12969 = ~w4864 & ~w2076;
assign w12970 = ~w1936 & ~w4176;
assign w12971 = a_13 & a_36;
assign w12972 = ~w14031 & w7770;
assign w12973 = ~w5168 & w18093;
assign w12974 = ~w1845 & ~w17104;
assign w12975 = (w10309 & w2849) | (w10309 & w14989) | (w2849 & w14989);
assign w12976 = w16481 & ~w9711;
assign w12977 = ~w11813 & ~w1192;
assign w12978 = ~w10765 & ~w3667;
assign w12979 = w941 & w5023;
assign w12980 = ~w3818 & ~w6916;
assign w12981 = w2876 & ~w2833;
assign w12982 = ~w14814 & w15287;
assign w12983 = ~w882 & ~w13330;
assign w12984 = ~w5623 & ~w16870;
assign w12985 = ~w17442 & ~w4469;
assign w12986 = w8930 & ~w27;
assign w12987 = a_42 & a_51;
assign w12988 = ~w12867 & w16614;
assign w12989 = w6163 & w6843;
assign w12990 = ~w2616 & ~w2231;
assign w12991 = ~w8089 & w2651;
assign w12992 = ~w296 & ~w9473;
assign w12993 = ~w3591 & w15093;
assign w12994 = ~w7942 & ~w12569;
assign w12995 = ~w977 & ~w5738;
assign w12996 = ~w2900 & ~w10750;
assign w12997 = a_25 & a_40;
assign w12998 = (~w17633 & ~w11178) | (~w17633 & w12729) | (~w11178 & w12729);
assign w12999 = ~w12430 & w7908;
assign w13000 = ~w6972 & ~w1479;
assign w13001 = ~w1873 & ~w13790;
assign w13002 = ~w13082 & w6957;
assign w13003 = a_14 & a_43;
assign w13004 = w2563 & ~w11206;
assign w13005 = ~w4193 & ~w4903;
assign w13006 = a_34 & a_62;
assign w13007 = w4367 & w19181;
assign w13008 = a_22 & a_27;
assign w13009 = (~w1610 & ~w15897) | (~w1610 & w8994) | (~w15897 & w8994);
assign w13010 = ~w10861 & w13845;
assign w13011 = a_41 & a_56;
assign w13012 = (~w4560 & ~w8101) | (~w4560 & w8898) | (~w8101 & w8898);
assign w13013 = ~w9376 & ~w11365;
assign w13014 = ~w14862 & ~w910;
assign w13015 = ~w5147 & ~w3983;
assign w13016 = a_19 & a_27;
assign w13017 = w12738 & ~w14791;
assign w13018 = (w13422 & w263) | (w13422 & w7315) | (w263 & w7315);
assign w13019 = w4546 & ~w18555;
assign w13020 = ~w14628 & ~w16711;
assign w13021 = ~w8861 & ~w4803;
assign w13022 = w8600 & ~w16586;
assign w13023 = ~w5397 & w18126;
assign w13024 = ~w5059 & ~w17390;
assign w13025 = ~w12235 & ~w9696;
assign w13026 = ~w4071 & ~w11678;
assign w13027 = ~w15530 & ~w8683;
assign w13028 = ~w3508 & ~w15391;
assign w13029 = ~w6207 & ~w4026;
assign w13030 = ~w3444 & ~w6483;
assign w13031 = ~w16615 & ~w17973;
assign w13032 = w116 & w8103;
assign w13033 = ~w8052 & w6693;
assign w13034 = ~w14364 & w15352;
assign w13035 = ~w3275 & ~w2944;
assign w13036 = a_24 & a_63;
assign w13037 = w15575 & w1003;
assign w13038 = ~w550 & ~w1245;
assign w13039 = ~w6133 & ~w15870;
assign w13040 = ~w7909 & ~w2476;
assign w13041 = ~w1661 & w17674;
assign w13042 = w14171 & ~w12779;
assign w13043 = ~w14998 & ~w8716;
assign w13044 = w6513 & w12911;
assign w13045 = ~w4180 & ~w3919;
assign w13046 = ~w15668 & ~w2539;
assign w13047 = w16389 & ~w10436;
assign w13048 = ~w5503 & ~w8526;
assign w13049 = ~w2938 & ~w1917;
assign w13050 = ~w2576 & ~w9577;
assign w13051 = ~w13840 & ~w1058;
assign w13052 = ~w14172 & w15463;
assign w13053 = ~w5943 & w6994;
assign w13054 = ~w15792 & ~w7478;
assign w13055 = w6786 & w9435;
assign w13056 = ~w15976 & ~w18778;
assign w13057 = ~w2716 & ~w17144;
assign w13058 = a_18 & a_38;
assign w13059 = ~w12583 & ~w4571;
assign w13060 = w12380 & w11560;
assign w13061 = a_44 & a_52;
assign w13062 = w2725 & w4478;
assign w13063 = ~w12547 & ~w9875;
assign w13064 = ~w5217 & ~w1645;
assign w13065 = ~w13078 & ~w16945;
assign w13066 = ~w4863 & w2347;
assign w13067 = ~w9681 & ~w17712;
assign w13068 = ~w14783 & w4146;
assign w13069 = ~w6864 & ~w2832;
assign w13070 = ~w14977 & ~w12875;
assign w13071 = w15397 & ~w10038;
assign w13072 = ~w5350 & ~w13638;
assign w13073 = (~w16365 & ~w286) | (~w16365 & w1491) | (~w286 & w1491);
assign w13074 = ~w8874 & w10690;
assign w13075 = a_12 & a_48;
assign w13076 = ~w11628 & ~w17447;
assign w13077 = ~w3799 & ~w12945;
assign w13078 = a_15 & a_44;
assign w13079 = ~w905 & ~w11500;
assign w13080 = (~w10271 & ~w8505) | (~w10271 & w11978) | (~w8505 & w11978);
assign w13081 = w15560 & w14460;
assign w13082 = ~w7409 & w16086;
assign w13083 = ~w5433 & ~w1342;
assign w13084 = w17657 & w16698;
assign w13085 = w14193 & ~w4953;
assign w13086 = a_24 & a_40;
assign w13087 = ~w12433 & w9182;
assign w13088 = ~w5771 & ~w743;
assign w13089 = w11192 & ~w3470;
assign w13090 = w16562 & ~w5509;
assign w13091 = ~w16140 & ~w5431;
assign w13092 = ~w4203 & ~w839;
assign w13093 = ~w267 & ~w12487;
assign w13094 = ~w15328 & ~w17771;
assign w13095 = (~w90 & ~w15074) | (~w90 & w13978) | (~w15074 & w13978);
assign w13096 = ~w1784 & ~w14148;
assign w13097 = w89 & ~w888;
assign w13098 = ~w9491 & ~w1550;
assign w13099 = ~w6709 & w18659;
assign w13100 = ~w9506 & w7296;
assign w13101 = ~w2043 & ~w4418;
assign w13102 = ~w5176 & w11590;
assign w13103 = ~w8551 & ~w7198;
assign w13104 = ~w13259 & ~w16520;
assign w13105 = ~w18468 & ~w5945;
assign w13106 = a_41 & a_48;
assign w13107 = ~w7554 & ~w2345;
assign w13108 = ~w4010 & ~w4183;
assign w13109 = ~w14534 & ~w8659;
assign w13110 = ~w11480 & ~w16894;
assign w13111 = ~w15532 & ~w1047;
assign w13112 = w8711 & w12289;
assign w13113 = ~w2053 & ~w18173;
assign w13114 = ~w18950 & ~w5634;
assign w13115 = ~w2950 & ~w988;
assign w13116 = ~w3840 & ~w15640;
assign w13117 = (~w5811 & w11532) | (~w5811 & w11572) | (w11532 & w11572);
assign w13118 = (~w15213 & w7979) | (~w15213 & w2890) | (w7979 & w2890);
assign w13119 = ~w12888 & ~w917;
assign w13120 = ~w7643 & ~w17494;
assign w13121 = ~w6564 & w13360;
assign w13122 = ~w194 & ~w11004;
assign w13123 = a_1 & a_16;
assign w13124 = ~w13498 & ~w1015;
assign w13125 = a_22 & a_29;
assign w13126 = (~w17101 & w17665) | (~w17101 & w13706) | (w17665 & w13706);
assign w13127 = ~w16235 & ~w15441;
assign w13128 = w2468 & ~w15634;
assign w13129 = w4553 & w10090;
assign w13130 = ~w17729 & ~w6107;
assign w13131 = ~w13433 & ~w881;
assign w13132 = ~w8312 & ~w6239;
assign w13133 = ~w17070 & ~w6508;
assign w13134 = ~w3168 & ~w4719;
assign w13135 = ~w14747 & ~w3723;
assign w13136 = ~w14134 & w15482;
assign w13137 = ~w7599 & ~w13209;
assign w13138 = ~w4171 & ~w15120;
assign w13139 = a_23 & a_44;
assign w13140 = ~w1099 & ~w8543;
assign w13141 = w14418 & ~w7913;
assign w13142 = a_48 & a_58;
assign w13143 = ~w1687 & w13590;
assign w13144 = ~w10594 & ~w17828;
assign w13145 = ~w14462 & ~w12568;
assign w13146 = ~w13073 & w3958;
assign w13147 = w9898 & w6137;
assign w13148 = a_23 & a_51;
assign w13149 = ~w5278 & ~w15805;
assign w13150 = ~w6656 & ~w18875;
assign w13151 = a_13 & w17557;
assign w13152 = ~w8148 & w18548;
assign w13153 = ~w126 & ~w12303;
assign w13154 = w13198 & ~w6054;
assign w13155 = ~w16798 & ~w19078;
assign w13156 = ~w14785 & ~w15839;
assign w13157 = ~w15265 & w1607;
assign w13158 = ~w569 & ~w2947;
assign w13159 = w10004 & ~w8661;
assign w13160 = ~w11168 & w18303;
assign w13161 = (~w11710 & ~w2348) | (~w11710 & w4095) | (~w2348 & w4095);
assign w13162 = ~w15701 & w11319;
assign w13163 = ~w2941 & ~w13042;
assign w13164 = a_7 & a_38;
assign w13165 = w696 & w6546;
assign w13166 = a_33 & a_42;
assign w13167 = ~w18430 & ~w15184;
assign w13168 = a_10 & a_24;
assign w13169 = a_32 & a_62;
assign w13170 = ~w5588 & ~w12674;
assign w13171 = ~w3708 & ~w14245;
assign w13172 = ~w8998 & w13977;
assign w13173 = ~w7377 & ~w12213;
assign w13174 = ~w7919 & ~w6206;
assign w13175 = (~w7768 & w16526) | (~w7768 & w9953) | (w16526 & w9953);
assign w13176 = w8350 & w9199;
assign w13177 = ~w11222 & ~w18738;
assign w13178 = ~w11352 & ~w15886;
assign w13179 = ~w13100 & w4129;
assign w13180 = w6111 & ~w19049;
assign w13181 = ~w6729 & ~w13250;
assign w13182 = ~w4758 & ~w5015;
assign w13183 = w15514 & w17493;
assign w13184 = w12229 & w157;
assign w13185 = (~w10273 & ~w53) | (~w10273 & w2147) | (~w53 & w2147);
assign w13186 = ~w7070 & w2663;
assign w13187 = ~w5680 & w4604;
assign w13188 = w11103 & ~w2312;
assign w13189 = w11413 & ~w18444;
assign w13190 = ~w5034 & ~w9054;
assign w13191 = w8264 & ~w1750;
assign w13192 = ~w75 & ~w3561;
assign w13193 = ~w12803 & ~w13109;
assign w13194 = ~w937 & ~w6404;
assign w13195 = ~w5163 & ~w10759;
assign w13196 = ~w6555 & ~w5049;
assign w13197 = ~w16326 & ~w6312;
assign w13198 = a_10 & w18633;
assign w13199 = ~w15827 & ~w7888;
assign w13200 = ~w11541 & ~w4293;
assign w13201 = ~w10240 & ~w18524;
assign w13202 = a_2 & a_50;
assign w13203 = ~w11043 & ~w10148;
assign w13204 = ~w8953 & ~w7319;
assign w13205 = w14751 & w6965;
assign w13206 = ~w16292 & ~w16434;
assign w13207 = a_15 & a_56;
assign w13208 = ~w9064 & ~w8040;
assign w13209 = w18327 & ~w6565;
assign w13210 = ~w11607 & ~w7064;
assign w13211 = ~w17986 & ~w15280;
assign w13212 = ~w11943 & w41;
assign w13213 = a_4 & a_20;
assign w13214 = ~w11752 & ~w6176;
assign w13215 = ~w14729 & ~w13146;
assign w13216 = w2577 & ~w990;
assign w13217 = ~w2980 & ~w2754;
assign w13218 = ~w5219 & ~w1038;
assign w13219 = a_8 & a_35;
assign w13220 = ~w16155 & ~w2508;
assign w13221 = a_1 & a_2;
assign w13222 = ~w15824 & ~w3282;
assign w13223 = a_1 & a_31;
assign w13224 = a_14 & a_41;
assign w13225 = ~w12990 & ~w16179;
assign w13226 = ~w17877 & ~w15687;
assign w13227 = a_9 & a_39;
assign w13228 = w11754 & ~w10253;
assign w13229 = ~w14827 & w9923;
assign w13230 = w2495 & ~w16960;
assign w13231 = ~w15797 & ~w11181;
assign w13232 = ~w12991 & ~w6245;
assign w13233 = ~w4091 & ~w13656;
assign w13234 = ~w11374 & w10123;
assign w13235 = ~w17655 & ~w14575;
assign w13236 = w7475 & w18105;
assign w13237 = ~w1302 & ~w2479;
assign w13238 = w7465 & ~w15865;
assign w13239 = w2319 & w6705;
assign w13240 = w10683 & w16350;
assign w13241 = ~w2496 & ~w1991;
assign w13242 = ~w4798 & ~w10105;
assign w13243 = w5365 & ~w7829;
assign w13244 = (~w963 & w1482) | (~w963 & ~w17701) | (w1482 & ~w17701);
assign w13245 = w14822 & ~w17509;
assign w13246 = ~w11833 & ~w5473;
assign w13247 = w576 & w304;
assign w13248 = ~w9388 & ~w2864;
assign w13249 = ~w18148 & ~w7245;
assign w13250 = ~w15175 & ~w17146;
assign w13251 = ~w10905 & ~w1856;
assign w13252 = a_55 & a_60;
assign w13253 = ~w8011 & ~w2787;
assign w13254 = w5632 & w5969;
assign w13255 = w8252 & w12891;
assign w13256 = w13801 & w6938;
assign w13257 = ~w4389 & w8774;
assign w13258 = ~w13859 & ~w5294;
assign w13259 = ~w15260 & ~w2036;
assign w13260 = w11982 & ~w1500;
assign w13261 = ~w14154 & ~w38;
assign w13262 = w18185 & ~w2879;
assign w13263 = w11826 & w14504;
assign w13264 = ~a_13 & w17557;
assign w13265 = w533 & w6592;
assign w13266 = a_11 & a_51;
assign w13267 = ~w4414 & ~w13188;
assign w13268 = a_46 & a_48;
assign w13269 = a_8 & a_13;
assign w13270 = ~w2727 & ~w15148;
assign w13271 = a_1 & a_49;
assign w13272 = ~w7237 & ~w11377;
assign w13273 = a_20 & a_36;
assign w13274 = ~w6177 & w18425;
assign w13275 = ~w8746 & ~w19139;
assign w13276 = w6057 & ~w8613;
assign w13277 = ~w6849 & w15784;
assign w13278 = w11278 & w5457;
assign w13279 = ~w19087 & ~w3778;
assign w13280 = w16493 & w19182;
assign w13281 = ~w8002 & ~w6512;
assign w13282 = ~w6315 & ~w6617;
assign w13283 = (w885 & w7034) | (w885 & w2650) | (w7034 & w2650);
assign w13284 = a_18 & a_54;
assign w13285 = w3932 & ~w7341;
assign w13286 = ~w985 & w2218;
assign w13287 = ~a_54 & a_55;
assign w13288 = ~w12904 & w15397;
assign w13289 = ~w2631 & ~w7542;
assign w13290 = a_31 & a_62;
assign w13291 = ~w12307 & ~w15709;
assign w13292 = ~w4778 & ~w8325;
assign w13293 = ~w5368 & ~w1521;
assign w13294 = ~w13076 & ~w9949;
assign w13295 = ~w8411 & ~w7554;
assign w13296 = ~w18150 & w8569;
assign w13297 = w17268 & ~w18038;
assign w13298 = ~w12618 & ~w8076;
assign w13299 = ~w16340 & ~w7223;
assign w13300 = ~w19143 & ~w17001;
assign w13301 = (~w27 & w593) | (~w27 & w12986) | (w593 & w12986);
assign w13302 = ~w12412 & ~w7403;
assign w13303 = a_5 & a_43;
assign w13304 = w18847 & w795;
assign w13305 = ~w16769 & w12422;
assign w13306 = ~w14633 & ~w1821;
assign w13307 = ~w4478 & ~w11854;
assign w13308 = w18485 & ~w8915;
assign w13309 = ~w17482 & ~w18735;
assign w13310 = ~w10943 & ~w4695;
assign w13311 = a_19 & a_57;
assign w13312 = ~w11372 & ~w10916;
assign w13313 = ~w7256 & ~w16571;
assign w13314 = ~w16749 & ~w6944;
assign w13315 = w18132 & w14828;
assign w13316 = w11492 & ~w11140;
assign w13317 = ~w10672 & ~w16898;
assign w13318 = w17956 & ~w4139;
assign w13319 = w15358 & w8627;
assign w13320 = a_1 & a_47;
assign w13321 = ~w9176 & ~w435;
assign w13322 = w14426 & w4639;
assign w13323 = ~w16399 & w14425;
assign w13324 = a_0 & a_23;
assign w13325 = ~w8201 & ~w1033;
assign w13326 = a_48 & a_59;
assign w13327 = ~w3235 & w375;
assign w13328 = ~w4645 & ~w8147;
assign w13329 = ~w17421 & w17757;
assign w13330 = w12894 & w12133;
assign w13331 = w12726 & ~w218;
assign w13332 = ~w3702 & ~w2360;
assign w13333 = a_10 & a_61;
assign w13334 = w7595 & w16878;
assign w13335 = ~w11119 & ~w4254;
assign w13336 = ~w4633 & ~w3126;
assign w13337 = w17980 & ~w5221;
assign w13338 = a_21 & a_28;
assign w13339 = ~w4033 & ~w4714;
assign w13340 = ~w4265 & w5767;
assign w13341 = (w15988 & w6740) | (w15988 & w3061) | (w6740 & w3061);
assign w13342 = ~w2042 & w4623;
assign w13343 = a_38 & a_52;
assign w13344 = ~w7560 & w8272;
assign w13345 = ~w9383 & ~w5364;
assign w13346 = a_9 & a_46;
assign w13347 = a_4 & a_35;
assign w13348 = w10838 & w18845;
assign w13349 = ~w5274 & ~w8470;
assign w13350 = a_26 & a_32;
assign w13351 = w11003 & ~w11231;
assign w13352 = ~w9882 & ~w1930;
assign w13353 = ~w17168 & ~w14272;
assign w13354 = (~w1525 & ~w321) | (~w1525 & w17756) | (~w321 & w17756);
assign w13355 = ~w17145 & ~w1623;
assign w13356 = w11944 & w13798;
assign w13357 = (w15306 & w13082) | (w15306 & w18265) | (w13082 & w18265);
assign w13358 = w15145 & w14553;
assign w13359 = w17379 & ~w3287;
assign w13360 = ~w7292 & ~w18231;
assign w13361 = ~w17800 & ~w12953;
assign w13362 = w18134 & w14166;
assign w13363 = w17115 & ~w2001;
assign w13364 = ~w15801 & ~w11872;
assign w13365 = ~w11591 & ~w12774;
assign w13366 = ~w17060 & w4506;
assign w13367 = ~w10786 & w767;
assign w13368 = ~w8735 & ~w12999;
assign w13369 = ~w4610 & ~w8359;
assign w13370 = ~w4840 & ~w8709;
assign w13371 = ~w5522 & ~w6352;
assign w13372 = w17218 & ~w11472;
assign w13373 = (~w9436 & ~w2423) | (~w9436 & w7547) | (~w2423 & w7547);
assign w13374 = w14547 & w15368;
assign w13375 = (w6279 & w2769) | (w6279 & w1197) | (w2769 & w1197);
assign w13376 = ~w1894 & ~w15618;
assign w13377 = (w10181 & ~w9201) | (w10181 & w12166) | (~w9201 & w12166);
assign w13378 = ~w5337 & w1869;
assign w13379 = (~w5999 & ~w3778) | (~w5999 & w3716) | (~w3778 & w3716);
assign w13380 = ~w15613 & ~w12338;
assign w13381 = w1962 & w11712;
assign w13382 = ~w1428 & ~w6240;
assign w13383 = ~w18437 & w14332;
assign w13384 = ~w16400 & ~w4401;
assign w13385 = ~w15394 & ~w6463;
assign w13386 = ~w1353 & w16614;
assign w13387 = w1298 & w1989;
assign w13388 = w4537 & ~w4715;
assign w13389 = ~w1954 & ~w6340;
assign w13390 = a_7 & a_35;
assign w13391 = ~w6951 & w15637;
assign w13392 = ~w8042 & ~w726;
assign w13393 = ~w3658 & w1382;
assign w13394 = ~w8439 & ~w10401;
assign w13395 = ~w2458 & ~w1171;
assign w13396 = ~w8688 & ~w15385;
assign w13397 = ~w5499 & w17846;
assign w13398 = ~w14510 & ~w18191;
assign w13399 = a_18 & a_62;
assign w13400 = ~w8896 & ~w6178;
assign w13401 = ~w4680 & ~w18142;
assign w13402 = w11528 & w8030;
assign w13403 = w8943 & ~w9118;
assign w13404 = (~w613 & ~w10577) | (~w613 & w14838) | (~w10577 & w14838);
assign w13405 = ~w10886 & ~w17403;
assign w13406 = ~w5944 & w15321;
assign w13407 = w18525 & w11056;
assign w13408 = a_8 & a_16;
assign w13409 = w12253 & ~w16082;
assign w13410 = w5349 & ~w13185;
assign w13411 = ~w12156 & w3532;
assign w13412 = ~w12123 & ~w6768;
assign w13413 = a_37 & a_53;
assign w13414 = ~w1711 & ~w10390;
assign w13415 = ~w15543 & w4156;
assign w13416 = w8870 & w5498;
assign w13417 = (~w10929 & ~w16016) | (~w10929 & w9967) | (~w16016 & w9967);
assign w13418 = w8718 & ~w15101;
assign w13419 = ~w17930 & ~w3558;
assign w13420 = (w5904 & ~w4766) | (w5904 & w15118) | (~w4766 & w15118);
assign w13421 = ~w2052 & ~w3953;
assign w13422 = ~w12297 & w8214;
assign w13423 = (~w12254 & w8854) | (~w12254 & w12920) | (w8854 & w12920);
assign w13424 = ~w6954 & ~w5922;
assign w13425 = w2182 & w2401;
assign w13426 = w13326 & ~w14040;
assign w13427 = ~w1965 & ~w10642;
assign w13428 = ~w3340 & ~w702;
assign w13429 = w15423 & w2543;
assign w13430 = ~w1635 & ~w6051;
assign w13431 = w6285 & ~w18969;
assign w13432 = a_44 & a_50;
assign w13433 = ~w6268 & ~w2488;
assign w13434 = ~w7696 & ~w3838;
assign w13435 = ~w7090 & w14915;
assign w13436 = ~w548 & ~w3374;
assign w13437 = ~w3800 & w2389;
assign w13438 = a_21 & a_61;
assign w13439 = ~w12027 & ~w10809;
assign w13440 = w10 & ~w11484;
assign w13441 = ~w10015 & ~w16043;
assign w13442 = w16951 & ~w18573;
assign w13443 = ~w14106 & w18556;
assign w13444 = w17946 & ~w17242;
assign w13445 = ~a_40 & ~w14868;
assign w13446 = w17858 & w15402;
assign w13447 = w15976 & ~w9451;
assign w13448 = ~w11323 & ~w10631;
assign w13449 = w15975 & ~w14711;
assign w13450 = ~w896 & ~w14739;
assign w13451 = w8761 & ~w13667;
assign w13452 = ~w15951 & ~w16171;
assign w13453 = ~w10734 & ~w10270;
assign w13454 = w16529 & ~w9179;
assign w13455 = ~w15548 & ~w18420;
assign w13456 = ~w8346 & ~w8415;
assign w13457 = ~w17502 & w7664;
assign w13458 = w17126 & w13697;
assign w13459 = ~w14160 & ~w13013;
assign w13460 = ~w6267 & w6236;
assign w13461 = ~w11567 & ~w3505;
assign w13462 = ~w19 & ~w16301;
assign w13463 = a_19 & a_63;
assign w13464 = ~w10466 & w17358;
assign w13465 = ~w18572 & ~w11359;
assign w13466 = a_39 & a_46;
assign w13467 = ~w9433 & ~w15683;
assign w13468 = w14006 & w8285;
assign w13469 = w6571 & ~w948;
assign w13470 = ~w17936 & ~w6854;
assign w13471 = w14359 & ~w15092;
assign w13472 = a_52 & a_60;
assign w13473 = ~w7582 & ~w13846;
assign w13474 = w6923 & w5642;
assign w13475 = ~w9437 & ~w16978;
assign w13476 = ~w18436 & ~w495;
assign w13477 = w9597 & ~w14769;
assign w13478 = a_11 & a_44;
assign w13479 = w1320 & w9799;
assign w13480 = a_21 & a_29;
assign w13481 = (~w7102 & w14021) | (~w7102 & w7876) | (w14021 & w7876);
assign w13482 = ~w10531 & ~w13184;
assign w13483 = (~w12299 & ~w15504) | (~w12299 & w2332) | (~w15504 & w2332);
assign w13484 = ~w2327 & ~w13550;
assign w13485 = ~w11475 & ~w14541;
assign w13486 = ~w14557 & ~w13084;
assign w13487 = a_41 & a_50;
assign w13488 = w3117 & ~w10020;
assign w13489 = a_14 & a_63;
assign w13490 = a_2 & a_48;
assign w13491 = ~w16600 & ~w4699;
assign w13492 = ~w9008 & w1598;
assign w13493 = ~w6225 & ~w18106;
assign w13494 = w94 & w169;
assign w13495 = ~w3228 & ~w3654;
assign w13496 = ~w6146 & w197;
assign w13497 = (~w10790 & w10770) | (~w10790 & w758) | (w10770 & w758);
assign w13498 = w16483 & ~w497;
assign w13499 = w8239 & w9914;
assign w13500 = ~w12750 & ~w1179;
assign w13501 = ~w5100 & ~w11796;
assign w13502 = w13140 & w488;
assign w13503 = ~w557 & w4489;
assign w13504 = a_18 & a_36;
assign w13505 = a_30 & a_31;
assign w13506 = w14982 & ~w186;
assign w13507 = w2637 & ~w4640;
assign w13508 = ~w4698 & ~w4817;
assign w13509 = (w7150 & ~w7586) | (w7150 & w7354) | (~w7586 & w7354);
assign w13510 = ~w9324 & ~w18384;
assign w13511 = ~w15384 & w2291;
assign w13512 = a_29 & a_63;
assign w13513 = ~w18069 & ~w3647;
assign w13514 = ~w7870 & ~w12128;
assign w13515 = ~w10243 & ~w933;
assign w13516 = ~w5194 & ~w13083;
assign w13517 = ~w12056 & ~w18044;
assign w13518 = w8551 & w7198;
assign w13519 = w5381 & w1026;
assign w13520 = ~w16626 & w6911;
assign w13521 = w8500 & w2685;
assign w13522 = a_2 & a_49;
assign w13523 = ~w2667 & ~w10161;
assign w13524 = ~w5692 & ~w6549;
assign w13525 = ~w6248 & ~w2501;
assign w13526 = ~w11344 & ~w7786;
assign w13527 = ~w2242 & w13829;
assign w13528 = ~w11562 & ~w18880;
assign w13529 = w697 & ~w11328;
assign w13530 = ~w14613 & ~w10021;
assign w13531 = ~w17052 & w10450;
assign w13532 = ~w5334 & ~w3617;
assign w13533 = (~w4517 & ~w6368) | (~w4517 & w1409) | (~w6368 & w1409);
assign w13534 = (~w14247 & ~w7976) | (~w14247 & w4175) | (~w7976 & w4175);
assign w13535 = w5176 & w17551;
assign w13536 = ~w5123 & ~w12339;
assign w13537 = ~w13432 & ~w5247;
assign w13538 = w6109 & w14176;
assign w13539 = w2876 & ~w18;
assign w13540 = ~w2714 & ~w9659;
assign w13541 = w17097 & w4373;
assign w13542 = w15149 & ~w4785;
assign w13543 = w1993 & w6068;
assign w13544 = ~w16976 & ~w16985;
assign w13545 = a_13 & a_21;
assign w13546 = w15274 & w15506;
assign w13547 = w16564 & ~w17947;
assign w13548 = w10926 & w2978;
assign w13549 = ~w10900 & ~w4239;
assign w13550 = ~w16741 & w10650;
assign w13551 = ~w2293 & ~w11524;
assign w13552 = ~w10853 & ~w7331;
assign w13553 = a_11 & a_35;
assign w13554 = w4367 & w19183;
assign w13555 = ~w5947 & w3856;
assign w13556 = ~w9315 & ~w9756;
assign w13557 = (~w411 & ~w1993) | (~w411 & w15892) | (~w1993 & w15892);
assign w13558 = (w152 & w3179) | (w152 & w19030) | (w3179 & w19030);
assign w13559 = (~w5035 & ~w14442) | (~w5035 & w163) | (~w14442 & w163);
assign w13560 = ~w4950 & w4245;
assign w13561 = ~w7630 & w7761;
assign w13562 = w3507 & w7027;
assign w13563 = ~w13168 & ~w18110;
assign w13564 = w4030 & ~w4875;
assign w13565 = (w13280 & w16428) | (w13280 & w15856) | (w16428 & w15856);
assign w13566 = ~w17538 & ~w8891;
assign w13567 = ~w7106 & ~w14197;
assign w13568 = ~w11674 & w4295;
assign w13569 = ~w6244 & ~w18050;
assign w13570 = ~w13281 & w2446;
assign w13571 = ~w9415 & ~w17125;
assign w13572 = ~w13164 & ~w17824;
assign w13573 = w6453 & ~w3909;
assign w13574 = (w17376 & ~w7299) | (w17376 & w122) | (~w7299 & w122);
assign w13575 = ~w14721 & ~w3700;
assign w13576 = ~w4800 & ~w18517;
assign w13577 = ~w17098 & ~w4602;
assign w13578 = w10206 & w16831;
assign w13579 = (~w17604 & w11644) | (~w17604 & w1618) | (w11644 & w1618);
assign w13580 = ~w5968 & ~w16875;
assign w13581 = a_9 & a_28;
assign w13582 = w15555 & w1700;
assign w13583 = ~w6853 & w9869;
assign w13584 = ~w7773 & w66;
assign w13585 = a_36 & a_60;
assign w13586 = ~w13116 & ~w14778;
assign w13587 = a_4 & a_54;
assign w13588 = ~w4137 & w17236;
assign w13589 = a_32 & a_42;
assign w13590 = ~w17581 & ~w12204;
assign w13591 = ~w2571 & ~w12276;
assign w13592 = w2921 & ~w6454;
assign w13593 = ~w5557 & ~w8132;
assign w13594 = w17955 & w2547;
assign w13595 = ~w6396 & w1553;
assign w13596 = ~w11317 & ~w3687;
assign w13597 = ~w237 & ~w17905;
assign w13598 = ~w11258 & ~w6606;
assign w13599 = ~w9458 & ~w805;
assign w13600 = w10121 & w1967;
assign w13601 = a_39 & a_59;
assign w13602 = w15686 & ~w12375;
assign w13603 = ~w14460 & ~w9776;
assign w13604 = ~w9135 & ~w18345;
assign w13605 = ~w7277 & ~w5748;
assign w13606 = w6383 & ~w3769;
assign w13607 = ~w11332 & ~w15601;
assign w13608 = (w15988 & w7023) | (w15988 & w7397) | (w7023 & w7397);
assign w13609 = ~w7177 & ~w13938;
assign w13610 = ~w2883 & ~w6978;
assign w13611 = ~w12051 & ~w2275;
assign w13612 = ~w8584 & w2806;
assign w13613 = ~w17659 & ~w13822;
assign w13614 = ~w2431 & ~w17159;
assign w13615 = ~w18700 & ~w16539;
assign w13616 = w7638 & ~w9468;
assign w13617 = ~w5483 & ~w15533;
assign w13618 = ~w12439 & ~w5131;
assign w13619 = ~w2915 & ~w17726;
assign w13620 = ~w11154 & ~w8082;
assign w13621 = ~w3160 & ~w16295;
assign w13622 = ~w14783 & ~w18677;
assign w13623 = w12038 & w1589;
assign w13624 = (w14792 & w16190) | (w14792 & w12530) | (w16190 & w12530);
assign w13625 = ~w3511 & ~w748;
assign w13626 = ~w5538 & ~w17144;
assign w13627 = w10082 & w4207;
assign w13628 = w13213 & w18098;
assign w13629 = ~w13771 & w5201;
assign w13630 = ~w11464 & ~w15525;
assign w13631 = w19134 & ~w8951;
assign w13632 = ~w261 & ~w18808;
assign w13633 = ~w16148 & ~w17158;
assign w13634 = ~w4894 & ~w115;
assign w13635 = ~w15095 & ~w6963;
assign w13636 = ~w1889 & ~w6544;
assign w13637 = ~w7941 & ~w8300;
assign w13638 = w16506 & w9887;
assign w13639 = w17581 & ~w9934;
assign w13640 = w15655 & w14266;
assign w13641 = w14786 & ~w8999;
assign w13642 = w18553 & ~w15772;
assign w13643 = ~w12641 & ~w7574;
assign w13644 = ~w5604 & ~w14094;
assign w13645 = ~w759 & w9888;
assign w13646 = ~w15609 & ~w15679;
assign w13647 = w11652 & w18462;
assign w13648 = ~w862 & ~w16446;
assign w13649 = ~w6901 & w6236;
assign w13650 = ~w10130 & ~w6175;
assign w13651 = ~w17554 & ~w5446;
assign w13652 = ~w17740 & ~w17020;
assign w13653 = a_1 & a_21;
assign w13654 = ~w6126 & ~w7364;
assign w13655 = a_5 & a_40;
assign w13656 = (w7596 & w2769) | (w7596 & w14766) | (w2769 & w14766);
assign w13657 = ~w14568 & ~w13277;
assign w13658 = ~w10770 & w7873;
assign w13659 = ~w374 & ~w3782;
assign w13660 = ~w10625 & ~w16411;
assign w13661 = ~w3772 & ~w5309;
assign w13662 = w6831 & ~w11396;
assign w13663 = w1320 & w3910;
assign w13664 = ~w15528 & ~w4685;
assign w13665 = ~w464 & ~w16682;
assign w13666 = ~w4586 & ~w5271;
assign w13667 = ~w13544 & ~w13368;
assign w13668 = ~w3082 & w15200;
assign w13669 = a_31 & a_47;
assign w13670 = ~w5782 & ~w6936;
assign w13671 = w2660 & ~w221;
assign w13672 = ~w6165 & w5496;
assign w13673 = ~w6381 & ~w13197;
assign w13674 = a_2 & a_22;
assign w13675 = w5435 & w6378;
assign w13676 = w562 & w6541;
assign w13677 = ~w2905 & w10815;
assign w13678 = w6360 & w8719;
assign w13679 = (w9208 & w14382) | (w9208 & w4059) | (w14382 & w4059);
assign w13680 = ~w7529 & ~w5757;
assign w13681 = ~w141 & ~w10727;
assign w13682 = ~w10030 & w14230;
assign w13683 = ~w17811 & w1420;
assign w13684 = a_26 & a_62;
assign w13685 = w14982 & ~w8164;
assign w13686 = ~w18383 & ~w7610;
assign w13687 = ~w17453 & ~w14962;
assign w13688 = ~w18437 & w9957;
assign w13689 = a_20 & a_25;
assign w13690 = ~w6760 & ~w4282;
assign w13691 = ~w3650 & ~w6508;
assign w13692 = w5022 & w1497;
assign w13693 = ~w10758 & ~w16339;
assign w13694 = w17359 & ~w10496;
assign w13695 = ~w993 & ~w16677;
assign w13696 = w3236 & ~w3556;
assign w13697 = ~w14222 & ~w15540;
assign w13698 = w16054 & w13910;
assign w13699 = a_13 & a_54;
assign w13700 = ~w18427 & ~w10636;
assign w13701 = ~w6583 & ~w7482;
assign w13702 = ~w2083 & ~w16233;
assign w13703 = ~w11309 & ~w8353;
assign w13704 = (w7102 & w14858) | (w7102 & w16561) | (w14858 & w16561);
assign w13705 = ~w13903 & ~w1639;
assign w13706 = w11748 & ~w17101;
assign w13707 = w4792 & w11681;
assign w13708 = w14367 & ~w1787;
assign w13709 = w4585 & w3431;
assign w13710 = w11533 & ~w16103;
assign w13711 = ~w10817 & ~w15438;
assign w13712 = w7630 & ~w7761;
assign w13713 = a_26 & a_49;
assign w13714 = a_6 & a_27;
assign w13715 = w17246 & w3867;
assign w13716 = w10363 & ~w2043;
assign w13717 = w8736 & ~w6471;
assign w13718 = a_20 & a_37;
assign w13719 = w4894 & w115;
assign w13720 = w11208 & w14441;
assign w13721 = a_2 & a_36;
assign w13722 = ~w8893 & ~w11677;
assign w13723 = ~w6130 & ~w11520;
assign w13724 = ~w10619 & ~w8149;
assign w13725 = w517 & ~w1579;
assign w13726 = w16546 & ~w18145;
assign w13727 = w6189 & w5030;
assign w13728 = w1316 & ~w7087;
assign w13729 = w3699 & ~w12064;
assign w13730 = a_8 & a_44;
assign w13731 = ~w8479 & w13194;
assign w13732 = a_27 & a_63;
assign w13733 = ~w19005 & w7969;
assign w13734 = ~w2022 & ~w6816;
assign w13735 = a_15 & a_29;
assign w13736 = a_19 & a_48;
assign w13737 = ~w969 & ~w15203;
assign w13738 = w960 & ~w16521;
assign w13739 = ~w7425 & w498;
assign w13740 = w5151 & ~w1045;
assign w13741 = ~w535 & w11037;
assign w13742 = ~w13021 & w17368;
assign w13743 = w1016 & w3194;
assign w13744 = ~w18762 & ~w2148;
assign w13745 = ~w5830 & ~w2854;
assign w13746 = w3121 & ~w15509;
assign w13747 = ~w16296 & ~w13824;
assign w13748 = ~w17449 & ~w16325;
assign w13749 = ~w10446 & ~w5717;
assign w13750 = w6741 & w4629;
assign w13751 = w4101 & ~w13776;
assign w13752 = (~w14630 & ~w7595) | (~w14630 & w997) | (~w7595 & w997);
assign w13753 = ~w12975 & ~w8124;
assign w13754 = w4053 & ~w17961;
assign w13755 = w12239 & ~w1094;
assign w13756 = ~w12262 & ~w10203;
assign w13757 = w4389 & ~w8774;
assign w13758 = (~w7102 & w18195) | (~w7102 & w16021) | (w18195 & w16021);
assign w13759 = ~w2235 & w17306;
assign w13760 = ~w15263 & ~w2640;
assign w13761 = a_7 & a_18;
assign w13762 = ~w3161 & w1152;
assign w13763 = ~w8941 & ~w12065;
assign w13764 = w4408 & w6063;
assign w13765 = a_4 & a_12;
assign w13766 = ~w12606 & w2037;
assign w13767 = ~w7190 & ~w3008;
assign w13768 = ~w83 & w12118;
assign w13769 = ~w11166 & w5886;
assign w13770 = ~w17193 & ~w13062;
assign w13771 = a_10 & a_15;
assign w13772 = ~w18998 & ~w7290;
assign w13773 = ~w10697 & ~w17294;
assign w13774 = w15744 & ~w10595;
assign w13775 = (w804 & ~w13082) | (w804 & w9628) | (~w13082 & w9628);
assign w13776 = ~w16364 & ~w1832;
assign w13777 = ~w12759 & ~w17044;
assign w13778 = w10338 & w2188;
assign w13779 = w18838 & ~w7259;
assign w13780 = ~w12374 & ~w6591;
assign w13781 = w11965 & ~w10958;
assign w13782 = w14985 & w11540;
assign w13783 = ~w18908 & ~w761;
assign w13784 = w6431 & ~w11603;
assign w13785 = ~w9844 & ~w13366;
assign w13786 = ~w7701 & w1225;
assign w13787 = ~w19072 & w17632;
assign w13788 = ~w9561 & ~w15339;
assign w13789 = ~w1752 & ~w1072;
assign w13790 = a_28 & a_46;
assign w13791 = ~w2243 & ~w7777;
assign w13792 = a_0 & a_40;
assign w13793 = a_22 & a_54;
assign w13794 = (~w7504 & ~w8786) | (~w7504 & w17594) | (~w8786 & w17594);
assign w13795 = ~w9243 & ~w15804;
assign w13796 = ~w17516 & ~w18436;
assign w13797 = ~w2906 & ~w14518;
assign w13798 = a_1 & a_17;
assign w13799 = ~w18027 & w2000;
assign w13800 = ~w15168 & ~w15682;
assign w13801 = ~w8695 & ~w3644;
assign w13802 = ~w18443 & ~w971;
assign w13803 = ~w11902 & ~w8139;
assign w13804 = ~w17930 & ~w17304;
assign w13805 = a_28 & a_41;
assign w13806 = (~w3856 & w11583) | (~w3856 & w10453) | (w11583 & w10453);
assign w13807 = a_26 & a_27;
assign w13808 = ~w7590 & w14734;
assign w13809 = ~w1212 & ~w8692;
assign w13810 = ~w1962 & w3238;
assign w13811 = ~w17949 & ~w15842;
assign w13812 = w18936 & w6479;
assign w13813 = a_12 & a_40;
assign w13814 = ~w11506 & w4513;
assign w13815 = ~w17850 & ~w10482;
assign w13816 = a_1 & a_52;
assign w13817 = ~w16220 & ~w14829;
assign w13818 = ~w2432 & ~w1310;
assign w13819 = ~w17171 & ~w8186;
assign w13820 = w10878 & w14764;
assign w13821 = ~w3612 & ~w1647;
assign w13822 = ~w13466 & w9563;
assign w13823 = ~w13326 & ~w11608;
assign w13824 = ~w1283 & w10513;
assign w13825 = a_49 & a_53;
assign w13826 = w508 & ~w17308;
assign w13827 = a_0 & a_45;
assign w13828 = ~w7652 & ~w7955;
assign w13829 = ~w15476 & ~w6785;
assign w13830 = ~w4375 & ~w17053;
assign w13831 = ~w5425 & w6296;
assign w13832 = ~w18285 & ~w342;
assign w13833 = ~w12879 & w4881;
assign w13834 = ~w7269 & ~w5709;
assign w13835 = ~w18675 & ~w2044;
assign w13836 = w11194 & ~w6971;
assign w13837 = (w1007 & w2769) | (w1007 & w516) | (w2769 & w516);
assign w13838 = ~w17999 & w11595;
assign w13839 = ~w3260 & ~w9797;
assign w13840 = ~w18510 & ~w4109;
assign w13841 = ~w1530 & ~w5674;
assign w13842 = ~w7501 & ~w12895;
assign w13843 = w4886 & w15089;
assign w13844 = a_12 & a_36;
assign w13845 = ~w10412 & ~w16872;
assign w13846 = ~w9873 & w17626;
assign w13847 = w12163 & w2368;
assign w13848 = (~w13179 & ~w17571) | (~w13179 & w3253) | (~w17571 & w3253);
assign w13849 = a_11 & a_50;
assign w13850 = ~w2843 & ~w11694;
assign w13851 = a_17 & a_58;
assign w13852 = ~w13379 & w7557;
assign w13853 = ~w9023 & ~w798;
assign w13854 = a_1 & a_60;
assign w13855 = ~w13442 & ~w1281;
assign w13856 = ~w10865 & w15341;
assign w13857 = ~w6525 & ~w10975;
assign w13858 = w2836 & ~w127;
assign w13859 = ~w3686 & ~w18426;
assign w13860 = ~w9494 & ~w14901;
assign w13861 = a_10 & a_63;
assign w13862 = w16807 & ~w16234;
assign w13863 = ~w9859 & w12882;
assign w13864 = a_31 & a_38;
assign w13865 = ~w11112 & w4274;
assign w13866 = ~w6424 & ~w18638;
assign w13867 = w5412 & w16806;
assign w13868 = ~w4418 & ~w13716;
assign w13869 = a_23 & a_35;
assign w13870 = ~w2942 & ~w3639;
assign w13871 = ~w3154 & ~w11584;
assign w13872 = (~w12281 & w1050) | (~w12281 & w18017) | (w1050 & w18017);
assign w13873 = a_39 & a_44;
assign w13874 = ~w13114 & ~w1835;
assign w13875 = w17418 & ~w14957;
assign w13876 = ~w13011 & ~w8631;
assign w13877 = w8737 & ~w8454;
assign w13878 = ~w7411 & ~w9660;
assign w13879 = ~w8609 & ~w3685;
assign w13880 = ~w10228 & w16977;
assign w13881 = ~w18179 & ~w7414;
assign w13882 = w11692 & w2381;
assign w13883 = w370 & ~w12057;
assign w13884 = ~w750 & ~w14037;
assign w13885 = w10350 & w10933;
assign w13886 = ~w5912 & ~w8253;
assign w13887 = (~w4884 & ~w10179) | (~w4884 & w6731) | (~w10179 & w6731);
assign w13888 = ~w1207 & ~w1188;
assign w13889 = ~w11339 & ~w18478;
assign w13890 = ~w10246 & ~w7458;
assign w13891 = ~w1191 & w16838;
assign w13892 = ~w13886 & ~w7422;
assign w13893 = ~w17475 & ~w10417;
assign w13894 = (~w9611 & w10337) | (~w9611 & w4178) | (w10337 & w4178);
assign w13895 = a_30 & a_55;
assign w13896 = ~w13418 & ~w1177;
assign w13897 = w2603 & ~w6193;
assign w13898 = (w10232 & w17132) | (w10232 & w16147) | (w17132 & w16147);
assign w13899 = ~w12238 & ~w11993;
assign w13900 = ~w18644 & w12261;
assign w13901 = ~w12098 & w1475;
assign w13902 = ~w563 & ~w18742;
assign w13903 = w11671 & w14908;
assign w13904 = w1050 | ~w12281;
assign w13905 = (~w9472 & ~w17185) | (~w9472 & w4127) | (~w17185 & w4127);
assign w13906 = ~w9593 & w10086;
assign w13907 = ~w16091 & ~w7203;
assign w13908 = ~w1035 & ~w12063;
assign w13909 = a_22 & a_45;
assign w13910 = ~w11188 & ~w16519;
assign w13911 = ~w11112 & ~w1779;
assign w13912 = w17362 & ~w12450;
assign w13913 = ~w8866 & ~w854;
assign w13914 = ~w19141 & ~w1240;
assign w13915 = ~w7369 & w18314;
assign w13916 = w6338 & ~w13963;
assign w13917 = (w10464 & w11313) | (w10464 & w11535) | (w11313 & w11535);
assign w13918 = ~w13444 & ~w14142;
assign w13919 = a_0 & a_22;
assign w13920 = ~w6825 & ~w14655;
assign w13921 = ~w12420 & ~w496;
assign w13922 = ~w16557 & ~w15819;
assign w13923 = (w10445 & w10330) | (w10445 & w16305) | (w10330 & w16305);
assign w13924 = (~w18554 & ~w4228) | (~w18554 & w17382) | (~w4228 & w17382);
assign w13925 = ~w942 & w6691;
assign w13926 = a_19 & a_44;
assign w13927 = (~w5745 & ~w8987) | (~w5745 & w2497) | (~w8987 & w2497);
assign w13928 = ~w8406 & ~w1185;
assign w13929 = ~w6853 & w1394;
assign w13930 = ~w677 & ~w12120;
assign w13931 = a_30 & a_46;
assign w13932 = ~w11465 & ~w3313;
assign w13933 = ~w17280 & ~w10915;
assign w13934 = ~w6264 & ~w9249;
assign w13935 = (w12404 & w6087) | (w12404 & w5882) | (w6087 & w5882);
assign w13936 = ~w8520 & ~w11682;
assign w13937 = w17622 & w1511;
assign w13938 = ~w9286 & w35;
assign w13939 = w8763 & ~w10491;
assign w13940 = (~w10092 & ~w18067) | (~w10092 & w17883) | (~w18067 & w17883);
assign w13941 = ~w18316 & w15961;
assign w13942 = ~w4208 & w4458;
assign w13943 = ~w18692 & ~w15857;
assign w13944 = w10922 & w12407;
assign w13945 = w7825 & w2352;
assign w13946 = w13605 & ~w7118;
assign w13947 = ~w7952 & ~w4755;
assign w13948 = ~w3259 & w93;
assign w13949 = ~w3786 & ~w14717;
assign w13950 = (w11243 & w13082) | (w11243 & w2784) | (w13082 & w2784);
assign w13951 = w17943 & w15932;
assign w13952 = w2837 & w5351;
assign w13953 = w394 & ~w18975;
assign w13954 = ~w4848 & ~w12478;
assign w13955 = w11736 & w10506;
assign w13956 = w279 & ~w3876;
assign w13957 = ~w1849 & ~w8656;
assign w13958 = a_10 & a_52;
assign w13959 = ~w17196 & ~w3692;
assign w13960 = w15443 & ~w10608;
assign w13961 = ~w4679 & ~w465;
assign w13962 = ~w11866 & w4789;
assign w13963 = ~w16625 & ~w4915;
assign w13964 = w5416 & w1949;
assign w13965 = ~w4083 & ~w2687;
assign w13966 = ~w13932 & ~w3163;
assign w13967 = w8039 & w14751;
assign w13968 = w9716 & ~w10235;
assign w13969 = (~w1953 & ~w15581) | (~w1953 & w9851) | (~w15581 & w9851);
assign w13970 = ~w8445 & ~w10886;
assign w13971 = (~w13060 & ~w7356) | (~w13060 & w11445) | (~w7356 & w11445);
assign w13972 = ~w11597 & w15652;
assign w13973 = a_3 & a_43;
assign w13974 = ~w7632 & ~w11384;
assign w13975 = w5697 & ~w14495;
assign w13976 = w3334 & ~w12856;
assign w13977 = ~w9187 & ~w2698;
assign w13978 = w4999 & ~w90;
assign w13979 = w4766 & ~w19035;
assign w13980 = ~w14171 & w2990;
assign w13981 = a_46 & a_63;
assign w13982 = ~w13300 & ~w16545;
assign w13983 = ~w8520 & ~w1334;
assign w13984 = ~w1633 & w3010;
assign w13985 = ~w963 & w1774;
assign w13986 = w18170 & w288;
assign w13987 = ~w2637 & w4640;
assign w13988 = w16792 & w3187;
assign w13989 = a_18 & a_42;
assign w13990 = ~w3381 & ~w12184;
assign w13991 = ~w9061 & ~w15390;
assign w13992 = ~w9753 & ~w7396;
assign w13993 = ~w15692 & w15612;
assign w13994 = ~w18205 & ~w12412;
assign w13995 = ~w3704 & ~w2823;
assign w13996 = w10650 & ~w10334;
assign w13997 = ~w2952 & ~w5265;
assign w13998 = a_3 & a_29;
assign w13999 = w14689 & w16489;
assign w14000 = w1208 & ~w10300;
assign w14001 = ~w8658 & ~w13520;
assign w14002 = w16836 & w9207;
assign w14003 = w2873 & w7226;
assign w14004 = w14699 & ~w12740;
assign w14005 = w8708 & w18634;
assign w14006 = ~w12199 & ~w9754;
assign w14007 = ~a_26 & ~w6141;
assign w14008 = (~w4062 & ~w8987) | (~w4062 & w5469) | (~w8987 & w5469);
assign w14009 = ~w11730 & ~w18700;
assign w14010 = ~w7591 & ~w8825;
assign w14011 = w9437 & w16978;
assign w14012 = a_37 & a_42;
assign w14013 = ~w17407 & ~w16019;
assign w14014 = ~w15557 & ~w10548;
assign w14015 = ~w1001 & ~w5390;
assign w14016 = ~w14000 & ~w4213;
assign w14017 = ~w7609 & ~w5998;
assign w14018 = ~w4298 & w12956;
assign w14019 = w10672 & w16898;
assign w14020 = ~w16153 & ~w18663;
assign w14021 = w8169 & ~w4766;
assign w14022 = ~w6002 & w4451;
assign w14023 = ~w18823 & w14937;
assign w14024 = (~w6886 & ~w1144) | (~w6886 & w133) | (~w1144 & w133);
assign w14025 = w811 & w9948;
assign w14026 = ~w10393 & ~w5182;
assign w14027 = ~w10044 & ~w13643;
assign w14028 = ~w16517 & ~w16502;
assign w14029 = w9567 & ~w5406;
assign w14030 = ~w16363 & ~w15703;
assign w14031 = ~w8840 & ~w9735;
assign w14032 = a_17 & a_40;
assign w14033 = ~w237 & ~w1372;
assign w14034 = a_14 & w14403;
assign w14035 = ~w6733 & ~w7386;
assign w14036 = w19130 & w13918;
assign w14037 = w12841 & w10384;
assign w14038 = w5682 & w5926;
assign w14039 = w4208 & ~w4458;
assign w14040 = ~w17351 & ~w11608;
assign w14041 = ~w10124 & ~w1205;
assign w14042 = w4662 & ~w3456;
assign w14043 = ~w17814 & w11037;
assign w14044 = ~w15472 & ~w1095;
assign w14045 = w14152 & ~w5405;
assign w14046 = ~w12446 & w6039;
assign w14047 = ~w8086 & ~w18976;
assign w14048 = ~w6756 & w13250;
assign w14049 = a_26 & a_40;
assign w14050 = a_46 & a_62;
assign w14051 = w9708 & w14949;
assign w14052 = ~w12777 & ~w11795;
assign w14053 = ~w12904 & ~w8639;
assign w14054 = ~w3731 & w4712;
assign w14055 = ~w17613 & ~w13536;
assign w14056 = w15782 & ~w1324;
assign w14057 = w16958 & w12535;
assign w14058 = (~w11104 & w1278) | (~w11104 & w18177) | (w1278 & w18177);
assign w14059 = ~w7185 & ~w16048;
assign w14060 = w2343 & ~w7093;
assign w14061 = ~w15225 & w18827;
assign w14062 = w9626 & ~w2442;
assign w14063 = (w2352 & w13558) | (w2352 & ~w1320) | (w13558 & ~w1320);
assign w14064 = ~w9446 & ~w3237;
assign w14065 = a_22 & a_47;
assign w14066 = ~w3646 & ~w13464;
assign w14067 = ~w6393 & ~w9846;
assign w14068 = (w15399 & w17780) | (w15399 & w19107) | (w17780 & w19107);
assign w14069 = ~w9708 & ~w6292;
assign w14070 = w785 & w10688;
assign w14071 = a_13 & a_59;
assign w14072 = ~w8799 & ~w8796;
assign w14073 = w13312 & ~w13134;
assign w14074 = w3006 & w13893;
assign w14075 = (~w18519 & ~w2743) | (~w18519 & w4596) | (~w2743 & w4596);
assign w14076 = w2888 & ~w3852;
assign w14077 = ~w6846 & ~w10014;
assign w14078 = a_21 & a_43;
assign w14079 = w11510 & ~w12614;
assign w14080 = w15624 & ~w9447;
assign w14081 = ~w16997 & ~w16298;
assign w14082 = a_31 & a_61;
assign w14083 = w10625 & w16411;
assign w14084 = ~w2260 & ~w13922;
assign w14085 = w14670 & w18559;
assign w14086 = ~w12429 & ~w10686;
assign w14087 = ~w7673 & w1621;
assign w14088 = ~w16517 & w5787;
assign w14089 = w2747 & w14224;
assign w14090 = ~w18695 & ~w9758;
assign w14091 = w6340 & w2746;
assign w14092 = w2573 & ~w6160;
assign w14093 = ~w15998 & ~w15075;
assign w14094 = (~w6390 & ~w16754) | (~w6390 & w12186) | (~w16754 & w12186);
assign w14095 = (w17513 & w5743) | (w17513 & w17920) | (w5743 & w17920);
assign w14096 = ~w14458 & w453;
assign w14097 = ~w5760 & w11675;
assign w14098 = w16063 & w5081;
assign w14099 = w15829 & ~w2929;
assign w14100 = w18764 & ~w2357;
assign w14101 = ~w8706 & ~w7769;
assign w14102 = w13003 & ~w18979;
assign w14103 = a_38 & a_39;
assign w14104 = w4381 & w5606;
assign w14105 = ~w12879 & ~w6179;
assign w14106 = a_19 & a_43;
assign w14107 = w817 & w14922;
assign w14108 = ~w18130 & w4874;
assign w14109 = ~w3588 & ~w15800;
assign w14110 = w13596 & w8572;
assign w14111 = ~w11565 & ~w6258;
assign w14112 = ~w11059 & w5419;
assign w14113 = w7049 & ~w17816;
assign w14114 = ~w18936 & ~w6479;
assign w14115 = ~w14209 & ~w19108;
assign w14116 = ~w10132 & ~w15651;
assign w14117 = w4143 & ~w11212;
assign w14118 = a_6 & a_28;
assign w14119 = ~w13365 & w7270;
assign w14120 = w2965 & ~w17792;
assign w14121 = ~w11846 & ~w17027;
assign w14122 = a_14 & a_42;
assign w14123 = ~w8421 & ~w14966;
assign w14124 = w12485 & ~w17843;
assign w14125 = ~w16211 & w11419;
assign w14126 = ~w9678 & ~w6894;
assign w14127 = a_0 & a_3;
assign w14128 = ~w17467 & ~w16466;
assign w14129 = w13332 & ~w2321;
assign w14130 = ~w15169 & ~w15186;
assign w14131 = w4250 & w14292;
assign w14132 = ~w6152 & ~w4853;
assign w14133 = (~w3852 & w12285) | (~w3852 & w14076) | (w12285 & w14076);
assign w14134 = a_7 & a_50;
assign w14135 = w18601 & ~w6524;
assign w14136 = ~w13 & w5817;
assign w14137 = w10909 & ~w18049;
assign w14138 = a_27 & a_52;
assign w14139 = ~w8782 & ~w1371;
assign w14140 = ~w502 & ~w14641;
assign w14141 = ~w6588 & w7622;
assign w14142 = ~w17946 & w17242;
assign w14143 = w10669 & ~w1709;
assign w14144 = ~w223 & ~w8133;
assign w14145 = ~w3500 & ~w8222;
assign w14146 = w1906 & w18431;
assign w14147 = a_26 & a_61;
assign w14148 = w246 & w8120;
assign w14149 = a_20 & a_53;
assign w14150 = a_14 & a_52;
assign w14151 = w17369 & ~w12848;
assign w14152 = (~w16175 & w2769) | (~w16175 & w11831) | (w2769 & w11831);
assign w14153 = (~w15953 & ~w8382) | (~w15953 & w15006) | (~w8382 & w15006);
assign w14154 = w17081 & ~w2865;
assign w14155 = w18313 & w11961;
assign w14156 = ~w2801 & w10802;
assign w14157 = w18829 & ~w7145;
assign w14158 = w1879 & ~w1665;
assign w14159 = w5686 & w467;
assign w14160 = w9376 & w11365;
assign w14161 = ~w12297 & ~w394;
assign w14162 = ~w14194 & w8935;
assign w14163 = w10231 & ~w3695;
assign w14164 = ~w3196 & w8622;
assign w14165 = a_34 & a_46;
assign w14166 = ~w5819 & ~w12158;
assign w14167 = a_16 & a_63;
assign w14168 = ~w1039 & ~w11499;
assign w14169 = ~w12029 & ~w17007;
assign w14170 = a_6 & a_9;
assign w14171 = a_14 & a_59;
assign w14172 = ~w1581 & ~w5445;
assign w14173 = ~w8525 & ~w12666;
assign w14174 = ~w16055 & ~w5534;
assign w14175 = ~w18188 & w16121;
assign w14176 = ~w8301 & ~w4876;
assign w14177 = ~w12275 & w17825;
assign w14178 = ~w10234 & w8048;
assign w14179 = ~w18831 & w7063;
assign w14180 = w6988 & w5296;
assign w14181 = a_3 & a_33;
assign w14182 = w15139 & w17552;
assign w14183 = a_38 & a_42;
assign w14184 = w17396 & w10432;
assign w14185 = (~w8486 & ~w15837) | (~w8486 & w618) | (~w15837 & w618);
assign w14186 = w15247 & ~w15256;
assign w14187 = ~w12268 & w15927;
assign w14188 = ~w1262 & ~w11051;
assign w14189 = ~w13807 & ~w5393;
assign w14190 = ~w1351 & w9743;
assign w14191 = w17489 & ~w8038;
assign w14192 = ~w14359 & w15092;
assign w14193 = ~w16289 & ~w3894;
assign w14194 = a_15 & a_34;
assign w14195 = w10933 & ~w12136;
assign w14196 = a_42 & a_60;
assign w14197 = a_20 & a_43;
assign w14198 = w4092 & ~w14396;
assign w14199 = a_18 & a_20;
assign w14200 = ~w5116 & ~w3587;
assign w14201 = a_0 & a_34;
assign w14202 = ~w4220 & ~w5246;
assign w14203 = w1212 & w8692;
assign w14204 = ~w229 & ~w4732;
assign w14205 = w9615 & ~w1926;
assign w14206 = (w17667 & w13082) | (w17667 & w10408) | (w13082 & w10408);
assign w14207 = ~w2782 & ~w4378;
assign w14208 = ~w13168 & w2204;
assign w14209 = ~w5571 & ~w1166;
assign w14210 = ~w14200 & ~w10536;
assign w14211 = (~w1551 & ~w1318) | (~w1551 & w16467) | (~w1318 & w16467);
assign w14212 = w10147 & w2713;
assign w14213 = ~w12552 & w137;
assign w14214 = w15984 & w18748;
assign w14215 = w13466 & w3491;
assign w14216 = a_33 & a_63;
assign w14217 = ~w16906 & ~w773;
assign w14218 = ~w16679 & ~w10628;
assign w14219 = w15594 & w15313;
assign w14220 = (~w12931 & w14031) | (~w12931 & w1059) | (w14031 & w1059);
assign w14221 = (~w12378 & ~w18170) | (~w12378 & w18114) | (~w18170 & w18114);
assign w14222 = w12222 & ~w6698;
assign w14223 = ~w11434 & ~w9241;
assign w14224 = (~w3475 & ~w8317) | (~w3475 & w319) | (~w8317 & w319);
assign w14225 = w2969 & w9323;
assign w14226 = w10468 & ~w428;
assign w14227 = w14551 & w10986;
assign w14228 = w13082 & ~w3175;
assign w14229 = ~w18134 & ~w14166;
assign w14230 = ~w15653 & ~w9144;
assign w14231 = a_8 & a_29;
assign w14232 = (~w8341 & w12897) | (~w8341 & w6956) | (w12897 & w6956);
assign w14233 = w15144 & w8628;
assign w14234 = w7621 & w772;
assign w14235 = w16238 & w11442;
assign w14236 = ~w16706 & w9467;
assign w14237 = w14831 & ~w416;
assign w14238 = ~w15833 & w5724;
assign w14239 = a_27 & a_32;
assign w14240 = ~w17482 & ~w15404;
assign w14241 = w8175 & ~w18670;
assign w14242 = w17549 & w551;
assign w14243 = ~w18192 & ~w16825;
assign w14244 = ~w1002 & ~w5994;
assign w14245 = ~w8950 & w11771;
assign w14246 = ~w4644 & ~w8333;
assign w14247 = ~w4895 & ~w4842;
assign w14248 = ~w7182 & ~w638;
assign w14249 = ~w13176 & ~w7437;
assign w14250 = ~w18847 & ~w795;
assign w14251 = a_1 & a_35;
assign w14252 = ~w10885 & ~w4336;
assign w14253 = ~w14112 & ~w9558;
assign w14254 = a_19 & a_47;
assign w14255 = ~w16905 & ~w5524;
assign w14256 = (~w18870 & w10330) | (~w18870 & w355) | (w10330 & w355);
assign w14257 = w15665 & w5175;
assign w14258 = ~w14771 & w4524;
assign w14259 = ~w1397 & ~w3408;
assign w14260 = w6438 & w4284;
assign w14261 = ~w1827 & ~w528;
assign w14262 = ~w15179 & ~w13802;
assign w14263 = w14384 & ~w5725;
assign w14264 = a_0 & a_50;
assign w14265 = ~w9791 & ~w7827;
assign w14266 = ~w10335 & ~w8805;
assign w14267 = ~w12670 & ~w17764;
assign w14268 = w6853 & w12456;
assign w14269 = ~w19005 & w17995;
assign w14270 = ~w11444 & ~w1055;
assign w14271 = w10542 & ~w7193;
assign w14272 = w4918 & ~w17703;
assign w14273 = (~w11396 & w5927) | (~w11396 & w13662) | (w5927 & w13662);
assign w14274 = ~w11180 & w4935;
assign w14275 = ~w8662 & ~w5228;
assign w14276 = w18364 & w1560;
assign w14277 = ~w2752 & ~w19048;
assign w14278 = ~w17326 & w1553;
assign w14279 = ~w6730 & ~w11475;
assign w14280 = ~w16282 & ~w10931;
assign w14281 = ~w11009 & w12041;
assign w14282 = ~w12385 & ~w1619;
assign w14283 = ~w6787 & w843;
assign w14284 = ~w17971 & ~w6073;
assign w14285 = ~w9963 & w8238;
assign w14286 = a_3 & a_38;
assign w14287 = ~w7336 & ~w9751;
assign w14288 = ~w17987 & ~w11936;
assign w14289 = w10534 & ~w6503;
assign w14290 = a_42 & a_55;
assign w14291 = w18150 & ~w8569;
assign w14292 = ~w11602 & ~w18111;
assign w14293 = w13008 & ~w17193;
assign w14294 = a_24 & a_36;
assign w14295 = ~w8357 & w11552;
assign w14296 = ~w12904 & w6136;
assign w14297 = ~w3886 & ~w456;
assign w14298 = (~w750 & ~w13884) | (~w750 & w10492) | (~w13884 & w10492);
assign w14299 = a_34 & w18633;
assign w14300 = ~w13315 & ~w6355;
assign w14301 = ~w5465 & w2624;
assign w14302 = ~w15303 & ~w12520;
assign w14303 = w17292 | w11523;
assign w14304 = ~w13302 & w16747;
assign w14305 = a_25 & a_56;
assign w14306 = ~w9448 & ~w4362;
assign w14307 = ~w11403 & w858;
assign w14308 = ~w17183 & ~w14927;
assign w14309 = w4083 & w2687;
assign w14310 = (~w5787 & w6688) | (~w5787 & w16459) | (w6688 & w16459);
assign w14311 = ~w16912 & w12638;
assign w14312 = w7545 & w7464;
assign w14313 = ~w5097 & w289;
assign w14314 = ~w15941 & ~w15180;
assign w14315 = w17054 & ~w8465;
assign w14316 = a_18 & a_37;
assign w14317 = w3975 & ~w9666;
assign w14318 = w17476 & ~w12828;
assign w14319 = ~w14374 & ~w4288;
assign w14320 = w14127 & w18528;
assign w14321 = ~w7067 & ~w254;
assign w14322 = ~w1567 & ~w15884;
assign w14323 = a_3 & a_10;
assign w14324 = ~w18553 & w15772;
assign w14325 = ~w1258 & ~w10342;
assign w14326 = (w3189 & w12) | (w3189 & w6489) | (w12 & w6489);
assign w14327 = w8362 & w15875;
assign w14328 = ~w2308 & ~w4283;
assign w14329 = (w6516 & w12398) | (w6516 & w6350) | (w12398 & w6350);
assign w14330 = a_21 & a_44;
assign w14331 = (~w16103 & ~w3360) | (~w16103 & w13710) | (~w3360 & w13710);
assign w14332 = ~w17344 & ~w1091;
assign w14333 = a_20 & a_55;
assign w14334 = w14204 & ~w3675;
assign w14335 = a_53 & a_54;
assign w14336 = w2420 & ~w6305;
assign w14337 = w11866 & ~w4789;
assign w14338 = ~w8765 & w7078;
assign w14339 = w15644 & ~w13232;
assign w14340 = ~w3469 & w17888;
assign w14341 = ~w17150 & ~w352;
assign w14342 = ~w12977 & ~w14925;
assign w14343 = w310 & ~w688;
assign w14344 = a_38 & a_50;
assign w14345 = ~w1747 & ~w17013;
assign w14346 = ~w5682 & ~w13206;
assign w14347 = ~w825 & ~w9828;
assign w14348 = a_13 & a_35;
assign w14349 = ~w10753 & ~w1129;
assign w14350 = w4998 & ~w1999;
assign w14351 = ~w17452 & ~w11293;
assign w14352 = ~w8352 & ~w15414;
assign w14353 = ~w3250 & ~w18631;
assign w14354 = ~w2627 & ~w7415;
assign w14355 = ~w4408 & ~w6063;
assign w14356 = a_11 & a_45;
assign w14357 = ~w13615 & ~w12076;
assign w14358 = w6969 & ~w19047;
assign w14359 = (~w2486 & ~w14598) | (~w2486 & w9237) | (~w14598 & w9237);
assign w14360 = ~w8767 & ~w6779;
assign w14361 = ~w7010 & ~w14844;
assign w14362 = a_44 & a_46;
assign w14363 = w13647 & ~w5191;
assign w14364 = ~w12947 & ~w2286;
assign w14365 = ~w3912 & ~w7707;
assign w14366 = w3658 & ~w18293;
assign w14367 = ~w3073 & ~w18256;
assign w14368 = w10624 & w3653;
assign w14369 = w16755 & ~w13261;
assign w14370 = w12331 & ~w1403;
assign w14371 = w11024 & ~w13108;
assign w14372 = a_2 & a_19;
assign w14373 = ~w1736 & ~w962;
assign w14374 = ~w5690 & ~w13322;
assign w14375 = ~w8578 & ~w6893;
assign w14376 = w4909 & ~w9253;
assign w14377 = w9390 & w3867;
assign w14378 = w15808 & ~w11057;
assign w14379 = w3861 & w11398;
assign w14380 = w3431 & w3077;
assign w14381 = (~w707 & ~w7915) | (~w707 & w7428) | (~w7915 & w7428);
assign w14382 = w9742 & ~w15754;
assign w14383 = a_4 & a_39;
assign w14384 = ~w16852 & ~w1814;
assign w14385 = ~w11118 & w13270;
assign w14386 = w10460 & w19184;
assign w14387 = a_9 & a_13;
assign w14388 = ~w15579 & w9969;
assign w14389 = w2304 & ~w1510;
assign w14390 = ~w3314 & w1279;
assign w14391 = ~w17681 & ~w3362;
assign w14392 = ~w16693 & w11281;
assign w14393 = ~w6780 & ~w11072;
assign w14394 = ~w10080 & ~w5560;
assign w14395 = ~w7990 & ~w11233;
assign w14396 = ~w8219 & ~w18021;
assign w14397 = w6752 & ~w17235;
assign w14398 = (~w6955 & ~w8611) | (~w6955 & w1156) | (~w8611 & w1156);
assign w14399 = ~w18494 & ~w6645;
assign w14400 = ~w6732 & ~w392;
assign w14401 = a_10 & a_62;
assign w14402 = w17466 & ~w15187;
assign w14403 = a_1 & a_26;
assign w14404 = ~w10199 & ~w761;
assign w14405 = ~w16727 & ~w7119;
assign w14406 = ~w1191 & ~w4933;
assign w14407 = ~w205 & w1605;
assign w14408 = ~w9707 & ~w10366;
assign w14409 = ~w15147 & ~w18617;
assign w14410 = a_4 & a_50;
assign w14411 = w4763 & w9850;
assign w14412 = (w5296 & w9337) | (w5296 & w159) | (w9337 & w159);
assign w14413 = w4566 & ~w215;
assign w14414 = ~w14961 & ~w13177;
assign w14415 = ~w1122 & ~w18299;
assign w14416 = ~w13221 & w9595;
assign w14417 = ~w5146 & ~w16734;
assign w14418 = a_2 & a_56;
assign w14419 = w13585 & w12656;
assign w14420 = ~w1724 & w16222;
assign w14421 = ~w13603 & w7038;
assign w14422 = ~w6568 & ~w14049;
assign w14423 = ~w2660 & w221;
assign w14424 = ~w18413 & w6828;
assign w14425 = (w4979 & w10330) | (w4979 & w4326) | (w10330 & w4326);
assign w14426 = ~w5690 & ~w2155;
assign w14427 = (~w4261 & ~w8819) | (~w4261 & w10707) | (~w8819 & w10707);
assign w14428 = a_33 & a_41;
assign w14429 = ~w17630 & w13143;
assign w14430 = w13377 & w13508;
assign w14431 = ~w2437 & ~w7359;
assign w14432 = ~w10155 & w4275;
assign w14433 = ~w6687 & ~w16065;
assign w14434 = w5378 & w3699;
assign w14435 = (~w16090 & ~w11056) | (~w16090 & w18075) | (~w11056 & w18075);
assign w14436 = ~w7344 & ~w1423;
assign w14437 = ~w8375 & ~w2821;
assign w14438 = ~w9614 & ~w16968;
assign w14439 = ~w15152 & ~w14846;
assign w14440 = ~w14382 & w7380;
assign w14441 = a_2 & a_12;
assign w14442 = ~w5035 & ~w15226;
assign w14443 = ~w11405 & ~w15613;
assign w14444 = ~w18930 & ~w10244;
assign w14445 = w15427 & ~w13364;
assign w14446 = w1738 & ~w9052;
assign w14447 = ~w12244 & ~w4215;
assign w14448 = ~w9615 & w1926;
assign w14449 = ~w7987 & ~w10369;
assign w14450 = ~w10034 & ~w11767;
assign w14451 = a_44 & a_47;
assign w14452 = ~w14156 & ~w15833;
assign w14453 = w12468 & ~w8851;
assign w14454 = ~w8617 & ~w7093;
assign w14455 = ~w6147 & ~w16030;
assign w14456 = (~w7555 & ~w10206) | (~w7555 & w16924) | (~w10206 & w16924);
assign w14457 = ~w13243 & ~w3035;
assign w14458 = ~w12410 & ~w11863;
assign w14459 = ~w17606 & ~w8823;
assign w14460 = ~w8471 & w4357;
assign w14461 = ~w15363 & ~w16752;
assign w14462 = ~w13141 & ~w3212;
assign w14463 = w13302 & ~w16747;
assign w14464 = (~w8543 & w488) | (~w8543 & w16330) | (w488 & w16330);
assign w14465 = ~w14993 & w1576;
assign w14466 = (~w14892 & ~w3059) | (~w14892 & w10458) | (~w3059 & w10458);
assign w14467 = w5189 & ~w2459;
assign w14468 = w18985 & ~w11555;
assign w14469 = ~w17043 & ~w10687;
assign w14470 = w8781 & ~w7953;
assign w14471 = w9700 & ~w95;
assign w14472 = a_0 & a_16;
assign w14473 = a_1 & a_33;
assign w14474 = ~w17635 & ~w17722;
assign w14475 = a_1 & a_12;
assign w14476 = w12222 & ~w7726;
assign w14477 = ~w10387 & ~w17846;
assign w14478 = ~w15904 & w17206;
assign w14479 = (~w10038 & w16242) | (~w10038 & w16480) | (w16242 & w16480);
assign w14480 = ~w1581 & ~w16837;
assign w14481 = ~w5501 & ~w14918;
assign w14482 = ~w11657 & ~w13824;
assign w14483 = w18813 & w7488;
assign w14484 = ~w8502 & ~w6198;
assign w14485 = ~w1142 & w13160;
assign w14486 = ~w559 & ~w10586;
assign w14487 = a_13 & a_27;
assign w14488 = (w15755 & w12168) | (w15755 & w13935) | (w12168 & w13935);
assign w14489 = ~w2925 & ~w16333;
assign w14490 = w6951 & ~w6719;
assign w14491 = ~w5443 & ~w3248;
assign w14492 = a_0 & a_55;
assign w14493 = ~w2921 & w6454;
assign w14494 = ~w17680 & ~w3284;
assign w14495 = ~w16243 & ~w3928;
assign w14496 = w17505 & w15958;
assign w14497 = w19122 & ~w1205;
assign w14498 = ~w853 & ~w17642;
assign w14499 = w2457 & ~w15161;
assign w14500 = ~w1573 & ~w16610;
assign w14501 = ~w15947 & ~w18971;
assign w14502 = ~w11973 & w15022;
assign w14503 = w14623 & ~w9663;
assign w14504 = ~w14291 & ~w1376;
assign w14505 = w1057 & ~w9705;
assign w14506 = ~w16735 & ~w501;
assign w14507 = ~w2725 & ~w16081;
assign w14508 = ~w3041 & ~w14749;
assign w14509 = ~w15705 & w5119;
assign w14510 = w8334 & ~w17079;
assign w14511 = ~w8293 & ~w2492;
assign w14512 = ~w15777 & w12148;
assign w14513 = ~w6943 & w15769;
assign w14514 = ~w6433 & ~w16371;
assign w14515 = w16362 & ~w11182;
assign w14516 = ~w12830 & ~w9759;
assign w14517 = ~w3769 & ~w11066;
assign w14518 = ~w1731 & ~w3577;
assign w14519 = (~w7341 & w9386) | (~w7341 & w11946) | (w9386 & w11946);
assign w14520 = a_20 & a_38;
assign w14521 = (~w7687 & ~w3775) | (~w7687 & w16470) | (~w3775 & w16470);
assign w14522 = ~w10410 & ~w13045;
assign w14523 = ~w15913 & ~w6861;
assign w14524 = (w3009 & w1142) | (w3009 & w1798) | (w1142 & w1798);
assign w14525 = (~w12801 & w8800) | (~w12801 & w7130) | (w8800 & w7130);
assign w14526 = ~w3341 & w13599;
assign w14527 = ~w7572 & ~w720;
assign w14528 = ~w3920 & ~w1478;
assign w14529 = ~w7545 & ~w8901;
assign w14530 = ~w2622 & w10877;
assign w14531 = ~w10045 & ~w16874;
assign w14532 = w139 & ~w44;
assign w14533 = ~w10610 & ~w6755;
assign w14534 = ~w7073 & ~w10944;
assign w14535 = ~w4153 & ~w16273;
assign w14536 = ~w2908 & ~w12630;
assign w14537 = ~w3057 & ~w17642;
assign w14538 = w760 & ~w2282;
assign w14539 = ~w4234 & ~w14829;
assign w14540 = ~w5085 & ~w14863;
assign w14541 = ~w10519 & ~w7957;
assign w14542 = (w7341 & w9069) | (w7341 & w6201) | (w9069 & w6201);
assign w14543 = ~w9716 & w10235;
assign w14544 = w6514 & w13666;
assign w14545 = ~w11092 & ~w4781;
assign w14546 = ~w7440 & ~w6608;
assign w14547 = ~w978 & ~w18599;
assign w14548 = ~w1890 & ~w792;
assign w14549 = w16785 & ~w472;
assign w14550 = ~w899 & ~w7217;
assign w14551 = a_7 & a_43;
assign w14552 = ~w53 & ~w7977;
assign w14553 = ~w9232 & ~w775;
assign w14554 = w14965 & ~w12970;
assign w14555 = w16121 & ~w14213;
assign w14556 = ~w12954 & w8549;
assign w14557 = ~w17657 & ~w16698;
assign w14558 = ~w1360 & ~w13540;
assign w14559 = ~w18056 & ~w6214;
assign w14560 = w12877 & w7578;
assign w14561 = w16849 & ~w8225;
assign w14562 = ~w6585 & ~w1028;
assign w14563 = ~w13724 & w8509;
assign w14564 = w14451 & w17246;
assign w14565 = w3236 & ~w18937;
assign w14566 = a_47 & a_55;
assign w14567 = w9698 & ~w1120;
assign w14568 = w6849 & ~w15784;
assign w14569 = ~w11349 & ~w3661;
assign w14570 = w15934 & w12490;
assign w14571 = w6030 & w3373;
assign w14572 = ~w5290 & ~w15729;
assign w14573 = w15350 & ~w9391;
assign w14574 = ~w1492 & ~w5478;
assign w14575 = ~w823 & w8783;
assign w14576 = w694 & ~w13105;
assign w14577 = ~w2579 & w15527;
assign w14578 = ~w3742 & ~w18590;
assign w14579 = ~w7507 & ~w1052;
assign w14580 = ~w8607 & ~w6722;
assign w14581 = w4948 & w4001;
assign w14582 = w12753 & ~w10680;
assign w14583 = w18678 & ~w9693;
assign w14584 = a_63 & a_1;
assign w14585 = ~w9289 & ~w10601;
assign w14586 = (~w1634 & w5541) | (~w1634 & w9720) | (w5541 & w9720);
assign w14587 = w5421 & w16582;
assign w14588 = ~w13765 & w10415;
assign w14589 = ~w6763 & ~w2939;
assign w14590 = ~w17840 & ~w16354;
assign w14591 = ~w8191 & ~w13014;
assign w14592 = w4542 & ~w12909;
assign w14593 = ~w14243 & ~w6851;
assign w14594 = w18396 & ~w960;
assign w14595 = a_7 & a_33;
assign w14596 = ~w9301 & ~w13336;
assign w14597 = ~w18313 & ~w11961;
assign w14598 = ~w2486 & ~w17875;
assign w14599 = w13749 & w16227;
assign w14600 = ~w1031 & ~w15403;
assign w14601 = ~w86 & w18078;
assign w14602 = ~w16794 & ~w4628;
assign w14603 = a_50 & a_59;
assign w14604 = ~w17983 & ~w5451;
assign w14605 = ~w8070 & ~w11497;
assign w14606 = ~w9260 & w17632;
assign w14607 = ~w6604 & ~w2721;
assign w14608 = a_45 & a_57;
assign w14609 = w17994 & ~w7233;
assign w14610 = w16178 & ~w261;
assign w14611 = w1320 & w2350;
assign w14612 = ~w7538 & w18172;
assign w14613 = ~w14038 & ~w2164;
assign w14614 = ~w10001 & ~w4480;
assign w14615 = ~w1740 & ~w4252;
assign w14616 = w8903 & w5212;
assign w14617 = a_30 & a_41;
assign w14618 = a_18 & a_21;
assign w14619 = w13049 & ~w13092;
assign w14620 = ~w14997 & ~w11841;
assign w14621 = ~w7180 & ~w14457;
assign w14622 = (~w5906 & ~w16693) | (~w5906 & w9879) | (~w16693 & w9879);
assign w14623 = ~w879 & ~w14246;
assign w14624 = w6277 & ~w11531;
assign w14625 = (~w5857 & ~w11182) | (~w5857 & w5671) | (~w11182 & w5671);
assign w14626 = ~w13585 & ~w10332;
assign w14627 = w15411 & ~w18780;
assign w14628 = ~w6372 & w10218;
assign w14629 = w16594 & w16885;
assign w14630 = ~w16087 & w4335;
assign w14631 = (w4355 & w5743) | (w4355 & w11179) | (w5743 & w11179);
assign w14632 = ~w14349 & ~w10328;
assign w14633 = w5043 & w14890;
assign w14634 = (~w11639 & ~w18152) | (~w11639 & w11347) | (~w18152 & w11347);
assign w14635 = w18492 & w437;
assign w14636 = (~w11827 & ~w10796) | (~w11827 & w7210) | (~w10796 & w7210);
assign w14637 = a_7 & a_49;
assign w14638 = ~w18558 & w3825;
assign w14639 = w12559 & ~w2643;
assign w14640 = w11062 & w3759;
assign w14641 = ~w3972 & ~w2866;
assign w14642 = ~w4983 & ~w1155;
assign w14643 = ~w14332 & w7755;
assign w14644 = ~w6047 & ~w6837;
assign w14645 = w6588 & ~w7622;
assign w14646 = ~w8844 & ~w2745;
assign w14647 = ~w16558 & ~w3812;
assign w14648 = w2622 & ~w10877;
assign w14649 = w14812 & w4921;
assign w14650 = ~w724 & w14221;
assign w14651 = ~w13111 & w17084;
assign w14652 = ~w7426 & ~w11411;
assign w14653 = a_21 & a_56;
assign w14654 = ~w2316 & ~w12661;
assign w14655 = w17551 & w6814;
assign w14656 = (~w3661 & ~w14569) | (~w3661 & w919) | (~w14569 & w919);
assign w14657 = ~w2980 & w1268;
assign w14658 = ~w15970 & w11737;
assign w14659 = ~w14239 & ~w3092;
assign w14660 = ~w9062 & ~w13262;
assign w14661 = ~w13579 & w6765;
assign w14662 = ~w11655 & ~w892;
assign w14663 = w12697 & w11638;
assign w14664 = ~w18544 & ~w1573;
assign w14665 = (w7610 & w6125) | (w7610 & w10424) | (w6125 & w10424);
assign w14666 = ~w3931 & ~w13474;
assign w14667 = (~w16855 & ~w15083) | (~w16855 & w15467) | (~w15083 & w15467);
assign w14668 = a_19 & a_31;
assign w14669 = ~w8296 & ~w3474;
assign w14670 = ~w5746 & w8005;
assign w14671 = w13182 & w4446;
assign w14672 = ~w10589 & ~w8818;
assign w14673 = w14123 & w8216;
assign w14674 = ~w17612 & ~w607;
assign w14675 = ~w5529 & ~w11766;
assign w14676 = ~w16321 & ~w8895;
assign w14677 = (w1962 & w452) | (w1962 & w3519) | (w452 & w3519);
assign w14678 = ~w12589 & ~w11885;
assign w14679 = ~w17536 & ~w8622;
assign w14680 = w3688 & ~w6010;
assign w14681 = w17899 & ~w212;
assign w14682 = ~w16915 & w12724;
assign w14683 = a_45 & a_58;
assign w14684 = ~w3438 & ~w12681;
assign w14685 = ~w8958 & ~w6930;
assign w14686 = ~w3652 & ~w19095;
assign w14687 = ~w18168 & ~w13132;
assign w14688 = w13024 & ~w14762;
assign w14689 = a_23 & a_50;
assign w14690 = a_30 & a_43;
assign w14691 = w3139 & ~w6993;
assign w14692 = ~w13501 & ~w4684;
assign w14693 = w2776 & ~w15864;
assign w14694 = ~w4182 & ~w7715;
assign w14695 = ~w17501 & ~w16507;
assign w14696 = w7985 & w12494;
assign w14697 = w634 & w5017;
assign w14698 = ~w9330 & w6874;
assign w14699 = ~w8737 & ~w10065;
assign w14700 = w11545 & ~w6559;
assign w14701 = a_15 & a_27;
assign w14702 = w14719 & w17732;
assign w14703 = ~w3121 & w12130;
assign w14704 = w15395 & w371;
assign w14705 = ~w7684 & ~w14271;
assign w14706 = ~w12652 & ~w249;
assign w14707 = ~w3293 & w14993;
assign w14708 = ~w7365 & ~w18104;
assign w14709 = ~w8677 & ~w13654;
assign w14710 = w3955 & w16847;
assign w14711 = (~w11660 & ~w2524) | (~w11660 & w17372) | (~w2524 & w17372);
assign w14712 = ~w1174 & w688;
assign w14713 = ~w12246 & w3719;
assign w14714 = a_15 & a_38;
assign w14715 = ~w8427 & ~w15874;
assign w14716 = ~w2797 & ~w9866;
assign w14717 = ~w12919 & w5712;
assign w14718 = w3570 & w3190;
assign w14719 = ~w9358 & ~w12190;
assign w14720 = w8382 & ~w1123;
assign w14721 = ~w7129 & w7235;
assign w14722 = a_29 & a_41;
assign w14723 = ~w73 & ~w13446;
assign w14724 = ~w16600 & ~w2212;
assign w14725 = a_48 & a_53;
assign w14726 = ~w7168 & ~w2749;
assign w14727 = ~w151 & ~w5162;
assign w14728 = w12562 & ~w16697;
assign w14729 = w13073 & ~w3958;
assign w14730 = ~w10175 & ~w11348;
assign w14731 = w12274 & ~w8585;
assign w14732 = w1097 & ~w5479;
assign w14733 = ~w16546 & w5356;
assign w14734 = ~w3733 & ~w6852;
assign w14735 = ~w6907 & ~w3052;
assign w14736 = w12390 & ~w6866;
assign w14737 = ~w5415 & w18222;
assign w14738 = w14830 & ~w12856;
assign w14739 = ~w1772 & w9853;
assign w14740 = ~w14323 & ~w11713;
assign w14741 = ~w11116 & ~w14988;
assign w14742 = ~w15713 & ~w16676;
assign w14743 = ~w427 & ~w4336;
assign w14744 = a_17 & a_50;
assign w14745 = w1488 & w13455;
assign w14746 = ~w13833 & ~w13085;
assign w14747 = ~w10469 & ~w5810;
assign w14748 = ~w14044 & ~w2517;
assign w14749 = ~w2975 & ~w1701;
assign w14750 = ~w5516 & w8281;
assign w14751 = a_8 & a_54;
assign w14752 = ~w4566 & w215;
assign w14753 = ~w14670 & ~w8267;
assign w14754 = a_14 & a_21;
assign w14755 = ~w7616 & ~w9100;
assign w14756 = a_26 & a_53;
assign w14757 = w11485 & ~w4545;
assign w14758 = ~w17779 & ~w2680;
assign w14759 = a_7 & a_56;
assign w14760 = ~w9913 & ~w16024;
assign w14761 = ~w1364 & w13681;
assign w14762 = ~w6599 & ~w8684;
assign w14763 = ~w3838 & ~w7108;
assign w14764 = ~w15132 & ~w11953;
assign w14765 = ~w8984 & ~w2673;
assign w14766 = ~w6853 & w7596;
assign w14767 = ~w6377 & ~w14878;
assign w14768 = ~w11136 & w1625;
assign w14769 = ~w61 & ~w4930;
assign w14770 = ~w18334 & ~w430;
assign w14771 = a_16 & a_33;
assign w14772 = ~w15642 & ~w7221;
assign w14773 = ~w8021 & ~w965;
assign w14774 = w5646 & w1392;
assign w14775 = ~w17285 & ~w7782;
assign w14776 = ~w6803 & ~w11338;
assign w14777 = ~w8341 & ~w11445;
assign w14778 = ~w7089 & ~w125;
assign w14779 = ~w13317 & ~w19089;
assign w14780 = w15796 & ~w10331;
assign w14781 = ~w18688 & w473;
assign w14782 = w10009 & ~w3336;
assign w14783 = a_2 & a_11;
assign w14784 = ~a_28 & ~w9010;
assign w14785 = w14240 & w18735;
assign w14786 = ~w12720 & w18492;
assign w14787 = ~w12904 & ~w11949;
assign w14788 = ~w7244 & ~w12748;
assign w14789 = ~w2664 & ~w6607;
assign w14790 = a_36 & a_52;
assign w14791 = ~w15373 & ~w10871;
assign w14792 = ~w7445 & w58;
assign w14793 = ~w1151 & ~w7176;
assign w14794 = ~a_23 & ~w7048;
assign w14795 = w9803 & w1871;
assign w14796 = ~w5329 & ~w18465;
assign w14797 = ~w13518 & ~w13103;
assign w14798 = a_28 & a_59;
assign w14799 = w2643 & ~w16966;
assign w14800 = ~w955 & ~w18472;
assign w14801 = w6249 & ~w17352;
assign w14802 = ~w906 & ~w11526;
assign w14803 = w4477 & ~w13201;
assign w14804 = w16092 & ~w3882;
assign w14805 = w13732 & ~w5076;
assign w14806 = w12436 & ~w6624;
assign w14807 = ~w1077 & ~w4464;
assign w14808 = w2075 & ~w10134;
assign w14809 = ~w18958 & ~w6232;
assign w14810 = w4790 & ~w4130;
assign w14811 = w13505 & w10047;
assign w14812 = a_12 & a_23;
assign w14813 = ~w16840 & ~w8913;
assign w14814 = ~w11023 & w4870;
assign w14815 = ~w11390 & w6085;
assign w14816 = ~w17337 & w4024;
assign w14817 = ~w17892 & w9329;
assign w14818 = w9415 & w17125;
assign w14819 = ~w9808 & ~w7460;
assign w14820 = ~w2134 & ~w17176;
assign w14821 = w5132 & w18322;
assign w14822 = ~w5636 & ~w18944;
assign w14823 = w7115 & w1508;
assign w14824 = w7576 & w19185;
assign w14825 = ~a_50 & a_51;
assign w14826 = ~w13016 & ~w14002;
assign w14827 = (~w16020 & ~w15283) | (~w16020 & w8376) | (~w15283 & w8376);
assign w14828 = (~w6152 & ~w14132) | (~w6152 & w4843) | (~w14132 & w4843);
assign w14829 = ~w13785 & w7339;
assign w14830 = ~w3424 & ~w3676;
assign w14831 = ~w9836 & w14972;
assign w14832 = ~w9009 & ~w6518;
assign w14833 = ~w13390 & ~w8211;
assign w14834 = ~w5825 & w9876;
assign w14835 = ~w11659 & w15578;
assign w14836 = ~w7153 & ~w18744;
assign w14837 = w16332 & w7928;
assign w14838 = ~w1533 & ~w613;
assign w14839 = w3938 & ~w1822;
assign w14840 = (~w2769 & w16242) | (~w2769 & w14479) | (w16242 & w14479);
assign w14841 = a_5 & a_46;
assign w14842 = ~w17483 & ~w768;
assign w14843 = ~w149 & ~w522;
assign w14844 = ~w10313 & ~w858;
assign w14845 = w8646 & w16993;
assign w14846 = ~w5980 & ~w7476;
assign w14847 = w1633 & ~w3010;
assign w14848 = w16562 & w19069;
assign w14849 = ~w3326 & ~w2244;
assign w14850 = ~w2150 & w756;
assign w14851 = ~w4050 & ~w7306;
assign w14852 = a_18 & a_23;
assign w14853 = ~w305 & ~w3917;
assign w14854 = w17285 & w7782;
assign w14855 = ~w18417 & ~w13784;
assign w14856 = ~w17586 & ~w3947;
assign w14857 = ~w11927 & w12845;
assign w14858 = (w7604 & w16136) | (w7604 & w13979) | (w16136 & w13979);
assign w14859 = ~w16537 & w5316;
assign w14860 = ~w14183 & ~w6413;
assign w14861 = ~w9 & w10186;
assign w14862 = ~w11190 & ~w17918;
assign w14863 = ~w2878 & w10141;
assign w14864 = ~w14395 & ~w17941;
assign w14865 = ~w6112 & w18063;
assign w14866 = ~w16672 & ~w13157;
assign w14867 = a_33 & a_60;
assign w14868 = a_17 & a_62;
assign w14869 = w3314 & ~w3380;
assign w14870 = w17524 & w12489;
assign w14871 = w5641 & w1639;
assign w14872 = a_15 & a_31;
assign w14873 = w17295 & w5362;
assign w14874 = (w2769 & w5156) | (w2769 & w14975) | (w5156 & w14975);
assign w14875 = ~w4237 & ~w6807;
assign w14876 = ~w6559 & ~w9211;
assign w14877 = (w2396 & w13082) | (w2396 & w5791) | (w13082 & w5791);
assign w14878 = ~w2144 & ~w13181;
assign w14879 = ~w10330 & w7905;
assign w14880 = ~w17712 & ~w11896;
assign w14881 = ~w15523 & ~w984;
assign w14882 = ~w18024 & w12745;
assign w14883 = ~w18985 & w11555;
assign w14884 = ~w11686 & w2996;
assign w14885 = ~w12447 & ~w14196;
assign w14886 = ~w5480 & w9524;
assign w14887 = ~w6853 & ~w11244;
assign w14888 = ~w1125 & ~w2440;
assign w14889 = ~w9150 & ~w2956;
assign w14890 = ~w2346 & ~w5250;
assign w14891 = ~w438 & ~w5364;
assign w14892 = w14144 & w6663;
assign w14893 = ~w7161 & ~w11035;
assign w14894 = w7902 & ~w12929;
assign w14895 = ~w10508 & ~w1812;
assign w14896 = a_38 & a_53;
assign w14897 = ~w18792 & ~w16416;
assign w14898 = a_9 & a_27;
assign w14899 = ~w18854 & ~w6342;
assign w14900 = w19069 & ~w949;
assign w14901 = ~w11290 & w13204;
assign w14902 = ~w10663 & ~w10161;
assign w14903 = w11143 & w970;
assign w14904 = ~w9413 & ~w11882;
assign w14905 = ~w18214 & ~w15359;
assign w14906 = ~w7105 & ~w7791;
assign w14907 = ~w17573 & w7978;
assign w14908 = ~w12855 & ~w15440;
assign w14909 = w16849 & ~w6922;
assign w14910 = a_2 & a_34;
assign w14911 = w13661 & w1153;
assign w14912 = w14374 & w4288;
assign w14913 = ~w3683 & ~w7154;
assign w14914 = ~w18014 & ~w8601;
assign w14915 = ~w3741 & ~w6086;
assign w14916 = ~w11084 & ~w9535;
assign w14917 = w3811 & ~w513;
assign w14918 = ~w7844 & w14607;
assign w14919 = ~w12457 & ~w16791;
assign w14920 = ~w10007 & ~w1433;
assign w14921 = (~w4676 & ~w5780) | (~w4676 & w4160) | (~w5780 & w4160);
assign w14922 = a_2 & a_44;
assign w14923 = w3796 & ~w16419;
assign w14924 = ~w11479 & ~w8581;
assign w14925 = w11813 & w1192;
assign w14926 = w2954 & ~w3595;
assign w14927 = ~w5058 & ~w4978;
assign w14928 = ~w2398 & ~w1013;
assign w14929 = ~w10897 & ~w14214;
assign w14930 = ~w2002 & ~w11388;
assign w14931 = ~w6971 & ~w198;
assign w14932 = ~w14756 & ~w8044;
assign w14933 = w16998 & w11070;
assign w14934 = ~w10812 & ~w4951;
assign w14935 = a_6 & a_14;
assign w14936 = a_54 & a_55;
assign w14937 = ~w12242 & ~w9393;
assign w14938 = ~w5435 & ~w6378;
assign w14939 = ~w7768 & w10155;
assign w14940 = (~w8170 & ~w12495) | (~w8170 & w4919) | (~w12495 & w4919);
assign w14941 = ~w2937 & ~w3256;
assign w14942 = ~w12562 & ~w9772;
assign w14943 = ~w12298 & ~w2986;
assign w14944 = ~w9489 & ~w3553;
assign w14945 = w18257 & ~w11868;
assign w14946 = ~w2216 & ~w16152;
assign w14947 = w6987 & ~w14001;
assign w14948 = ~w2281 & ~w1582;
assign w14949 = ~w12487 & ~w2867;
assign w14950 = ~w13140 & ~w488;
assign w14951 = w9045 & ~w4000;
assign w14952 = ~w6027 & w1561;
assign w14953 = ~w13672 & ~w11885;
assign w14954 = ~w18784 & ~w10925;
assign w14955 = ~w11177 & ~w14227;
assign w14956 = ~w14341 & ~w2926;
assign w14957 = ~w636 & ~w3903;
assign w14958 = ~w7508 & ~w6251;
assign w14959 = w8717 & w10939;
assign w14960 = ~w7043 & ~w3098;
assign w14961 = ~a_54 & w11222;
assign w14962 = w6836 & ~w7628;
assign w14963 = ~w13849 & ~w6861;
assign w14964 = ~w16911 & w5585;
assign w14965 = (~w16835 & ~w124) | (~w16835 & w6582) | (~w124 & w6582);
assign w14966 = ~w13684 & w17142;
assign w14967 = ~w9347 & ~w10671;
assign w14968 = ~w13782 & ~w1702;
assign w14969 = ~w2533 & w3863;
assign w14970 = ~w6798 & w5404;
assign w14971 = w18369 & ~w18164;
assign w14972 = ~w6797 & ~w18888;
assign w14973 = ~w12486 & ~w3758;
assign w14974 = ~w1365 & w9017;
assign w14975 = (w12904 & w7133) | (w12904 & w5156) | (w7133 & w5156);
assign w14976 = ~w11926 & ~w3751;
assign w14977 = ~w3502 & ~w5324;
assign w14978 = a_4 & a_57;
assign w14979 = w372 & w6396;
assign w14980 = (a_60 & w10984) | (a_60 & w16116) | (w10984 & w16116);
assign w14981 = w13164 & w15567;
assign w14982 = a_46 & a_59;
assign w14983 = ~w9574 & w6265;
assign w14984 = ~w16930 & ~w16300;
assign w14985 = a_56 & a_60;
assign w14986 = (a_51 & w1138) | (a_51 & w7031) | (w1138 & w7031);
assign w14987 = ~w9320 & ~w13701;
assign w14988 = ~w11202 & ~w12988;
assign w14989 = w16822 & w10309;
assign w14990 = ~w4400 & ~w12839;
assign w14991 = w14185 & ~w11227;
assign w14992 = ~w9805 & w11807;
assign w14993 = ~w19001 & w7848;
assign w14994 = ~w16544 & w735;
assign w14995 = ~w18025 & w1748;
assign w14996 = a_24 & a_30;
assign w14997 = ~w15591 & ~w9591;
assign w14998 = w13465 & w7167;
assign w14999 = ~w11977 & w3933;
assign w15000 = ~w15792 & ~w4671;
assign w15001 = w5365 & ~w8307;
assign w15002 = ~w17454 & w14625;
assign w15003 = ~w14837 & ~w11589;
assign w15004 = ~w2007 & ~w1438;
assign w15005 = ~w812 & ~w7014;
assign w15006 = w1123 & ~w15953;
assign w15007 = ~w16659 & w18359;
assign w15008 = w1958 & ~w12532;
assign w15009 = (~w18863 & ~w16601) | (~w18863 & w16464) | (~w16601 & w16464);
assign w15010 = a_14 & a_57;
assign w15011 = w16272 & ~w14993;
assign w15012 = ~w10623 & w18394;
assign w15013 = ~w3030 & w13780;
assign w15014 = ~w11672 & ~w13087;
assign w15015 = w11277 & ~w5824;
assign w15016 = ~w2393 & ~w10459;
assign w15017 = ~w16585 & w13860;
assign w15018 = a_16 & a_51;
assign w15019 = a_26 & a_45;
assign w15020 = a_34 & a_49;
assign w15021 = a_51 & a_59;
assign w15022 = ~w6819 & ~w7444;
assign w15023 = ~w3713 & w14111;
assign w15024 = ~w12982 & w17147;
assign w15025 = a_20 & a_58;
assign w15026 = ~w6620 & ~w10985;
assign w15027 = ~w7409 & w6840;
assign w15028 = ~w6742 & ~w14842;
assign w15029 = w422 & ~w10486;
assign w15030 = ~w2965 & w17792;
assign w15031 = w1217 & ~w10326;
assign w15032 = ~w14633 & ~w12506;
assign w15033 = ~w2362 & ~w9367;
assign w15034 = ~w10081 & ~w1609;
assign w15035 = ~w2588 & ~w5504;
assign w15036 = ~w7137 & ~w5428;
assign w15037 = w9330 & ~w6874;
assign w15038 = w16447 & ~w12526;
assign w15039 = ~w5973 & ~w6553;
assign w15040 = w14745 & w19014;
assign w15041 = ~w11263 & ~w1176;
assign w15042 = ~w5140 & ~w7635;
assign w15043 = ~w18017 & w6426;
assign w15044 = w5173 & ~w9519;
assign w15045 = a_13 & a_14;
assign w15046 = w8021 & w965;
assign w15047 = ~w11221 & ~w16645;
assign w15048 = ~w6670 & ~w8366;
assign w15049 = ~w10328 & ~w10753;
assign w15050 = ~w12842 & ~w6945;
assign w15051 = a_8 & a_21;
assign w15052 = a_17 & a_29;
assign w15053 = w2838 & ~w8068;
assign w15054 = ~w10540 & ~w317;
assign w15055 = ~w4387 & ~w8827;
assign w15056 = ~w17932 & ~w1376;
assign w15057 = w10057 & ~w10400;
assign w15058 = w6534 & ~w8208;
assign w15059 = ~w4485 & ~w12870;
assign w15060 = ~w4386 & ~w4086;
assign w15061 = w1386 & w10803;
assign w15062 = (~w8636 & w2175) | (~w8636 & w8665) | (w2175 & w8665);
assign w15063 = ~w7076 & ~w16378;
assign w15064 = ~w8544 & ~w1110;
assign w15065 = ~w8252 & ~w12891;
assign w15066 = w12804 & ~w16642;
assign w15067 = w3143 & ~w8006;
assign w15068 = a_12 & a_32;
assign w15069 = w6349 & ~w5001;
assign w15070 = w9929 & ~w348;
assign w15071 = w5260 & ~w309;
assign w15072 = ~w1202 & w9091;
assign w15073 = ~w7091 & ~w4368;
assign w15074 = ~w90 & ~w7274;
assign w15075 = ~w5017 & w3351;
assign w15076 = ~w2531 & ~w3614;
assign w15077 = a_10 & a_33;
assign w15078 = ~w10956 & ~w17783;
assign w15079 = (~w2769 & w9102) | (~w2769 & w10825) | (w9102 & w10825);
assign w15080 = w15399 & ~w983;
assign w15081 = a_5 & a_6;
assign w15082 = w5507 & w4673;
assign w15083 = ~w16855 & ~w16352;
assign w15084 = (~w1582 & ~w6476) | (~w1582 & w14948) | (~w6476 & w14948);
assign w15085 = ~w1115 & ~w12395;
assign w15086 = ~w14773 & ~w15046;
assign w15087 = w15969 & ~w18551;
assign w15088 = ~w9766 & ~w3214;
assign w15089 = ~w7126 & ~w10493;
assign w15090 = ~w18521 & ~w12582;
assign w15091 = ~w18017 & w18853;
assign w15092 = (~w9443 & ~w16767) | (~w9443 & w16887) | (~w16767 & w16887);
assign w15093 = ~w10420 & ~w18207;
assign w15094 = w10056 & w12224;
assign w15095 = a_27 & a_28;
assign w15096 = w12305 & ~w3891;
assign w15097 = ~w4433 & ~w5584;
assign w15098 = ~w16686 & ~w8952;
assign w15099 = a_6 & a_34;
assign w15100 = a_24 & a_35;
assign w15101 = ~w650 & ~w14697;
assign w15102 = a_35 & a_57;
assign w15103 = w4075 & w17649;
assign w15104 = ~w1755 & ~w9938;
assign w15105 = w4989 & w10033;
assign w15106 = ~w5506 & w17197;
assign w15107 = w3196 & ~w8622;
assign w15108 = a_11 & a_12;
assign w15109 = w927 & ~w8612;
assign w15110 = a_24 & a_27;
assign w15111 = ~w10739 & ~w9624;
assign w15112 = ~w672 & ~w3154;
assign w15113 = ~w2917 & w5607;
assign w15114 = a_0 & a_46;
assign w15115 = (~w17596 & ~w1758) | (~w17596 & w3329) | (~w1758 & w3329);
assign w15116 = a_8 & a_57;
assign w15117 = ~w16768 & ~w10245;
assign w15118 = w19035 & w5904;
assign w15119 = w15711 & ~w18007;
assign w15120 = w11995 & ~w7489;
assign w15121 = a_18 & a_47;
assign w15122 = ~w11648 & ~w17281;
assign w15123 = ~w586 & ~w23;
assign w15124 = ~w13850 & ~w5819;
assign w15125 = w16074 & w5959;
assign w15126 = ~w1237 & w56;
assign w15127 = ~w8236 & w10528;
assign w15128 = a_9 & a_20;
assign w15129 = ~w13275 & w4594;
assign w15130 = w5025 & ~w18423;
assign w15131 = ~w17489 & w8038;
assign w15132 = w15084 & ~w3526;
assign w15133 = ~w19053 & w17539;
assign w15134 = ~w2398 & ~w5664;
assign w15135 = ~w2013 & ~w14186;
assign w15136 = ~w269 & ~w19088;
assign w15137 = ~w6862 & w3394;
assign w15138 = w4045 & ~w18274;
assign w15139 = ~w9431 & ~w14826;
assign w15140 = ~w17781 & ~w9640;
assign w15141 = w271 & ~w8987;
assign w15142 = ~w11683 & w13462;
assign w15143 = ~w2015 & ~w325;
assign w15144 = ~w8534 & ~w10368;
assign w15145 = ~w827 & ~w11034;
assign w15146 = w16731 & w5038;
assign w15147 = ~w7113 & ~w14208;
assign w15148 = ~w18469 & ~w10024;
assign w15149 = ~w5732 & ~w9110;
assign w15150 = ~w2594 & ~w16456;
assign w15151 = a_31 & a_48;
assign w15152 = ~w12522 & ~w17254;
assign w15153 = ~w13938 & ~w9906;
assign w15154 = ~w18636 & w1294;
assign w15155 = w6481 & ~w3540;
assign w15156 = ~w815 & w15765;
assign w15157 = w15018 & w16262;
assign w15158 = (w15306 & w10330) | (w15306 & w13357) | (w10330 & w13357);
assign w15159 = (w1386 & w5527) | (w1386 & w1532) | (w5527 & w1532);
assign w15160 = ~w17511 & ~w4865;
assign w15161 = ~w4984 & ~w14811;
assign w15162 = ~w10607 & ~w12091;
assign w15163 = (~w7102 & w1659) | (~w7102 & w17639) | (w1659 & w17639);
assign w15164 = ~w6514 & ~w4586;
assign w15165 = ~w18449 & ~w9763;
assign w15166 = ~w10738 & ~w7613;
assign w15167 = a_26 & a_31;
assign w15168 = a_25 & a_63;
assign w15169 = w12940 & ~w18903;
assign w15170 = ~w8235 & ~w4231;
assign w15171 = w2034 & w18705;
assign w15172 = ~w17122 & ~w485;
assign w15173 = ~w16497 & w16436;
assign w15174 = ~w6042 & ~w18348;
assign w15175 = w18774 & w3489;
assign w15176 = w1119 | w11949;
assign w15177 = a_15 & a_32;
assign w15178 = ~w16949 & w10319;
assign w15179 = ~w10629 & ~w8036;
assign w15180 = ~a_30 & ~w11865;
assign w15181 = ~w15453 & ~w11670;
assign w15182 = ~w6145 & ~w13820;
assign w15183 = ~w15963 & ~w11114;
assign w15184 = ~w7875 & ~w7831;
assign w15185 = ~w13213 & ~w18098;
assign w15186 = w16820 & w9952;
assign w15187 = ~w12597 & ~w15635;
assign w15188 = ~w2257 & w13108;
assign w15189 = ~a_18 & ~w15994;
assign w15190 = ~w16513 & ~w8379;
assign w15191 = ~w9020 & w16999;
assign w15192 = ~w12968 & ~w13999;
assign w15193 = ~w11083 & ~w10130;
assign w15194 = a_59 & a_63;
assign w15195 = w14924 & w18574;
assign w15196 = w12561 & ~w3525;
assign w15197 = w7117 & w13873;
assign w15198 = ~w18388 & ~w17332;
assign w15199 = ~w16663 & ~w18686;
assign w15200 = ~w2402 & w6975;
assign w15201 = w8250 & w17693;
assign w15202 = ~w18017 & w11002;
assign w15203 = a_32 & a_47;
assign w15204 = ~w14600 & ~w18949;
assign w15205 = (~w10170 & ~w11454) | (~w10170 & w10067) | (~w11454 & w10067);
assign w15206 = ~w17017 & ~w17290;
assign w15207 = ~w16868 & ~w18921;
assign w15208 = ~w6272 & ~w18645;
assign w15209 = a_51 & a_61;
assign w15210 = ~w6884 & ~w793;
assign w15211 = (~w2769 & w3519) | (~w2769 & w14677) | (w3519 & w14677);
assign w15212 = ~w5328 & w1415;
assign w15213 = ~w13712 & ~w13561;
assign w15214 = ~w2017 & w14695;
assign w15215 = ~w17897 & ~w8541;
assign w15216 = w8673 & ~w16222;
assign w15217 = w15935 & ~w9620;
assign w15218 = a_43 & a_46;
assign w15219 = ~w17727 & ~w10202;
assign w15220 = ~w9299 & ~w14865;
assign w15221 = w2572 & ~w17317;
assign w15222 = ~w4940 & ~w5277;
assign w15223 = w6385 & ~w12822;
assign w15224 = ~a_47 & a_48;
assign w15225 = ~w5360 & ~w1004;
assign w15226 = w16198 & w15498;
assign w15227 = a_40 & a_57;
assign w15228 = a_28 & a_31;
assign w15229 = w6650 & ~w16156;
assign w15230 = a_45 & a_51;
assign w15231 = ~w11582 & ~w17569;
assign w15232 = w4373 & w13512;
assign w15233 = w8633 & w5126;
assign w15234 = ~w14670 & ~w1287;
assign w15235 = a_2 & a_43;
assign w15236 = w11782 & ~w12488;
assign w15237 = ~w5475 & ~w18470;
assign w15238 = ~w9710 & ~w14036;
assign w15239 = (~w2330 & w1540) | (~w2330 & w5882) | (w1540 & w5882);
assign w15240 = ~w6392 & ~w6139;
assign w15241 = ~w3321 & ~w9504;
assign w15242 = w3993 & w11900;
assign w15243 = w6426 & w15693;
assign w15244 = ~w17804 & w18226;
assign w15245 = ~w8840 & ~w8899;
assign w15246 = w14047 & w4300;
assign w15247 = ~w5526 & ~w18680;
assign w15248 = a_34 & a_60;
assign w15249 = ~w15990 & ~w15491;
assign w15250 = a_42 & a_54;
assign w15251 = a_38 & a_57;
assign w15252 = ~w5400 & ~w9365;
assign w15253 = ~w9533 & ~w5627;
assign w15254 = w8029 & ~w1367;
assign w15255 = w17653 & ~w18382;
assign w15256 = ~w9363 & ~w14117;
assign w15257 = w5934 & ~w15273;
assign w15258 = ~w9679 & w5391;
assign w15259 = w18993 & ~w14352;
assign w15260 = w15083 & w18320;
assign w15261 = a_17 & a_31;
assign w15262 = ~w17018 & ~w12787;
assign w15263 = w5105 & ~w16869;
assign w15264 = w861 & w17782;
assign w15265 = ~w5669 & ~w13881;
assign w15266 = ~w10502 & ~w14680;
assign w15267 = ~w4544 & ~w17510;
assign w15268 = ~w791 & ~w822;
assign w15269 = ~w13955 & w7;
assign w15270 = ~w13531 & ~w2500;
assign w15271 = ~w3762 & ~w1578;
assign w15272 = ~w9307 & ~w4664;
assign w15273 = ~w16281 & ~w11699;
assign w15274 = ~w4128 & ~w17181;
assign w15275 = ~w11122 & ~w15746;
assign w15276 = ~w14151 & ~w5388;
assign w15277 = ~w5651 & ~w5055;
assign w15278 = ~w7060 & w19052;
assign w15279 = a_44 & a_56;
assign w15280 = ~w11394 & w611;
assign w15281 = ~w679 & ~w17817;
assign w15282 = w12534 & ~w5115;
assign w15283 = ~w16020 & ~w12831;
assign w15284 = w7314 & ~w14820;
assign w15285 = ~w4244 & ~w12896;
assign w15286 = ~w12427 & w4470;
assign w15287 = ~w9886 & ~w8256;
assign w15288 = ~w15566 & ~w5567;
assign w15289 = a_49 & a_62;
assign w15290 = w1284 & w3992;
assign w15291 = a_46 & a_61;
assign w15292 = w14323 & ~w1134;
assign w15293 = w7529 & ~w17948;
assign w15294 = ~w9657 & ~w8190;
assign w15295 = w16563 & ~w1863;
assign w15296 = w713 & ~w8526;
assign w15297 = ~w7039 & w18446;
assign w15298 = ~w4450 & ~w474;
assign w15299 = ~w8433 & w14986;
assign w15300 = w13803 & w15298;
assign w15301 = ~w8645 & w4307;
assign w15302 = ~w6462 & w8809;
assign w15303 = w19022 & w1523;
assign w15304 = ~w11545 & ~w14876;
assign w15305 = w19027 & w1706;
assign w15306 = (w2254 & w13665) | (w2254 & w2400) | (w13665 & w2400);
assign w15307 = (~w15399 & w9270) | (~w15399 & w17151) | (w9270 & w17151);
assign w15308 = ~w11594 & ~w13079;
assign w15309 = ~w7879 & ~w5684;
assign w15310 = ~w11337 & ~w4724;
assign w15311 = w10345 & ~w10644;
assign w15312 = (w12904 & w5657) | (w12904 & w17715) | (w5657 & w17715);
assign w15313 = a_21 & a_24;
assign w15314 = w14714 & w4677;
assign w15315 = ~w2201 & w1640;
assign w15316 = a_0 & a_28;
assign w15317 = w7154 & w7691;
assign w15318 = w18647 & ~w9674;
assign w15319 = ~w12487 & w15535;
assign w15320 = a_29 & a_57;
assign w15321 = ~w7246 & ~w8919;
assign w15322 = ~w584 & ~w7018;
assign w15323 = ~w8083 & w14275;
assign w15324 = w16497 & ~w16436;
assign w15325 = a_27 & a_31;
assign w15326 = ~w6537 & ~w11823;
assign w15327 = ~w3224 & ~w199;
assign w15328 = w11845 & w2882;
assign w15329 = (w7102 & w18651) | (w7102 & w258) | (w18651 & w258);
assign w15330 = ~w18476 & ~w5905;
assign w15331 = ~w4296 & w18720;
assign w15332 = a_17 & a_34;
assign w15333 = ~w2963 & ~w7808;
assign w15334 = w7322 & w10993;
assign w15335 = ~w15453 & ~w17774;
assign w15336 = ~w14020 & ~w17043;
assign w15337 = (~w11001 & w10330) | (~w11001 & w6892) | (w10330 & w6892);
assign w15338 = ~w10574 & ~w13406;
assign w15339 = w17347 & w185;
assign w15340 = ~w16947 & ~w14651;
assign w15341 = ~w13567 & ~w2555;
assign w15342 = ~w2390 & ~w18237;
assign w15343 = w17950 & ~w13156;
assign w15344 = ~w3476 & ~w5125;
assign w15345 = ~w9822 & w2771;
assign w15346 = ~w7304 & ~w5779;
assign w15347 = a_26 & a_52;
assign w15348 = ~w10904 & ~w11815;
assign w15349 = ~w934 & ~w1955;
assign w15350 = ~w13407 & ~w15716;
assign w15351 = ~w1694 & ~w13356;
assign w15352 = ~w7172 & ~w6290;
assign w15353 = (~w803 & ~w8385) | (~w803 & w9056) | (~w8385 & w9056);
assign w15354 = ~w5961 & ~w3307;
assign w15355 = w10765 & w3667;
assign w15356 = w16086 & w5882;
assign w15357 = (~w16641 & ~w11485) | (~w16641 & w5653) | (~w11485 & w5653);
assign w15358 = ~w10251 & ~w4630;
assign w15359 = w3276 & w12077;
assign w15360 = ~w15910 & ~w7817;
assign w15361 = ~w645 & ~w10181;
assign w15362 = ~w13604 & w6132;
assign w15363 = a_41 & a_52;
assign w15364 = w17840 & ~w6510;
assign w15365 = ~w4922 & ~w10682;
assign w15366 = a_47 & a_49;
assign w15367 = ~w5696 & ~w3156;
assign w15368 = ~w18017 & w14976;
assign w15369 = (w10099 & ~w1320) | (w10099 & w1036) | (~w1320 & w1036);
assign w15370 = w13909 & ~w4554;
assign w15371 = ~w13613 & ~w15437;
assign w15372 = ~w14071 & w11770;
assign w15373 = ~w4169 & ~w11837;
assign w15374 = w7408 & w2556;
assign w15375 = ~w18182 & w11714;
assign w15376 = w4965 & ~w10444;
assign w15377 = w4611 & ~w4166;
assign w15378 = ~w13402 & ~w14420;
assign w15379 = w12941 & ~w17964;
assign w15380 = ~w5615 & ~w11958;
assign w15381 = ~w23 & ~w7797;
assign w15382 = w1351 & ~w9743;
assign w15383 = w17481 & w16391;
assign w15384 = ~w15178 & ~w16701;
assign w15385 = ~w18914 & ~w18424;
assign w15386 = ~w1287 & w18559;
assign w15387 = w15894 & w18620;
assign w15388 = w6388 & ~w8671;
assign w15389 = ~w7685 & ~w16351;
assign w15390 = ~w12634 & ~w3451;
assign w15391 = w18672 & ~w18954;
assign w15392 = ~w4530 & ~w16312;
assign w15393 = ~w11402 & ~w802;
assign w15394 = w4692 & ~w6037;
assign w15395 = a_16 & a_17;
assign w15396 = a_4 & a_29;
assign w15397 = (~w10149 & ~w16101) | (~w10149 & w7989) | (~w16101 & w7989);
assign w15398 = w7800 & ~w6314;
assign w15399 = ~w7610 & w11742;
assign w15400 = ~w18607 & ~w4573;
assign w15401 = ~w17033 & ~w4782;
assign w15402 = a_14 & a_28;
assign w15403 = ~w17840 & ~w6374;
assign w15404 = w16813 & ~w16750;
assign w15405 = ~w13011 & ~w10343;
assign w15406 = ~w9278 & w14796;
assign w15407 = ~w5809 & ~w2140;
assign w15408 = (~w5526 & ~w15247) | (~w5526 & w9488) | (~w15247 & w9488);
assign w15409 = w8909 & ~w5644;
assign w15410 = w323 & ~w19075;
assign w15411 = a_14 & a_32;
assign w15412 = w5973 & w6553;
assign w15413 = ~w12703 & ~w18315;
assign w15414 = ~w17260 & ~w334;
assign w15415 = (~w8452 & w12398) | (~w8452 & w2566) | (w12398 & w2566);
assign w15416 = w1113 & ~w15659;
assign w15417 = w7492 & ~w17891;
assign w15418 = ~w2495 & ~w16960;
assign w15419 = w5239 & w14348;
assign w15420 = (~w9253 & w12982) | (~w9253 & w14376) | (w12982 & w14376);
assign w15421 = ~w11776 & w2444;
assign w15422 = a_16 & a_32;
assign w15423 = ~w9224 & ~w13740;
assign w15424 = (w17995 & w10330) | (w17995 & w16) | (w10330 & w16);
assign w15425 = ~w7013 & ~w18612;
assign w15426 = ~w10845 & w9903;
assign w15427 = ~w1401 & ~w12455;
assign w15428 = a_12 & a_35;
assign w15429 = (~w11814 & ~w7538) | (~w11814 & w5242) | (~w7538 & w5242);
assign w15430 = ~w3466 & ~w6437;
assign w15431 = ~w4187 & w5396;
assign w15432 = w9452 & w3504;
assign w15433 = (~w74 & ~w8996) | (~w74 & w7045) | (~w8996 & w7045);
assign w15434 = a_2 & a_60;
assign w15435 = w17886 & w12649;
assign w15436 = ~w11009 & ~w5714;
assign w15437 = w17088 & w13292;
assign w15438 = w7910 & w368;
assign w15439 = w2075 & ~w740;
assign w15440 = ~w9434 & ~w10528;
assign w15441 = ~w5302 & ~w3902;
assign w15442 = ~w12374 & ~w16182;
assign w15443 = a_21 & a_54;
assign w15444 = w9859 & ~w12882;
assign w15445 = w942 & ~w6691;
assign w15446 = w13131 & ~w1226;
assign w15447 = (~w3160 & ~w13621) | (~w3160 & w7648) | (~w13621 & w7648);
assign w15448 = ~w16920 & w10698;
assign w15449 = w5545 & ~w11069;
assign w15450 = w5532 & ~w857;
assign w15451 = ~w1721 & ~w14502;
assign w15452 = ~w14841 & ~w1;
assign w15453 = w406 & w14669;
assign w15454 = ~w10651 & ~w6879;
assign w15455 = w7860 & w9387;
assign w15456 = ~w17316 & ~w248;
assign w15457 = w16172 & w13585;
assign w15458 = ~w6218 & ~w13618;
assign w15459 = w14375 & w6166;
assign w15460 = ~w5384 & w13874;
assign w15461 = w3167 & w2813;
assign w15462 = ~w11150 & w15181;
assign w15463 = ~w5978 & w1164;
assign w15464 = a_1 & a_6;
assign w15465 = ~w17982 & w2931;
assign w15466 = w10660 & ~w18674;
assign w15467 = ~w18320 & ~w16855;
assign w15468 = ~w8507 & ~w5286;
assign w15469 = ~w4522 & w3690;
assign w15470 = ~w8955 & w11096;
assign w15471 = w2457 & w8201;
assign w15472 = ~w13457 & ~w16290;
assign w15473 = a_35 & a_36;
assign w15474 = ~w16532 & ~w2232;
assign w15475 = w12001 & w588;
assign w15476 = w19003 & w16674;
assign w15477 = w17185 & ~w7657;
assign w15478 = ~w1158 & ~w3449;
assign w15479 = ~w7940 & ~w9423;
assign w15480 = w14028 & ~w463;
assign w15481 = ~w10813 & ~w9571;
assign w15482 = ~w7631 & ~w65;
assign w15483 = ~w1745 & ~w15917;
assign w15484 = ~w11251 & ~w10250;
assign w15485 = w1678 & ~w5630;
assign w15486 = ~w17284 & ~w10520;
assign w15487 = ~w13552 & ~w1218;
assign w15488 = w11506 & ~w4513;
assign w15489 = ~w14831 & w416;
assign w15490 = ~w16427 & ~w10476;
assign w15491 = ~w12963 & ~w17935;
assign w15492 = a_16 & a_34;
assign w15493 = w7029 & w9781;
assign w15494 = (~w13679 & ~w11594) | (~w13679 & w15891) | (~w11594 & w15891);
assign w15495 = ~w3776 & ~w1756;
assign w15496 = w10639 & ~w10238;
assign w15497 = w16959 & w16109;
assign w15498 = ~w13885 & ~w16268;
assign w15499 = ~a_56 & a_57;
assign w15500 = w9598 & ~w15896;
assign w15501 = ~w8353 & ~w2800;
assign w15502 = ~w13221 & ~w3826;
assign w15503 = (~w10330 & w17646) | (~w10330 & w13775) | (w17646 & w13775);
assign w15504 = ~w15096 & ~w12299;
assign w15505 = ~w18773 & w6678;
assign w15506 = ~w4595 & ~w10263;
assign w15507 = a_4 & a_60;
assign w15508 = w5981 & w683;
assign w15509 = ~w836 & ~w12416;
assign w15510 = ~w7967 & ~w10685;
assign w15511 = (~w12541 & ~w18636) | (~w12541 & w2628) | (~w18636 & w2628);
assign w15512 = w7355 & ~w17867;
assign w15513 = ~w17218 & w11472;
assign w15514 = a_12 & a_13;
assign w15515 = ~w7632 & ~w10694;
assign w15516 = ~w3187 & ~w3789;
assign w15517 = a_1 & a_23;
assign w15518 = ~w11041 & ~w5429;
assign w15519 = ~w3048 & ~w4422;
assign w15520 = ~w10921 & ~w1180;
assign w15521 = w4347 & w4797;
assign w15522 = ~w15807 & ~w9490;
assign w15523 = w1778 & ~w15429;
assign w15524 = ~w31 & w12818;
assign w15525 = a_16 & a_23;
assign w15526 = ~w7605 & ~w492;
assign w15527 = ~w6880 & ~w8694;
assign w15528 = w4421 & w14047;
assign w15529 = ~w12477 & ~w12388;
assign w15530 = w15595 & ~w1306;
assign w15531 = a_39 & a_52;
assign w15532 = ~w3308 & ~w12169;
assign w15533 = ~w4549 & w18566;
assign w15534 = w555 & w5170;
assign w15535 = ~w6178 & w14893;
assign w15536 = w12906 & w15569;
assign w15537 = w8243 & ~w9269;
assign w15538 = ~w2769 & w11790;
assign w15539 = ~w1253 & w12315;
assign w15540 = ~w12222 & w6698;
assign w15541 = a_18 & a_22;
assign w15542 = (~w9332 & ~w10487) | (~w9332 & w12173) | (~w10487 & w12173);
assign w15543 = ~w8426 & w14282;
assign w15544 = ~w15030 & ~w14120;
assign w15545 = ~w2534 & ~w18009;
assign w15546 = ~w1902 & ~w18729;
assign w15547 = ~w14837 & ~w8348;
assign w15548 = ~w18336 & w13650;
assign w15549 = w10614 & ~w9483;
assign w15550 = ~w10377 & ~w14527;
assign w15551 = ~w13295 & w2345;
assign w15552 = a_36 & a_38;
assign w15553 = w11549 & w3123;
assign w15554 = a_17 & a_36;
assign w15555 = a_41 & a_60;
assign w15556 = w1408 & ~w13756;
assign w15557 = ~w15205 & w7250;
assign w15558 = ~w5161 & ~w17541;
assign w15559 = ~w3693 & ~w3067;
assign w15560 = ~w8604 & ~w13242;
assign w15561 = w1661 & ~w3523;
assign w15562 = ~w7505 & ~w7923;
assign w15563 = ~w9493 & ~w13173;
assign w15564 = a_38 & a_61;
assign w15565 = w17359 & ~w3619;
assign w15566 = w6782 & w7427;
assign w15567 = a_8 & a_39;
assign w15568 = ~w14194 & ~w8571;
assign w15569 = ~w13100 & ~w6522;
assign w15570 = w5439 & ~w2173;
assign w15571 = ~w13501 & ~w10771;
assign w15572 = ~w16505 & ~w11338;
assign w15573 = ~w17654 & ~w13307;
assign w15574 = ~w15236 & ~w8152;
assign w15575 = (~w16284 & ~w994) | (~w16284 & w9380) | (~w994 & w9380);
assign w15576 = w4598 & ~w3350;
assign w15577 = ~w18000 & ~w2180;
assign w15578 = ~w13089 & w12347;
assign w15579 = ~w8991 & ~w8869;
assign w15580 = ~w4790 & w4130;
assign w15581 = ~w8817 & ~w6077;
assign w15582 = ~w3014 & ~w8934;
assign w15583 = w3858 & w3586;
assign w15584 = (~w8307 & ~w7829) | (~w8307 & w15001) | (~w7829 & w15001);
assign w15585 = ~w895 & w5227;
assign w15586 = w5868 & w18468;
assign w15587 = w14134 & w9598;
assign w15588 = ~w11687 & ~w617;
assign w15589 = w13169 & ~w9275;
assign w15590 = w13291 & ~w4173;
assign w15591 = ~w973 & ~w7347;
assign w15592 = ~w6100 & ~w6306;
assign w15593 = a_35 & a_46;
assign w15594 = a_22 & a_23;
assign w15595 = ~w10549 & ~w15383;
assign w15596 = ~w7945 & ~w256;
assign w15597 = ~w9780 & ~w7007;
assign w15598 = ~w5889 & ~w5476;
assign w15599 = w5738 & w16232;
assign w15600 = w4556 & ~w1948;
assign w15601 = a_30 & a_39;
assign w15602 = ~w10154 & ~w4012;
assign w15603 = w18350 & ~w13723;
assign w15604 = w4107 & ~w13225;
assign w15605 = ~w2837 & ~w5351;
assign w15606 = w18958 & w6232;
assign w15607 = w13295 & ~w2345;
assign w15608 = ~w3476 & ~w18166;
assign w15609 = w8503 & w257;
assign w15610 = w5859 & w5112;
assign w15611 = ~w1267 & ~w3302;
assign w15612 = ~w18978 & ~w17719;
assign w15613 = ~w6708 & ~w2415;
assign w15614 = w16475 & w5133;
assign w15615 = ~w11189 & ~w9787;
assign w15616 = ~w5900 & ~w17114;
assign w15617 = w7722 & ~w15625;
assign w15618 = ~w11017 & ~w13969;
assign w15619 = a_22 & a_36;
assign w15620 = w9814 & w10074;
assign w15621 = ~w10000 & ~w15665;
assign w15622 = a_6 & a_60;
assign w15623 = ~w10995 & ~w13252;
assign w15624 = ~w6045 & ~w9411;
assign w15625 = ~w5118 & ~w8254;
assign w15626 = w18147 & ~w2933;
assign w15627 = ~w482 & ~w3868;
assign w15628 = ~w15423 & w17400;
assign w15629 = a_9 & a_23;
assign w15630 = a_0 & a_19;
assign w15631 = ~w16071 & ~w15300;
assign w15632 = w18562 & ~w7149;
assign w15633 = ~w17310 & ~w980;
assign w15634 = ~w8241 & ~w1359;
assign w15635 = w1935 & w17161;
assign w15636 = a_26 & a_59;
assign w15637 = ~w6719 & ~w15587;
assign w15638 = ~w4713 & ~w16811;
assign w15639 = w8034 & w16035;
assign w15640 = w9512 & ~w5376;
assign w15641 = ~w9154 & w15845;
assign w15642 = ~w5895 & ~w16311;
assign w15643 = ~w13003 & ~w4955;
assign w15644 = ~w999 & w13150;
assign w15645 = ~w6214 & ~w13981;
assign w15646 = w8597 & ~w9498;
assign w15647 = (~w13577 & w16916) | (~w13577 & w5114) | (w16916 & w5114);
assign w15648 = ~w13534 & ~w17255;
assign w15649 = a_13 & a_39;
assign w15650 = ~w3493 & ~w15069;
assign w15651 = ~w409 & ~w10757;
assign w15652 = ~w18321 & ~w15878;
assign w15653 = ~w690 & ~w11765;
assign w15654 = ~a_6 & ~w7098;
assign w15655 = ~w18759 & ~w8689;
assign w15656 = ~w3780 & ~w5245;
assign w15657 = a_10 & a_40;
assign w15658 = ~w10516 & w6863;
assign w15659 = ~w13060 & ~w11379;
assign w15660 = w15225 & ~w18827;
assign w15661 = ~w18866 & ~w13989;
assign w15662 = w8896 & w6178;
assign w15663 = a_9 & a_34;
assign w15664 = w3059 & w8428;
assign w15665 = ~w16200 & ~w15983;
assign w15666 = ~w6420 & w14188;
assign w15667 = w16206 & ~w11089;
assign w15668 = (~w15026 & w10693) | (~w15026 & w7208) | (w10693 & w7208);
assign w15669 = ~w2917 & ~w6116;
assign w15670 = w19055 & ~w14885;
assign w15671 = ~w11742 & w1596;
assign w15672 = w16546 & w3839;
assign w15673 = w18085 & ~w5698;
assign w15674 = ~w381 & ~w9587;
assign w15675 = ~w7825 & ~w19001;
assign w15676 = ~w587 & ~w6282;
assign w15677 = ~w6293 & w9157;
assign w15678 = ~w13882 & ~w8995;
assign w15679 = ~w8503 & ~w257;
assign w15680 = ~w17310 & ~w12312;
assign w15681 = w15010 & w7705;
assign w15682 = (a_44 & w11965) | (a_44 & w10716) | (w11965 & w10716);
assign w15683 = (~w12255 & w11985) | (~w12255 & w6255) | (w11985 & w6255);
assign w15684 = ~w1025 & ~w10423;
assign w15685 = a_5 & a_9;
assign w15686 = ~w211 & ~w9145;
assign w15687 = ~w18696 & ~w19111;
assign w15688 = ~w3335 & ~w11155;
assign w15689 = w4208 & ~w1641;
assign w15690 = w14734 & ~w13964;
assign w15691 = ~w16942 & ~w7629;
assign w15692 = ~w14845 & ~w887;
assign w15693 = ~w7610 & w12104;
assign w15694 = (w8045 & w2769) | (w8045 & w10265) | (w2769 & w10265);
assign w15695 = w5919 & ~w2329;
assign w15696 = ~w8054 & ~w9255;
assign w15697 = ~w11644 & w15424;
assign w15698 = ~w7821 & ~w6019;
assign w15699 = w676 & ~w15516;
assign w15700 = w6511 & w10742;
assign w15701 = a_15 & a_54;
assign w15702 = (w5743 & w3465) | (w5743 & w9706) | (w3465 & w9706);
assign w15703 = w13861 & w18813;
assign w15704 = ~w7320 & ~w15966;
assign w15705 = w7881 & w7309;
assign w15706 = a_31 & a_32;
assign w15707 = ~w1506 & ~w976;
assign w15708 = ~w12798 & ~w6625;
assign w15709 = ~w3064 & ~w16029;
assign w15710 = ~w464 & ~w7802;
assign w15711 = w9648 & ~w10125;
assign w15712 = ~w5484 & ~w13112;
assign w15713 = (~w2657 & w18646) | (~w2657 & w10976) | (w18646 & w10976);
assign w15714 = ~w811 & ~w9948;
assign w15715 = ~w1696 & ~w1322;
assign w15716 = ~w18525 & ~w11056;
assign w15717 = w1489 & ~w9947;
assign w15718 = w4491 & ~w16152;
assign w15719 = ~w8370 & ~w16608;
assign w15720 = ~w15861 & w2526;
assign w15721 = a_48 & a_50;
assign w15722 = ~w6184 & ~w705;
assign w15723 = ~w17576 & w1242;
assign w15724 = ~w3459 & w17694;
assign w15725 = a_13 & a_58;
assign w15726 = a_25 & a_60;
assign w15727 = ~w7064 & ~w5171;
assign w15728 = a_42 & a_49;
assign w15729 = w2374 & w12052;
assign w15730 = ~w12325 & ~w2773;
assign w15731 = w1679 & ~w11629;
assign w15732 = ~w10896 & w16681;
assign w15733 = ~w1877 & ~w4701;
assign w15734 = ~w3128 & ~w18039;
assign w15735 = w2413 & ~w1127;
assign w15736 = ~w11146 & w11174;
assign w15737 = w4502 & ~w12009;
assign w15738 = w18702 & ~w14578;
assign w15739 = ~w9580 & w824;
assign w15740 = ~w8124 & ~w17014;
assign w15741 = ~w11081 & ~w14704;
assign w15742 = (~w14429 & w9396) | (~w14429 & w5474) | (w9396 & w5474);
assign w15743 = ~w11106 & w7142;
assign w15744 = w6102 & ~w11653;
assign w15745 = ~w10262 & w13651;
assign w15746 = w16900 & w2961;
assign w15747 = ~w10846 & ~w383;
assign w15748 = ~w4368 & ~w332;
assign w15749 = (~w1145 & ~w1057) | (~w1145 & w8914) | (~w1057 & w8914);
assign w15750 = ~w9267 & w3986;
assign w15751 = ~w14566 & ~w9854;
assign w15752 = w9014 & w826;
assign w15753 = a_11 & a_58;
assign w15754 = ~w13873 & ~w11401;
assign w15755 = ~w18272 & w18128;
assign w15756 = w5929 & ~w1765;
assign w15757 = w14302 & ~w6675;
assign w15758 = w2925 & w16333;
assign w15759 = ~w16413 & ~w10857;
assign w15760 = ~w9226 & ~w14732;
assign w15761 = ~w5629 & w4486;
assign w15762 = w10697 & ~w16515;
assign w15763 = ~w7129 & w5706;
assign w15764 = ~w17067 & ~w10829;
assign w15765 = ~w8757 & ~w1530;
assign w15766 = w16826 & w7857;
assign w15767 = ~w11791 & ~w11137;
assign w15768 = ~w13962 & ~w14337;
assign w15769 = ~w3829 & ~w19029;
assign w15770 = ~w3136 & w13549;
assign w15771 = ~w15620 & w1537;
assign w15772 = ~w12905 & ~w5083;
assign w15773 = ~w1038 & ~w3728;
assign w15774 = ~w9461 & w19186;
assign w15775 = ~w1904 & w18639;
assign w15776 = (~w11789 & w8143) | (~w11789 & w10194) | (w8143 & w10194);
assign w15777 = (~w7854 & ~w9557) | (~w7854 & w10579) | (~w9557 & w10579);
assign w15778 = w19057 & w9004;
assign w15779 = ~w9616 & ~w14664;
assign w15780 = ~w18151 & ~w18403;
assign w15781 = ~w15030 & w14287;
assign w15782 = ~w18721 & ~w3914;
assign w15783 = w31 & ~w12818;
assign w15784 = ~w11463 & ~w12129;
assign w15785 = a_13 & a_22;
assign w15786 = ~w7714 & ~w10655;
assign w15787 = w7086 & ~w18087;
assign w15788 = ~w9946 & ~w11299;
assign w15789 = a_19 & a_53;
assign w15790 = ~w9476 & w17157;
assign w15791 = ~w2243 & ~w957;
assign w15792 = ~w6095 & ~w2692;
assign w15793 = ~w282 & ~w7966;
assign w15794 = ~w6595 & ~w14696;
assign w15795 = (~w19046 & ~w1320) | (~w19046 & w8497) | (~w1320 & w8497);
assign w15796 = (~w1644 & ~w11235) | (~w1644 & w4508) | (~w11235 & w4508);
assign w15797 = ~w848 & ~w9499;
assign w15798 = a_62 & w14032;
assign w15799 = w11340 & w14985;
assign w15800 = ~w13522 & w5315;
assign w15801 = ~w3033 & ~w10777;
assign w15802 = ~w11040 & w12125;
assign w15803 = ~w15576 & ~w2920;
assign w15804 = ~w15626 & ~w5248;
assign w15805 = (~w8542 & ~w2593) | (~w8542 & w6129) | (~w2593 & w6129);
assign w15806 = (~w17699 & ~w11076) | (~w17699 & w9800) | (~w11076 & w9800);
assign w15807 = w9348 & ~w7516;
assign w15808 = ~w13797 & ~w4564;
assign w15809 = ~w11579 & ~w16139;
assign w15810 = w18496 & ~w3624;
assign w15811 = w6453 & ~w1597;
assign w15812 = (~w8967 & ~w18433) | (~w8967 & w12806) | (~w18433 & w12806);
assign w15813 = ~w12751 & w5695;
assign w15814 = ~w15114 & ~w17435;
assign w15815 = ~w8433 & ~w14380;
assign w15816 = w2988 & w4856;
assign w15817 = ~w8264 & w1750;
assign w15818 = ~a_4 & ~w15464;
assign w15819 = ~w8013 & w18076;
assign w15820 = w11194 & ~w14931;
assign w15821 = a_20 & a_31;
assign w15822 = ~w16246 & ~w14138;
assign w15823 = ~w11881 & ~w9589;
assign w15824 = ~w17970 & ~w3282;
assign w15825 = w19063 & w11667;
assign w15826 = w12805 & ~w6061;
assign w15827 = ~w94 & ~w169;
assign w15828 = w13164 & ~w17535;
assign w15829 = ~w2233 & ~w4879;
assign w15830 = a_47 & a_52;
assign w15831 = ~w18430 & ~w7831;
assign w15832 = ~w3790 & w18508;
assign w15833 = w2801 & ~w10802;
assign w15834 = ~w18096 & ~w13385;
assign w15835 = ~a_22 & ~w12083;
assign w15836 = a_26 & a_47;
assign w15837 = ~w244 & ~w8486;
assign w15838 = ~w8643 & w8854;
assign w15839 = ~w14240 & ~w18735;
assign w15840 = w16131 & w259;
assign w15841 = a_2 & a_63;
assign w15842 = ~w13581 & w2850;
assign w15843 = a_1 & a_22;
assign w15844 = w6229 & ~w14436;
assign w15845 = ~w16901 & ~w10837;
assign w15846 = w14071 & ~w11770;
assign w15847 = ~w10465 & ~w7265;
assign w15848 = ~w3635 & ~w11951;
assign w15849 = ~w13919 & ~w3485;
assign w15850 = ~w11391 & w19187;
assign w15851 = ~w13229 & ~w12927;
assign w15852 = w11014 & w13619;
assign w15853 = w17855 & w3534;
assign w15854 = ~w14812 & ~w4921;
assign w15855 = ~w13630 & ~w4526;
assign w15856 = w413 & ~w17770;
assign w15857 = ~w13273 & ~w4431;
assign w15858 = ~w8960 & ~w7283;
assign w15859 = ~w7447 & ~w11778;
assign w15860 = w5384 & ~w13874;
assign w15861 = w7594 & w14053;
assign w15862 = (~w18980 & w8635) | (~w18980 & w18041) | (w8635 & w18041);
assign w15863 = ~w18623 & ~w8821;
assign w15864 = ~w17224 & w6598;
assign w15865 = ~w5839 & ~w6783;
assign w15866 = ~w7800 & w6314;
assign w15867 = ~w15439 & ~w5995;
assign w15868 = ~w1464 & ~w15545;
assign w15869 = ~w6500 & w665;
assign w15870 = ~w15818 & ~w6481;
assign w15871 = ~w5515 & ~w11729;
assign w15872 = a_40 & a_60;
assign w15873 = ~w2655 & ~w3678;
assign w15874 = ~w8834 & ~w16454;
assign w15875 = a_27 & a_59;
assign w15876 = w16097 & ~w2759;
assign w15877 = (~w3840 & ~w13116) | (~w3840 & w10799) | (~w13116 & w10799);
assign w15878 = ~w4950 & ~w16573;
assign w15879 = ~w12255 & w7015;
assign w15880 = w9201 & w15361;
assign w15881 = w15495 & w8949;
assign w15882 = (~w12227 & ~w18645) | (~w12227 & w12013) | (~w18645 & w12013);
assign w15883 = w11883 & w7972;
assign w15884 = w20 & w14075;
assign w15885 = ~w4344 & ~w16516;
assign w15886 = ~w4037 & w1825;
assign w15887 = ~w12673 & w18993;
assign w15888 = w13700 & w1715;
assign w15889 = ~w14309 & ~w13215;
assign w15890 = ~w4456 & ~w2744;
assign w15891 = ~w13079 & ~w13679;
assign w15892 = ~w6068 & ~w411;
assign w15893 = ~w1320 & ~w4766;
assign w15894 = a_7 & a_9;
assign w15895 = ~w5845 & ~w3205;
assign w15896 = ~w8305 & ~w17993;
assign w15897 = ~w10367 & ~w1610;
assign w15898 = a_21 & a_34;
assign w15899 = a_4 & a_37;
assign w15900 = w10984 & ~w10454;
assign w15901 = ~w10834 & ~w5318;
assign w15902 = a_38 & a_60;
assign w15903 = ~w8283 & ~w10021;
assign w15904 = ~w15426 & ~w14800;
assign w15905 = w7965 & w616;
assign w15906 = w3603 & ~w16481;
assign w15907 = w227 & ~w1137;
assign w15908 = ~w2192 & w8945;
assign w15909 = (~w6428 & ~w7561) | (~w6428 & w17900) | (~w7561 & w17900);
assign w15910 = a_11 & a_37;
assign w15911 = a_19 & a_50;
assign w15912 = w1441 & ~w7448;
assign w15913 = ~w3051 & ~w12286;
assign w15914 = ~w9598 & w15896;
assign w15915 = w3087 & ~w9349;
assign w15916 = w6521 & w8100;
assign w15917 = ~w5562 & w11661;
assign w15918 = ~w12853 & ~w10911;
assign w15919 = w16585 & ~w13860;
assign w15920 = w7134 & ~w10531;
assign w15921 = ~w11395 & ~w8403;
assign w15922 = w927 & w945;
assign w15923 = ~w6212 & ~w7519;
assign w15924 = w3996 & w17404;
assign w15925 = w9840 & ~w4495;
assign w15926 = ~w393 & ~w9760;
assign w15927 = ~w4831 & ~w7200;
assign w15928 = (~w1956 & ~w7022) | (~w1956 & w10006) | (~w7022 & w10006);
assign w15929 = (w12616 & w2769) | (w12616 & w605) | (w2769 & w605);
assign w15930 = ~w13080 & ~w17110;
assign w15931 = ~w17653 & w18382;
assign w15932 = ~w6557 & ~w1932;
assign w15933 = ~w15084 & ~w18154;
assign w15934 = (~w17569 & ~w8189) | (~w17569 & w15231) | (~w8189 & w15231);
assign w15935 = ~w4354 & ~w14369;
assign w15936 = ~w7445 & w16241;
assign w15937 = ~w17473 & ~w5783;
assign w15938 = w15123 & ~w14013;
assign w15939 = ~w16159 & w8671;
assign w15940 = ~w6362 & ~w2118;
assign w15941 = a_58 & w2249;
assign w15942 = w16188 & ~w17378;
assign w15943 = w627 & w14754;
assign w15944 = ~w6332 & ~w15388;
assign w15945 = w9547 & w15034;
assign w15946 = ~w8043 & ~w12593;
assign w15947 = ~w63 & w13497;
assign w15948 = ~w14295 & ~w814;
assign w15949 = ~w18186 & ~w6592;
assign w15950 = ~w9926 & ~w8073;
assign w15951 = ~w8905 & ~w1305;
assign w15952 = ~w1048 & ~w8921;
assign w15953 = ~w1493 & ~w4822;
assign w15954 = ~w11290 & ~w7319;
assign w15955 = ~w1093 & ~w3118;
assign w15956 = ~w5610 & ~w874;
assign w15957 = ~w11391 & w9130;
assign w15958 = a_21 & a_31;
assign w15959 = (~w1503 & w5270) | (~w1503 & w18238) | (w5270 & w18238);
assign w15960 = w10851 & ~w12512;
assign w15961 = ~w13377 & ~w13508;
assign w15962 = ~w8673 & w16222;
assign w15963 = (w17557 & w6208) | (w17557 & w13264) | (w6208 & w13264);
assign w15964 = w2529 & w2149;
assign w15965 = ~w1124 & ~w12777;
assign w15966 = ~w7066 & ~w18318;
assign w15967 = w5220 & w10187;
assign w15968 = w13428 & ~w11300;
assign w15969 = ~w11792 & w4577;
assign w15970 = (~w3264 & ~w582) | (~w3264 & w4728) | (~w582 & w4728);
assign w15971 = a_12 & a_51;
assign w15972 = ~w16394 & ~w3732;
assign w15973 = ~w8450 & ~w4482;
assign w15974 = w8651 & ~w2145;
assign w15975 = ~w12206 & ~w1581;
assign w15976 = a_32 & a_40;
assign w15977 = w17169 & ~w12853;
assign w15978 = w15598 & w1327;
assign w15979 = ~w13884 & ~w12820;
assign w15980 = w16162 & w14450;
assign w15981 = ~w17793 & w4295;
assign w15982 = w1850 & ~w7258;
assign w15983 = ~w3912 & ~w7534;
assign w15984 = ~w2261 & ~w10692;
assign w15985 = ~w10150 & ~w2469;
assign w15986 = ~w16916 & w2473;
assign w15987 = ~w14860 & ~w973;
assign w15988 = ~w10198 & w2429;
assign w15989 = w7447 & w11778;
assign w15990 = ~w11587 & ~w7804;
assign w15991 = ~w16788 & w15805;
assign w15992 = (~w922 & ~w2217) | (~w922 & w2371) | (~w2217 & w2371);
assign w15993 = ~w17555 & ~w2213;
assign w15994 = a_1 & a_34;
assign w15995 = ~w14309 & ~w13965;
assign w15996 = ~w14751 & ~w6965;
assign w15997 = ~w10351 & ~w12721;
assign w15998 = w5017 & ~w3351;
assign w15999 = w8777 & w9040;
assign w16000 = ~w4759 & ~w12913;
assign w16001 = ~w6229 & ~w1365;
assign w16002 = w4332 & w16218;
assign w16003 = ~w16563 & w1863;
assign w16004 = ~w12232 & ~w10474;
assign w16005 = w16018 & ~w2116;
assign w16006 = a_12 & a_37;
assign w16007 = ~w7636 & ~w3026;
assign w16008 = w14249 & ~w9339;
assign w16009 = ~w14333 & ~w5614;
assign w16010 = ~w10147 & ~w12463;
assign w16011 = w11061 & w3185;
assign w16012 = ~w6523 & ~w17391;
assign w16013 = ~w6628 & w2611;
assign w16014 = ~w13831 & ~w8018;
assign w16015 = w1507 & ~w11550;
assign w16016 = ~w938 & ~w10929;
assign w16017 = ~w3543 & ~w1883;
assign w16018 = ~w18818 & ~w3808;
assign w16019 = w734 & ~w17050;
assign w16020 = ~w14101 & w18616;
assign w16021 = w17701 & w13033;
assign w16022 = ~w2016 & ~w19068;
assign w16023 = ~w2828 & ~w13393;
assign w16024 = w13958 & w5462;
assign w16025 = w18128 & w19188;
assign w16026 = ~w7043 & ~w12054;
assign w16027 = ~w6019 & w9773;
assign w16028 = ~w15639 & ~w816;
assign w16029 = ~w6665 & ~w8035;
assign w16030 = ~w11062 & ~w18157;
assign w16031 = ~w1505 & ~w3301;
assign w16032 = a_3 & a_11;
assign w16033 = (~w11958 & w5527) | (~w11958 & w3247) | (w5527 & w3247);
assign w16034 = ~w18951 & ~w2953;
assign w16035 = a_4 & a_58;
assign w16036 = a_53 & a_56;
assign w16037 = ~w9742 & w10659;
assign w16038 = ~w12410 & ~w453;
assign w16039 = (~w17964 & ~w1568) | (~w17964 & w15379) | (~w1568 & w15379);
assign w16040 = w1679 & ~w4251;
assign w16041 = ~w10615 & ~w19174;
assign w16042 = w8318 & ~w15638;
assign w16043 = w16699 & w16596;
assign w16044 = ~w9403 & ~w3412;
assign w16045 = (w15061 & w5527) | (w15061 & w561) | (w5527 & w561);
assign w16046 = ~w8306 & ~w16407;
assign w16047 = ~w3961 & ~w19025;
assign w16048 = w2308 & w15291;
assign w16049 = ~w2861 & w9820;
assign w16050 = ~w13592 & ~w14493;
assign w16051 = ~w7293 & ~w11033;
assign w16052 = ~w12755 & ~w1149;
assign w16053 = ~w17643 & w8251;
assign w16054 = ~w6506 & ~w3312;
assign w16055 = a_9 & a_37;
assign w16056 = ~w18714 & ~w14027;
assign w16057 = ~w14745 & ~w19014;
assign w16058 = ~w7246 & w2657;
assign w16059 = w13829 & ~w17276;
assign w16060 = (w18357 & w12669) | (w18357 & w2474) | (w12669 & w2474);
assign w16061 = ~w9802 & w14819;
assign w16062 = (~w999 & w7863) | (~w999 & w9550) | (w7863 & w9550);
assign w16063 = w10234 & w11601;
assign w16064 = w12560 & ~w17383;
assign w16065 = w4692 & ~w2810;
assign w16066 = ~w8234 & ~w7027;
assign w16067 = w15726 & ~w16708;
assign w16068 = ~w14516 & ~w7711;
assign w16069 = a_25 & a_46;
assign w16070 = ~w954 & ~w12471;
assign w16071 = ~w1098 & ~w19067;
assign w16072 = ~w15311 & ~w10890;
assign w16073 = w3230 & ~w4511;
assign w16074 = ~w5839 & ~w455;
assign w16075 = ~w10542 & w1311;
assign w16076 = w17335 & w4222;
assign w16077 = w13971 & w13020;
assign w16078 = ~w15582 & ~w686;
assign w16079 = (w1524 & w12846) | (w1524 & w7729) | (w12846 & w7729);
assign w16080 = ~w11006 & ~w4507;
assign w16081 = w6519 & w15422;
assign w16082 = ~w4347 & ~w4797;
assign w16083 = ~w18260 & ~w5128;
assign w16084 = ~w4421 & ~w15246;
assign w16085 = ~w16946 & ~w5295;
assign w16086 = (w375 & w16269) | (w375 & w13327) | (w16269 & w13327);
assign w16087 = ~w4659 & ~w17386;
assign w16088 = w14713 & w18095;
assign w16089 = ~w7404 & ~w3581;
assign w16090 = w3116 & w2951;
assign w16091 = w5144 & w1051;
assign w16092 = w18943 & ~w17462;
assign w16093 = ~w7812 & ~w5561;
assign w16094 = ~w2590 & ~w13956;
assign w16095 = a_26 & a_46;
assign w16096 = ~w4219 & w11527;
assign w16097 = ~w7571 & ~w18013;
assign w16098 = a_3 & a_4;
assign w16099 = ~w19016 & ~w14821;
assign w16100 = ~w1838 & ~w13263;
assign w16101 = ~w6102 & w11653;
assign w16102 = ~w18020 & ~w13611;
assign w16103 = w8380 & w14788;
assign w16104 = a_43 & a_56;
assign w16105 = ~w11309 & ~w15501;
assign w16106 = ~w753 & ~w18183;
assign w16107 = w16095 & ~w11084;
assign w16108 = ~w6786 & ~w9435;
assign w16109 = ~w2739 & ~w18291;
assign w16110 = a_2 & a_57;
assign w16111 = ~w12687 & ~w4632;
assign w16112 = ~w3000 & ~w3597;
assign w16113 = ~w2769 & w3019;
assign w16114 = w3152 & w678;
assign w16115 = ~w6226 & w14800;
assign w16116 = a_59 & a_60;
assign w16117 = ~w6764 & ~w2656;
assign w16118 = ~w13754 & ~w8071;
assign w16119 = (w15415 & w10553) | (w15415 & w711) | (w10553 & w711);
assign w16120 = ~w18356 & ~w10312;
assign w16121 = ~w15410 & ~w17202;
assign w16122 = a_8 & a_60;
assign w16123 = w12803 & w13109;
assign w16124 = ~w7496 & ~w11431;
assign w16125 = ~w6985 & w2675;
assign w16126 = ~w14667 & ~w8070;
assign w16127 = ~w1460 & ~w679;
assign w16128 = ~w12651 & ~w2788;
assign w16129 = ~w3616 & ~w18424;
assign w16130 = w14930 & ~w6321;
assign w16131 = a_16 & a_53;
assign w16132 = ~w9777 & ~w16037;
assign w16133 = w9461 & ~w262;
assign w16134 = ~w6444 & ~w9195;
assign w16135 = ~w13812 & ~w14114;
assign w16136 = (w7604 & w8052) | (w7604 & w11914) | (w8052 & w11914);
assign w16137 = ~w3492 & w18561;
assign w16138 = w16891 & w1375;
assign w16139 = ~w1063 & w16460;
assign w16140 = w8824 & w12304;
assign w16141 = ~w16590 & w12279;
assign w16142 = (~w1696 & ~w15715) | (~w1696 & w18439) | (~w15715 & w18439);
assign w16143 = ~w12372 & ~w18801;
assign w16144 = (~w10834 & ~w15901) | (~w10834 & w10439) | (~w15901 & w10439);
assign w16145 = (~w8195 & ~w7446) | (~w8195 & w5117) | (~w7446 & w5117);
assign w16146 = ~w15377 & ~w3575;
assign w16147 = ~w963 & w4067;
assign w16148 = w15160 & w18610;
assign w16149 = w8369 & ~w6696;
assign w16150 = ~w4615 & ~w9424;
assign w16151 = ~w17990 & ~w2003;
assign w16152 = ~w18335 & ~w7197;
assign w16153 = ~w4609 & ~w6058;
assign w16154 = ~w3327 & ~w11681;
assign w16155 = ~w10699 & ~w8294;
assign w16156 = w17928 & w12251;
assign w16157 = w10254 & w15036;
assign w16158 = ~w6111 & w19049;
assign w16159 = w9980 & w15848;
assign w16160 = ~w9117 & ~w12735;
assign w16161 = ~w9518 & ~w2542;
assign w16162 = ~w15233 & ~w17244;
assign w16163 = ~w17409 & ~w4801;
assign w16164 = w10697 & w8240;
assign w16165 = w7912 & w1767;
assign w16166 = a_2 & a_27;
assign w16167 = w13752 & w9068;
assign w16168 = ~w16193 & ~w10775;
assign w16169 = w10234 & ~w13957;
assign w16170 = w10119 & ~w13959;
assign w16171 = ~w5582 & ~w16827;
assign w16172 = a_35 & a_59;
assign w16173 = w2758 & ~w6848;
assign w16174 = ~w15264 & w2524;
assign w16175 = (w9337 & w17297) | (w9337 & w778) | (w17297 & w778);
assign w16176 = w7456 & ~w12363;
assign w16177 = w8504 & ~w10599;
assign w16178 = ~w5942 & ~w14514;
assign w16179 = ~w13151 & ~w5178;
assign w16180 = w13153 & w17650;
assign w16181 = w3629 & w9728;
assign w16182 = ~w3030 & ~w6591;
assign w16183 = ~w10591 & w3672;
assign w16184 = ~w636 & ~w7964;
assign w16185 = (w8618 & w13275) | (w8618 & w4625) | (w13275 & w4625);
assign w16186 = a_13 & a_44;
assign w16187 = a_34 & a_52;
assign w16188 = ~w16360 & ~w8739;
assign w16189 = ~w1387 & ~w12808;
assign w16190 = ~w7576 & ~w2977;
assign w16191 = w15544 & w4349;
assign w16192 = ~w1307 & ~w6460;
assign w16193 = w15344 & w18166;
assign w16194 = ~w9692 & w894;
assign w16195 = ~w1274 & ~w18851;
assign w16196 = ~w413 & w19189;
assign w16197 = w2448 & ~w17474;
assign w16198 = ~w3108 & ~w18225;
assign w16199 = (~w18069 & ~w13513) | (~w18069 & w8959) | (~w13513 & w8959);
assign w16200 = ~w11404 & ~w6093;
assign w16201 = a_6 & w7098;
assign w16202 = ~w19004 & w4364;
assign w16203 = ~w13610 & ~w979;
assign w16204 = ~w6153 & ~w9228;
assign w16205 = w16174 & ~w19116;
assign w16206 = (~w7378 & ~w12558) | (~w7378 & w18542) | (~w12558 & w18542);
assign w16207 = w2089 & ~w483;
assign w16208 = ~w13172 & ~w16411;
assign w16209 = ~w12226 & ~w4569;
assign w16210 = ~w4025 & ~w6018;
assign w16211 = ~w11942 & ~w16807;
assign w16212 = ~w17684 & ~w19039;
assign w16213 = ~w13308 & ~w158;
assign w16214 = ~w7164 & ~w11468;
assign w16215 = ~w9774 & ~w6964;
assign w16216 = w3189 & w15150;
assign w16217 = (~w4979 & w16399) | (~w4979 & w1165) | (w16399 & w1165);
assign w16218 = ~w9565 & ~w13751;
assign w16219 = ~w16251 & ~w6771;
assign w16220 = ~w16040 & ~w9024;
assign w16221 = ~w9300 & w12542;
assign w16222 = ~w9018 & ~w751;
assign w16223 = ~w6671 & ~w8093;
assign w16224 = ~w779 & ~w1024;
assign w16225 = ~w2142 & w17874;
assign w16226 = ~w15974 & ~w8386;
assign w16227 = ~w10255 & ~w13099;
assign w16228 = a_24 & a_41;
assign w16229 = a_3 & a_13;
assign w16230 = a_9 & a_54;
assign w16231 = (~w428 & ~w1448) | (~w428 & w14226) | (~w1448 & w14226);
assign w16232 = a_30 & a_53;
assign w16233 = a_18 & a_59;
assign w16234 = ~w5856 & ~w42;
assign w16235 = ~w17718 & w11247;
assign w16236 = (~w15050 & w2150) | (~w15050 & w1104) | (w2150 & w1104);
assign w16237 = ~w6784 & ~w5314;
assign w16238 = ~w4697 & ~w1377;
assign w16239 = ~w4812 & ~w6925;
assign w16240 = ~w3725 & ~w17760;
assign w16241 = ~w6249 & w17352;
assign w16242 = ~w6653 & w13071;
assign w16243 = ~w10302 & ~w8759;
assign w16244 = ~w3770 & w1570;
assign w16245 = ~w3659 & ~w19117;
assign w16246 = a_23 & a_56;
assign w16247 = (~w900 & ~w4009) | (~w900 & w3317) | (~w4009 & w3317);
assign w16248 = (~w3630 & ~w18831) | (~w3630 & w1241) | (~w18831 & w1241);
assign w16249 = (~w19034 & ~w17031) | (~w19034 & w11433) | (~w17031 & w11433);
assign w16250 = a_36 & a_51;
assign w16251 = ~w17735 & ~w1860;
assign w16252 = a_25 & a_31;
assign w16253 = w13290 & ~w9962;
assign w16254 = a_30 & a_57;
assign w16255 = ~w6006 & ~w13815;
assign w16256 = ~w7086 & ~w1838;
assign w16257 = ~w7929 & w13171;
assign w16258 = w3592 & ~w1380;
assign w16259 = ~w4679 & ~w17427;
assign w16260 = w5692 & w6549;
assign w16261 = ~w9144 & ~w11986;
assign w16262 = a_30 & a_37;
assign w16263 = ~w16001 & ~w9017;
assign w16264 = ~w1567 & ~w8802;
assign w16265 = ~w5422 & ~w8583;
assign w16266 = ~w11292 & ~w8019;
assign w16267 = ~w11031 & ~w10554;
assign w16268 = w2583 & ~w2414;
assign w16269 = ~w2330 & w11312;
assign w16270 = (~w9620 & ~w17102) | (~w9620 & w15217) | (~w17102 & w15217);
assign w16271 = ~w5637 & ~w4928;
assign w16272 = ~w963 & w12394;
assign w16273 = a_10 & a_51;
assign w16274 = ~w16636 & ~w6989;
assign w16275 = ~w8332 & ~w14050;
assign w16276 = ~a_20 & ~w5914;
assign w16277 = a_6 & a_39;
assign w16278 = (~w494 & ~w7250) | (~w494 & w1293) | (~w7250 & w1293);
assign w16279 = w12229 & ~w4102;
assign w16280 = a_46 & w17557;
assign w16281 = ~w10532 & w8883;
assign w16282 = w3109 & w16444;
assign w16283 = ~w397 & ~w9233;
assign w16284 = ~w6065 & w5441;
assign w16285 = w6237 & ~w7458;
assign w16286 = ~w3803 & ~w9838;
assign w16287 = a_10 & a_53;
assign w16288 = ~w9410 & ~w18370;
assign w16289 = ~w914 & w10292;
assign w16290 = w17502 & ~w7664;
assign w16291 = w2870 & ~w13979;
assign w16292 = (~w15300 & ~w11133) | (~w15300 & w15631) | (~w11133 & w15631);
assign w16293 = ~w16996 & ~w12829;
assign w16294 = w4567 & ~w381;
assign w16295 = ~w3721 & ~w6842;
assign w16296 = (~w16555 & ~w309) | (~w16555 & w18138) | (~w309 & w18138);
assign w16297 = w7295 & ~w6243;
assign w16298 = ~a_11 & ~w10055;
assign w16299 = a_9 & a_26;
assign w16300 = ~w17028 & w18461;
assign w16301 = ~w2227 & w15499;
assign w16302 = ~w12343 & w14417;
assign w16303 = ~w4995 & ~w18800;
assign w16304 = ~w3846 & ~w5459;
assign w16305 = (w10445 & w13082) | (w10445 & w16797) | (w13082 & w16797);
assign w16306 = ~w11021 & w6072;
assign w16307 = ~w201 & w11588;
assign w16308 = ~w12105 & ~w3074;
assign w16309 = w14506 & w4020;
assign w16310 = w285 & ~w12757;
assign w16311 = a_0 & a_17;
assign w16312 = ~w1906 & w19190;
assign w16313 = ~w17610 & ~w18368;
assign w16314 = a_15 & a_53;
assign w16315 = a_20 & a_47;
assign w16316 = w1253 & ~w12315;
assign w16317 = ~w13661 & ~w1153;
assign w16318 = ~w18756 & ~w7637;
assign w16319 = w2260 & w13922;
assign w16320 = a_5 & a_17;
assign w16321 = ~w3996 & ~w17404;
assign w16322 = ~w3930 & ~w11906;
assign w16323 = ~w12994 & ~w7720;
assign w16324 = ~w2127 & ~w7107;
assign w16325 = w15009 & w12267;
assign w16326 = w7205 & w4267;
assign w16327 = ~w11725 & ~w11343;
assign w16328 = ~w17406 & ~w6690;
assign w16329 = w12693 & ~w18864;
assign w16330 = w1099 & ~w8543;
assign w16331 = a_5 & w12021;
assign w16332 = ~w17232 & ~w12518;
assign w16333 = (~w13616 & ~w2123) | (~w13616 & w11793) | (~w2123 & w11793);
assign w16334 = w13082 & w13160;
assign w16335 = ~w6182 & ~w11741;
assign w16336 = w916 & ~w17241;
assign w16337 = w5837 & w12733;
assign w16338 = ~w19066 & ~w6126;
assign w16339 = w12256 & w3506;
assign w16340 = ~w12900 & ~w19017;
assign w16341 = ~w1631 & ~w8297;
assign w16342 = w5337 & w8928;
assign w16343 = ~w9116 & ~w12860;
assign w16344 = ~w12975 & ~w15740;
assign w16345 = w6487 & w7419;
assign w16346 = ~w11626 & ~w14177;
assign w16347 = a_19 & a_23;
assign w16348 = ~w7085 & ~w12451;
assign w16349 = ~w18552 & ~w700;
assign w16350 = ~w11517 & ~w2999;
assign w16351 = ~w5102 & w10362;
assign w16352 = w434 & w6110;
assign w16353 = ~w9402 & ~w15906;
assign w16354 = w5870 & w13202;
assign w16355 = w7430 & ~w4580;
assign w16356 = ~w7177 & w240;
assign w16357 = a_16 & a_25;
assign w16358 = ~w14530 & ~w14648;
assign w16359 = (~w18365 & w10070) | (~w18365 & w9617) | (w10070 & w9617);
assign w16360 = ~w5739 & ~w308;
assign w16361 = ~w10036 & ~w2901;
assign w16362 = (~w17495 & ~w6285) | (~w17495 & w19135) | (~w6285 & w19135);
assign w16363 = a_25 & a_48;
assign w16364 = w429 & ~w13580;
assign w16365 = w12960 & ~w5333;
assign w16366 = ~w8156 & ~w15517;
assign w16367 = w8793 & ~w12444;
assign w16368 = ~w13545 & w3153;
assign w16369 = w14167 & ~w16729;
assign w16370 = ~w13646 & ~w1411;
assign w16371 = ~w12531 & ~w2829;
assign w16372 = a_6 & a_35;
assign w16373 = ~w10679 & ~w5752;
assign w16374 = ~w10858 & ~w4448;
assign w16375 = w16174 & w14480;
assign w16376 = w4089 & ~w8437;
assign w16377 = ~w10772 & ~w10323;
assign w16378 = w6398 & w14852;
assign w16379 = a_16 & w2249;
assign w16380 = ~w10859 & ~w17560;
assign w16381 = w17814 & ~w11037;
assign w16382 = ~w12337 & ~w12539;
assign w16383 = w1845 & w19099;
assign w16384 = ~w3207 & ~w16809;
assign w16385 = ~w7013 & ~w12548;
assign w16386 = ~w1785 & ~w6757;
assign w16387 = ~w2874 & ~w9606;
assign w16388 = ~w13737 & ~w19013;
assign w16389 = a_13 & a_51;
assign w16390 = ~w14254 & ~w5179;
assign w16391 = ~w8925 & ~w18991;
assign w16392 = w15000 & w18297;
assign w16393 = w4421 & ~w18878;
assign w16394 = ~w2545 & ~w114;
assign w16395 = ~w3305 & ~w9295;
assign w16396 = ~w4408 & ~w10136;
assign w16397 = ~w11212 & ~w9363;
assign w16398 = a_50 & a_57;
assign w16399 = ~w2769 & w8933;
assign w16400 = w11457 & w9665;
assign w16401 = ~w9058 & w13400;
assign w16402 = ~w8399 & ~w3410;
assign w16403 = w7594 & w14787;
assign w16404 = ~w12295 & w2835;
assign w16405 = (~w4021 & ~w18837) | (~w4021 & w3656) | (~w18837 & w3656);
assign w16406 = ~w7652 & ~w8877;
assign w16407 = w14254 & w5179;
assign w16408 = ~w15646 & ~w11693;
assign w16409 = ~w9019 & ~w15490;
assign w16410 = (~w896 & ~w10257) | (~w896 & w8916) | (~w10257 & w8916);
assign w16411 = ~w6138 & ~w12215;
assign w16412 = ~w10162 & ~w3007;
assign w16413 = a_24 & a_37;
assign w16414 = ~w11392 & ~w9194;
assign w16415 = ~w97 & w9003;
assign w16416 = ~w4637 & ~w12006;
assign w16417 = ~w6412 & ~w9991;
assign w16418 = ~w7232 & ~w5301;
assign w16419 = ~w17182 & ~w8177;
assign w16420 = ~w18696 & ~w17877;
assign w16421 = (~w2369 & ~w11495) | (~w2369 & w7391) | (~w11495 & w7391);
assign w16422 = a_17 & a_61;
assign w16423 = ~w11631 & ~w11529;
assign w16424 = ~w255 & ~w10863;
assign w16425 = w11547 & ~w11075;
assign w16426 = ~w4184 & ~w4666;
assign w16427 = a_5 & a_10;
assign w16428 = w413 & ~w10544;
assign w16429 = w16214 & w17094;
assign w16430 = w9574 & ~w6265;
assign w16431 = ~w9079 & w10061;
assign w16432 = (~w12487 & w464) | (~w12487 & w13093) | (w464 & w13093);
assign w16433 = ~w5343 & ~w479;
assign w16434 = (~w5909 & ~w2537) | (~w5909 & w8605) | (~w2537 & w8605);
assign w16435 = w17061 & w967;
assign w16436 = ~w7988 & ~w7405;
assign w16437 = (w18128 & w5882) | (w18128 & w15755) | (w5882 & w15755);
assign w16438 = ~a_7 & ~w14475;
assign w16439 = ~w10169 & ~w9878;
assign w16440 = ~w85 & ~w15950;
assign w16441 = ~w18440 & ~w172;
assign w16442 = w7711 & ~w5320;
assign w16443 = ~w1336 & w16508;
assign w16444 = ~w12265 & ~w17318;
assign w16445 = (~w17779 & ~w5492) | (~w17779 & w8276) | (~w5492 & w8276);
assign w16446 = w6903 & w12886;
assign w16447 = (~w1579 & ~w12664) | (~w1579 & w13725) | (~w12664 & w13725);
assign w16448 = ~w11583 & w13555;
assign w16449 = ~w5558 & ~w9904;
assign w16450 = w11662 & ~w14261;
assign w16451 = ~w1594 & w15287;
assign w16452 = w11316 & ~w4081;
assign w16453 = w1061 & ~w6650;
assign w16454 = ~w4404 & ~w4825;
assign w16455 = w7412 & ~w1433;
assign w16456 = ~w321 & w6622;
assign w16457 = ~w10291 & ~w13271;
assign w16458 = w18866 & w13989;
assign w16459 = w16517 & ~w5787;
assign w16460 = ~w10710 & ~w18691;
assign w16461 = ~w13597 & w12626;
assign w16462 = ~w17122 & ~w3563;
assign w16463 = ~w9649 & w3411;
assign w16464 = w1834 & ~w18863;
assign w16465 = ~w15194 & ~w16717;
assign w16466 = ~w9155 & w7438;
assign w16467 = ~w14447 & ~w1551;
assign w16468 = ~w17128 & ~w837;
assign w16469 = w17960 & ~w2067;
assign w16470 = w9570 & ~w7687;
assign w16471 = ~w2111 & ~w11404;
assign w16472 = w11374 & w17886;
assign w16473 = ~w18165 & ~w11341;
assign w16474 = ~w6092 & ~w9536;
assign w16475 = a_10 & a_29;
assign w16476 = ~w15445 & ~w13925;
assign w16477 = (a_41 & w7435) | (a_41 & w11191) | (w7435 & w11191);
assign w16478 = ~w6789 & ~w2106;
assign w16479 = ~w6482 & ~w9416;
assign w16480 = w7594 & w13288;
assign w16481 = ~w366 & ~w3565;
assign w16482 = ~w10990 & ~w11382;
assign w16483 = ~w12660 & ~w7021;
assign w16484 = ~w4804 & w13287;
assign w16485 = ~w3298 & ~w11625;
assign w16486 = ~w5072 & ~w16925;
assign w16487 = w16379 & ~w1732;
assign w16488 = ~w18533 & ~w14955;
assign w16489 = a_24 & a_51;
assign w16490 = w15821 & w9456;
assign w16491 = ~w14973 & ~w16796;
assign w16492 = ~w13428 & w11300;
assign w16493 = ~w8871 & w2699;
assign w16494 = ~w3980 & ~w14865;
assign w16495 = a_14 & a_26;
assign w16496 = ~w11540 & ~w12857;
assign w16497 = ~w11922 & ~w16975;
assign w16498 = a_36 & a_49;
assign w16499 = ~w12717 & ~w4756;
assign w16500 = ~w3452 & w2521;
assign w16501 = w7747 & ~w19006;
assign w16502 = w14899 & w7146;
assign w16503 = a_23 & a_58;
assign w16504 = ~w12228 & ~w16902;
assign w16505 = a_22 & a_49;
assign w16506 = ~w13062 & ~w14293;
assign w16507 = ~w6266 & w3100;
assign w16508 = ~w16009 & ~w3140;
assign w16509 = ~w3955 & ~w16847;
assign w16510 = ~w17645 & w13293;
assign w16511 = w833 & ~w15474;
assign w16512 = a_24 & a_45;
assign w16513 = w5051 & w3943;
assign w16514 = a_0 & a_57;
assign w16515 = w347 & ~w16445;
assign w16516 = w3410 & w1809;
assign w16517 = ~w14899 & ~w7146;
assign w16518 = ~w9513 & w5261;
assign w16519 = w5176 & ~w12346;
assign w16520 = ~w6939 & ~w14570;
assign w16521 = w12737 & w10358;
assign w16522 = w13706 & ~w17101;
assign w16523 = ~w16903 & ~w10485;
assign w16524 = w11552 & ~w10003;
assign w16525 = ~w2074 & ~w7011;
assign w16526 = w9524 & w3455;
assign w16527 = ~w4472 & ~w18414;
assign w16528 = w6275 & w153;
assign w16529 = a_27 & a_48;
assign w16530 = ~w11269 & ~w12141;
assign w16531 = w3433 & w5089;
assign w16532 = ~w9219 & ~w14390;
assign w16533 = a_14 & a_39;
assign w16534 = ~w4105 & w4546;
assign w16535 = w1041 & ~w6446;
assign w16536 = ~w16229 & ~w2516;
assign w16537 = ~w6257 & ~w1569;
assign w16538 = ~w3936 & ~w11158;
assign w16539 = w1054 & ~w11730;
assign w16540 = w10428 & w14603;
assign w16541 = ~w17909 & w16970;
assign w16542 = ~a_1 & ~a_2;
assign w16543 = ~w5214 & w14259;
assign w16544 = ~w11873 & ~w11665;
assign w16545 = w19143 & w17001;
assign w16546 = a_31 & a_42;
assign w16547 = ~w13255 & ~w15065;
assign w16548 = ~w19036 & w10571;
assign w16549 = ~w6127 & w15111;
assign w16550 = ~w18755 & ~w15972;
assign w16551 = ~w8324 & ~w16845;
assign w16552 = w11392 & w9194;
assign w16553 = w1750 & ~w11835;
assign w16554 = ~w7660 & ~w14552;
assign w16555 = w18124 & w11635;
assign w16556 = w18494 & w8299;
assign w16557 = w8013 & ~w18076;
assign w16558 = ~w149 & ~w5986;
assign w16559 = w13818 & ~w3296;
assign w16560 = ~w17754 & ~w6196;
assign w16561 = (w1320 & w757) | (w1320 & w14858) | (w757 & w14858);
assign w16562 = a_7 & a_60;
assign w16563 = (~w15355 & ~w18244) | (~w15355 & w18060) | (~w18244 & w18060);
assign w16564 = (~w19028 & ~w11439) | (~w19028 & w17064) | (~w11439 & w17064);
assign w16565 = a_35 & a_62;
assign w16566 = ~w9122 & w14958;
assign w16567 = (~w9799 & w6857) | (~w9799 & w3293) | (w6857 & w3293);
assign w16568 = ~w6277 & w11531;
assign w16569 = a_42 & a_45;
assign w16570 = w14253 & ~w14347;
assign w16571 = (~w6502 & ~w11910) | (~w6502 & w18456) | (~w11910 & w18456);
assign w16572 = ~w10338 & ~w2188;
assign w16573 = w2287 & w12698;
assign w16574 = ~w419 & w8187;
assign w16575 = w3134 & ~w16142;
assign w16576 = ~w3216 & ~w8748;
assign w16577 = ~w16571 & ~w18217;
assign w16578 = ~w14450 & ~w15233;
assign w16579 = w2927 & ~w7718;
assign w16580 = ~w10890 & w2894;
assign w16581 = w12795 & ~w893;
assign w16582 = (a_39 & w5654) | (a_39 & w14103) | (w5654 & w14103);
assign w16583 = ~w11620 & ~w17547;
assign w16584 = w17282 & ~w2084;
assign w16585 = ~w9067 & ~w9351;
assign w16586 = ~w16570 & ~w3147;
assign w16587 = a_24 & a_49;
assign w16588 = w10291 & w13271;
assign w16589 = ~w2976 & w9833;
assign w16590 = ~w13762 & ~w12659;
assign w16591 = w3652 & w19095;
assign w16592 = w9368 & w1286;
assign w16593 = ~w8341 & w13060;
assign w16594 = ~w9458 & ~w7850;
assign w16595 = ~w15925 & ~w7222;
assign w16596 = a_7 & a_57;
assign w16597 = (~w16552 & ~w1202) | (~w16552 & w4174) | (~w1202 & w4174);
assign w16598 = ~w12485 & w5394;
assign w16599 = ~w17246 & ~w3867;
assign w16600 = ~w12221 & ~w8847;
assign w16601 = ~w18863 & ~w907;
assign w16602 = w7570 & w2855;
assign w16603 = ~w5888 & ~w6234;
assign w16604 = (~w18217 & ~w7256) | (~w18217 & w16577) | (~w7256 & w16577);
assign w16605 = w12219 & w5848;
assign w16606 = w16918 & w1225;
assign w16607 = ~w13678 & ~w5110;
assign w16608 = (~w18263 & ~w17600) | (~w18263 & w7000) | (~w17600 & w7000);
assign w16609 = ~w12924 & w11209;
assign w16610 = w9616 & ~w18544;
assign w16611 = ~w13041 & ~w2688;
assign w16612 = ~w8651 & w2145;
assign w16613 = ~w708 & ~w16167;
assign w16614 = ~w7567 & ~w10098;
assign w16615 = ~w1844 & w4519;
assign w16616 = w1246 & w11621;
assign w16617 = ~w13044 & ~w6809;
assign w16618 = (w4195 & w13082) | (w4195 & w1362) | (w13082 & w1362);
assign w16619 = ~w13278 & ~w11282;
assign w16620 = w9154 & ~w15845;
assign w16621 = ~w11785 & ~w13669;
assign w16622 = ~w14484 & ~w317;
assign w16623 = ~w16954 & ~w7543;
assign w16624 = ~w422 & ~w1650;
assign w16625 = w5097 & ~w289;
assign w16626 = a_42 & a_48;
assign w16627 = ~w577 & ~w14840;
assign w16628 = a_29 & a_61;
assign w16629 = ~w12873 & ~w3970;
assign w16630 = ~w14205 & ~w14448;
assign w16631 = ~w4663 & ~w10151;
assign w16632 = w1601 & ~w17859;
assign w16633 = w17593 & ~w13593;
assign w16634 = ~w11788 & w6962;
assign w16635 = ~w1480 & ~w4014;
assign w16636 = (~w12880 & ~w164) | (~w12880 & w5996) | (~w164 & w5996);
assign w16637 = ~w10289 & ~w4330;
assign w16638 = ~w12480 & ~w119;
assign w16639 = a_14 & a_61;
assign w16640 = a_32 & a_38;
assign w16641 = ~w15624 & w9447;
assign w16642 = ~w9373 & ~w7641;
assign w16643 = ~w17321 & ~w4264;
assign w16644 = w13909 & w4996;
assign w16645 = ~w16971 & ~w14590;
assign w16646 = ~w7897 & ~w18179;
assign w16647 = ~w14202 & ~w7997;
assign w16648 = ~w6182 & ~w5229;
assign w16649 = ~w18085 & w5698;
assign w16650 = ~w7793 & ~w10661;
assign w16651 = (~w3497 & ~w2604) | (~w3497 & w18746) | (~w2604 & w18746);
assign w16652 = ~w17258 & ~w3068;
assign w16653 = w5879 & w12623;
assign w16654 = w4412 & w9486;
assign w16655 = ~w13915 & ~w8226;
assign w16656 = ~w13869 & ~w11935;
assign w16657 = ~w19086 & ~w7586;
assign w16658 = ~w16381 & ~w14043;
assign w16659 = ~w6450 & ~w11928;
assign w16660 = w14462 & w12568;
assign w16661 = ~w3645 & w4075;
assign w16662 = ~w1092 & ~w18262;
assign w16663 = ~w12096 & ~w1872;
assign w16664 = ~w9782 & ~w16816;
assign w16665 = ~w3194 & w7699;
assign w16666 = w8974 & w4075;
assign w16667 = ~w11960 & w16648;
assign w16668 = ~w10634 & ~w4099;
assign w16669 = ~w9104 & ~w6697;
assign w16670 = ~w8473 & ~w13068;
assign w16671 = w1320 & w983;
assign w16672 = w5669 & w13881;
assign w16673 = a_12 & w15843;
assign w16674 = a_34 & a_45;
assign w16675 = a_34 & a_59;
assign w16676 = ~w18646 & w16058;
assign w16677 = a_40 & a_46;
assign w16678 = ~w12766 & ~w18353;
assign w16679 = ~w2564 & ~w17725;
assign w16680 = ~w9737 & ~w3895;
assign w16681 = ~w15635 & ~w3613;
assign w16682 = ~w14069 & w9103;
assign w16683 = ~w8884 & ~w9775;
assign w16684 = ~w5763 & ~w1853;
assign w16685 = ~w168 & ~w2050;
assign w16686 = w11939 & w15911;
assign w16687 = w11331 & w5707;
assign w16688 = ~w16342 & ~w15556;
assign w16689 = (w11252 & w13962) | (w11252 & w9302) | (w13962 & w9302);
assign w16690 = ~w227 & w1137;
assign w16691 = (w10727 & w1364) | (w10727 & w6440) | (w1364 & w6440);
assign w16692 = ~w5159 & ~w13878;
assign w16693 = ~w5906 & ~w17508;
assign w16694 = w7462 & ~w2977;
assign w16695 = ~w4342 & w14919;
assign w16696 = ~w15483 & ~w1704;
assign w16697 = ~w11132 & ~w9772;
assign w16698 = ~w10348 & ~w4131;
assign w16699 = a_17 & a_47;
assign w16700 = (w14161 & w1566) | (w14161 & w3608) | (w1566 & w3608);
assign w16701 = w16949 & ~w10319;
assign w16702 = w16247 & w9734;
assign w16703 = a_10 & a_16;
assign w16704 = ~w10701 & ~w873;
assign w16705 = w14830 & w12856;
assign w16706 = a_6 & a_53;
assign w16707 = w13864 & ~w5568;
assign w16708 = ~w17156 & ~w14327;
assign w16709 = ~w2960 & w6396;
assign w16710 = ~w7235 & w9902;
assign w16711 = w923 & w2136;
assign w16712 = a_27 & a_53;
assign w16713 = w13886 & w7422;
assign w16714 = ~w295 & ~w15105;
assign w16715 = ~w10330 & w17056;
assign w16716 = (w18718 & ~w1320) | (w18718 & w484) | (~w1320 & w484);
assign w16717 = a_60 & a_62;
assign w16718 = w6485 & w6368;
assign w16719 = ~w17982 & ~w12903;
assign w16720 = (w17022 & w2769) | (w17022 & w17320) | (w2769 & w17320);
assign w16721 = ~w4332 & ~w16218;
assign w16722 = w124 & w15346;
assign w16723 = ~w10354 & ~w7611;
assign w16724 = ~w11580 & w11640;
assign w16725 = ~w13683 & ~w18788;
assign w16726 = ~w491 & ~w16463;
assign w16727 = ~w6386 & ~w14483;
assign w16728 = ~w10103 & ~w9023;
assign w16729 = ~w11486 & ~w15317;
assign w16730 = ~w14014 & ~w8650;
assign w16731 = a_3 & a_17;
assign w16732 = (~w5191 & w18650) | (~w5191 & w14363) | (w18650 & w14363);
assign w16733 = w14746 & ~w14325;
assign w16734 = w17214 & ~w12320;
assign w16735 = w17149 & ~w36;
assign w16736 = (~w7432 & ~w17543) | (~w7432 & w3290) | (~w17543 & w3290);
assign w16737 = ~w2857 & w2275;
assign w16738 = a_4 & a_10;
assign w16739 = ~w13809 & ~w14203;
assign w16740 = ~w6318 & w13348;
assign w16741 = ~w10334 & ~w5373;
assign w16742 = (w18733 & w18239) | (w18733 & w619) | (w18239 & w619);
assign w16743 = ~w754 & ~w15315;
assign w16744 = ~w8317 & w3718;
assign w16745 = ~w703 & ~w1708;
assign w16746 = w694 & ~w3368;
assign w16747 = ~w15592 & ~w3643;
assign w16748 = w139 & ~w9718;
assign w16749 = ~w15919 & ~w15017;
assign w16750 = ~w6130 & ~w17066;
assign w16751 = w1667 & w9675;
assign w16752 = a_40 & a_53;
assign w16753 = a_53 & a_63;
assign w16754 = ~w6390 & ~w12359;
assign w16755 = (~w7124 & ~w6792) | (~w7124 & w16927) | (~w6792 & w16927);
assign w16756 = w11504 & ~w17713;
assign w16757 = ~w3975 & w9666;
assign w16758 = ~w13847 & ~w8902;
assign w16759 = (~w9337 & w17906) | (~w9337 & w17426) | (w17906 & w17426);
assign w16760 = a_5 & a_26;
assign w16761 = ~w11436 & ~w9290;
assign w16762 = ~w6140 & ~w1564;
assign w16763 = ~w760 & w2282;
assign w16764 = ~w4763 & ~w9850;
assign w16765 = (w6794 & w10330) | (w6794 & w11735) | (w10330 & w11735);
assign w16766 = ~w12576 & ~w7452;
assign w16767 = ~w9443 & ~w1900;
assign w16768 = ~w10011 & w16100;
assign w16769 = ~w4297 & ~w8400;
assign w16770 = ~w330 & w12092;
assign w16771 = ~w6341 & ~w3485;
assign w16772 = ~w11183 & ~w12401;
assign w16773 = ~w4280 & w4935;
assign w16774 = w3862 & ~w17442;
assign w16775 = w96 & w16315;
assign w16776 = ~w7790 & ~w11402;
assign w16777 = ~w9359 & ~w12590;
assign w16778 = ~w3924 & ~w8239;
assign w16779 = ~w15066 & ~w17127;
assign w16780 = w15902 & ~w7212;
assign w16781 = ~w2638 & ~w5701;
assign w16782 = a_13 & a_57;
assign w16783 = w9134 & ~w13110;
assign w16784 = w8043 & w12593;
assign w16785 = ~w17504 & ~w13104;
assign w16786 = w13887 & w17887;
assign w16787 = ~w16958 & ~w12535;
assign w16788 = ~w9860 & ~w5278;
assign w16789 = w10615 & w19191;
assign w16790 = a_33 & a_49;
assign w16791 = ~w5598 & ~w15447;
assign w16792 = a_46 & a_55;
assign w16793 = ~w17751 & ~w13573;
assign w16794 = ~w13354 & w251;
assign w16795 = w12612 & ~w16380;
assign w16796 = w12486 & w3758;
assign w16797 = ~w19005 & w10445;
assign w16798 = w13463 & w16477;
assign w16799 = ~w14508 & ~w5836;
assign w16800 = ~w4868 & ~w16921;
assign w16801 = ~w11283 & ~w12469;
assign w16802 = (w17711 & w10330) | (w17711 & w16815) | (w10330 & w16815);
assign w16803 = ~w6441 & w926;
assign w16804 = w16261 & ~w13570;
assign w16805 = ~w8198 & w11218;
assign w16806 = a_2 & a_15;
assign w16807 = ~w5195 & ~w12771;
assign w16808 = ~w16798 & ~w5584;
assign w16809 = ~w2185 & ~w12650;
assign w16810 = ~w3796 & w16419;
assign w16811 = ~w9540 & ~w6222;
assign w16812 = w8039 & ~w18719;
assign w16813 = ~w18224 & ~w439;
assign w16814 = ~w558 & ~w5013;
assign w16815 = (w17711 & w13082) | (w17711 & w11964) | (w13082 & w11964);
assign w16816 = w15674 & ~w4567;
assign w16817 = w7298 & ~w16776;
assign w16818 = ~w18501 & ~w6674;
assign w16819 = w16607 & ~w19112;
assign w16820 = ~w8163 & ~w15169;
assign w16821 = ~w9307 & w4664;
assign w16822 = w7639 & ~w8292;
assign w16823 = ~w8577 & ~w17430;
assign w16824 = w7838 & w16514;
assign w16825 = a_21 & a_42;
assign w16826 = ~w12835 & ~w9202;
assign w16827 = ~w3200 & ~w9771;
assign w16828 = w14299 & w7891;
assign w16829 = ~w8507 & w4949;
assign w16830 = ~w5505 & ~w5880;
assign w16831 = ~w14191 & ~w15131;
assign w16832 = ~w18287 & w6773;
assign w16833 = ~w11728 & w16635;
assign w16834 = ~w4099 & ~w3813;
assign w16835 = w15215 & w1381;
assign w16836 = a_20 & a_26;
assign w16837 = w2960 & ~w17326;
assign w16838 = ~w12609 & ~w4933;
assign w16839 = (w13018 & w19124) | (w13018 & w18017) | (w19124 & w18017);
assign w16840 = w9880 & w10945;
assign w16841 = ~w14464 & ~w6703;
assign w16842 = (w7102 & w15307) | (w7102 & w9296) | (w15307 & w9296);
assign w16843 = ~w13535 & ~w13539;
assign w16844 = w3878 & w4528;
assign w16845 = a_9 & a_41;
assign w16846 = ~w6934 & w2654;
assign w16847 = ~w15318 & ~w8812;
assign w16848 = a_47 & a_63;
assign w16849 = a_21 & a_63;
assign w16850 = ~w13065 & ~w9084;
assign w16851 = w10470 & ~w4718;
assign w16852 = ~w14572 & w4309;
assign w16853 = w13051 & ~w15546;
assign w16854 = ~w2174 & ~w4561;
assign w16855 = ~w434 & ~w6110;
assign w16856 = ~w14642 & ~w6575;
assign w16857 = ~w1845 & w7615;
assign w16858 = ~w3102 & ~w4866;
assign w16859 = a_36 & a_57;
assign w16860 = ~w15737 & w12153;
assign w16861 = ~w581 & w2659;
assign w16862 = w5897 & ~w8097;
assign w16863 = w13186 & ~w2541;
assign w16864 = w9697 & w18266;
assign w16865 = ~w9691 & w7072;
assign w16866 = w8236 & ~w10528;
assign w16867 = a_7 & a_54;
assign w16868 = a_3 & a_36;
assign w16869 = ~w15512 & ~w11113;
assign w16870 = ~w1354 & ~w15478;
assign w16871 = ~w15593 & w5726;
assign w16872 = w7705 & w7981;
assign w16873 = a_22 & a_43;
assign w16874 = ~w14613 & ~w15903;
assign w16875 = ~w675 & ~w799;
assign w16876 = ~w17758 & ~w7298;
assign w16877 = w2123 & ~w5063;
assign w16878 = ~w9277 & ~w5021;
assign w16879 = w5919 & w7732;
assign w16880 = (~w12255 & w11418) | (~w12255 & w18637) | (w11418 & w18637);
assign w16881 = w3763 & w8150;
assign w16882 = ~w12620 & ~w18210;
assign w16883 = ~w8374 & ~w17117;
assign w16884 = ~w685 & ~w1668;
assign w16885 = ~w5898 & ~w11663;
assign w16886 = ~w8824 & ~w12304;
assign w16887 = w3797 & ~w9443;
assign w16888 = (w11667 & w2769) | (w11667 & w664) | (w2769 & w664);
assign w16889 = ~w13150 & w666;
assign w16890 = ~w9614 & w18508;
assign w16891 = ~w15603 & ~w10649;
assign w16892 = ~w7825 & w14221;
assign w16893 = w7446 & ~w15867;
assign w16894 = w17809 & ~w5264;
assign w16895 = ~w12236 & ~w15872;
assign w16896 = w10803 & w14934;
assign w16897 = ~w15504 & w2949;
assign w16898 = a_0 & a_63;
assign w16899 = w2674 & ~w16617;
assign w16900 = a_28 & a_34;
assign w16901 = ~w12691 & w7749;
assign w16902 = ~w1983 & w5728;
assign w16903 = w9076 & ~w11162;
assign w16904 = (w6917 & w10330) | (w6917 & w303) | (w10330 & w303);
assign w16905 = w228 & w16441;
assign w16906 = ~w10072 & w3576;
assign w16907 = w4125 & ~w12892;
assign w16908 = ~w9569 & ~w3229;
assign w16909 = a_19 & a_22;
assign w16910 = w623 & ~w16409;
assign w16911 = w4904 & w52;
assign w16912 = ~w5137 & ~w4727;
assign w16913 = w1603 & w1651;
assign w16914 = ~w7595 & ~w16878;
assign w16915 = ~w4808 & ~w2461;
assign w16916 = ~w9177 & ~w11518;
assign w16917 = (~w11396 & w13422) | (~w11396 & w14273) | (w13422 & w14273);
assign w16918 = (~w12991 & ~w13232) | (~w12991 & w12505) | (~w13232 & w12505);
assign w16919 = w18375 & ~w388;
assign w16920 = ~w11731 & ~w11820;
assign w16921 = ~w15567 & w3365;
assign w16922 = ~w7868 & w13514;
assign w16923 = (a_50 & w11889) | (a_50 & w4315) | (w11889 & w4315);
assign w16924 = ~w16831 & ~w7555;
assign w16925 = ~w9155 & ~w11199;
assign w16926 = a_0 & a_51;
assign w16927 = ~w18236 & ~w7124;
assign w16928 = ~w16035 & ~w7869;
assign w16929 = ~w8146 & ~w13931;
assign w16930 = w17028 & ~w18461;
assign w16931 = a_27 & a_51;
assign w16932 = ~w7962 & ~w12524;
assign w16933 = ~w18027 & ~w9073;
assign w16934 = w10890 & ~w2894;
assign w16935 = ~w1026 & ~w5078;
assign w16936 = w8362 & ~w5048;
assign w16937 = ~w16469 & ~w8368;
assign w16938 = ~w18310 & ~w1232;
assign w16939 = w19098 & w15473;
assign w16940 = ~w18442 & w18109;
assign w16941 = ~w16201 & ~w15654;
assign w16942 = (w399 & w844) | (w399 & w4177) | (w844 & w4177);
assign w16943 = ~w3583 & w17370;
assign w16944 = w13324 & w17622;
assign w16945 = a_10 & a_49;
assign w16946 = w13736 & ~w7662;
assign w16947 = w13111 & ~w17084;
assign w16948 = a_11 & a_16;
assign w16949 = ~w4132 & ~w1383;
assign w16950 = ~w5239 & ~w14348;
assign w16951 = ~w8373 & ~w11214;
assign w16952 = w7601 & ~w17666;
assign w16953 = ~w13838 & ~w11690;
assign w16954 = a_2 & a_32;
assign w16955 = w11003 & ~w18181;
assign w16956 = w4211 & ~w13528;
assign w16957 = w9917 & w3267;
assign w16958 = ~w13494 & ~w15827;
assign w16959 = ~w3495 & ~w12993;
assign w16960 = ~w5683 & ~w12762;
assign w16961 = ~w14702 & ~w11721;
assign w16962 = ~w4749 & w14954;
assign w16963 = ~w17065 & w16762;
assign w16964 = ~w17311 & ~w18655;
assign w16965 = ~w5012 & ~w10769;
assign w16966 = ~w16486 & ~w7051;
assign w16967 = ~w12175 & ~w5616;
assign w16968 = ~w11893 & ~w2323;
assign w16969 = ~w2274 & ~w10200;
assign w16970 = ~w2057 & ~w8141;
assign w16971 = ~w14264 & ~w13490;
assign w16972 = ~w12330 & ~w9921;
assign w16973 = ~w8575 & ~w1931;
assign w16974 = ~w12562 & w16697;
assign w16975 = ~w18867 & ~w12712;
assign w16976 = w5797 & ~w10847;
assign w16977 = ~w11013 & ~w12928;
assign w16978 = ~w3122 & ~w17802;
assign w16979 = ~w16895 & ~w2638;
assign w16980 = ~w15274 & ~w15506;
assign w16981 = ~w5388 & ~w9788;
assign w16982 = ~w11857 & ~w10023;
assign w16983 = ~w16873 & ~w14330;
assign w16984 = (~w11421 & w5743) | (~w11421 & w19033) | (w5743 & w19033);
assign w16985 = ~w5797 & w10847;
assign w16986 = w17611 & ~w12534;
assign w16987 = ~w612 & ~w7746;
assign w16988 = a_12 & a_14;
assign w16989 = ~w13082 & w10293;
assign w16990 = w653 & ~w18965;
assign w16991 = ~w18740 & w16630;
assign w16992 = ~w9608 & ~w11184;
assign w16993 = ~w787 & ~w10089;
assign w16994 = (~w16521 & ~w18396) | (~w16521 & w13738) | (~w18396 & w13738);
assign w16995 = w1939 & w14255;
assign w16996 = w6363 & w14759;
assign w16997 = a_11 & w10055;
assign w16998 = (~w5290 & ~w14572) | (~w5290 & w17736) | (~w14572 & w17736);
assign w16999 = ~w1978 & ~w18089;
assign w17000 = ~w5512 & w5187;
assign w17001 = ~w7541 & ~w4672;
assign w17002 = ~w15972 & ~w18513;
assign w17003 = ~w10333 & ~w5185;
assign w17004 = ~w999 & ~w6402;
assign w17005 = w3396 & w12575;
assign w17006 = a_39 & a_40;
assign w17007 = w5009 & w1224;
assign w17008 = ~w15199 & w13163;
assign w17009 = ~w12032 & ~w13321;
assign w17010 = ~w14006 & ~w8285;
assign w17011 = ~w11044 & ~w15435;
assign w17012 = w10052 & w6560;
assign w17013 = ~w15724 & ~w5506;
assign w17014 = ~w1884 & ~w16473;
assign w17015 = a_8 & a_50;
assign w17016 = w6291 & ~w6834;
assign w17017 = (~w10566 & ~w12042) | (~w10566 & w17975) | (~w12042 & w17975);
assign w17018 = w6108 & ~w12582;
assign w17019 = a_16 & a_50;
assign w17020 = ~w12433 & ~w10115;
assign w17021 = ~w17425 & ~w14055;
assign w17022 = (w9025 & w10330) | (w9025 & w4258) | (w10330 & w4258);
assign w17023 = ~w17270 & ~w6515;
assign w17024 = ~w9535 & ~w16107;
assign w17025 = w16814 & w8789;
assign w17026 = ~w8057 & w513;
assign w17027 = ~w10487 & ~w18874;
assign w17028 = a_31 & a_52;
assign w17029 = ~w11637 & ~w6611;
assign w17030 = ~w11644 & w18455;
assign w17031 = ~w19034 & ~w4563;
assign w17032 = ~w17476 & w12828;
assign w17033 = ~w15005 & ~w10113;
assign w17034 = a_3 & a_19;
assign w17035 = ~w10704 & ~w11734;
assign w17036 = w13979 & w744;
assign w17037 = ~w17530 & ~w5581;
assign w17038 = w6811 & ~w13796;
assign w17039 = (w12904 & w8944) | (w12904 & w3345) | (w8944 & w3345);
assign w17040 = w2491 & w16981;
assign w17041 = (~w3745 & ~w18222) | (~w3745 & w5517) | (~w18222 & w5517);
assign w17042 = ~w14608 & w11802;
assign w17043 = w16153 & w18663;
assign w17044 = ~w6656 & ~w13232;
assign w17045 = ~w16494 & ~w9299;
assign w17046 = ~w5091 & ~w6720;
assign w17047 = a_62 & w11297;
assign w17048 = w16398 & ~w14288;
assign w17049 = ~w5978 & w17658;
assign w17050 = ~w8423 & ~w13730;
assign w17051 = ~w3059 & ~w8428;
assign w17052 = ~w3047 & ~w14104;
assign w17053 = w6915 & ~w1221;
assign w17054 = a_2 & a_18;
assign w17055 = ~w4535 & w5018;
assign w17056 = ~w13082 & w12201;
assign w17057 = ~w3397 & ~w10253;
assign w17058 = ~w11899 & ~w4427;
assign w17059 = ~w15074 & w4999;
assign w17060 = w9039 & ~w4198;
assign w17061 = ~w12653 & ~w2460;
assign w17062 = ~w575 & ~w8586;
assign w17063 = ~w14744 & ~w1555;
assign w17064 = w3904 & ~w19028;
assign w17065 = (~w7221 & ~w14772) | (~w7221 & w10434) | (~w14772 & w10434);
assign w17066 = ~w18350 & ~w11520;
assign w17067 = w3862 & ~w12985;
assign w17068 = ~w2226 & ~w15067;
assign w17069 = ~w9244 & ~w1239;
assign w17070 = w10907 & w1608;
assign w17071 = ~w13178 & w9234;
assign w17072 = ~w697 & w11328;
assign w17073 = ~w15113 & w18294;
assign w17074 = ~w4468 & ~w11151;
assign w17075 = w5629 & ~w4486;
assign w17076 = w12137 & ~w5821;
assign w17077 = w11333 & ~w11470;
assign w17078 = w4764 & w6419;
assign w17079 = ~w5386 & ~w11318;
assign w17080 = ~w728 & ~w11895;
assign w17081 = ~w11806 & ~w18079;
assign w17082 = ~w2924 & ~w1781;
assign w17083 = ~w11177 & w19064;
assign w17084 = ~w13529 & ~w17072;
assign w17085 = w5337 & ~w7387;
assign w17086 = ~w13849 & w14523;
assign w17087 = ~w2543 & ~w17940;
assign w17088 = ~w8927 & ~w9082;
assign w17089 = w13558 & w2352;
assign w17090 = ~w18244 & w4376;
assign w17091 = ~w1357 & ~w15876;
assign w17092 = ~w2959 & ~w3893;
assign w17093 = w17585 & ~w11849;
assign w17094 = ~w5065 & ~w7321;
assign w17095 = ~w12508 & w714;
assign w17096 = ~w4399 & ~w14536;
assign w17097 = a_32 & a_58;
assign w17098 = w11429 & ~w14027;
assign w17099 = ~w1410 & ~w16955;
assign w17100 = w13849 & ~w14523;
assign w17101 = ~w13089 & ~w8756;
assign w17102 = ~w9620 & ~w17073;
assign w17103 = ~w394 & ~w6716;
assign w17104 = ~w1653 & ~w8837;
assign w17105 = ~w9338 & ~w875;
assign w17106 = ~w17148 & ~w2677;
assign w17107 = w7961 & w1260;
assign w17108 = a_44 & a_53;
assign w17109 = a_9 & a_40;
assign w17110 = (~w14865 & ~w16494) | (~w14865 & w15220) | (~w16494 & w15220);
assign w17111 = (w14321 & w2517) | (w14321 & w189) | (w2517 & w189);
assign w17112 = a_8 & a_40;
assign w17113 = ~w18514 & ~w15214;
assign w17114 = ~w6541 & w1132;
assign w17115 = ~w18342 & ~w1272;
assign w17116 = a_20 & a_40;
assign w17117 = ~w4243 & ~w6747;
assign w17118 = ~w8303 & ~w17199;
assign w17119 = ~w11703 & ~w9169;
assign w17120 = ~w9293 & ~w15929;
assign w17121 = (~w8669 & ~w4798) | (~w8669 & w12914) | (~w4798 & w12914);
assign w17122 = (w14675 & w14509) | (w14675 & w9438) | (w14509 & w9438);
assign w17123 = a_7 & a_31;
assign w17124 = ~w8800 & w12214;
assign w17125 = ~w4286 & ~w12496;
assign w17126 = ~w17741 & ~w5485;
assign w17127 = w10459 & ~w11580;
assign w17128 = ~w11848 & ~w11022;
assign w17129 = w15483 & w1704;
assign w17130 = w4739 & ~w11322;
assign w17131 = w12594 & ~w731;
assign w17132 = w14221 & w10232;
assign w17133 = w6064 & w11413;
assign w17134 = w9120 & ~w16723;
assign w17135 = w12010 & ~w4864;
assign w17136 = ~w9395 & ~w8725;
assign w17137 = a_10 & a_26;
assign w17138 = ~w7909 & ~w17278;
assign w17139 = (~w18087 & ~w5191) | (~w18087 & w8533) | (~w5191 & w8533);
assign w17140 = w4776 & w10073;
assign w17141 = ~w979 & ~w17257;
assign w17142 = ~w7627 & ~w10901;
assign w17143 = ~w17588 & ~w17868;
assign w17144 = ~w3810 & w10684;
assign w17145 = ~w15868 & ~w18242;
assign w17146 = w12693 & ~w6700;
assign w17147 = ~w4909 & w9253;
assign w17148 = w5592 & ~w642;
assign w17149 = ~w17365 & ~w9930;
assign w17150 = a_11 & a_52;
assign w17151 = (w13979 & w17132) | (w13979 & w13898) | (w17132 & w13898);
assign w17152 = ~w11671 & ~w14908;
assign w17153 = ~w8462 & ~w4482;
assign w17154 = w6066 & w9356;
assign w17155 = w10723 & w10695;
assign w17156 = ~w18261 & ~w15636;
assign w17157 = ~w9277 & ~w3546;
assign w17158 = ~w15160 & ~w18610;
assign w17159 = w15108 & w1891;
assign w17160 = ~w11623 & w8761;
assign w17161 = a_45 & a_56;
assign w17162 = a_45 & a_53;
assign w17163 = ~w3971 & ~w15438;
assign w17164 = a_3 & a_58;
assign w17165 = w11126 & ~w9932;
assign w17166 = w7091 & w4368;
assign w17167 = ~w3781 & ~w5304;
assign w17168 = ~w4918 & w17703;
assign w17169 = ~w9294 & ~w12386;
assign w17170 = ~w818 & ~w12827;
assign w17171 = ~w16313 & w12211;
assign w17172 = ~w12063 & ~w13015;
assign w17173 = ~w8564 & w1658;
assign w17174 = ~w6299 & ~w782;
assign w17175 = w19055 & ~w4126;
assign w17176 = ~w4965 & w10444;
assign w17177 = ~w16695 & ~w17788;
assign w17178 = w5993 & w7337;
assign w17179 = ~w7160 & ~w3205;
assign w17180 = w18567 & w4987;
assign w17181 = ~w17827 & w15678;
assign w17182 = ~w7337 & ~w15320;
assign w17183 = ~w16085 & ~w2584;
assign w17184 = ~w4731 & ~w17880;
assign w17185 = ~w9472 & ~w9465;
assign w17186 = ~w16643 & ~w16353;
assign w17187 = ~w8145 & ~w6576;
assign w17188 = w14797 & w8863;
assign w17189 = ~w5491 & ~w16122;
assign w17190 = a_47 & a_48;
assign w17191 = ~w15763 & w4979;
assign w17192 = w5881 & w17111;
assign w17193 = ~w2163 & ~w790;
assign w17194 = ~w4390 & ~w4144;
assign w17195 = ~w15018 & ~w16262;
assign w17196 = (~w14415 & w16513) | (~w14415 & w657) | (w16513 & w657);
assign w17197 = ~w17216 & ~w14917;
assign w17198 = ~w203 & ~w6873;
assign w17199 = w12725 & w6736;
assign w17200 = w15492 & ~w9162;
assign w17201 = ~w13696 & ~w12792;
assign w17202 = ~w323 & w19075;
assign w17203 = ~w10615 & ~w19173;
assign w17204 = ~w14839 & ~w4090;
assign w17205 = w2220 & w18404;
assign w17206 = ~w12100 & w5967;
assign w17207 = ~w18017 & w10737;
assign w17208 = ~w525 & ~w12585;
assign w17209 = w16931 & ~w8289;
assign w17210 = w604 & w7238;
assign w17211 = ~w5086 & ~w18900;
assign w17212 = a_50 & a_62;
assign w17213 = w13615 & w12076;
assign w17214 = w8410 & ~w8515;
assign w17215 = ~w10581 & ~w13715;
assign w17216 = ~w3811 & w513;
assign w17217 = w9235 & w9653;
assign w17218 = a_48 & a_63;
assign w17219 = w12924 & ~w11209;
assign w17220 = ~w11460 & w17954;
assign w17221 = w13 & ~w5817;
assign w17222 = w4035 & ~w5834;
assign w17223 = ~w14896 & ~w15531;
assign w17224 = ~w16225 & ~w3371;
assign w17225 = w11689 & ~w14221;
assign w17226 = ~w8033 & ~w7121;
assign w17227 = a_15 & a_33;
assign w17228 = w17310 & w12312;
assign w17229 = ~w17753 & w8265;
assign w17230 = w3925 & ~w1434;
assign w17231 = ~w4983 & ~w302;
assign w17232 = ~w14517 & w6383;
assign w17233 = ~w2240 & w13070;
assign w17234 = (w2396 & w10330) | (w2396 & w14877) | (w10330 & w14877);
assign w17235 = ~w11097 & ~w11248;
assign w17236 = (~w11320 & ~w4541) | (~w11320 & w2205) | (~w4541 & w2205);
assign w17237 = a_37 & a_61;
assign w17238 = ~w15877 & w7299;
assign w17239 = (w5790 & w12446) | (w5790 & w3490) | (w12446 & w3490);
assign w17240 = w10139 & w14652;
assign w17241 = (~w13667 & ~w11623) | (~w13667 & w13451) | (~w11623 & w13451);
assign w17242 = ~w16275 & ~w9105;
assign w17243 = w18244 & ~w4376;
assign w17244 = ~w8633 & ~w5126;
assign w17245 = w3289 & ~w1554;
assign w17246 = a_45 & a_48;
assign w17247 = ~w286 & ~w13027;
assign w17248 = a_2 & a_40;
assign w17249 = ~w7892 & ~w12149;
assign w17250 = ~w17088 & ~w13292;
assign w17251 = ~w14241 & ~w10570;
assign w17252 = a_6 & a_61;
assign w17253 = (~w1069 & ~w8987) | (~w1069 & w10551) | (~w8987 & w10551);
assign w17254 = ~w3966 & w8096;
assign w17255 = ~w10080 & ~w8330;
assign w17256 = ~w7598 & ~w14947;
assign w17257 = w11483 & ~w13610;
assign w17258 = ~w4225 & ~w5490;
assign w17259 = ~w7012 & ~w8941;
assign w17260 = ~w13434 & w7108;
assign w17261 = ~w9827 & ~w11810;
assign w17262 = ~w15060 & w5811;
assign w17263 = w5680 & ~w4604;
assign w17264 = a_18 & a_57;
assign w17265 = w11537 & w3202;
assign w17266 = ~w9929 & w4110;
assign w17267 = w18904 & w4372;
assign w17268 = ~w379 & ~w9282;
assign w17269 = ~w18247 & w12599;
assign w17270 = ~w304 & ~w1331;
assign w17271 = ~w842 & w14008;
assign w17272 = ~w15474 & ~w3584;
assign w17273 = ~w16014 & ~w9453;
assign w17274 = ~w12554 & ~w5167;
assign w17275 = w2193 & w13587;
assign w17276 = ~w9868 & ~w7995;
assign w17277 = w3560 & ~w231;
assign w17278 = ~w13921 & ~w16530;
assign w17279 = ~w12572 & ~w7880;
assign w17280 = a_2 & a_28;
assign w17281 = w2005 & w12282;
assign w17282 = a_12 & a_50;
assign w17283 = a_39 & a_54;
assign w17284 = a_39 & a_58;
assign w17285 = a_8 & w19009;
assign w17286 = ~w17761 & ~w9212;
assign w17287 = (w13934 & w4477) | (w13934 & w1332) | (w4477 & w1332);
assign w17288 = ~w10789 & ~w9673;
assign w17289 = w5398 & ~w6547;
assign w17290 = w8843 & w8545;
assign w17291 = ~w14689 & ~w4985;
assign w17292 = (w16917 & w16606) | (w16917 & w7441) | (w16606 & w7441);
assign w17293 = w6736 & w10095;
assign w17294 = ~w11859 & ~w16515;
assign w17295 = ~w2422 & ~w9005;
assign w17296 = w11874 & w7080;
assign w17297 = w6396 & ~w1553;
assign w17298 = ~w3794 & ~w18398;
assign w17299 = ~w14132 & w9995;
assign w17300 = w13879 & ~w10784;
assign w17301 = ~w10169 & ~w6469;
assign w17302 = w8462 & w4482;
assign w17303 = w1908 & w16954;
assign w17304 = ~w16997 & ~w18498;
assign w17305 = ~w10709 & ~w2162;
assign w17306 = ~w16794 & ~w11176;
assign w17307 = (~w4150 & ~w8874) | (~w4150 & w9264) | (~w8874 & w9264);
assign w17308 = ~w16987 & ~w13208;
assign w17309 = ~w6269 & ~w14434;
assign w17310 = ~w16331 & ~w4771;
assign w17311 = ~w531 & ~w15301;
assign w17312 = ~w3180 & ~w1219;
assign w17313 = ~w929 & ~w5279;
assign w17314 = a_45 & a_52;
assign w17315 = w11545 & w14876;
assign w17316 = w11109 & w17631;
assign w17317 = ~w4430 & ~w12695;
assign w17318 = ~w18837 & w10419;
assign w17319 = w11696 & w10640;
assign w17320 = ~w6853 & w17022;
assign w17321 = w13267 & ~w8448;
assign w17322 = ~w8369 & w6696;
assign w17323 = ~w1286 & w11855;
assign w17324 = ~w9603 & w2306;
assign w17325 = w5758 & ~w18252;
assign w17326 = ~w861 & ~w17782;
assign w17327 = ~w16911 & ~w6333;
assign w17328 = w12997 & w7910;
assign w17329 = ~w12249 & ~w2441;
assign w17330 = w1158 & ~w4735;
assign w17331 = ~w1746 & ~w7138;
assign w17332 = w5795 & ~w18681;
assign w17333 = a_19 & a_36;
assign w17334 = ~w13521 & ~w2170;
assign w17335 = ~w8253 & ~w12672;
assign w17336 = ~w10214 & ~w5511;
assign w17337 = ~w11242 & ~w17180;
assign w17338 = ~w9999 & ~w16796;
assign w17339 = (~w9549 & ~w8747) | (~w9549 & w2936) | (~w8747 & w2936);
assign w17340 = ~w7357 & ~w4638;
assign w17341 = w104 & w5288;
assign w17342 = ~w4460 & ~w18029;
assign w17343 = w9141 & ~w16969;
assign w17344 = w11011 & w12967;
assign w17345 = ~w4148 & ~w8624;
assign w17346 = ~w16310 & ~w7285;
assign w17347 = ~w17071 & ~w9561;
assign w17348 = ~w14585 & ~w8226;
assign w17349 = ~w4106 & ~w14832;
assign w17350 = ~w11972 & w5714;
assign w17351 = ~w10428 & ~w18953;
assign w17352 = ~w7462 & ~w14233;
assign w17353 = (w10529 & w961) | (w10529 & w5882) | (w961 & w5882);
assign w17354 = ~w9142 & ~w1481;
assign w17355 = w10620 & ~w3881;
assign w17356 = w18781 & w13832;
assign w17357 = w12150 & ~w9326;
assign w17358 = ~w9485 & ~w5736;
assign w17359 = (~w12744 & ~w18203) | (~w12744 & w6867) | (~w18203 & w6867);
assign w17360 = ~w4697 & ~w1771;
assign w17361 = a_13 & a_28;
assign w17362 = ~w4317 & ~w16215;
assign w17363 = w16163 & ~w3783;
assign w17364 = w6267 & ~w6236;
assign w17365 = w13115 & w15028;
assign w17366 = ~w14248 & ~w4163;
assign w17367 = ~w10148 & ~w4741;
assign w17368 = ~w6327 & ~w5054;
assign w17369 = (~w5345 & ~w4278) | (~w5345 & w913) | (~w4278 & w913);
assign w17370 = ~w7500 & ~w1718;
assign w17371 = ~w11897 & w16017;
assign w17372 = w15264 & ~w11660;
assign w17373 = ~w14770 & w19032;
assign w17374 = ~w9236 & ~w4054;
assign w17375 = ~w11580 & ~w7373;
assign w17376 = ~w2753 & ~w8387;
assign w17377 = (w804 & w6416) | (w804 & w6853) | (w6416 & w6853);
assign w17378 = ~w15746 & ~w6379;
assign w17379 = a_21 & a_62;
assign w17380 = ~w11409 & ~w15497;
assign w17381 = ~w13060 & ~w14628;
assign w17382 = ~w16346 & ~w18554;
assign w17383 = ~w8565 & ~w7744;
assign w17384 = w8098 & w5720;
assign w17385 = ~w18398 & ~w7019;
assign w17386 = w16931 & ~w11314;
assign w17387 = ~w14602 & w18716;
assign w17388 = w2963 & ~w17533;
assign w17389 = ~w7363 & ~w18618;
assign w17390 = w3425 & ~w15574;
assign w17391 = ~w10656 & ~w13403;
assign w17392 = w2131 & w314;
assign w17393 = ~w5514 & ~w5206;
assign w17394 = w10623 & ~w18394;
assign w17395 = ~w3746 & ~w8079;
assign w17396 = ~w5927 & ~w6831;
assign w17397 = ~w9422 & ~w15841;
assign w17398 = w13338 & w8682;
assign w17399 = ~w3833 & ~w17431;
assign w17400 = ~w4826 & ~w3665;
assign w17401 = ~w8559 & ~w17598;
assign w17402 = (~w7102 & w9316) | (~w7102 & w3631) | (w9316 & w3631);
assign w17403 = ~w8445 & ~w17301;
assign w17404 = a_29 & a_55;
assign w17405 = ~w6610 & ~w8550;
assign w17406 = ~w7399 & w10764;
assign w17407 = w3514 & w18350;
assign w17408 = a_29 & a_48;
assign w17409 = ~w9712 & ~w128;
assign w17410 = ~w14684 & ~w4829;
assign w17411 = ~w14875 & w6329;
assign w17412 = ~w16656 & ~w8188;
assign w17413 = ~w7563 & ~w13680;
assign w17414 = ~w10059 & w15124;
assign w17415 = ~w11434 & ~w165;
assign w17416 = ~w729 & w18053;
assign w17417 = ~w1506 & ~w14285;
assign w17418 = a_17 & a_43;
assign w17419 = a_5 & a_54;
assign w17420 = w9544 & w4929;
assign w17421 = ~w12245 & ~w5911;
assign w17422 = ~w10791 & ~w14709;
assign w17423 = a_8 & a_38;
assign w17424 = w3030 & ~w13780;
assign w17425 = ~w11542 & ~w701;
assign w17426 = w15975 & w9932;
assign w17427 = w13961 & ~w14880;
assign w17428 = ~w16702 & ~w4786;
assign w17429 = ~w13284 & ~w6458;
assign w17430 = w10793 & w16347;
assign w17431 = a_22 & a_37;
assign w17432 = ~w2536 & ~w106;
assign w17433 = ~w11315 & ~w8548;
assign w17434 = ~w443 & ~w6239;
assign w17435 = a_4 & a_42;
assign w17436 = ~w11446 & ~w13948;
assign w17437 = ~w19106 & ~w17776;
assign w17438 = a_8 & a_20;
assign w17439 = (w13462 & w17258) | (w13462 & w10028) | (w17258 & w10028);
assign w17440 = ~w15975 & w14711;
assign w17441 = ~w8271 & w4873;
assign w17442 = ~w13095 & ~w17998;
assign w17443 = ~w15000 & ~w18297;
assign w17444 = ~w1128 & ~w1077;
assign w17445 = ~w16036 & ~w9897;
assign w17446 = ~w8897 & ~w16031;
assign w17447 = ~w11030 & ~w11451;
assign w17448 = ~w16907 & ~w18387;
assign w17449 = ~w15009 & ~w12267;
assign w17450 = w14121 & ~w16994;
assign w17451 = ~w13584 & ~w18328;
assign w17452 = a_6 & a_49;
assign w17453 = ~w6836 & w7628;
assign w17454 = ~w9251 & ~w998;
assign w17455 = ~w17392 & ~w17406;
assign w17456 = ~w7971 & ~w7677;
assign w17457 = w1553 & w2960;
assign w17458 = ~w10580 & ~w14025;
assign w17459 = ~w3066 & ~w6970;
assign w17460 = w2710 & ~w11957;
assign w17461 = ~w18725 & ~w13649;
assign w17462 = ~w7228 & ~w4572;
assign w17463 = ~w8989 & w14354;
assign w17464 = w4989 & ~w16343;
assign w17465 = w2930 & w9661;
assign w17466 = a_43 & a_57;
assign w17467 = w9155 & ~w7438;
assign w17468 = ~w17362 & ~w13577;
assign w17469 = (w17914 & w9765) | (w17914 & w17222) | (w9765 & w17222);
assign w17470 = w4180 & ~w4799;
assign w17471 = a_2 & a_41;
assign w17472 = ~w16833 & ~w9406;
assign w17473 = ~w14792 & w4574;
assign w17474 = w4029 & ~w1558;
assign w17475 = ~w3582 & ~w5907;
assign w17476 = a_57 & a_63;
assign w17477 = a_30 & a_62;
assign w17478 = ~w2120 & ~w12631;
assign w17479 = ~w11906 & ~w2161;
assign w17480 = ~w1620 & ~w8512;
assign w17481 = ~w11732 & ~w1909;
assign w17482 = ~w16813 & w16750;
assign w17483 = a_7 & a_21;
assign w17484 = w506 & w7579;
assign w17485 = a_18 & a_35;
assign w17486 = ~w9558 & ~w14347;
assign w17487 = w6225 & w18106;
assign w17488 = w16890 & w18804;
assign w17489 = a_24 & a_57;
assign w17490 = w4575 & w3420;
assign w17491 = ~w13342 & ~w3266;
assign w17492 = w5590 & w13841;
assign w17493 = a_11 & a_14;
assign w17494 = ~w13664 & ~w12025;
assign w17495 = (w9049 & w5220) | (w9049 & w11129) | (w5220 & w11129);
assign w17496 = ~w8644 & ~w16856;
assign w17497 = ~w3088 & ~w193;
assign w17498 = ~w7352 & ~w11777;
assign w17499 = w3583 & ~w17370;
assign w17500 = w12850 & w13954;
assign w17501 = w6266 & ~w3100;
assign w17502 = ~w418 & ~w12800;
assign w17503 = ~w2888 & w3852;
assign w17504 = w13259 & w16520;
assign w17505 = a_20 & a_32;
assign w17506 = (w16857 & w2896) | (w16857 & w12700) | (w2896 & w12700);
assign w17507 = ~w1135 & ~w13719;
assign w17508 = w11717 & w10422;
assign w17509 = (~w18286 & ~w111) | (~w18286 & w1435) | (~w111 & w1435);
assign w17510 = ~w6529 & w14559;
assign w17511 = ~w7284 & w17455;
assign w17512 = ~w5579 & ~w17405;
assign w17513 = ~w9153 & ~w12212;
assign w17514 = w11123 & w5200;
assign w17515 = a_6 & a_8;
assign w17516 = ~w7661 & ~w9492;
assign w17517 = w15959 & w6323;
assign w17518 = w11215 & w4689;
assign w17519 = ~w9284 & w18460;
assign w17520 = w9938 & w11822;
assign w17521 = ~w18751 & ~w1801;
assign w17522 = ~w4512 & ~w5847;
assign w17523 = ~w14356 & w16266;
assign w17524 = a_6 & a_21;
assign w17525 = a_54 & a_62;
assign w17526 = ~w4892 & ~w14471;
assign w17527 = w5667 & w5259;
assign w17528 = ~w8745 & ~w18915;
assign w17529 = w15560 & ~w410;
assign w17530 = w2228 & ~w1243;
assign w17531 = (w8836 & w14429) | (w8836 & w1308) | (w14429 & w1308);
assign w17532 = (w16174 & w4170) | (w16174 & w18536) | (w4170 & w18536);
assign w17533 = ~w9812 & ~w7808;
assign w17534 = ~w6741 & ~w4629;
assign w17535 = ~w18927 & ~w17824;
assign w17536 = ~w1733 & w17884;
assign w17537 = w14106 & ~w18556;
assign w17538 = w18277 & w15507;
assign w17539 = ~w19053 & w1786;
assign w17540 = w8725 & ~w11406;
assign w17541 = a_7 & a_32;
assign w17542 = ~w4325 & ~w18012;
assign w17543 = ~w7432 & ~w18090;
assign w17544 = (~w9711 & ~w3603) | (~w9711 & w12976) | (~w3603 & w12976);
assign w17545 = w4664 & ~w18767;
assign w17546 = ~w2875 & ~w15475;
assign w17547 = (w17788 & w9931) | (w17788 & w6324) | (w9931 & w6324);
assign w17548 = ~w6322 & ~w1261;
assign w17549 = a_10 & a_59;
assign w17550 = ~w2625 & ~w17893;
assign w17551 = a_21 & a_57;
assign w17552 = ~w4847 & ~w11727;
assign w17553 = ~w16214 & ~w17094;
assign w17554 = ~w16587 & ~w12503;
assign w17555 = ~w11105 & ~w8576;
assign w17556 = ~w16106 & ~w14564;
assign w17557 = a_1 & a_24;
assign w17558 = ~w16018 & w2116;
assign w17559 = w12495 & ~w7617;
assign w17560 = w11106 & w2799;
assign w17561 = w3221 & w13207;
assign w17562 = ~w18938 & ~w18652;
assign w17563 = ~w17030 & ~w9905;
assign w17564 = w2541 & w7612;
assign w17565 = ~w9994 & ~w13492;
assign w17566 = a_53 & a_58;
assign w17567 = w8175 & ~w10898;
assign w17568 = ~w11839 & ~w18968;
assign w17569 = w8271 & ~w4873;
assign w17570 = ~w13131 & w1226;
assign w17571 = ~w327 & ~w13179;
assign w17572 = ~w7150 & ~w5166;
assign w17573 = ~w959 & ~w13787;
assign w17574 = ~w13313 & ~w11962;
assign w17575 = ~w14034 & ~w10818;
assign w17576 = ~w11574 & ~w9583;
assign w17577 = ~w8077 & ~w1664;
assign w17578 = w109 & ~w11156;
assign w17579 = ~w1673 & w12680;
assign w17580 = (~w17322 & ~w6571) | (~w17322 & w5799) | (~w6571 & w5799);
assign w17581 = ~w13423 & w270;
assign w17582 = ~w12849 & ~w18531;
assign w17583 = w2274 & w10200;
assign w17584 = ~w4932 & ~w5991;
assign w17585 = a_15 & a_42;
assign w17586 = w3542 & ~w4723;
assign w17587 = w18151 & w18403;
assign w17588 = a_26 & a_42;
assign w17589 = w16917 & w9132;
assign w17590 = ~w16789 & ~w8972;
assign w17591 = w9609 & w16303;
assign w17592 = (~w10619 & ~w13724) | (~w10619 & w10612) | (~w13724 & w10612);
assign w17593 = a_2 & a_62;
assign w17594 = w7814 & ~w7504;
assign w17595 = ~w13353 & ~w3990;
assign w17596 = w10267 & w6247;
assign w17597 = w6988 & ~w2960;
assign w17598 = ~w10648 & w18995;
assign w17599 = (~w1669 & ~w4905) | (~w1669 & w9839) | (~w4905 & w9839);
assign w17600 = ~w18263 & ~w2158;
assign w17601 = ~w2489 & ~w5903;
assign w17602 = ~w17710 & w6565;
assign w17603 = w4005 & ~w11842;
assign w17604 = ~w14665 & ~w2087;
assign w17605 = w11403 & ~w858;
assign w17606 = a_0 & a_11;
assign w17607 = w3172 & w14978;
assign w17608 = ~w10267 & ~w6247;
assign w17609 = ~w13051 & w15546;
assign w17610 = w16588 & w16926;
assign w17611 = ~w8813 & ~w5115;
assign w17612 = w10933 & ~w12121;
assign w17613 = ~w10290 & ~w2504;
assign w17614 = ~w11271 & w9503;
assign w17615 = (w16603 & ~w5836) | (w16603 & w6336) | (~w5836 & w6336);
assign w17616 = ~w18272 & w794;
assign w17617 = ~w1942 & ~w17290;
assign w17618 = a_25 & a_51;
assign w17619 = w18025 & ~w1748;
assign w17620 = ~w8436 & w14452;
assign w17621 = ~w9530 & ~w1782;
assign w17622 = a_2 & a_25;
assign w17623 = w16006 & w8652;
assign w17624 = ~w17773 & w16979;
assign w17625 = ~w11141 & w6461;
assign w17626 = ~w15959 & ~w3428;
assign w17627 = ~w7562 & ~w17972;
assign w17628 = ~w10796 & w14298;
assign w17629 = w9250 & ~w8636;
assign w17630 = w17910 & ~w2402;
assign w17631 = ~w15558 & ~w6050;
assign w17632 = ~w17852 & ~w7005;
assign w17633 = ~w2548 & ~w18267;
assign w17634 = ~w1046 & ~w10883;
assign w17635 = w18984 & ~w16827;
assign w17636 = w3806 & w12578;
assign w17637 = w18354 & ~w14839;
assign w17638 = a_49 & a_55;
assign w17639 = (w15080 & w7366) | (w15080 & w7473) | (w7366 & w7473);
assign w17640 = w17909 & ~w16970;
assign w17641 = w8286 & ~w5809;
assign w17642 = w13311 & w786;
assign w17643 = ~w3670 & ~w8790;
assign w17644 = ~w14418 & ~w17275;
assign w17645 = ~w15487 & ~w7487;
assign w17646 = w804 & w9628;
assign w17647 = w6397 & ~w4316;
assign w17648 = w16808 & ~w8392;
assign w17649 = ~w10767 & w4209;
assign w17650 = ~w12674 & ~w17720;
assign w17651 = ~w742 & ~w16984;
assign w17652 = ~w13371 & ~w5948;
assign w17653 = ~w19080 & ~w16510;
assign w17654 = ~w18459 & ~w7267;
assign w17655 = w823 & ~w8783;
assign w17656 = ~w14312 & ~w18516;
assign w17657 = ~w17200 & ~w11647;
assign w17658 = ~w6988 & ~w5296;
assign w17659 = w13466 & ~w9563;
assign w17660 = w14168 & w6357;
assign w17661 = w10737 & w15091;
assign w17662 = w12452 & w15151;
assign w17663 = ~w6237 & w7458;
assign w17664 = ~w12194 & ~w14097;
assign w17665 = w13830 & ~w553;
assign w17666 = ~w6367 & ~w6260;
assign w17667 = (w1638 & w3807) | (w1638 & w4455) | (w3807 & w4455);
assign w17668 = w6294 & ~w15059;
assign w17669 = ~w11876 & ~w18945;
assign w17670 = w18775 & ~w7738;
assign w17671 = ~w11602 & ~w10998;
assign w17672 = ~w12560 & w17383;
assign w17673 = w15974 & w8386;
assign w17674 = ~w3523 & ~w14301;
assign w17675 = ~w10516 & ~w1230;
assign w17676 = ~w5177 & ~w11019;
assign w17677 = a_9 & a_24;
assign w17678 = w1852 & w5655;
assign w17679 = w15251 & w17284;
assign w17680 = ~w8817 & ~w681;
assign w17681 = ~w17926 & ~w14594;
assign w17682 = ~w9814 & ~w10074;
assign w17683 = w15352 & ~w12947;
assign w17684 = w16127 & ~w17817;
assign w17685 = a_29 & a_58;
assign w17686 = (w2092 & ~w17111) | (w2092 & w18453) | (~w17111 & w18453);
assign w17687 = ~w17062 & ~w3191;
assign w17688 = ~w10484 & ~w1807;
assign w17689 = (w6407 & w2769) | (w6407 & w8663) | (w2769 & w8663);
assign w17690 = ~w12782 & w9703;
assign w17691 = ~w17000 & ~w18796;
assign w17692 = ~w2491 & ~w16981;
assign w17693 = w11295 & w8250;
assign w17694 = ~w17315 & ~w15304;
assign w17695 = w13029 & ~w3300;
assign w17696 = ~w1195 & ~w1851;
assign w17697 = w5852 & w2052;
assign w17698 = ~w999 & ~w19124;
assign w17699 = (~w14287 & w16191) | (~w14287 & w2763) | (w16191 & w2763);
assign w17700 = ~w13533 & w2277;
assign w17701 = (w2870 & ~w1320) | (w2870 & w16291) | (~w1320 & w16291);
assign w17702 = ~w8834 & ~w8427;
assign w17703 = ~w5970 & ~w16044;
assign w17704 = ~w17496 & w1920;
assign w17705 = w13830 & w2964;
assign w17706 = a_40 & a_49;
assign w17707 = ~w1416 & ~w6646;
assign w17708 = ~w18494 & ~w8299;
assign w17709 = ~w1867 & ~w72;
assign w17710 = w11334 & w2742;
assign w17711 = (w7102 & w17036) | (w7102 & w1837) | (w17036 & w1837);
assign w17712 = ~w16843 & w4823;
assign w17713 = ~w17445 & ~w8476;
assign w17714 = w15336 & ~w10687;
assign w17715 = (w13037 & w10397) | (w13037 & w10231) | (w10397 & w10231);
assign w17716 = (w8836 & w8122) | (w8836 & ~w1074) | (w8122 & ~w1074);
assign w17717 = ~w8602 & ~w147;
assign w17718 = ~w8431 & w12078;
assign w17719 = ~w18059 & ~w4001;
assign w17720 = w12797 & ~w5588;
assign w17721 = a_4 & a_15;
assign w17722 = ~w18984 & w16827;
assign w17723 = ~w11822 & w16728;
assign w17724 = ~w14789 & w14802;
assign w17725 = ~w7040 & ~w4836;
assign w17726 = ~w11889 & w17848;
assign w17727 = ~w9131 & w2798;
assign w17728 = ~w1894 & w14592;
assign w17729 = w10645 & ~w18697;
assign w17730 = w1494 & w15923;
assign w17731 = w13771 & ~w1404;
assign w17732 = ~w7002 & ~w13124;
assign w17733 = (~w7768 & w16077) | (~w7768 & w17831) | (w16077 & w17831);
assign w17734 = (~w8437 & w8121) | (~w8437 & w16376) | (w8121 & w16376);
assign w17735 = w11976 & ~w16423;
assign w17736 = w4309 & ~w5290;
assign w17737 = ~w2573 & ~w4185;
assign w17738 = ~w11662 & w14261;
assign w17739 = w8215 & ~w10462;
assign w17740 = ~w13268 & ~w10930;
assign w17741 = w18397 & ~w14169;
assign w17742 = w12612 & ~w10859;
assign w17743 = a_48 & a_57;
assign w17744 = ~w9529 & ~w5440;
assign w17745 = w15074 & ~w4999;
assign w17746 = ~w18737 & ~w1907;
assign w17747 = w7488 & ~w19129;
assign w17748 = ~w4151 & ~w14023;
assign w17749 = ~w10774 & ~w14326;
assign w17750 = ~w5220 & w10301;
assign w17751 = ~w6453 & w3909;
assign w17752 = ~w11987 & ~w5842;
assign w17753 = a_6 & a_63;
assign w17754 = ~w6484 & ~w17400;
assign w17755 = w651 & w14265;
assign w17756 = w6622 & ~w1525;
assign w17757 = ~w11596 & ~w2290;
assign w17758 = ~w1027 & ~w10483;
assign w17759 = ~w16602 & ~w5111;
assign w17760 = ~w294 & ~w10379;
assign w17761 = w13664 & w4371;
assign w17762 = ~w4784 & ~w5721;
assign w17763 = ~w10097 & ~w2852;
assign w17764 = ~w14231 & w15993;
assign w17765 = ~w18473 & w9201;
assign w17766 = w12576 & w7452;
assign w17767 = ~w13480 & ~w11164;
assign w17768 = ~w11726 & ~w15898;
assign w17769 = w13219 & w15077;
assign w17770 = (~w11906 & ~w11107) | (~w11906 & w10544) | (~w11107 & w10544);
assign w17771 = ~w11845 & ~w2882;
assign w17772 = ~w1612 & ~w271;
assign w17773 = a_38 & a_62;
assign w17774 = ~w406 & ~w14669;
assign w17775 = ~w14433 & w18167;
assign w17776 = ~w6434 & ~w4466;
assign w17777 = ~w2631 & ~w402;
assign w17778 = ~w17543 & ~w2478;
assign w17779 = ~w10653 & w11498;
assign w17780 = w2352 & ~w1596;
assign w17781 = w18125 & w6205;
assign w17782 = ~w7495 & ~w12316;
assign w17783 = ~w5890 & w10996;
assign w17784 = w4155 & w7350;
assign w17785 = (~w18796 & ~w17691) | (~w18796 & w2011) | (~w17691 & w2011);
assign w17786 = a_12 & a_28;
assign w17787 = ~w4092 & w14396;
assign w17788 = ~w9714 & ~w13448;
assign w17789 = w6887 & ~w1613;
assign w17790 = ~w12919 & ~w6036;
assign w17791 = ~a_24 & w6208;
assign w17792 = ~w8731 & ~w11966;
assign w17793 = ~w18251 & ~w11630;
assign w17794 = ~w16812 & ~w7750;
assign w17795 = ~w7416 & w7721;
assign w17796 = w4288 & w11782;
assign w17797 = (~w15956 & w10330) | (~w15956 & w17870) | (w10330 & w17870);
assign w17798 = ~w11040 & ~w14616;
assign w17799 = ~w17068 & ~w16328;
assign w17800 = ~w12355 & w12055;
assign w17801 = w8088 & ~w14984;
assign w17802 = ~w16095 & w14916;
assign w17803 = w2775 & ~w1032;
assign w17804 = ~w4073 & ~w3384;
assign w17805 = ~w17928 & ~w12251;
assign w17806 = ~w8600 & w16586;
assign w17807 = w16036 & w5793;
assign w17808 = ~w16923 & ~w1444;
assign w17809 = a_43 & a_45;
assign w17810 = ~w18715 & w3736;
assign w17811 = ~w8890 & ~w18849;
assign w17812 = ~w11705 & ~w13223;
assign w17813 = w6702 & ~w4882;
assign w17814 = ~w535 & ~w14310;
assign w17815 = w16546 & ~w5356;
assign w17816 = ~w2551 & ~w16865;
assign w17817 = ~w10779 & ~w3055;
assign w17818 = ~w18234 & w16670;
assign w17819 = a_28 & a_52;
assign w17820 = ~w6496 & ~w14704;
assign w17821 = a_28 & a_45;
assign w17822 = (~w15399 & w3338) | (~w15399 & w11706) | (w3338 & w11706);
assign w17823 = ~w8287 & ~w16263;
assign w17824 = w1378 & w6252;
assign w17825 = ~w15037 & ~w11695;
assign w17826 = ~w17927 & ~w4656;
assign w17827 = ~w5317 & ~w4218;
assign w17828 = ~w8878 & w17866;
assign w17829 = ~w2897 & ~w9516;
assign w17830 = ~w16008 & ~w8451;
assign w17831 = w1501 & ~w6956;
assign w17832 = ~w14444 & ~w1400;
assign w17833 = ~w7673 & ~w1977;
assign w17834 = ~w17728 & w12707;
assign w17835 = w16278 & w11453;
assign w17836 = ~w10979 & ~w6808;
assign w17837 = ~w7433 & ~w14560;
assign w17838 = w11277 & ~w17528;
assign w17839 = w15812 & ~w5928;
assign w17840 = a_48 & w3299;
assign w17841 = w12382 & ~w597;
assign w17842 = ~w3934 & ~w16191;
assign w17843 = ~w3949 & ~w6017;
assign w17844 = w13459 & ~w1539;
assign w17845 = ~w15002 & ~w7401;
assign w17846 = ~w12291 & ~w1031;
assign w17847 = w4267 & ~w18260;
assign w17848 = ~a_49 & a_50;
assign w17849 = ~w17939 & w18252;
assign w17850 = w17137 & ~w1790;
assign w17851 = ~w7812 & ~w8262;
assign w17852 = w4852 & ~w167;
assign w17853 = ~w12371 & ~w5822;
assign w17854 = ~w19063 & ~w11667;
assign w17855 = a_19 & a_39;
assign w17856 = a_3 & a_26;
assign w17857 = ~w16112 & w18215;
assign w17858 = a_4 & a_38;
assign w17859 = ~w880 & ~w11240;
assign w17860 = ~w2590 & ~w8249;
assign w17861 = ~w11026 & ~w6631;
assign w17862 = ~w5 & ~w9761;
assign w17863 = w3029 & w8814;
assign w17864 = ~w16016 & ~w8619;
assign w17865 = ~w8623 & w8014;
assign w17866 = ~w8393 & ~w4963;
assign w17867 = ~w17182 & ~w716;
assign w17868 = a_25 & a_43;
assign w17869 = ~w2251 & ~w13430;
assign w17870 = w13082 & ~w15956;
assign w17871 = w16808 & ~w17801;
assign w17872 = ~w6181 & ~w15809;
assign w17873 = ~w12772 & ~w18084;
assign w17874 = ~w11073 & ~w2096;
assign w17875 = ~w9631 & ~w11217;
assign w17876 = ~w1855 & ~w326;
assign w17877 = w441 & ~w15727;
assign w17878 = ~w8777 & ~w9040;
assign w17879 = a_28 & a_62;
assign w17880 = ~w7020 & w16714;
assign w17881 = (w8250 & w12086) | (w8250 & w6853) | (w12086 & w6853);
assign w17882 = ~w12230 & w11716;
assign w17883 = w14522 & ~w10092;
assign w17884 = ~w7775 & ~w15334;
assign w17885 = a_26 & a_34;
assign w17886 = a_15 & a_51;
assign w17887 = ~w8432 & ~w13906;
assign w17888 = ~w10329 & ~w1682;
assign w17889 = ~w9532 & ~w18086;
assign w17890 = a_24 & a_61;
assign w17891 = ~w3835 & ~w2344;
assign w17892 = (~w15297 & ~w7419) | (~w15297 & w4579) | (~w7419 & w4579);
assign w17893 = a_6 & a_29;
assign w17894 = w5019 & ~w15172;
assign w17895 = ~w13082 & w7413;
assign w17896 = w10075 & ~w18243;
assign w17897 = w18908 & ~w14404;
assign w17898 = ~w5358 & ~w6787;
assign w17899 = ~w8263 & ~w9686;
assign w17900 = ~w1705 & ~w6428;
assign w17901 = w8284 & ~w4912;
assign w17902 = ~w1595 & w17253;
assign w17903 = w18495 & ~w18474;
assign w17904 = ~w18045 & ~w15570;
assign w17905 = w6079 & w6429;
assign w17906 = w9806 & w9971;
assign w17907 = ~w9919 & ~w1102;
assign w17908 = a_3 & a_16;
assign w17909 = ~w7424 & ~w8784;
assign w17910 = ~w307 & w8434;
assign w17911 = ~w15860 & ~w15460;
assign w17912 = a_1 & a_46;
assign w17913 = w11662 & ~w1827;
assign w17914 = ~w1074 & ~w4559;
assign w17915 = w2950 & w1908;
assign w17916 = ~w10817 & w17163;
assign w17917 = ~w868 & w17907;
assign w17918 = w8384 & w3625;
assign w17919 = w9750 & ~w10143;
assign w17920 = ~w18005 & w17513;
assign w17921 = ~w11170 & w10043;
assign w17922 = ~w10578 & ~w1130;
assign w17923 = w3014 & w8934;
assign w17924 = ~w15542 & w16973;
assign w17925 = w18184 & w10104;
assign w17926 = ~w18396 & w960;
assign w17927 = w17762 & ~w1547;
assign w17928 = (~w17230 & ~w5452) | (~w17230 & w11999) | (~w5452 & w11999);
assign w17929 = w11044 & ~w5768;
assign w17930 = w16997 & w18498;
assign w17931 = ~w6422 & ~w3677;
assign w17932 = w17574 & ~w6465;
assign w17933 = ~w808 & ~w13926;
assign w17934 = w947 & ~w12023;
assign w17935 = ~w9604 & ~w265;
assign w17936 = ~w9990 & w8754;
assign w17937 = ~w10522 & ~w10835;
assign w17938 = ~w13139 & ~w18275;
assign w17939 = ~w3044 & ~w3822;
assign w17940 = w15423 & w17400;
assign w17941 = ~w3364 & ~w1343;
assign w17942 = ~w998 & ~w681;
assign w17943 = ~w17464 & ~w9189;
assign w17944 = ~w13596 & ~w8572;
assign w17945 = ~w8327 & ~w10494;
assign w17946 = a_45 & a_63;
assign w17947 = ~w3987 & ~w18301;
assign w17948 = ~w7563 & ~w5757;
assign w17949 = w13581 & ~w2850;
assign w17950 = ~w5398 & ~w6590;
assign w17951 = ~w14978 & ~w17164;
assign w17952 = ~w15234 & w18187;
assign w17953 = ~w11024 & w13108;
assign w17954 = ~w3370 & ~w9680;
assign w17955 = a_33 & a_47;
assign w17956 = w6003 & w7241;
assign w17957 = w717 & ~w7213;
assign w17958 = ~w3186 & ~w766;
assign w17959 = ~w7067 & ~w6494;
assign w17960 = ~w8993 & ~w8286;
assign w17961 = ~w12933 & ~w15964;
assign w17962 = ~w13601 & ~w6421;
assign w17963 = a_12 & a_56;
assign w17964 = ~a_6 & w6133;
assign w17965 = ~w11556 & ~w4302;
assign w17966 = w4996 & ~w6269;
assign w17967 = ~w11641 & ~w9785;
assign w17968 = ~w7506 & ~w3660;
assign w17969 = ~w17522 & ~w9787;
assign w17970 = w1865 & ~w9223;
assign w17971 = ~w2270 & w1879;
assign w17972 = (~w16667 & ~w12098) | (~w16667 & w10233) | (~w12098 & w10233);
assign w17973 = w1844 & ~w4519;
assign w17974 = ~w7444 & ~w2751;
assign w17975 = ~w7568 & ~w10566;
assign w17976 = ~w8132 & ~w7384;
assign w17977 = ~w6619 & ~w11423;
assign w17978 = a_6 & a_56;
assign w17979 = a_3 & a_40;
assign w17980 = ~w11863 & ~w16038;
assign w17981 = (~w9291 & ~w11017) | (~w9291 & w12668) | (~w11017 & w12668);
assign w17982 = a_16 & a_31;
assign w17983 = ~w9629 & w15032;
assign w17984 = w11416 & ~w17433;
assign w17985 = ~w10810 & ~w3170;
assign w17986 = w11394 & ~w611;
assign w17987 = ~w18346 & ~w10920;
assign w17988 = ~w8258 & w4287;
assign w17989 = ~w14102 & ~w7787;
assign w17990 = ~w14620 & ~w9870;
assign w17991 = ~w11340 & ~w1546;
assign w17992 = ~w2385 & ~w17759;
assign w17993 = w5351 & w17418;
assign w17994 = ~w3443 & ~w12019;
assign w17995 = (w7102 & w9579) | (w7102 & w7187) | (w9579 & w7187);
assign w17996 = w7671 & ~w17069;
assign w17997 = w88 & w4409;
assign w17998 = (~w16764 & ~w12751) | (~w16764 & w3369) | (~w12751 & w3369);
assign w17999 = ~w14658 & ~w5770;
assign w18000 = ~w7830 & w15427;
assign w18001 = ~w8205 & ~w17217;
assign w18002 = w6853 & w7608;
assign w18003 = w17892 & ~w9329;
assign w18004 = ~w4267 & w16083;
assign w18005 = ~w16015 & w9849;
assign w18006 = ~w16896 & ~w11270;
assign w18007 = ~w13322 & ~w6942;
assign w18008 = ~w13973 & w5053;
assign w18009 = ~w7899 & w2065;
assign w18010 = w7160 & ~w15895;
assign w18011 = w110 & w6369;
assign w18012 = w4804 & w17218;
assign w18013 = w13220 & ~w7268;
assign w18014 = ~w15 & ~w8893;
assign w18015 = a_37 & a_38;
assign w18016 = ~w978 & w10376;
assign w18017 = w9085 & ~w15319;
assign w18018 = w940 & ~w11275;
assign w18019 = w4896 & ~w14654;
assign w18020 = ~w10747 & ~w4165;
assign w18021 = w5033 & ~w16349;
assign w18022 = w10002 & ~w2039;
assign w18023 = w11997 & w19126;
assign w18024 = ~w9469 & ~w2404;
assign w18025 = a_39 & a_51;
assign w18026 = ~w12248 & ~w2600;
assign w18027 = a_12 & a_33;
assign w18028 = ~w11815 & ~w7983;
assign w18029 = w15610 & ~w18624;
assign w18030 = w353 & w3276;
assign w18031 = ~w10621 & ~w9559;
assign w18032 = ~w15552 & w15192;
assign w18033 = (~w4190 & ~w4878) | (~w4190 & w9375) | (~w4878 & w9375);
assign w18034 = a_28 & a_49;
assign w18035 = w17489 & ~w16120;
assign w18036 = ~w8939 & w9195;
assign w18037 = a_11 & a_15;
assign w18038 = ~w9618 & ~w13424;
assign w18039 = w2540 & ~w10373;
assign w18040 = ~w9140 & ~w10807;
assign w18041 = (w14221 & w8635) | (w14221 & w11689) | (w8635 & w11689);
assign w18042 = (w10004 & ~w5720) | (w10004 & w12159) | (~w5720 & w12159);
assign w18043 = w12862 & w16230;
assign w18044 = ~w7533 & ~w5241;
assign w18045 = ~w5439 & w2173;
assign w18046 = ~w12648 & w2184;
assign w18047 = w11516 & ~w12995;
assign w18048 = ~w9278 & ~w18465;
assign w18049 = ~w10635 & ~w2246;
assign w18050 = ~w1836 & ~w11888;
assign w18051 = a_18 & a_26;
assign w18052 = ~w2127 & ~w2984;
assign w18053 = ~w3928 & ~w17890;
assign w18054 = ~w18369 & w18164;
assign w18055 = ~w2778 & ~w17041;
assign w18056 = ~w9044 & ~w18783;
assign w18057 = w3078 & ~w14662;
assign w18058 = w16675 & ~w14461;
assign w18059 = ~w5232 & w5379;
assign w18060 = w4376 & ~w15355;
assign w18061 = w11322 & ~w13769;
assign w18062 = ~w11931 & ~w10005;
assign w18063 = ~w17554 & ~w10507;
assign w18064 = ~w4750 & w13439;
assign w18065 = w10132 & w15651;
assign w18066 = w5439 & ~w7033;
assign w18067 = ~w10092 & ~w2298;
assign w18068 = ~w4667 & ~w18311;
assign w18069 = w15873 & w6778;
assign w18070 = ~w6253 & ~w17261;
assign w18071 = ~w5693 & ~w9658;
assign w18072 = ~w5130 & w8281;
assign w18073 = (~w9701 & ~w12595) | (~w9701 & w19200) | (~w12595 & w19200);
assign w18074 = (~w16072 & w175) | (~w16072 & w5969) | (w175 & w5969);
assign w18075 = ~w18525 & ~w16090;
assign w18076 = ~w10399 & ~w1143;
assign w18077 = ~w5740 & ~w11954;
assign w18078 = ~w12588 & ~w17434;
assign w18079 = w16529 & ~w16935;
assign w18080 = ~w10666 & ~w925;
assign w18081 = w15554 & w17485;
assign w18082 = ~w5849 & w5897;
assign w18083 = ~w8668 & w5864;
assign w18084 = w8873 & ~w992;
assign w18085 = ~w4484 & ~w9573;
assign w18086 = ~w13767 & w14017;
assign w18087 = w13379 & ~w7557;
assign w18088 = ~w18819 & ~w3471;
assign w18089 = ~w11374 & ~w7642;
assign w18090 = w15357 & ~w6910;
assign w18091 = ~w11704 & ~w6242;
assign w18092 = ~w2315 & ~w18376;
assign w18093 = w17620 & w6399;
assign w18094 = ~w4693 & ~w4457;
assign w18095 = w923 & w6339;
assign w18096 = ~w11838 & ~w11145;
assign w18097 = w10844 & w8763;
assign w18098 = a_5 & a_19;
assign w18099 = ~w17233 & ~w5209;
assign w18100 = w9061 & w15390;
assign w18101 = a_18 & a_50;
assign w18102 = ~w10534 & w6503;
assign w18103 = (a_35 & w18485) | (a_35 & w4423) | (w18485 & w4423);
assign w18104 = ~w13576 & ~w9929;
assign w18105 = ~w16501 & ~w12608;
assign w18106 = ~w7882 & ~w9717;
assign w18107 = w17691 & w3141;
assign w18108 = (~w1962 & w12059) | (~w1962 & w16759) | (w12059 & w16759);
assign w18109 = ~w6149 & ~w160;
assign w18110 = w12105 & w3074;
assign w18111 = ~w10998 & w15174;
assign w18112 = a_12 & w4923;
assign w18113 = w3795 & ~w556;
assign w18114 = ~w8135 & ~w12378;
assign w18115 = ~w9632 & ~w3989;
assign w18116 = ~w3021 & ~w1944;
assign w18117 = ~w8326 & ~w10561;
assign w18118 = w4641 & ~w15940;
assign w18119 = ~w4011 & w7302;
assign w18120 = ~w4144 & ~w135;
assign w18121 = w4653 & ~w3387;
assign w18122 = ~w10270 & ~w2095;
assign w18123 = w8251 & ~w3670;
assign w18124 = ~w16559 & ~w1840;
assign w18125 = (~w16960 & ~w9528) | (~w16960 & w13230) | (~w9528 & w13230);
assign w18126 = ~w12694 & ~w7325;
assign w18127 = ~w16689 & ~w6104;
assign w18128 = ~w1535 & w9815;
assign w18129 = w6278 & ~w14553;
assign w18130 = (~w11181 & ~w6820) | (~w11181 & w13231) | (~w6820 & w13231);
assign w18131 = a_3 & a_35;
assign w18132 = ~w6504 & ~w10040;
assign w18133 = ~w111 & w4141;
assign w18134 = ~w17388 & ~w9975;
assign w18135 = ~w17010 & w8422;
assign w18136 = ~w8284 & w4912;
assign w18137 = w3968 & w13200;
assign w18138 = w5260 & ~w16555;
assign w18139 = ~w3429 & ~w5236;
assign w18140 = a_18 & a_53;
assign w18141 = (~w5830 & ~w13745) | (~w5830 & w3820) | (~w13745 & w3820);
assign w18142 = ~w10392 & w18638;
assign w18143 = ~w15179 & ~w971;
assign w18144 = ~w7970 & ~w17623;
assign w18145 = ~w2418 & ~w337;
assign w18146 = w2591 & ~w15793;
assign w18147 = w7240 & w13653;
assign w18148 = w12641 & ~w1514;
assign w18149 = ~w16725 & ~w7745;
assign w18150 = (~w9036 & ~w1170) | (~w9036 & w12414) | (~w1170 & w12414);
assign w18151 = ~w16574 & ~w5057;
assign w18152 = ~w11639 & ~w9972;
assign w18153 = ~w16599 & ~w13715;
assign w18154 = w16199 & w18606;
assign w18155 = w8897 & w16031;
assign w18156 = (~w9497 & ~w8603) | (~w9497 & w9097) | (~w8603 & w9097);
assign w18157 = w1897 & ~w2200;
assign w18158 = w17785 & ~w4840;
assign w18159 = w18277 & ~w6344;
assign w18160 = w9090 & w8310;
assign w18161 = ~w16676 & w1368;
assign w18162 = w16525 & ~w444;
assign w18163 = ~w682 & ~w2587;
assign w18164 = ~w15076 & ~w9032;
assign w18165 = ~w18895 & ~w8703;
assign w18166 = ~w15925 & ~w8246;
assign w18167 = ~w5329 & ~w18048;
assign w18168 = w8312 & w6239;
assign w18169 = ~w15514 & ~w17493;
assign w18170 = ~w5120 & ~w16861;
assign w18171 = ~w999 & ~w5939;
assign w18172 = ~w16633 & ~w7999;
assign w18173 = ~w12635 & ~w9203;
assign w18174 = ~w15010 & w9562;
assign w18175 = ~w17921 & ~w13180;
assign w18176 = (~w13831 & ~w16014) | (~w13831 & w7140) | (~w16014 & w7140);
assign w18177 = ~w11789 & ~w11104;
assign w18178 = ~w11210 & ~w4055;
assign w18179 = w16523 & ~w6602;
assign w18180 = ~w17326 & ~w2524;
assign w18181 = ~w15250 & ~w3310;
assign w18182 = a_39 & a_53;
assign w18183 = a_45 & a_47;
assign w18184 = w1307 & w10995;
assign w18185 = ~w11745 & ~w18248;
assign w18186 = w18884 & ~w17861;
assign w18187 = ~w14670 & ~w18559;
assign w18188 = ~w6902 & ~w14213;
assign w18189 = ~w5104 & w3255;
assign w18190 = ~w12696 & ~w4850;
assign w18191 = ~w8334 & w17079;
assign w18192 = a_22 & a_41;
assign w18193 = ~w13267 & ~w16353;
assign w18194 = w14539 & w16220;
assign w18195 = w18718 & w9316;
assign w18196 = ~w4590 & w8554;
assign w18197 = w3737 & w4923;
assign w18198 = ~w4576 & ~w1213;
assign w18199 = (~w15080 & w40) | (~w15080 & w5230) | (w40 & w5230);
assign w18200 = a_18 & a_61;
assign w18201 = ~w4758 & ~w4446;
assign w18202 = (~w3806 & ~w6295) | (~w3806 & w12684) | (~w6295 & w12684);
assign w18203 = ~w8078 & ~w13325;
assign w18204 = ~w2721 & ~w7585;
assign w18205 = ~w658 & ~w13792;
assign w18206 = ~w7493 & ~w3032;
assign w18207 = w17743 & w10428;
assign w18208 = ~w7631 & ~w12571;
assign w18209 = (~w2602 & ~w4665) | (~w2602 & w4017) | (~w4665 & w4017);
assign w18210 = w13298 & w12756;
assign w18211 = ~w11755 & ~w18040;
assign w18212 = ~w11266 & w5591;
assign w18213 = w13911 & ~w4274;
assign w18214 = ~w13487 & ~w11829;
assign w18215 = (~w17449 & ~w13748) | (~w17449 & w9111) | (~w13748 & w9111);
assign w18216 = (w13422 & w2493) | (w13422 & w1181) | (w2493 & w1181);
assign w18217 = w6106 & ~w4613;
assign w18218 = (w9221 & w15176) | (w9221 & w9322) | (w15176 & w9322);
assign w18219 = ~w14951 & ~w10019;
assign w18220 = w1345 & w4438;
assign w18221 = a_25 & a_57;
assign w18222 = ~w3745 & ~w13538;
assign w18223 = w11594 & w13079;
assign w18224 = w13202 & w3054;
assign w18225 = w4138 & ~w12633;
assign w18226 = a_30 & a_60;
assign w18227 = ~w17167 & ~w14546;
assign w18228 = ~w336 & ~w17841;
assign w18229 = ~w12080 & w3129;
assign w18230 = ~w2480 & ~w7323;
assign w18231 = ~w8381 & ~w6351;
assign w18232 = ~w16673 & ~w1222;
assign w18233 = a_35 & a_39;
assign w18234 = ~w16274 & ~w4809;
assign w18235 = a_11 & a_53;
assign w18236 = a_30 & a_45;
assign w18237 = ~w7748 & w15559;
assign w18238 = w13768 & ~w1503;
assign w18239 = w14339 & ~w19124;
assign w18240 = (~w10401 & w3984) | (~w10401 & w13394) | (w3984 & w13394);
assign w18241 = w1688 & ~w18679;
assign w18242 = w305 & w3917;
assign w18243 = ~w6123 & ~w15770;
assign w18244 = ~w12978 & ~w15355;
assign w18245 = ~w13627 & ~w5103;
assign w18246 = ~w18207 & ~w9268;
assign w18247 = ~w8830 & ~w12097;
assign w18248 = w16651 & w15078;
assign w18249 = ~w13073 & ~w1066;
assign w18250 = ~w11559 & ~w18347;
assign w18251 = ~w3851 & ~w11360;
assign w18252 = ~w869 & ~w8457;
assign w18253 = w5771 & w743;
assign w18254 = ~w6853 & w11173;
assign w18255 = w6961 & w13470;
assign w18256 = ~w15734 & w16223;
assign w18257 = ~w4346 & ~w17924;
assign w18258 = ~w13735 & ~w10297;
assign w18259 = (~w12631 & ~w4770) | (~w12631 & w17478) | (~w4770 & w17478);
assign w18260 = ~w9480 & ~w5423;
assign w18261 = a_27 & a_58;
assign w18262 = w220 & w16488;
assign w18263 = w16224 & w13485;
assign w18264 = ~w28 & ~w550;
assign w18265 = ~w12456 & w15306;
assign w18266 = ~w17021 & ~w11345;
assign w18267 = ~w3954 & ~w7828;
assign w18268 = ~w18211 & w10735;
assign w18269 = w3221 & ~w2774;
assign w18270 = ~w14244 & ~w14856;
assign w18271 = ~w8323 & ~w13952;
assign w18272 = w15578 & w3304;
assign w18273 = a_20 & a_45;
assign w18274 = ~w13445 & ~w15798;
assign w18275 = a_24 & a_43;
assign w18276 = ~w17697 & ~w3442;
assign w18277 = a_3 & a_59;
assign w18278 = w1464 & w15545;
assign w18279 = (~w11446 & w11949) | (~w11446 & w18128) | (w11949 & w18128);
assign w18280 = ~w6752 & w17235;
assign w18281 = ~w2679 & ~w8954;
assign w18282 = ~w15644 & w13150;
assign w18283 = w2807 & w3832;
assign w18284 = w14689 & ~w6517;
assign w18285 = w17599 & ~w6584;
assign w18286 = ~w3450 & ~w12884;
assign w18287 = ~w15672 & ~w3815;
assign w18288 = ~w11485 & w4545;
assign w18289 = a_40 & a_61;
assign w18290 = ~w6218 & ~w12058;
assign w18291 = ~w11483 & w16203;
assign w18292 = ~w15311 & w58;
assign w18293 = ~w10560 & ~w1436;
assign w18294 = ~w6116 & w2794;
assign w18295 = w18543 & ~w656;
assign w18296 = a_49 & a_60;
assign w18297 = ~w14060 & ~w510;
assign w18298 = ~w2284 & ~w14732;
assign w18299 = ~w9651 & w4523;
assign w18300 = ~w13564 & w15213;
assign w18301 = w10664 & w1379;
assign w18302 = w5311 & w13982;
assign w18303 = (~w16432 & w15662) | (~w16432 & w8556) | (w15662 & w8556);
assign w18304 = ~w13442 & ~w12851;
assign w18305 = ~w708 & ~w445;
assign w18306 = a_38 & a_58;
assign w18307 = ~w13911 & w4274;
assign w18308 = w5816 & ~w17548;
assign w18309 = ~w9184 & ~w15648;
assign w18310 = ~w17505 & ~w15958;
assign w18311 = ~w6844 & ~w5225;
assign w18312 = ~w19004 & ~w1875;
assign w18313 = a_28 & a_32;
assign w18314 = (~w15268 & w3208) | (~w15268 & w4201) | (w3208 & w4201);
assign w18315 = ~w16405 & ~w18467;
assign w18316 = ~w15880 & w17744;
assign w18317 = ~w18385 & w1459;
assign w18318 = ~w11131 & ~w12000;
assign w18319 = w12334 & ~w12992;
assign w18320 = ~w15757 & ~w3294;
assign w18321 = ~w2287 & ~w12698;
assign w18322 = a_17 & a_35;
assign w18323 = ~w17126 & ~w13697;
assign w18324 = w14715 & ~w5374;
assign w18325 = ~w12617 & w3651;
assign w18326 = w13345 & w438;
assign w18327 = ~w11505 & ~w17710;
assign w18328 = w7773 & ~w66;
assign w18329 = ~w8697 & ~w10776;
assign w18330 = ~w8727 & ~w11228;
assign w18331 = ~w8230 & ~w399;
assign w18332 = ~w1571 & ~w7313;
assign w18333 = w18487 & ~w5052;
assign w18334 = w15285 & w2649;
assign w18335 = w1030 & ~w4738;
assign w18336 = ~w5372 & ~w18809;
assign w18337 = a_6 & a_26;
assign w18338 = ~w3552 & ~w1683;
assign w18339 = ~w10254 & ~w15036;
assign w18340 = ~w5560 & w16685;
assign w18341 = ~w2012 & ~w15055;
assign w18342 = w10732 & w7459;
assign w18343 = ~w5216 & w7976;
assign w18344 = ~w245 & w367;
assign w18345 = ~w958 & w8729;
assign w18346 = a_52 & a_55;
assign w18347 = w18607 & w4573;
assign w18348 = ~w12810 & w13983;
assign w18349 = ~w8602 & ~w17484;
assign w18350 = a_8 & a_45;
assign w18351 = ~w18792 & ~w14716;
assign w18352 = ~w18067 & w14522;
assign w18353 = ~w14512 & ~w4968;
assign w18354 = ~w9522 & ~w10678;
assign w18355 = ~w18131 & ~w4055;
assign w18356 = a_33 & a_48;
assign w18357 = ~w63 & w9252;
assign w18358 = ~w15489 & ~w14237;
assign w18359 = ~w17977 & ~w456;
assign w18360 = w10449 & ~w18219;
assign w18361 = ~w8349 & ~w10391;
assign w18362 = w19011 & w6907;
assign w18363 = ~w11992 & ~w5853;
assign w18364 = a_5 & a_38;
assign w18365 = (w4559 & w15742) | (w4559 & w18073) | (w15742 & w18073);
assign w18366 = ~w6701 & ~w18273;
assign w18367 = ~w4073 & w18226;
assign w18368 = ~w16588 & ~w16926;
assign w18369 = a_5 & a_33;
assign w18370 = ~w432 & w11844;
assign w18371 = ~w5164 & ~w3689;
assign w18372 = w9679 & ~w5391;
assign w18373 = w13106 & ~w3579;
assign w18374 = ~w912 & ~w8161;
assign w18375 = (~w701 & ~w17425) | (~w701 & w9978) | (~w17425 & w9978);
assign w18376 = w7469 & w14270;
assign w18377 = ~w18715 & ~w9240;
assign w18378 = ~w5390 & w5148;
assign w18379 = w2923 & ~w8351;
assign w18380 = ~w4793 & ~w4838;
assign w18381 = ~w9996 & ~w15045;
assign w18382 = ~w3478 & ~w7820;
assign w18383 = w10473 & ~w11955;
assign w18384 = ~w10252 & ~w16105;
assign w18385 = ~w12354 & ~w6183;
assign w18386 = ~w12340 & ~w15432;
assign w18387 = ~w4125 & w12892;
assign w18388 = ~w5795 & w18681;
assign w18389 = ~w11058 & ~w6121;
assign w18390 = ~w10053 & w6570;
assign w18391 = ~w11492 & w11140;
assign w18392 = a_50 & a_58;
assign w18393 = a_35 & a_43;
assign w18394 = ~w12208 & ~w6806;
assign w18395 = w13545 & ~w3153;
assign w18396 = ~w16521 & ~w11482;
assign w18397 = a_22 & a_52;
assign w18398 = w10172 & w16622;
assign w18399 = ~w11296 & ~w13006;
assign w18400 = ~w15443 & ~w298;
assign w18401 = ~w4386 & ~w13117;
assign w18402 = w7070 & ~w2663;
assign w18403 = ~w8841 & ~w196;
assign w18404 = (a_53 & w3227) | (a_53 & w8298) | (w3227 & w8298);
assign w18405 = ~w7474 & ~w1957;
assign w18406 = w18306 & w13601;
assign w18407 = a_3 & a_7;
assign w18408 = ~w11470 & ~w4034;
assign w18409 = ~w10437 & ~w7026;
assign w18410 = ~w10873 & w9549;
assign w18411 = w12606 & ~w15486;
assign w18412 = ~w2858 & ~w5359;
assign w18413 = (w15159 & w2769) | (w15159 & w1552) | (w2769 & w1552);
assign w18414 = ~w14716 & ~w14897;
assign w18415 = w5769 & w4388;
assign w18416 = w10320 & w2223;
assign w18417 = ~w7001 & ~w9479;
assign w18418 = ~w13085 & ~w11074;
assign w18419 = ~w18017 & ~w14161;
assign w18420 = ~w18520 & w18421;
assign w18421 = ~w3524 & ~w5639;
assign w18422 = a_6 & a_25;
assign w18423 = ~w785 & ~w10688;
assign w18424 = ~w4358 & ~w10689;
assign w18425 = ~w6941 & ~w13258;
assign w18426 = ~w8469 & w8560;
assign w18427 = ~w7230 & w6661;
assign w18428 = a_17 & a_52;
assign w18429 = ~w5132 & ~w18322;
assign w18430 = ~w7550 & ~w18814;
assign w18431 = (~w7341 & ~w1962) | (~w7341 & w13285) | (~w1962 & w13285);
assign w18432 = ~w3245 & ~w1870;
assign w18433 = ~w4366 & ~w8967;
assign w18434 = ~w16245 & ~w10866;
assign w18435 = ~w15104 & ~w11274;
assign w18436 = w16498 & w10030;
assign w18437 = ~w16008 & ~w8922;
assign w18438 = w7501 & ~w3942;
assign w18439 = w1636 & ~w1696;
assign w18440 = w8304 & ~w1418;
assign w18441 = ~w17665 & w6890;
assign w18442 = ~w4589 & ~w7491;
assign w18443 = a_4 & a_63;
assign w18444 = ~w15722 & ~w5710;
assign w18445 = w5763 & w5640;
assign w18446 = (~w7968 & ~w11148) | (~w7968 & w18795) | (~w11148 & w18795);
assign w18447 = ~w19140 & ~w6833;
assign w18448 = w12124 & ~w12357;
assign w18449 = ~w834 & ~w6283;
assign w18450 = ~w12317 & w17184;
assign w18451 = a_57 & a_60;
assign w18452 = ~w11879 & w6238;
assign w18453 = ~w5881 & w2092;
assign w18454 = ~w7485 & w10438;
assign w18455 = (w7969 & w10330) | (w7969 & w5407) | (w10330 & w5407);
assign w18456 = w278 & ~w6502;
assign w18457 = ~w18175 & w7758;
assign w18458 = a_12 & a_60;
assign w18459 = a_4 & a_46;
assign w18460 = (w3580 & w17506) | (w3580 & w4210) | (w17506 & w4210);
assign w18461 = ~w905 & ~w4049;
assign w18462 = ~w5804 & ~w17818;
assign w18463 = w8052 & ~w17833;
assign w18464 = ~w12012 & ~w11871;
assign w18465 = w2961 & w9331;
assign w18466 = ~w13958 & ~w5462;
assign w18467 = (~w1699 & ~w1958) | (~w1699 & w12387) | (~w1958 & w12387);
assign w18468 = a_44 & a_51;
assign w18469 = w14034 & w6981;
assign w18470 = ~w5702 & ~w7679;
assign w18471 = ~w1454 & ~w7982;
assign w18472 = ~w6035 & ~w17816;
assign w18473 = ~w18904 & ~w9093;
assign w18474 = ~w8099 & ~w6525;
assign w18475 = ~w9034 & ~w7247;
assign w18476 = ~w73 & ~w11925;
assign w18477 = w2868 & ~w8535;
assign w18478 = ~w17898 & w843;
assign w18479 = ~w14140 & ~w6686;
assign w18480 = (~w7102 & w19132) | (~w7102 & w6142) | (w19132 & w6142);
assign w18481 = ~w8670 & ~w1593;
assign w18482 = ~w4666 & ~w9696;
assign w18483 = ~w17777 & ~w7542;
assign w18484 = w9347 & ~w6877;
assign w18485 = a_7 & a_62;
assign w18486 = ~w6950 & ~w7147;
assign w18487 = ~w13676 & ~w17093;
assign w18488 = ~w5084 & ~w16309;
assign w18489 = ~w10852 & ~w10783;
assign w18490 = ~w4312 & ~w11958;
assign w18491 = w9929 & ~w4110;
assign w18492 = ~w7165 & ~w4377;
assign w18493 = w6491 & ~w10558;
assign w18494 = ~w15820 & ~w5940;
assign w18495 = a_36 & a_47;
assign w18496 = ~w4533 & ~w11975;
assign w18497 = ~a_8 & ~w19009;
assign w18498 = ~w18512 & ~w18147;
assign w18499 = (w17667 & w10330) | (w17667 & w14206) | (w10330 & w14206);
assign w18500 = w2598 & w19193;
assign w18501 = ~w6001 & w2562;
assign w18502 = ~w18323 & w1421;
assign w18503 = a_10 & a_36;
assign w18504 = ~w6982 & ~w16440;
assign w18505 = ~w12905 & ~w1815;
assign w18506 = w2116 & ~w18818;
assign w18507 = w7891 & w658;
assign w18508 = ~w13692 & ~w749;
assign w18509 = ~w17416 & w14676;
assign w18510 = ~w5838 & ~w2957;
assign w18511 = w10080 & w5560;
assign w18512 = ~w7240 & ~w13653;
assign w18513 = ~w18755 & ~w10451;
assign w18514 = w2017 & ~w14695;
assign w18515 = w18418 & ~w5953;
assign w18516 = ~w7545 & ~w7464;
assign w18517 = a_1 & a_57;
assign w18518 = ~w18184 & ~w10104;
assign w18519 = w15135 & ~w2166;
assign w18520 = w18336 & ~w13650;
assign w18521 = w12683 & w6271;
assign w18522 = w11788 & ~w6962;
assign w18523 = ~w13627 & w4742;
assign w18524 = w1103 & ~w9832;
assign w18525 = a_25 & a_58;
assign w18526 = w1700 & ~w8303;
assign w18527 = w6193 & ~w2597;
assign w18528 = a_2 & a_6;
assign w18529 = w11927 & ~w12845;
assign w18530 = ~w17610 & ~w12211;
assign w18531 = w2269 & ~w10027;
assign w18532 = w15871 & ~w17748;
assign w18533 = ~w14551 & ~w10986;
assign w18534 = ~w4228 & ~w16346;
assign w18535 = w4168 & w7367;
assign w18536 = ~w11408 & w16174;
assign w18537 = a_36 & a_45;
assign w18538 = ~w10893 & w18230;
assign w18539 = ~w678 & ~w8979;
assign w18540 = w7562 & w17972;
assign w18541 = a_48 & a_62;
assign w18542 = w3318 & ~w7378;
assign w18543 = a_4 & a_25;
assign w18544 = ~w8838 & w9694;
assign w18545 = ~w1246 & ~w11621;
assign w18546 = ~w13830 & w11659;
assign w18547 = w13544 & w13368;
assign w18548 = ~w1291 & ~w3464;
assign w18549 = ~w11888 & ~w293;
assign w18550 = (~w8900 & w3850) | (~w8900 & w2198) | (w3850 & w2198);
assign w18551 = ~w11762 & w5044;
assign w18552 = w5654 & ~w18865;
assign w18553 = ~w2171 & ~w4444;
assign w18554 = ~w16344 & ~w5774;
assign w18555 = ~w4603 & ~w328;
assign w18556 = ~w15996 & ~w13205;
assign w18557 = w15068 & w11196;
assign w18558 = a_55 & a_62;
assign w18559 = ~w8267 & ~w4787;
assign w18560 = ~w15833 & ~w18907;
assign w18561 = ~w18869 & ~w4199;
assign w18562 = ~w477 & ~w17835;
assign w18563 = ~w15516 & ~w10041;
assign w18564 = ~w99 & ~w3574;
assign w18565 = ~w14595 & w5281;
assign w18566 = ~w11940 & ~w1309;
assign w18567 = ~w415 & ~w7525;
assign w18568 = w10589 & w8818;
assign w18569 = w10534 & ~w12791;
assign w18570 = w4820 & ~w11450;
assign w18571 = ~w5916 & ~w12457;
assign w18572 = w2408 & w7816;
assign w18573 = ~w8443 & ~w11984;
assign w18574 = ~w10501 & ~w173;
assign w18575 = ~w5099 & ~w13382;
assign w18576 = w9514 & ~w18932;
assign w18577 = w13489 & w11400;
assign w18578 = ~w7760 & ~w943;
assign w18579 = a_3 & a_23;
assign w18580 = w11491 & w9582;
assign w18581 = w3897 & ~w14968;
assign w18582 = ~w1740 & ~w14629;
assign w18583 = w16014 & w9453;
assign w18584 = ~w10285 & w8573;
assign w18585 = w15789 & ~w11522;
assign w18586 = ~w14447 & ~w1318;
assign w18587 = w16954 & ~w789;
assign w18588 = ~w8442 & w923;
assign w18589 = ~w17923 & ~w16078;
assign w18590 = ~w4138 & w5041;
assign w18591 = w15193 & w931;
assign w18592 = a_20 & a_21;
assign w18593 = w13328 & ~w12024;
assign w18594 = ~w2818 & ~w4514;
assign w18595 = w11041 & w5429;
assign w18596 = a_27 & a_61;
assign w18597 = ~w3514 & w18630;
assign w18598 = (~w7047 & ~w2660) | (~w7047 & w1064) | (~w2660 & w1064);
assign w18599 = w394 & w8214;
assign w18600 = a_23 & a_45;
assign w18601 = ~w14289 & ~w18102;
assign w18602 = ~w16782 & ~w12675;
assign w18603 = w10705 & ~w10864;
assign w18604 = w9909 & w10427;
assign w18605 = (w14695 & ~w6223) | (w14695 & w19144) | (~w6223 & w19144);
assign w18606 = (~w5364 & ~w13345) | (~w5364 & w14891) | (~w13345 & w14891);
assign w18607 = a_4 & a_26;
assign w18608 = ~w17450 & ~w11904;
assign w18609 = ~w18655 & ~w15301;
assign w18610 = ~w11366 & ~w16581;
assign w18611 = ~w13345 & ~w438;
assign w18612 = ~w14492 & ~w12548;
assign w18613 = w10223 & w5806;
assign w18614 = ~w7322 & ~w1406;
assign w18615 = a_41 & a_49;
assign w18616 = ~w10131 & ~w15949;
assign w18617 = ~w18395 & ~w16368;
assign w18618 = ~w14229 & ~w2848;
assign w18619 = ~w9252 & w4900;
assign w18620 = a_1 & a_15;
assign w18621 = ~w11654 & ~w7776;
assign w18622 = (~w10430 & w13701) | (~w10430 & w9861) | (w13701 & w9861);
assign w18623 = ~w15971 & ~w5196;
assign w18624 = ~w18794 & ~w16166;
assign w18625 = w4970 & ~w1919;
assign w18626 = w3239 & ~w9940;
assign w18627 = ~w521 & ~w7810;
assign w18628 = ~w1889 & w7549;
assign w18629 = ~w17221 & ~w14136;
assign w18630 = ~w3729 & ~w4221;
assign w18631 = a_48 & a_56;
assign w18632 = ~w18582 & w1425;
assign w18633 = a_1 & a_18;
assign w18634 = ~w16329 & ~w4085;
assign w18635 = ~w10294 & ~w18475;
assign w18636 = ~w6586 & ~w12541;
assign w18637 = (~w8182 & w7015) | (~w8182 & w11418) | (w7015 & w11418);
assign w18638 = ~w8629 & ~w11673;
assign w18639 = ~w1847 & ~w16996;
assign w18640 = ~w15066 & ~w11580;
assign w18641 = w15698 & ~w9773;
assign w18642 = w18882 & w5160;
assign w18643 = ~w3201 & ~w1447;
assign w18644 = (w6052 & w2769) | (w6052 & w5601) | (w2769 & w5601);
assign w18645 = ~w12227 & ~w12074;
assign w18646 = ~w5944 & ~w8919;
assign w18647 = a_36 & a_56;
assign w18648 = ~w3145 & ~w1992;
assign w18649 = ~w2117 & ~w13746;
assign w18650 = (w10838 & w17728) | (w10838 & w9960) | (w17728 & w9960);
assign w18651 = (~w15399 & w14465) | (~w15399 & w8975) | (w14465 & w8975);
assign w18652 = w14122 & w3225;
assign w18653 = ~w11198 & ~w3286;
assign w18654 = ~w13948 & ~w7513;
assign w18655 = ~w8130 & ~w5353;
assign w18656 = w16151 & ~w16265;
assign w18657 = w14433 & ~w18167;
assign w18658 = ~w4653 & w3387;
assign w18659 = ~w6805 & ~w6199;
assign w18660 = ~w17121 & w15995;
assign w18661 = ~w10005 & ~w6632;
assign w18662 = (~w14854 & ~w9376) | (~w14854 & w10318) | (~w9376 & w10318);
assign w18663 = ~w9812 & ~w15333;
assign w18664 = ~w16551 & ~w2550;
assign w18665 = w16544 & ~w735;
assign w18666 = ~w9368 & ~w1716;
assign w18667 = ~w14375 & ~w6166;
assign w18668 = ~w3664 & ~w10185;
assign w18669 = w12671 & w7282;
assign w18670 = ~w10898 & ~w4277;
assign w18671 = ~w12909 & ~w15153;
assign w18672 = (~w780 & ~w2908) | (~w780 & w5322) | (~w2908 & w5322);
assign w18673 = ~w14585 & ~w16655;
assign w18674 = ~w3473 & ~w8200;
assign w18675 = w15911 & ~w8347;
assign w18676 = ~w6248 & w7077;
assign w18677 = w9843 & w19060;
assign w18678 = ~w7008 & ~w2452;
assign w18679 = ~w11232 & ~w7822;
assign w18680 = (~w14986 & w396) | (~w14986 & w12314) | (w396 & w12314);
assign w18681 = ~w12520 & ~w7511;
assign w18682 = (~w3769 & ~w14517) | (~w3769 & w13606) | (~w14517 & w13606);
assign w18683 = ~w9368 & ~w1286;
assign w18684 = w3966 & ~w17336;
assign w18685 = a_56 & a_57;
assign w18686 = w12096 & w1872;
assign w18687 = ~w17768 & ~w8020;
assign w18688 = a_34 & a_55;
assign w18689 = w18247 & ~w12599;
assign w18690 = a_7 & a_24;
assign w18691 = w8626 & w3615;
assign w18692 = ~w290 & ~w3316;
assign w18693 = ~w10216 & ~w7451;
assign w18694 = ~w16824 & ~w100;
assign w18695 = w3080 & ~w18687;
assign w18696 = ~w441 & w15727;
assign w18697 = ~w17488 & ~w3467;
assign w18698 = a_38 & a_45;
assign w18699 = ~w1648 & w10268;
assign w18700 = w18261 & w14798;
assign w18701 = ~w1776 & ~w18669;
assign w18702 = ~w1037 & ~w17154;
assign w18703 = ~w7160 & w15895;
assign w18704 = ~w316 & ~w677;
assign w18705 = ~w14057 & ~w16787;
assign w18706 = ~w6356 & w2537;
assign w18707 = w14171 & ~w2990;
assign w18708 = w3664 & w4471;
assign w18709 = w4700 & w5455;
assign w18710 = w19115 & ~w3291;
assign w18711 = a_40 & a_52;
assign w18712 = w17461 & ~w18576;
assign w18713 = ~w7102 & w15893;
assign w18714 = w6059 & w8418;
assign w18715 = a_4 & a_17;
assign w18716 = ~w14727 & ~w16763;
assign w18717 = w15630 & ~w16854;
assign w18718 = ~w8052 & w2211;
assign w18719 = ~w15661 & ~w16458;
assign w18720 = ~w17198 & ~w2581;
assign w18721 = w2620 & w17346;
assign w18722 = w16604 & ~w1517;
assign w18723 = a_13 & a_38;
assign w18724 = w13603 & ~w7038;
assign w18725 = w16249 & ~w16023;
assign w18726 = w13082 & w8008;
assign w18727 = ~w2900 & ~w8523;
assign w18728 = ~w6655 & ~w12574;
assign w18729 = ~w13408 & w2629;
assign w18730 = ~w12460 & w8951;
assign w18731 = a_12 & a_18;
assign w18732 = (~w14213 & ~w18188) | (~w14213 & w14555) | (~w18188 & w14555);
assign w18733 = ~w18017 & ~w1566;
assign w18734 = w16800 & w8181;
assign w18735 = ~w9813 & ~w12938;
assign w18736 = w2948 & w9043;
assign w18737 = a_23 & a_57;
assign w18738 = ~w9917 & ~w14784;
assign w18739 = a_20 & a_24;
assign w18740 = ~w13941 & ~w11481;
assign w18741 = w1320 & w4766;
assign w18742 = a_4 & a_59;
assign w18743 = ~w481 & ~w1670;
assign w18744 = ~w11719 & w7682;
assign w18745 = ~w16183 & ~w2132;
assign w18746 = ~w1901 & ~w3497;
assign w18747 = ~w5743 & w382;
assign w18748 = ~w4555 & ~w2259;
assign w18749 = ~w14131 & ~w4166;
assign w18750 = (~w10343 & ~w8631) | (~w10343 & w15405) | (~w8631 & w15405);
assign w18751 = w6887 & ~w10924;
assign w18752 = ~w15780 & ~w17587;
assign w18753 = a_10 & a_21;
assign w18754 = w10817 & w6216;
assign w18755 = w16394 & w3732;
assign w18756 = ~w1144 & w4993;
assign w18757 = ~w10330 & w9245;
assign w18758 = w17497 & ~w9749;
assign w18759 = w6899 & w14953;
assign w18760 = ~w17956 & ~w12523;
assign w18761 = w17065 & ~w16762;
assign w18762 = w16972 & w417;
assign w18763 = ~a_37 & ~w11203;
assign w18764 = ~w11514 & ~w15249;
assign w18765 = ~w12809 & ~w7527;
assign w18766 = ~w14983 & ~w15997;
assign w18767 = ~w3852 & ~w1604;
assign w18768 = w14414 & ~w17974;
assign w18769 = ~w11115 & ~w8930;
assign w18770 = ~w6626 & ~w2518;
assign w18771 = ~w11169 & ~w18995;
assign w18772 = (~w11446 & w11949) | (~w11446 & w5882) | (w11949 & w5882);
assign w18773 = ~w5741 & ~w6868;
assign w18774 = a_28 & a_37;
assign w18775 = ~w11773 & ~w4119;
assign w18776 = ~w12648 & ~w14155;
assign w18777 = (a_38 & w7488) | (a_38 & w18015) | (w7488 & w18015);
assign w18778 = w3757 & w10037;
assign w18779 = w9278 & ~w14796;
assign w18780 = ~w11157 & ~w12584;
assign w18781 = ~w1692 & ~w4807;
assign w18782 = ~w10936 & ~w1882;
assign w18783 = a_53 & a_55;
assign w18784 = ~w16069 & ~w15019;
assign w18785 = ~w10307 & ~w3039;
assign w18786 = a_3 & a_12;
assign w18787 = ~w4944 & w8151;
assign w18788 = w17811 & ~w1420;
assign w18789 = ~w15345 & w6667;
assign w18790 = ~w13486 & ~w2860;
assign w18791 = w15619 & ~w16656;
assign w18792 = w2797 & w9866;
assign w18793 = ~w9646 & ~w8260;
assign w18794 = a_0 & a_29;
assign w18795 = ~w15014 & ~w7968;
assign w18796 = w5512 & ~w5187;
assign w18797 = (~w8341 & w12897) | (~w8341 & w16711) | (w12897 & w16711);
assign w18798 = ~w3001 & ~w17679;
assign w18799 = ~w3418 & w386;
assign w18800 = w9390 & ~w17223;
assign w18801 = (w19083 & w2809) | (w19083 & w11676) | (w2809 & w11676);
assign w18802 = a_13 & a_49;
assign w18803 = w5087 & ~w4747;
assign w18804 = ~w16968 & ~w11108;
assign w18805 = ~w14746 & w14325;
assign w18806 = ~w5453 & ~w12319;
assign w18807 = ~w11044 & w5768;
assign w18808 = ~w935 & ~w6406;
assign w18809 = ~w4428 & ~w10641;
assign w18810 = ~w16733 & ~w18805;
assign w18811 = a_30 & a_33;
assign w18812 = w5754 & ~w8215;
assign w18813 = a_12 & a_61;
assign w18814 = a_34 & a_61;
assign w18815 = ~w4872 & w9164;
assign w18816 = w9603 & ~w2306;
assign w18817 = w8606 & ~w13532;
assign w18818 = ~w511 & w12533;
assign w18819 = (w19046 & w11644) | (w19046 & w14879) | (w11644 & w14879);
assign w18820 = ~w4056 & ~w6156;
assign w18821 = (w19005 & w13758) | (w19005 & w11327) | (w13758 & w11327);
assign w18822 = ~w1034 & ~w12843;
assign w18823 = ~w17553 & ~w16429;
assign w18824 = w933 & w14418;
assign w18825 = ~w2881 & w18152;
assign w18826 = w12060 & ~w16052;
assign w18827 = ~w12519 & ~w17572;
assign w18828 = a_19 & a_30;
assign w18829 = a_49 & a_56;
assign w18830 = w12606 & ~w2037;
assign w18831 = ~w3630 & ~w14601;
assign w18832 = ~w6662 & ~w3530;
assign w18833 = w11357 & ~w15241;
assign w18834 = ~w978 & w4660;
assign w18835 = w10516 & ~w6863;
assign w18836 = ~w109 & w11156;
assign w18837 = ~w5121 & ~w4021;
assign w18838 = a_19 & a_42;
assign w18839 = w2689 & ~w16818;
assign w18840 = ~w12128 & w2691;
assign w18841 = a_37 & a_46;
assign w18842 = (~w6834 & w6291) | (~w6834 & w16147) | (w6291 & w16147);
assign w18843 = ~w963 & w13186;
assign w18844 = w2080 & ~w4636;
assign w18845 = ~w18087 & ~w7581;
assign w18846 = w16398 & ~w17987;
assign w18847 = ~w12521 & ~w5293;
assign w18848 = (w2769 & w10622) | (w2769 & w3114) | (w10622 & w3114);
assign w18849 = w13030 & ~w14081;
assign w18850 = a_5 & a_62;
assign w18851 = ~w15471 & ~w16584;
assign w18852 = ~w14980 & ~w2508;
assign w18853 = w6426 & ~w10266;
assign w18854 = ~w14016 & ~w13772;
assign w18855 = ~w9605 & ~w6642;
assign w18856 = ~w10330 & w13002;
assign w18857 = ~w14961 & w17974;
assign w18858 = a_11 & a_61;
assign w18859 = a_11 & a_27;
assign w18860 = w7472 & w13613;
assign w18861 = w14127 & w19065;
assign w18862 = ~w17750 & ~w15967;
assign w18863 = ~w1811 & ~w18931;
assign w18864 = ~w6700 & ~w15175;
assign w18865 = ~a_38 & a_39;
assign w18866 = a_8 & a_52;
assign w18867 = ~w3382 & ~w2913;
assign w18868 = w6529 & ~w18056;
assign w18869 = w17428 & ~w12958;
assign w18870 = w6347 & w19194;
assign w18871 = ~w15108 & ~w1891;
assign w18872 = a_5 & a_63;
assign w18873 = ~w18588 & w7809;
assign w18874 = ~w272 & ~w5218;
assign w18875 = w4161 & ~w15210;
assign w18876 = ~w1234 & ~w4722;
assign w18877 = w3864 & ~w8864;
assign w18878 = ~w14047 & w4300;
assign w18879 = ~w10613 & w14556;
assign w18880 = w11306 & w1490;
assign w18881 = ~w10922 & ~w12407;
assign w18882 = a_9 & a_31;
assign w18883 = ~w5769 & ~w4388;
assign w18884 = ~w5710 & ~w11804;
assign w18885 = w2053 & w18173;
assign w18886 = w11081 & ~w17820;
assign w18887 = w5176 & ~w11590;
assign w18888 = ~w3334 & w14738;
assign w18889 = a_9 & a_16;
assign w18890 = w7863 & w17004;
assign w18891 = a_8 & a_59;
assign w18892 = w10302 & w4989;
assign w18893 = ~w15620 & ~w17682;
assign w18894 = w16174 & ~w14278;
assign w18895 = ~w8803 & w5240;
assign w18896 = a_42 & a_43;
assign w18897 = w13735 & w10297;
assign w18898 = a_10 & a_44;
assign w18899 = ~w2507 & ~w911;
assign w18900 = ~w3491 & ~w15700;
assign w18901 = ~w12893 & w9259;
assign w18902 = w2068 & w13432;
assign w18903 = ~w1941 & ~w806;
assign w18904 = ~w1548 & ~w15477;
assign w18905 = w13718 & w3833;
assign w18906 = ~w5014 & ~w18859;
assign w18907 = ~w8488 & w1112;
assign w18908 = a_29 & a_36;
assign w18909 = w7971 & w7677;
assign w18910 = ~w2113 & ~w7244;
assign w18911 = ~w14277 & ~w8907;
assign w18912 = ~w11711 & ~w13130;
assign w18913 = ~w13605 & w7118;
assign w18914 = w18820 & w6389;
assign w18915 = a_33 & a_58;
assign w18916 = ~w14755 & w1693;
assign w18917 = ~w13191 & ~w15817;
assign w18918 = ~w7593 & ~w4483;
assign w18919 = (w2093 & ~w13966) | (w2093 & w46) | (~w13966 & w46);
assign w18920 = ~w18112 & ~w16438;
assign w18921 = a_13 & a_26;
assign w18922 = ~w14645 & ~w14141;
assign w18923 = (a_48 & w8371) | (a_48 & w17190) | (w8371 & w17190);
assign w18924 = ~w1763 & ~w6280;
assign w18925 = w16254 & w313;
assign w18926 = w9297 & ~w17256;
assign w18927 = ~w1378 & ~w6252;
assign w18928 = ~w5183 & w17584;
assign w18929 = ~w13768 & w1503;
assign w18930 = w1170 & w13417;
assign w18931 = ~w13743 & ~w3788;
assign w18932 = ~w526 & ~w1735;
assign w18933 = w4327 & ~w15890;
assign w18934 = w8637 & ~w17546;
assign w18935 = ~w697 & ~w7480;
assign w18936 = ~w2135 & ~w7320;
assign w18937 = ~w8928 & ~w19003;
assign w18938 = ~w14122 & ~w3225;
assign w18939 = ~w5831 & ~w17187;
assign w18940 = ~w13647 & ~w13852;
assign w18941 = ~w4672 & ~w12472;
assign w18942 = ~w3243 & ~w8961;
assign w18943 = ~w1256 & ~w10237;
assign w18944 = w15511 & ~w15378;
assign w18945 = w9585 & ~w9556;
assign w18946 = ~w2450 & w18200;
assign w18947 = a_58 & a_59;
assign w18948 = ~w8475 & ~w4334;
assign w18949 = ~a_48 & w1031;
assign w18950 = a_6 & a_45;
assign w18951 = ~w10824 & w640;
assign w18952 = ~w18774 & ~w3398;
assign w18953 = a_44 & a_63;
assign w18954 = ~w14083 & ~w13660;
assign w18955 = w13082 & ~w1798;
assign w18956 = ~w1584 & ~w2294;
assign w18957 = w1719 & ~w2278;
assign w18958 = ~w14062 & ~w8908;
assign w18959 = ~w12654 & w13436;
assign w18960 = ~w7311 & ~w10658;
assign w18961 = (w5296 & w1962) | (w5296 & w14412) | (w1962 & w14412);
assign w18962 = ~w16931 & w8289;
assign w18963 = ~w1093 & ~w16042;
assign w18964 = w1956 & ~w17173;
assign w18965 = ~w18602 & ~w9063;
assign w18966 = w11271 & ~w9503;
assign w18967 = w8488 & ~w1112;
assign w18968 = w13834 & ~w5764;
assign w18969 = (~w1885 & ~w3826) | (~w1885 & w732) | (~w3826 & w732);
assign w18970 = ~w250 & ~w9421;
assign w18971 = (w10790 & w63) | (w10790 & w13658) | (w63 & w13658);
assign w18972 = w6420 & ~w14188;
assign w18973 = a_62 & w5133;
assign w18974 = ~w15251 & ~w8771;
assign w18975 = ~w8519 & ~w7863;
assign w18976 = w17231 & ~w16683;
assign w18977 = (~w3624 & w8747) | (~w3624 & w7708) | (w8747 & w7708);
assign w18978 = w5232 & ~w5379;
assign w18979 = ~w4096 & ~w4955;
assign w18980 = w14521 & w5113;
assign w18981 = w8763 & w6550;
assign w18982 = ~w12464 & w2614;
assign w18983 = w7484 & w13936;
assign w18984 = ~w5582 & ~w15951;
assign w18985 = a_24 & a_55;
assign w18986 = ~w17991 & ~w18184;
assign w18987 = ~w6315 & w1452;
assign w18988 = ~w8056 & ~w13622;
assign w18989 = w12268 & ~w15927;
assign w18990 = ~w2621 & ~w4057;
assign w18991 = ~w10350 & w1249;
assign w18992 = a_3 & a_49;
assign w18993 = ~w8522 & ~w8751;
assign w18994 = ~w3770 & ~w15614;
assign w18995 = ~w12786 & ~w11253;
assign w18996 = ~w11387 & ~w15756;
assign w18997 = a_43 & a_58;
assign w18998 = w5387 & ~w15855;
assign w18999 = ~w9388 & ~w3261;
assign w19000 = ~w1574 & w315;
assign w19001 = w16124 & ~w18202;
assign w19002 = ~w4269 & ~w16686;
assign w19003 = a_33 & a_44;
assign w19004 = a_12 & a_38;
assign w19005 = ~w7129 & w11884;
assign w19006 = ~w13065 & ~w2981;
assign w19007 = ~w5468 & ~w5875;
assign w19008 = (~w2769 & w7885) | (~w2769 & w12146) | (w7885 & w12146);
assign w19009 = a_1 & a_14;
assign w19010 = ~w16404 & w15087;
assign w19011 = ~w3052 & ~w9148;
assign w19012 = ~w2009 & ~w5122;
assign w19013 = w3800 & w17955;
assign w19014 = ~w14179 & ~w11055;
assign w19015 = w3009 & ~w15662;
assign w19016 = a_0 & a_52;
assign w19017 = a_38 & a_47;
assign w19018 = ~w13004 & ~w6231;
assign w19019 = ~w17356 & w2114;
assign w19020 = ~w16950 & ~w11757;
assign w19021 = ~w17670 & ~w3192;
assign w19022 = ~w9015 & ~w9225;
assign w19023 = a_45 & a_50;
assign w19024 = w3880 & ~w13476;
assign w19025 = (~w13917 & ~w6001) | (~w13917 & w9723) | (~w6001 & w9723);
assign w19026 = ~w567 & ~w14859;
assign w19027 = a_25 & a_37;
assign w19028 = ~w5590 & ~w13841;
assign w19029 = w18537 & w18841;
assign w19030 = (w2352 & w13945) | (w2352 & w19001) | (w13945 & w19001);
assign w19031 = w8765 & ~w7078;
assign w19032 = ~w19119 & ~w5413;
assign w19033 = (~w11421 & w16015) | (~w11421 & w7530) | (w16015 & w7530);
assign w19034 = w13853 & ~w17354;
assign w19035 = ~w3303 & w4901;
assign w19036 = ~w2769 & w7055;
assign w19037 = ~w9514 & w18932;
assign w19038 = ~w15650 & ~w5138;
assign w19039 = ~w16127 & w17817;
assign w19040 = ~w9911 & ~w3107;
assign w19041 = w6619 & w11423;
assign w19042 = w13061 & ~w18798;
assign w19043 = ~w6527 & w18486;
assign w19044 = ~w6485 & ~w6368;
assign w19045 = (w5410 & w2769) | (w5410 & w6776) | (w2769 & w6776);
assign w19046 = ~w18463 & ~w7805;
assign w19047 = ~w19123 & ~w11381;
assign w19048 = ~w17984 & ~w10166;
assign w19049 = ~w8876 & ~w12345;
assign w19050 = ~w17901 & ~w18136;
assign w19051 = ~w2405 & ~w7924;
assign w19052 = ~w6671 & ~w9444;
assign w19053 = ~w4375 & ~w8062;
assign w19054 = a_58 & a_62;
assign w19055 = a_39 & a_63;
assign w19056 = ~w7962 & w5565;
assign w19057 = ~w11139 & ~w3401;
assign w19058 = w15059 & w17256;
assign w19059 = ~w2626 & w17575;
assign w19060 = a_5 & a_8;
assign w19061 = w12717 & w4756;
assign w19062 = ~w5102 & ~w18043;
assign w19063 = ~w13624 & ~w14824;
assign w19064 = ~w18533 & ~w14227;
assign w19065 = a_1 & a_4;
assign w19066 = ~w1888 & w8615;
assign w19067 = w15252 & ~w8721;
assign w19068 = ~w7588 & ~w7442;
assign w19069 = a_8 & a_61;
assign w19070 = (~w14260 & ~w1773) | (~w14260 & w3747) | (~w1773 & w3747);
assign w19071 = ~w10029 & w17744;
assign w19072 = ~w5335 & w16743;
assign w19073 = ~w12586 & ~w1614;
assign w19074 = w15273 & ~w14903;
assign w19075 = ~w2386 & ~w6676;
assign w19076 = ~w402 & ~w13289;
assign w19077 = ~w9917 & ~w3267;
assign w19078 = ~w13463 & ~w16477;
assign w19079 = ~w18710 & ~w12644;
assign w19080 = w17645 & ~w13293;
assign w19081 = w16725 & w7745;
assign w19082 = ~w1141 & ~w18581;
assign w19083 = ~w18957 & ~w9699;
assign w19084 = ~w2757 & ~w12516;
assign w19085 = ~w12237 & ~w11610;
assign w19086 = ~w6799 & ~w6456;
assign w19087 = ~w5999 & ~w16687;
assign w19088 = w870 & w7104;
assign w19089 = ~w2762 & ~w14019;
assign w19090 = (w11782 & w14374) | (w11782 & w17796) | (w14374 & w17796);
assign w19091 = w11914 & w7604;
assign w19092 = ~w8041 & ~w1734;
assign w19093 = ~w6003 & ~w7241;
assign w19094 = w16681 & ~w1805;
assign w19095 = (a_59 & w18558) | (a_59 & w18947) | (w18558 & w18947);
assign w19096 = (~w7341 & w10046) | (~w7341 & w540) | (w10046 & w540);
assign w19097 = ~w16124 & w18202;
assign w19098 = a_34 & a_37;
assign w19099 = ~w8060 & w12295;
assign w19100 = ~w4114 & ~w9454;
assign w19101 = ~w16390 & ~w16046;
assign w19102 = ~w7129 & w12602;
assign w19103 = w11879 & ~w6238;
assign w19104 = w17856 & w15051;
assign w19105 = w12640 & ~w4006;
assign w19106 = ~w10620 & w3881;
assign w19107 = (w2352 & ~w13979) | (w2352 & w6197) | (~w13979 & w6197);
assign w19108 = w786 & w12761;
assign w19109 = w15199 & ~w13163;
assign w19110 = ~w17296 & ~w34;
assign w19111 = ~w10435 & ~w13066;
assign w19112 = ~w1009 & ~w7785;
assign w19113 = ~w6742 & ~w768;
assign w19114 = ~w537 & ~w4587;
assign w19115 = a_18 & a_43;
assign w19116 = w2960 & w11408;
assign w19117 = ~w3516 & w17342;
assign w19118 = w6101 & ~w11981;
assign w19119 = ~w13219 & ~w15077;
assign w19120 = ~w8637 & w17546;
assign w19121 = w11166 & ~w5886;
assign w19122 = ~w13988 & ~w5000;
assign w19123 = w6311 & w864;
assign w19124 = (w16917 & w13786) | (w16917 & w6493) | (w13786 & w6493);
assign w19125 = w13011 & w11600;
assign w19126 = ~w2820 & ~w6694;
assign w19127 = ~w16111 & ~w14011;
assign w19128 = a_10 & a_47;
assign w19129 = ~a_37 & a_38;
assign w19130 = (~w6897 & w17141) | (~w6897 & w2366) | (w17141 & w2366);
assign w19131 = w14904 & ~w14267;
assign w19132 = (w15399 & w17089) | (w15399 & w2914) | (w17089 & w2914);
assign w19133 = (~w10549 & ~w15595) | (~w10549 & w654) | (~w15595 & w654);
assign w19134 = ~w12460 & ~w113;
assign w19135 = w18969 & ~w17495;
assign w19136 = ~w1367 & ~w15599;
assign w19137 = ~w12229 & w4102;
assign w19138 = ~w11756 & ~w16115;
assign w19139 = ~w12609 & ~w14406;
assign w19140 = ~w4905 & ~w12819;
assign w19141 = a_6 & a_20;
assign w19142 = ~w10632 & ~w2738;
assign w19143 = ~w3948 & ~w15550;
assign w19144 = ~w13404 & w14695;
assign w19145 = ~w14646 & ~w15691;
assign w19146 = (~w1225 & ~w5939) | (~w1225 & ~w16917) | (~w5939 & ~w16917);
assign w19147 = (~w4075 & ~w16661) | (~w4075 & ~w15988) | (~w16661 & ~w15988);
assign w19148 = (w410 & ~w14460) | (w410 & ~w13603) | (~w14460 & ~w13603);
assign w19149 = (~w7612 & ~w19001) | (~w7612 & ~w152) | (~w19001 & ~w152);
assign w19150 = (w1606 & ~w3640) | (w1606 & ~w3601) | (~w3640 & ~w3601);
assign w19151 = (w13938 & ~w240) | (w13938 & ~w1894) | (~w240 & ~w1894);
assign w19152 = (w14532 & ~w668) | (w14532 & ~w7102) | (~w668 & ~w7102);
assign w19153 = ~w16410 | w896;
assign w19154 = (w2508 & ~w11585) | (w2508 & ~w7268) | (~w11585 & ~w7268);
assign w19155 = (w2433 & ~w5464) | (w2433 & ~w15988) | (~w5464 & ~w15988);
assign w19156 = (w17910 & ~w5720) | (w17910 & ~w5495) | (~w5720 & ~w5495);
assign w19157 = (w11320 & ~w17236) | (w11320 & ~w1648) | (~w17236 & ~w1648);
assign w19158 = (w1956 & ~w15928) | (w1956 & ~w7768) | (~w15928 & ~w7768);
assign w19159 = w1621 & w14087;
assign w19160 = (~w3695 & ~w4420) | (~w3695 & w3417) | (~w4420 & w3417);
assign w19161 = (w8436 & ~w7759) | (w8436 & ~w12095) | (~w7759 & ~w12095);
assign w19162 = (~w18272 & w16086) | (~w18272 & w15356) | (w16086 & w15356);
assign w19163 = (w18967 & ~w9065) | (w18967 & ~w3182) | (~w9065 & ~w3182);
assign w19164 = (~w1558 & ~w10349) | (~w1558 & ~w7768) | (~w10349 & ~w7768);
assign w19165 = (w8678 & ~w12297) | (w8678 & w18017) | (~w12297 & w18017);
assign w19166 = (w9291 & ~w17981) | (w9291 & ~w6775) | (~w17981 & ~w6775);
assign w19167 = (~w10459 & w10970) | (~w10459 & ~w15415) | (w10970 & ~w15415);
assign w19168 = (w896 & ~w16410) | (w896 & ~w12887) | (~w16410 & ~w12887);
assign w19169 = (~w1786 & w9641) | (~w1786 & ~w7341) | (w9641 & ~w7341);
assign w19170 = w8080 & w19196;
assign w19171 = (w12440 & ~w10073) | (w12440 & ~w10390) | (~w10073 & ~w10390);
assign w19172 = (~w16370 & w2143) | (~w16370 & ~w18365) | (w2143 & ~w18365);
assign w19173 = (~w13059 & w7544) | (~w13059 & w9252) | (w7544 & w9252);
assign w19174 = w7544 & ~w13059;
assign w19175 = ~w12297 | w8678;
assign w19176 = (w6734 & ~w1468) | (w6734 & ~w6475) | (~w1468 & ~w6475);
assign w19177 = (~w8983 & ~w13422) | (~w8983 & ~w18017) | (~w13422 & ~w18017);
assign w19178 = (~w11270 & w7772) | (~w11270 & ~w5527) | (w7772 & ~w5527);
assign w19179 = (~w1838 & w16256) | (~w1838 & ~w11864) | (w16256 & ~w11864);
assign w19180 = (w2960 & ~w4170) | (w2960 & ~w9337) | (~w4170 & ~w9337);
assign w19181 = ~w10382 | w1876;
assign w19182 = (~w832 & ~w12040) | (~w832 & ~w18357) | (~w12040 & ~w18357);
assign w19183 = (w1876 & ~w10382) | (w1876 & ~w195) | (~w10382 & ~w195);
assign w19184 = (~w16711 & ~w6956) | (~w16711 & ~w7768) | (~w6956 & ~w7768);
assign w19185 = (w2977 & ~w12513) | (w2977 & ~w14792) | (~w12513 & ~w14792);
assign w19186 = (w262 & ~w6242) | (w262 & ~w18091) | (~w6242 & ~w18091);
assign w19187 = (~w6832 & w10946) | (~w6832 & ~w7341) | (w10946 & ~w7341);
assign w19188 = (~w18272 & ~w4312) | (~w18272 & w7886) | (~w4312 & w7886);
assign w19189 = (w10544 & w17770) | (w10544 & ~w13280) | (w17770 & ~w13280);
assign w19190 = (w7341 & ~w18431) | (w7341 & ~w2769) | (~w18431 & ~w2769);
assign w19191 = (~w13059 & w7544) | (~w13059 & w18357) | (w7544 & w18357);
assign w19192 = (w994 & ~w10231) | (w994 & ~w1728) | (~w10231 & ~w1728);
assign w19193 = (~w4275 & ~w14432) | (~w4275 & ~w7768) | (~w14432 & ~w7768);
assign w19194 = (~w983 & ~w16671) | (~w983 & ~w7102) | (~w16671 & ~w7102);
assign w19195 = w10385 & ~w14429;
assign w19196 = (~w8836 & ~w8122) | (~w8836 & ~w17914) | (~w8122 & ~w17914);
assign w19197 = (~w896 & w16410) | (~w896 & w742) | (w16410 & w742);
assign w19198 = (~w11733 & w19177) | (~w11733 & ~w1566) | (w19177 & ~w1566);
assign w19199 = (w19192 & w994) | (w19192 & ~w12904) | (w994 & ~w12904);
assign w19200 = (w10385 & w19195) | (w10385 & w1074) | (w19195 & w1074);
assign one = 1;
assign asquared_0 = a_0;// level 0
assign asquared_1 = ~one;// level 0
assign asquared_2 = w255;// level 1
assign asquared_3 = w14416;// level 3
assign asquared_4 = w5326;// level 4
assign asquared_5 = w12017;// level 7
assign asquared_6 = w2605;// level 7
assign asquared_7 = w10700;// level 9
assign asquared_8 = w17845;// level 11
assign asquared_9 = ~w10512;// level 12
assign asquared_10 = w2112;// level 14
assign asquared_11 = ~w13376;// level 15
assign asquared_12 = w18948;// level 16
assign asquared_13 = w11276;// level 17
assign asquared_14 = w8667;// level 17
assign asquared_15 = ~w7083;// level 18
assign asquared_16 = w10778;// level 19
assign asquared_17 = ~w4678;// level 20
assign asquared_18 = w12409;// level 20
assign asquared_19 = ~w12948;// level 21
assign asquared_20 = w18621;// level 21
assign asquared_21 = w12140;// level 22
assign asquared_22 = w14748;// level 22
assign asquared_23 = ~w3865;// level 23
assign asquared_24 = w9229;// level 23
assign asquared_25 = w4076;// level 24
assign asquared_26 = w7620;// level 24
assign asquared_27 = w2194;// level 24
assign asquared_28 = ~w18077;// level 25
assign asquared_29 = w12004;// level 26
assign asquared_30 = w13069;// level 25
assign asquared_31 = w16937;// level 26
assign asquared_32 = w14501;// level 26
assign asquared_33 = w15365;// level 26
assign asquared_34 = ~w17590;// level 28
assign asquared_35 = ~w18409;// level 27
assign asquared_36 = ~w18481;// level 28
assign asquared_37 = w6664;// level 29
assign asquared_38 = w5284;// level 30
assign asquared_39 = w3899;// level 29
assign asquared_40 = w51;// level 29
assign asquared_41 = ~w15326;// level 29
assign asquared_42 = w3132;// level 30
assign asquared_43 = w3435;// level 29
assign asquared_44 = w19040;// level 30
assign asquared_45 = w13097;// level 30
assign asquared_46 = ~w7936;// level 30
assign asquared_47 = w9792;// level 31
assign asquared_48 = w6850;// level 30
assign asquared_49 = w704;// level 30
assign asquared_50 = ~w17074;// level 32
assign asquared_51 = w13251;// level 33
assign asquared_52 = w2301;// level 32
assign asquared_53 = w10543;// level 33
assign asquared_54 = ~w17651;// level 32
assign asquared_55 = w11225;// level 33
assign asquared_56 = w4204;// level 34
assign asquared_57 = w1947;// level 33
assign asquared_58 = w9385;// level 33
assign asquared_59 = ~w12507;// level 33
assign asquared_60 = w166;// level 33
assign asquared_61 = w13467;// level 33
assign asquared_62 = w6040;// level 34
assign asquared_63 = ~w5252;// level 34
assign asquared_64 = w16210;// level 35
assign asquared_65 = w7421;// level 35
assign asquared_66 = w2214;// level 34
assign asquared_67 = w6464;// level 35
assign asquared_68 = ~w16080;// level 34
assign asquared_69 = w4;// level 35
assign asquared_70 = ~w10583;// level 36
assign asquared_71 = ~w17271;// level 35
assign asquared_72 = w17902;// level 35
assign asquared_73 = w4249;// level 35
assign asquared_74 = ~w17519;// level 35
assign asquared_75 = w9361;// level 35
assign asquared_76 = w6303;// level 35
assign asquared_77 = ~w8259;// level 35
assign asquared_78 = ~w18163;// level 36
assign asquared_79 = ~w1741;// level 36
assign asquared_80 = ~w12570;// level 35
assign asquared_81 = w7383;// level 35
assign asquared_82 = w17577;// level 35
assign asquared_83 = w14045;// level 35
assign asquared_84 = w7402;// level 35
assign asquared_85 = ~w1346;// level 35
assign asquared_86 = ~w15392;// level 36
assign asquared_87 = ~w8495;// level 35
assign asquared_88 = w16348;// level 36
assign asquared_89 = ~w9408;// level 35
assign asquared_90 = w2032;// level 35
assign asquared_91 = ~w11213;// level 35
assign asquared_92 = w2632;// level 36
assign asquared_93 = w9149;// level 36
assign asquared_94 = w10876;// level 36
assign asquared_95 = ~w16627;// level 35
assign asquared_96 = w17120;// level 35
assign asquared_97 = ~w16068;// level 36
assign asquared_98 = w12962;// level 36
assign asquared_99 = ~w9186;// level 36
assign asquared_100 = ~w4737;// level 36
assign asquared_101 = w18855;// level 36
assign asquared_102 = ~w6298;// level 36
assign asquared_103 = w8388;// level 36
assign asquared_104 = w7752;// level 36
assign asquared_105 = w9000;// level 36
assign asquared_106 = ~w12424;// level 36
assign asquared_107 = w9655;// level 36
assign asquared_108 = w15309;// level 36
assign asquared_109 = w9845;// level 36
assign asquared_110 = w9895;// level 36
assign asquared_111 = ~w6281;// level 36
assign asquared_112 = w3662;// level 36
assign asquared_113 = w389;// level 36
assign asquared_114 = ~w6120;// level 36
assign asquared_115 = w11553;// level 36
assign asquared_116 = ~w8136;// level 36
assign asquared_117 = w3963;// level 36
assign asquared_118 = ~w1630;// level 36
assign asquared_119 = ~w18088;// level 36
assign asquared_120 = w16566;// level 36
assign asquared_121 = ~w18879;// level 36
assign asquared_122 = ~w17563;// level 36
assign asquared_123 = ~w14661;// level 36
assign asquared_124 = w7231;// level 36
assign asquared_125 = ~w3885;// level 36
assign asquared_126 = ~w13690;// level 36
assign asquared_127 = w7867;// level 36
endmodule

// written by CirKit Wed Nov  2 14:26:17 2016

module router_best_speed.blif_ (
        pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, 
        po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112;
assign w0 = ~pi05 & ~pi06;
assign w1 = ~pi07 & ~pi08;
assign w2 = w0 & w1;
assign w3 = ~pi01 & ~pi02;
assign w4 = ~pi03 & ~pi04;
assign w5 = w3 & w4;
assign w6 = w2 & w5;
assign w7 = pi09 & ~w6;
assign w8 = ~pi12 & ~pi13;
assign w9 = pi14 & pi15;
assign w10 = ~w8 & w9;
assign w11 = ~pi16 & ~pi18;
assign w12 = ~w10 & w11;
assign w13 = ~pi10 & ~pi21;
assign w14 = ~pi22 & w13;
assign w15 = w12 & w14;
assign w16 = ~w7 & w15;
assign w17 = pi23 & pi24;
assign w18 = pi25 & pi27;
assign w19 = w17 & w18;
assign w20 = pi28 & pi29;
assign w21 = w19 & w20;
assign w22 = ~pi17 & ~pi18;
assign w23 = pi19 & pi20;
assign w24 = ~w22 & w23;
assign w25 = pi11 & pi14;
assign w26 = pi15 & w25;
assign w27 = w24 & w26;
assign w28 = (~w12 & w24) | (~w12 & w27) | (w24 & w27);
assign w29 = ~pi21 & ~pi22;
assign w30 = w20 & ~w29;
assign w31 = w19 & w30;
assign w32 = (w21 & w28) | (w21 & w31) | (w28 & w31);
assign w33 = w16 & w32;
assign w34 = pi03 & pi04;
assign w35 = pi05 & pi06;
assign w36 = w34 & w35;
assign w37 = pi07 & pi08;
assign w38 = pi02 & w37;
assign w39 = w36 & w38;
assign w40 = pi00 & pi01;
assign w41 = ~pi09 & ~w40;
assign w42 = (~pi09 & ~w39) | (~pi09 & w41) | (~w39 & w41);
assign w43 = ~pi26 & ~w42;
assign w44 = w33 & w43;
assign w45 = pi58 & pi59;
assign w46 = pi09 & pi57;
assign w47 = w45 & w46;
assign w48 = (pi57 & w40) | (pi57 & w46) | (w40 & w46);
assign w49 = w45 & w48;
assign w50 = (w39 & w47) | (w39 & w49) | (w47 & w49);
assign w51 = ~pi41 & ~pi42;
assign w52 = pi43 & pi55;
assign w53 = (pi55 & ~w51) | (pi55 & w52) | (~w51 & w52);
assign w54 = pi53 & pi54;
assign w55 = pi44 & w54;
assign w56 = w53 & w55;
assign w57 = pi45 & pi47;
assign w58 = pi49 & pi50;
assign w59 = w57 & w58;
assign w60 = w56 & w59;
assign w61 = ~pi35 & ~pi36;
assign w62 = ~pi37 & ~pi38;
assign w63 = w61 & w62;
assign w64 = ~pi30 & w63;
assign w65 = ~pi31 & ~pi32;
assign w66 = ~pi33 & ~pi34;
assign w67 = w65 & w66;
assign w68 = ~pi00 & w67;
assign w69 = w64 & w68;
assign w70 = pi39 & ~w69;
assign w71 = ~pi40 & ~pi42;
assign w72 = ~pi43 & w71;
assign w73 = pi33 & pi34;
assign w74 = pi35 & pi36;
assign w75 = w73 & w74;
assign w76 = pi37 & pi38;
assign w77 = ~pi00 & w76;
assign w78 = w75 & w77;
assign w79 = pi31 & pi32;
assign w80 = pi30 & w79;
assign w81 = w72 & ~w80;
assign w82 = (w72 & ~w78) | (w72 & w81) | (~w78 & w81);
assign w83 = w60 & ~w82;
assign w84 = (w60 & w70) | (w60 & w83) | (w70 & w83);
assign w85 = ~pi51 & ~pi52;
assign w86 = pi46 & pi47;
assign w87 = pi48 & pi50;
assign w88 = (pi50 & w86) | (pi50 & w87) | (w86 & w87);
assign w89 = ~pi49 & w85;
assign w90 = (w85 & ~w88) | (w85 & w89) | (~w88 & w89);
assign w91 = ~pi55 & ~pi56;
assign w92 = (~pi56 & ~w54) | (~pi56 & w91) | (~w54 & w91);
assign w93 = (~pi56 & w90) | (~pi56 & w92) | (w90 & w92);
assign w94 = w50 & ~w93;
assign w95 = (w50 & w84) | (w50 & w94) | (w84 & w94);
assign w96 = ~w16 & w32;
assign w97 = (w32 & w95) | (w32 & w96) | (w95 & w96);
assign w98 = pi26 & pi27;
assign w99 = w20 & w98;
assign w100 = ~w97 & ~w99;
assign w101 = w63 & w67;
assign w102 = ~pi39 & w72;
assign w103 = pi00 & pi30;
assign w104 = pi39 & w103;
assign w105 = w72 & ~w104;
assign w106 = (w101 & w102) | (w101 & w105) | (w102 & w105);
assign w107 = w60 & ~w106;
assign w108 = pi59 & ~w93;
assign w109 = (pi59 & w107) | (pi59 & w108) | (w107 & w108);
assign w110 = pi57 & pi58;
assign w111 = w109 & w110;
assign w112 = w44 & w111;
assign one = 1;
assign po00 = ~w44;
assign po01 = w100;
assign po02 = w112;
assign po03 = ~one;
assign po04 = ~one;
assign po05 = ~one;
assign po06 = ~one;
assign po07 = ~one;
assign po08 = ~one;
assign po09 = ~one;
assign po10 = ~one;
assign po11 = ~one;
assign po12 = ~one;
assign po13 = ~one;
assign po14 = ~one;
assign po15 = ~one;
assign po16 = ~one;
assign po17 = ~one;
assign po18 = ~one;
assign po19 = ~one;
assign po20 = ~one;
assign po21 = ~one;
assign po22 = ~one;
assign po23 = ~one;
assign po24 = ~one;
assign po25 = ~one;
assign po26 = ~one;
assign po27 = ~one;
assign po28 = ~one;
assign po29 = ~one;
endmodule

// Benchmark "apex6" written by ABC on Sun Apr 22 21:42:57 2018

module apex6 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83,
    po84, po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95,
    po96, po97, po98  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82,
    po83, po84, po85, po86, po87, po88, po89, po90, po91, po92, po93, po94,
    po95, po96, po97, po98;
  wire n236, n237, n238, n239, n240, n241, n242, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n288, n289, n291, n292, n293, n294, n295, n297, n298, n300,
    n301, n303, n304, n306, n307, n309, n310, n312, n313, n315, n316, n318,
    n319, n320, n321, n322, n324, n325, n327, n328, n330, n331, n333, n334,
    n336, n337, n339, n340, n342, n343, n345, n346, n347, n348, n349, n351,
    n352, n354, n355, n357, n358, n360, n361, n363, n364, n366, n367, n369,
    n370, n372, n373, n374, n375, n376, n378, n379, n381, n382, n384, n385,
    n387, n388, n390, n391, n393, n394, n396, n397, n399, n400, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n459, n460, n461, n462, n463, n464, n465, n467,
    n468, n469, n470, n471, n472, n474, n475, n476, n477, n478, n481, n482,
    n483, n484, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n531, n532,
    n533, n534, n535, n536, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n563, n564, n565, n566, n567, n568, n569, n570, n572,
    n573, n574, n576, n577, n578, n579, n580, n582, n583, n584, n585, n586,
    n587, n589, n590, n591, n592, n593, n595, n596, n597, n598, n599, n600,
    n602, n603, n604, n605, n606, n608, n609, n610, n611, n613, n614, n615,
    n616, n617, n619, n620, n622, n623, n625, n626, n628, n629, n631, n632,
    n634, n635, n637, n638, n640, n641, n642, n643, n644, n646, n647, n649,
    n650, n652, n653, n655, n656, n658, n659, n661, n662, n664, n665, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n833, n834, n835, n836, n837, n838,
    n839, n841, n842, n844, n845, n846, n847, n848, n850, n851, n852, n853,
    n854, n856, n857, n858, n859, n860, n861, n863, n864, n865, n866, n868,
    n869, n870, n871, n873, n874, n875, n876, n877, n878, n879, n881, n882,
    n883, n884, n885, n886, n887, n889, n890, n891, n892;
  assign po00 = ~pi072 | pi075;
  assign n236 = ~pi002 & ~pi003;
  assign n237 = ~pi072 & pi091;
  assign n238 = pi092 & n237;
  assign n239 = pi083 & n238;
  assign n240 = ~pi039 & ~n239;
  assign n241 = n236 & ~n240;
  assign n242 = ~pi001 & n241;
  assign po01 = pi073 | n242;
  assign n244 = pi034 & pi086;
  assign n245 = pi035 & ~pi086;
  assign n246 = ~n244 & ~n245;
  assign n247 = pi033 & ~pi086;
  assign n248 = pi032 & pi086;
  assign n249 = ~n247 & ~n248;
  assign n250 = pi088 & ~n249;
  assign n251 = ~pi087 & n250;
  assign n252 = ~pi088 & ~n246;
  assign n253 = pi087 & n252;
  assign n254 = ~n251 & ~n253;
  assign n255 = pi028 & ~pi091;
  assign n256 = ~pi074 & pi091;
  assign n257 = ~n255 & ~n256;
  assign n258 = pi092 & ~n257;
  assign n259 = pi091 & ~pi092;
  assign n260 = ~pi027 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = ~pi084 & ~pi085;
  assign n263 = ~pi091 & ~pi092;
  assign n264 = pi083 & ~n263;
  assign n265 = pi083 & ~n261;
  assign n266 = pi109 & ~n264;
  assign n267 = ~n262 & n266;
  assign n268 = ~n265 & ~n267;
  assign n269 = n262 & ~n264;
  assign n270 = ~pi075 & n269;
  assign n271 = po00 & ~n270;
  assign n272 = pi079 & ~pi080;
  assign n273 = ~pi028 & n272;
  assign n274 = ~pi079 & pi080;
  assign n275 = pi028 & n274;
  assign n276 = ~n273 & ~n275;
  assign n277 = pi037 & ~n276;
  assign n278 = pi075 & n277;
  assign n279 = ~pi072 & ~n268;
  assign n280 = ~pi075 & n279;
  assign n281 = ~pi089 & ~n254;
  assign n282 = ~pi090 & ~n271;
  assign n283 = n281 & n282;
  assign n284 = ~n280 & ~n283;
  assign n285 = ~n278 & n284;
  assign po02 = ~pi073 & ~n285;
  assign po45 = ~pi038 & pi082;
  assign n288 = pi081 & po45;
  assign n289 = ~pi038 & pi077;
  assign po03 = n288 | n289;
  assign n291 = pi007 & ~pi016;
  assign n292 = ~pi073 & ~n291;
  assign n293 = ~pi073 & n291;
  assign n294 = pi040 & n292;
  assign n295 = pi008 & n293;
  assign po04 = n294 | n295;
  assign n297 = pi041 & n292;
  assign n298 = pi009 & n293;
  assign po05 = n297 | n298;
  assign n300 = pi042 & n292;
  assign n301 = pi010 & n293;
  assign po06 = n300 | n301;
  assign n303 = pi043 & n292;
  assign n304 = pi011 & n293;
  assign po07 = n303 | n304;
  assign n306 = pi044 & n292;
  assign n307 = pi012 & n293;
  assign po08 = n306 | n307;
  assign n309 = pi045 & n292;
  assign n310 = pi013 & n293;
  assign po09 = n309 | n310;
  assign n312 = pi046 & n292;
  assign n313 = pi014 & n293;
  assign po10 = n312 | n313;
  assign n315 = pi047 & n292;
  assign n316 = pi015 & n293;
  assign po11 = n315 | n316;
  assign n318 = pi007 & pi016;
  assign n319 = ~pi073 & ~n318;
  assign n320 = ~pi073 & n318;
  assign n321 = pi048 & n319;
  assign n322 = pi008 & n320;
  assign po12 = n321 | n322;
  assign n324 = pi049 & n319;
  assign n325 = pi009 & n320;
  assign po13 = n324 | n325;
  assign n327 = pi050 & n319;
  assign n328 = pi010 & n320;
  assign po14 = n327 | n328;
  assign n330 = pi051 & n319;
  assign n331 = pi011 & n320;
  assign po15 = n330 | n331;
  assign n333 = pi052 & n319;
  assign n334 = pi012 & n320;
  assign po16 = n333 | n334;
  assign n336 = pi053 & n319;
  assign n337 = pi013 & n320;
  assign po17 = n336 | n337;
  assign n339 = pi054 & n319;
  assign n340 = pi014 & n320;
  assign po18 = n339 | n340;
  assign n342 = pi055 & n319;
  assign n343 = pi015 & n320;
  assign po19 = n342 | n343;
  assign n345 = pi017 & ~pi026;
  assign n346 = ~pi073 & ~n345;
  assign n347 = ~pi073 & n345;
  assign n348 = pi056 & n346;
  assign n349 = pi018 & n347;
  assign po20 = n348 | n349;
  assign n351 = pi057 & n346;
  assign n352 = pi019 & n347;
  assign po21 = n351 | n352;
  assign n354 = pi058 & n346;
  assign n355 = pi020 & n347;
  assign po22 = n354 | n355;
  assign n357 = pi059 & n346;
  assign n358 = pi021 & n347;
  assign po23 = n357 | n358;
  assign n360 = pi060 & n346;
  assign n361 = pi022 & n347;
  assign po24 = n360 | n361;
  assign n363 = pi061 & n346;
  assign n364 = pi023 & n347;
  assign po25 = n363 | n364;
  assign n366 = pi062 & n346;
  assign n367 = pi024 & n347;
  assign po26 = n366 | n367;
  assign n369 = pi063 & n346;
  assign n370 = pi025 & n347;
  assign po27 = n369 | n370;
  assign n372 = pi017 & pi026;
  assign n373 = ~pi073 & ~n372;
  assign n374 = ~pi073 & n372;
  assign n375 = pi064 & n373;
  assign n376 = pi018 & n374;
  assign po28 = n375 | n376;
  assign n378 = pi065 & n373;
  assign n379 = pi019 & n374;
  assign po29 = n378 | n379;
  assign n381 = pi066 & n373;
  assign n382 = pi020 & n374;
  assign po30 = n381 | n382;
  assign n384 = pi067 & n373;
  assign n385 = pi021 & n374;
  assign po31 = n384 | n385;
  assign n387 = pi068 & n373;
  assign n388 = pi022 & n374;
  assign po32 = n387 | n388;
  assign n390 = pi069 & n373;
  assign n391 = pi023 & n374;
  assign po33 = n390 | n391;
  assign n393 = pi070 & n373;
  assign n394 = pi024 & n374;
  assign po34 = n393 | n394;
  assign n396 = pi071 & n373;
  assign n397 = pi025 & n374;
  assign po35 = n396 | n397;
  assign n399 = ~pi001 & pi072;
  assign n400 = n236 & n399;
  assign po36 = pi073 | n400;
  assign po37 = pi038 | n239;
  assign n403 = pi109 & ~n262;
  assign n404 = ~pi090 & ~n254;
  assign n405 = ~pi089 & n262;
  assign n406 = n404 & n405;
  assign n407 = ~n403 & ~n406;
  assign n408 = pi028 & pi092;
  assign n409 = ~pi027 & pi091;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~pi028 & pi092;
  assign n412 = pi027 & pi091;
  assign n413 = ~n411 & ~n412;
  assign n414 = pi074 & ~n413;
  assign n415 = ~pi072 & ~pi074;
  assign n416 = ~n410 & n415;
  assign n417 = ~n414 & ~n416;
  assign n418 = ~n238 & n417;
  assign n419 = ~n264 & n407;
  assign n420 = ~pi072 & ~n419;
  assign n421 = pi074 & ~n420;
  assign n422 = pi083 & ~n418;
  assign n423 = ~n264 & ~n407;
  assign n424 = n415 & n423;
  assign n425 = ~n422 & ~n424;
  assign n426 = ~n421 & n425;
  assign po38 = ~pi073 & ~n426;
  assign n428 = pi079 & pi080;
  assign n429 = pi036 & pi078;
  assign n430 = ~pi034 & ~pi035;
  assign n431 = n429 & n430;
  assign n432 = pi126 & pi127;
  assign n433 = pi125 & pi128;
  assign n434 = n432 & n433;
  assign n435 = ~pi035 & ~pi133;
  assign n436 = pi035 & pi133;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~pi034 & ~pi132;
  assign n439 = pi034 & pi132;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n437 & ~n440;
  assign n442 = ~pi033 & ~pi131;
  assign n443 = pi033 & pi131;
  assign n444 = ~n442 & ~n443;
  assign n445 = ~pi032 & pi130;
  assign n446 = pi032 & ~pi130;
  assign n447 = ~n445 & ~n446;
  assign n448 = pi129 & pi134;
  assign n449 = n434 & n448;
  assign n450 = n441 & n449;
  assign n451 = ~n444 & n450;
  assign n452 = ~n447 & n451;
  assign n453 = pi075 & ~n428;
  assign n454 = ~pi033 & n431;
  assign n455 = ~pi032 & n454;
  assign n456 = ~n453 & ~n455;
  assign n457 = ~n452 & n456;
  assign po39 = ~pi073 & ~n457;
  assign n459 = pi128 & pi129;
  assign n460 = n432 & n459;
  assign n461 = ~pi133 & n460;
  assign n462 = pi130 & ~pi131;
  assign n463 = ~pi132 & n462;
  assign n464 = n461 & n463;
  assign n465 = ~pi036 & ~pi038;
  assign po89 = ~pi125 & n465;
  assign n467 = ~n464 & n465;
  assign n468 = ~po89 & ~n467;
  assign n469 = pi125 & n465;
  assign n470 = pi076 & ~n468;
  assign n471 = n464 & n469;
  assign n472 = ~pi076 & n471;
  assign po40 = n470 | n472;
  assign n474 = ~pi076 & n465;
  assign n475 = n468 & ~n474;
  assign n476 = pi077 & ~n475;
  assign n477 = pi076 & ~pi077;
  assign n478 = n471 & n477;
  assign po41 = n476 | n478;
  assign po46 = pi036 & ~pi038;
  assign n481 = ~pi038 & pi078;
  assign n482 = ~po46 & ~n481;
  assign n483 = pi081 & pi082;
  assign n484 = pi000 & ~n482;
  assign po42 = ~n483 & n484;
  assign n486 = ~pi075 & ~n452;
  assign n487 = ~pi038 & ~n486;
  assign n488 = ~pi032 & pi078;
  assign n489 = po46 & n488;
  assign n490 = ~pi033 & n430;
  assign n491 = n489 & n490;
  assign n492 = ~n487 & ~n491;
  assign n493 = ~pi034 & pi132;
  assign n494 = pi133 & ~n493;
  assign n495 = pi125 & n494;
  assign n496 = ~pi035 & pi133;
  assign n497 = pi132 & ~n496;
  assign n498 = pi125 & n497;
  assign n499 = ~pi032 & ~pi130;
  assign n500 = n460 & ~n499;
  assign n501 = ~n493 & ~n496;
  assign n502 = pi125 & n501;
  assign n503 = pi131 & pi134;
  assign n504 = n500 & n502;
  assign n505 = n503 & n504;
  assign n506 = ~pi033 & pi131;
  assign n507 = pi134 & ~n506;
  assign n508 = n500 & n507;
  assign n509 = ~pi130 & n460;
  assign n510 = n507 & n509;
  assign n511 = n502 & n510;
  assign n512 = ~pi078 & ~n502;
  assign n513 = pi032 & ~n511;
  assign n514 = ~n431 & ~n508;
  assign n515 = ~n513 & ~n514;
  assign n516 = ~n512 & n515;
  assign n517 = ~pi036 & ~n501;
  assign n518 = pi035 & ~n495;
  assign n519 = ~n517 & ~n518;
  assign n520 = pi034 & ~n498;
  assign n521 = pi033 & ~n505;
  assign n522 = ~n520 & ~n521;
  assign n523 = n519 & n522;
  assign n524 = n516 & n523;
  assign n525 = ~pi038 & ~n524;
  assign n526 = ~po89 & ~n525;
  assign n527 = ~pi079 & ~n492;
  assign n528 = pi079 & ~n526;
  assign n529 = ~pi075 & n528;
  assign po43 = n527 | n529;
  assign n531 = ~pi038 & ~pi079;
  assign n532 = ~pi075 & ~n526;
  assign n533 = ~n531 & ~n532;
  assign n534 = pi080 & ~n533;
  assign n535 = ~pi080 & ~n492;
  assign n536 = pi079 & n535;
  assign po44 = n534 | n536;
  assign n538 = pi086 & ~pi087;
  assign n539 = pi088 & n538;
  assign n540 = pi031 & ~pi090;
  assign n541 = pi084 & ~pi090;
  assign n542 = ~pi089 & ~n540;
  assign n543 = pi089 & n541;
  assign n544 = ~n542 & ~n543;
  assign n545 = n539 & ~n544;
  assign n546 = ~pi072 & n545;
  assign n547 = ~pi083 & ~n546;
  assign po47 = ~pi073 & ~n547;
  assign n549 = ~pi029 & ~pi030;
  assign n550 = pi031 & ~n549;
  assign n551 = ~pi090 & n539;
  assign n552 = ~pi089 & ~n550;
  assign n553 = ~pi072 & ~n552;
  assign n554 = n551 & n553;
  assign n555 = pi084 & ~n554;
  assign n556 = ~pi084 & n539;
  assign n557 = n550 & n556;
  assign n558 = ~pi072 & ~pi090;
  assign n559 = ~pi089 & n558;
  assign n560 = n557 & n559;
  assign n561 = ~n555 & ~n560;
  assign po48 = ~pi073 & ~n561;
  assign n563 = pi031 & n549;
  assign n564 = ~pi072 & ~pi089;
  assign n565 = ~pi090 & ~n563;
  assign n566 = n539 & ~n565;
  assign n567 = n564 & n566;
  assign n568 = ~pi085 & n567;
  assign n569 = pi085 & ~n567;
  assign n570 = ~n568 & ~n569;
  assign po49 = ~pi073 & ~n570;
  assign n572 = pi086 & n400;
  assign n573 = ~pi073 & n572;
  assign n574 = ~pi086 & ~po36;
  assign po50 = n573 | n574;
  assign n576 = pi086 & ~n400;
  assign n577 = ~pi073 & ~n576;
  assign n578 = pi087 & n577;
  assign n579 = ~pi087 & ~po36;
  assign n580 = pi086 & n579;
  assign po51 = n578 | n580;
  assign n582 = pi087 & n576;
  assign n583 = pi086 & pi087;
  assign n584 = ~po36 & n583;
  assign n585 = ~pi088 & n584;
  assign n586 = ~pi073 & ~n582;
  assign n587 = pi088 & n586;
  assign po52 = n585 | n587;
  assign n589 = pi088 & n582;
  assign n590 = ~pi089 & n584;
  assign n591 = pi088 & n590;
  assign n592 = ~pi073 & ~n589;
  assign n593 = pi089 & n592;
  assign po53 = n591 | n593;
  assign n595 = pi089 & n589;
  assign n596 = ~pi073 & pi090;
  assign n597 = ~n595 & n596;
  assign n598 = pi088 & pi089;
  assign n599 = ~pi090 & n584;
  assign n600 = n598 & n599;
  assign po54 = n597 | n600;
  assign n602 = ~pi083 & ~n545;
  assign n603 = ~pi072 & ~n602;
  assign n604 = ~pi091 & n603;
  assign n605 = pi091 & ~n603;
  assign n606 = ~n604 & ~n605;
  assign po55 = ~pi073 & ~n606;
  assign n608 = pi091 & n603;
  assign n609 = pi092 & ~n608;
  assign n610 = n259 & n603;
  assign n611 = ~n609 & ~n610;
  assign po56 = ~pi073 & ~n611;
  assign n613 = pi004 & ~pi006;
  assign n614 = ~pi073 & ~n613;
  assign n615 = ~pi073 & n613;
  assign n616 = pi094 & n615;
  assign n617 = pi093 & n614;
  assign po57 = n616 | n617;
  assign n619 = pi095 & n615;
  assign n620 = pi094 & n614;
  assign po58 = n619 | n620;
  assign n622 = pi096 & n615;
  assign n623 = pi095 & n614;
  assign po59 = n622 | n623;
  assign n625 = pi097 & n615;
  assign n626 = pi096 & n614;
  assign po60 = n625 | n626;
  assign n628 = pi098 & n615;
  assign n629 = pi097 & n614;
  assign po61 = n628 | n629;
  assign n631 = pi099 & n615;
  assign n632 = pi098 & n614;
  assign po62 = n631 | n632;
  assign n634 = pi100 & n615;
  assign n635 = pi099 & n614;
  assign po63 = n634 | n635;
  assign n637 = pi100 & n614;
  assign n638 = pi005 & n615;
  assign po64 = n637 | n638;
  assign n640 = pi004 & pi006;
  assign n641 = ~pi073 & ~n640;
  assign n642 = ~pi073 & n640;
  assign n643 = pi102 & n642;
  assign n644 = pi101 & n641;
  assign po65 = n643 | n644;
  assign n646 = pi103 & n642;
  assign n647 = pi102 & n641;
  assign po66 = n646 | n647;
  assign n649 = pi104 & n642;
  assign n650 = pi103 & n641;
  assign po67 = n649 | n650;
  assign n652 = pi105 & n642;
  assign n653 = pi104 & n641;
  assign po68 = n652 | n653;
  assign n655 = pi106 & n642;
  assign n656 = pi105 & n641;
  assign po69 = n655 | n656;
  assign n658 = pi107 & n642;
  assign n659 = pi106 & n641;
  assign po70 = n658 | n659;
  assign n661 = pi108 & n642;
  assign n662 = pi107 & n641;
  assign po71 = n661 | n662;
  assign n664 = pi108 & n641;
  assign n665 = pi005 & n642;
  assign po72 = n664 | n665;
  assign n667 = pi002 & ~pi003;
  assign n668 = ~pi072 & ~n262;
  assign n669 = ~pi001 & ~n668;
  assign n670 = ~pi001 & n668;
  assign n671 = pi110 & n670;
  assign n672 = pi001 & pi093;
  assign n673 = pi109 & n669;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n671 & n674;
  assign n676 = pi040 & n667;
  assign n677 = pi003 & pi056;
  assign n678 = n236 & ~n675;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n676 & n679;
  assign po73 = ~pi073 & ~n680;
  assign n682 = ~pi003 & ~pi073;
  assign n683 = pi003 & ~pi073;
  assign n684 = ~pi002 & n669;
  assign n685 = ~pi002 & n670;
  assign n686 = pi001 & ~pi002;
  assign n687 = pi094 & n686;
  assign n688 = pi111 & n685;
  assign n689 = ~n687 & ~n688;
  assign n690 = pi002 & pi041;
  assign n691 = pi110 & n684;
  assign n692 = ~n690 & ~n691;
  assign n693 = n689 & n692;
  assign n694 = pi057 & n683;
  assign n695 = n682 & ~n693;
  assign po74 = n694 | n695;
  assign n697 = pi095 & n686;
  assign n698 = pi112 & n685;
  assign n699 = ~n697 & ~n698;
  assign n700 = pi002 & pi042;
  assign n701 = pi111 & n684;
  assign n702 = ~n700 & ~n701;
  assign n703 = n699 & n702;
  assign n704 = pi058 & n683;
  assign n705 = n682 & ~n703;
  assign po75 = n704 | n705;
  assign n707 = pi002 & n682;
  assign n708 = pi113 & n670;
  assign n709 = pi001 & pi096;
  assign n710 = pi112 & n669;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n708 & n711;
  assign n713 = ~pi002 & n682;
  assign n714 = ~n712 & n713;
  assign n715 = pi059 & n683;
  assign n716 = pi043 & n707;
  assign n717 = ~n715 & ~n716;
  assign po76 = n714 | ~n717;
  assign n719 = pi114 & n670;
  assign n720 = pi001 & pi097;
  assign n721 = pi113 & n669;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~n719 & n722;
  assign n724 = n713 & ~n723;
  assign n725 = pi060 & n683;
  assign n726 = pi044 & n707;
  assign n727 = ~n725 & ~n726;
  assign po77 = n724 | ~n727;
  assign n729 = pi115 & n670;
  assign n730 = pi001 & pi098;
  assign n731 = pi114 & n669;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n729 & n732;
  assign n734 = n713 & ~n733;
  assign n735 = pi061 & n683;
  assign n736 = pi045 & n707;
  assign n737 = ~n735 & ~n736;
  assign po78 = n734 | ~n737;
  assign n739 = pi116 & n670;
  assign n740 = pi001 & pi099;
  assign n741 = pi115 & n669;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~n739 & n742;
  assign n744 = n713 & ~n743;
  assign n745 = pi062 & n683;
  assign n746 = pi046 & n707;
  assign n747 = ~n745 & ~n746;
  assign po79 = n744 | ~n747;
  assign n749 = pi117 & n670;
  assign n750 = pi001 & pi100;
  assign n751 = pi116 & n669;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~n749 & n752;
  assign n754 = pi047 & n667;
  assign n755 = n236 & ~n753;
  assign n756 = pi003 & pi063;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n754 & n757;
  assign po80 = ~pi073 & ~n758;
  assign n760 = pi118 & n670;
  assign n761 = pi001 & pi101;
  assign n762 = pi117 & n669;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n760 & n763;
  assign n765 = n713 & ~n764;
  assign n766 = pi064 & n683;
  assign n767 = pi048 & n707;
  assign n768 = ~n766 & ~n767;
  assign po81 = n765 | ~n768;
  assign n770 = pi102 & n686;
  assign n771 = pi119 & n685;
  assign n772 = ~n770 & ~n771;
  assign n773 = pi002 & pi049;
  assign n774 = pi118 & n684;
  assign n775 = ~n773 & ~n774;
  assign n776 = n772 & n775;
  assign n777 = pi065 & n683;
  assign n778 = n682 & ~n776;
  assign po82 = n777 | n778;
  assign n780 = pi120 & n670;
  assign n781 = pi001 & pi103;
  assign n782 = pi119 & n669;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n780 & n783;
  assign n785 = pi003 & pi066;
  assign n786 = pi050 & n667;
  assign n787 = n236 & ~n784;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~n785 & n788;
  assign po83 = ~pi073 & ~n789;
  assign n791 = pi121 & n670;
  assign n792 = pi001 & pi104;
  assign n793 = pi120 & n669;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~n791 & n794;
  assign n796 = pi003 & pi067;
  assign n797 = pi051 & n667;
  assign n798 = n236 & ~n795;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n796 & n799;
  assign po84 = ~pi073 & ~n800;
  assign n802 = pi122 & n670;
  assign n803 = pi001 & pi105;
  assign n804 = pi121 & n669;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n802 & n805;
  assign n807 = pi003 & pi068;
  assign n808 = pi052 & n667;
  assign n809 = n236 & ~n806;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~n807 & n810;
  assign po85 = ~pi073 & ~n811;
  assign n813 = pi123 & n670;
  assign n814 = pi001 & pi106;
  assign n815 = pi122 & n669;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~n813 & n816;
  assign n818 = n713 & ~n817;
  assign n819 = pi053 & n707;
  assign n820 = pi069 & n683;
  assign n821 = ~n819 & ~n820;
  assign po86 = n818 | ~n821;
  assign n823 = pi124 & n670;
  assign n824 = pi001 & pi107;
  assign n825 = pi123 & n669;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~n823 & n826;
  assign n828 = pi070 & n683;
  assign n829 = pi054 & n707;
  assign n830 = ~n828 & ~n829;
  assign n831 = n713 & ~n827;
  assign po87 = ~n830 | n831;
  assign n833 = pi108 & n686;
  assign n834 = pi002 & pi055;
  assign n835 = pi124 & n684;
  assign n836 = ~n834 & ~n835;
  assign n837 = ~n833 & n836;
  assign n838 = pi071 & n683;
  assign n839 = n682 & ~n837;
  assign po88 = n838 | n839;
  assign n841 = ~pi126 & n469;
  assign n842 = pi126 & po89;
  assign po90 = n841 | n842;
  assign n844 = ~pi126 & n465;
  assign n845 = ~po89 & ~n844;
  assign n846 = pi127 & ~n845;
  assign n847 = ~pi127 & n469;
  assign n848 = pi126 & n847;
  assign po91 = n846 | n848;
  assign n850 = ~pi127 & n465;
  assign n851 = n845 & ~n850;
  assign n852 = n432 & n469;
  assign n853 = ~pi128 & n852;
  assign n854 = pi128 & ~n851;
  assign po92 = n853 | n854;
  assign n856 = pi127 & pi128;
  assign n857 = n465 & ~n856;
  assign n858 = n845 & ~n857;
  assign n859 = n434 & n465;
  assign n860 = ~pi129 & n859;
  assign n861 = pi129 & ~n858;
  assign po93 = n860 | n861;
  assign n863 = ~n460 & n465;
  assign n864 = ~po89 & ~n863;
  assign n865 = pi130 & ~n864;
  assign n866 = n469 & n509;
  assign po94 = n865 | n866;
  assign n868 = n465 & ~n509;
  assign n869 = ~po89 & ~n868;
  assign n870 = pi131 & ~n869;
  assign n871 = ~pi131 & n866;
  assign po95 = n870 | n871;
  assign n873 = pi125 & pi131;
  assign n874 = n509 & n873;
  assign n875 = ~pi131 & n465;
  assign n876 = n869 & ~n875;
  assign n877 = pi132 & ~n876;
  assign n878 = ~pi132 & n465;
  assign n879 = n874 & n878;
  assign po96 = n877 | n879;
  assign n881 = pi131 & pi132;
  assign n882 = n465 & ~n881;
  assign n883 = n869 & ~n882;
  assign n884 = pi133 & ~n883;
  assign n885 = pi132 & n874;
  assign n886 = ~pi133 & n465;
  assign n887 = n885 & n886;
  assign po97 = n884 | n887;
  assign n889 = pi078 & po46;
  assign n890 = ~pi038 & pi134;
  assign n891 = ~n889 & ~n890;
  assign n892 = pi000 & ~n891;
  assign po98 = ~n483 & n892;
endmodule



// Benchmark "frg2" written by ABC on Sun Apr 22 21:43:04 2018

module frg2 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138;
  wire n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n343, n344, n345,
    n346, n347, n348, n349, n351, n352, n353, n354, n356, n357, n358, n359,
    n361, n362, n363, n364, n366, n367, n368, n369, n371, n372, n373, n374,
    n376, n377, n378, n379, n381, n382, n383, n384, n395, n397, n399, n401,
    n403, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n416,
    n427, n428, n430, n431, n432, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n498, n499, n500, n501, n502, n503, n504,
    n506, n507, n508, n509, n510, n511, n512, n514, n515, n516, n517, n518,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1227, n1228, n1229, n1230, n1231, n1232, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1430, n1431, n1432, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444;
  assign n283 = pi037 & pi114;
  assign n284 = ~pi106 & ~n283;
  assign n285 = pi037 & ~pi114;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~pi037 & pi114;
  assign n288 = ~pi106 & ~n287;
  assign n289 = ~pi037 & ~pi114;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~pi038 & ~pi122;
  assign n292 = pi036 & ~n290;
  assign n293 = n286 & ~n292;
  assign n294 = pi036 & n290;
  assign n295 = pi038 & ~n294;
  assign n296 = ~n293 & n295;
  assign po001 = ~n291 & ~n296;
  assign n298 = pi037 & pi113;
  assign n299 = ~pi105 & ~n298;
  assign n300 = pi037 & ~pi113;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~pi037 & pi113;
  assign n303 = ~pi105 & ~n302;
  assign n304 = ~pi037 & ~pi113;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~pi038 & ~pi121;
  assign n307 = pi036 & ~n305;
  assign n308 = n301 & ~n307;
  assign n309 = pi036 & n305;
  assign n310 = pi038 & ~n309;
  assign n311 = ~n308 & n310;
  assign po002 = ~n306 & ~n311;
  assign n313 = pi037 & pi112;
  assign n314 = ~pi104 & ~n313;
  assign n315 = pi037 & ~pi112;
  assign n316 = ~n314 & ~n315;
  assign n317 = ~pi037 & pi112;
  assign n318 = ~pi104 & ~n317;
  assign n319 = ~pi037 & ~pi112;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~pi038 & ~pi120;
  assign n322 = pi036 & ~n320;
  assign n323 = n316 & ~n322;
  assign n324 = pi036 & n320;
  assign n325 = pi038 & ~n324;
  assign n326 = ~n323 & n325;
  assign po003 = ~n321 & ~n326;
  assign n328 = pi037 & pi111;
  assign n329 = ~pi103 & ~n328;
  assign n330 = pi037 & ~pi111;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~pi037 & pi111;
  assign n333 = ~pi103 & ~n332;
  assign n334 = ~pi037 & ~pi111;
  assign n335 = ~n333 & ~n334;
  assign n336 = ~pi038 & ~pi119;
  assign n337 = pi036 & ~n335;
  assign n338 = n331 & ~n337;
  assign n339 = pi036 & n335;
  assign n340 = pi038 & ~n339;
  assign n341 = ~n338 & n340;
  assign po004 = ~n336 & ~n341;
  assign n343 = pi036 & pi037;
  assign n344 = ~pi036 & ~pi037;
  assign n345 = ~n343 & ~n344;
  assign n346 = ~pi107 & ~n345;
  assign n347 = pi038 & ~n346;
  assign n348 = ~pi115 & ~n344;
  assign n349 = ~n343 & n348;
  assign po007 = n347 & ~n349;
  assign n351 = ~pi108 & ~n345;
  assign n352 = pi038 & ~n351;
  assign n353 = ~pi116 & ~n344;
  assign n354 = ~n343 & n353;
  assign po008 = n352 & ~n354;
  assign n356 = ~pi109 & ~n345;
  assign n357 = pi038 & ~n356;
  assign n358 = ~pi117 & ~n344;
  assign n359 = ~n343 & n358;
  assign po009 = n357 & ~n359;
  assign n361 = ~pi110 & ~n345;
  assign n362 = pi038 & ~n361;
  assign n363 = ~pi118 & ~n344;
  assign n364 = ~n343 & n363;
  assign po010 = n362 & ~n364;
  assign n366 = ~pi111 & ~n345;
  assign n367 = pi038 & ~n366;
  assign n368 = ~pi119 & ~n344;
  assign n369 = ~n343 & n368;
  assign po011 = n367 & ~n369;
  assign n371 = ~pi112 & ~n345;
  assign n372 = pi038 & ~n371;
  assign n373 = ~pi120 & ~n344;
  assign n374 = ~n343 & n373;
  assign po012 = n372 & ~n374;
  assign n376 = ~pi113 & ~n345;
  assign n377 = pi038 & ~n376;
  assign n378 = ~pi121 & ~n344;
  assign n379 = ~n343 & n378;
  assign po013 = n377 & ~n379;
  assign n381 = ~pi114 & ~n345;
  assign n382 = pi038 & ~n381;
  assign n383 = ~pi122 & ~n344;
  assign n384 = ~n343 & n383;
  assign po014 = n382 & ~n384;
  assign po015 = pi038 & pi115;
  assign po016 = pi038 & pi116;
  assign po017 = pi038 & pi117;
  assign po018 = pi038 & pi118;
  assign po019 = pi038 & pi119;
  assign po020 = pi038 & pi120;
  assign po021 = pi038 & pi121;
  assign po022 = pi038 & pi122;
  assign po023 = pi057 & ~pi138;
  assign n395 = pi058 & ~pi139;
  assign po025 = pi039 | ~n395;
  assign n397 = pi059 & ~pi139;
  assign po026 = pi039 | ~n397;
  assign n399 = pi060 & ~pi139;
  assign po027 = pi039 | ~n399;
  assign n401 = pi061 & ~pi139;
  assign po028 = pi039 | ~n401;
  assign n403 = pi062 & ~pi139;
  assign po029 = pi039 | ~n403;
  assign n405 = pi127 & pi128;
  assign n406 = ~pi130 & ~pi131;
  assign n407 = ~pi129 & n406;
  assign n408 = ~pi056 & pi137;
  assign n409 = pi056 & ~pi137;
  assign n410 = ~n408 & ~n409;
  assign n411 = n405 & n407;
  assign n412 = ~pi064 & ~n411;
  assign n413 = n407 & ~n410;
  assign n414 = n405 & n413;
  assign po030 = ~n412 & ~n414;
  assign n416 = pi063 & ~pi139;
  assign po035 = ~pi058 | ~n416;
  assign po036 = ~pi059 | ~n416;
  assign po037 = ~pi060 | ~n416;
  assign po038 = ~pi061 | ~n416;
  assign po039 = ~pi062 | ~n416;
  assign po040 = ~pi058 | ~pi140;
  assign po041 = ~pi059 | ~pi140;
  assign po042 = ~pi060 | ~pi140;
  assign po043 = ~pi061 | ~pi140;
  assign po044 = ~pi062 | ~pi140;
  assign n427 = pi056 & pi137;
  assign n428 = ~pi056 & ~pi137;
  assign po051 = n427 | n428;
  assign n430 = pi128 & ~pi129;
  assign n431 = pi126 & pi127;
  assign n432 = n430 & n431;
  assign po052 = n406 & n432;
  assign n434 = ~pi135 & ~pi136;
  assign n435 = pi133 & pi134;
  assign n436 = n434 & n435;
  assign n437 = ~pi057 & pi132;
  assign n438 = n435 & n437;
  assign n439 = n434 & n438;
  assign n440 = ~pi052 & pi062;
  assign n441 = ~n436 & ~n440;
  assign n442 = pi142 & n441;
  assign n443 = ~n439 & ~n442;
  assign n444 = ~pi050 & pi060;
  assign n445 = ~pi051 & pi061;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n436 & ~n446;
  assign n448 = ~n443 & ~n447;
  assign n449 = ~pi048 & pi058;
  assign n450 = ~pi049 & pi059;
  assign n451 = ~n449 & ~n450;
  assign n452 = ~n436 & ~n451;
  assign n453 = n448 & ~n452;
  assign n454 = ~pi042 & n453;
  assign po053 = pi040 & n454;
  assign n456 = ~pi042 & ~pi053;
  assign n457 = pi040 & n456;
  assign n458 = ~pi059 & ~pi060;
  assign n459 = ~pi058 & n458;
  assign n460 = ~pi061 & ~pi062;
  assign n461 = n459 & n460;
  assign n462 = ~pi055 & n461;
  assign n463 = ~pi054 & n462;
  assign n464 = ~pi057 & pi058;
  assign n465 = ~pi042 & n464;
  assign n466 = ~pi053 & ~pi054;
  assign n467 = pi055 & ~n466;
  assign n468 = ~pi039 & n461;
  assign n469 = ~n467 & n468;
  assign n470 = n465 & ~n469;
  assign n471 = pi040 & n470;
  assign n472 = n457 & n463;
  assign n473 = ~pi039 & n472;
  assign po054 = n471 | n473;
  assign n475 = pi054 & pi055;
  assign n476 = ~pi053 & ~n475;
  assign n477 = pi054 & ~pi055;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~pi039 & n462;
  assign n480 = ~pi059 & ~n479;
  assign n481 = pi040 & ~pi042;
  assign n482 = ~n480 & n481;
  assign n483 = pi057 & ~n479;
  assign n484 = ~pi039 & ~n478;
  assign n485 = n461 & n484;
  assign n486 = ~n483 & ~n485;
  assign po055 = n482 & n486;
  assign n488 = pi053 & pi055;
  assign n489 = ~pi054 & ~n488;
  assign n490 = pi053 & ~pi055;
  assign n491 = ~n489 & ~n490;
  assign n492 = ~pi060 & ~n479;
  assign n493 = n481 & ~n492;
  assign n494 = ~pi039 & ~n491;
  assign n495 = n461 & n494;
  assign n496 = ~n483 & ~n495;
  assign po056 = n493 & n496;
  assign n498 = ~pi054 & ~pi055;
  assign n499 = ~n476 & ~n498;
  assign n500 = ~pi061 & ~n479;
  assign n501 = n481 & ~n500;
  assign n502 = ~pi039 & ~n499;
  assign n503 = n461 & n502;
  assign n504 = ~n483 & ~n503;
  assign po057 = n501 & n504;
  assign n506 = ~pi054 & n461;
  assign n507 = ~pi039 & ~pi053;
  assign n508 = n506 & n507;
  assign n509 = ~pi042 & ~n479;
  assign n510 = pi040 & n509;
  assign n511 = ~pi057 & pi062;
  assign n512 = ~n508 & ~n511;
  assign po058 = n510 & ~n512;
  assign n514 = pi063 & n453;
  assign n515 = ~pi042 & ~n514;
  assign n516 = pi040 & n515;
  assign n517 = ~pi039 & pi041;
  assign n518 = ~pi063 & ~n517;
  assign po059 = n516 & ~n518;
  assign n520 = ~pi126 & pi127;
  assign n521 = n430 & n520;
  assign n522 = n406 & n521;
  assign n523 = ~pi065 & pi140;
  assign n524 = pi140 & ~n522;
  assign n525 = ~pi035 & n468;
  assign n526 = ~pi042 & ~n525;
  assign n527 = pi040 & n526;
  assign n528 = ~n461 & ~n524;
  assign n529 = ~pi064 & n528;
  assign n530 = n527 & ~n529;
  assign n531 = pi039 & ~n524;
  assign n532 = ~pi064 & n531;
  assign n533 = ~n468 & n523;
  assign n534 = ~n522 & n533;
  assign n535 = ~n532 & ~n534;
  assign po060 = n530 & n535;
  assign n537 = ~pi066 & pi140;
  assign n538 = ~pi034 & n468;
  assign n539 = ~pi042 & ~n538;
  assign n540 = pi040 & n539;
  assign n541 = ~pi065 & n528;
  assign n542 = n540 & ~n541;
  assign n543 = ~pi065 & n531;
  assign n544 = ~n468 & n537;
  assign n545 = ~n522 & n544;
  assign n546 = ~n543 & ~n545;
  assign po061 = n542 & n546;
  assign n548 = ~pi067 & pi140;
  assign n549 = ~pi033 & n468;
  assign n550 = ~pi042 & ~n549;
  assign n551 = pi040 & n550;
  assign n552 = ~pi066 & n528;
  assign n553 = n551 & ~n552;
  assign n554 = ~pi066 & n531;
  assign n555 = ~n468 & n548;
  assign n556 = ~n522 & n555;
  assign n557 = ~n554 & ~n556;
  assign po062 = n553 & n557;
  assign n559 = ~pi068 & pi140;
  assign n560 = ~pi032 & n468;
  assign n561 = ~pi042 & ~n560;
  assign n562 = pi040 & n561;
  assign n563 = ~pi067 & n528;
  assign n564 = n562 & ~n563;
  assign n565 = ~pi067 & n531;
  assign n566 = ~n468 & n559;
  assign n567 = ~n522 & n566;
  assign n568 = ~n565 & ~n567;
  assign po063 = n564 & n568;
  assign n570 = ~pi069 & pi140;
  assign n571 = ~pi031 & n468;
  assign n572 = ~pi042 & ~n571;
  assign n573 = pi040 & n572;
  assign n574 = ~pi068 & n528;
  assign n575 = n573 & ~n574;
  assign n576 = ~pi068 & n531;
  assign n577 = ~n468 & n570;
  assign n578 = ~n522 & n577;
  assign n579 = ~n576 & ~n578;
  assign po064 = n575 & n579;
  assign n581 = ~pi070 & pi140;
  assign n582 = ~pi030 & n468;
  assign n583 = ~pi042 & ~n582;
  assign n584 = pi040 & n583;
  assign n585 = ~pi069 & n528;
  assign n586 = n584 & ~n585;
  assign n587 = ~pi069 & n531;
  assign n588 = ~n468 & n581;
  assign n589 = ~n522 & n588;
  assign n590 = ~n587 & ~n589;
  assign po065 = n586 & n590;
  assign n592 = ~pi071 & pi140;
  assign n593 = ~pi029 & n468;
  assign n594 = ~pi042 & ~n593;
  assign n595 = pi040 & n594;
  assign n596 = ~pi070 & n528;
  assign n597 = n595 & ~n596;
  assign n598 = ~pi070 & n531;
  assign n599 = ~n468 & n592;
  assign n600 = ~n522 & n599;
  assign n601 = ~n598 & ~n600;
  assign po066 = n597 & n601;
  assign n603 = ~pi072 & pi140;
  assign n604 = ~pi038 & n468;
  assign n605 = ~pi042 & ~n604;
  assign n606 = pi040 & n605;
  assign n607 = ~pi071 & n528;
  assign n608 = n606 & ~n607;
  assign n609 = ~pi071 & n531;
  assign n610 = ~n468 & n603;
  assign n611 = ~n522 & n610;
  assign n612 = ~n609 & ~n611;
  assign po067 = n608 & n612;
  assign n614 = ~pi073 & pi140;
  assign n615 = ~pi036 & n468;
  assign n616 = ~pi042 & ~n615;
  assign n617 = pi040 & n616;
  assign n618 = ~pi072 & n528;
  assign n619 = n617 & ~n618;
  assign n620 = ~pi072 & n531;
  assign n621 = ~n468 & n614;
  assign n622 = ~n522 & n621;
  assign n623 = ~n620 & ~n622;
  assign po068 = n619 & n623;
  assign n625 = ~pi074 & pi140;
  assign n626 = ~pi037 & n468;
  assign n627 = ~pi042 & ~n626;
  assign n628 = pi040 & n627;
  assign n629 = ~pi073 & n528;
  assign n630 = n628 & ~n629;
  assign n631 = ~pi073 & n531;
  assign n632 = ~n468 & n625;
  assign n633 = ~n522 & n632;
  assign n634 = ~n631 & ~n633;
  assign po069 = n630 & n634;
  assign n636 = ~pi075 & pi140;
  assign n637 = ~pi016 & n468;
  assign n638 = ~pi042 & ~n637;
  assign n639 = pi040 & n638;
  assign n640 = ~pi074 & n528;
  assign n641 = n639 & ~n640;
  assign n642 = ~pi074 & n531;
  assign n643 = ~n468 & n636;
  assign n644 = ~n522 & n643;
  assign n645 = ~n642 & ~n644;
  assign po070 = n641 & n645;
  assign n647 = ~pi076 & pi140;
  assign n648 = ~pi017 & n468;
  assign n649 = ~pi042 & ~n648;
  assign n650 = pi040 & n649;
  assign n651 = ~pi075 & n528;
  assign n652 = n650 & ~n651;
  assign n653 = ~pi075 & n531;
  assign n654 = ~n468 & n647;
  assign n655 = ~n522 & n654;
  assign n656 = ~n653 & ~n655;
  assign po071 = n652 & n656;
  assign n658 = ~pi077 & pi140;
  assign n659 = ~pi018 & n468;
  assign n660 = ~pi042 & ~n659;
  assign n661 = pi040 & n660;
  assign n662 = ~pi076 & n528;
  assign n663 = n661 & ~n662;
  assign n664 = ~pi076 & n531;
  assign n665 = ~n468 & n658;
  assign n666 = ~n522 & n665;
  assign n667 = ~n664 & ~n666;
  assign po072 = n663 & n667;
  assign n669 = ~pi078 & pi140;
  assign n670 = ~pi019 & n468;
  assign n671 = ~pi042 & ~n670;
  assign n672 = pi040 & n671;
  assign n673 = ~pi077 & n528;
  assign n674 = n672 & ~n673;
  assign n675 = ~pi077 & n531;
  assign n676 = ~n468 & n669;
  assign n677 = ~n522 & n676;
  assign n678 = ~n675 & ~n677;
  assign po073 = n674 & n678;
  assign n680 = ~pi079 & pi140;
  assign n681 = ~pi020 & n468;
  assign n682 = ~pi042 & ~n681;
  assign n683 = pi040 & n682;
  assign n684 = ~pi078 & n528;
  assign n685 = n683 & ~n684;
  assign n686 = ~pi078 & n531;
  assign n687 = ~n468 & n680;
  assign n688 = ~n522 & n687;
  assign n689 = ~n686 & ~n688;
  assign po074 = n685 & n689;
  assign n691 = ~pi080 & pi140;
  assign n692 = ~pi021 & n468;
  assign n693 = ~pi042 & ~n692;
  assign n694 = pi040 & n693;
  assign n695 = ~pi079 & n528;
  assign n696 = n694 & ~n695;
  assign n697 = ~pi079 & n531;
  assign n698 = ~n468 & n691;
  assign n699 = ~n522 & n698;
  assign n700 = ~n697 & ~n699;
  assign po075 = n696 & n700;
  assign n702 = ~pi081 & pi140;
  assign n703 = ~pi022 & n468;
  assign n704 = ~pi042 & ~n703;
  assign n705 = pi040 & n704;
  assign n706 = ~pi080 & n528;
  assign n707 = n705 & ~n706;
  assign n708 = ~pi080 & n531;
  assign n709 = ~n468 & n702;
  assign n710 = ~n522 & n709;
  assign n711 = ~n708 & ~n710;
  assign po076 = n707 & n711;
  assign n713 = ~pi082 & pi140;
  assign n714 = ~pi023 & n468;
  assign n715 = ~pi042 & ~n714;
  assign n716 = pi040 & n715;
  assign n717 = ~pi081 & n528;
  assign n718 = n716 & ~n717;
  assign n719 = ~pi081 & n531;
  assign n720 = ~n468 & n713;
  assign n721 = ~n522 & n720;
  assign n722 = ~n719 & ~n721;
  assign po077 = n718 & n722;
  assign n724 = ~pi083 & pi140;
  assign n725 = ~pi024 & n468;
  assign n726 = ~pi042 & ~n725;
  assign n727 = pi040 & n726;
  assign n728 = ~pi082 & n528;
  assign n729 = n727 & ~n728;
  assign n730 = ~pi082 & n531;
  assign n731 = ~n468 & n724;
  assign n732 = ~n522 & n731;
  assign n733 = ~n730 & ~n732;
  assign po078 = n729 & n733;
  assign n735 = ~pi084 & pi140;
  assign n736 = ~pi025 & n468;
  assign n737 = ~pi042 & ~n736;
  assign n738 = pi040 & n737;
  assign n739 = ~pi083 & n528;
  assign n740 = n738 & ~n739;
  assign n741 = ~pi083 & n531;
  assign n742 = ~n468 & n735;
  assign n743 = ~n522 & n742;
  assign n744 = ~n741 & ~n743;
  assign po079 = n740 & n744;
  assign n746 = ~pi085 & pi140;
  assign n747 = ~pi026 & n468;
  assign n748 = ~pi042 & ~n747;
  assign n749 = pi040 & n748;
  assign n750 = ~pi084 & n528;
  assign n751 = n749 & ~n750;
  assign n752 = ~pi084 & n531;
  assign n753 = ~n468 & n746;
  assign n754 = ~n522 & n753;
  assign n755 = ~n752 & ~n754;
  assign po080 = n751 & n755;
  assign n757 = ~pi086 & pi140;
  assign n758 = ~pi027 & n468;
  assign n759 = ~pi042 & ~n758;
  assign n760 = pi040 & n759;
  assign n761 = ~pi085 & n528;
  assign n762 = n760 & ~n761;
  assign n763 = ~pi085 & n531;
  assign n764 = ~n468 & n757;
  assign n765 = ~n522 & n764;
  assign n766 = ~n763 & ~n765;
  assign po081 = n762 & n766;
  assign n768 = ~pi087 & pi140;
  assign n769 = ~pi028 & n468;
  assign n770 = ~pi042 & ~n769;
  assign n771 = pi040 & n770;
  assign n772 = ~pi086 & n528;
  assign n773 = n771 & ~n772;
  assign n774 = ~pi086 & n531;
  assign n775 = ~n468 & n768;
  assign n776 = ~n522 & n775;
  assign n777 = ~n774 & ~n776;
  assign po082 = n773 & n777;
  assign n779 = pi008 & ~pi037;
  assign n780 = pi036 & n779;
  assign n781 = pi036 & ~pi037;
  assign n782 = pi000 & ~n781;
  assign n783 = ~n780 & ~n782;
  assign n784 = ~pi088 & pi140;
  assign n785 = ~n524 & ~n604;
  assign n786 = ~pi087 & n785;
  assign n787 = n468 & n783;
  assign n788 = ~pi038 & n787;
  assign n789 = ~n604 & n784;
  assign n790 = ~n522 & n789;
  assign n791 = ~n788 & ~n790;
  assign n792 = ~n786 & n791;
  assign po083 = n481 & n792;
  assign n794 = pi009 & ~pi037;
  assign n795 = pi036 & n794;
  assign n796 = pi001 & ~n781;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~pi089 & pi140;
  assign n799 = ~pi088 & n785;
  assign n800 = n468 & n797;
  assign n801 = ~pi038 & n800;
  assign n802 = ~n604 & n798;
  assign n803 = ~n522 & n802;
  assign n804 = ~n801 & ~n803;
  assign n805 = ~n799 & n804;
  assign po084 = n481 & n805;
  assign n807 = pi010 & ~pi037;
  assign n808 = pi036 & n807;
  assign n809 = pi002 & ~n781;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~pi090 & pi140;
  assign n812 = ~pi089 & n785;
  assign n813 = n468 & n810;
  assign n814 = ~pi038 & n813;
  assign n815 = ~n604 & n811;
  assign n816 = ~n522 & n815;
  assign n817 = ~n814 & ~n816;
  assign n818 = ~n812 & n817;
  assign po085 = n481 & n818;
  assign n820 = pi011 & ~pi037;
  assign n821 = pi036 & n820;
  assign n822 = pi003 & ~n781;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~pi091 & pi140;
  assign n825 = ~pi090 & n785;
  assign n826 = n468 & n823;
  assign n827 = ~pi038 & n826;
  assign n828 = ~n604 & n824;
  assign n829 = ~n522 & n828;
  assign n830 = ~n827 & ~n829;
  assign n831 = ~n825 & n830;
  assign po086 = n481 & n831;
  assign n833 = pi012 & ~pi037;
  assign n834 = pi036 & n833;
  assign n835 = pi004 & ~n781;
  assign n836 = ~n834 & ~n835;
  assign n837 = ~pi092 & pi140;
  assign n838 = ~pi091 & n785;
  assign n839 = n468 & n836;
  assign n840 = ~pi038 & n839;
  assign n841 = ~n604 & n837;
  assign n842 = ~n522 & n841;
  assign n843 = ~n840 & ~n842;
  assign n844 = ~n838 & n843;
  assign po087 = n481 & n844;
  assign n846 = pi013 & ~pi037;
  assign n847 = pi036 & n846;
  assign n848 = pi005 & ~n781;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~pi093 & pi140;
  assign n851 = ~pi092 & n785;
  assign n852 = n468 & n849;
  assign n853 = ~pi038 & n852;
  assign n854 = ~n604 & n850;
  assign n855 = ~n522 & n854;
  assign n856 = ~n853 & ~n855;
  assign n857 = ~n851 & n856;
  assign po088 = n481 & n857;
  assign n859 = pi014 & ~pi037;
  assign n860 = pi036 & n859;
  assign n861 = pi006 & ~n781;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~pi094 & pi140;
  assign n864 = ~pi093 & n785;
  assign n865 = n468 & n862;
  assign n866 = ~pi038 & n865;
  assign n867 = ~n604 & n863;
  assign n868 = ~n522 & n867;
  assign n869 = ~n866 & ~n868;
  assign n870 = ~n864 & n869;
  assign po089 = n481 & n870;
  assign n872 = pi015 & ~pi037;
  assign n873 = pi036 & n872;
  assign n874 = pi007 & ~n781;
  assign n875 = ~n873 & ~n874;
  assign n876 = ~pi095 & pi140;
  assign n877 = ~pi094 & n785;
  assign n878 = n468 & n875;
  assign n879 = ~pi038 & n878;
  assign n880 = ~n604 & n876;
  assign n881 = ~n522 & n880;
  assign n882 = ~n879 & ~n881;
  assign n883 = ~n877 & n882;
  assign po090 = n481 & n883;
  assign n885 = pi096 & pi140;
  assign n886 = ~n345 & n461;
  assign n887 = ~pi038 & ~pi039;
  assign n888 = n886 & n887;
  assign n889 = ~pi036 & pi037;
  assign n890 = ~n781 & ~n889;
  assign n891 = n461 & n890;
  assign n892 = n887 & n891;
  assign n893 = pi095 & ~n892;
  assign n894 = ~pi140 & n893;
  assign n895 = n604 & n890;
  assign n896 = pi008 & n895;
  assign n897 = ~n894 & ~n896;
  assign n898 = ~n522 & n885;
  assign n899 = ~pi095 & ~n898;
  assign n900 = ~n522 & ~n885;
  assign n901 = ~n888 & ~n900;
  assign n902 = ~n899 & n901;
  assign n903 = n897 & ~n902;
  assign po091 = n481 & ~n903;
  assign n905 = pi097 & pi140;
  assign n906 = pi096 & ~n892;
  assign n907 = ~pi140 & n906;
  assign n908 = pi009 & n895;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n522 & n905;
  assign n911 = ~pi096 & ~n910;
  assign n912 = ~n522 & ~n905;
  assign n913 = ~n888 & ~n912;
  assign n914 = ~n911 & n913;
  assign n915 = n909 & ~n914;
  assign po092 = n481 & ~n915;
  assign n917 = pi098 & pi140;
  assign n918 = pi097 & ~n892;
  assign n919 = ~pi140 & n918;
  assign n920 = pi010 & n895;
  assign n921 = ~n919 & ~n920;
  assign n922 = ~n522 & n917;
  assign n923 = ~pi097 & ~n922;
  assign n924 = ~n522 & ~n917;
  assign n925 = ~n888 & ~n924;
  assign n926 = ~n923 & n925;
  assign n927 = n921 & ~n926;
  assign po093 = n481 & ~n927;
  assign n929 = pi099 & pi140;
  assign n930 = pi098 & ~n892;
  assign n931 = ~pi140 & n930;
  assign n932 = pi011 & n895;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~n522 & n929;
  assign n935 = ~pi098 & ~n934;
  assign n936 = ~n522 & ~n929;
  assign n937 = ~n888 & ~n936;
  assign n938 = ~n935 & n937;
  assign n939 = n933 & ~n938;
  assign po094 = n481 & ~n939;
  assign n941 = pi100 & pi140;
  assign n942 = pi099 & ~n892;
  assign n943 = ~pi140 & n942;
  assign n944 = pi012 & n895;
  assign n945 = ~n943 & ~n944;
  assign n946 = ~n522 & n941;
  assign n947 = ~pi099 & ~n946;
  assign n948 = ~n522 & ~n941;
  assign n949 = ~n888 & ~n948;
  assign n950 = ~n947 & n949;
  assign n951 = n945 & ~n950;
  assign po095 = n481 & ~n951;
  assign n953 = pi101 & pi140;
  assign n954 = pi100 & ~n892;
  assign n955 = ~pi140 & n954;
  assign n956 = pi013 & n895;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n522 & n953;
  assign n959 = ~pi100 & ~n958;
  assign n960 = ~n522 & ~n953;
  assign n961 = ~n888 & ~n960;
  assign n962 = ~n959 & n961;
  assign n963 = n957 & ~n962;
  assign po096 = n481 & ~n963;
  assign n965 = pi102 & pi140;
  assign n966 = pi101 & ~n892;
  assign n967 = ~pi140 & n966;
  assign n968 = pi014 & n895;
  assign n969 = ~n967 & ~n968;
  assign n970 = ~n522 & n965;
  assign n971 = ~pi101 & ~n970;
  assign n972 = ~n522 & ~n965;
  assign n973 = ~n888 & ~n972;
  assign n974 = ~n971 & n973;
  assign n975 = n969 & ~n974;
  assign po097 = n481 & ~n975;
  assign n977 = pi015 & n887;
  assign n978 = ~pi042 & n461;
  assign n979 = pi040 & n978;
  assign n980 = ~pi042 & pi102;
  assign n981 = n468 & n890;
  assign n982 = ~pi038 & n981;
  assign n983 = ~n524 & ~n982;
  assign n984 = n980 & n983;
  assign n985 = pi040 & n984;
  assign n986 = n890 & n979;
  assign n987 = n977 & n986;
  assign po098 = n985 | n987;
  assign n989 = ~n440 & n446;
  assign n990 = n451 & n989;
  assign n991 = ~pi042 & ~n990;
  assign n992 = pi040 & n991;
  assign n993 = pi134 & ~pi135;
  assign n994 = pi133 & n993;
  assign n995 = ~pi136 & n994;
  assign n996 = pi104 & pi139;
  assign n997 = ~n995 & n996;
  assign n998 = n458 & n460;
  assign n999 = ~pi060 & n460;
  assign n1000 = pi061 & pi062;
  assign n1001 = pi060 & ~n460;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~pi058 & n999;
  assign n1004 = ~pi059 & n1003;
  assign n1005 = n1002 & ~n1004;
  assign n1006 = pi058 & ~n998;
  assign n1007 = pi059 & ~n999;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = n1005 & n1008;
  assign n1010 = ~pi042 & pi103;
  assign n1011 = pi060 & pi061;
  assign n1012 = ~n990 & ~n1011;
  assign n1013 = ~n461 & n1012;
  assign n1014 = pi060 & pi062;
  assign n1015 = n1013 & ~n1014;
  assign n1016 = ~n995 & n1015;
  assign n1017 = pi139 & ~n1000;
  assign n1018 = n1016 & n1017;
  assign n1019 = n1008 & n1018;
  assign n1020 = n1010 & ~n1019;
  assign n1021 = pi040 & n1020;
  assign n1022 = n997 & n1009;
  assign n1023 = n992 & n1022;
  assign po099 = n1021 | n1023;
  assign n1025 = pi105 & pi139;
  assign n1026 = ~n995 & n1025;
  assign n1027 = ~pi042 & pi104;
  assign n1028 = ~n1019 & n1027;
  assign n1029 = pi040 & n1028;
  assign n1030 = n1009 & n1026;
  assign n1031 = n992 & n1030;
  assign po100 = n1029 | n1031;
  assign n1033 = pi106 & pi139;
  assign n1034 = ~n995 & n1033;
  assign n1035 = ~pi042 & pi105;
  assign n1036 = ~n1019 & n1035;
  assign n1037 = pi040 & n1036;
  assign n1038 = n1009 & n1034;
  assign n1039 = n992 & n1038;
  assign po101 = n1037 | n1039;
  assign n1041 = pi107 & pi139;
  assign n1042 = ~n995 & n1041;
  assign n1043 = ~pi042 & pi106;
  assign n1044 = ~n1019 & n1043;
  assign n1045 = pi040 & n1044;
  assign n1046 = n1009 & n1042;
  assign n1047 = n992 & n1046;
  assign po102 = n1045 | n1047;
  assign n1049 = pi108 & pi139;
  assign n1050 = ~n995 & n1049;
  assign n1051 = ~pi042 & pi107;
  assign n1052 = ~n1019 & n1051;
  assign n1053 = pi040 & n1052;
  assign n1054 = n1009 & n1050;
  assign n1055 = n992 & n1054;
  assign po103 = n1053 | n1055;
  assign n1057 = pi109 & pi139;
  assign n1058 = ~n995 & n1057;
  assign n1059 = ~pi042 & pi108;
  assign n1060 = ~n1019 & n1059;
  assign n1061 = pi040 & n1060;
  assign n1062 = n1009 & n1058;
  assign n1063 = n992 & n1062;
  assign po104 = n1061 | n1063;
  assign n1065 = pi110 & pi139;
  assign n1066 = ~n995 & n1065;
  assign n1067 = ~pi042 & pi109;
  assign n1068 = ~n1019 & n1067;
  assign n1069 = pi040 & n1068;
  assign n1070 = n1009 & n1066;
  assign n1071 = n992 & n1070;
  assign po105 = n1069 | n1071;
  assign n1073 = pi111 & pi139;
  assign n1074 = ~n995 & n1073;
  assign n1075 = ~pi042 & pi110;
  assign n1076 = ~n1019 & n1075;
  assign n1077 = pi040 & n1076;
  assign n1078 = n1009 & n1074;
  assign n1079 = n992 & n1078;
  assign po106 = n1077 | n1079;
  assign n1081 = pi112 & pi139;
  assign n1082 = ~n995 & n1081;
  assign n1083 = ~pi042 & pi111;
  assign n1084 = ~n1019 & n1083;
  assign n1085 = pi040 & n1084;
  assign n1086 = n1009 & n1082;
  assign n1087 = n992 & n1086;
  assign po107 = n1085 | n1087;
  assign n1089 = pi113 & pi139;
  assign n1090 = ~n995 & n1089;
  assign n1091 = ~pi042 & pi112;
  assign n1092 = ~n1019 & n1091;
  assign n1093 = pi040 & n1092;
  assign n1094 = n1009 & n1090;
  assign n1095 = n992 & n1094;
  assign po108 = n1093 | n1095;
  assign n1097 = pi114 & pi139;
  assign n1098 = ~n995 & n1097;
  assign n1099 = ~pi042 & pi113;
  assign n1100 = ~n1019 & n1099;
  assign n1101 = pi040 & n1100;
  assign n1102 = n1009 & n1098;
  assign n1103 = n992 & n1102;
  assign po109 = n1101 | n1103;
  assign n1105 = pi115 & pi139;
  assign n1106 = ~n995 & n1105;
  assign n1107 = ~pi042 & pi114;
  assign n1108 = ~n1019 & n1107;
  assign n1109 = pi040 & n1108;
  assign n1110 = n1009 & n1106;
  assign n1111 = n992 & n1110;
  assign po110 = n1109 | n1111;
  assign n1113 = pi116 & pi139;
  assign n1114 = ~n995 & n1113;
  assign n1115 = ~pi042 & pi115;
  assign n1116 = ~n1019 & n1115;
  assign n1117 = pi040 & n1116;
  assign n1118 = n1009 & n1114;
  assign n1119 = n992 & n1118;
  assign po111 = n1117 | n1119;
  assign n1121 = pi117 & pi139;
  assign n1122 = ~n995 & n1121;
  assign n1123 = ~pi042 & pi116;
  assign n1124 = ~n1019 & n1123;
  assign n1125 = pi040 & n1124;
  assign n1126 = n1009 & n1122;
  assign n1127 = n992 & n1126;
  assign po112 = n1125 | n1127;
  assign n1129 = pi118 & pi139;
  assign n1130 = ~n995 & n1129;
  assign n1131 = ~pi042 & pi117;
  assign n1132 = ~n1019 & n1131;
  assign n1133 = pi040 & n1132;
  assign n1134 = n1009 & n1130;
  assign n1135 = n992 & n1134;
  assign po113 = n1133 | n1135;
  assign n1137 = pi119 & pi139;
  assign n1138 = ~n995 & n1137;
  assign n1139 = ~pi042 & pi118;
  assign n1140 = ~n1019 & n1139;
  assign n1141 = pi040 & n1140;
  assign n1142 = n1009 & n1138;
  assign n1143 = n992 & n1142;
  assign po114 = n1141 | n1143;
  assign n1145 = pi120 & pi139;
  assign n1146 = ~n995 & n1145;
  assign n1147 = ~pi042 & pi119;
  assign n1148 = ~n1019 & n1147;
  assign n1149 = pi040 & n1148;
  assign n1150 = n1009 & n1146;
  assign n1151 = n992 & n1150;
  assign po115 = n1149 | n1151;
  assign n1153 = pi121 & pi139;
  assign n1154 = ~n995 & n1153;
  assign n1155 = ~pi042 & pi120;
  assign n1156 = ~n1019 & n1155;
  assign n1157 = pi040 & n1156;
  assign n1158 = n1009 & n1154;
  assign n1159 = n992 & n1158;
  assign po116 = n1157 | n1159;
  assign n1161 = pi122 & pi139;
  assign n1162 = ~n995 & n1161;
  assign n1163 = ~pi042 & pi121;
  assign n1164 = ~n1019 & n1163;
  assign n1165 = pi040 & n1164;
  assign n1166 = n1009 & n1162;
  assign n1167 = n992 & n1166;
  assign po117 = n1165 | n1167;
  assign n1169 = pi123 & pi139;
  assign n1170 = ~n995 & n1169;
  assign n1171 = ~pi042 & pi122;
  assign n1172 = ~n1019 & n1171;
  assign n1173 = pi040 & n1172;
  assign n1174 = n1009 & n1170;
  assign n1175 = n992 & n1174;
  assign po118 = n1173 | n1175;
  assign n1177 = pi124 & pi139;
  assign n1178 = ~n995 & n1177;
  assign n1179 = ~pi042 & pi123;
  assign n1180 = ~n1019 & n1179;
  assign n1181 = pi040 & n1180;
  assign n1182 = n1009 & n1178;
  assign n1183 = n992 & n1182;
  assign po119 = n1181 | n1183;
  assign n1185 = pi125 & pi139;
  assign n1186 = ~n995 & n1185;
  assign n1187 = ~pi042 & pi124;
  assign n1188 = ~n1019 & n1187;
  assign n1189 = pi040 & n1188;
  assign n1190 = n1009 & n1186;
  assign n1191 = n992 & n1190;
  assign po120 = n1189 | n1191;
  assign n1193 = pi139 & ~n995;
  assign n1194 = ~n990 & n1193;
  assign n1195 = pi058 & ~pi059;
  assign n1196 = ~pi061 & pi062;
  assign n1197 = ~pi060 & pi061;
  assign n1198 = pi046 & n1197;
  assign n1199 = ~pi062 & n1198;
  assign n1200 = pi045 & n460;
  assign n1201 = ~pi060 & n1196;
  assign n1202 = pi047 & n1201;
  assign n1203 = ~n1200 & ~n1202;
  assign n1204 = pi047 & n1196;
  assign n1205 = ~pi060 & ~n1204;
  assign n1206 = ~n1203 & ~n1205;
  assign n1207 = ~n1199 & ~n1206;
  assign n1208 = pi044 & n999;
  assign n1209 = pi059 & n1208;
  assign n1210 = ~pi059 & ~n1207;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~pi058 & ~n1211;
  assign n1213 = n999 & n1195;
  assign n1214 = pi043 & n1213;
  assign n1215 = ~n1212 & ~n1214;
  assign n1216 = ~pi042 & pi125;
  assign n1217 = ~n1001 & ~n1004;
  assign n1218 = ~n1000 & n1217;
  assign n1219 = ~n990 & n1218;
  assign n1220 = n1193 & n1219;
  assign n1221 = n1008 & n1220;
  assign n1222 = n1216 & ~n1221;
  assign n1223 = pi040 & n1222;
  assign n1224 = n1194 & ~n1215;
  assign n1225 = n481 & n1224;
  assign po121 = n1223 | n1225;
  assign n1227 = ~pi042 & ~n468;
  assign n1228 = pi040 & n1227;
  assign n1229 = pi126 & ~n522;
  assign n1230 = pi140 & n1229;
  assign n1231 = n1228 & ~n1230;
  assign n1232 = ~pi126 & ~n524;
  assign po122 = n1231 & ~n1232;
  assign n1234 = ~pi126 & pi140;
  assign n1235 = ~n522 & n1234;
  assign n1236 = ~pi126 & ~pi127;
  assign n1237 = ~n522 & n1236;
  assign n1238 = pi140 & n1237;
  assign n1239 = ~n468 & ~n1238;
  assign n1240 = ~pi042 & n1239;
  assign n1241 = pi127 & ~n1235;
  assign n1242 = pi040 & ~n1241;
  assign po123 = ~n1240 | ~n1242;
  assign n1244 = pi127 & pi140;
  assign n1245 = ~pi126 & ~n522;
  assign n1246 = n1244 & n1245;
  assign n1247 = n520 & ~n522;
  assign n1248 = ~pi128 & pi140;
  assign n1249 = n1247 & n1248;
  assign n1250 = ~n468 & ~n1249;
  assign n1251 = ~pi042 & n1250;
  assign n1252 = pi128 & ~n1246;
  assign n1253 = pi040 & ~n1252;
  assign po124 = ~n1251 | ~n1253;
  assign n1255 = ~pi129 & pi140;
  assign n1256 = pi128 & n1255;
  assign n1257 = pi128 & pi140;
  assign n1258 = pi127 & n1257;
  assign n1259 = n1245 & n1258;
  assign n1260 = pi039 & n461;
  assign n1261 = ~n461 & n1259;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = pi129 & ~n461;
  assign n1264 = ~pi129 & ~n461;
  assign n1265 = ~pi038 & ~n890;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1263 & ~n1266;
  assign n1268 = n1262 & ~n1267;
  assign n1269 = ~n468 & n1256;
  assign n1270 = n1247 & n1269;
  assign n1271 = pi039 & ~n1259;
  assign n1272 = pi129 & n1271;
  assign n1273 = ~n1270 & ~n1272;
  assign n1274 = ~n1268 & n1273;
  assign po125 = n481 & ~n1274;
  assign n1276 = ~pi130 & pi140;
  assign n1277 = ~pi129 & n1276;
  assign n1278 = pi040 & n405;
  assign n1279 = n1277 & n1278;
  assign n1280 = ~pi042 & n1245;
  assign n1281 = ~pi042 & pi130;
  assign n1282 = n520 & n1256;
  assign n1283 = ~n522 & n1282;
  assign n1284 = ~n468 & ~n1283;
  assign n1285 = ~pi039 & pi040;
  assign n1286 = pi038 & n1285;
  assign n1287 = n978 & n1286;
  assign n1288 = n1281 & n1284;
  assign n1289 = pi040 & n1288;
  assign n1290 = ~n468 & n1280;
  assign n1291 = n1279 & n1290;
  assign n1292 = ~n1289 & ~n1291;
  assign po126 = n1287 | ~n1292;
  assign n1294 = pi127 & n430;
  assign n1295 = ~pi131 & pi140;
  assign n1296 = ~pi130 & n1295;
  assign n1297 = pi040 & n1294;
  assign n1298 = n1296 & n1297;
  assign n1299 = ~pi042 & pi131;
  assign n1300 = ~pi126 & n405;
  assign n1301 = n1277 & n1300;
  assign n1302 = ~n522 & n1301;
  assign n1303 = ~n468 & ~n1302;
  assign n1304 = ~pi038 & n1285;
  assign n1305 = n978 & n1304;
  assign n1306 = n1299 & n1303;
  assign n1307 = pi040 & n1306;
  assign n1308 = n1290 & n1298;
  assign n1309 = ~n1307 & ~n1308;
  assign po127 = n1305 | ~n1309;
  assign n1311 = ~pi042 & ~pi057;
  assign n1312 = pi132 & pi139;
  assign n1313 = ~pi132 & ~n1194;
  assign n1314 = ~n990 & n1312;
  assign n1315 = ~n995 & n1314;
  assign n1316 = ~n1313 & ~n1315;
  assign n1317 = n1311 & n1316;
  assign n1318 = ~pi039 & n978;
  assign n1319 = ~n1317 & ~n1318;
  assign po128 = pi040 & ~n1319;
  assign n1321 = ~pi132 & pi139;
  assign n1322 = ~n990 & ~n995;
  assign n1323 = n1321 & n1322;
  assign n1324 = ~pi133 & pi139;
  assign n1325 = ~pi132 & n1324;
  assign n1326 = ~n990 & n1325;
  assign n1327 = ~n995 & n1326;
  assign n1328 = ~n468 & ~n1327;
  assign n1329 = n1311 & n1328;
  assign n1330 = pi133 & ~n1323;
  assign n1331 = pi040 & ~n1330;
  assign po129 = ~n1329 | ~n1331;
  assign n1333 = pi133 & pi139;
  assign n1334 = ~pi132 & n1333;
  assign n1335 = n1322 & n1334;
  assign n1336 = ~pi132 & ~n995;
  assign n1337 = ~pi134 & pi139;
  assign n1338 = pi133 & n1337;
  assign n1339 = n1336 & n1338;
  assign n1340 = ~n990 & n1339;
  assign n1341 = ~n468 & ~n1340;
  assign n1342 = n1311 & n1341;
  assign n1343 = pi134 & ~n1335;
  assign n1344 = pi040 & ~n1343;
  assign po130 = ~n1342 | ~n1344;
  assign n1346 = ~pi132 & pi133;
  assign n1347 = ~pi057 & n1346;
  assign n1348 = ~pi135 & pi139;
  assign n1349 = pi134 & n1348;
  assign n1350 = pi040 & n1347;
  assign n1351 = n1349 & n1350;
  assign n1352 = ~pi042 & n1322;
  assign n1353 = ~pi057 & pi135;
  assign n1354 = ~pi042 & n1353;
  assign n1355 = pi134 & pi139;
  assign n1356 = pi133 & n1355;
  assign n1357 = n1336 & n1356;
  assign n1358 = ~n990 & n1357;
  assign n1359 = ~n468 & ~n1358;
  assign n1360 = pi038 & ~n890;
  assign n1361 = ~pi039 & ~n1360;
  assign n1362 = pi040 & n1361;
  assign n1363 = n978 & n1362;
  assign n1364 = n1354 & n1359;
  assign n1365 = pi040 & n1364;
  assign n1366 = ~n468 & n1352;
  assign n1367 = n1351 & n1366;
  assign n1368 = ~n1365 & ~n1367;
  assign po131 = n1363 | ~n1368;
  assign n1370 = ~pi057 & ~n995;
  assign n1371 = ~pi132 & n435;
  assign n1372 = ~pi136 & pi139;
  assign n1373 = ~pi135 & n1372;
  assign n1374 = n1370 & n1371;
  assign n1375 = n1373 & n1374;
  assign n1376 = ~pi057 & pi136;
  assign n1377 = ~pi042 & n1376;
  assign n1378 = ~n995 & n1346;
  assign n1379 = n1349 & n1378;
  assign n1380 = ~n990 & n1379;
  assign n1381 = ~n468 & ~n1380;
  assign n1382 = n1377 & n1381;
  assign n1383 = pi040 & n1382;
  assign n1384 = ~n468 & n992;
  assign n1385 = n1375 & n1384;
  assign n1386 = ~n1383 & ~n1385;
  assign po132 = n1287 | ~n1386;
  assign n1388 = ~pi042 & ~n522;
  assign n1389 = pi040 & n1388;
  assign n1390 = pi064 & pi137;
  assign n1391 = n1389 & ~n1390;
  assign n1392 = ~pi064 & ~pi137;
  assign n1393 = n1391 & ~n1392;
  assign po133 = pi140 & n1393;
  assign n1395 = pi139 & pi142;
  assign n1396 = ~pi138 & n1395;
  assign n1397 = n481 & n1396;
  assign n1398 = ~n990 & n1370;
  assign n1399 = ~pi057 & pi138;
  assign n1400 = ~pi042 & n1399;
  assign n1401 = ~pi046 & ~pi062;
  assign n1402 = pi047 & pi062;
  assign n1403 = ~pi061 & ~n1402;
  assign n1404 = ~n1401 & ~n1403;
  assign n1405 = pi043 & ~pi059;
  assign n1406 = n999 & n1405;
  assign n1407 = ~pi059 & n460;
  assign n1408 = pi044 & ~pi060;
  assign n1409 = n460 & n1408;
  assign n1410 = ~n995 & ~n1001;
  assign n1411 = ~n990 & ~n1000;
  assign n1412 = n1410 & n1411;
  assign n1413 = n1395 & n1412;
  assign n1414 = ~pi045 & n1407;
  assign n1415 = ~pi058 & n1414;
  assign n1416 = pi059 & ~n1409;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = n1413 & n1417;
  assign n1419 = pi058 & n1406;
  assign n1420 = pi058 & ~n1406;
  assign n1421 = n458 & ~n1404;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1419 & ~n1422;
  assign n1424 = n1418 & ~n1423;
  assign n1425 = n1400 & ~n1424;
  assign n1426 = pi040 & n1425;
  assign n1427 = ~n1215 & n1398;
  assign n1428 = n1397 & n1427;
  assign po134 = n1426 | n1428;
  assign n1430 = ~pi042 & pi063;
  assign n1431 = pi040 & n1430;
  assign n1432 = n1294 & n1431;
  assign po135 = n406 & n1432;
  assign po136 = pi063 & n1389;
  assign n1435 = ~n440 & ~n445;
  assign n1436 = ~n995 & n1435;
  assign n1437 = ~n444 & ~n450;
  assign n1438 = n1436 & n1437;
  assign n1439 = pi142 & ~n449;
  assign n1440 = n1438 & n1439;
  assign n1441 = n990 & ~n1440;
  assign n1442 = ~pi042 & ~n1441;
  assign n1443 = pi040 & n1442;
  assign n1444 = ~n453 & ~n1440;
  assign po137 = n1443 & ~n1444;
  assign po138 = pi139 & n992;
  assign po000 = ~pi057;
  assign po045 = ~pi058;
  assign po046 = ~pi059;
  assign po047 = ~pi060;
  assign po048 = ~pi061;
  assign po049 = ~pi062;
  assign po005 = pi123;
  assign po006 = pi124;
  assign po024 = pi141;
  assign po031 = po030;
  assign po032 = po030;
  assign po033 = po030;
  assign po034 = po030;
  assign po050 = pi139;
endmodule



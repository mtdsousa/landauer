// Benchmark "pair" written by ABC on Sun Apr 22 21:43:11 2018

module pair ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136;
  wire n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554, n555, n556, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n652, n653, n654, n656, n657, n658, n659, n660, n662,
    n663, n664, n665, n666, n668, n669, n670, n671, n672, n673, n675, n676,
    n677, n678, n679, n681, n682, n683, n684, n685, n687, n688, n689, n690,
    n691, n692, n693, n695, n696, n697, n698, n699, n701, n702, n703, n705,
    n706, n707, n709, n710, n711, n712, n713, n714, n715, n716, n718, n719,
    n720, n721, n722, n723, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n746, n747, n748, n749, n750, n751, n752, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n942, n943, n945, n946, n948, n949, n950, n951, n952, n953,
    n954, n955, n957, n958, n959, n960, n961, n962, n963, n965, n966, n968,
    n969, n970, n971, n972, n973, n974, n975, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n987, n988, n989, n990, n991, n992, n993, n994,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1042, n1043, n1044, n1046, n1047, n1048, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1091, n1092, n1093, n1094, n1095,
    n1096, n1098, n1099, n1100, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1213, n1214, n1215, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1261, n1262, n1263, n1264, n1265, n1266, n1268, n1269, n1270, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1533, n1534, n1536, n1537, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1559, n1560, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1648, n1649, n1650, n1652, n1653, n1654, n1655, n1656,
    n1658, n1659, n1660, n1661, n1662, n1664, n1665, n1666, n1667, n1668,
    n1669, n1671, n1672, n1673, n1674, n1675, n1677, n1678, n1679, n1680,
    n1681, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1691, n1692,
    n1693, n1694, n1695, n1697, n1698, n1699, n1701, n1702, n1703, n1705,
    n1706, n1707, n1708, n1709, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1719, n1720, n1721, n1722, n1723, n1725, n1726, n1727, n1728,
    n1730, n1731, n1732, n1734, n1735, n1736, n1737, n1738, n1739, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809;
  assign n311 = pi022 & pi049;
  assign n312 = pi021 & pi054;
  assign n313 = pi020 & pi083;
  assign n314 = pi019 & pi086;
  assign n315 = ~n311 & ~n312;
  assign n316 = ~n313 & ~n314;
  assign n317 = n315 & n316;
  assign n318 = pi018 & pi091;
  assign n319 = pi017 & pi071;
  assign n320 = pi016 & pi074;
  assign n321 = pi015 & pi077;
  assign n322 = ~n318 & ~n319;
  assign n323 = ~n320 & ~n321;
  assign n324 = n322 & n323;
  assign n325 = pi014 & pi096;
  assign n326 = pi013 & pi103;
  assign n327 = pi012 & pi107;
  assign n328 = ~n325 & ~n326;
  assign n329 = ~n327 & n328;
  assign n330 = n317 & n324;
  assign po000 = ~n329 | ~n330;
  assign n332 = pi022 & pi048;
  assign n333 = pi021 & pi053;
  assign n334 = pi020 & pi080;
  assign n335 = pi019 & pi085;
  assign n336 = ~n332 & ~n333;
  assign n337 = ~n334 & ~n335;
  assign n338 = n336 & n337;
  assign n339 = pi018 & pi089;
  assign n340 = pi017 & pi070;
  assign n341 = pi016 & pi073;
  assign n342 = pi015 & pi076;
  assign n343 = ~n339 & ~n340;
  assign n344 = ~n341 & ~n342;
  assign n345 = n343 & n344;
  assign n346 = pi014 & pi095;
  assign n347 = pi013 & pi102;
  assign n348 = pi012 & pi106;
  assign n349 = ~n346 & ~n347;
  assign n350 = ~n348 & n349;
  assign n351 = n338 & n345;
  assign po001 = ~n350 | ~n351;
  assign n353 = pi022 & pi047;
  assign n354 = pi021 & pi052;
  assign n355 = pi020 & pi079;
  assign n356 = pi019 & pi084;
  assign n357 = ~n353 & ~n354;
  assign n358 = ~n355 & ~n356;
  assign n359 = n357 & n358;
  assign n360 = pi018 & pi088;
  assign n361 = pi017 & pi069;
  assign n362 = pi016 & pi072;
  assign n363 = pi015 & pi075;
  assign n364 = ~n360 & ~n361;
  assign n365 = ~n362 & ~n363;
  assign n366 = n364 & n365;
  assign n367 = pi014 & pi094;
  assign n368 = pi013 & pi101;
  assign n369 = pi012 & pi105;
  assign n370 = ~n367 & ~n368;
  assign n371 = ~n369 & n370;
  assign n372 = n359 & n366;
  assign po002 = ~n371 | ~n372;
  assign n374 = pi022 & pi046;
  assign n375 = pi021 & pi051;
  assign n376 = pi020 & pi078;
  assign n377 = pi019 & pi082;
  assign n378 = ~n374 & ~n375;
  assign n379 = ~n376 & ~n377;
  assign n380 = n378 & n379;
  assign n381 = pi018 & pi087;
  assign n382 = pi017 & pi063;
  assign n383 = pi016 & pi068;
  assign n384 = pi015 & pi066;
  assign n385 = ~n381 & ~n382;
  assign n386 = ~n383 & ~n384;
  assign n387 = n385 & n386;
  assign n388 = pi014 & pi093;
  assign n389 = pi013 & pi100;
  assign n390 = pi012 & pi104;
  assign n391 = ~n388 & ~n389;
  assign n392 = ~n390 & n391;
  assign n393 = n380 & n387;
  assign po003 = ~n392 | ~n393;
  assign n395 = pi022 & pi062;
  assign n396 = pi021 & pi050;
  assign n397 = ~pi058 & ~pi059;
  assign n398 = pi055 & ~pi056;
  assign n399 = ~pi061 & pi065;
  assign n400 = ~pi060 & ~pi065;
  assign n401 = ~n399 & ~n400;
  assign n402 = pi060 & ~n401;
  assign n403 = ~n398 & n402;
  assign n404 = n398 & ~n402;
  assign n405 = ~n403 & ~n404;
  assign n406 = n397 & ~n405;
  assign n407 = n402 & n406;
  assign n408 = ~pi058 & ~n407;
  assign n409 = n398 & ~n405;
  assign n410 = n397 & n409;
  assign po021 = pi059 | n410;
  assign n412 = ~pi057 & ~po021;
  assign n413 = ~pi048 & ~pi049;
  assign n414 = ~pi050 & n413;
  assign n415 = ~pi051 & n414;
  assign n416 = ~pi052 & n415;
  assign n417 = ~pi053 & n416;
  assign n418 = ~pi047 & n417;
  assign n419 = ~pi054 & n418;
  assign n420 = ~pi046 & n419;
  assign n421 = n408 & n412;
  assign n422 = n420 & ~n421;
  assign n423 = pi062 & pi063;
  assign n424 = ~pi001 & ~pi064;
  assign n425 = n423 & n424;
  assign n426 = ~pi062 & ~pi063;
  assign n427 = ~pi064 & n426;
  assign po029 = pi001 | n427;
  assign n429 = n422 & po029;
  assign n430 = ~pi046 & pi068;
  assign n431 = n425 & ~n430;
  assign n432 = ~n429 & ~n431;
  assign n433 = ~pi005 & n432;
  assign n434 = pi020 & n433;
  assign n435 = pi019 & pi081;
  assign n436 = ~n395 & ~n396;
  assign n437 = ~n434 & ~n435;
  assign n438 = n436 & n437;
  assign n439 = ~pi011 & pi067;
  assign n440 = pi078 & pi079;
  assign n441 = pi080 & n440;
  assign n442 = ~n439 & ~n441;
  assign n443 = pi083 & ~n442;
  assign n444 = ~pi011 & ~pi066;
  assign n445 = ~n443 & n444;
  assign n446 = pi081 & ~n445;
  assign n447 = pi090 & n446;
  assign n448 = pi018 & n447;
  assign n449 = pi017 & pi064;
  assign n450 = ~pi062 & pi063;
  assign n451 = ~pi064 & n450;
  assign n452 = ~pi001 & n451;
  assign n453 = ~pi001 & ~n452;
  assign n454 = pi016 & ~n453;
  assign n455 = pi015 & pi067;
  assign n456 = ~n448 & ~n449;
  assign n457 = ~n454 & ~n455;
  assign n458 = n456 & n457;
  assign n459 = pi106 & pi107;
  assign n460 = pi105 & n459;
  assign n461 = pi014 & n460;
  assign n462 = pi013 & pi099;
  assign n463 = pi101 & ~pi102;
  assign n464 = ~pi103 & n463;
  assign n465 = ~pi104 & ~pi105;
  assign n466 = ~pi106 & ~pi107;
  assign n467 = n465 & n466;
  assign n468 = n464 & n467;
  assign n469 = pi012 & n468;
  assign n470 = ~n461 & ~n462;
  assign n471 = ~n469 & n470;
  assign n472 = n438 & n458;
  assign po004 = ~n471 | ~n472;
  assign n474 = pi045 & pi149;
  assign n475 = pi044 & pi154;
  assign n476 = pi043 & pi137;
  assign n477 = pi042 & pi140;
  assign n478 = ~n474 & ~n475;
  assign n479 = ~n476 & ~n477;
  assign n480 = n478 & n479;
  assign n481 = pi041 & pi145;
  assign n482 = pi040 & pi125;
  assign n483 = pi039 & pi128;
  assign n484 = pi038 & pi131;
  assign n485 = ~n481 & ~n482;
  assign n486 = ~n483 & ~n484;
  assign n487 = n485 & n486;
  assign n488 = pi037 & pi111;
  assign n489 = pi036 & pi118;
  assign n490 = pi035 & pi122;
  assign n491 = ~n488 & ~n489;
  assign n492 = ~n490 & n491;
  assign n493 = n480 & n487;
  assign po005 = ~n492 | ~n493;
  assign n495 = pi045 & pi148;
  assign n496 = pi044 & pi153;
  assign n497 = pi043 & pi134;
  assign n498 = pi042 & pi139;
  assign n499 = ~n495 & ~n496;
  assign n500 = ~n497 & ~n498;
  assign n501 = n499 & n500;
  assign n502 = pi041 & pi143;
  assign n503 = pi040 & pi124;
  assign n504 = pi039 & pi127;
  assign n505 = pi038 & pi130;
  assign n506 = ~n502 & ~n503;
  assign n507 = ~n504 & ~n505;
  assign n508 = n506 & n507;
  assign n509 = pi037 & pi110;
  assign n510 = pi036 & pi117;
  assign n511 = pi035 & pi121;
  assign n512 = ~n509 & ~n510;
  assign n513 = ~n511 & n512;
  assign n514 = n501 & n508;
  assign po006 = ~n513 | ~n514;
  assign n516 = pi045 & pi147;
  assign n517 = pi044 & pi152;
  assign n518 = pi043 & pi133;
  assign n519 = pi042 & pi138;
  assign n520 = ~n516 & ~n517;
  assign n521 = ~n518 & ~n519;
  assign n522 = n520 & n521;
  assign n523 = pi041 & pi142;
  assign n524 = pi040 & pi123;
  assign n525 = pi039 & pi126;
  assign n526 = pi038 & pi129;
  assign n527 = ~n523 & ~n524;
  assign n528 = ~n525 & ~n526;
  assign n529 = n527 & n528;
  assign n530 = pi037 & pi109;
  assign n531 = pi036 & pi116;
  assign n532 = pi035 & pi120;
  assign n533 = ~n530 & ~n531;
  assign n534 = ~n532 & n533;
  assign n535 = n522 & n529;
  assign po007 = ~n534 | ~n535;
  assign n537 = pi045 & pi146;
  assign n538 = pi044 & pi151;
  assign n539 = pi043 & pi132;
  assign n540 = pi042 & pi136;
  assign n541 = ~n537 & ~n538;
  assign n542 = ~n539 & ~n540;
  assign n543 = n541 & n542;
  assign n544 = pi041 & pi141;
  assign n545 = pi040 & pi167;
  assign n546 = pi039 & pi172;
  assign n547 = pi038 & pi170;
  assign n548 = ~n544 & ~n545;
  assign n549 = ~n546 & ~n547;
  assign n550 = n548 & n549;
  assign n551 = pi037 & pi108;
  assign n552 = pi036 & pi115;
  assign n553 = pi035 & pi119;
  assign n554 = ~n551 & ~n552;
  assign n555 = ~n553 & n554;
  assign n556 = n543 & n550;
  assign po008 = ~n555 | ~n556;
  assign n558 = pi045 & pi166;
  assign n559 = pi044 & pi150;
  assign n560 = ~pi164 & pi165;
  assign n561 = ~pi158 & ~pi159;
  assign n562 = pi155 & ~pi156;
  assign n563 = ~pi163 & pi169;
  assign n564 = ~pi161 & ~pi169;
  assign n565 = ~n563 & ~n564;
  assign n566 = pi161 & ~n565;
  assign n567 = ~n562 & n566;
  assign n568 = n562 & ~n566;
  assign n569 = ~n567 & ~n568;
  assign n570 = n561 & ~n569;
  assign n571 = n566 & n570;
  assign n572 = ~pi158 & ~n571;
  assign n573 = n562 & ~n569;
  assign n574 = n561 & n573;
  assign po121 = pi159 | n574;
  assign n576 = ~pi157 & ~po121;
  assign n577 = ~pi148 & ~pi149;
  assign n578 = ~pi150 & n577;
  assign n579 = ~pi151 & n578;
  assign n580 = ~pi152 & n579;
  assign n581 = ~pi153 & n580;
  assign n582 = ~pi147 & n581;
  assign n583 = ~pi154 & n582;
  assign n584 = ~pi146 & n583;
  assign n585 = n572 & n576;
  assign n586 = n584 & ~n585;
  assign n587 = ~pi166 & ~pi167;
  assign n588 = ~pi168 & n587;
  assign po133 = pi024 | n588;
  assign n590 = n586 & po133;
  assign n591 = ~pi146 & pi172;
  assign n592 = n560 & ~n591;
  assign n593 = ~n590 & ~n592;
  assign n594 = ~pi028 & n593;
  assign n595 = pi043 & n594;
  assign n596 = pi042 & pi135;
  assign n597 = ~n558 & ~n559;
  assign n598 = ~n595 & ~n596;
  assign n599 = n597 & n598;
  assign n600 = ~pi034 & pi171;
  assign n601 = pi132 & pi133;
  assign n602 = pi134 & n601;
  assign n603 = ~n600 & ~n602;
  assign n604 = pi137 & ~n603;
  assign n605 = ~pi034 & ~pi170;
  assign n606 = ~n604 & n605;
  assign n607 = pi135 & ~n606;
  assign n608 = pi144 & n607;
  assign n609 = pi041 & n608;
  assign n610 = pi040 & pi168;
  assign n611 = ~pi166 & pi167;
  assign n612 = ~pi168 & n611;
  assign n613 = ~pi024 & n612;
  assign n614 = ~pi024 & ~n613;
  assign n615 = pi039 & ~n614;
  assign n616 = pi038 & pi171;
  assign n617 = ~n609 & ~n610;
  assign n618 = ~n615 & ~n616;
  assign n619 = n617 & n618;
  assign n620 = pi118 & pi119;
  assign n621 = pi121 & pi122;
  assign n622 = pi120 & n621;
  assign n623 = n620 & n622;
  assign n624 = pi037 & n623;
  assign n625 = pi036 & pi114;
  assign n626 = pi116 & ~pi117;
  assign n627 = ~pi118 & n626;
  assign n628 = ~pi119 & ~pi120;
  assign n629 = ~pi121 & ~pi122;
  assign n630 = n628 & n629;
  assign n631 = n627 & n630;
  assign n632 = pi035 & n631;
  assign n633 = ~n624 & ~n625;
  assign n634 = ~n632 & n633;
  assign n635 = n599 & n619;
  assign po009 = ~n634 | ~n635;
  assign n637 = pi068 & n425;
  assign n638 = n412 & ~n637;
  assign n639 = n408 & n638;
  assign n640 = ~pi046 & n639;
  assign n641 = pi046 & ~n639;
  assign n642 = ~n640 & ~n641;
  assign n643 = n421 & po029;
  assign n644 = pi046 & n637;
  assign n645 = ~pi063 & pi064;
  assign n646 = ~pi001 & pi062;
  assign n647 = n645 & n646;
  assign n648 = ~n643 & ~n644;
  assign n649 = ~pi001 & ~n647;
  assign n650 = n648 & n649;
  assign po010 = n642 & n650;
  assign n652 = ~pi047 & ~n641;
  assign n653 = pi047 & n641;
  assign n654 = ~n652 & ~n653;
  assign po011 = n650 & n654;
  assign n656 = pi046 & pi047;
  assign n657 = ~n639 & n656;
  assign n658 = ~pi048 & ~n657;
  assign n659 = pi048 & n657;
  assign n660 = ~n658 & ~n659;
  assign po012 = n650 & n660;
  assign n662 = pi048 & n656;
  assign n663 = ~n639 & n662;
  assign n664 = ~pi049 & ~n663;
  assign n665 = pi049 & n663;
  assign n666 = ~n664 & ~n665;
  assign po013 = n650 & n666;
  assign n668 = pi048 & pi049;
  assign n669 = n656 & n668;
  assign n670 = ~n639 & n669;
  assign n671 = ~pi050 & ~n670;
  assign n672 = pi050 & n670;
  assign n673 = ~n671 & ~n672;
  assign po014 = n650 & n673;
  assign n675 = pi050 & n669;
  assign n676 = ~n639 & n675;
  assign n677 = ~pi051 & ~n676;
  assign n678 = pi051 & n676;
  assign n679 = ~n677 & ~n678;
  assign po015 = n650 & n679;
  assign n681 = pi051 & n675;
  assign n682 = ~n639 & n681;
  assign n683 = ~pi052 & ~n682;
  assign n684 = pi052 & n682;
  assign n685 = ~n683 & ~n684;
  assign po016 = n650 & n685;
  assign n687 = pi050 & pi051;
  assign n688 = pi052 & n687;
  assign n689 = n669 & n688;
  assign n690 = ~n639 & n689;
  assign n691 = ~pi053 & ~n690;
  assign n692 = pi053 & n690;
  assign n693 = ~n691 & ~n692;
  assign po017 = n650 & n693;
  assign n695 = pi053 & ~n639;
  assign n696 = n689 & n695;
  assign n697 = pi054 & n696;
  assign n698 = ~pi054 & ~n696;
  assign n699 = ~n697 & ~n698;
  assign po018 = n650 & n699;
  assign n701 = pi058 & n398;
  assign n702 = n649 & ~n701;
  assign n703 = pi058 & n702;
  assign po022 = n407 | n703;
  assign n705 = pi059 & n402;
  assign n706 = n649 & ~n705;
  assign n707 = pi059 & n706;
  assign po023 = n410 | n707;
  assign n709 = pi060 & n447;
  assign n710 = ~pi060 & ~n447;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~pi001 & n711;
  assign n713 = pi062 & ~pi063;
  assign n714 = ~pi064 & n713;
  assign n715 = ~pi001 & n714;
  assign n716 = ~n647 & ~n715;
  assign po024 = n712 | ~n716;
  assign n718 = n398 & ~n468;
  assign n719 = n460 & n718;
  assign n720 = n425 & ~n719;
  assign n721 = n398 & n452;
  assign n722 = ~n715 & ~n720;
  assign n723 = ~n721 & n722;
  assign po026 = ~pi001 & ~n723;
  assign n725 = pi068 & ~n697;
  assign n726 = pi068 & n697;
  assign n727 = ~pi054 & ~n726;
  assign n728 = ~n725 & ~n727;
  assign n729 = ~pi002 & ~n728;
  assign n730 = po029 & ~n729;
  assign n731 = n425 & n468;
  assign n732 = ~n730 & ~n731;
  assign n733 = pi064 & n426;
  assign n734 = ~pi001 & n733;
  assign n735 = ~n452 & n732;
  assign n736 = ~n734 & n735;
  assign n737 = pi064 & n423;
  assign n738 = ~pi001 & n737;
  assign n739 = pi063 & pi064;
  assign n740 = ~n398 & ~n468;
  assign n741 = n425 & n740;
  assign n742 = ~n739 & ~n741;
  assign n743 = ~n738 & n742;
  assign n744 = n736 & n743;
  assign po027 = ~pi001 & ~n744;
  assign n746 = ~n731 & ~n734;
  assign n747 = ~n715 & n746;
  assign n748 = n398 & n425;
  assign n749 = n460 & ~n468;
  assign n750 = n748 & n749;
  assign n751 = ~n738 & ~n750;
  assign n752 = n747 & n751;
  assign po028 = ~pi001 & ~n752;
  assign n754 = pi067 & pi068;
  assign n755 = ~pi066 & ~n754;
  assign n756 = ~pi067 & ~pi068;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~pi066 & n756;
  assign n759 = ~pi001 & ~n758;
  assign n760 = ~n757 & n759;
  assign n761 = ~pi004 & ~n738;
  assign n762 = ~pi003 & ~n734;
  assign n763 = pi067 & ~n762;
  assign n764 = pi068 & ~n761;
  assign n765 = ~pi066 & ~n764;
  assign n766 = ~pi068 & ~n761;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n763 & ~n767;
  assign n769 = ~n762 & ~n764;
  assign n770 = ~pi067 & n769;
  assign n771 = ~n768 & ~n770;
  assign po030 = ~n760 | n771;
  assign n773 = pi068 & ~n762;
  assign n774 = pi067 & n761;
  assign n775 = ~pi066 & ~n774;
  assign n776 = ~pi067 & n761;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~n773 & ~n777;
  assign n779 = pi066 & ~n761;
  assign n780 = ~n762 & ~n779;
  assign n781 = ~pi068 & n780;
  assign n782 = ~n778 & ~n781;
  assign po031 = n760 & n782;
  assign n784 = pi066 & ~n762;
  assign n785 = ~pi068 & n761;
  assign n786 = pi068 & n761;
  assign n787 = ~pi067 & ~n786;
  assign n788 = ~n785 & ~n787;
  assign n789 = ~n784 & ~n788;
  assign n790 = pi067 & ~n761;
  assign n791 = ~n762 & ~n790;
  assign n792 = ~pi066 & n791;
  assign n793 = ~n789 & ~n792;
  assign po032 = n760 & n793;
  assign n795 = pi046 & n419;
  assign n796 = po029 & n795;
  assign n797 = ~n715 & ~n796;
  assign n798 = ~pi046 & pi047;
  assign n799 = pi067 & n414;
  assign n800 = pi068 & n417;
  assign n801 = pi066 & n413;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~n799 & n802;
  assign n804 = n798 & ~n803;
  assign n805 = po029 & n804;
  assign n806 = ~pi007 & ~n805;
  assign n807 = ~pi069 & ~n806;
  assign n808 = pi069 & n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = n797 & n809;
  assign n811 = n797 & ~n809;
  assign n812 = ~pi099 & ~n811;
  assign n813 = ~n810 & ~n812;
  assign po033 = ~pi001 & n813;
  assign n815 = ~pi008 & n412;
  assign n816 = ~pi069 & ~n815;
  assign n817 = pi069 & n815;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n806 & n818;
  assign n820 = ~pi070 & n819;
  assign n821 = pi070 & ~n819;
  assign n822 = ~n820 & ~n821;
  assign n823 = n797 & n822;
  assign n824 = n797 & ~n822;
  assign n825 = ~pi100 & ~n824;
  assign n826 = ~n823 & ~n825;
  assign po034 = ~pi001 & n826;
  assign n828 = ~pi069 & ~pi070;
  assign n829 = pi069 & pi070;
  assign n830 = ~n815 & n829;
  assign n831 = ~n828 & ~n830;
  assign n832 = ~n815 & ~n829;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n806 & n833;
  assign n835 = ~pi071 & n834;
  assign n836 = pi071 & ~n834;
  assign n837 = ~n835 & ~n836;
  assign n838 = n797 & n837;
  assign n839 = n797 & ~n837;
  assign n840 = ~pi101 & ~n839;
  assign n841 = ~n838 & ~n840;
  assign po035 = ~pi001 & n841;
  assign n843 = ~pi071 & n828;
  assign n844 = ~pi010 & ~n843;
  assign n845 = pi071 & n829;
  assign n846 = ~pi010 & ~n845;
  assign n847 = ~n815 & ~n846;
  assign n848 = n844 & ~n847;
  assign n849 = ~n815 & n846;
  assign n850 = ~n848 & ~n849;
  assign n851 = ~n806 & n850;
  assign n852 = ~pi072 & n851;
  assign n853 = pi072 & ~n851;
  assign n854 = ~n852 & ~n853;
  assign n855 = n797 & n854;
  assign n856 = n797 & ~n854;
  assign n857 = ~pi102 & ~n856;
  assign n858 = ~n855 & ~n857;
  assign po036 = pi001 | n858;
  assign n860 = ~pi072 & ~n844;
  assign n861 = pi072 & ~n846;
  assign n862 = ~n815 & n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = ~n815 & ~n861;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~n806 & n865;
  assign n867 = ~pi073 & n866;
  assign n868 = pi073 & ~n866;
  assign n869 = ~n867 & ~n868;
  assign n870 = n797 & n869;
  assign n871 = n797 & ~n869;
  assign n872 = ~pi103 & ~n871;
  assign n873 = ~n870 & ~n872;
  assign po037 = pi001 | n873;
  assign n875 = ~pi073 & n860;
  assign n876 = pi072 & pi073;
  assign n877 = ~n846 & n876;
  assign n878 = ~n815 & n877;
  assign n879 = ~n875 & ~n878;
  assign n880 = ~n815 & ~n877;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n806 & n881;
  assign n883 = ~pi074 & n882;
  assign n884 = pi074 & ~n882;
  assign n885 = ~n883 & ~n884;
  assign n886 = n797 & n885;
  assign n887 = n797 & ~n885;
  assign n888 = ~pi104 & ~n887;
  assign n889 = ~n886 & ~n888;
  assign po038 = pi001 | n889;
  assign n891 = ~pi073 & ~pi074;
  assign n892 = n860 & n891;
  assign n893 = ~pi010 & ~n892;
  assign n894 = pi073 & pi074;
  assign n895 = n861 & n894;
  assign n896 = ~pi010 & ~n895;
  assign n897 = ~n815 & ~n896;
  assign n898 = n893 & ~n897;
  assign n899 = ~n815 & n896;
  assign n900 = ~n898 & ~n899;
  assign n901 = ~n806 & n900;
  assign n902 = ~pi075 & n901;
  assign n903 = pi075 & ~n901;
  assign n904 = ~n902 & ~n903;
  assign n905 = n797 & n904;
  assign n906 = n797 & ~n904;
  assign n907 = ~pi105 & ~n906;
  assign n908 = ~n905 & ~n907;
  assign po039 = ~pi001 & n908;
  assign n910 = ~pi075 & ~n893;
  assign n911 = pi075 & ~n896;
  assign n912 = ~n815 & n911;
  assign n913 = ~n910 & ~n912;
  assign n914 = ~n815 & ~n911;
  assign n915 = ~n913 & ~n914;
  assign n916 = ~n806 & n915;
  assign n917 = ~pi076 & n916;
  assign n918 = pi076 & ~n916;
  assign n919 = ~n917 & ~n918;
  assign n920 = n797 & n919;
  assign n921 = n797 & ~n919;
  assign n922 = ~pi106 & ~n921;
  assign n923 = ~n920 & ~n922;
  assign po040 = pi001 | n923;
  assign n925 = ~pi076 & n910;
  assign n926 = pi075 & pi076;
  assign n927 = ~n896 & n926;
  assign n928 = ~n815 & n927;
  assign n929 = ~n925 & ~n928;
  assign n930 = ~n815 & ~n927;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n806 & n931;
  assign n933 = ~pi077 & n932;
  assign n934 = pi077 & ~n932;
  assign n935 = ~n933 & ~n934;
  assign n936 = n797 & n935;
  assign n937 = n797 & ~n935;
  assign n938 = ~pi107 & ~n937;
  assign n939 = ~n936 & ~n938;
  assign po041 = pi001 | n939;
  assign po042 = pi001 | ~pi078;
  assign n942 = ~pi078 & ~pi079;
  assign n943 = ~n440 & ~n942;
  assign po043 = pi001 | n943;
  assign n945 = ~pi080 & ~n440;
  assign n946 = ~n441 & ~n945;
  assign po044 = pi001 | n946;
  assign n948 = ~n447 & ~n647;
  assign n949 = ~pi081 & ~n445;
  assign n950 = pi081 & n445;
  assign n951 = ~n949 & ~n950;
  assign n952 = n948 & ~n951;
  assign n953 = ~pi069 & ~n952;
  assign n954 = n948 & n951;
  assign n955 = ~n953 & ~n954;
  assign po045 = pi001 | n955;
  assign n957 = ~pi082 & n446;
  assign n958 = pi082 & ~n446;
  assign n959 = ~n957 & ~n958;
  assign n960 = n948 & ~n959;
  assign n961 = ~pi070 & ~n960;
  assign n962 = n948 & n959;
  assign n963 = ~n961 & ~n962;
  assign po046 = pi001 | n963;
  assign n965 = ~pi083 & n442;
  assign n966 = ~n443 & ~n965;
  assign po047 = pi001 | n966;
  assign n968 = pi082 & n446;
  assign n969 = ~pi084 & n968;
  assign n970 = pi084 & ~n968;
  assign n971 = ~n969 & ~n970;
  assign n972 = n948 & ~n971;
  assign n973 = ~pi071 & ~n972;
  assign n974 = n948 & n971;
  assign n975 = ~n973 & ~n974;
  assign po048 = pi001 | n975;
  assign n977 = pi082 & pi084;
  assign n978 = n446 & n977;
  assign n979 = ~pi085 & n978;
  assign n980 = pi085 & ~n978;
  assign n981 = ~n979 & ~n980;
  assign n982 = n948 & ~n981;
  assign n983 = ~pi072 & ~n982;
  assign n984 = n948 & n981;
  assign n985 = ~n983 & ~n984;
  assign po049 = pi001 | n985;
  assign n987 = pi085 & n978;
  assign n988 = ~pi086 & n987;
  assign n989 = pi086 & ~n987;
  assign n990 = ~n988 & ~n989;
  assign n991 = n948 & ~n990;
  assign n992 = ~pi073 & ~n991;
  assign n993 = n948 & n990;
  assign n994 = ~n992 & ~n993;
  assign po050 = pi001 | n994;
  assign n996 = pi086 & n987;
  assign n997 = ~pi011 & ~n996;
  assign n998 = ~pi087 & ~n997;
  assign n999 = pi087 & n997;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = n948 & ~n1000;
  assign n1002 = ~pi074 & ~n1001;
  assign n1003 = n948 & n1000;
  assign n1004 = ~n1002 & ~n1003;
  assign po051 = pi001 | n1004;
  assign n1006 = pi087 & ~n997;
  assign n1007 = ~pi088 & n1006;
  assign n1008 = pi088 & ~n1006;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = n948 & ~n1009;
  assign n1011 = ~pi075 & ~n1010;
  assign n1012 = n948 & n1009;
  assign n1013 = ~n1011 & ~n1012;
  assign po052 = pi001 | n1013;
  assign n1015 = pi087 & pi088;
  assign n1016 = ~n997 & n1015;
  assign n1017 = ~pi089 & n1016;
  assign n1018 = pi089 & ~n1016;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n948 & ~n1019;
  assign n1021 = ~pi076 & ~n1020;
  assign n1022 = n948 & n1019;
  assign n1023 = ~n1021 & ~n1022;
  assign po053 = pi001 | n1023;
  assign n1025 = pi089 & pi091;
  assign n1026 = pi088 & n1025;
  assign n1027 = pi086 & pi087;
  assign n1028 = pi085 & n1027;
  assign n1029 = ~pi001 & ~n948;
  assign n1030 = n1026 & n1028;
  assign n1031 = n977 & n1030;
  assign po054 = ~n1029 & n1031;
  assign n1033 = pi089 & n1016;
  assign n1034 = ~pi091 & n1033;
  assign n1035 = pi091 & ~n1033;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = n948 & ~n1036;
  assign n1038 = ~pi077 & ~n1037;
  assign n1039 = n948 & n1036;
  assign n1040 = ~n1038 & ~n1039;
  assign po055 = pi001 | n1040;
  assign n1042 = ~pi092 & ~n709;
  assign n1043 = ~pi000 & ~n1042;
  assign n1044 = pi092 & ~n709;
  assign po056 = n1043 | n1044;
  assign n1046 = ~pi093 & n433;
  assign n1047 = pi093 & ~n433;
  assign n1048 = ~n1046 & ~n1047;
  assign po057 = n453 & n1048;
  assign n1050 = ~n412 & po029;
  assign n1051 = ~pi006 & ~n1050;
  assign n1052 = ~pi093 & ~n1051;
  assign n1053 = pi093 & n1051;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = ~n433 & n1054;
  assign n1056 = ~pi094 & ~n1055;
  assign n1057 = pi094 & n1055;
  assign n1058 = ~n1056 & ~n1057;
  assign po058 = n453 & n1058;
  assign n1060 = pi067 & n425;
  assign n1061 = ~pi009 & n1060;
  assign n1062 = ~pi093 & ~pi094;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = pi093 & pi094;
  assign n1065 = ~n1061 & ~n1064;
  assign n1066 = ~n1051 & ~n1065;
  assign n1067 = n1063 & ~n1066;
  assign n1068 = ~n1051 & n1065;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = ~n433 & n1069;
  assign n1071 = ~pi095 & ~n1070;
  assign n1072 = pi095 & n1070;
  assign n1073 = ~n1071 & ~n1072;
  assign po059 = n453 & n1073;
  assign n1075 = pi066 & n425;
  assign n1076 = ~pi009 & n1075;
  assign n1077 = ~pi095 & ~n1063;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = pi095 & ~n1065;
  assign n1080 = ~n1076 & ~n1079;
  assign n1081 = n1051 & ~n1078;
  assign n1082 = ~n1051 & ~n1080;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n433 & ~n1083;
  assign n1085 = ~pi096 & n1084;
  assign n1086 = pi096 & ~n1084;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = n453 & ~n1087;
  assign n1089 = ~n453 & ~n1051;
  assign po060 = n1088 | n1089;
  assign n1091 = ~pi099 & ~pi100;
  assign n1092 = ~pi101 & ~pi102;
  assign n1093 = n1091 & n1092;
  assign n1094 = n453 & ~n1093;
  assign n1095 = n1051 & ~n1094;
  assign n1096 = n453 & n1093;
  assign po061 = n1095 | n1096;
  assign n1098 = pi099 & pi100;
  assign n1099 = pi101 & pi102;
  assign n1100 = n1098 & n1099;
  assign po062 = n453 & n1100;
  assign n1102 = ~pi096 & ~n1078;
  assign n1103 = ~pi009 & ~n1102;
  assign n1104 = pi096 & ~n1080;
  assign n1105 = ~pi009 & ~n1104;
  assign n1106 = ~n1051 & ~n1105;
  assign n1107 = n1103 & ~n1106;
  assign n1108 = ~n1051 & n1105;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~n433 & n1109;
  assign n1111 = ~pi099 & ~n1110;
  assign n1112 = pi099 & n1110;
  assign n1113 = ~n1111 & ~n1112;
  assign po063 = n453 & n1113;
  assign n1115 = ~pi099 & ~n1103;
  assign n1116 = pi099 & ~n1105;
  assign n1117 = ~n1051 & n1116;
  assign n1118 = ~n1115 & ~n1117;
  assign n1119 = ~n1051 & ~n1116;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~n433 & n1120;
  assign n1122 = ~pi100 & ~n1121;
  assign n1123 = pi100 & n1121;
  assign n1124 = ~n1122 & ~n1123;
  assign po064 = n453 & n1124;
  assign n1126 = ~pi100 & n1115;
  assign n1127 = n1098 & ~n1105;
  assign n1128 = ~n1051 & n1127;
  assign n1129 = ~n1126 & ~n1128;
  assign n1130 = ~n1051 & ~n1127;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = ~n433 & n1131;
  assign n1133 = ~pi101 & ~n1132;
  assign n1134 = pi101 & n1132;
  assign n1135 = ~n1133 & ~n1134;
  assign po065 = n453 & n1135;
  assign n1137 = ~pi101 & n1126;
  assign n1138 = pi100 & pi101;
  assign n1139 = pi099 & n1138;
  assign n1140 = ~n1105 & n1139;
  assign n1141 = ~n1051 & n1140;
  assign n1142 = ~n1137 & ~n1141;
  assign n1143 = ~n1051 & ~n1140;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = ~n433 & n1144;
  assign n1146 = ~pi102 & n1145;
  assign n1147 = pi102 & ~n1145;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = n453 & ~n1148;
  assign po066 = n1089 | n1149;
  assign n1151 = pi097 & ~n1103;
  assign n1152 = pi098 & ~n1105;
  assign n1153 = ~n1051 & n1152;
  assign n1154 = ~n1151 & ~n1153;
  assign n1155 = ~n1051 & ~n1152;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = ~n433 & n1156;
  assign n1158 = ~pi103 & n1157;
  assign n1159 = pi103 & ~n1157;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = n453 & ~n1160;
  assign po067 = n1089 | n1161;
  assign n1163 = ~pi103 & n1151;
  assign n1164 = ~pi009 & ~n1163;
  assign n1165 = pi103 & n1152;
  assign n1166 = ~pi009 & ~n1165;
  assign n1167 = ~n1051 & ~n1166;
  assign n1168 = n1164 & ~n1167;
  assign n1169 = ~n1051 & n1166;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n433 & n1170;
  assign n1172 = ~pi104 & n1171;
  assign n1173 = pi104 & ~n1171;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = n453 & ~n1174;
  assign po068 = n1089 | n1175;
  assign n1177 = ~pi104 & ~n1164;
  assign n1178 = pi104 & ~n1166;
  assign n1179 = ~n1051 & ~n1178;
  assign n1180 = ~n1051 & n1178;
  assign n1181 = ~n1177 & ~n1180;
  assign n1182 = ~n1179 & ~n1181;
  assign n1183 = ~n433 & n1182;
  assign n1184 = ~pi105 & ~n1183;
  assign n1185 = pi105 & n1183;
  assign n1186 = ~n1184 & ~n1185;
  assign po069 = n453 & n1186;
  assign n1188 = ~pi105 & n1177;
  assign n1189 = pi105 & n1178;
  assign n1190 = ~n1051 & n1189;
  assign n1191 = ~n1188 & ~n1190;
  assign n1192 = ~n1051 & ~n1189;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n433 & n1193;
  assign n1195 = ~pi106 & n1194;
  assign n1196 = pi106 & ~n1194;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = n453 & ~n1197;
  assign po070 = n1089 | n1198;
  assign n1200 = ~pi106 & n1188;
  assign n1201 = pi105 & pi106;
  assign n1202 = n1178 & n1201;
  assign n1203 = ~n1051 & n1202;
  assign n1204 = ~n1200 & ~n1203;
  assign n1205 = ~n1051 & ~n1202;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n433 & n1206;
  assign n1208 = ~pi107 & n1207;
  assign n1209 = pi107 & ~n1207;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = n453 & ~n1210;
  assign po071 = n1089 | n1211;
  assign n1213 = ~pi108 & n594;
  assign n1214 = pi108 & ~n594;
  assign n1215 = ~n1213 & ~n1214;
  assign po072 = n614 & n1215;
  assign n1217 = ~n576 & po133;
  assign n1218 = ~pi029 & ~n1217;
  assign n1219 = ~pi108 & ~n1218;
  assign n1220 = pi108 & n1218;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n594 & n1221;
  assign n1223 = ~pi109 & ~n1222;
  assign n1224 = pi109 & n1222;
  assign n1225 = ~n1223 & ~n1224;
  assign po073 = n614 & n1225;
  assign n1227 = pi166 & pi167;
  assign n1228 = ~pi024 & ~pi168;
  assign n1229 = n1227 & n1228;
  assign n1230 = pi171 & n1229;
  assign n1231 = ~pi032 & n1230;
  assign n1232 = ~pi108 & ~pi109;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = pi108 & pi109;
  assign n1235 = ~n1231 & ~n1234;
  assign n1236 = ~n1218 & n1235;
  assign n1237 = ~n1218 & ~n1235;
  assign n1238 = n1233 & ~n1237;
  assign n1239 = ~n1236 & ~n1238;
  assign n1240 = ~n594 & n1239;
  assign n1241 = ~pi110 & ~n1240;
  assign n1242 = pi110 & n1240;
  assign n1243 = ~n1241 & ~n1242;
  assign po074 = n614 & n1243;
  assign n1245 = pi170 & n1229;
  assign n1246 = ~pi032 & n1245;
  assign n1247 = ~pi110 & ~n1233;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = pi110 & ~n1235;
  assign n1250 = ~n1246 & ~n1249;
  assign n1251 = n1218 & ~n1248;
  assign n1252 = ~n1218 & ~n1250;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n594 & ~n1253;
  assign n1255 = ~pi111 & n1254;
  assign n1256 = pi111 & ~n1254;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = n614 & ~n1257;
  assign n1259 = ~n614 & ~n1218;
  assign po075 = n1258 | n1259;
  assign n1261 = ~pi114 & ~pi115;
  assign n1262 = ~pi116 & ~pi117;
  assign n1263 = n1261 & n1262;
  assign n1264 = n614 & n1263;
  assign n1265 = n614 & ~n1263;
  assign n1266 = n1218 & ~n1265;
  assign po076 = n1264 | n1266;
  assign n1268 = pi114 & pi115;
  assign n1269 = pi116 & pi117;
  assign n1270 = n1268 & n1269;
  assign po077 = n614 & n1270;
  assign n1272 = ~pi111 & ~n1248;
  assign n1273 = ~pi032 & ~n1272;
  assign n1274 = pi111 & ~n1250;
  assign n1275 = ~pi032 & ~n1274;
  assign n1276 = ~n1218 & n1275;
  assign n1277 = ~n1218 & ~n1275;
  assign n1278 = n1273 & ~n1277;
  assign n1279 = ~n1276 & ~n1278;
  assign n1280 = ~n594 & n1279;
  assign n1281 = ~pi114 & ~n1280;
  assign n1282 = pi114 & n1280;
  assign n1283 = ~n1281 & ~n1282;
  assign po078 = n614 & n1283;
  assign n1285 = ~pi114 & ~n1273;
  assign n1286 = pi114 & ~n1275;
  assign n1287 = ~n1218 & ~n1286;
  assign n1288 = ~n1218 & n1286;
  assign n1289 = ~n1285 & ~n1288;
  assign n1290 = ~n1287 & ~n1289;
  assign n1291 = ~n594 & n1290;
  assign n1292 = ~pi115 & ~n1291;
  assign n1293 = pi115 & n1291;
  assign n1294 = ~n1292 & ~n1293;
  assign po079 = n614 & n1294;
  assign n1296 = ~pi115 & n1285;
  assign n1297 = n1268 & ~n1275;
  assign n1298 = ~n1218 & ~n1297;
  assign n1299 = ~n1218 & n1297;
  assign n1300 = ~n1296 & ~n1299;
  assign n1301 = ~n1298 & ~n1300;
  assign n1302 = ~n594 & n1301;
  assign n1303 = ~pi116 & ~n1302;
  assign n1304 = pi116 & n1302;
  assign n1305 = ~n1303 & ~n1304;
  assign po080 = n614 & n1305;
  assign n1307 = ~pi116 & n1296;
  assign n1308 = pi115 & pi116;
  assign n1309 = pi114 & n1308;
  assign n1310 = ~n1275 & n1309;
  assign n1311 = ~n1218 & ~n1310;
  assign n1312 = ~n1218 & n1310;
  assign n1313 = ~n1307 & ~n1312;
  assign n1314 = ~n1311 & ~n1313;
  assign n1315 = ~n594 & n1314;
  assign n1316 = ~pi117 & n1315;
  assign n1317 = pi117 & ~n1315;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = n614 & ~n1318;
  assign po081 = n1259 | n1319;
  assign n1321 = pi112 & ~n1273;
  assign n1322 = pi113 & ~n1275;
  assign n1323 = ~n1218 & ~n1322;
  assign n1324 = ~n1218 & n1322;
  assign n1325 = ~n1321 & ~n1324;
  assign n1326 = ~n1323 & ~n1325;
  assign n1327 = ~n594 & n1326;
  assign n1328 = ~pi118 & n1327;
  assign n1329 = pi118 & ~n1327;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = n614 & ~n1330;
  assign po082 = n1259 | n1331;
  assign n1333 = ~pi118 & n1321;
  assign n1334 = ~pi032 & ~n1333;
  assign n1335 = pi118 & n1322;
  assign n1336 = ~pi032 & ~n1335;
  assign n1337 = ~n1218 & n1336;
  assign n1338 = ~n1218 & ~n1336;
  assign n1339 = n1334 & ~n1338;
  assign n1340 = ~n1337 & ~n1339;
  assign n1341 = ~n594 & n1340;
  assign n1342 = ~pi119 & n1341;
  assign n1343 = pi119 & ~n1341;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = n614 & ~n1344;
  assign po083 = n1259 | n1345;
  assign n1347 = ~pi119 & ~n1334;
  assign n1348 = pi119 & ~n1336;
  assign n1349 = ~n1218 & ~n1348;
  assign n1350 = ~n1218 & n1348;
  assign n1351 = ~n1347 & ~n1350;
  assign n1352 = ~n1349 & ~n1351;
  assign n1353 = ~n594 & n1352;
  assign n1354 = ~pi120 & ~n1353;
  assign n1355 = pi120 & n1353;
  assign n1356 = ~n1354 & ~n1355;
  assign po084 = n614 & n1356;
  assign n1358 = ~pi120 & n1347;
  assign n1359 = pi120 & n1348;
  assign n1360 = ~n1218 & ~n1359;
  assign n1361 = ~n1218 & n1359;
  assign n1362 = ~n1358 & ~n1361;
  assign n1363 = ~n1360 & ~n1362;
  assign n1364 = ~n594 & n1363;
  assign n1365 = ~pi121 & n1364;
  assign n1366 = pi121 & ~n1364;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = n614 & ~n1367;
  assign po085 = n1259 | n1368;
  assign n1370 = ~pi121 & n1358;
  assign n1371 = pi120 & pi121;
  assign n1372 = n1348 & n1371;
  assign n1373 = ~n1218 & ~n1372;
  assign n1374 = ~n1218 & n1372;
  assign n1375 = ~n1370 & ~n1374;
  assign n1376 = ~n1373 & ~n1375;
  assign n1377 = ~n594 & n1376;
  assign n1378 = ~pi122 & n1377;
  assign n1379 = pi122 & ~n1377;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = n614 & ~n1380;
  assign po086 = n1259 | n1381;
  assign n1383 = ~pi146 & pi147;
  assign n1384 = pi172 & n581;
  assign n1385 = pi170 & n577;
  assign n1386 = pi171 & n578;
  assign n1387 = ~n1385 & ~n1386;
  assign n1388 = ~n1384 & n1387;
  assign n1389 = n1383 & ~n1388;
  assign n1390 = po133 & n1389;
  assign n1391 = ~pi030 & ~n1390;
  assign n1392 = ~pi123 & ~n1391;
  assign n1393 = pi123 & n1391;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = pi146 & n583;
  assign n1396 = pi166 & ~pi167;
  assign n1397 = ~pi168 & n1396;
  assign n1398 = ~pi024 & n1397;
  assign n1399 = po133 & n1395;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = n1394 & n1400;
  assign n1402 = ~n1394 & n1400;
  assign n1403 = ~pi114 & ~n1402;
  assign n1404 = ~n1401 & ~n1403;
  assign po087 = ~pi024 & n1404;
  assign n1406 = ~pi031 & n576;
  assign n1407 = ~pi123 & ~n1406;
  assign n1408 = pi123 & n1406;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = ~n1391 & n1409;
  assign n1411 = ~pi124 & n1410;
  assign n1412 = pi124 & ~n1410;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = n1400 & n1413;
  assign n1415 = n1400 & ~n1413;
  assign n1416 = ~pi115 & ~n1415;
  assign n1417 = ~n1414 & ~n1416;
  assign po088 = ~pi024 & n1417;
  assign n1419 = ~pi123 & ~pi124;
  assign n1420 = pi123 & pi124;
  assign n1421 = ~n1406 & ~n1420;
  assign n1422 = ~n1406 & n1420;
  assign n1423 = ~n1419 & ~n1422;
  assign n1424 = ~n1421 & ~n1423;
  assign n1425 = ~n1391 & n1424;
  assign n1426 = ~pi125 & n1425;
  assign n1427 = pi125 & ~n1425;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = n1400 & n1428;
  assign n1430 = n1400 & ~n1428;
  assign n1431 = ~pi116 & ~n1430;
  assign n1432 = ~n1429 & ~n1431;
  assign po089 = ~pi024 & n1432;
  assign n1434 = ~pi125 & n1419;
  assign n1435 = ~pi033 & ~n1434;
  assign n1436 = pi125 & n1420;
  assign n1437 = ~pi033 & ~n1436;
  assign n1438 = ~n1406 & n1437;
  assign n1439 = ~n1406 & ~n1437;
  assign n1440 = n1435 & ~n1439;
  assign n1441 = ~n1438 & ~n1440;
  assign n1442 = ~n1391 & n1441;
  assign n1443 = ~pi126 & n1442;
  assign n1444 = pi126 & ~n1442;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = n1400 & n1445;
  assign n1447 = n1400 & ~n1445;
  assign n1448 = ~pi117 & ~n1447;
  assign n1449 = ~n1446 & ~n1448;
  assign po090 = pi024 | n1449;
  assign n1451 = ~pi126 & ~n1435;
  assign n1452 = pi126 & ~n1437;
  assign n1453 = ~n1406 & ~n1452;
  assign n1454 = ~n1406 & n1452;
  assign n1455 = ~n1451 & ~n1454;
  assign n1456 = ~n1453 & ~n1455;
  assign n1457 = ~n1391 & n1456;
  assign n1458 = ~pi127 & n1457;
  assign n1459 = pi127 & ~n1457;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = n1400 & n1460;
  assign n1462 = n1400 & ~n1460;
  assign n1463 = ~pi118 & ~n1462;
  assign n1464 = ~n1461 & ~n1463;
  assign po091 = pi024 | n1464;
  assign n1466 = ~pi127 & n1451;
  assign n1467 = pi126 & pi127;
  assign n1468 = ~n1437 & n1467;
  assign n1469 = ~n1406 & ~n1468;
  assign n1470 = ~n1406 & n1468;
  assign n1471 = ~n1466 & ~n1470;
  assign n1472 = ~n1469 & ~n1471;
  assign n1473 = ~n1391 & n1472;
  assign n1474 = ~pi128 & n1473;
  assign n1475 = pi128 & ~n1473;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = n1400 & n1476;
  assign n1478 = n1400 & ~n1476;
  assign n1479 = ~pi119 & ~n1478;
  assign n1480 = ~n1477 & ~n1479;
  assign po092 = pi024 | n1480;
  assign n1482 = ~pi127 & ~pi128;
  assign n1483 = n1451 & n1482;
  assign n1484 = ~pi033 & ~n1483;
  assign n1485 = pi127 & pi128;
  assign n1486 = n1452 & n1485;
  assign n1487 = ~pi033 & ~n1486;
  assign n1488 = ~n1406 & n1487;
  assign n1489 = ~n1406 & ~n1487;
  assign n1490 = n1484 & ~n1489;
  assign n1491 = ~n1488 & ~n1490;
  assign n1492 = ~n1391 & n1491;
  assign n1493 = ~pi129 & n1492;
  assign n1494 = pi129 & ~n1492;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = n1400 & n1495;
  assign n1497 = n1400 & ~n1495;
  assign n1498 = ~pi120 & ~n1497;
  assign n1499 = ~n1496 & ~n1498;
  assign po093 = ~pi024 & n1499;
  assign n1501 = ~pi129 & ~n1484;
  assign n1502 = pi129 & ~n1487;
  assign n1503 = ~n1406 & ~n1502;
  assign n1504 = ~n1406 & n1502;
  assign n1505 = ~n1501 & ~n1504;
  assign n1506 = ~n1503 & ~n1505;
  assign n1507 = ~n1391 & n1506;
  assign n1508 = ~pi130 & n1507;
  assign n1509 = pi130 & ~n1507;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = n1400 & n1510;
  assign n1512 = n1400 & ~n1510;
  assign n1513 = ~pi121 & ~n1512;
  assign n1514 = ~n1511 & ~n1513;
  assign po094 = pi024 | n1514;
  assign n1516 = ~pi130 & n1501;
  assign n1517 = pi129 & pi130;
  assign n1518 = ~n1487 & n1517;
  assign n1519 = ~n1406 & ~n1518;
  assign n1520 = ~n1406 & n1518;
  assign n1521 = ~n1516 & ~n1520;
  assign n1522 = ~n1519 & ~n1521;
  assign n1523 = ~n1391 & n1522;
  assign n1524 = ~pi131 & n1523;
  assign n1525 = pi131 & ~n1523;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = n1400 & n1526;
  assign n1528 = n1400 & ~n1526;
  assign n1529 = ~pi122 & ~n1528;
  assign n1530 = ~n1527 & ~n1529;
  assign po095 = pi024 | n1530;
  assign po096 = pi024 | ~pi132;
  assign n1533 = ~pi132 & ~pi133;
  assign n1534 = ~n601 & ~n1533;
  assign po097 = pi024 | n1534;
  assign n1536 = ~pi134 & ~n601;
  assign n1537 = ~n602 & ~n1536;
  assign po098 = pi024 | n1537;
  assign n1539 = ~pi135 & ~n606;
  assign n1540 = pi135 & n606;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~pi167 & pi168;
  assign n1543 = ~pi024 & pi166;
  assign n1544 = n1542 & n1543;
  assign n1545 = ~n608 & ~n1544;
  assign n1546 = n1541 & n1545;
  assign n1547 = ~n1541 & n1545;
  assign n1548 = ~pi123 & ~n1547;
  assign n1549 = ~n1546 & ~n1548;
  assign po099 = pi024 | n1549;
  assign n1551 = ~pi136 & n607;
  assign n1552 = pi136 & ~n607;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = n1545 & n1553;
  assign n1555 = n1545 & ~n1553;
  assign n1556 = ~pi124 & ~n1555;
  assign n1557 = ~n1554 & ~n1556;
  assign po100 = pi024 | n1557;
  assign n1559 = ~pi137 & n603;
  assign n1560 = ~n604 & ~n1559;
  assign po101 = pi024 | n1560;
  assign n1562 = pi136 & n607;
  assign n1563 = ~pi138 & n1562;
  assign n1564 = pi138 & ~n1562;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = n1545 & n1565;
  assign n1567 = n1545 & ~n1565;
  assign n1568 = ~pi125 & ~n1567;
  assign n1569 = ~n1566 & ~n1568;
  assign po102 = pi024 | n1569;
  assign n1571 = pi136 & pi138;
  assign n1572 = n607 & n1571;
  assign n1573 = ~pi139 & n1572;
  assign n1574 = pi139 & ~n1572;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = n1545 & n1575;
  assign n1577 = n1545 & ~n1575;
  assign n1578 = ~pi126 & ~n1577;
  assign n1579 = ~n1576 & ~n1578;
  assign po103 = pi024 | n1579;
  assign n1581 = pi139 & n1572;
  assign n1582 = ~pi140 & n1581;
  assign n1583 = pi140 & ~n1581;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n1545 & n1584;
  assign n1586 = n1545 & ~n1584;
  assign n1587 = ~pi127 & ~n1586;
  assign n1588 = ~n1585 & ~n1587;
  assign po104 = pi024 | n1588;
  assign n1590 = pi140 & n1581;
  assign n1591 = ~pi034 & ~n1590;
  assign n1592 = ~pi141 & ~n1591;
  assign n1593 = pi141 & n1591;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = n1545 & n1594;
  assign n1596 = n1545 & ~n1594;
  assign n1597 = ~pi128 & ~n1596;
  assign n1598 = ~n1595 & ~n1597;
  assign po105 = pi024 | n1598;
  assign n1600 = pi141 & ~n1591;
  assign n1601 = ~pi142 & n1600;
  assign n1602 = pi142 & ~n1600;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = n1545 & n1603;
  assign n1605 = n1545 & ~n1603;
  assign n1606 = ~pi129 & ~n1605;
  assign n1607 = ~n1604 & ~n1606;
  assign po106 = pi024 | n1607;
  assign n1609 = pi141 & pi142;
  assign n1610 = ~n1591 & n1609;
  assign n1611 = ~pi143 & n1610;
  assign n1612 = pi143 & ~n1610;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = n1545 & n1613;
  assign n1615 = n1545 & ~n1613;
  assign n1616 = ~pi130 & ~n1615;
  assign n1617 = ~n1614 & ~n1616;
  assign po107 = pi024 | n1617;
  assign n1619 = pi143 & pi145;
  assign n1620 = pi142 & n1619;
  assign n1621 = pi140 & pi141;
  assign n1622 = pi139 & n1621;
  assign n1623 = ~pi024 & ~n1545;
  assign n1624 = n1620 & n1622;
  assign n1625 = n1571 & n1624;
  assign po108 = ~n1623 & n1625;
  assign n1627 = pi143 & n1610;
  assign n1628 = ~pi145 & n1627;
  assign n1629 = pi145 & ~n1627;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n1545 & n1630;
  assign n1632 = n1545 & ~n1630;
  assign n1633 = ~pi131 & ~n1632;
  assign n1634 = ~n1631 & ~n1633;
  assign po109 = pi024 | n1634;
  assign n1636 = pi172 & n1229;
  assign n1637 = n576 & ~n1636;
  assign n1638 = n572 & n1637;
  assign n1639 = ~pi146 & n1638;
  assign n1640 = pi146 & ~n1638;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = n585 & po133;
  assign n1643 = pi146 & n1636;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = ~pi024 & ~n1544;
  assign n1646 = n1644 & n1645;
  assign po110 = n1641 & n1646;
  assign n1648 = ~pi147 & ~n1640;
  assign n1649 = pi147 & n1640;
  assign n1650 = ~n1648 & ~n1649;
  assign po111 = n1646 & n1650;
  assign n1652 = pi146 & pi147;
  assign n1653 = ~n1638 & n1652;
  assign n1654 = ~pi148 & ~n1653;
  assign n1655 = pi148 & n1653;
  assign n1656 = ~n1654 & ~n1655;
  assign po112 = n1646 & n1656;
  assign n1658 = pi148 & n1652;
  assign n1659 = ~n1638 & n1658;
  assign n1660 = ~pi149 & ~n1659;
  assign n1661 = pi149 & n1659;
  assign n1662 = ~n1660 & ~n1661;
  assign po113 = n1646 & n1662;
  assign n1664 = pi148 & pi149;
  assign n1665 = n1652 & n1664;
  assign n1666 = ~n1638 & n1665;
  assign n1667 = ~pi150 & ~n1666;
  assign n1668 = pi150 & n1666;
  assign n1669 = ~n1667 & ~n1668;
  assign po114 = n1646 & n1669;
  assign n1671 = pi150 & n1665;
  assign n1672 = ~n1638 & n1671;
  assign n1673 = ~pi151 & ~n1672;
  assign n1674 = pi151 & n1672;
  assign n1675 = ~n1673 & ~n1674;
  assign po115 = n1646 & n1675;
  assign n1677 = pi151 & n1671;
  assign n1678 = ~n1638 & n1677;
  assign n1679 = ~pi152 & ~n1678;
  assign n1680 = pi152 & n1678;
  assign n1681 = ~n1679 & ~n1680;
  assign po116 = n1646 & n1681;
  assign n1683 = pi150 & pi151;
  assign n1684 = pi152 & n1683;
  assign n1685 = n1665 & n1684;
  assign n1686 = ~n1638 & n1685;
  assign n1687 = ~pi153 & ~n1686;
  assign n1688 = pi153 & n1686;
  assign n1689 = ~n1687 & ~n1688;
  assign po117 = n1646 & n1689;
  assign n1691 = pi153 & ~n1638;
  assign n1692 = n1685 & n1691;
  assign n1693 = pi154 & n1692;
  assign n1694 = ~pi154 & ~n1692;
  assign n1695 = ~n1693 & ~n1694;
  assign po118 = n1646 & n1695;
  assign n1697 = pi158 & n562;
  assign n1698 = n1645 & ~n1697;
  assign n1699 = pi158 & n1698;
  assign po122 = n571 | n1699;
  assign n1701 = pi159 & n566;
  assign n1702 = n1645 & ~n1701;
  assign n1703 = pi159 & n1702;
  assign po123 = n574 | n1703;
  assign n1705 = pi162 & n608;
  assign n1706 = ~pi162 & ~n608;
  assign n1707 = ~n1705 & ~n1706;
  assign n1708 = ~pi024 & n1707;
  assign n1709 = ~n1398 & ~n1544;
  assign po126 = n1708 | ~n1709;
  assign n1711 = ~pi162 & po126;
  assign n1712 = ~pi160 & ~pi161;
  assign n1713 = n1711 & ~n1712;
  assign n1714 = n1711 & n1712;
  assign n1715 = ~pi160 & ~n1714;
  assign n1716 = ~n1713 & ~n1715;
  assign n1717 = ~pi024 & ~n1716;
  assign po124 = n1709 & ~n1717;
  assign n1719 = ~pi161 & ~n1711;
  assign n1720 = pi161 & ~n1711;
  assign n1721 = ~pi160 & ~n1720;
  assign n1722 = ~n1719 & ~n1721;
  assign n1723 = n1709 & ~n1722;
  assign po125 = ~pi024 & ~n1723;
  assign n1725 = pi164 & n1229;
  assign n1726 = ~pi164 & ~n1229;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~pi024 & ~n560;
  assign po128 = n1727 & n1728;
  assign n1730 = ~pi165 & ~n1725;
  assign n1731 = pi165 & n1725;
  assign n1732 = ~n1730 & ~n1731;
  assign po129 = n1728 & n1732;
  assign n1734 = n562 & ~n631;
  assign n1735 = n623 & n1734;
  assign n1736 = n1229 & ~n1735;
  assign n1737 = n562 & n613;
  assign n1738 = ~n1398 & ~n1736;
  assign n1739 = ~n1737 & n1738;
  assign po130 = ~pi024 & ~n1739;
  assign n1741 = pi172 & ~n1693;
  assign n1742 = pi172 & n1693;
  assign n1743 = ~pi154 & ~n1742;
  assign n1744 = ~n1741 & ~n1743;
  assign n1745 = ~pi025 & ~n1744;
  assign n1746 = po133 & ~n1745;
  assign n1747 = n631 & n1229;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = pi168 & n587;
  assign n1750 = ~pi024 & n1749;
  assign n1751 = ~n613 & n1748;
  assign n1752 = ~n1750 & n1751;
  assign n1753 = pi168 & n1227;
  assign n1754 = ~pi024 & n1753;
  assign n1755 = pi167 & pi168;
  assign n1756 = ~n562 & ~n631;
  assign n1757 = n1229 & n1756;
  assign n1758 = ~n1755 & ~n1757;
  assign n1759 = ~n1754 & n1758;
  assign n1760 = n1752 & n1759;
  assign po131 = ~pi024 & ~n1760;
  assign n1762 = ~n1747 & ~n1750;
  assign n1763 = ~n1398 & n1762;
  assign n1764 = n562 & n1229;
  assign n1765 = n623 & ~n631;
  assign n1766 = n1764 & n1765;
  assign n1767 = ~n1754 & ~n1766;
  assign n1768 = n1763 & n1767;
  assign po132 = ~pi024 & ~n1768;
  assign n1770 = pi171 & pi172;
  assign n1771 = ~pi170 & ~n1770;
  assign n1772 = ~pi171 & ~pi172;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = ~pi170 & n1772;
  assign n1775 = ~pi024 & ~n1774;
  assign n1776 = ~n1773 & n1775;
  assign n1777 = ~pi027 & ~n1754;
  assign n1778 = ~pi026 & ~n1750;
  assign n1779 = pi171 & ~n1778;
  assign n1780 = pi172 & ~n1777;
  assign n1781 = ~pi170 & ~n1780;
  assign n1782 = ~pi172 & ~n1777;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1779 & ~n1783;
  assign n1785 = ~n1778 & ~n1780;
  assign n1786 = ~pi171 & n1785;
  assign n1787 = ~n1784 & ~n1786;
  assign po134 = ~n1776 | n1787;
  assign n1789 = pi172 & ~n1778;
  assign n1790 = pi171 & n1777;
  assign n1791 = ~pi170 & ~n1790;
  assign n1792 = ~pi171 & n1777;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = ~n1789 & ~n1793;
  assign n1795 = pi170 & ~n1777;
  assign n1796 = ~n1778 & ~n1795;
  assign n1797 = ~pi172 & n1796;
  assign n1798 = ~n1794 & ~n1797;
  assign po135 = n1776 & n1798;
  assign n1800 = pi170 & ~n1778;
  assign n1801 = ~pi172 & n1777;
  assign n1802 = pi172 & n1777;
  assign n1803 = ~pi171 & ~n1802;
  assign n1804 = ~n1801 & ~n1803;
  assign n1805 = ~n1800 & ~n1804;
  assign n1806 = pi171 & ~n1777;
  assign n1807 = ~n1778 & ~n1806;
  assign n1808 = ~pi170 & n1807;
  assign n1809 = ~n1805 & ~n1808;
  assign po136 = n1776 & n1809;
  assign po019 = pi000;
  assign po020 = pi055;
  assign po025 = pi060;
  assign po119 = pi023;
  assign po120 = pi155;
  assign po127 = pi161;
endmodule



// Benchmark "DES" written by ABC on Sun Apr 22 21:43:02 2018

module DES ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244;
  wire n502, n503, n504, n505, n506, n507, n509, n510, n511, n513, n514,
    n515, n517, n518, n519, n521, n522, n523, n525, n526, n527, n529, n530,
    n531, n533, n534, n535, n537, n538, n539, n541, n542, n543, n545, n546,
    n547, n549, n550, n551, n553, n554, n555, n557, n558, n559, n561, n562,
    n563, n565, n566, n567, n569, n570, n571, n573, n574, n575, n577, n578,
    n579, n581, n582, n583, n585, n586, n587, n589, n590, n591, n593, n594,
    n595, n597, n598, n599, n601, n602, n603, n605, n606, n607, n609, n610,
    n611, n613, n614, n615, n617, n618, n619, n621, n622, n623, n625, n626,
    n627, n629, n630, n631, n633, n634, n635, n637, n638, n639, n641, n642,
    n643, n645, n646, n647, n649, n650, n651, n653, n654, n655, n657, n658,
    n659, n661, n662, n663, n665, n666, n667, n669, n670, n671, n673, n674,
    n675, n677, n678, n679, n681, n682, n683, n685, n686, n687, n689, n690,
    n691, n693, n694, n695, n697, n698, n699, n701, n702, n703, n705, n706,
    n707, n709, n710, n711, n713, n714, n715, n717, n718, n719, n721, n722,
    n723, n725, n726, n727, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n872, n873, n874, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1022,
    n1023, n1024, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1088, n1089, n1090, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1235, n1236,
    n1237, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1309, n1310, n1311, n1312, n1313, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1466, n1467, n1468, n1469, n1470,
    n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1524, n1525, n1526, n1527, n1528, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1600, n1601, n1602, n1603, n1604,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1758, n1759, n1760, n1761, n1762, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1917, n1918,
    n1919, n1920, n1921, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1983, n1984, n1985, n1986, n1987, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2061, n2062,
    n2063, n2064, n2065, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2118, n2119, n2120, n2121, n2122, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2168, n2169, n2170, n2171, n2172, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2318,
    n2319, n2320, n2321, n2322, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2379, n2380,
    n2381, n2382, n2383, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
    n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2432,
    n2433, n2434, n2435, n2436, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2505, n2506, n2507, n2508, n2509, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2559, n2560, n2561, n2562, n2563, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613, n2615, n2616, n2617, n2618,
    n2619, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2768, n2769, n2770,
    n2771, n2772, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2845, n2846, n2847, n2848, n2849, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2911, n2912, n2913, n2914,
    n2915, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2987, n2988, n2989, n2990, n2991, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3044, n3045, n3046, n3047, n3048,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3096, n3097, n3098, n3099, n3100,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
    n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3154, n3155, n3156, n3157, n3158, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3214,
    n3215, n3216, n3217, n3218, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
    n3267, n3268, n3269, n3270, n3271, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3326, n3327, n3328,
    n3329, n3330, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3380,
    n3381, n3382, n3383, n3384, n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
    n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3432, n3434, n3435, n3436, n3437, n3438, n3440, n3441, n3443, n3444,
    n3446, n3447, n3449, n3450, n3452, n3453, n3455, n3456, n3458, n3459,
    n3461, n3462, n3464, n3465, n3467, n3468, n3470, n3471, n3473, n3474,
    n3476, n3477, n3479, n3480, n3482, n3483, n3485, n3486, n3488, n3489,
    n3491, n3492, n3494, n3495, n3497, n3498, n3500, n3501, n3503, n3504,
    n3506, n3507, n3509, n3510, n3512, n3513, n3515, n3516, n3518, n3519,
    n3521, n3522, n3524, n3525, n3527, n3528, n3530, n3531, n3533, n3534,
    n3536, n3537, n3539, n3540, n3542, n3543, n3545, n3546, n3548, n3549,
    n3551, n3552, n3554, n3555, n3557, n3558, n3560, n3561, n3563, n3564,
    n3566, n3567, n3569, n3570, n3572, n3573, n3575, n3576, n3578, n3579,
    n3581, n3582, n3584, n3585, n3587, n3588, n3590, n3591, n3593, n3594,
    n3596, n3597, n3599, n3600, n3602, n3603, n3605, n3606, n3608, n3609,
    n3611, n3612, n3614, n3615, n3617, n3618, n3620, n3621, n3623, n3624,
    n3626, n3627, n3629, n3630, n3632, n3633, n3634, n3635, n3636, n3637,
    n3639, n3640, n3641, n3642, n3644, n3645, n3646, n3647, n3649, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
    n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
    n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3859, n3860, n3861, n3862,
    n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
    n3905, n3906, n3907, n3908, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942, n3944, n3945, n3946, n3947,
    n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
    n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
    n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
    n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4505, n4506, n4507, n4508, n4509, n4510,
    n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
    n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
    n4553, n4554, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4603, n4604, n4605, n4606,
    n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
    n4618, n4619, n4620, n4621, n4622, n4623;
  assign n502 = pi197 & pi198;
  assign n503 = pi196 & n502;
  assign n504 = pi195 & n503;
  assign n505 = pi019 & pi198;
  assign n506 = pi011 & ~pi198;
  assign n507 = ~n505 & ~n506;
  assign po000 = ~n504 & ~n507;
  assign n509 = pi020 & pi198;
  assign n510 = pi012 & ~pi198;
  assign n511 = ~n509 & ~n510;
  assign po001 = ~n504 & ~n511;
  assign n513 = pi021 & pi198;
  assign n514 = pi013 & ~pi198;
  assign n515 = ~n513 & ~n514;
  assign po002 = ~n504 & ~n515;
  assign n517 = pi022 & pi198;
  assign n518 = pi014 & ~pi198;
  assign n519 = ~n517 & ~n518;
  assign po003 = ~n504 & ~n519;
  assign n521 = pi023 & pi198;
  assign n522 = pi015 & ~pi198;
  assign n523 = ~n521 & ~n522;
  assign po004 = ~n504 & ~n523;
  assign n525 = pi024 & pi198;
  assign n526 = pi016 & ~pi198;
  assign n527 = ~n525 & ~n526;
  assign po005 = ~n504 & ~n527;
  assign n529 = pi025 & pi198;
  assign n530 = pi017 & ~pi198;
  assign n531 = ~n529 & ~n530;
  assign po006 = ~n504 & ~n531;
  assign n533 = pi026 & pi198;
  assign n534 = pi018 & ~pi198;
  assign n535 = ~n533 & ~n534;
  assign po007 = ~n504 & ~n535;
  assign n537 = pi027 & pi198;
  assign n538 = pi019 & ~pi198;
  assign n539 = ~n537 & ~n538;
  assign po008 = ~n504 & ~n539;
  assign n541 = pi028 & pi198;
  assign n542 = pi020 & ~pi198;
  assign n543 = ~n541 & ~n542;
  assign po009 = ~n504 & ~n543;
  assign n545 = pi029 & pi198;
  assign n546 = pi021 & ~pi198;
  assign n547 = ~n545 & ~n546;
  assign po010 = ~n504 & ~n547;
  assign n549 = pi030 & pi198;
  assign n550 = pi022 & ~pi198;
  assign n551 = ~n549 & ~n550;
  assign po011 = ~n504 & ~n551;
  assign n553 = pi031 & pi198;
  assign n554 = pi023 & ~pi198;
  assign n555 = ~n553 & ~n554;
  assign po012 = ~n504 & ~n555;
  assign n557 = pi032 & pi198;
  assign n558 = pi024 & ~pi198;
  assign n559 = ~n557 & ~n558;
  assign po013 = ~n504 & ~n559;
  assign n561 = pi033 & pi198;
  assign n562 = pi025 & ~pi198;
  assign n563 = ~n561 & ~n562;
  assign po014 = ~n504 & ~n563;
  assign n565 = pi034 & pi198;
  assign n566 = pi026 & ~pi198;
  assign n567 = ~n565 & ~n566;
  assign po015 = ~n504 & ~n567;
  assign n569 = pi035 & pi198;
  assign n570 = pi027 & ~pi198;
  assign n571 = ~n569 & ~n570;
  assign po016 = ~n504 & ~n571;
  assign n573 = pi036 & pi198;
  assign n574 = pi028 & ~pi198;
  assign n575 = ~n573 & ~n574;
  assign po017 = ~n504 & ~n575;
  assign n577 = pi037 & pi198;
  assign n578 = pi029 & ~pi198;
  assign n579 = ~n577 & ~n578;
  assign po018 = ~n504 & ~n579;
  assign n581 = pi038 & pi198;
  assign n582 = pi030 & ~pi198;
  assign n583 = ~n581 & ~n582;
  assign po019 = ~n504 & ~n583;
  assign n585 = pi039 & pi198;
  assign n586 = pi031 & ~pi198;
  assign n587 = ~n585 & ~n586;
  assign po020 = ~n504 & ~n587;
  assign n589 = pi040 & pi198;
  assign n590 = pi032 & ~pi198;
  assign n591 = ~n589 & ~n590;
  assign po021 = ~n504 & ~n591;
  assign n593 = pi041 & pi198;
  assign n594 = pi033 & ~pi198;
  assign n595 = ~n593 & ~n594;
  assign po022 = ~n504 & ~n595;
  assign n597 = pi042 & pi198;
  assign n598 = pi034 & ~pi198;
  assign n599 = ~n597 & ~n598;
  assign po023 = ~n504 & ~n599;
  assign n601 = pi043 & pi198;
  assign n602 = pi035 & ~pi198;
  assign n603 = ~n601 & ~n602;
  assign po024 = ~n504 & ~n603;
  assign n605 = pi044 & pi198;
  assign n606 = pi036 & ~pi198;
  assign n607 = ~n605 & ~n606;
  assign po025 = ~n504 & ~n607;
  assign n609 = pi045 & pi198;
  assign n610 = pi037 & ~pi198;
  assign n611 = ~n609 & ~n610;
  assign po026 = ~n504 & ~n611;
  assign n613 = pi046 & pi198;
  assign n614 = pi038 & ~pi198;
  assign n615 = ~n613 & ~n614;
  assign po027 = ~n504 & ~n615;
  assign n617 = pi047 & pi198;
  assign n618 = pi039 & ~pi198;
  assign n619 = ~n617 & ~n618;
  assign po028 = ~n504 & ~n619;
  assign n621 = pi048 & pi198;
  assign n622 = pi040 & ~pi198;
  assign n623 = ~n621 & ~n622;
  assign po029 = ~n504 & ~n623;
  assign n625 = pi049 & pi198;
  assign n626 = pi041 & ~pi198;
  assign n627 = ~n625 & ~n626;
  assign po030 = ~n504 & ~n627;
  assign n629 = pi050 & pi198;
  assign n630 = pi042 & ~pi198;
  assign n631 = ~n629 & ~n630;
  assign po031 = ~n504 & ~n631;
  assign n633 = pi051 & pi198;
  assign n634 = pi043 & ~pi198;
  assign n635 = ~n633 & ~n634;
  assign po032 = ~n504 & ~n635;
  assign n637 = pi052 & pi198;
  assign n638 = pi044 & ~pi198;
  assign n639 = ~n637 & ~n638;
  assign po033 = ~n504 & ~n639;
  assign n641 = pi053 & pi198;
  assign n642 = pi045 & ~pi198;
  assign n643 = ~n641 & ~n642;
  assign po034 = ~n504 & ~n643;
  assign n645 = pi054 & pi198;
  assign n646 = pi046 & ~pi198;
  assign n647 = ~n645 & ~n646;
  assign po035 = ~n504 & ~n647;
  assign n649 = pi055 & pi198;
  assign n650 = pi047 & ~pi198;
  assign n651 = ~n649 & ~n650;
  assign po036 = ~n504 & ~n651;
  assign n653 = pi056 & pi198;
  assign n654 = pi048 & ~pi198;
  assign n655 = ~n653 & ~n654;
  assign po037 = ~n504 & ~n655;
  assign n657 = pi049 & ~pi198;
  assign n658 = pi057 & pi198;
  assign n659 = ~n657 & ~n658;
  assign po038 = ~n504 & ~n659;
  assign n661 = pi050 & ~pi198;
  assign n662 = pi058 & pi198;
  assign n663 = ~n661 & ~n662;
  assign po039 = ~n504 & ~n663;
  assign n665 = pi051 & ~pi198;
  assign n666 = pi059 & pi198;
  assign n667 = ~n665 & ~n666;
  assign po040 = ~n504 & ~n667;
  assign n669 = pi052 & ~pi198;
  assign n670 = pi060 & pi198;
  assign n671 = ~n669 & ~n670;
  assign po041 = ~n504 & ~n671;
  assign n673 = pi053 & ~pi198;
  assign n674 = pi061 & pi198;
  assign n675 = ~n673 & ~n674;
  assign po042 = ~n504 & ~n675;
  assign n677 = pi054 & ~pi198;
  assign n678 = pi062 & pi198;
  assign n679 = ~n677 & ~n678;
  assign po043 = ~n504 & ~n679;
  assign n681 = pi055 & ~pi198;
  assign n682 = pi063 & pi198;
  assign n683 = ~n681 & ~n682;
  assign po044 = ~n504 & ~n683;
  assign n685 = pi056 & ~pi198;
  assign n686 = pi064 & pi198;
  assign n687 = ~n685 & ~n686;
  assign po045 = ~n504 & ~n687;
  assign n689 = pi065 & pi198;
  assign n690 = pi057 & ~pi198;
  assign n691 = ~n689 & ~n690;
  assign po046 = ~n504 & ~n691;
  assign n693 = pi066 & pi198;
  assign n694 = pi058 & ~pi198;
  assign n695 = ~n693 & ~n694;
  assign po047 = ~n504 & ~n695;
  assign n697 = pi000 & pi198;
  assign n698 = pi059 & ~pi198;
  assign n699 = ~n697 & ~n698;
  assign po048 = ~n504 & ~n699;
  assign n701 = pi001 & pi198;
  assign n702 = pi060 & ~pi198;
  assign n703 = ~n701 & ~n702;
  assign po049 = ~n504 & ~n703;
  assign n705 = pi002 & pi198;
  assign n706 = pi061 & ~pi198;
  assign n707 = ~n705 & ~n706;
  assign po050 = ~n504 & ~n707;
  assign n709 = pi003 & pi198;
  assign n710 = pi062 & ~pi198;
  assign n711 = ~n709 & ~n710;
  assign po051 = ~n504 & ~n711;
  assign n713 = pi004 & pi198;
  assign n714 = pi063 & ~pi198;
  assign n715 = ~n713 & ~n714;
  assign po052 = ~n504 & ~n715;
  assign n717 = pi005 & pi198;
  assign n718 = pi064 & ~pi198;
  assign n719 = ~n717 & ~n718;
  assign po053 = ~n504 & ~n719;
  assign n721 = pi006 & pi198;
  assign n722 = pi065 & ~pi198;
  assign n723 = ~n721 & ~n722;
  assign po054 = ~n504 & ~n723;
  assign n725 = pi007 & pi198;
  assign n726 = pi066 & ~pi198;
  assign n727 = ~n725 & ~n726;
  assign po055 = ~n504 & ~n727;
  assign n729 = pi147 & ~pi242;
  assign n730 = ~pi147 & pi242;
  assign n731 = ~n729 & ~n730;
  assign n732 = pi146 & ~pi231;
  assign n733 = ~pi146 & pi231;
  assign n734 = ~n732 & ~n733;
  assign n735 = pi145 & ~pi252;
  assign n736 = ~pi145 & pi252;
  assign n737 = ~n735 & ~n736;
  assign n738 = pi144 & ~pi246;
  assign n739 = ~pi144 & pi246;
  assign n740 = ~n738 & ~n739;
  assign n741 = pi143 & ~pi236;
  assign n742 = ~pi143 & pi236;
  assign n743 = ~n741 & ~n742;
  assign n744 = pi142 & ~pi228;
  assign n745 = ~pi142 & pi228;
  assign n746 = ~n744 & ~n745;
  assign n747 = n731 & n734;
  assign n748 = ~n737 & n747;
  assign n749 = n740 & n748;
  assign n750 = n743 & n749;
  assign n751 = n746 & n750;
  assign n752 = ~n743 & n749;
  assign n753 = n746 & n752;
  assign n754 = ~n740 & n748;
  assign n755 = n743 & n754;
  assign n756 = n746 & n755;
  assign n757 = ~n743 & n754;
  assign n758 = n746 & n757;
  assign n759 = n731 & ~n734;
  assign n760 = n737 & n759;
  assign n761 = ~n740 & n760;
  assign n762 = n743 & n761;
  assign n763 = n746 & n762;
  assign n764 = ~n743 & n761;
  assign n765 = n746 & n764;
  assign n766 = ~n737 & n759;
  assign n767 = ~n740 & n766;
  assign n768 = n743 & n767;
  assign n769 = n746 & n768;
  assign n770 = n737 & n747;
  assign n771 = n740 & n770;
  assign n772 = n743 & n771;
  assign n773 = ~n746 & n772;
  assign n774 = ~n743 & n771;
  assign n775 = ~n746 & n774;
  assign n776 = ~n746 & n752;
  assign n777 = ~n746 & n762;
  assign n778 = ~n746 & n764;
  assign n779 = n740 & n766;
  assign n780 = n743 & n779;
  assign n781 = ~n746 & n780;
  assign n782 = ~n743 & n767;
  assign n783 = ~n746 & n782;
  assign n784 = ~n731 & n734;
  assign n785 = n737 & n784;
  assign n786 = ~n740 & n785;
  assign n787 = ~n743 & n786;
  assign n788 = n746 & n787;
  assign n789 = ~n737 & n784;
  assign n790 = n740 & n789;
  assign n791 = n743 & n790;
  assign n792 = n746 & n791;
  assign n793 = ~n740 & n789;
  assign n794 = n743 & n793;
  assign n795 = n746 & n794;
  assign n796 = ~n731 & ~n734;
  assign n797 = n737 & n796;
  assign n798 = n740 & n797;
  assign n799 = n743 & n798;
  assign n800 = n746 & n799;
  assign n801 = ~n737 & n796;
  assign n802 = n740 & n801;
  assign n803 = n743 & n802;
  assign n804 = n746 & n803;
  assign n805 = ~n743 & n802;
  assign n806 = n746 & n805;
  assign n807 = ~n740 & n801;
  assign n808 = ~n743 & n807;
  assign n809 = n746 & n808;
  assign n810 = n740 & n785;
  assign n811 = n743 & n810;
  assign n812 = ~n746 & n811;
  assign n813 = ~n746 & n787;
  assign n814 = ~n743 & n790;
  assign n815 = ~n746 & n814;
  assign n816 = ~n746 & n799;
  assign n817 = ~n743 & n798;
  assign n818 = ~n746 & n817;
  assign n819 = ~n746 & n803;
  assign n820 = ~n746 & n808;
  assign n821 = ~n753 & ~n756;
  assign n822 = ~n751 & n821;
  assign n823 = ~n758 & ~n763;
  assign n824 = ~n765 & ~n769;
  assign n825 = n823 & n824;
  assign n826 = n822 & n825;
  assign n827 = ~n775 & ~n776;
  assign n828 = ~n773 & n827;
  assign n829 = ~n777 & ~n778;
  assign n830 = ~n781 & ~n783;
  assign n831 = n829 & n830;
  assign n832 = n828 & n831;
  assign n833 = n826 & n832;
  assign n834 = ~n792 & ~n795;
  assign n835 = ~n788 & n834;
  assign n836 = ~n800 & ~n804;
  assign n837 = ~n806 & ~n809;
  assign n838 = n836 & n837;
  assign n839 = n835 & n838;
  assign n840 = ~n813 & ~n815;
  assign n841 = ~n812 & n840;
  assign n842 = ~n816 & ~n818;
  assign n843 = ~n819 & ~n820;
  assign n844 = n842 & n843;
  assign n845 = n841 & n844;
  assign n846 = n839 & n845;
  assign n847 = n833 & n846;
  assign n848 = n743 & ~n746;
  assign n849 = ~n737 & ~n740;
  assign n850 = n848 & n849;
  assign n851 = n737 & n740;
  assign n852 = ~n743 & n746;
  assign n853 = n851 & n852;
  assign n854 = ~n850 & ~n853;
  assign n855 = ~n731 & ~n854;
  assign n856 = ~n740 & ~n746;
  assign n857 = n740 & n746;
  assign n858 = ~n856 & ~n857;
  assign n859 = n743 & ~n858;
  assign n860 = n737 & n859;
  assign n861 = n731 & n860;
  assign n862 = ~n855 & ~n861;
  assign n863 = n734 & ~n862;
  assign n864 = n847 & ~n863;
  assign n865 = ~pi170 & ~n864;
  assign n866 = pi170 & n864;
  assign n867 = ~n865 & ~n866;
  assign n868 = n504 & ~n867;
  assign n869 = pi067 & ~pi198;
  assign n870 = ~n504 & n869;
  assign po056 = n868 | n870;
  assign n872 = pi138 & n504;
  assign n873 = pi068 & ~pi198;
  assign n874 = ~n504 & n873;
  assign po057 = n872 | n874;
  assign n876 = pi131 & ~pi213;
  assign n877 = ~pi131 & pi213;
  assign n878 = ~n876 & ~n877;
  assign n879 = pi162 & ~pi210;
  assign n880 = ~pi162 & pi210;
  assign n881 = ~n879 & ~n880;
  assign n882 = pi161 & ~pi216;
  assign n883 = ~pi161 & pi216;
  assign n884 = ~n882 & ~n883;
  assign n885 = pi160 & ~pi203;
  assign n886 = ~pi160 & pi203;
  assign n887 = ~n885 & ~n886;
  assign n888 = pi159 & ~pi226;
  assign n889 = ~pi159 & pi226;
  assign n890 = ~n888 & ~n889;
  assign n891 = pi158 & ~pi222;
  assign n892 = ~pi158 & pi222;
  assign n893 = ~n891 & ~n892;
  assign n894 = n878 & n881;
  assign n895 = n884 & n894;
  assign n896 = n887 & n895;
  assign n897 = n890 & n896;
  assign n898 = n893 & n897;
  assign n899 = n878 & ~n881;
  assign n900 = n884 & n899;
  assign n901 = ~n887 & n900;
  assign n902 = n890 & n901;
  assign n903 = n893 & n902;
  assign n904 = ~n890 & n901;
  assign n905 = n893 & n904;
  assign n906 = ~n884 & n899;
  assign n907 = n887 & n906;
  assign n908 = n890 & n907;
  assign n909 = n893 & n908;
  assign n910 = ~n887 & n906;
  assign n911 = ~n890 & n910;
  assign n912 = n893 & n911;
  assign n913 = ~n890 & n896;
  assign n914 = ~n893 & n913;
  assign n915 = ~n887 & n895;
  assign n916 = n890 & n915;
  assign n917 = ~n893 & n916;
  assign n918 = ~n884 & n894;
  assign n919 = n887 & n918;
  assign n920 = n890 & n919;
  assign n921 = ~n893 & n920;
  assign n922 = ~n887 & n918;
  assign n923 = n890 & n922;
  assign n924 = ~n893 & n923;
  assign n925 = n887 & n900;
  assign n926 = ~n890 & n925;
  assign n927 = ~n893 & n926;
  assign n928 = ~n893 & n902;
  assign n929 = ~n890 & n907;
  assign n930 = ~n893 & n929;
  assign n931 = n893 & n916;
  assign n932 = ~n878 & n881;
  assign n933 = n884 & n932;
  assign n934 = ~n887 & n933;
  assign n935 = n890 & n934;
  assign n936 = n893 & n935;
  assign n937 = ~n884 & n932;
  assign n938 = n887 & n937;
  assign n939 = n890 & n938;
  assign n940 = n893 & n939;
  assign n941 = ~n890 & n938;
  assign n942 = n893 & n941;
  assign n943 = ~n878 & ~n881;
  assign n944 = n884 & n943;
  assign n945 = n887 & n944;
  assign n946 = n890 & n945;
  assign n947 = n893 & n946;
  assign n948 = ~n890 & n945;
  assign n949 = n893 & n948;
  assign n950 = ~n887 & n944;
  assign n951 = ~n890 & n950;
  assign n952 = n893 & n951;
  assign n953 = ~n884 & n943;
  assign n954 = ~n887 & n953;
  assign n955 = n890 & n954;
  assign n956 = n893 & n955;
  assign n957 = n887 & n933;
  assign n958 = n890 & n957;
  assign n959 = ~n893 & n958;
  assign n960 = ~n890 & n957;
  assign n961 = ~n893 & n960;
  assign n962 = ~n887 & n937;
  assign n963 = ~n890 & n962;
  assign n964 = ~n893 & n963;
  assign n965 = ~n893 & n946;
  assign n966 = ~n893 & n951;
  assign n967 = ~n890 & n919;
  assign n968 = n893 & n967;
  assign n969 = ~n893 & n955;
  assign n970 = ~n890 & n954;
  assign n971 = ~n893 & n970;
  assign n972 = ~n903 & ~n905;
  assign n973 = ~n898 & n972;
  assign n974 = ~n909 & ~n912;
  assign n975 = ~n914 & ~n917;
  assign n976 = n974 & n975;
  assign n977 = n973 & n976;
  assign n978 = ~n924 & ~n927;
  assign n979 = ~n921 & n978;
  assign n980 = ~n928 & ~n930;
  assign n981 = ~n931 & ~n936;
  assign n982 = n980 & n981;
  assign n983 = n979 & n982;
  assign n984 = n977 & n983;
  assign n985 = ~n942 & ~n947;
  assign n986 = ~n940 & n985;
  assign n987 = ~n949 & ~n952;
  assign n988 = ~n956 & ~n959;
  assign n989 = n987 & n988;
  assign n990 = n986 & n989;
  assign n991 = ~n964 & ~n965;
  assign n992 = ~n961 & n991;
  assign n993 = ~n966 & ~n968;
  assign n994 = ~n969 & ~n971;
  assign n995 = n993 & n994;
  assign n996 = n992 & n995;
  assign n997 = n990 & n996;
  assign n998 = n984 & n997;
  assign n999 = ~n884 & ~n893;
  assign n1000 = n884 & n893;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = n890 & ~n1001;
  assign n1003 = ~n878 & n1002;
  assign n1004 = ~n890 & n893;
  assign n1005 = n878 & n884;
  assign n1006 = n1004 & n1005;
  assign n1007 = ~n1003 & ~n1006;
  assign n1008 = n887 & ~n1007;
  assign n1009 = ~n890 & ~n893;
  assign n1010 = ~n887 & n1009;
  assign n1011 = n1005 & n1010;
  assign n1012 = ~n1008 & ~n1011;
  assign n1013 = n881 & ~n1012;
  assign n1014 = n998 & ~n1013;
  assign n1015 = ~pi178 & ~n1014;
  assign n1016 = pi178 & n1014;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = n504 & ~n1017;
  assign n1019 = pi069 & ~pi198;
  assign n1020 = ~n504 & n1019;
  assign po058 = n1018 | n1020;
  assign n1022 = pi146 & n504;
  assign n1023 = pi070 & ~pi198;
  assign n1024 = ~n504 & n1023;
  assign po059 = n1022 | n1024;
  assign n1026 = n893 & n929;
  assign n1027 = n890 & n925;
  assign n1028 = ~n893 & n1027;
  assign n1029 = ~n893 & n904;
  assign n1030 = ~n893 & n908;
  assign n1031 = n893 & n963;
  assign n1032 = n890 & n950;
  assign n1033 = n893 & n1032;
  assign n1034 = n887 & n953;
  assign n1035 = ~n890 & n1034;
  assign n1036 = n893 & n1035;
  assign n1037 = ~n893 & n941;
  assign n1038 = ~n893 & n948;
  assign n1039 = n890 & n1034;
  assign n1040 = ~n893 & n1039;
  assign n1041 = n893 & n923;
  assign n1042 = n893 & n926;
  assign n1043 = ~n905 & ~n1026;
  assign n1044 = ~n898 & n1043;
  assign n1045 = ~n914 & ~n921;
  assign n1046 = ~n924 & ~n1028;
  assign n1047 = n1045 & n1046;
  assign n1048 = n1044 & n1047;
  assign n1049 = ~n1029 & ~n1030;
  assign n1050 = ~n928 & n1049;
  assign n1051 = ~n940 & ~n1031;
  assign n1052 = n981 & n1051;
  assign n1053 = n1050 & n1052;
  assign n1054 = n1048 & n1053;
  assign n1055 = ~n949 & ~n1033;
  assign n1056 = ~n947 & n1055;
  assign n1057 = ~n959 & ~n1036;
  assign n1058 = ~n961 & ~n1037;
  assign n1059 = n1057 & n1058;
  assign n1060 = n1056 & n1059;
  assign n1061 = n993 & ~n1038;
  assign n1062 = ~n971 & ~n1040;
  assign n1063 = ~n1041 & ~n1042;
  assign n1064 = n1062 & n1063;
  assign n1065 = n1061 & n1064;
  assign n1066 = n1060 & n1065;
  assign n1067 = n1054 & n1066;
  assign n1068 = n890 & ~n893;
  assign n1069 = ~n1004 & ~n1068;
  assign n1070 = n884 & ~n1069;
  assign n1071 = ~n878 & n1070;
  assign n1072 = n878 & ~n884;
  assign n1073 = n1004 & n1072;
  assign n1074 = ~n1071 & ~n1073;
  assign n1075 = n881 & ~n1074;
  assign n1076 = ~n884 & n1009;
  assign n1077 = n899 & n1076;
  assign n1078 = ~n1075 & ~n1077;
  assign n1079 = ~n887 & ~n1078;
  assign n1080 = n1067 & ~n1079;
  assign n1081 = ~pi186 & ~n1080;
  assign n1082 = pi186 & n1080;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = n504 & ~n1083;
  assign n1085 = pi071 & ~pi198;
  assign n1086 = ~n504 & n1085;
  assign po060 = n1084 | n1086;
  assign n1088 = pi154 & n504;
  assign n1089 = pi072 & ~pi198;
  assign n1090 = ~n504 & n1089;
  assign po061 = n1088 | n1090;
  assign n1092 = pi151 & ~pi211;
  assign n1093 = ~pi151 & pi211;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = pi150 & ~pi220;
  assign n1096 = ~pi150 & pi220;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = pi149 & ~pi200;
  assign n1099 = ~pi149 & pi200;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = pi148 & ~pi207;
  assign n1102 = ~pi148 & pi207;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = pi147 & ~pi214;
  assign n1105 = ~pi147 & pi214;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = pi146 & ~pi225;
  assign n1108 = ~pi146 & pi225;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = n1094 & n1097;
  assign n1111 = n1100 & n1110;
  assign n1112 = n1103 & n1111;
  assign n1113 = n1106 & n1112;
  assign n1114 = n1109 & n1113;
  assign n1115 = ~n1106 & n1112;
  assign n1116 = n1109 & n1115;
  assign n1117 = ~n1103 & n1111;
  assign n1118 = ~n1106 & n1117;
  assign n1119 = n1109 & n1118;
  assign n1120 = ~n1100 & n1110;
  assign n1121 = ~n1103 & n1120;
  assign n1122 = n1106 & n1121;
  assign n1123 = n1109 & n1122;
  assign n1124 = n1094 & ~n1097;
  assign n1125 = n1100 & n1124;
  assign n1126 = ~n1103 & n1125;
  assign n1127 = ~n1106 & n1126;
  assign n1128 = n1109 & n1127;
  assign n1129 = ~n1100 & n1124;
  assign n1130 = n1103 & n1129;
  assign n1131 = n1106 & n1130;
  assign n1132 = n1109 & n1131;
  assign n1133 = ~n1103 & n1129;
  assign n1134 = ~n1106 & n1133;
  assign n1135 = n1109 & n1134;
  assign n1136 = ~n1109 & n1113;
  assign n1137 = n1106 & n1117;
  assign n1138 = ~n1109 & n1137;
  assign n1139 = ~n1109 & n1118;
  assign n1140 = n1103 & n1120;
  assign n1141 = ~n1106 & n1140;
  assign n1142 = ~n1109 & n1141;
  assign n1143 = ~n1106 & n1121;
  assign n1144 = ~n1109 & n1143;
  assign n1145 = n1103 & n1125;
  assign n1146 = ~n1106 & n1145;
  assign n1147 = ~n1109 & n1146;
  assign n1148 = ~n1109 & n1134;
  assign n1149 = ~n1094 & n1097;
  assign n1150 = n1100 & n1149;
  assign n1151 = ~n1103 & n1150;
  assign n1152 = n1106 & n1151;
  assign n1153 = n1109 & n1152;
  assign n1154 = ~n1100 & n1149;
  assign n1155 = n1103 & n1154;
  assign n1156 = ~n1106 & n1155;
  assign n1157 = n1109 & n1156;
  assign n1158 = ~n1103 & n1154;
  assign n1159 = n1106 & n1158;
  assign n1160 = n1109 & n1159;
  assign n1161 = ~n1106 & n1158;
  assign n1162 = n1109 & n1161;
  assign n1163 = ~n1094 & ~n1097;
  assign n1164 = n1100 & n1163;
  assign n1165 = n1103 & n1164;
  assign n1166 = n1106 & n1165;
  assign n1167 = n1109 & n1166;
  assign n1168 = ~n1103 & n1164;
  assign n1169 = n1106 & n1168;
  assign n1170 = n1109 & n1169;
  assign n1171 = ~n1100 & n1163;
  assign n1172 = n1103 & n1171;
  assign n1173 = n1106 & n1172;
  assign n1174 = n1109 & n1173;
  assign n1175 = n1103 & n1150;
  assign n1176 = n1106 & n1175;
  assign n1177 = ~n1109 & n1176;
  assign n1178 = ~n1106 & n1175;
  assign n1179 = ~n1109 & n1178;
  assign n1180 = ~n1109 & n1159;
  assign n1181 = ~n1109 & n1166;
  assign n1182 = ~n1109 & n1169;
  assign n1183 = ~n1106 & n1168;
  assign n1184 = ~n1109 & n1183;
  assign n1185 = ~n1106 & n1172;
  assign n1186 = ~n1109 & n1185;
  assign n1187 = ~n1116 & ~n1119;
  assign n1188 = ~n1114 & n1187;
  assign n1189 = ~n1123 & ~n1128;
  assign n1190 = ~n1132 & ~n1135;
  assign n1191 = n1189 & n1190;
  assign n1192 = n1188 & n1191;
  assign n1193 = ~n1138 & ~n1139;
  assign n1194 = ~n1136 & n1193;
  assign n1195 = ~n1142 & ~n1144;
  assign n1196 = ~n1147 & ~n1148;
  assign n1197 = n1195 & n1196;
  assign n1198 = n1194 & n1197;
  assign n1199 = n1192 & n1198;
  assign n1200 = ~n1157 & ~n1160;
  assign n1201 = ~n1153 & n1200;
  assign n1202 = ~n1162 & ~n1167;
  assign n1203 = ~n1170 & ~n1174;
  assign n1204 = n1202 & n1203;
  assign n1205 = n1201 & n1204;
  assign n1206 = ~n1179 & ~n1180;
  assign n1207 = ~n1177 & n1206;
  assign n1208 = ~n1181 & ~n1182;
  assign n1209 = ~n1184 & ~n1186;
  assign n1210 = n1208 & n1209;
  assign n1211 = n1207 & n1210;
  assign n1212 = n1205 & n1211;
  assign n1213 = n1199 & n1212;
  assign n1214 = ~n1100 & ~n1109;
  assign n1215 = n1097 & n1214;
  assign n1216 = n1100 & n1109;
  assign n1217 = ~n1097 & n1216;
  assign n1218 = ~n1215 & ~n1217;
  assign n1219 = ~n1106 & ~n1218;
  assign n1220 = ~n1094 & n1219;
  assign n1221 = ~n1214 & ~n1216;
  assign n1222 = n1106 & ~n1221;
  assign n1223 = ~n1097 & n1222;
  assign n1224 = n1094 & n1223;
  assign n1225 = ~n1220 & ~n1224;
  assign n1226 = n1103 & ~n1225;
  assign n1227 = n1213 & ~n1226;
  assign n1228 = ~pi194 & ~n1227;
  assign n1229 = pi194 & n1227;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = n504 & ~n1230;
  assign n1232 = pi073 & ~pi198;
  assign n1233 = ~n504 & n1232;
  assign po062 = n1231 | n1233;
  assign n1235 = pi162 & n504;
  assign n1236 = pi074 & ~pi198;
  assign n1237 = ~n504 & n1236;
  assign po063 = n1235 | n1237;
  assign n1239 = n1109 & n1137;
  assign n1240 = n1109 & n1143;
  assign n1241 = ~n1106 & n1130;
  assign n1242 = n1109 & n1241;
  assign n1243 = ~n1109 & n1127;
  assign n1244 = ~n1109 & n1241;
  assign n1245 = n1106 & n1133;
  assign n1246 = ~n1109 & n1245;
  assign n1247 = n1109 & n1176;
  assign n1248 = n1106 & n1155;
  assign n1249 = n1109 & n1248;
  assign n1250 = n1109 & n1183;
  assign n1251 = ~n1109 & n1248;
  assign n1252 = ~n1109 & n1173;
  assign n1253 = ~n1103 & n1171;
  assign n1254 = ~n1106 & n1253;
  assign n1255 = ~n1109 & n1254;
  assign n1256 = ~n1106 & ~n1109;
  assign n1257 = n1097 & n1256;
  assign n1258 = n1106 & n1109;
  assign n1259 = ~n1097 & n1258;
  assign n1260 = ~n1257 & ~n1259;
  assign n1261 = ~n1100 & ~n1260;
  assign n1262 = ~n1094 & n1261;
  assign n1263 = n1100 & n1258;
  assign n1264 = n1124 & n1263;
  assign n1265 = ~n1262 & ~n1264;
  assign n1266 = ~n1103 & ~n1265;
  assign n1267 = ~n1123 & ~n1239;
  assign n1268 = ~n1116 & n1267;
  assign n1269 = ~n1132 & ~n1240;
  assign n1270 = ~n1135 & ~n1242;
  assign n1271 = n1269 & n1270;
  assign n1272 = n1268 & n1271;
  assign n1273 = ~n1138 & ~n1142;
  assign n1274 = ~n1136 & n1273;
  assign n1275 = ~n1243 & ~n1244;
  assign n1276 = ~n1148 & ~n1246;
  assign n1277 = n1275 & n1276;
  assign n1278 = n1274 & n1277;
  assign n1279 = n1272 & n1278;
  assign n1280 = ~n1153 & ~n1249;
  assign n1281 = ~n1247 & n1280;
  assign n1282 = ~n1157 & ~n1162;
  assign n1283 = ~n1167 & ~n1250;
  assign n1284 = n1282 & n1283;
  assign n1285 = n1281 & n1284;
  assign n1286 = ~n1179 & ~n1251;
  assign n1287 = ~n1180 & ~n1181;
  assign n1288 = n1286 & n1287;
  assign n1289 = ~n1184 & ~n1252;
  assign n1290 = n1097 & n1100;
  assign n1291 = n1094 & n1290;
  assign n1292 = n1103 & n1256;
  assign n1293 = n1291 & n1292;
  assign n1294 = ~n1255 & ~n1293;
  assign n1295 = n1289 & n1294;
  assign n1296 = n1288 & n1295;
  assign n1297 = n1285 & n1296;
  assign n1298 = n1279 & n1297;
  assign n1299 = ~n1266 & n1298;
  assign n1300 = ~pi169 & ~n1299;
  assign n1301 = pi169 & n1299;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = n504 & ~n1302;
  assign n1304 = pi075 & ~pi198;
  assign n1305 = pi067 & pi198;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = ~n504 & ~n1306;
  assign po064 = n1303 | n1307;
  assign n1309 = pi137 & n504;
  assign n1310 = pi076 & ~pi198;
  assign n1311 = pi068 & pi198;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = ~n504 & ~n1312;
  assign po065 = n1309 | n1313;
  assign n1315 = pi155 & ~pi206;
  assign n1316 = ~pi155 & pi206;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = pi154 & ~pi217;
  assign n1319 = ~pi154 & pi217;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = pi159 & ~pi224;
  assign n1322 = ~pi159 & pi224;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = pi158 & ~pi199;
  assign n1325 = ~pi158 & pi199;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = pi157 & ~pi212;
  assign n1328 = ~pi157 & pi212;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = pi156 & ~pi221;
  assign n1331 = ~pi156 & pi221;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = ~n1317 & n1320;
  assign n1334 = ~n1323 & n1333;
  assign n1335 = n1326 & n1334;
  assign n1336 = n1329 & n1335;
  assign n1337 = ~n1332 & n1336;
  assign n1338 = n1317 & n1320;
  assign n1339 = ~n1323 & n1338;
  assign n1340 = n1326 & n1339;
  assign n1341 = ~n1329 & n1340;
  assign n1342 = ~n1332 & n1341;
  assign n1343 = ~n1326 & n1339;
  assign n1344 = n1329 & n1343;
  assign n1345 = n1332 & n1344;
  assign n1346 = ~n1329 & n1343;
  assign n1347 = n1332 & n1346;
  assign n1348 = ~n1326 & n1334;
  assign n1349 = ~n1329 & n1348;
  assign n1350 = n1332 & n1349;
  assign n1351 = ~n1332 & n1349;
  assign n1352 = n1317 & ~n1320;
  assign n1353 = ~n1323 & n1352;
  assign n1354 = n1326 & n1353;
  assign n1355 = n1329 & n1354;
  assign n1356 = n1332 & n1355;
  assign n1357 = ~n1329 & n1354;
  assign n1358 = n1332 & n1357;
  assign n1359 = ~n1317 & ~n1320;
  assign n1360 = ~n1323 & n1359;
  assign n1361 = n1326 & n1360;
  assign n1362 = ~n1329 & n1361;
  assign n1363 = n1332 & n1362;
  assign n1364 = ~n1326 & n1353;
  assign n1365 = n1329 & n1364;
  assign n1366 = n1332 & n1365;
  assign n1367 = ~n1332 & n1365;
  assign n1368 = ~n1326 & n1360;
  assign n1369 = ~n1329 & n1368;
  assign n1370 = n1332 & n1369;
  assign n1371 = ~n1332 & n1369;
  assign n1372 = n1323 & n1338;
  assign n1373 = n1326 & n1372;
  assign n1374 = n1329 & n1373;
  assign n1375 = n1332 & n1374;
  assign n1376 = n1323 & n1333;
  assign n1377 = n1326 & n1376;
  assign n1378 = ~n1329 & n1377;
  assign n1379 = n1332 & n1378;
  assign n1380 = ~n1329 & n1373;
  assign n1381 = ~n1332 & n1380;
  assign n1382 = ~n1326 & n1372;
  assign n1383 = n1329 & n1382;
  assign n1384 = n1332 & n1383;
  assign n1385 = ~n1326 & n1376;
  assign n1386 = n1329 & n1385;
  assign n1387 = n1332 & n1386;
  assign n1388 = ~n1332 & n1386;
  assign n1389 = ~n1329 & n1382;
  assign n1390 = ~n1332 & n1389;
  assign n1391 = n1323 & n1352;
  assign n1392 = n1326 & n1391;
  assign n1393 = n1329 & n1392;
  assign n1394 = n1332 & n1393;
  assign n1395 = n1323 & n1359;
  assign n1396 = n1326 & n1395;
  assign n1397 = n1329 & n1396;
  assign n1398 = n1332 & n1397;
  assign n1399 = ~n1332 & n1397;
  assign n1400 = ~n1329 & n1392;
  assign n1401 = n1332 & n1400;
  assign n1402 = ~n1326 & n1395;
  assign n1403 = ~n1329 & n1402;
  assign n1404 = n1332 & n1403;
  assign n1405 = ~n1326 & n1391;
  assign n1406 = ~n1329 & n1405;
  assign n1407 = ~n1332 & n1406;
  assign n1408 = ~n1332 & n1403;
  assign n1409 = n1329 & n1340;
  assign n1410 = ~n1332 & n1409;
  assign n1411 = ~n1323 & ~n1332;
  assign n1412 = ~n1320 & n1411;
  assign n1413 = n1323 & n1332;
  assign n1414 = n1320 & n1413;
  assign n1415 = ~n1412 & ~n1414;
  assign n1416 = n1326 & ~n1415;
  assign n1417 = ~n1317 & n1416;
  assign n1418 = ~n1326 & ~n1332;
  assign n1419 = n1323 & n1418;
  assign n1420 = n1352 & n1419;
  assign n1421 = ~n1417 & ~n1420;
  assign n1422 = n1329 & ~n1421;
  assign n1423 = ~n1342 & ~n1345;
  assign n1424 = ~n1337 & n1423;
  assign n1425 = ~n1347 & ~n1350;
  assign n1426 = ~n1351 & ~n1356;
  assign n1427 = n1425 & n1426;
  assign n1428 = n1424 & n1427;
  assign n1429 = ~n1363 & ~n1366;
  assign n1430 = ~n1358 & n1429;
  assign n1431 = ~n1367 & ~n1370;
  assign n1432 = ~n1371 & ~n1375;
  assign n1433 = n1431 & n1432;
  assign n1434 = n1430 & n1433;
  assign n1435 = n1428 & n1434;
  assign n1436 = ~n1381 & ~n1384;
  assign n1437 = ~n1379 & n1436;
  assign n1438 = ~n1387 & ~n1388;
  assign n1439 = ~n1390 & ~n1394;
  assign n1440 = n1438 & n1439;
  assign n1441 = n1437 & n1440;
  assign n1442 = ~n1398 & ~n1399;
  assign n1443 = ~n1401 & ~n1404;
  assign n1444 = n1442 & n1443;
  assign n1445 = ~n1407 & ~n1408;
  assign n1446 = ~n1329 & ~n1332;
  assign n1447 = n1326 & n1446;
  assign n1448 = n1320 & ~n1323;
  assign n1449 = ~n1317 & n1448;
  assign n1450 = n1447 & n1449;
  assign n1451 = ~n1410 & ~n1450;
  assign n1452 = n1445 & n1451;
  assign n1453 = n1444 & n1452;
  assign n1454 = n1441 & n1453;
  assign n1455 = n1435 & n1454;
  assign n1456 = ~n1422 & n1455;
  assign n1457 = ~pi177 & ~n1456;
  assign n1458 = pi177 & n1456;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = n504 & ~n1459;
  assign n1461 = pi077 & ~pi198;
  assign n1462 = pi069 & pi198;
  assign n1463 = ~n1461 & ~n1462;
  assign n1464 = ~n504 & ~n1463;
  assign po066 = n1460 | n1464;
  assign n1466 = pi145 & n504;
  assign n1467 = pi078 & ~pi198;
  assign n1468 = pi070 & pi198;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = ~n504 & ~n1469;
  assign po067 = n1466 | n1470;
  assign n1472 = n1109 & n1141;
  assign n1473 = n1106 & n1140;
  assign n1474 = ~n1109 & n1473;
  assign n1475 = n1109 & n1178;
  assign n1476 = ~n1106 & n1151;
  assign n1477 = ~n1109 & n1476;
  assign n1478 = ~n1119 & ~n1239;
  assign n1479 = ~n1114 & n1478;
  assign n1480 = ~n1240 & ~n1472;
  assign n1481 = n1190 & n1480;
  assign n1482 = n1479 & n1481;
  assign n1483 = ~n1142 & ~n1474;
  assign n1484 = ~n1138 & n1483;
  assign n1485 = ~n1144 & ~n1147;
  assign n1486 = ~n1244 & ~n1246;
  assign n1487 = n1485 & n1486;
  assign n1488 = n1484 & n1487;
  assign n1489 = n1482 & n1488;
  assign n1490 = ~n1157 & ~n1475;
  assign n1491 = ~n1247 & n1490;
  assign n1492 = ~n1160 & ~n1167;
  assign n1493 = ~n1170 & ~n1250;
  assign n1494 = n1492 & n1493;
  assign n1495 = n1491 & n1494;
  assign n1496 = ~n1179 & ~n1477;
  assign n1497 = ~n1177 & n1496;
  assign n1498 = ~n1184 & ~n1251;
  assign n1499 = ~n1186 & ~n1255;
  assign n1500 = n1498 & n1499;
  assign n1501 = n1497 & n1500;
  assign n1502 = n1495 & n1501;
  assign n1503 = n1489 & n1502;
  assign n1504 = ~n1106 & n1109;
  assign n1505 = n1103 & n1504;
  assign n1506 = n1106 & ~n1109;
  assign n1507 = ~n1103 & n1506;
  assign n1508 = ~n1505 & ~n1507;
  assign n1509 = n1094 & n1100;
  assign n1510 = ~n1094 & ~n1100;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n1508 & ~n1511;
  assign n1513 = ~n1097 & n1512;
  assign n1514 = n1503 & ~n1513;
  assign n1515 = ~pi185 & ~n1514;
  assign n1516 = pi185 & n1514;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = n504 & ~n1517;
  assign n1519 = pi079 & ~pi198;
  assign n1520 = pi071 & pi198;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n504 & ~n1521;
  assign po068 = n1518 | n1522;
  assign n1524 = pi153 & n504;
  assign n1525 = pi080 & ~pi198;
  assign n1526 = pi072 & pi198;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = ~n504 & ~n1527;
  assign po069 = n1524 | n1528;
  assign n1530 = n1332 & n1341;
  assign n1531 = n1329 & n1348;
  assign n1532 = ~n1332 & n1531;
  assign n1533 = ~n1332 & n1355;
  assign n1534 = n1329 & n1368;
  assign n1535 = n1332 & n1534;
  assign n1536 = ~n1329 & n1364;
  assign n1537 = ~n1332 & n1536;
  assign n1538 = n1329 & n1377;
  assign n1539 = ~n1332 & n1538;
  assign n1540 = n1332 & n1380;
  assign n1541 = ~n1329 & n1385;
  assign n1542 = ~n1332 & n1541;
  assign n1543 = ~n1329 & n1396;
  assign n1544 = ~n1332 & n1543;
  assign n1545 = n1329 & n1402;
  assign n1546 = ~n1332 & n1545;
  assign n1547 = n1332 & n1406;
  assign n1548 = n1332 & n1336;
  assign n1549 = ~n1411 & ~n1413;
  assign n1550 = n1326 & ~n1549;
  assign n1551 = ~n1320 & n1550;
  assign n1552 = ~n1317 & n1551;
  assign n1553 = ~n1323 & n1418;
  assign n1554 = n1338 & n1553;
  assign n1555 = ~n1552 & ~n1554;
  assign n1556 = ~n1329 & ~n1555;
  assign n1557 = ~n1530 & ~n1532;
  assign n1558 = ~n1337 & n1557;
  assign n1559 = ~n1350 & ~n1351;
  assign n1560 = ~n1358 & ~n1533;
  assign n1561 = n1559 & n1560;
  assign n1562 = n1558 & n1561;
  assign n1563 = ~n1366 & ~n1535;
  assign n1564 = ~n1363 & n1563;
  assign n1565 = ~n1367 & ~n1537;
  assign n1566 = ~n1375 & ~n1539;
  assign n1567 = n1565 & n1566;
  assign n1568 = n1564 & n1567;
  assign n1569 = n1562 & n1568;
  assign n1570 = ~n1379 & ~n1381;
  assign n1571 = ~n1540 & n1570;
  assign n1572 = ~n1387 & ~n1542;
  assign n1573 = ~n1394 & ~n1399;
  assign n1574 = n1572 & n1573;
  assign n1575 = n1571 & n1574;
  assign n1576 = ~n1401 & ~n1544;
  assign n1577 = ~n1546 & ~n1547;
  assign n1578 = n1576 & n1577;
  assign n1579 = ~n1407 & ~n1548;
  assign n1580 = n1320 & n1323;
  assign n1581 = n1317 & n1580;
  assign n1582 = n1329 & ~n1332;
  assign n1583 = ~n1326 & n1582;
  assign n1584 = n1581 & n1583;
  assign n1585 = ~n1410 & ~n1584;
  assign n1586 = n1579 & n1585;
  assign n1587 = n1578 & n1586;
  assign n1588 = n1575 & n1587;
  assign n1589 = n1569 & n1588;
  assign n1590 = ~n1556 & n1589;
  assign n1591 = ~pi193 & ~n1590;
  assign n1592 = pi193 & n1590;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = n504 & ~n1593;
  assign n1595 = pi081 & ~pi198;
  assign n1596 = pi073 & pi198;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n504 & ~n1597;
  assign po070 = n1594 | n1598;
  assign n1600 = pi161 & n504;
  assign n1601 = pi082 & ~pi198;
  assign n1602 = pi074 & pi198;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n504 & ~n1603;
  assign po071 = n1600 | n1604;
  assign n1606 = pi135 & ~pi237;
  assign n1607 = ~pi135 & pi237;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = pi134 & ~pi241;
  assign n1610 = ~pi134 & pi241;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = pi133 & ~pi233;
  assign n1613 = ~pi133 & pi233;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = pi132 & ~pi247;
  assign n1616 = ~pi132 & pi247;
  assign n1617 = ~n1615 & ~n1616;
  assign n1618 = pi131 & ~pi254;
  assign n1619 = ~pi131 & pi254;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = pi162 & ~pi251;
  assign n1622 = ~pi162 & pi251;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = n1608 & n1611;
  assign n1625 = n1614 & n1624;
  assign n1626 = n1617 & n1625;
  assign n1627 = n1620 & n1626;
  assign n1628 = n1623 & n1627;
  assign n1629 = ~n1614 & n1624;
  assign n1630 = n1617 & n1629;
  assign n1631 = n1620 & n1630;
  assign n1632 = n1623 & n1631;
  assign n1633 = ~n1620 & n1630;
  assign n1634 = n1623 & n1633;
  assign n1635 = n1608 & ~n1611;
  assign n1636 = n1614 & n1635;
  assign n1637 = ~n1617 & n1636;
  assign n1638 = ~n1620 & n1637;
  assign n1639 = n1623 & n1638;
  assign n1640 = ~n1614 & n1635;
  assign n1641 = n1617 & n1640;
  assign n1642 = n1620 & n1641;
  assign n1643 = n1623 & n1642;
  assign n1644 = ~n1617 & n1640;
  assign n1645 = n1620 & n1644;
  assign n1646 = n1623 & n1645;
  assign n1647 = ~n1620 & n1644;
  assign n1648 = n1623 & n1647;
  assign n1649 = ~n1620 & n1626;
  assign n1650 = ~n1623 & n1649;
  assign n1651 = ~n1617 & n1625;
  assign n1652 = n1620 & n1651;
  assign n1653 = ~n1623 & n1652;
  assign n1654 = ~n1617 & n1629;
  assign n1655 = n1620 & n1654;
  assign n1656 = ~n1623 & n1655;
  assign n1657 = n1617 & n1636;
  assign n1658 = n1620 & n1657;
  assign n1659 = ~n1623 & n1658;
  assign n1660 = ~n1620 & n1657;
  assign n1661 = ~n1623 & n1660;
  assign n1662 = n1620 & n1637;
  assign n1663 = ~n1623 & n1662;
  assign n1664 = ~n1620 & n1641;
  assign n1665 = ~n1623 & n1664;
  assign n1666 = ~n1608 & n1611;
  assign n1667 = n1614 & n1666;
  assign n1668 = n1617 & n1667;
  assign n1669 = n1620 & n1668;
  assign n1670 = n1623 & n1669;
  assign n1671 = ~n1614 & n1666;
  assign n1672 = n1617 & n1671;
  assign n1673 = ~n1620 & n1672;
  assign n1674 = n1623 & n1673;
  assign n1675 = ~n1617 & n1671;
  assign n1676 = n1620 & n1675;
  assign n1677 = n1623 & n1676;
  assign n1678 = ~n1608 & ~n1611;
  assign n1679 = n1614 & n1678;
  assign n1680 = n1617 & n1679;
  assign n1681 = ~n1620 & n1680;
  assign n1682 = n1623 & n1681;
  assign n1683 = ~n1617 & n1679;
  assign n1684 = ~n1620 & n1683;
  assign n1685 = n1623 & n1684;
  assign n1686 = ~n1614 & n1678;
  assign n1687 = n1617 & n1686;
  assign n1688 = n1620 & n1687;
  assign n1689 = n1623 & n1688;
  assign n1690 = ~n1617 & n1686;
  assign n1691 = n1620 & n1690;
  assign n1692 = n1623 & n1691;
  assign n1693 = ~n1617 & n1667;
  assign n1694 = n1620 & n1693;
  assign n1695 = ~n1623 & n1694;
  assign n1696 = ~n1620 & n1693;
  assign n1697 = ~n1623 & n1696;
  assign n1698 = ~n1620 & n1675;
  assign n1699 = ~n1623 & n1698;
  assign n1700 = n1620 & n1680;
  assign n1701 = ~n1623 & n1700;
  assign n1702 = ~n1623 & n1681;
  assign n1703 = ~n1620 & n1687;
  assign n1704 = ~n1623 & n1703;
  assign n1705 = ~n1623 & n1691;
  assign n1706 = n1617 & ~n1623;
  assign n1707 = ~n1614 & n1706;
  assign n1708 = ~n1617 & n1623;
  assign n1709 = n1614 & n1708;
  assign n1710 = ~n1707 & ~n1709;
  assign n1711 = n1620 & ~n1710;
  assign n1712 = ~n1608 & n1711;
  assign n1713 = ~n1614 & ~n1623;
  assign n1714 = n1614 & n1623;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n1620 & ~n1715;
  assign n1717 = ~n1617 & n1716;
  assign n1718 = n1608 & n1717;
  assign n1719 = ~n1712 & ~n1718;
  assign n1720 = n1611 & ~n1719;
  assign n1721 = ~n1632 & ~n1634;
  assign n1722 = ~n1628 & n1721;
  assign n1723 = ~n1639 & ~n1643;
  assign n1724 = ~n1646 & ~n1648;
  assign n1725 = n1723 & n1724;
  assign n1726 = n1722 & n1725;
  assign n1727 = ~n1653 & ~n1656;
  assign n1728 = ~n1650 & n1727;
  assign n1729 = ~n1659 & ~n1661;
  assign n1730 = ~n1663 & ~n1665;
  assign n1731 = n1729 & n1730;
  assign n1732 = n1728 & n1731;
  assign n1733 = n1726 & n1732;
  assign n1734 = ~n1674 & ~n1677;
  assign n1735 = ~n1670 & n1734;
  assign n1736 = ~n1682 & ~n1685;
  assign n1737 = ~n1689 & ~n1692;
  assign n1738 = n1736 & n1737;
  assign n1739 = n1735 & n1738;
  assign n1740 = ~n1697 & ~n1699;
  assign n1741 = ~n1695 & n1740;
  assign n1742 = ~n1701 & ~n1702;
  assign n1743 = ~n1704 & ~n1705;
  assign n1744 = n1742 & n1743;
  assign n1745 = n1741 & n1744;
  assign n1746 = n1739 & n1745;
  assign n1747 = n1733 & n1746;
  assign n1748 = ~n1720 & n1747;
  assign n1749 = ~pi168 & ~n1748;
  assign n1750 = pi168 & n1748;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = n504 & ~n1751;
  assign n1753 = pi083 & ~pi198;
  assign n1754 = pi075 & pi198;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n504 & ~n1755;
  assign po072 = n1752 | n1756;
  assign n1758 = pi136 & n504;
  assign n1759 = pi084 & ~pi198;
  assign n1760 = pi076 & pi198;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = ~n504 & ~n1761;
  assign po073 = n1758 | n1762;
  assign n1764 = pi143 & ~pi253;
  assign n1765 = ~pi143 & pi253;
  assign n1766 = ~n1764 & ~n1765;
  assign n1767 = pi142 & ~pi243;
  assign n1768 = ~pi142 & pi243;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = pi141 & ~pi232;
  assign n1771 = ~pi141 & pi232;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = pi140 & ~pi238;
  assign n1774 = ~pi140 & pi238;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = pi139 & ~pi250;
  assign n1777 = ~pi139 & pi250;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = pi138 & ~pi235;
  assign n1780 = ~pi138 & pi235;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = n1766 & n1769;
  assign n1783 = n1772 & n1782;
  assign n1784 = ~n1775 & n1783;
  assign n1785 = ~n1778 & n1784;
  assign n1786 = n1781 & n1785;
  assign n1787 = ~n1772 & n1782;
  assign n1788 = n1775 & n1787;
  assign n1789 = n1778 & n1788;
  assign n1790 = n1781 & n1789;
  assign n1791 = n1766 & ~n1769;
  assign n1792 = n1772 & n1791;
  assign n1793 = n1775 & n1792;
  assign n1794 = ~n1778 & n1793;
  assign n1795 = n1781 & n1794;
  assign n1796 = ~n1775 & n1792;
  assign n1797 = n1778 & n1796;
  assign n1798 = n1781 & n1797;
  assign n1799 = ~n1772 & n1791;
  assign n1800 = n1775 & n1799;
  assign n1801 = ~n1778 & n1800;
  assign n1802 = n1781 & n1801;
  assign n1803 = ~n1775 & n1799;
  assign n1804 = n1778 & n1803;
  assign n1805 = n1781 & n1804;
  assign n1806 = ~n1778 & n1803;
  assign n1807 = n1781 & n1806;
  assign n1808 = n1775 & n1783;
  assign n1809 = ~n1778 & n1808;
  assign n1810 = ~n1781 & n1809;
  assign n1811 = ~n1781 & n1789;
  assign n1812 = ~n1775 & n1787;
  assign n1813 = n1778 & n1812;
  assign n1814 = ~n1781 & n1813;
  assign n1815 = ~n1778 & n1812;
  assign n1816 = ~n1781 & n1815;
  assign n1817 = ~n1781 & n1797;
  assign n1818 = ~n1781 & n1801;
  assign n1819 = ~n1781 & n1804;
  assign n1820 = ~n1766 & n1769;
  assign n1821 = n1772 & n1820;
  assign n1822 = n1775 & n1821;
  assign n1823 = n1778 & n1822;
  assign n1824 = n1781 & n1823;
  assign n1825 = ~n1775 & n1821;
  assign n1826 = n1778 & n1825;
  assign n1827 = n1781 & n1826;
  assign n1828 = ~n1778 & n1825;
  assign n1829 = n1781 & n1828;
  assign n1830 = ~n1772 & n1820;
  assign n1831 = ~n1775 & n1830;
  assign n1832 = ~n1778 & n1831;
  assign n1833 = n1781 & n1832;
  assign n1834 = ~n1766 & ~n1769;
  assign n1835 = n1772 & n1834;
  assign n1836 = n1775 & n1835;
  assign n1837 = n1778 & n1836;
  assign n1838 = n1781 & n1837;
  assign n1839 = ~n1772 & n1834;
  assign n1840 = n1775 & n1839;
  assign n1841 = ~n1778 & n1840;
  assign n1842 = n1781 & n1841;
  assign n1843 = ~n1775 & n1839;
  assign n1844 = n1778 & n1843;
  assign n1845 = n1781 & n1844;
  assign n1846 = ~n1778 & n1822;
  assign n1847 = ~n1781 & n1846;
  assign n1848 = n1775 & n1830;
  assign n1849 = n1778 & n1848;
  assign n1850 = ~n1781 & n1849;
  assign n1851 = ~n1778 & n1848;
  assign n1852 = ~n1781 & n1851;
  assign n1853 = n1778 & n1831;
  assign n1854 = ~n1781 & n1853;
  assign n1855 = ~n1781 & n1837;
  assign n1856 = ~n1775 & n1835;
  assign n1857 = ~n1778 & n1856;
  assign n1858 = ~n1781 & n1857;
  assign n1859 = ~n1778 & n1843;
  assign n1860 = ~n1781 & n1859;
  assign n1861 = ~n1775 & ~n1781;
  assign n1862 = n1772 & n1861;
  assign n1863 = n1775 & n1781;
  assign n1864 = ~n1772 & n1863;
  assign n1865 = ~n1862 & ~n1864;
  assign n1866 = n1778 & ~n1865;
  assign n1867 = ~n1766 & n1866;
  assign n1868 = n1766 & n1772;
  assign n1869 = ~n1778 & ~n1781;
  assign n1870 = n1775 & n1869;
  assign n1871 = n1868 & n1870;
  assign n1872 = ~n1867 & ~n1871;
  assign n1873 = ~n1769 & ~n1872;
  assign n1874 = ~n1790 & ~n1795;
  assign n1875 = ~n1786 & n1874;
  assign n1876 = ~n1798 & ~n1802;
  assign n1877 = ~n1805 & ~n1807;
  assign n1878 = n1876 & n1877;
  assign n1879 = n1875 & n1878;
  assign n1880 = ~n1811 & ~n1814;
  assign n1881 = ~n1810 & n1880;
  assign n1882 = ~n1816 & ~n1817;
  assign n1883 = ~n1818 & ~n1819;
  assign n1884 = n1882 & n1883;
  assign n1885 = n1881 & n1884;
  assign n1886 = n1879 & n1885;
  assign n1887 = ~n1827 & ~n1829;
  assign n1888 = ~n1824 & n1887;
  assign n1889 = ~n1833 & ~n1838;
  assign n1890 = ~n1842 & ~n1845;
  assign n1891 = n1889 & n1890;
  assign n1892 = n1888 & n1891;
  assign n1893 = ~n1847 & ~n1850;
  assign n1894 = ~n1852 & ~n1854;
  assign n1895 = n1893 & n1894;
  assign n1896 = ~n1855 & ~n1858;
  assign n1897 = ~n1778 & n1781;
  assign n1898 = n1775 & n1897;
  assign n1899 = n1769 & n1772;
  assign n1900 = n1766 & n1899;
  assign n1901 = n1898 & n1900;
  assign n1902 = ~n1860 & ~n1901;
  assign n1903 = n1896 & n1902;
  assign n1904 = n1895 & n1903;
  assign n1905 = n1892 & n1904;
  assign n1906 = n1886 & n1905;
  assign n1907 = ~n1873 & n1906;
  assign n1908 = ~pi176 & ~n1907;
  assign n1909 = pi176 & n1907;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n504 & ~n1910;
  assign n1912 = pi085 & ~pi198;
  assign n1913 = pi077 & pi198;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n504 & ~n1914;
  assign po074 = n1911 | n1915;
  assign n1917 = pi144 & n504;
  assign n1918 = pi086 & ~pi198;
  assign n1919 = pi078 & pi198;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n504 & ~n1920;
  assign po075 = n1917 | n1921;
  assign n1923 = n1778 & n1784;
  assign n1924 = n1781 & n1923;
  assign n1925 = n1781 & n1813;
  assign n1926 = n1778 & n1800;
  assign n1927 = n1781 & n1926;
  assign n1928 = n1778 & n1808;
  assign n1929 = ~n1781 & n1928;
  assign n1930 = n1778 & n1793;
  assign n1931 = ~n1781 & n1930;
  assign n1932 = ~n1778 & n1796;
  assign n1933 = ~n1781 & n1932;
  assign n1934 = n1781 & n1846;
  assign n1935 = n1781 & n1857;
  assign n1936 = n1781 & n1859;
  assign n1937 = ~n1781 & n1832;
  assign n1938 = ~n1778 & n1836;
  assign n1939 = ~n1781 & n1938;
  assign n1940 = n1778 & n1840;
  assign n1941 = ~n1781 & n1940;
  assign n1942 = ~n1786 & ~n1925;
  assign n1943 = ~n1924 & n1942;
  assign n1944 = ~n1798 & ~n1927;
  assign n1945 = ~n1802 & ~n1807;
  assign n1946 = n1944 & n1945;
  assign n1947 = n1943 & n1946;
  assign n1948 = ~n1810 & ~n1811;
  assign n1949 = ~n1929 & n1948;
  assign n1950 = ~n1931 & ~n1933;
  assign n1951 = n1883 & n1950;
  assign n1952 = n1949 & n1951;
  assign n1953 = n1947 & n1952;
  assign n1954 = ~n1827 & ~n1833;
  assign n1955 = ~n1934 & n1954;
  assign n1956 = ~n1838 & ~n1935;
  assign n1957 = ~n1845 & ~n1936;
  assign n1958 = n1956 & n1957;
  assign n1959 = n1955 & n1958;
  assign n1960 = ~n1854 & ~n1937;
  assign n1961 = ~n1847 & n1960;
  assign n1962 = ~n1855 & ~n1939;
  assign n1963 = ~n1858 & ~n1941;
  assign n1964 = n1962 & n1963;
  assign n1965 = n1961 & n1964;
  assign n1966 = n1959 & n1965;
  assign n1967 = n1953 & n1966;
  assign n1968 = n1766 & ~n1778;
  assign n1969 = ~n1766 & n1778;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~n1865 & ~n1970;
  assign n1972 = n1769 & n1971;
  assign n1973 = n1967 & ~n1972;
  assign n1974 = ~pi184 & ~n1973;
  assign n1975 = pi184 & n1973;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = n504 & ~n1976;
  assign n1978 = pi087 & ~pi198;
  assign n1979 = pi079 & pi198;
  assign n1980 = ~n1978 & ~n1979;
  assign n1981 = ~n504 & ~n1980;
  assign po076 = n1977 | n1981;
  assign n1983 = pi152 & n504;
  assign n1984 = pi088 & ~pi198;
  assign n1985 = pi080 & pi198;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~n504 & ~n1986;
  assign po077 = n1983 | n1987;
  assign n1989 = n740 & n760;
  assign n1990 = ~n743 & n1989;
  assign n1991 = n746 & n1990;
  assign n1992 = n746 & n780;
  assign n1993 = n746 & n782;
  assign n1994 = ~n746 & n755;
  assign n1995 = n743 & n1989;
  assign n1996 = ~n746 & n1995;
  assign n1997 = ~n743 & n779;
  assign n1998 = ~n746 & n1997;
  assign n1999 = n746 & n814;
  assign n2000 = n746 & n817;
  assign n2001 = ~n740 & n797;
  assign n2002 = ~n743 & n2001;
  assign n2003 = n746 & n2002;
  assign n2004 = ~n743 & n793;
  assign n2005 = ~n746 & n2004;
  assign n2006 = ~n746 & n2002;
  assign n2007 = n743 & n807;
  assign n2008 = ~n746 & n2007;
  assign n2009 = n740 & ~n746;
  assign n2010 = ~n737 & n2009;
  assign n2011 = ~n740 & n746;
  assign n2012 = n737 & n2011;
  assign n2013 = ~n2010 & ~n2012;
  assign n2014 = n743 & ~n2013;
  assign n2015 = ~n731 & n2014;
  assign n2016 = ~n737 & ~n746;
  assign n2017 = n737 & n746;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = ~n743 & ~n2018;
  assign n2020 = ~n740 & n2019;
  assign n2021 = n731 & n2020;
  assign n2022 = ~n2015 & ~n2021;
  assign n2023 = n734 & ~n2022;
  assign n2024 = ~n756 & ~n1991;
  assign n2025 = ~n751 & n2024;
  assign n2026 = ~n763 & ~n765;
  assign n2027 = ~n1992 & ~n1993;
  assign n2028 = n2026 & n2027;
  assign n2029 = n2025 & n2028;
  assign n2030 = ~n776 & ~n1994;
  assign n2031 = ~n775 & n2030;
  assign n2032 = ~n777 & ~n1996;
  assign n2033 = ~n781 & ~n1998;
  assign n2034 = n2032 & n2033;
  assign n2035 = n2031 & n2034;
  assign n2036 = n2029 & n2035;
  assign n2037 = ~n795 & ~n1999;
  assign n2038 = ~n788 & n2037;
  assign n2039 = ~n800 & ~n2000;
  assign n2040 = ~n806 & ~n2003;
  assign n2041 = n2039 & n2040;
  assign n2042 = n2038 & n2041;
  assign n2043 = ~n813 & ~n2005;
  assign n2044 = ~n812 & n2043;
  assign n2045 = ~n818 & ~n2006;
  assign n2046 = ~n820 & ~n2008;
  assign n2047 = n2045 & n2046;
  assign n2048 = n2044 & n2047;
  assign n2049 = n2042 & n2048;
  assign n2050 = n2036 & n2049;
  assign n2051 = ~n2023 & n2050;
  assign n2052 = ~pi192 & ~n2051;
  assign n2053 = pi192 & n2051;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n504 & ~n2054;
  assign n2056 = pi089 & ~pi198;
  assign n2057 = pi081 & pi198;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n504 & ~n2058;
  assign po078 = n2055 | n2059;
  assign n2061 = pi160 & n504;
  assign n2062 = pi090 & ~pi198;
  assign n2063 = pi082 & pi198;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = ~n504 & ~n2064;
  assign po079 = n2061 | n2065;
  assign n2067 = ~n1332 & n1344;
  assign n2068 = ~n1332 & n1534;
  assign n2069 = n1332 & n1389;
  assign n2070 = n1329 & n1405;
  assign n2071 = n1332 & n2070;
  assign n2072 = ~n1345 & ~n2067;
  assign n2073 = ~n1342 & n2072;
  assign n2074 = ~n1351 & ~n1532;
  assign n2075 = ~n1356 & ~n1363;
  assign n2076 = n2074 & n2075;
  assign n2077 = n2073 & n2076;
  assign n2078 = ~n1367 & ~n2068;
  assign n2079 = ~n1535 & n2078;
  assign n2080 = ~n1370 & ~n1537;
  assign n2081 = n1566 & n2080;
  assign n2082 = n2079 & n2081;
  assign n2083 = n2077 & n2082;
  assign n2084 = n1438 & ~n1540;
  assign n2085 = ~n1390 & ~n2069;
  assign n2086 = n1442 & n2085;
  assign n2087 = n2084 & n2086;
  assign n2088 = ~n1544 & ~n2071;
  assign n2089 = ~n1401 & n2088;
  assign n2090 = ~n1408 & ~n1547;
  assign n2091 = ~n1410 & ~n1548;
  assign n2092 = n2090 & n2091;
  assign n2093 = n2089 & n2092;
  assign n2094 = n2087 & n2093;
  assign n2095 = n2083 & n2094;
  assign n2096 = ~n1323 & n1332;
  assign n2097 = n1323 & ~n1332;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = n1320 & ~n2098;
  assign n2100 = ~n1317 & n2099;
  assign n2101 = n1352 & n1411;
  assign n2102 = ~n2100 & ~n2101;
  assign n2103 = ~n1329 & ~n2102;
  assign n2104 = n1323 & n1582;
  assign n2105 = n1352 & n2104;
  assign n2106 = ~n2103 & ~n2105;
  assign n2107 = n1326 & ~n2106;
  assign n2108 = n2095 & ~n2107;
  assign n2109 = ~pi167 & ~n2108;
  assign n2110 = pi167 & n2108;
  assign n2111 = ~n2109 & ~n2110;
  assign n2112 = n504 & ~n2111;
  assign n2113 = pi091 & ~pi198;
  assign n2114 = pi083 & pi198;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = ~n504 & ~n2115;
  assign po080 = n2112 | n2116;
  assign n2118 = pi135 & n504;
  assign n2119 = pi092 & ~pi198;
  assign n2120 = pi084 & pi198;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = ~n504 & ~n2121;
  assign po081 = n2118 | n2122;
  assign n2124 = ~n1116 & ~n1239;
  assign n2125 = ~n1114 & n2124;
  assign n2126 = ~n1128 & ~n1472;
  assign n2127 = n1270 & n2126;
  assign n2128 = n2125 & n2127;
  assign n2129 = ~n1139 & ~n1474;
  assign n2130 = ~n1136 & n2129;
  assign n2131 = ~n1142 & ~n1147;
  assign n2132 = ~n1243 & ~n1246;
  assign n2133 = n2131 & n2132;
  assign n2134 = n2130 & n2133;
  assign n2135 = n2128 & n2134;
  assign n2136 = ~n1160 & ~n1249;
  assign n2137 = ~n1475 & n2136;
  assign n2138 = ~n1174 & ~n1250;
  assign n2139 = n1202 & n2138;
  assign n2140 = n2137 & n2139;
  assign n2141 = ~n1180 & ~n1477;
  assign n2142 = ~n1179 & n2141;
  assign n2143 = ~n1182 & ~n1252;
  assign n2144 = n1499 & n2143;
  assign n2145 = n2142 & n2144;
  assign n2146 = n2140 & n2145;
  assign n2147 = n2135 & n2146;
  assign n2148 = ~n1094 & ~n1106;
  assign n2149 = n1094 & n1106;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = n1103 & ~n1109;
  assign n2152 = n1100 & n2151;
  assign n2153 = ~n1103 & n1109;
  assign n2154 = ~n1100 & n2153;
  assign n2155 = ~n2152 & ~n2154;
  assign n2156 = ~n2150 & ~n2155;
  assign n2157 = ~n1097 & n2156;
  assign n2158 = n2147 & ~n2157;
  assign n2159 = ~pi175 & ~n2158;
  assign n2160 = pi175 & n2158;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = n504 & ~n2161;
  assign n2163 = pi093 & ~pi198;
  assign n2164 = pi085 & pi198;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = ~n504 & ~n2165;
  assign po082 = n2162 | n2166;
  assign n2168 = pi143 & n504;
  assign n2169 = pi094 & ~pi198;
  assign n2170 = pi086 & pi198;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = ~n504 & ~n2171;
  assign po083 = n2168 | n2172;
  assign n2174 = pi139 & ~pi239;
  assign n2175 = ~pi139 & pi239;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = pi138 & ~pi234;
  assign n2178 = ~pi138 & pi234;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = pi137 & ~pi244;
  assign n2181 = ~pi137 & pi244;
  assign n2182 = ~n2180 & ~n2181;
  assign n2183 = pi136 & ~pi227;
  assign n2184 = ~pi136 & pi227;
  assign n2185 = ~n2183 & ~n2184;
  assign n2186 = pi135 & ~pi249;
  assign n2187 = ~pi135 & pi249;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = pi134 & ~pi230;
  assign n2190 = ~pi134 & pi230;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = n2176 & n2179;
  assign n2193 = n2182 & n2192;
  assign n2194 = ~n2185 & n2193;
  assign n2195 = ~n2188 & n2194;
  assign n2196 = n2191 & n2195;
  assign n2197 = ~n2182 & n2192;
  assign n2198 = n2185 & n2197;
  assign n2199 = n2188 & n2198;
  assign n2200 = n2191 & n2199;
  assign n2201 = ~n2185 & n2197;
  assign n2202 = ~n2188 & n2201;
  assign n2203 = n2191 & n2202;
  assign n2204 = n2176 & ~n2179;
  assign n2205 = n2182 & n2204;
  assign n2206 = n2185 & n2205;
  assign n2207 = ~n2188 & n2206;
  assign n2208 = n2191 & n2207;
  assign n2209 = ~n2185 & n2205;
  assign n2210 = ~n2188 & n2209;
  assign n2211 = n2191 & n2210;
  assign n2212 = ~n2182 & n2204;
  assign n2213 = n2185 & n2212;
  assign n2214 = n2188 & n2213;
  assign n2215 = n2191 & n2214;
  assign n2216 = ~n2185 & n2212;
  assign n2217 = n2188 & n2216;
  assign n2218 = n2191 & n2217;
  assign n2219 = n2185 & n2193;
  assign n2220 = n2188 & n2219;
  assign n2221 = ~n2191 & n2220;
  assign n2222 = ~n2191 & n2195;
  assign n2223 = n2188 & n2206;
  assign n2224 = ~n2191 & n2223;
  assign n2225 = n2188 & n2209;
  assign n2226 = ~n2191 & n2225;
  assign n2227 = ~n2191 & n2210;
  assign n2228 = ~n2188 & n2213;
  assign n2229 = ~n2191 & n2228;
  assign n2230 = ~n2188 & n2216;
  assign n2231 = ~n2191 & n2230;
  assign n2232 = ~n2176 & n2179;
  assign n2233 = n2182 & n2232;
  assign n2234 = ~n2185 & n2233;
  assign n2235 = ~n2188 & n2234;
  assign n2236 = n2191 & n2235;
  assign n2237 = ~n2182 & n2232;
  assign n2238 = n2185 & n2237;
  assign n2239 = n2188 & n2238;
  assign n2240 = n2191 & n2239;
  assign n2241 = ~n2185 & n2237;
  assign n2242 = n2188 & n2241;
  assign n2243 = n2191 & n2242;
  assign n2244 = ~n2188 & n2241;
  assign n2245 = n2191 & n2244;
  assign n2246 = ~n2176 & ~n2179;
  assign n2247 = n2182 & n2246;
  assign n2248 = n2185 & n2247;
  assign n2249 = ~n2188 & n2248;
  assign n2250 = n2191 & n2249;
  assign n2251 = ~n2185 & n2247;
  assign n2252 = n2188 & n2251;
  assign n2253 = n2191 & n2252;
  assign n2254 = ~n2182 & n2246;
  assign n2255 = n2185 & n2254;
  assign n2256 = ~n2188 & n2255;
  assign n2257 = n2191 & n2256;
  assign n2258 = n2185 & n2233;
  assign n2259 = n2188 & n2258;
  assign n2260 = ~n2191 & n2259;
  assign n2261 = n2188 & n2234;
  assign n2262 = ~n2191 & n2261;
  assign n2263 = ~n2191 & n2244;
  assign n2264 = ~n2191 & n2249;
  assign n2265 = ~n2188 & n2251;
  assign n2266 = ~n2191 & n2265;
  assign n2267 = n2188 & n2255;
  assign n2268 = ~n2191 & n2267;
  assign n2269 = ~n2185 & n2254;
  assign n2270 = ~n2188 & n2269;
  assign n2271 = ~n2191 & n2270;
  assign n2272 = ~n2200 & ~n2203;
  assign n2273 = ~n2196 & n2272;
  assign n2274 = ~n2208 & ~n2211;
  assign n2275 = ~n2215 & ~n2218;
  assign n2276 = n2274 & n2275;
  assign n2277 = n2273 & n2276;
  assign n2278 = ~n2222 & ~n2224;
  assign n2279 = ~n2221 & n2278;
  assign n2280 = ~n2226 & ~n2227;
  assign n2281 = ~n2229 & ~n2231;
  assign n2282 = n2280 & n2281;
  assign n2283 = n2279 & n2282;
  assign n2284 = n2277 & n2283;
  assign n2285 = ~n2240 & ~n2243;
  assign n2286 = ~n2236 & n2285;
  assign n2287 = ~n2245 & ~n2250;
  assign n2288 = ~n2253 & ~n2257;
  assign n2289 = n2287 & n2288;
  assign n2290 = n2286 & n2289;
  assign n2291 = ~n2262 & ~n2263;
  assign n2292 = ~n2260 & n2291;
  assign n2293 = ~n2264 & ~n2266;
  assign n2294 = ~n2268 & ~n2271;
  assign n2295 = n2293 & n2294;
  assign n2296 = n2292 & n2295;
  assign n2297 = n2290 & n2296;
  assign n2298 = n2284 & n2297;
  assign n2299 = ~n2182 & ~n2191;
  assign n2300 = n2182 & n2191;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2176 & ~n2188;
  assign n2303 = n2176 & n2188;
  assign n2304 = ~n2302 & ~n2303;
  assign n2305 = ~n2301 & ~n2304;
  assign n2306 = n2185 & n2305;
  assign n2307 = n2179 & n2306;
  assign n2308 = n2298 & ~n2307;
  assign n2309 = ~pi183 & ~n2308;
  assign n2310 = pi183 & n2308;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = n504 & ~n2311;
  assign n2313 = pi095 & ~pi198;
  assign n2314 = pi087 & pi198;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~n504 & ~n2315;
  assign po084 = n2312 | n2316;
  assign n2318 = pi151 & n504;
  assign n2319 = pi096 & ~pi198;
  assign n2320 = pi088 & pi198;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = ~n504 & ~n2321;
  assign po085 = n2318 | n2322;
  assign n2324 = n1781 & n1928;
  assign n2325 = ~n1778 & n1788;
  assign n2326 = ~n1781 & n2325;
  assign n2327 = n1781 & n1853;
  assign n2328 = ~n1781 & n1828;
  assign n2329 = ~n1786 & ~n1924;
  assign n2330 = ~n2324 & n2329;
  assign n2331 = ~n1807 & ~n1927;
  assign n2332 = n1874 & n2331;
  assign n2333 = n2330 & n2332;
  assign n2334 = ~n1810 & ~n2326;
  assign n2335 = ~n1929 & n2334;
  assign n2336 = ~n1814 & ~n1817;
  assign n2337 = ~n1818 & ~n1933;
  assign n2338 = n2336 & n2337;
  assign n2339 = n2335 & n2338;
  assign n2340 = n2333 & n2339;
  assign n2341 = ~n1827 & ~n1934;
  assign n2342 = ~n1824 & n2341;
  assign n2343 = ~n1935 & ~n2327;
  assign n2344 = n1890 & n2343;
  assign n2345 = n2342 & n2344;
  assign n2346 = ~n1850 & ~n1854;
  assign n2347 = ~n2328 & n2346;
  assign n2348 = ~n1855 & ~n1937;
  assign n2349 = ~n1860 & ~n1939;
  assign n2350 = n2348 & n2349;
  assign n2351 = n2347 & n2350;
  assign n2352 = n2345 & n2351;
  assign n2353 = n2340 & n2352;
  assign n2354 = n1778 & ~n1781;
  assign n2355 = ~n1769 & ~n1775;
  assign n2356 = n2354 & n2355;
  assign n2357 = n1769 & n1775;
  assign n2358 = n1897 & n2357;
  assign n2359 = ~n2356 & ~n2358;
  assign n2360 = ~n1766 & ~n2359;
  assign n2361 = ~n1769 & ~n1781;
  assign n2362 = n1769 & n1781;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~n1778 & ~n2363;
  assign n2365 = ~n1775 & n2364;
  assign n2366 = n1766 & n2365;
  assign n2367 = ~n2360 & ~n2366;
  assign n2368 = ~n1772 & ~n2367;
  assign n2369 = n2353 & ~n2368;
  assign n2370 = ~pi191 & ~n2369;
  assign n2371 = pi191 & n2369;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = n504 & ~n2372;
  assign n2374 = pi097 & ~pi198;
  assign n2375 = pi089 & pi198;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = ~n504 & ~n2376;
  assign po086 = n2373 | n2377;
  assign n2379 = pi159 & n504;
  assign n2380 = pi098 & ~pi198;
  assign n2381 = pi090 & pi198;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = ~n504 & ~n2382;
  assign po087 = n2379 | n2383;
  assign n2385 = n1942 & ~n2324;
  assign n2386 = ~n1795 & ~n1927;
  assign n2387 = ~n1802 & ~n1805;
  assign n2388 = n2386 & n2387;
  assign n2389 = n2385 & n2388;
  assign n2390 = ~n1811 & ~n2326;
  assign n2391 = ~n1810 & n2390;
  assign n2392 = ~n1816 & ~n1931;
  assign n2393 = ~n1817 & ~n1933;
  assign n2394 = n2392 & n2393;
  assign n2395 = n2391 & n2394;
  assign n2396 = n2389 & n2395;
  assign n2397 = n1887 & ~n1934;
  assign n2398 = ~n1838 & ~n2327;
  assign n2399 = ~n1842 & ~n1936;
  assign n2400 = n2398 & n2399;
  assign n2401 = n2397 & n2400;
  assign n2402 = n1894 & ~n2328;
  assign n2403 = ~n1858 & ~n1939;
  assign n2404 = ~n1860 & ~n1941;
  assign n2405 = n2403 & n2404;
  assign n2406 = n2402 & n2405;
  assign n2407 = n2401 & n2406;
  assign n2408 = n2396 & n2407;
  assign n2409 = n1775 & ~n1781;
  assign n2410 = n1769 & n2409;
  assign n2411 = ~n1775 & n1781;
  assign n2412 = ~n1769 & n2411;
  assign n2413 = ~n2410 & ~n2412;
  assign n2414 = ~n1766 & ~n2413;
  assign n2415 = n1782 & n1861;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = n1778 & ~n2416;
  assign n2418 = ~n1775 & n1897;
  assign n2419 = n1791 & n2418;
  assign n2420 = ~n2417 & ~n2419;
  assign n2421 = n1772 & ~n2420;
  assign n2422 = n2408 & ~n2421;
  assign n2423 = ~pi166 & ~n2422;
  assign n2424 = pi166 & n2422;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = n504 & ~n2425;
  assign n2427 = pi099 & ~pi198;
  assign n2428 = pi091 & pi198;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n504 & ~n2429;
  assign po088 = n2426 | n2430;
  assign n2432 = pi134 & n504;
  assign n2433 = pi100 & ~pi198;
  assign n2434 = pi092 & pi198;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = ~n504 & ~n2435;
  assign po089 = n2432 | n2436;
  assign n2438 = n1623 & n1655;
  assign n2439 = n1623 & n1660;
  assign n2440 = n1623 & n1662;
  assign n2441 = ~n1623 & n1633;
  assign n2442 = ~n1623 & n1638;
  assign n2443 = ~n1623 & n1645;
  assign n2444 = ~n1620 & n1668;
  assign n2445 = n1623 & n2444;
  assign n2446 = n1620 & n1672;
  assign n2447 = n1623 & n2446;
  assign n2448 = n1623 & n1703;
  assign n2449 = n1620 & n1683;
  assign n2450 = ~n1623 & n2449;
  assign n2451 = ~n1623 & n1688;
  assign n2452 = ~n1620 & n1690;
  assign n2453 = ~n1623 & n2452;
  assign n2454 = ~n1634 & ~n2438;
  assign n2455 = ~n1628 & n2454;
  assign n2456 = ~n2439 & ~n2440;
  assign n2457 = ~n1643 & ~n1648;
  assign n2458 = n2456 & n2457;
  assign n2459 = n2455 & n2458;
  assign n2460 = ~n1653 & ~n2441;
  assign n2461 = ~n1650 & n2460;
  assign n2462 = ~n1656 & ~n1661;
  assign n2463 = ~n2442 & ~n2443;
  assign n2464 = n2462 & n2463;
  assign n2465 = n2461 & n2464;
  assign n2466 = n2459 & n2465;
  assign n2467 = ~n2445 & ~n2447;
  assign n2468 = ~n1670 & n2467;
  assign n2469 = ~n1685 & ~n1689;
  assign n2470 = ~n1692 & ~n2448;
  assign n2471 = n2469 & n2470;
  assign n2472 = n2468 & n2471;
  assign n2473 = ~n1699 & ~n1701;
  assign n2474 = ~n1697 & n2473;
  assign n2475 = ~n2450 & ~n2451;
  assign n2476 = ~n1704 & ~n2453;
  assign n2477 = n2475 & n2476;
  assign n2478 = n2474 & n2477;
  assign n2479 = n2472 & n2478;
  assign n2480 = n2466 & n2479;
  assign n2481 = ~n1706 & ~n1708;
  assign n2482 = ~n1620 & ~n2481;
  assign n2483 = ~n1608 & n2482;
  assign n2484 = n1620 & ~n1623;
  assign n2485 = n1608 & n1617;
  assign n2486 = n2484 & n2485;
  assign n2487 = ~n2483 & ~n2486;
  assign n2488 = n1614 & ~n2487;
  assign n2489 = n1608 & ~n1614;
  assign n2490 = ~n1620 & n1623;
  assign n2491 = ~n1617 & n2490;
  assign n2492 = n2489 & n2491;
  assign n2493 = ~n2488 & ~n2492;
  assign n2494 = n1611 & ~n2493;
  assign n2495 = n2480 & ~n2494;
  assign n2496 = ~pi174 & ~n2495;
  assign n2497 = pi174 & n2495;
  assign n2498 = ~n2496 & ~n2497;
  assign n2499 = n504 & ~n2498;
  assign n2500 = pi101 & ~pi198;
  assign n2501 = pi093 & pi198;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = ~n504 & ~n2502;
  assign po090 = n2499 | n2503;
  assign n2505 = pi142 & n504;
  assign n2506 = pi102 & ~pi198;
  assign n2507 = pi094 & pi198;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = ~n504 & ~n2508;
  assign po091 = n2505 | n2509;
  assign n2511 = n1320 & ~n1326;
  assign n2512 = ~n1320 & n1326;
  assign n2513 = ~n2511 & ~n2512;
  assign n2514 = n1332 & ~n2513;
  assign n2515 = ~n1323 & n2514;
  assign n2516 = ~n1317 & n2515;
  assign n2517 = n1326 & ~n1332;
  assign n2518 = n1323 & n2517;
  assign n2519 = n1338 & n2518;
  assign n2520 = ~n2516 & ~n2519;
  assign n2521 = n1329 & ~n2520;
  assign n2522 = ~n1342 & ~n1530;
  assign n2523 = ~n1337 & n2522;
  assign n2524 = ~n1347 & ~n2067;
  assign n2525 = n1426 & n2524;
  assign n2526 = n2523 & n2525;
  assign n2527 = n1429 & ~n1533;
  assign n2528 = ~n1537 & ~n2068;
  assign n2529 = n1432 & n2528;
  assign n2530 = n2527 & n2529;
  assign n2531 = n2526 & n2530;
  assign n2532 = ~n1379 & ~n1384;
  assign n2533 = ~n1539 & n2532;
  assign n2534 = ~n1388 & ~n2069;
  assign n2535 = ~n1398 & ~n1542;
  assign n2536 = n2534 & n2535;
  assign n2537 = n2533 & n2536;
  assign n2538 = ~n1546 & ~n2071;
  assign n2539 = n1576 & n2538;
  assign n2540 = ~n1404 & ~n1407;
  assign n2541 = ~n1320 & n1323;
  assign n2542 = n1317 & n2541;
  assign n2543 = n1447 & n2542;
  assign n2544 = ~n1548 & ~n2543;
  assign n2545 = n2540 & n2544;
  assign n2546 = n2539 & n2545;
  assign n2547 = n2537 & n2546;
  assign n2548 = n2531 & n2547;
  assign n2549 = ~n2521 & n2548;
  assign n2550 = ~pi182 & ~n2549;
  assign n2551 = pi182 & n2549;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = n504 & ~n2552;
  assign n2554 = pi103 & ~pi198;
  assign n2555 = pi095 & pi198;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n504 & ~n2556;
  assign po092 = n2553 | n2557;
  assign n2559 = pi150 & n504;
  assign n2560 = pi104 & ~pi198;
  assign n2561 = pi096 & pi198;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~n504 & ~n2562;
  assign po093 = n2559 | n2563;
  assign n2565 = n1623 & n1658;
  assign n2566 = ~n1623 & n1631;
  assign n2567 = n1623 & n2449;
  assign n2568 = ~n1623 & n1673;
  assign n2569 = ~n2439 & ~n2565;
  assign n2570 = ~n1639 & ~n1646;
  assign n2571 = n2569 & n2570;
  assign n2572 = n2455 & n2571;
  assign n2573 = ~n1653 & ~n2566;
  assign n2574 = ~n1650 & n2573;
  assign n2575 = ~n1659 & ~n2442;
  assign n2576 = ~n1665 & ~n2443;
  assign n2577 = n2575 & n2576;
  assign n2578 = n2574 & n2577;
  assign n2579 = n2572 & n2578;
  assign n2580 = ~n1674 & ~n2447;
  assign n2581 = ~n2445 & n2580;
  assign n2582 = ~n1677 & ~n2567;
  assign n2583 = n2469 & n2582;
  assign n2584 = n2581 & n2583;
  assign n2585 = ~n1699 & ~n2568;
  assign n2586 = ~n1695 & n2585;
  assign n2587 = ~n2450 & ~n2453;
  assign n2588 = n1742 & n2587;
  assign n2589 = n2586 & n2588;
  assign n2590 = n2584 & n2589;
  assign n2591 = n2579 & n2590;
  assign n2592 = n1611 & n2484;
  assign n2593 = ~n1611 & n2490;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n1614 & ~n2594;
  assign n2596 = ~n1608 & n2595;
  assign n2597 = ~n1620 & ~n1623;
  assign n2598 = n1620 & n1623;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = n1614 & ~n2599;
  assign n2601 = n1611 & n2600;
  assign n2602 = n1608 & n2601;
  assign n2603 = ~n2596 & ~n2602;
  assign n2604 = ~n1617 & ~n2603;
  assign n2605 = n2591 & ~n2604;
  assign n2606 = ~pi190 & ~n2605;
  assign n2607 = pi190 & n2605;
  assign n2608 = ~n2606 & ~n2607;
  assign n2609 = n504 & ~n2608;
  assign n2610 = pi105 & ~pi198;
  assign n2611 = pi097 & pi198;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n504 & ~n2612;
  assign po094 = n2609 | n2613;
  assign n2615 = pi158 & n504;
  assign n2616 = pi106 & ~pi198;
  assign n2617 = pi098 & pi198;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n504 & ~n2618;
  assign po095 = n2615 | n2619;
  assign n2621 = pi155 & ~pi204;
  assign n2622 = ~pi155 & pi204;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = pi154 & ~pi208;
  assign n2625 = ~pi154 & pi208;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = pi153 & ~pi215;
  assign n2628 = ~pi153 & pi215;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = pi152 & ~pi223;
  assign n2631 = ~pi152 & pi223;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = pi151 & ~pi201;
  assign n2634 = ~pi151 & pi201;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = pi150 & ~pi219;
  assign n2637 = ~pi150 & pi219;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = n2623 & n2626;
  assign n2640 = n2629 & n2639;
  assign n2641 = n2632 & n2640;
  assign n2642 = n2635 & n2641;
  assign n2643 = n2638 & n2642;
  assign n2644 = ~n2632 & n2640;
  assign n2645 = ~n2635 & n2644;
  assign n2646 = n2638 & n2645;
  assign n2647 = ~n2629 & n2639;
  assign n2648 = n2632 & n2647;
  assign n2649 = n2635 & n2648;
  assign n2650 = n2638 & n2649;
  assign n2651 = ~n2635 & n2648;
  assign n2652 = n2638 & n2651;
  assign n2653 = ~n2632 & n2647;
  assign n2654 = n2635 & n2653;
  assign n2655 = n2638 & n2654;
  assign n2656 = n2623 & ~n2626;
  assign n2657 = n2629 & n2656;
  assign n2658 = ~n2632 & n2657;
  assign n2659 = ~n2635 & n2658;
  assign n2660 = n2638 & n2659;
  assign n2661 = ~n2629 & n2656;
  assign n2662 = n2632 & n2661;
  assign n2663 = n2635 & n2662;
  assign n2664 = n2638 & n2663;
  assign n2665 = ~n2635 & n2641;
  assign n2666 = ~n2638 & n2665;
  assign n2667 = ~n2638 & n2649;
  assign n2668 = ~n2638 & n2654;
  assign n2669 = ~n2635 & n2653;
  assign n2670 = ~n2638 & n2669;
  assign n2671 = ~n2638 & n2659;
  assign n2672 = ~n2635 & n2662;
  assign n2673 = ~n2638 & n2672;
  assign n2674 = ~n2632 & n2661;
  assign n2675 = n2635 & n2674;
  assign n2676 = ~n2638 & n2675;
  assign n2677 = ~n2623 & n2626;
  assign n2678 = n2629 & n2677;
  assign n2679 = n2632 & n2678;
  assign n2680 = ~n2635 & n2679;
  assign n2681 = n2638 & n2680;
  assign n2682 = ~n2629 & n2677;
  assign n2683 = n2632 & n2682;
  assign n2684 = ~n2635 & n2683;
  assign n2685 = n2638 & n2684;
  assign n2686 = ~n2632 & n2682;
  assign n2687 = n2635 & n2686;
  assign n2688 = n2638 & n2687;
  assign n2689 = ~n2623 & ~n2626;
  assign n2690 = n2629 & n2689;
  assign n2691 = n2632 & n2690;
  assign n2692 = n2635 & n2691;
  assign n2693 = n2638 & n2692;
  assign n2694 = ~n2629 & n2689;
  assign n2695 = n2632 & n2694;
  assign n2696 = ~n2635 & n2695;
  assign n2697 = n2638 & n2696;
  assign n2698 = ~n2632 & n2694;
  assign n2699 = n2635 & n2698;
  assign n2700 = n2638 & n2699;
  assign n2701 = ~n2635 & n2698;
  assign n2702 = n2638 & n2701;
  assign n2703 = ~n2638 & n2680;
  assign n2704 = n2635 & n2683;
  assign n2705 = ~n2638 & n2704;
  assign n2706 = ~n2635 & n2686;
  assign n2707 = ~n2638 & n2706;
  assign n2708 = ~n2635 & n2691;
  assign n2709 = ~n2638 & n2708;
  assign n2710 = ~n2632 & n2690;
  assign n2711 = n2635 & n2710;
  assign n2712 = ~n2638 & n2711;
  assign n2713 = ~n2635 & n2710;
  assign n2714 = ~n2638 & n2713;
  assign n2715 = n2635 & n2695;
  assign n2716 = ~n2638 & n2715;
  assign n2717 = ~n2646 & ~n2650;
  assign n2718 = ~n2643 & n2717;
  assign n2719 = ~n2652 & ~n2655;
  assign n2720 = ~n2660 & ~n2664;
  assign n2721 = n2719 & n2720;
  assign n2722 = n2718 & n2721;
  assign n2723 = ~n2667 & ~n2668;
  assign n2724 = ~n2666 & n2723;
  assign n2725 = ~n2670 & ~n2671;
  assign n2726 = ~n2673 & ~n2676;
  assign n2727 = n2725 & n2726;
  assign n2728 = n2724 & n2727;
  assign n2729 = n2722 & n2728;
  assign n2730 = ~n2685 & ~n2688;
  assign n2731 = ~n2681 & n2730;
  assign n2732 = ~n2693 & ~n2697;
  assign n2733 = ~n2700 & ~n2702;
  assign n2734 = n2732 & n2733;
  assign n2735 = n2731 & n2734;
  assign n2736 = ~n2705 & ~n2707;
  assign n2737 = ~n2703 & n2736;
  assign n2738 = ~n2709 & ~n2712;
  assign n2739 = ~n2714 & ~n2716;
  assign n2740 = n2738 & n2739;
  assign n2741 = n2737 & n2740;
  assign n2742 = n2735 & n2741;
  assign n2743 = n2729 & n2742;
  assign n2744 = ~n2629 & ~n2638;
  assign n2745 = n2629 & n2638;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = ~n2623 & ~n2746;
  assign n2748 = ~n2629 & n2638;
  assign n2749 = n2623 & n2748;
  assign n2750 = ~n2747 & ~n2749;
  assign n2751 = ~n2632 & ~n2750;
  assign n2752 = n2632 & ~n2638;
  assign n2753 = n2623 & n2629;
  assign n2754 = n2752 & n2753;
  assign n2755 = ~n2751 & ~n2754;
  assign n2756 = n2635 & ~n2755;
  assign n2757 = ~n2626 & n2756;
  assign n2758 = n2743 & ~n2757;
  assign n2759 = ~pi165 & ~n2758;
  assign n2760 = pi165 & n2758;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = n504 & ~n2761;
  assign n2763 = pi107 & ~pi198;
  assign n2764 = pi099 & pi198;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = ~n504 & ~n2765;
  assign po096 = n2762 | n2766;
  assign n2768 = pi133 & n504;
  assign n2769 = pi108 & ~pi198;
  assign n2770 = pi100 & pi198;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = ~n504 & ~n2771;
  assign po097 = n2768 | n2772;
  assign n2774 = ~n2188 & n2219;
  assign n2775 = n2191 & n2774;
  assign n2776 = n2191 & n2223;
  assign n2777 = n2191 & n2228;
  assign n2778 = n2188 & n2194;
  assign n2779 = ~n2191 & n2778;
  assign n2780 = ~n2191 & n2202;
  assign n2781 = ~n2191 & n2207;
  assign n2782 = n2191 & n2261;
  assign n2783 = ~n2188 & n2238;
  assign n2784 = n2191 & n2783;
  assign n2785 = n2188 & n2248;
  assign n2786 = n2191 & n2785;
  assign n2787 = ~n2188 & n2258;
  assign n2788 = ~n2191 & n2787;
  assign n2789 = ~n2191 & n2242;
  assign n2790 = n2188 & n2269;
  assign n2791 = ~n2191 & n2790;
  assign n2792 = n2185 & ~n2191;
  assign n2793 = ~n2185 & n2191;
  assign n2794 = ~n2792 & ~n2793;
  assign n2795 = ~n2188 & ~n2794;
  assign n2796 = ~n2176 & n2795;
  assign n2797 = n2188 & ~n2191;
  assign n2798 = n2176 & n2185;
  assign n2799 = n2797 & n2798;
  assign n2800 = ~n2796 & ~n2799;
  assign n2801 = ~n2182 & ~n2800;
  assign n2802 = ~n2179 & n2801;
  assign n2803 = ~n2196 & ~n2200;
  assign n2804 = ~n2775 & n2803;
  assign n2805 = ~n2211 & ~n2776;
  assign n2806 = ~n2218 & ~n2777;
  assign n2807 = n2805 & n2806;
  assign n2808 = n2804 & n2807;
  assign n2809 = ~n2222 & ~n2780;
  assign n2810 = ~n2779 & n2809;
  assign n2811 = ~n2224 & ~n2781;
  assign n2812 = n2281 & n2811;
  assign n2813 = n2810 & n2812;
  assign n2814 = n2808 & n2813;
  assign n2815 = ~n2243 & ~n2784;
  assign n2816 = ~n2782 & n2815;
  assign n2817 = ~n2245 & ~n2786;
  assign n2818 = ~n2250 & ~n2253;
  assign n2819 = n2817 & n2818;
  assign n2820 = n2816 & n2819;
  assign n2821 = ~n2260 & ~n2788;
  assign n2822 = ~n2263 & ~n2789;
  assign n2823 = n2821 & n2822;
  assign n2824 = ~n2266 & ~n2268;
  assign n2825 = n2179 & n2182;
  assign n2826 = n2176 & n2825;
  assign n2827 = n2188 & n2191;
  assign n2828 = ~n2185 & n2827;
  assign n2829 = n2826 & n2828;
  assign n2830 = ~n2791 & ~n2829;
  assign n2831 = n2824 & n2830;
  assign n2832 = n2823 & n2831;
  assign n2833 = n2820 & n2832;
  assign n2834 = n2814 & n2833;
  assign n2835 = ~n2802 & n2834;
  assign n2836 = ~pi173 & ~n2835;
  assign n2837 = pi173 & n2835;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = n504 & ~n2838;
  assign n2840 = pi109 & ~pi198;
  assign n2841 = pi101 & pi198;
  assign n2842 = ~n2840 & ~n2841;
  assign n2843 = ~n504 & ~n2842;
  assign po098 = n2839 | n2843;
  assign n2845 = pi141 & n504;
  assign n2846 = pi110 & ~pi198;
  assign n2847 = pi102 & pi198;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = ~n504 & ~n2848;
  assign po099 = n2845 | n2849;
  assign n2851 = n746 & n774;
  assign n2852 = ~n740 & n770;
  assign n2853 = ~n743 & n2852;
  assign n2854 = ~n746 & n2853;
  assign n2855 = n743 & n2001;
  assign n2856 = n746 & n2855;
  assign n2857 = n743 & n786;
  assign n2858 = ~n746 & n2857;
  assign n2859 = ~n751 & ~n758;
  assign n2860 = ~n2851 & n2859;
  assign n2861 = ~n765 & ~n1991;
  assign n2862 = ~n769 & ~n1992;
  assign n2863 = n2861 & n2862;
  assign n2864 = n2860 & n2863;
  assign n2865 = ~n776 & ~n2854;
  assign n2866 = ~n773 & n2865;
  assign n2867 = ~n1994 & ~n1996;
  assign n2868 = ~n777 & ~n783;
  assign n2869 = n2867 & n2868;
  assign n2870 = n2866 & n2869;
  assign n2871 = n2864 & n2870;
  assign n2872 = ~n795 & ~n800;
  assign n2873 = ~n1999 & n2872;
  assign n2874 = ~n2003 & ~n2856;
  assign n2875 = ~n804 & ~n809;
  assign n2876 = n2874 & n2875;
  assign n2877 = n2873 & n2876;
  assign n2878 = ~n813 & ~n2858;
  assign n2879 = ~n815 & ~n2005;
  assign n2880 = n2878 & n2879;
  assign n2881 = n734 & n737;
  assign n2882 = n731 & n2881;
  assign n2883 = n743 & n746;
  assign n2884 = ~n740 & n2883;
  assign n2885 = n2882 & n2884;
  assign n2886 = ~n2008 & ~n2885;
  assign n2887 = n842 & n2886;
  assign n2888 = n2880 & n2887;
  assign n2889 = n2877 & n2888;
  assign n2890 = n2871 & n2889;
  assign n2891 = ~n734 & ~n737;
  assign n2892 = ~n743 & ~n746;
  assign n2893 = n2891 & n2892;
  assign n2894 = n2881 & n2883;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = ~n731 & ~n2895;
  assign n2897 = ~n737 & n848;
  assign n2898 = n747 & n2897;
  assign n2899 = ~n2896 & ~n2898;
  assign n2900 = n740 & ~n2899;
  assign n2901 = n2890 & ~n2900;
  assign n2902 = ~pi181 & ~n2901;
  assign n2903 = pi181 & n2901;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = n504 & ~n2904;
  assign n2906 = pi111 & ~pi198;
  assign n2907 = pi103 & pi198;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = ~n504 & ~n2908;
  assign po100 = n2905 | n2909;
  assign n2911 = pi149 & n504;
  assign n2912 = pi112 & ~pi198;
  assign n2913 = pi104 & pi198;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = ~n504 & ~n2914;
  assign po101 = n2911 | n2915;
  assign n2917 = n2635 & n2644;
  assign n2918 = n2638 & n2917;
  assign n2919 = n2638 & n2669;
  assign n2920 = n2632 & n2657;
  assign n2921 = ~n2635 & n2920;
  assign n2922 = n2638 & n2921;
  assign n2923 = ~n2638 & n2642;
  assign n2924 = ~n2638 & n2645;
  assign n2925 = n2635 & n2658;
  assign n2926 = ~n2638 & n2925;
  assign n2927 = n2635 & n2679;
  assign n2928 = n2638 & n2927;
  assign n2929 = ~n2632 & n2678;
  assign n2930 = ~n2635 & n2929;
  assign n2931 = n2638 & n2930;
  assign n2932 = n2638 & n2715;
  assign n2933 = n2635 & n2929;
  assign n2934 = ~n2638 & n2933;
  assign n2935 = ~n2638 & n2684;
  assign n2936 = ~n2638 & n2696;
  assign n2937 = n2719 & ~n2918;
  assign n2938 = ~n2919 & ~n2922;
  assign n2939 = n2720 & n2938;
  assign n2940 = n2937 & n2939;
  assign n2941 = ~n2666 & ~n2924;
  assign n2942 = ~n2923 & n2941;
  assign n2943 = ~n2667 & ~n2926;
  assign n2944 = n2726 & n2943;
  assign n2945 = n2942 & n2944;
  assign n2946 = n2940 & n2945;
  assign n2947 = ~n2685 & ~n2931;
  assign n2948 = ~n2928 & n2947;
  assign n2949 = ~n2688 & ~n2693;
  assign n2950 = ~n2702 & ~n2932;
  assign n2951 = n2949 & n2950;
  assign n2952 = n2948 & n2951;
  assign n2953 = ~n2934 & ~n2935;
  assign n2954 = ~n2707 & ~n2709;
  assign n2955 = n2953 & n2954;
  assign n2956 = ~n2626 & ~n2629;
  assign n2957 = n2623 & n2956;
  assign n2958 = ~n2635 & ~n2638;
  assign n2959 = ~n2632 & n2958;
  assign n2960 = n2957 & n2959;
  assign n2961 = ~n2936 & ~n2960;
  assign n2962 = n2739 & n2961;
  assign n2963 = n2955 & n2962;
  assign n2964 = n2952 & n2963;
  assign n2965 = n2946 & n2964;
  assign n2966 = n2635 & ~n2638;
  assign n2967 = n2626 & n2966;
  assign n2968 = ~n2635 & n2638;
  assign n2969 = ~n2626 & n2968;
  assign n2970 = ~n2967 & ~n2969;
  assign n2971 = ~n2623 & ~n2970;
  assign n2972 = n2635 & n2638;
  assign n2973 = n2656 & n2972;
  assign n2974 = ~n2971 & ~n2973;
  assign n2975 = n2632 & ~n2974;
  assign n2976 = n2629 & n2975;
  assign n2977 = n2965 & ~n2976;
  assign n2978 = ~pi189 & ~n2977;
  assign n2979 = pi189 & n2977;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = n504 & ~n2980;
  assign n2982 = pi113 & ~pi198;
  assign n2983 = pi105 & pi198;
  assign n2984 = ~n2982 & ~n2983;
  assign n2985 = ~n504 & ~n2984;
  assign po102 = n2981 | n2985;
  assign n2987 = pi157 & n504;
  assign n2988 = pi114 & ~pi198;
  assign n2989 = pi106 & pi198;
  assign n2990 = ~n2988 & ~n2989;
  assign n2991 = ~n504 & ~n2990;
  assign po103 = n2987 | n2991;
  assign n2993 = n890 & n910;
  assign n2994 = ~n893 & n2993;
  assign n2995 = n893 & n1039;
  assign n2996 = ~n893 & n1032;
  assign n2997 = n893 & n1027;
  assign n2998 = ~n912 & ~n1026;
  assign n2999 = ~n909 & n2998;
  assign n3000 = ~n924 & ~n1029;
  assign n3001 = n975 & n3000;
  assign n3002 = n2999 & n3001;
  assign n3003 = ~n930 & ~n931;
  assign n3004 = ~n1030 & n3003;
  assign n3005 = ~n940 & ~n2994;
  assign n3006 = ~n947 & ~n1031;
  assign n3007 = n3005 & n3006;
  assign n3008 = n3004 & n3007;
  assign n3009 = n3002 & n3008;
  assign n3010 = ~n952 & ~n2995;
  assign n3011 = ~n1033 & n3010;
  assign n3012 = ~n964 & ~n1037;
  assign n3013 = n988 & n3012;
  assign n3014 = n3011 & n3013;
  assign n3015 = ~n1038 & ~n2996;
  assign n3016 = ~n965 & n3015;
  assign n3017 = ~n968 & ~n971;
  assign n3018 = ~n1041 & ~n2997;
  assign n3019 = n3017 & n3018;
  assign n3020 = n3016 & n3019;
  assign n3021 = n3014 & n3020;
  assign n3022 = n3009 & n3021;
  assign n3023 = ~n890 & ~n1001;
  assign n3024 = ~n887 & n3023;
  assign n3025 = n878 & n3024;
  assign n3026 = ~n884 & ~n887;
  assign n3027 = n1068 & n3026;
  assign n3028 = n884 & n887;
  assign n3029 = n1004 & n3028;
  assign n3030 = ~n3027 & ~n3029;
  assign n3031 = ~n878 & ~n3030;
  assign n3032 = ~n3025 & ~n3031;
  assign n3033 = n881 & ~n3032;
  assign n3034 = n3022 & ~n3033;
  assign n3035 = ~pi164 & ~n3034;
  assign n3036 = pi164 & n3034;
  assign n3037 = ~n3035 & ~n3036;
  assign n3038 = n504 & ~n3037;
  assign n3039 = pi115 & ~pi198;
  assign n3040 = pi107 & pi198;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n504 & ~n3041;
  assign po104 = n3038 | n3042;
  assign n3044 = pi132 & n504;
  assign n3045 = pi116 & ~pi198;
  assign n3046 = pi108 & pi198;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = ~n504 & ~n3047;
  assign po105 = n3044 | n3048;
  assign n3050 = ~n903 & ~n912;
  assign n3051 = ~n898 & n3050;
  assign n3052 = ~n921 & ~n1028;
  assign n3053 = n975 & n3052;
  assign n3054 = n3051 & n3053;
  assign n3055 = ~n1029 & ~n2994;
  assign n3056 = ~n927 & n3055;
  assign n3057 = ~n936 & ~n942;
  assign n3058 = n3006 & n3057;
  assign n3059 = n3056 & n3058;
  assign n3060 = n3054 & n3059;
  assign n3061 = ~n1036 & ~n2995;
  assign n3062 = ~n952 & n3061;
  assign n3063 = ~n959 & ~n964;
  assign n3064 = n3015 & n3063;
  assign n3065 = n3062 & n3064;
  assign n3066 = ~n968 & ~n1040;
  assign n3067 = ~n966 & n3066;
  assign n3068 = ~n969 & ~n1041;
  assign n3069 = ~n1042 & ~n2997;
  assign n3070 = n3068 & n3069;
  assign n3071 = n3067 & n3070;
  assign n3072 = n3065 & n3071;
  assign n3073 = n3060 & n3072;
  assign n3074 = n884 & n1009;
  assign n3075 = n890 & n893;
  assign n3076 = ~n884 & n3075;
  assign n3077 = ~n3074 & ~n3076;
  assign n3078 = ~n887 & ~n3077;
  assign n3079 = ~n878 & n3078;
  assign n3080 = ~n1009 & ~n3075;
  assign n3081 = n887 & ~n3080;
  assign n3082 = ~n884 & n3081;
  assign n3083 = n878 & n3082;
  assign n3084 = ~n3079 & ~n3083;
  assign n3085 = n881 & ~n3084;
  assign n3086 = n3073 & ~n3085;
  assign n3087 = ~pi172 & ~n3086;
  assign n3088 = pi172 & n3086;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = n504 & ~n3089;
  assign n3091 = pi117 & ~pi198;
  assign n3092 = pi109 & pi198;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = ~n504 & ~n3093;
  assign po106 = n3090 | n3094;
  assign n3096 = pi140 & n504;
  assign n3097 = pi118 & ~pi198;
  assign n3098 = pi110 & pi198;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = ~n504 & ~n3099;
  assign po107 = n3096 | n3100;
  assign n3102 = n1614 & n1617;
  assign n3103 = n2484 & n3102;
  assign n3104 = ~n1614 & ~n1617;
  assign n3105 = n2490 & n3104;
  assign n3106 = ~n3103 & ~n3105;
  assign n3107 = ~n1608 & ~n3106;
  assign n3108 = n1608 & n1614;
  assign n3109 = n1617 & n2490;
  assign n3110 = n3108 & n3109;
  assign n3111 = ~n3107 & ~n3110;
  assign n3112 = n1611 & ~n3111;
  assign n3113 = ~n1632 & n2454;
  assign n3114 = ~n2440 & ~n2565;
  assign n3115 = ~n1639 & ~n1648;
  assign n3116 = n3114 & n3115;
  assign n3117 = n3113 & n3116;
  assign n3118 = ~n2441 & ~n2566;
  assign n3119 = ~n1650 & n3118;
  assign n3120 = ~n1656 & ~n1663;
  assign n3121 = ~n1665 & ~n2442;
  assign n3122 = n3120 & n3121;
  assign n3123 = n3119 & n3122;
  assign n3124 = n3117 & n3123;
  assign n3125 = ~n1677 & ~n2445;
  assign n3126 = ~n1670 & n3125;
  assign n3127 = ~n1682 & ~n2567;
  assign n3128 = ~n1689 & ~n2448;
  assign n3129 = n3127 & n3128;
  assign n3130 = n3126 & n3129;
  assign n3131 = ~n1695 & ~n1697;
  assign n3132 = ~n1701 & ~n2568;
  assign n3133 = n3131 & n3132;
  assign n3134 = ~n1705 & ~n2451;
  assign n3135 = ~n1611 & ~n1614;
  assign n3136 = n1608 & n3135;
  assign n3137 = ~n1617 & n2597;
  assign n3138 = n3136 & n3137;
  assign n3139 = ~n2453 & ~n3138;
  assign n3140 = n3134 & n3139;
  assign n3141 = n3133 & n3140;
  assign n3142 = n3130 & n3141;
  assign n3143 = n3124 & n3142;
  assign n3144 = ~n3112 & n3143;
  assign n3145 = ~pi180 & ~n3144;
  assign n3146 = pi180 & n3144;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = n504 & ~n3147;
  assign n3149 = pi119 & ~pi198;
  assign n3150 = pi111 & pi198;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = ~n504 & ~n3151;
  assign po108 = n3148 | n3152;
  assign n3154 = pi148 & n504;
  assign n3155 = pi120 & ~pi198;
  assign n3156 = pi112 & pi198;
  assign n3157 = ~n3155 & ~n3156;
  assign n3158 = ~n504 & ~n3157;
  assign po109 = n3154 | n3158;
  assign n3160 = n2191 & n2225;
  assign n3161 = ~n2188 & n2198;
  assign n3162 = ~n2191 & n3161;
  assign n3163 = n2191 & n2790;
  assign n3164 = ~n2191 & n2785;
  assign n3165 = n2185 & ~n2301;
  assign n3166 = ~n2176 & n3165;
  assign n3167 = n2176 & ~n2182;
  assign n3168 = ~n2185 & ~n2191;
  assign n3169 = n3167 & n3168;
  assign n3170 = ~n3166 & ~n3169;
  assign n3171 = n2188 & ~n3170;
  assign n3172 = n2179 & n3171;
  assign n3173 = n2272 & ~n2775;
  assign n3174 = ~n2776 & ~n3160;
  assign n3175 = ~n2211 & ~n2215;
  assign n3176 = n3174 & n3175;
  assign n3177 = n3173 & n3176;
  assign n3178 = ~n2222 & ~n2779;
  assign n3179 = ~n2221 & n3178;
  assign n3180 = ~n2781 & ~n3162;
  assign n3181 = ~n2226 & ~n2229;
  assign n3182 = n3180 & n3181;
  assign n3183 = n3179 & n3182;
  assign n3184 = n3177 & n3183;
  assign n3185 = ~n2236 & ~n2784;
  assign n3186 = ~n2782 & n3185;
  assign n3187 = ~n2243 & ~n2250;
  assign n3188 = ~n2257 & ~n3163;
  assign n3189 = n3187 & n3188;
  assign n3190 = n3186 & n3189;
  assign n3191 = ~n2262 & ~n2788;
  assign n3192 = ~n2263 & ~n3164;
  assign n3193 = n3191 & n3192;
  assign n3194 = ~n2179 & ~n2182;
  assign n3195 = n2176 & n3194;
  assign n3196 = ~n2188 & n2191;
  assign n3197 = ~n2185 & n3196;
  assign n3198 = n3195 & n3197;
  assign n3199 = ~n2791 & ~n3198;
  assign n3200 = n2293 & n3199;
  assign n3201 = n3193 & n3200;
  assign n3202 = n3190 & n3201;
  assign n3203 = n3184 & n3202;
  assign n3204 = ~n3172 & n3203;
  assign n3205 = ~pi188 & ~n3204;
  assign n3206 = pi188 & n3204;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = n504 & ~n3207;
  assign n3209 = pi113 & pi198;
  assign n3210 = pi121 & ~pi198;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = ~n504 & ~n3211;
  assign po110 = n3208 | n3212;
  assign n3214 = pi156 & n504;
  assign n3215 = pi114 & pi198;
  assign n3216 = pi122 & ~pi198;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = ~n504 & ~n3217;
  assign po111 = n3214 | n3218;
  assign n3220 = ~n2203 & ~n2208;
  assign n3221 = ~n2777 & ~n3160;
  assign n3222 = n3220 & n3221;
  assign n3223 = n2804 & n3222;
  assign n3224 = ~n2779 & ~n3162;
  assign n3225 = ~n2221 & n3224;
  assign n3226 = ~n2224 & ~n2780;
  assign n3227 = ~n2227 & ~n2229;
  assign n3228 = n3226 & n3227;
  assign n3229 = n3225 & n3228;
  assign n3230 = n3223 & n3229;
  assign n3231 = ~n2236 & ~n2240;
  assign n3232 = ~n2782 & n3231;
  assign n3233 = ~n2250 & ~n3163;
  assign n3234 = n2817 & n3233;
  assign n3235 = n3232 & n3234;
  assign n3236 = ~n2262 & ~n2789;
  assign n3237 = ~n2788 & n3236;
  assign n3238 = ~n2266 & ~n3164;
  assign n3239 = n2294 & n3238;
  assign n3240 = n3237 & n3239;
  assign n3241 = n3235 & n3240;
  assign n3242 = n3230 & n3241;
  assign n3243 = n2179 & ~n2191;
  assign n3244 = ~n2179 & n2191;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n2188 & ~n3245;
  assign n3247 = n2182 & n3246;
  assign n3248 = ~n2176 & n3247;
  assign n3249 = ~n2179 & ~n2191;
  assign n3250 = n2179 & n2191;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = n2188 & ~n3251;
  assign n3253 = ~n2182 & n3252;
  assign n3254 = n2176 & n3253;
  assign n3255 = ~n3248 & ~n3254;
  assign n3256 = ~n2185 & ~n3255;
  assign n3257 = n3242 & ~n3256;
  assign n3258 = ~pi163 & ~n3257;
  assign n3259 = pi163 & n3257;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = n504 & ~n3260;
  assign n3262 = pi115 & pi198;
  assign n3263 = pi123 & ~pi198;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = ~n504 & ~n3264;
  assign po112 = n3261 | n3265;
  assign n3267 = pi131 & n504;
  assign n3268 = pi116 & pi198;
  assign n3269 = pi124 & ~pi198;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~n504 & ~n3270;
  assign po113 = n3267 | n3271;
  assign n3273 = n2638 & n2925;
  assign n3274 = ~n2638 & n2663;
  assign n3275 = n2638 & n2713;
  assign n3276 = ~n2638 & n2701;
  assign n3277 = ~n2646 & ~n2918;
  assign n3278 = ~n2643 & n3277;
  assign n3279 = ~n2655 & ~n2922;
  assign n3280 = ~n2664 & ~n3273;
  assign n3281 = n3279 & n3280;
  assign n3282 = n3278 & n3281;
  assign n3283 = ~n2670 & ~n2924;
  assign n3284 = ~n2923 & n3283;
  assign n3285 = ~n2671 & ~n3274;
  assign n3286 = n2726 & n3285;
  assign n3287 = n3284 & n3286;
  assign n3288 = n3282 & n3287;
  assign n3289 = ~n2693 & ~n3275;
  assign n3290 = ~n2697 & ~n2700;
  assign n3291 = n3289 & n3290;
  assign n3292 = n2948 & n3291;
  assign n3293 = ~n2703 & ~n2934;
  assign n3294 = ~n2709 & ~n2935;
  assign n3295 = n3293 & n3294;
  assign n3296 = ~n2712 & ~n2716;
  assign n3297 = n2632 & n2958;
  assign n3298 = ~n2626 & n2629;
  assign n3299 = n2623 & n3298;
  assign n3300 = n3297 & n3299;
  assign n3301 = ~n3276 & ~n3300;
  assign n3302 = n3296 & n3301;
  assign n3303 = n3295 & n3302;
  assign n3304 = n3292 & n3303;
  assign n3305 = n3288 & n3304;
  assign n3306 = ~n2632 & n2968;
  assign n3307 = n2656 & n3306;
  assign n3308 = ~n2632 & ~n2638;
  assign n3309 = n2632 & n2638;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = n2635 & ~n3310;
  assign n3312 = n2626 & n3311;
  assign n3313 = ~n2623 & n3312;
  assign n3314 = ~n3307 & ~n3313;
  assign n3315 = ~n2629 & ~n3314;
  assign n3316 = n3305 & ~n3315;
  assign n3317 = ~pi171 & ~n3316;
  assign n3318 = pi171 & n3316;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = n504 & ~n3319;
  assign n3321 = pi117 & pi198;
  assign n3322 = pi125 & ~pi198;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n504 & ~n3323;
  assign po114 = n3320 | n3324;
  assign n3326 = pi139 & n504;
  assign n3327 = pi118 & pi198;
  assign n3328 = pi126 & ~pi198;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = ~n504 & ~n3329;
  assign po115 = n3326 | n3330;
  assign n3332 = ~n2626 & n2752;
  assign n3333 = ~n2632 & n2638;
  assign n3334 = n2626 & n3333;
  assign n3335 = ~n3332 & ~n3334;
  assign n3336 = n2635 & ~n3335;
  assign n3337 = n2629 & n3336;
  assign n3338 = ~n2623 & n3337;
  assign n3339 = ~n2650 & ~n2655;
  assign n3340 = ~n2646 & n3339;
  assign n3341 = ~n2660 & ~n3273;
  assign n3342 = n2938 & n3341;
  assign n3343 = n3340 & n3342;
  assign n3344 = ~n2666 & ~n2668;
  assign n3345 = ~n2923 & n3344;
  assign n3346 = ~n2671 & ~n2926;
  assign n3347 = ~n2676 & ~n3274;
  assign n3348 = n3346 & n3347;
  assign n3349 = n3345 & n3348;
  assign n3350 = n3343 & n3349;
  assign n3351 = ~n2681 & ~n2685;
  assign n3352 = ~n2928 & n3351;
  assign n3353 = ~n2932 & ~n3275;
  assign n3354 = n2733 & n3353;
  assign n3355 = n3352 & n3354;
  assign n3356 = n2736 & ~n2934;
  assign n3357 = ~n2936 & ~n3276;
  assign n3358 = n2738 & n3357;
  assign n3359 = n3356 & n3358;
  assign n3360 = n3355 & n3359;
  assign n3361 = n3350 & n3360;
  assign n3362 = n2626 & ~n2638;
  assign n3363 = ~n2626 & n2638;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n2635 & ~n3364;
  assign n3366 = n2632 & n3365;
  assign n3367 = ~n2629 & n3366;
  assign n3368 = n2623 & n3367;
  assign n3369 = n3361 & ~n3368;
  assign n3370 = ~n3338 & n3369;
  assign n3371 = ~pi179 & ~n3370;
  assign n3372 = pi179 & n3370;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = n504 & ~n3373;
  assign n3375 = pi119 & pi198;
  assign n3376 = pi127 & ~pi198;
  assign n3377 = ~n3375 & ~n3376;
  assign n3378 = ~n504 & ~n3377;
  assign po116 = n3374 | n3378;
  assign n3380 = pi147 & n504;
  assign n3381 = pi120 & pi198;
  assign n3382 = pi128 & ~pi198;
  assign n3383 = ~n3381 & ~n3382;
  assign n3384 = ~n504 & ~n3383;
  assign po117 = n3380 | n3384;
  assign n3386 = n737 & n2009;
  assign n3387 = ~n737 & n2011;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = ~n743 & ~n3388;
  assign n3390 = n734 & n3389;
  assign n3391 = ~n731 & n3390;
  assign n3392 = n821 & ~n2851;
  assign n3393 = ~n765 & ~n1992;
  assign n3394 = ~n769 & ~n1993;
  assign n3395 = n3393 & n3394;
  assign n3396 = n3392 & n3395;
  assign n3397 = ~n775 & ~n2854;
  assign n3398 = ~n773 & n3397;
  assign n3399 = ~n777 & ~n1994;
  assign n3400 = ~n778 & ~n1998;
  assign n3401 = n3399 & n3400;
  assign n3402 = n3398 & n3401;
  assign n3403 = n3396 & n3402;
  assign n3404 = ~n792 & ~n1999;
  assign n3405 = ~n788 & n3404;
  assign n3406 = ~n809 & ~n2856;
  assign n3407 = n2039 & n3406;
  assign n3408 = n3405 & n3407;
  assign n3409 = ~n815 & ~n2858;
  assign n3410 = ~n812 & n3409;
  assign n3411 = ~n818 & ~n2005;
  assign n3412 = ~n819 & ~n2006;
  assign n3413 = n3411 & n3412;
  assign n3414 = n3410 & n3413;
  assign n3415 = n3408 & n3414;
  assign n3416 = n3403 & n3415;
  assign n3417 = ~n737 & n856;
  assign n3418 = n737 & n857;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = n743 & ~n3419;
  assign n3421 = ~n734 & n3420;
  assign n3422 = n731 & n3421;
  assign n3423 = n3416 & ~n3422;
  assign n3424 = ~n3391 & n3423;
  assign n3425 = ~pi187 & ~n3424;
  assign n3426 = pi187 & n3424;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = n504 & ~n3427;
  assign n3429 = pi129 & ~pi198;
  assign n3430 = pi121 & pi198;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = ~n504 & ~n3431;
  assign po118 = n3428 | n3432;
  assign n3434 = pi155 & n504;
  assign n3435 = pi130 & ~pi198;
  assign n3436 = pi122 & pi198;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = ~n504 & ~n3437;
  assign po119 = n3434 | n3438;
  assign n3440 = ~n504 & ~n3260;
  assign n3441 = pi001 & n504;
  assign po120 = n3440 | n3441;
  assign n3443 = ~n504 & ~n3037;
  assign n3444 = pi060 & n504;
  assign po121 = n3443 | n3444;
  assign n3446 = ~n504 & ~n2761;
  assign n3447 = pi052 & n504;
  assign po122 = n3446 | n3447;
  assign n3449 = ~n504 & ~n2425;
  assign n3450 = pi044 & n504;
  assign po123 = n3449 | n3450;
  assign n3452 = ~n504 & ~n2111;
  assign n3453 = pi036 & n504;
  assign po124 = n3452 | n3453;
  assign n3455 = ~n504 & ~n1751;
  assign n3456 = pi028 & n504;
  assign po125 = n3455 | n3456;
  assign n3458 = ~n504 & ~n1302;
  assign n3459 = pi020 & n504;
  assign po126 = n3458 | n3459;
  assign n3461 = ~n504 & ~n867;
  assign n3462 = pi012 & n504;
  assign po127 = n3461 | n3462;
  assign n3464 = ~n504 & ~n3319;
  assign n3465 = pi003 & n504;
  assign po128 = n3464 | n3465;
  assign n3467 = ~n504 & ~n3089;
  assign n3468 = pi062 & n504;
  assign po129 = n3467 | n3468;
  assign n3470 = ~n504 & ~n2838;
  assign n3471 = pi054 & n504;
  assign po130 = n3470 | n3471;
  assign n3473 = ~n504 & ~n2498;
  assign n3474 = pi046 & n504;
  assign po131 = n3473 | n3474;
  assign n3476 = ~n504 & ~n2161;
  assign n3477 = pi038 & n504;
  assign po132 = n3476 | n3477;
  assign n3479 = ~n504 & ~n1910;
  assign n3480 = pi030 & n504;
  assign po133 = n3479 | n3480;
  assign n3482 = ~n504 & ~n1459;
  assign n3483 = pi022 & n504;
  assign po134 = n3482 | n3483;
  assign n3485 = ~n504 & ~n1017;
  assign n3486 = pi014 & n504;
  assign po135 = n3485 | n3486;
  assign n3488 = ~n504 & ~n3373;
  assign n3489 = pi005 & n504;
  assign po136 = n3488 | n3489;
  assign n3491 = ~n504 & ~n3147;
  assign n3492 = pi064 & n504;
  assign po137 = n3491 | n3492;
  assign n3494 = ~n504 & ~n2904;
  assign n3495 = pi056 & n504;
  assign po138 = n3494 | n3495;
  assign n3497 = ~n504 & ~n2552;
  assign n3498 = pi048 & n504;
  assign po139 = n3497 | n3498;
  assign n3500 = ~n504 & ~n2311;
  assign n3501 = pi040 & n504;
  assign po140 = n3500 | n3501;
  assign n3503 = ~n504 & ~n1976;
  assign n3504 = pi032 & n504;
  assign po141 = n3503 | n3504;
  assign n3506 = ~n504 & ~n1517;
  assign n3507 = pi024 & n504;
  assign po142 = n3506 | n3507;
  assign n3509 = ~n504 & ~n1083;
  assign n3510 = pi016 & n504;
  assign po143 = n3509 | n3510;
  assign n3512 = ~n504 & ~n3427;
  assign n3513 = pi007 & n504;
  assign po144 = n3512 | n3513;
  assign n3515 = ~n504 & ~n3207;
  assign n3516 = pi066 & n504;
  assign po145 = n3515 | n3516;
  assign n3518 = ~n504 & ~n2980;
  assign n3519 = pi058 & n504;
  assign po146 = n3518 | n3519;
  assign n3521 = ~n504 & ~n2608;
  assign n3522 = pi050 & n504;
  assign po147 = n3521 | n3522;
  assign n3524 = ~n504 & ~n2372;
  assign n3525 = pi042 & n504;
  assign po148 = n3524 | n3525;
  assign n3527 = ~n504 & ~n2054;
  assign n3528 = pi034 & n504;
  assign po149 = n3527 | n3528;
  assign n3530 = ~n504 & ~n1593;
  assign n3531 = pi026 & n504;
  assign po150 = n3530 | n3531;
  assign n3533 = ~n504 & ~n1230;
  assign n3534 = pi018 & n504;
  assign po151 = n3533 | n3534;
  assign n3536 = pi131 & ~n504;
  assign n3537 = pi000 & n504;
  assign po152 = n3536 | n3537;
  assign n3539 = pi132 & ~n504;
  assign n3540 = pi059 & n504;
  assign po153 = n3539 | n3540;
  assign n3542 = pi133 & ~n504;
  assign n3543 = pi051 & n504;
  assign po154 = n3542 | n3543;
  assign n3545 = pi134 & ~n504;
  assign n3546 = pi043 & n504;
  assign po155 = n3545 | n3546;
  assign n3548 = pi135 & ~n504;
  assign n3549 = pi035 & n504;
  assign po156 = n3548 | n3549;
  assign n3551 = pi136 & ~n504;
  assign n3552 = pi027 & n504;
  assign po157 = n3551 | n3552;
  assign n3554 = pi137 & ~n504;
  assign n3555 = pi019 & n504;
  assign po158 = n3554 | n3555;
  assign n3557 = pi138 & ~n504;
  assign n3558 = pi011 & n504;
  assign po159 = n3557 | n3558;
  assign n3560 = pi139 & ~n504;
  assign n3561 = pi002 & n504;
  assign po160 = n3560 | n3561;
  assign n3563 = pi140 & ~n504;
  assign n3564 = pi061 & n504;
  assign po161 = n3563 | n3564;
  assign n3566 = pi141 & ~n504;
  assign n3567 = pi053 & n504;
  assign po162 = n3566 | n3567;
  assign n3569 = pi142 & ~n504;
  assign n3570 = pi045 & n504;
  assign po163 = n3569 | n3570;
  assign n3572 = pi143 & ~n504;
  assign n3573 = pi037 & n504;
  assign po164 = n3572 | n3573;
  assign n3575 = pi144 & ~n504;
  assign n3576 = pi029 & n504;
  assign po165 = n3575 | n3576;
  assign n3578 = pi145 & ~n504;
  assign n3579 = pi021 & n504;
  assign po166 = n3578 | n3579;
  assign n3581 = pi146 & ~n504;
  assign n3582 = pi013 & n504;
  assign po167 = n3581 | n3582;
  assign n3584 = pi147 & ~n504;
  assign n3585 = pi004 & n504;
  assign po168 = n3584 | n3585;
  assign n3587 = pi148 & ~n504;
  assign n3588 = pi063 & n504;
  assign po169 = n3587 | n3588;
  assign n3590 = pi149 & ~n504;
  assign n3591 = pi055 & n504;
  assign po170 = n3590 | n3591;
  assign n3593 = pi150 & ~n504;
  assign n3594 = pi047 & n504;
  assign po171 = n3593 | n3594;
  assign n3596 = pi151 & ~n504;
  assign n3597 = pi039 & n504;
  assign po172 = n3596 | n3597;
  assign n3599 = pi152 & ~n504;
  assign n3600 = pi031 & n504;
  assign po173 = n3599 | n3600;
  assign n3602 = pi153 & ~n504;
  assign n3603 = pi023 & n504;
  assign po174 = n3602 | n3603;
  assign n3605 = pi154 & ~n504;
  assign n3606 = pi015 & n504;
  assign po175 = n3605 | n3606;
  assign n3608 = pi155 & ~n504;
  assign n3609 = pi006 & n504;
  assign po176 = n3608 | n3609;
  assign n3611 = pi156 & ~n504;
  assign n3612 = pi065 & n504;
  assign po177 = n3611 | n3612;
  assign n3614 = pi157 & ~n504;
  assign n3615 = pi057 & n504;
  assign po178 = n3614 | n3615;
  assign n3617 = pi158 & ~n504;
  assign n3618 = pi049 & n504;
  assign po179 = n3617 | n3618;
  assign n3620 = pi159 & ~n504;
  assign n3621 = pi041 & n504;
  assign po180 = n3620 | n3621;
  assign n3623 = pi160 & ~n504;
  assign n3624 = pi033 & n504;
  assign po181 = n3623 | n3624;
  assign n3626 = pi161 & ~n504;
  assign n3627 = pi025 & n504;
  assign po182 = n3626 | n3627;
  assign n3629 = pi162 & ~n504;
  assign n3630 = pi017 & n504;
  assign po183 = n3629 | n3630;
  assign n3632 = pi010 & n504;
  assign n3633 = pi195 & ~n503;
  assign n3634 = ~pi195 & pi196;
  assign n3635 = n502 & n3634;
  assign n3636 = ~n3633 & ~n3635;
  assign n3637 = ~pi008 & ~n3636;
  assign po184 = ~n3632 & n3637;
  assign n3639 = pi196 & ~n502;
  assign n3640 = ~pi196 & n502;
  assign n3641 = ~n3639 & ~n3640;
  assign n3642 = ~pi008 & ~n3641;
  assign po185 = ~n3632 & n3642;
  assign n3644 = pi197 & ~pi198;
  assign n3645 = ~pi197 & pi198;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = ~pi008 & ~n3646;
  assign po186 = ~n3632 & n3647;
  assign n3649 = ~pi008 & ~n3632;
  assign po187 = ~pi198 & n3649;
  assign n3651 = ~pi009 & pi255;
  assign n3652 = pi009 & ~pi255;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = pi195 & ~n3653;
  assign n3655 = pi196 & n3654;
  assign n3656 = pi197 & n3655;
  assign n3657 = pi198 & n3656;
  assign n3658 = pi195 & ~pi198;
  assign n3659 = ~pi198 & ~n3658;
  assign n3660 = pi196 & ~n3659;
  assign n3661 = pi197 & n3660;
  assign n3662 = ~pi197 & ~pi198;
  assign n3663 = ~pi195 & ~pi196;
  assign n3664 = n3662 & n3663;
  assign n3665 = ~n3661 & ~n3664;
  assign n3666 = ~pi009 & pi039;
  assign n3667 = pi009 & pi018;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = n3632 & ~n3668;
  assign n3670 = pi226 & ~n3665;
  assign n3671 = pi225 & n3665;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = pi255 & ~n3672;
  assign n3674 = pi200 & ~n3665;
  assign n3675 = pi201 & n3665;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = ~pi255 & ~n3676;
  assign n3678 = ~n3673 & ~n3677;
  assign n3679 = ~n3657 & ~n3678;
  assign n3680 = pi199 & n3657;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = ~n3632 & ~n3681;
  assign n3683 = ~n3669 & ~n3682;
  assign po188 = ~pi008 & ~n3683;
  assign n3685 = pi009 & pi039;
  assign n3686 = ~pi009 & pi031;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = n3632 & ~n3687;
  assign n3689 = pi199 & ~n3665;
  assign n3690 = pi226 & n3665;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = pi255 & ~n3691;
  assign n3693 = pi201 & ~n3665;
  assign n3694 = pi202 & n3665;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = ~pi255 & ~n3695;
  assign n3697 = ~n3692 & ~n3696;
  assign n3698 = ~n3657 & ~n3697;
  assign n3699 = pi200 & n3657;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~n3632 & ~n3700;
  assign n3702 = ~n3688 & ~n3701;
  assign po189 = ~pi008 & ~n3702;
  assign n3704 = pi199 & n3665;
  assign n3705 = ~n3674 & ~n3704;
  assign n3706 = pi255 & ~n3705;
  assign n3707 = pi202 & ~n3665;
  assign n3708 = pi203 & n3665;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = ~pi255 & ~n3709;
  assign n3711 = ~n3706 & ~n3710;
  assign n3712 = ~n3657 & ~n3711;
  assign n3713 = pi201 & n3657;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = ~n3632 & ~n3714;
  assign n3716 = pi009 & pi031;
  assign n3717 = ~pi009 & pi023;
  assign n3718 = ~n3716 & ~n3717;
  assign n3719 = n3632 & ~n3718;
  assign n3720 = ~n3715 & ~n3719;
  assign po190 = ~pi008 & ~n3720;
  assign n3722 = pi200 & n3665;
  assign n3723 = ~n3693 & ~n3722;
  assign n3724 = pi255 & ~n3723;
  assign n3725 = pi203 & ~n3665;
  assign n3726 = pi204 & n3665;
  assign n3727 = ~n3725 & ~n3726;
  assign n3728 = ~pi255 & ~n3727;
  assign n3729 = ~n3724 & ~n3728;
  assign n3730 = ~n3657 & ~n3729;
  assign n3731 = pi202 & n3657;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = ~n3632 & ~n3732;
  assign n3734 = pi009 & pi023;
  assign n3735 = ~pi009 & pi015;
  assign n3736 = ~n3734 & ~n3735;
  assign n3737 = n3632 & ~n3736;
  assign n3738 = ~n3733 & ~n3737;
  assign po191 = ~pi008 & ~n3738;
  assign n3740 = pi005 & ~pi009;
  assign n3741 = pi009 & pi015;
  assign n3742 = ~n3740 & ~n3741;
  assign n3743 = n3632 & ~n3742;
  assign n3744 = ~n3675 & ~n3707;
  assign n3745 = pi255 & ~n3744;
  assign n3746 = pi205 & n3665;
  assign n3747 = pi204 & ~n3665;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = ~pi255 & ~n3748;
  assign n3750 = ~n3745 & ~n3749;
  assign n3751 = ~n3657 & ~n3750;
  assign n3752 = pi203 & n3657;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = ~n3632 & ~n3753;
  assign n3755 = ~n3743 & ~n3754;
  assign po192 = ~pi008 & ~n3755;
  assign n3757 = pi005 & pi009;
  assign n3758 = ~pi009 & pi064;
  assign n3759 = ~n3757 & ~n3758;
  assign n3760 = n3632 & ~n3759;
  assign n3761 = ~n3694 & ~n3725;
  assign n3762 = pi255 & ~n3761;
  assign n3763 = pi206 & n3665;
  assign n3764 = pi205 & ~n3665;
  assign n3765 = ~n3763 & ~n3764;
  assign n3766 = ~pi255 & ~n3765;
  assign n3767 = ~n3762 & ~n3766;
  assign n3768 = ~n3657 & ~n3767;
  assign n3769 = pi204 & n3657;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = ~n3632 & ~n3770;
  assign n3772 = ~n3760 & ~n3771;
  assign po193 = ~pi008 & ~n3772;
  assign n3774 = ~pi009 & pi056;
  assign n3775 = pi009 & pi064;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = n3632 & ~n3776;
  assign n3778 = ~n3708 & ~n3747;
  assign n3779 = pi255 & ~n3778;
  assign n3780 = pi206 & ~n3665;
  assign n3781 = pi207 & n3665;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~pi255 & ~n3782;
  assign n3784 = ~n3779 & ~n3783;
  assign n3785 = ~n3657 & ~n3784;
  assign n3786 = pi205 & n3657;
  assign n3787 = ~n3785 & ~n3786;
  assign n3788 = ~n3632 & ~n3787;
  assign n3789 = ~n3777 & ~n3788;
  assign po194 = ~pi008 & ~n3789;
  assign n3791 = ~n3726 & ~n3764;
  assign n3792 = pi255 & ~n3791;
  assign n3793 = pi207 & ~n3665;
  assign n3794 = pi208 & n3665;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = ~pi255 & ~n3795;
  assign n3797 = ~n3792 & ~n3796;
  assign n3798 = ~n3657 & ~n3797;
  assign n3799 = pi206 & n3657;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = ~n3632 & ~n3800;
  assign n3802 = pi009 & pi056;
  assign n3803 = ~pi009 & pi048;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = n3632 & ~n3804;
  assign n3806 = ~n3801 & ~n3805;
  assign po195 = ~pi008 & ~n3806;
  assign n3808 = ~n3746 & ~n3780;
  assign n3809 = pi255 & ~n3808;
  assign n3810 = pi208 & ~n3665;
  assign n3811 = pi209 & n3665;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~pi255 & ~n3812;
  assign n3814 = ~n3809 & ~n3813;
  assign n3815 = ~n3657 & ~n3814;
  assign n3816 = pi207 & n3657;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n3632 & ~n3817;
  assign n3819 = pi009 & pi048;
  assign n3820 = ~pi009 & pi040;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = n3632 & ~n3821;
  assign n3823 = ~n3818 & ~n3822;
  assign po196 = ~pi008 & ~n3823;
  assign n3825 = ~n3763 & ~n3793;
  assign n3826 = pi255 & ~n3825;
  assign n3827 = pi209 & ~n3665;
  assign n3828 = pi210 & n3665;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = ~pi255 & ~n3829;
  assign n3831 = ~n3826 & ~n3830;
  assign n3832 = ~n3657 & ~n3831;
  assign n3833 = pi208 & n3657;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = ~n3632 & ~n3834;
  assign n3836 = pi009 & pi040;
  assign n3837 = ~pi009 & pi032;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = n3632 & ~n3838;
  assign n3840 = ~n3835 & ~n3839;
  assign po197 = ~pi008 & ~n3840;
  assign n3842 = ~n3781 & ~n3810;
  assign n3843 = pi255 & ~n3842;
  assign n3844 = pi210 & ~n3665;
  assign n3845 = pi211 & n3665;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = ~pi255 & ~n3846;
  assign n3848 = ~n3843 & ~n3847;
  assign n3849 = ~n3657 & ~n3848;
  assign n3850 = pi209 & n3657;
  assign n3851 = ~n3849 & ~n3850;
  assign n3852 = ~n3632 & ~n3851;
  assign n3853 = pi009 & pi032;
  assign n3854 = ~pi009 & pi024;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = n3632 & ~n3855;
  assign n3857 = ~n3852 & ~n3856;
  assign po198 = ~pi008 & ~n3857;
  assign n3859 = ~n3794 & ~n3827;
  assign n3860 = pi255 & ~n3859;
  assign n3861 = pi211 & ~n3665;
  assign n3862 = pi212 & n3665;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~pi255 & ~n3863;
  assign n3865 = ~n3860 & ~n3864;
  assign n3866 = ~n3657 & ~n3865;
  assign n3867 = pi210 & n3657;
  assign n3868 = ~n3866 & ~n3867;
  assign n3869 = ~n3632 & ~n3868;
  assign n3870 = pi009 & pi024;
  assign n3871 = ~pi009 & pi016;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = n3632 & ~n3872;
  assign n3874 = ~n3869 & ~n3873;
  assign po199 = ~pi008 & ~n3874;
  assign n3876 = pi006 & ~pi009;
  assign n3877 = pi009 & pi016;
  assign n3878 = ~n3876 & ~n3877;
  assign n3879 = n3632 & ~n3878;
  assign n3880 = ~n3811 & ~n3844;
  assign n3881 = pi255 & ~n3880;
  assign n3882 = pi213 & n3665;
  assign n3883 = pi212 & ~n3665;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = ~pi255 & ~n3884;
  assign n3886 = ~n3881 & ~n3885;
  assign n3887 = ~n3657 & ~n3886;
  assign n3888 = pi211 & n3657;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = ~n3632 & ~n3889;
  assign n3891 = ~n3879 & ~n3890;
  assign po200 = ~pi008 & ~n3891;
  assign n3893 = pi006 & pi009;
  assign n3894 = ~pi009 & pi065;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = n3632 & ~n3895;
  assign n3897 = ~n3828 & ~n3861;
  assign n3898 = pi255 & ~n3897;
  assign n3899 = pi214 & n3665;
  assign n3900 = pi213 & ~n3665;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = ~pi255 & ~n3901;
  assign n3903 = ~n3898 & ~n3902;
  assign n3904 = ~n3657 & ~n3903;
  assign n3905 = pi212 & n3657;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3632 & ~n3906;
  assign n3908 = ~n3896 & ~n3907;
  assign po201 = ~pi008 & ~n3908;
  assign n3910 = ~n3845 & ~n3883;
  assign n3911 = pi255 & ~n3910;
  assign n3912 = pi214 & ~n3665;
  assign n3913 = pi215 & n3665;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = ~pi255 & ~n3914;
  assign n3916 = ~n3911 & ~n3915;
  assign n3917 = ~n3657 & ~n3916;
  assign n3918 = pi213 & n3657;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n3632 & ~n3919;
  assign n3921 = pi009 & pi065;
  assign n3922 = ~pi009 & pi057;
  assign n3923 = ~n3921 & ~n3922;
  assign n3924 = n3632 & ~n3923;
  assign n3925 = ~n3920 & ~n3924;
  assign po202 = ~pi008 & ~n3925;
  assign n3927 = ~pi009 & pi049;
  assign n3928 = pi009 & pi057;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = n3632 & ~n3929;
  assign n3931 = ~n3862 & ~n3900;
  assign n3932 = pi255 & ~n3931;
  assign n3933 = pi215 & ~n3665;
  assign n3934 = pi216 & n3665;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = ~pi255 & ~n3935;
  assign n3937 = ~n3932 & ~n3936;
  assign n3938 = ~n3657 & ~n3937;
  assign n3939 = pi214 & n3657;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = ~n3632 & ~n3940;
  assign n3942 = ~n3930 & ~n3941;
  assign po203 = ~pi008 & ~n3942;
  assign n3944 = pi009 & pi049;
  assign n3945 = ~pi009 & pi041;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n3632 & ~n3946;
  assign n3948 = ~n3882 & ~n3912;
  assign n3949 = pi255 & ~n3948;
  assign n3950 = pi217 & n3665;
  assign n3951 = pi216 & ~n3665;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = ~pi255 & ~n3952;
  assign n3954 = ~n3949 & ~n3953;
  assign n3955 = ~n3657 & ~n3954;
  assign n3956 = pi215 & n3657;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = ~n3632 & ~n3957;
  assign n3959 = ~n3947 & ~n3958;
  assign po204 = ~pi008 & ~n3959;
  assign n3961 = pi009 & pi041;
  assign n3962 = ~pi009 & pi033;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = n3632 & ~n3963;
  assign n3965 = ~n3899 & ~n3933;
  assign n3966 = pi255 & ~n3965;
  assign n3967 = pi217 & ~n3665;
  assign n3968 = pi218 & n3665;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = ~pi255 & ~n3969;
  assign n3971 = ~n3966 & ~n3970;
  assign n3972 = ~n3657 & ~n3971;
  assign n3973 = pi216 & n3657;
  assign n3974 = ~n3972 & ~n3973;
  assign n3975 = ~n3632 & ~n3974;
  assign n3976 = ~n3964 & ~n3975;
  assign po205 = ~pi008 & ~n3976;
  assign n3978 = pi009 & pi033;
  assign n3979 = ~pi009 & pi025;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = n3632 & ~n3980;
  assign n3982 = ~n3913 & ~n3951;
  assign n3983 = pi255 & ~n3982;
  assign n3984 = pi218 & ~n3665;
  assign n3985 = pi219 & n3665;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = ~pi255 & ~n3986;
  assign n3988 = ~n3983 & ~n3987;
  assign n3989 = ~n3657 & ~n3988;
  assign n3990 = pi217 & n3657;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = ~n3632 & ~n3991;
  assign n3993 = ~n3981 & ~n3992;
  assign po206 = ~pi008 & ~n3993;
  assign n3995 = pi009 & pi025;
  assign n3996 = ~pi009 & pi017;
  assign n3997 = ~n3995 & ~n3996;
  assign n3998 = n3632 & ~n3997;
  assign n3999 = ~n3934 & ~n3967;
  assign n4000 = pi255 & ~n3999;
  assign n4001 = pi219 & ~n3665;
  assign n4002 = pi220 & n3665;
  assign n4003 = ~n4001 & ~n4002;
  assign n4004 = ~pi255 & ~n4003;
  assign n4005 = ~n4000 & ~n4004;
  assign n4006 = ~n3657 & ~n4005;
  assign n4007 = pi218 & n3657;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = ~n3632 & ~n4008;
  assign n4010 = ~n3998 & ~n4009;
  assign po207 = ~pi008 & ~n4010;
  assign n4012 = pi007 & ~pi009;
  assign n4013 = pi009 & pi017;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = n3632 & ~n4014;
  assign n4016 = ~n3950 & ~n3984;
  assign n4017 = pi255 & ~n4016;
  assign n4018 = pi221 & n3665;
  assign n4019 = pi220 & ~n3665;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = ~pi255 & ~n4020;
  assign n4022 = ~n4017 & ~n4021;
  assign n4023 = ~n3657 & ~n4022;
  assign n4024 = pi219 & n3657;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = ~n3632 & ~n4025;
  assign n4027 = ~n4015 & ~n4026;
  assign po208 = ~pi008 & ~n4027;
  assign n4029 = pi007 & pi009;
  assign n4030 = ~pi009 & pi066;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = n3632 & ~n4031;
  assign n4033 = ~n3968 & ~n4001;
  assign n4034 = pi255 & ~n4033;
  assign n4035 = pi222 & n3665;
  assign n4036 = pi221 & ~n3665;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = ~pi255 & ~n4037;
  assign n4039 = ~n4034 & ~n4038;
  assign n4040 = ~n3657 & ~n4039;
  assign n4041 = pi220 & n3657;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = ~n3632 & ~n4042;
  assign n4044 = ~n4032 & ~n4043;
  assign po209 = ~pi008 & ~n4044;
  assign n4046 = ~n3985 & ~n4019;
  assign n4047 = pi255 & ~n4046;
  assign n4048 = pi222 & ~n3665;
  assign n4049 = pi223 & n3665;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = ~pi255 & ~n4050;
  assign n4052 = ~n4047 & ~n4051;
  assign n4053 = ~n3657 & ~n4052;
  assign n4054 = pi221 & n3657;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = ~n3632 & ~n4055;
  assign n4057 = pi009 & pi066;
  assign n4058 = ~pi009 & pi058;
  assign n4059 = ~n4057 & ~n4058;
  assign n4060 = n3632 & ~n4059;
  assign n4061 = ~n4056 & ~n4060;
  assign po210 = ~pi008 & ~n4061;
  assign n4063 = ~pi009 & pi050;
  assign n4064 = pi009 & pi058;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = n3632 & ~n4065;
  assign n4067 = ~n4002 & ~n4036;
  assign n4068 = pi255 & ~n4067;
  assign n4069 = pi223 & ~n3665;
  assign n4070 = pi224 & n3665;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = ~pi255 & ~n4071;
  assign n4073 = ~n4068 & ~n4072;
  assign n4074 = ~n3657 & ~n4073;
  assign n4075 = pi222 & n3657;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~n3632 & ~n4076;
  assign n4078 = ~n4066 & ~n4077;
  assign po211 = ~pi008 & ~n4078;
  assign n4080 = ~n4018 & ~n4048;
  assign n4081 = pi255 & ~n4080;
  assign n4082 = pi224 & ~n3665;
  assign n4083 = ~n3671 & ~n4082;
  assign n4084 = ~pi255 & ~n4083;
  assign n4085 = ~n4081 & ~n4084;
  assign n4086 = ~n3657 & ~n4085;
  assign n4087 = pi223 & n3657;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = ~n3632 & ~n4088;
  assign n4090 = pi009 & pi050;
  assign n4091 = ~pi009 & pi042;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = n3632 & ~n4092;
  assign n4094 = ~n4089 & ~n4093;
  assign po212 = ~pi008 & ~n4094;
  assign n4096 = ~n4035 & ~n4069;
  assign n4097 = pi255 & ~n4096;
  assign n4098 = pi225 & ~n3665;
  assign n4099 = ~n3690 & ~n4098;
  assign n4100 = ~pi255 & ~n4099;
  assign n4101 = ~n4097 & ~n4100;
  assign n4102 = ~n3657 & ~n4101;
  assign n4103 = pi224 & n3657;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n3632 & ~n4104;
  assign n4106 = pi009 & pi042;
  assign n4107 = ~pi009 & pi034;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = n3632 & ~n4108;
  assign n4110 = ~n4105 & ~n4109;
  assign po213 = ~pi008 & ~n4110;
  assign n4112 = pi009 & pi034;
  assign n4113 = ~pi009 & pi026;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = n3632 & ~n4114;
  assign n4116 = pi225 & n3657;
  assign n4117 = ~n4049 & ~n4082;
  assign n4118 = pi255 & ~n4117;
  assign n4119 = ~n3670 & ~n3704;
  assign n4120 = ~pi255 & ~n4119;
  assign n4121 = ~n4118 & ~n4120;
  assign n4122 = ~n3657 & ~n4121;
  assign n4123 = ~n4116 & ~n4122;
  assign n4124 = ~n3632 & ~n4123;
  assign n4125 = ~n4115 & ~n4124;
  assign po214 = ~pi008 & ~n4125;
  assign n4127 = pi009 & pi026;
  assign n4128 = ~pi009 & pi018;
  assign n4129 = ~n4127 & ~n4128;
  assign n4130 = n3632 & ~n4129;
  assign n4131 = pi226 & n3657;
  assign n4132 = ~n3689 & ~n3722;
  assign n4133 = ~pi255 & ~n4132;
  assign n4134 = ~n4070 & ~n4098;
  assign n4135 = pi255 & ~n4134;
  assign n4136 = ~n4133 & ~n4135;
  assign n4137 = ~n3657 & ~n4136;
  assign n4138 = ~n4131 & ~n4137;
  assign n4139 = ~n3632 & ~n4138;
  assign n4140 = ~n4130 & ~n4139;
  assign po215 = ~pi008 & ~n4140;
  assign n4142 = pi004 & ~pi009;
  assign n4143 = pi009 & pi012;
  assign n4144 = ~n4142 & ~n4143;
  assign n4145 = n3632 & ~n4144;
  assign n4146 = pi254 & ~n3665;
  assign n4147 = pi253 & n3665;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = pi255 & ~n4148;
  assign n4150 = pi228 & ~n3665;
  assign n4151 = pi229 & n3665;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = ~pi255 & ~n4152;
  assign n4154 = ~n4149 & ~n4153;
  assign n4155 = ~n3657 & ~n4154;
  assign n4156 = pi227 & n3657;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n3632 & ~n4157;
  assign n4159 = ~n4145 & ~n4158;
  assign po216 = ~pi008 & ~n4159;
  assign n4161 = pi004 & pi009;
  assign n4162 = ~pi009 & pi063;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = n3632 & ~n4163;
  assign n4165 = pi227 & ~n3665;
  assign n4166 = pi254 & n3665;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = pi255 & ~n4167;
  assign n4169 = pi230 & n3665;
  assign n4170 = pi229 & ~n3665;
  assign n4171 = ~n4169 & ~n4170;
  assign n4172 = ~pi255 & ~n4171;
  assign n4173 = ~n4168 & ~n4172;
  assign n4174 = ~n3657 & ~n4173;
  assign n4175 = pi228 & n3657;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = ~n3632 & ~n4176;
  assign n4178 = ~n4164 & ~n4177;
  assign po217 = ~pi008 & ~n4178;
  assign n4180 = ~pi009 & pi055;
  assign n4181 = pi009 & pi063;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = n3632 & ~n4182;
  assign n4184 = pi227 & n3665;
  assign n4185 = ~n4150 & ~n4184;
  assign n4186 = pi255 & ~n4185;
  assign n4187 = pi230 & ~n3665;
  assign n4188 = pi231 & n3665;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~pi255 & ~n4189;
  assign n4191 = ~n4186 & ~n4190;
  assign n4192 = ~n3657 & ~n4191;
  assign n4193 = pi229 & n3657;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n3632 & ~n4194;
  assign n4196 = ~n4183 & ~n4195;
  assign po218 = ~pi008 & ~n4196;
  assign n4198 = pi228 & n3665;
  assign n4199 = ~n4170 & ~n4198;
  assign n4200 = pi255 & ~n4199;
  assign n4201 = pi231 & ~n3665;
  assign n4202 = pi232 & n3665;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = ~pi255 & ~n4203;
  assign n4205 = ~n4200 & ~n4204;
  assign n4206 = ~n3657 & ~n4205;
  assign n4207 = pi230 & n3657;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = ~n3632 & ~n4208;
  assign n4210 = pi009 & pi055;
  assign n4211 = ~pi009 & pi047;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = n3632 & ~n4212;
  assign n4214 = ~n4209 & ~n4213;
  assign po219 = ~pi008 & ~n4214;
  assign n4216 = pi003 & ~pi009;
  assign n4217 = pi009 & pi047;
  assign n4218 = ~n4216 & ~n4217;
  assign n4219 = n3632 & ~n4218;
  assign n4220 = ~n4151 & ~n4187;
  assign n4221 = pi255 & ~n4220;
  assign n4222 = pi233 & n3665;
  assign n4223 = pi232 & ~n3665;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~pi255 & ~n4224;
  assign n4226 = ~n4221 & ~n4225;
  assign n4227 = ~n3657 & ~n4226;
  assign n4228 = pi231 & n3657;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n3632 & ~n4229;
  assign n4231 = ~n4219 & ~n4230;
  assign po220 = ~pi008 & ~n4231;
  assign n4233 = pi003 & pi009;
  assign n4234 = ~pi009 & pi062;
  assign n4235 = ~n4233 & ~n4234;
  assign n4236 = n3632 & ~n4235;
  assign n4237 = ~n4169 & ~n4201;
  assign n4238 = pi255 & ~n4237;
  assign n4239 = pi234 & n3665;
  assign n4240 = pi233 & ~n3665;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = ~pi255 & ~n4241;
  assign n4243 = ~n4238 & ~n4242;
  assign n4244 = ~n3657 & ~n4243;
  assign n4245 = pi232 & n3657;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n3632 & ~n4246;
  assign n4248 = ~n4236 & ~n4247;
  assign po221 = ~pi008 & ~n4248;
  assign n4250 = ~pi009 & pi054;
  assign n4251 = pi009 & pi062;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = n3632 & ~n4252;
  assign n4254 = ~n4188 & ~n4223;
  assign n4255 = pi255 & ~n4254;
  assign n4256 = pi234 & ~n3665;
  assign n4257 = pi235 & n3665;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = ~pi255 & ~n4258;
  assign n4260 = ~n4255 & ~n4259;
  assign n4261 = ~n3657 & ~n4260;
  assign n4262 = pi233 & n3657;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = ~n3632 & ~n4263;
  assign n4265 = ~n4253 & ~n4264;
  assign po222 = ~pi008 & ~n4265;
  assign n4267 = ~n4202 & ~n4240;
  assign n4268 = pi255 & ~n4267;
  assign n4269 = pi235 & ~n3665;
  assign n4270 = pi236 & n3665;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~pi255 & ~n4271;
  assign n4273 = ~n4268 & ~n4272;
  assign n4274 = ~n3657 & ~n4273;
  assign n4275 = pi234 & n3657;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~n3632 & ~n4276;
  assign n4278 = pi009 & pi054;
  assign n4279 = ~pi009 & pi046;
  assign n4280 = ~n4278 & ~n4279;
  assign n4281 = n3632 & ~n4280;
  assign n4282 = ~n4277 & ~n4281;
  assign po223 = ~pi008 & ~n4282;
  assign n4284 = ~n4222 & ~n4256;
  assign n4285 = pi255 & ~n4284;
  assign n4286 = pi236 & ~n3665;
  assign n4287 = pi237 & n3665;
  assign n4288 = ~n4286 & ~n4287;
  assign n4289 = ~pi255 & ~n4288;
  assign n4290 = ~n4285 & ~n4289;
  assign n4291 = ~n3657 & ~n4290;
  assign n4292 = pi235 & n3657;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = ~n3632 & ~n4293;
  assign n4295 = pi009 & pi046;
  assign n4296 = ~pi009 & pi038;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = n3632 & ~n4297;
  assign n4299 = ~n4294 & ~n4298;
  assign po224 = ~pi008 & ~n4299;
  assign n4301 = ~n4239 & ~n4269;
  assign n4302 = pi255 & ~n4301;
  assign n4303 = pi237 & ~n3665;
  assign n4304 = pi238 & n3665;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = ~pi255 & ~n4305;
  assign n4307 = ~n4302 & ~n4306;
  assign n4308 = ~n3657 & ~n4307;
  assign n4309 = pi236 & n3657;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = ~n3632 & ~n4310;
  assign n4312 = pi009 & pi038;
  assign n4313 = ~pi009 & pi030;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = n3632 & ~n4314;
  assign n4316 = ~n4311 & ~n4315;
  assign po225 = ~pi008 & ~n4316;
  assign n4318 = ~n4257 & ~n4286;
  assign n4319 = pi255 & ~n4318;
  assign n4320 = pi238 & ~n3665;
  assign n4321 = pi239 & n3665;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = ~pi255 & ~n4322;
  assign n4324 = ~n4319 & ~n4323;
  assign n4325 = ~n3657 & ~n4324;
  assign n4326 = pi237 & n3657;
  assign n4327 = ~n4325 & ~n4326;
  assign n4328 = ~n3632 & ~n4327;
  assign n4329 = pi009 & pi030;
  assign n4330 = ~pi009 & pi022;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = n3632 & ~n4331;
  assign n4333 = ~n4328 & ~n4332;
  assign po226 = ~pi008 & ~n4333;
  assign n4335 = ~n4270 & ~n4303;
  assign n4336 = pi255 & ~n4335;
  assign n4337 = pi239 & ~n3665;
  assign n4338 = pi240 & n3665;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = ~pi255 & ~n4339;
  assign n4341 = ~n4336 & ~n4340;
  assign n4342 = ~n3657 & ~n4341;
  assign n4343 = pi238 & n3657;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = ~n3632 & ~n4344;
  assign n4346 = pi009 & pi022;
  assign n4347 = ~pi009 & pi014;
  assign n4348 = ~n4346 & ~n4347;
  assign n4349 = n3632 & ~n4348;
  assign n4350 = ~n4345 & ~n4349;
  assign po227 = ~pi008 & ~n4350;
  assign n4352 = pi002 & ~pi009;
  assign n4353 = pi009 & pi014;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = n3632 & ~n4354;
  assign n4356 = ~n4287 & ~n4320;
  assign n4357 = pi255 & ~n4356;
  assign n4358 = pi241 & n3665;
  assign n4359 = pi240 & ~n3665;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~pi255 & ~n4360;
  assign n4362 = ~n4357 & ~n4361;
  assign n4363 = ~n3657 & ~n4362;
  assign n4364 = pi239 & n3657;
  assign n4365 = ~n4363 & ~n4364;
  assign n4366 = ~n3632 & ~n4365;
  assign n4367 = ~n4355 & ~n4366;
  assign po228 = ~pi008 & ~n4367;
  assign n4369 = pi002 & pi009;
  assign n4370 = ~pi009 & pi061;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = n3632 & ~n4371;
  assign n4373 = ~n4304 & ~n4337;
  assign n4374 = pi255 & ~n4373;
  assign n4375 = pi242 & n3665;
  assign n4376 = pi241 & ~n3665;
  assign n4377 = ~n4375 & ~n4376;
  assign n4378 = ~pi255 & ~n4377;
  assign n4379 = ~n4374 & ~n4378;
  assign n4380 = ~n3657 & ~n4379;
  assign n4381 = pi240 & n3657;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = ~n3632 & ~n4382;
  assign n4384 = ~n4372 & ~n4383;
  assign po229 = ~pi008 & ~n4384;
  assign n4386 = ~pi009 & pi053;
  assign n4387 = pi009 & pi061;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = n3632 & ~n4388;
  assign n4390 = ~n4321 & ~n4359;
  assign n4391 = pi255 & ~n4390;
  assign n4392 = pi242 & ~n3665;
  assign n4393 = pi243 & n3665;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = ~pi255 & ~n4394;
  assign n4396 = ~n4391 & ~n4395;
  assign n4397 = ~n3657 & ~n4396;
  assign n4398 = pi241 & n3657;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n3632 & ~n4399;
  assign n4401 = ~n4389 & ~n4400;
  assign po230 = ~pi008 & ~n4401;
  assign n4403 = ~n4338 & ~n4376;
  assign n4404 = pi255 & ~n4403;
  assign n4405 = pi243 & ~n3665;
  assign n4406 = pi244 & n3665;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = ~pi255 & ~n4407;
  assign n4409 = ~n4404 & ~n4408;
  assign n4410 = ~n3657 & ~n4409;
  assign n4411 = pi242 & n3657;
  assign n4412 = ~n4410 & ~n4411;
  assign n4413 = ~n3632 & ~n4412;
  assign n4414 = pi009 & pi053;
  assign n4415 = ~pi009 & pi045;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = n3632 & ~n4416;
  assign n4418 = ~n4413 & ~n4417;
  assign po231 = ~pi008 & ~n4418;
  assign n4420 = pi009 & pi045;
  assign n4421 = ~pi009 & pi037;
  assign n4422 = ~n4420 & ~n4421;
  assign n4423 = n3632 & ~n4422;
  assign n4424 = ~n4358 & ~n4392;
  assign n4425 = pi255 & ~n4424;
  assign n4426 = pi245 & n3665;
  assign n4427 = pi244 & ~n3665;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = ~pi255 & ~n4428;
  assign n4430 = ~n4425 & ~n4429;
  assign n4431 = ~n3657 & ~n4430;
  assign n4432 = pi243 & n3657;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = ~n3632 & ~n4433;
  assign n4435 = ~n4423 & ~n4434;
  assign po232 = ~pi008 & ~n4435;
  assign n4437 = pi009 & pi037;
  assign n4438 = ~pi009 & pi029;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = n3632 & ~n4439;
  assign n4441 = ~n4375 & ~n4405;
  assign n4442 = pi255 & ~n4441;
  assign n4443 = pi245 & ~n3665;
  assign n4444 = pi246 & n3665;
  assign n4445 = ~n4443 & ~n4444;
  assign n4446 = ~pi255 & ~n4445;
  assign n4447 = ~n4442 & ~n4446;
  assign n4448 = ~n3657 & ~n4447;
  assign n4449 = pi244 & n3657;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = ~n3632 & ~n4450;
  assign n4452 = ~n4440 & ~n4451;
  assign po233 = ~pi008 & ~n4452;
  assign n4454 = pi009 & pi029;
  assign n4455 = ~pi009 & pi021;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = n3632 & ~n4456;
  assign n4458 = ~n4393 & ~n4427;
  assign n4459 = pi255 & ~n4458;
  assign n4460 = pi246 & ~n3665;
  assign n4461 = pi247 & n3665;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = ~pi255 & ~n4462;
  assign n4464 = ~n4459 & ~n4463;
  assign n4465 = ~n3657 & ~n4464;
  assign n4466 = pi245 & n3657;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = ~n3632 & ~n4467;
  assign n4469 = ~n4457 & ~n4468;
  assign po234 = ~pi008 & ~n4469;
  assign n4471 = pi009 & pi021;
  assign n4472 = ~pi009 & pi013;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = n3632 & ~n4473;
  assign n4475 = ~n4406 & ~n4443;
  assign n4476 = pi255 & ~n4475;
  assign n4477 = pi247 & ~n3665;
  assign n4478 = pi248 & n3665;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = ~pi255 & ~n4479;
  assign n4481 = ~n4476 & ~n4480;
  assign n4482 = ~n3657 & ~n4481;
  assign n4483 = pi246 & n3657;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~n3632 & ~n4484;
  assign n4486 = ~n4474 & ~n4485;
  assign po235 = ~pi008 & ~n4486;
  assign n4488 = pi001 & ~pi009;
  assign n4489 = pi009 & pi013;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = n3632 & ~n4490;
  assign n4492 = ~n4426 & ~n4460;
  assign n4493 = pi255 & ~n4492;
  assign n4494 = pi249 & n3665;
  assign n4495 = pi248 & ~n3665;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = ~pi255 & ~n4496;
  assign n4498 = ~n4493 & ~n4497;
  assign n4499 = ~n3657 & ~n4498;
  assign n4500 = pi247 & n3657;
  assign n4501 = ~n4499 & ~n4500;
  assign n4502 = ~n3632 & ~n4501;
  assign n4503 = ~n4491 & ~n4502;
  assign po236 = ~pi008 & ~n4503;
  assign n4505 = pi001 & pi009;
  assign n4506 = ~pi009 & pi060;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = n3632 & ~n4507;
  assign n4509 = ~n4444 & ~n4477;
  assign n4510 = pi255 & ~n4509;
  assign n4511 = pi250 & n3665;
  assign n4512 = pi249 & ~n3665;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = ~pi255 & ~n4513;
  assign n4515 = ~n4510 & ~n4514;
  assign n4516 = ~n3657 & ~n4515;
  assign n4517 = pi248 & n3657;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = ~n3632 & ~n4518;
  assign n4520 = ~n4508 & ~n4519;
  assign po237 = ~pi008 & ~n4520;
  assign n4522 = ~pi009 & pi052;
  assign n4523 = pi009 & pi060;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n3632 & ~n4524;
  assign n4526 = ~n4461 & ~n4495;
  assign n4527 = pi255 & ~n4526;
  assign n4528 = pi250 & ~n3665;
  assign n4529 = pi251 & n3665;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = ~pi255 & ~n4530;
  assign n4532 = ~n4527 & ~n4531;
  assign n4533 = ~n3657 & ~n4532;
  assign n4534 = pi249 & n3657;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = ~n3632 & ~n4535;
  assign n4537 = ~n4525 & ~n4536;
  assign po238 = ~pi008 & ~n4537;
  assign n4539 = ~n4478 & ~n4512;
  assign n4540 = pi255 & ~n4539;
  assign n4541 = pi251 & ~n3665;
  assign n4542 = pi252 & n3665;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = ~pi255 & ~n4543;
  assign n4545 = ~n4540 & ~n4544;
  assign n4546 = ~n3657 & ~n4545;
  assign n4547 = pi250 & n3657;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n3632 & ~n4548;
  assign n4550 = pi009 & pi052;
  assign n4551 = ~pi009 & pi044;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = n3632 & ~n4552;
  assign n4554 = ~n4549 & ~n4553;
  assign po239 = ~pi008 & ~n4554;
  assign n4556 = ~n4494 & ~n4528;
  assign n4557 = pi255 & ~n4556;
  assign n4558 = pi252 & ~n3665;
  assign n4559 = ~n4147 & ~n4558;
  assign n4560 = ~pi255 & ~n4559;
  assign n4561 = ~n4557 & ~n4560;
  assign n4562 = ~n3657 & ~n4561;
  assign n4563 = pi251 & n3657;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = ~n3632 & ~n4564;
  assign n4566 = pi009 & pi044;
  assign n4567 = ~pi009 & pi036;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = n3632 & ~n4568;
  assign n4570 = ~n4565 & ~n4569;
  assign po240 = ~pi008 & ~n4570;
  assign n4572 = ~n4511 & ~n4541;
  assign n4573 = pi255 & ~n4572;
  assign n4574 = pi253 & ~n3665;
  assign n4575 = ~n4166 & ~n4574;
  assign n4576 = ~pi255 & ~n4575;
  assign n4577 = ~n4573 & ~n4576;
  assign n4578 = ~n3657 & ~n4577;
  assign n4579 = pi252 & n3657;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~n3632 & ~n4580;
  assign n4582 = pi009 & pi036;
  assign n4583 = ~pi009 & pi028;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = n3632 & ~n4584;
  assign n4586 = ~n4581 & ~n4585;
  assign po241 = ~pi008 & ~n4586;
  assign n4588 = pi009 & pi028;
  assign n4589 = ~pi009 & pi020;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = n3632 & ~n4590;
  assign n4592 = pi253 & n3657;
  assign n4593 = ~n4529 & ~n4558;
  assign n4594 = pi255 & ~n4593;
  assign n4595 = ~n4146 & ~n4184;
  assign n4596 = ~pi255 & ~n4595;
  assign n4597 = ~n4594 & ~n4596;
  assign n4598 = ~n3657 & ~n4597;
  assign n4599 = ~n4592 & ~n4598;
  assign n4600 = ~n3632 & ~n4599;
  assign n4601 = ~n4591 & ~n4600;
  assign po242 = ~pi008 & ~n4601;
  assign n4603 = pi009 & pi020;
  assign n4604 = ~pi009 & pi012;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = n3632 & ~n4605;
  assign n4607 = pi254 & n3657;
  assign n4608 = ~n4165 & ~n4198;
  assign n4609 = ~pi255 & ~n4608;
  assign n4610 = ~n4542 & ~n4574;
  assign n4611 = pi255 & ~n4610;
  assign n4612 = ~n4609 & ~n4611;
  assign n4613 = ~n3657 & ~n4612;
  assign n4614 = ~n4607 & ~n4613;
  assign n4615 = ~n3632 & ~n4614;
  assign n4616 = ~n4606 & ~n4615;
  assign po243 = ~pi008 & ~n4616;
  assign n4618 = pi195 & pi196;
  assign n4619 = n502 & n4618;
  assign n4620 = pi255 & ~n4619;
  assign n4621 = pi197 & n4618;
  assign n4622 = pi009 & pi198;
  assign n4623 = n4621 & n4622;
  assign po244 = n4620 | n4623;
endmodule



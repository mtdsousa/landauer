// Benchmark "rot" written by ABC on Sun Apr 22 21:43:12 2018

module rot ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106;
  wire n243, n244, n245, n247, n248, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n276, n277, n278, n279, n280, n281,
    n283, n284, n285, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n369, n370,
    n371, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n402, n403, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n441, n442, n443, n445, n446, n447, n448,
    n449, n451, n452, n453, n454, n455, n456, n457, n459, n462, n463, n465,
    n466, n467, n468, n470, n471, n472, n473, n474, n476, n478, n479, n481,
    n483, n484, n486, n488, n490, n491, n493, n495, n496, n497, n499, n501,
    n502, n503, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n575,
    n576, n577, n578, n579, n580, n581, n583, n584, n585, n587, n588, n590,
    n591, n592, n593, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n607, n608, n610, n611, n613, n614, n616, n617, n618, n620, n621,
    n623, n624, n626, n627, n629, n630, n632, n633, n634, n635, n636, n638,
    n639, n640, n641, n642, n645, n646, n647, n650, n651, n652, n654, n655,
    n656, n657, n659, n660, n661, n662, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n688, n689, n690, n691, n692, n694, n695, n696,
    n697, n698, n700, n701, n702, n704, n709, n710, n711, n712, n713, n714,
    n715, n717, n718, n719, n720, n721, n723, n724, n725, n727, n729, n730,
    n731, n732, n733, n734, n736, n737, n738, n739, n740, n745, n746, n747,
    n749, n752, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n771, n772, n773, n775, n777, n778,
    n779, n782, n783, n786, n787, n789, n791;
  assign n243 = pi023 & ~pi024;
  assign n244 = pi030 & ~n243;
  assign n245 = pi061 & n243;
  assign po000 = n244 | n245;
  assign n247 = pi041 & ~pi076;
  assign n248 = pi062 & pi076;
  assign po001 = n247 | n248;
  assign n250 = pi075 & pi090;
  assign n251 = pi076 & n250;
  assign n252 = ~pi020 & pi044;
  assign n253 = ~pi033 & ~pi044;
  assign n254 = ~n252 & ~n253;
  assign n255 = ~pi010 & pi029;
  assign n256 = ~pi012 & ~pi029;
  assign n257 = ~n255 & ~n256;
  assign n258 = pi101 & ~n257;
  assign n259 = ~pi100 & n258;
  assign n260 = ~pi007 & pi124;
  assign n261 = ~n259 & ~n260;
  assign n262 = ~n254 & ~n261;
  assign n263 = pi098 & n262;
  assign n264 = ~pi008 & pi124;
  assign n265 = pi006 & ~n264;
  assign n266 = ~pi009 & pi029;
  assign n267 = ~pi011 & ~pi029;
  assign n268 = ~n266 & ~n267;
  assign n269 = n265 & n268;
  assign n270 = ~n263 & n269;
  assign n271 = pi101 & ~n251;
  assign n272 = pi101 & ~n270;
  assign n273 = pi100 & ~n272;
  assign po102 = n271 | n273;
  assign po002 = pi099 | po102;
  assign n276 = pi020 & pi044;
  assign n277 = ~pi019 & n276;
  assign n278 = pi033 & ~pi044;
  assign n279 = ~pi032 & n278;
  assign n280 = ~n277 & ~n279;
  assign n281 = pi098 & ~n280;
  assign po003 = po102 | n281;
  assign n283 = ~n276 & ~n278;
  assign n284 = pi098 & ~n283;
  assign n285 = pi080 & po102;
  assign po004 = n284 | n285;
  assign n287 = pi093 & pi094;
  assign n288 = pi090 & ~n287;
  assign n289 = ~pi076 & n288;
  assign n290 = pi075 & n289;
  assign n291 = pi043 & n290;
  assign n292 = ~pi075 & pi076;
  assign n293 = pi090 & n292;
  assign n294 = pi055 & pi056;
  assign n295 = pi054 & n294;
  assign n296 = pi013 & ~n295;
  assign n297 = n293 & ~n296;
  assign n298 = ~pi074 & n251;
  assign n299 = ~n291 & ~n298;
  assign po008 = n297 | ~n299;
  assign po009 = pi074 & n251;
  assign n302 = pi079 & ~po102;
  assign n303 = ~pi070 & n302;
  assign n304 = pi044 & ~n303;
  assign n305 = ~pi069 & pi070;
  assign n306 = n302 & n305;
  assign n307 = pi065 & ~n306;
  assign n308 = pi083 & ~pi085;
  assign n309 = ~pi083 & pi085;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~pi084 & ~n310;
  assign n312 = ~pi083 & ~pi085;
  assign n313 = pi069 & ~pi070;
  assign n314 = ~n305 & ~n313;
  assign n315 = pi089 & n311;
  assign n316 = ~pi077 & ~n315;
  assign n317 = ~n314 & ~n316;
  assign n318 = ~n312 & n317;
  assign n319 = pi092 & n318;
  assign n320 = ~pi067 & n319;
  assign n321 = pi069 & n320;
  assign n322 = pi073 & pi079;
  assign n323 = ~po102 & n322;
  assign n324 = ~pi112 & pi116;
  assign n325 = pi111 & n324;
  assign n326 = ~pi108 & ~n325;
  assign n327 = ~n323 & ~n326;
  assign n328 = pi112 & pi116;
  assign n329 = ~pi111 & n328;
  assign n330 = ~pi109 & ~n329;
  assign n331 = ~n323 & ~n330;
  assign n332 = ~n327 & ~n331;
  assign n333 = pi110 & ~n323;
  assign n334 = ~n321 & n333;
  assign n335 = ~n332 & n334;
  assign n336 = ~pi018 & ~pi115;
  assign n337 = ~n304 & ~n336;
  assign n338 = pi098 & ~n337;
  assign n339 = pi128 & ~n307;
  assign n340 = pi099 & ~n339;
  assign n341 = pi102 & ~n321;
  assign n342 = ~n332 & n335;
  assign n343 = n341 & n342;
  assign n344 = ~n340 & ~n343;
  assign n345 = ~n338 & n344;
  assign n346 = ~pi129 & ~n345;
  assign n347 = ~po102 & n346;
  assign n348 = n251 & n270;
  assign n349 = pi101 & ~n348;
  assign n350 = pi100 & ~n349;
  assign n351 = ~n347 & ~n350;
  assign n352 = pi000 & pi031;
  assign n353 = ~po004 & n320;
  assign n354 = ~n352 & ~n353;
  assign n355 = pi095 & n354;
  assign n356 = n351 & ~n355;
  assign n357 = ~pi071 & pi097;
  assign n358 = pi083 & pi085;
  assign n359 = ~pi084 & pi089;
  assign n360 = ~pi077 & ~n359;
  assign n361 = ~n358 & ~n360;
  assign n362 = pi084 & pi089;
  assign n363 = pi077 & ~n362;
  assign n364 = ~n312 & ~n363;
  assign n365 = ~n361 & n364;
  assign n366 = ~n357 & ~n365;
  assign n367 = ~n356 & n366;
  assign po010 = ~pi000 & n367;
  assign n369 = ~pi000 & ~pi071;
  assign n370 = n312 & n369;
  assign n371 = ~pi052 & ~n370;
  assign po011 = pi097 & ~n371;
  assign n373 = pi000 & ~pi085;
  assign n374 = ~pi069 & ~pi070;
  assign n375 = ~pi068 & n374;
  assign n376 = n373 & n375;
  assign n377 = ~pi014 & pi085;
  assign n378 = ~pi015 & ~pi016;
  assign n379 = n377 & n378;
  assign n380 = ~n376 & ~n379;
  assign n381 = ~pi040 & n380;
  assign n382 = ~pi089 & ~n381;
  assign n383 = ~pi057 & ~pi058;
  assign n384 = ~pi059 & pi084;
  assign n385 = n383 & n384;
  assign n386 = ~pi068 & ~pi069;
  assign n387 = ~pi070 & ~pi084;
  assign n388 = n386 & n387;
  assign n389 = ~n385 & ~n388;
  assign n390 = ~pi040 & ~n379;
  assign n391 = ~n389 & ~n390;
  assign n392 = pi084 & ~n385;
  assign n393 = ~pi070 & ~n392;
  assign n394 = ~pi069 & n393;
  assign n395 = ~pi068 & n394;
  assign n396 = ~pi085 & n395;
  assign n397 = ~n391 & ~n396;
  assign n398 = pi000 & ~n397;
  assign n399 = ~n311 & n391;
  assign n400 = ~n398 & ~n399;
  assign po012 = n382 | ~n400;
  assign n402 = po004 & n320;
  assign n403 = ~pi031 & ~n402;
  assign po013 = ~pi000 & ~n403;
  assign n405 = ~n351 & ~n355;
  assign n406 = pi004 & pi005;
  assign n407 = pi003 & n406;
  assign n408 = ~pi069 & ~n407;
  assign n409 = pi013 & pi070;
  assign n410 = n408 & n409;
  assign n411 = pi000 & ~n410;
  assign n412 = ~pi091 & ~pi092;
  assign n413 = n411 & ~n412;
  assign n414 = ~pi091 & n413;
  assign n415 = pi091 & ~n413;
  assign n416 = ~n414 & ~n415;
  assign n417 = ~n405 & ~n416;
  assign n418 = pi021 & pi044;
  assign n419 = pi034 & ~pi044;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~po002 & n420;
  assign n422 = ~po003 & ~n421;
  assign n423 = ~po002 & po003;
  assign n424 = pi102 & ~n332;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~n422 & n425;
  assign n427 = n405 & ~n426;
  assign po014 = n417 | n427;
  assign n429 = pi092 & ~n414;
  assign n430 = ~pi092 & n413;
  assign n431 = ~pi091 & n430;
  assign n432 = ~n429 & ~n431;
  assign n433 = ~n405 & ~n432;
  assign n434 = po002 & ~po003;
  assign n435 = n327 & n331;
  assign n436 = pi102 & n435;
  assign n437 = ~n423 & ~n436;
  assign n438 = ~n434 & n437;
  assign n439 = n405 & ~n438;
  assign po015 = n433 | n439;
  assign n441 = ~pi095 & n351;
  assign n442 = n411 & n412;
  assign n443 = ~n441 & ~n442;
  assign po016 = n354 & n443;
  assign n445 = pi081 & n405;
  assign n446 = pi001 & ~n411;
  assign n447 = ~pi001 & n411;
  assign n448 = ~n446 & ~n447;
  assign n449 = ~n405 & ~n448;
  assign po017 = n445 | n449;
  assign n451 = pi082 & n405;
  assign n452 = pi001 & n411;
  assign n453 = pi002 & ~n452;
  assign n454 = ~pi002 & n411;
  assign n455 = pi001 & n454;
  assign n456 = ~n453 & ~n455;
  assign n457 = ~n405 & ~n456;
  assign po018 = n451 | n457;
  assign n459 = pi047 & ~pi127;
  assign po019 = pi000 | n459;
  assign po020 = pi047 & pi131;
  assign n462 = ~pi054 & pi055;
  assign n463 = pi054 & ~pi055;
  assign po022 = n462 | n463;
  assign n465 = pi054 & pi055;
  assign n466 = pi056 & ~n465;
  assign n467 = pi055 & ~pi056;
  assign n468 = pi054 & n467;
  assign po023 = n466 | n468;
  assign n470 = pi013 & ~pi015;
  assign n471 = pi016 & n470;
  assign n472 = ~pi055 & ~pi056;
  assign n473 = ~pi054 & n472;
  assign n474 = n471 & ~n473;
  assign po024 = pi089 & ~n474;
  assign n476 = n471 & ~n472;
  assign po025 = pi089 & ~n476;
  assign n478 = ~pi054 & ~pi056;
  assign n479 = n471 & ~n478;
  assign po026 = pi089 & ~n479;
  assign n481 = pi056 & n471;
  assign po027 = pi089 & ~n481;
  assign n483 = ~pi054 & ~pi055;
  assign n484 = n471 & ~n483;
  assign po028 = pi089 & ~n484;
  assign n486 = pi055 & n471;
  assign po029 = pi089 & ~n486;
  assign n488 = pi054 & n471;
  assign po030 = pi089 & ~n488;
  assign n490 = pi013 & pi054;
  assign n491 = pi055 & n490;
  assign po032 = pi056 & n491;
  assign n493 = ~pi053 & ~n305;
  assign po033 = ~n407 & ~n493;
  assign n495 = ~pi083 & pi084;
  assign n496 = pi085 & ~pi089;
  assign n497 = n495 & n496;
  assign po034 = pi000 | n497;
  assign n499 = ~pi089 & ~n495;
  assign po035 = pi085 & n499;
  assign n501 = ~pi085 & ~pi089;
  assign n502 = ~pi083 & ~pi084;
  assign n503 = ~n496 & ~n502;
  assign po036 = n501 | n503;
  assign n505 = pi014 & ~pi015;
  assign n506 = ~pi016 & n505;
  assign n507 = ~pi103 & ~pi104;
  assign n508 = ~pi105 & ~pi107;
  assign n509 = pi040 & pi089;
  assign n510 = pi105 & n509;
  assign n511 = ~n508 & ~n510;
  assign n512 = ~pi106 & ~n511;
  assign n513 = pi107 & n509;
  assign n514 = ~n512 & ~n513;
  assign n515 = pi104 & n321;
  assign n516 = ~pi103 & n515;
  assign n517 = ~n514 & ~n516;
  assign n518 = n507 & n517;
  assign n519 = pi116 & ~n321;
  assign n520 = pi111 & pi112;
  assign n521 = ~n519 & ~n520;
  assign n522 = n507 & ~n521;
  assign n523 = ~n518 & n522;
  assign n524 = pi048 & pi051;
  assign n525 = ~pi049 & pi050;
  assign n526 = pi049 & ~pi050;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~pi051 & ~n527;
  assign n529 = ~pi048 & n528;
  assign n530 = ~n524 & ~n529;
  assign n531 = ~pi049 & ~pi051;
  assign n532 = pi049 & pi051;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~pi048 & ~pi050;
  assign n535 = pi048 & pi050;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n533 & ~n536;
  assign n538 = pi072 & n537;
  assign n539 = n530 & ~n538;
  assign n540 = pi087 & ~n539;
  assign n541 = ~pi111 & pi112;
  assign n542 = pi111 & ~pi112;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~pi117 & ~pi118;
  assign n545 = ~pi123 & n544;
  assign n546 = pi078 & ~n545;
  assign n547 = pi032 & pi045;
  assign n548 = ~pi089 & n547;
  assign n549 = n538 & n548;
  assign n550 = ~pi129 & ~po102;
  assign n551 = ~n254 & ~n550;
  assign n552 = n506 & ~n530;
  assign n553 = pi089 & n552;
  assign n554 = n540 & ~n553;
  assign n555 = ~pi033 & n507;
  assign n556 = ~n355 & ~n555;
  assign n557 = pi098 & n556;
  assign n558 = pi045 & ~n557;
  assign n559 = ~pi115 & n558;
  assign n560 = ~n549 & ~n559;
  assign n561 = n546 & ~n560;
  assign n562 = ~n523 & ~n543;
  assign n563 = ~n561 & ~n562;
  assign n564 = ~n554 & n563;
  assign n565 = ~n551 & n564;
  assign n566 = pi036 & pi037;
  assign n567 = pi038 & n566;
  assign n568 = ~n540 & n567;
  assign n569 = ~pi033 & pi045;
  assign n570 = pi117 & n569;
  assign n571 = ~pi035 & ~n546;
  assign n572 = n568 & ~n570;
  assign n573 = n565 & n572;
  assign po037 = ~n571 & ~n573;
  assign n575 = ~pi032 & pi033;
  assign n576 = pi045 & n575;
  assign n577 = ~pi115 & n576;
  assign n578 = n546 & ~n570;
  assign n579 = ~pi035 & ~n578;
  assign n580 = n568 & ~n579;
  assign n581 = n565 & ~n577;
  assign po038 = n580 & n581;
  assign n583 = pi087 & n530;
  assign n584 = ~n538 & n583;
  assign n585 = ~pi118 & n546;
  assign po039 = n584 | n585;
  assign n587 = n546 & n555;
  assign n588 = pi036 & ~n587;
  assign po040 = pi089 | n588;
  assign n590 = pi098 & ~n355;
  assign n591 = n546 & ~n590;
  assign n592 = pi044 & n591;
  assign n593 = pi037 & ~n592;
  assign po041 = ~n316 | n593;
  assign n595 = ~pi014 & ~n541;
  assign n596 = ~pi093 & ~n595;
  assign n597 = pi089 & ~n596;
  assign n598 = ~pi016 & n597;
  assign n599 = pi015 & n598;
  assign n600 = ~pi076 & pi090;
  assign n601 = ~pi074 & pi075;
  assign n602 = n600 & n601;
  assign n603 = ~pi038 & ~n602;
  assign n604 = ~n599 & n603;
  assign po042 = ~n577 & ~n604;
  assign po043 = pi117 & n580;
  assign n607 = pi089 & n506;
  assign n608 = pi088 & ~n607;
  assign po044 = n549 | n608;
  assign n610 = pi045 & pi115;
  assign n611 = pi032 & n610;
  assign po045 = n540 | n611;
  assign n613 = ~pi086 & ~pi088;
  assign n614 = ~po102 & ~n570;
  assign po046 = ~n613 | ~n614;
  assign n616 = ~pi023 & pi024;
  assign n617 = pi039 & ~n616;
  assign n618 = pi030 & n616;
  assign po047 = n617 | n618;
  assign n620 = ~pi064 & ~pi094;
  assign n621 = ~pi043 & n620;
  assign po048 = pi090 & ~n621;
  assign n623 = pi074 & pi075;
  assign n624 = ~pi076 & n623;
  assign po049 = pi090 & n624;
  assign n626 = ~pi093 & pi094;
  assign n627 = pi093 & ~pi094;
  assign po051 = n626 | n627;
  assign n629 = ~pi093 & ~pi094;
  assign n630 = ~pi043 & n629;
  assign po052 = pi090 & ~n630;
  assign n632 = pi015 & ~pi090;
  assign n633 = n287 & n632;
  assign n634 = ~n291 & ~n633;
  assign n635 = ~pi041 & ~n634;
  assign n636 = pi125 & n634;
  assign po053 = n635 | n636;
  assign n638 = pi126 & n634;
  assign n639 = pi041 & ~pi042;
  assign n640 = ~pi041 & pi042;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n634 & ~n641;
  assign po054 = n638 | n642;
  assign po055 = pi115 & n580;
  assign n645 = pi089 & n287;
  assign n646 = ~n321 & ~n645;
  assign n647 = pi043 & n646;
  assign po056 = n577 | n647;
  assign po057 = ~pi038 & ~pi088;
  assign n650 = pi038 & ~pi093;
  assign n651 = pi090 & ~n541;
  assign n652 = n650 & ~n651;
  assign po058 = ~pi088 & ~n652;
  assign n654 = ~n518 & n569;
  assign n655 = n507 & n654;
  assign n656 = pi111 & n523;
  assign n657 = ~n577 & ~n656;
  assign po059 = n655 | ~n657;
  assign n659 = pi112 & n523;
  assign n660 = ~pi112 & ~n523;
  assign n661 = pi111 & n660;
  assign n662 = ~n659 & ~n661;
  assign po060 = n655 | ~n662;
  assign n664 = n507 & ~n518;
  assign n665 = ~n321 & ~n543;
  assign n666 = pi116 & n665;
  assign n667 = ~n655 & ~n666;
  assign n668 = ~n520 & n667;
  assign n669 = ~n664 & ~n668;
  assign n670 = n518 & ~n669;
  assign n671 = n543 & ~n670;
  assign n672 = ~n518 & ~n669;
  assign n673 = ~n671 & ~n672;
  assign n674 = pi103 & ~n673;
  assign n675 = ~n254 & n669;
  assign po061 = n674 | n675;
  assign n677 = ~pi103 & n321;
  assign n678 = ~n283 & ~n670;
  assign n679 = ~n672 & ~n678;
  assign n680 = ~n677 & ~n679;
  assign n681 = pi104 & n680;
  assign n682 = ~pi020 & n418;
  assign n683 = ~pi033 & n419;
  assign n684 = ~n682 & ~n683;
  assign n685 = n543 & n684;
  assign n686 = n669 & ~n685;
  assign po062 = n681 | n686;
  assign n688 = ~pi105 & ~pi106;
  assign n689 = pi040 & ~n688;
  assign n690 = pi103 & n518;
  assign n691 = ~n518 & ~n689;
  assign n692 = pi105 & n691;
  assign po063 = n690 | n692;
  assign n694 = ~pi105 & n321;
  assign n695 = ~n518 & ~n694;
  assign n696 = ~n689 & n695;
  assign n697 = pi106 & n696;
  assign n698 = pi104 & n518;
  assign po064 = n697 | n698;
  assign n700 = pi106 & n689;
  assign n701 = ~pi040 & ~n518;
  assign n702 = pi107 & n701;
  assign po065 = n700 | n702;
  assign n704 = ~pi088 & n607;
  assign po066 = n584 | n704;
  assign po067 = ~n538 & n547;
  assign po068 = ~pi050 & ~pi051;
  assign po070 = ~pi048 & ~pi049;
  assign n709 = pi016 & pi089;
  assign n710 = pi093 & n709;
  assign n711 = pi094 & n710;
  assign n712 = pi070 & n320;
  assign n713 = pi066 & ~pi128;
  assign n714 = ~pi064 & ~n713;
  assign n715 = ~n712 & ~n714;
  assign po075 = ~n711 & n715;
  assign n717 = ~pi060 & ~n713;
  assign n718 = pi064 & ~n712;
  assign n719 = n629 & n709;
  assign n720 = ~n718 & n719;
  assign n721 = ~n717 & ~n720;
  assign po076 = ~n711 & n721;
  assign n723 = pi060 & pi134;
  assign n724 = pi129 & ~n336;
  assign n725 = pi128 & n724;
  assign po077 = n723 & n725;
  assign n727 = ~pi064 & n629;
  assign po078 = pi090 & ~n727;
  assign n729 = ~n287 & n293;
  assign n730 = pi016 & ~pi090;
  assign n731 = n287 & n730;
  assign n732 = ~n729 & ~n731;
  assign n733 = ~pi062 & ~n732;
  assign n734 = pi120 & n732;
  assign po079 = n733 | n734;
  assign n736 = pi121 & n732;
  assign n737 = pi062 & ~pi063;
  assign n738 = ~pi062 & pi063;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n732 & ~n739;
  assign po080 = n736 | n740;
  assign po081 = pi128 & n723;
  assign po082 = ~pi064 & ~po102;
  assign po083 = pi060 | n293;
  assign n745 = pi018 & ~pi115;
  assign n746 = pi098 & n405;
  assign n747 = ~n745 & ~n746;
  assign po084 = n335 | ~n747;
  assign n749 = ~n307 & ~n545;
  assign po085 = ~n335 & n749;
  assign po086 = ~n307 & n335;
  assign n752 = ~n335 & n545;
  assign po087 = n307 | n752;
  assign n754 = pi099 & n355;
  assign n755 = n307 & ~n754;
  assign n756 = ~n580 & ~n723;
  assign n757 = ~n338 & ~n756;
  assign n758 = ~n335 & n757;
  assign n759 = ~n321 & ~n332;
  assign n760 = pi102 & n759;
  assign n761 = n335 & ~n760;
  assign n762 = ~n758 & ~n761;
  assign n763 = ~n340 & ~n762;
  assign n764 = ~n335 & ~n723;
  assign n765 = ~n580 & n764;
  assign n766 = ~n355 & ~n765;
  assign n767 = ~n763 & ~n766;
  assign n768 = ~n755 & n767;
  assign n769 = pi130 & ~n768;
  assign po088 = ~po102 & n769;
  assign n771 = n251 & ~n270;
  assign n772 = ~pi133 & ~n771;
  assign n773 = ~po102 & n772;
  assign po089 = ~pi070 & ~n773;
  assign n775 = pi070 & ~n773;
  assign po090 = ~pi069 & n775;
  assign n777 = pi046 & pi096;
  assign n778 = ~pi114 & pi119;
  assign n779 = pi017 & ~n778;
  assign po096 = n777 | n779;
  assign po097 = pi113 & pi119;
  assign n782 = pi010 & ~pi029;
  assign n783 = pi012 & pi029;
  assign po098 = n782 | n783;
  assign po099 = pi132 | n771;
  assign n786 = ~pi100 & pi101;
  assign n787 = n251 & n786;
  assign po100 = n270 & n787;
  assign n789 = pi100 & ~n251;
  assign po101 = ~pi130 | n789;
  assign n791 = pi101 & ~po102;
  assign po106 = ~pi100 & ~n791;
  assign po006 = ~pi118;
  assign po050 = ~pi093;
  assign po005 = pi122;
  assign po007 = pi123;
  assign po021 = pi090;
  assign po031 = pi089;
  assign po069 = pi050;
  assign po071 = pi048;
  assign po072 = po068;
  assign po073 = pi050;
  assign po074 = pi051;
  assign po091 = pi022;
  assign po092 = pi025;
  assign po093 = pi026;
  assign po094 = pi027;
  assign po095 = pi028;
  assign po103 = po070;
  assign po104 = pi048;
  assign po105 = pi049;
endmodule



// Benchmark "too_large" written by ABC on Sun Apr 22 21:43:15 2018

module too_large ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37,
    po0, po1, po2  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37;
  output po0, po1, po2;
  wire n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864;
  assign n42 = pi02 & ~pi12;
  assign n43 = ~pi14 & n42;
  assign n44 = ~pi15 & n43;
  assign n45 = ~pi19 & n44;
  assign n46 = ~pi20 & n45;
  assign n47 = ~pi22 & n46;
  assign n48 = ~pi23 & n47;
  assign n49 = ~pi25 & n48;
  assign n50 = ~pi26 & n49;
  assign n51 = ~pi27 & n50;
  assign n52 = pi28 & n51;
  assign n53 = ~pi13 & n42;
  assign n54 = ~pi15 & n53;
  assign n55 = ~pi19 & n54;
  assign n56 = ~pi20 & n55;
  assign n57 = ~pi22 & n56;
  assign n58 = ~pi23 & n57;
  assign n59 = ~pi25 & n58;
  assign n60 = ~pi26 & n59;
  assign n61 = ~pi27 & n60;
  assign n62 = pi28 & n61;
  assign n63 = ~pi12 & ~pi14;
  assign n64 = ~pi15 & n63;
  assign n65 = ~pi22 & n64;
  assign n66 = pi24 & n65;
  assign n67 = ~pi26 & n66;
  assign n68 = ~pi27 & n67;
  assign n69 = ~pi28 & n68;
  assign n70 = pi32 & n69;
  assign n71 = ~pi33 & n70;
  assign n72 = pi34 & n71;
  assign n73 = ~pi14 & ~pi15;
  assign n74 = ~pi16 & n73;
  assign n75 = ~pi22 & n74;
  assign n76 = pi24 & n75;
  assign n77 = ~pi26 & n76;
  assign n78 = ~pi27 & n77;
  assign n79 = ~pi28 & n78;
  assign n80 = pi32 & n79;
  assign n81 = ~pi33 & n80;
  assign n82 = pi34 & n81;
  assign n83 = pi19 & n64;
  assign n84 = ~pi20 & n83;
  assign n85 = ~pi21 & n84;
  assign n86 = ~pi22 & n85;
  assign n87 = ~pi23 & n86;
  assign n88 = ~pi25 & n87;
  assign n89 = ~pi26 & n88;
  assign n90 = ~pi27 & n89;
  assign n91 = pi28 & n90;
  assign n92 = pi19 & n74;
  assign n93 = ~pi20 & n92;
  assign n94 = ~pi21 & n93;
  assign n95 = ~pi22 & n94;
  assign n96 = ~pi23 & n95;
  assign n97 = ~pi25 & n96;
  assign n98 = ~pi26 & n97;
  assign n99 = ~pi27 & n98;
  assign n100 = pi28 & n99;
  assign n101 = ~pi12 & ~pi13;
  assign n102 = ~pi15 & n101;
  assign n103 = pi19 & n102;
  assign n104 = ~pi20 & n103;
  assign n105 = ~pi21 & n104;
  assign n106 = ~pi22 & n105;
  assign n107 = ~pi23 & n106;
  assign n108 = ~pi25 & n107;
  assign n109 = ~pi26 & n108;
  assign n110 = ~pi27 & n109;
  assign n111 = pi28 & n110;
  assign n112 = ~pi13 & ~pi15;
  assign n113 = ~pi16 & n112;
  assign n114 = pi19 & n113;
  assign n115 = ~pi20 & n114;
  assign n116 = ~pi21 & n115;
  assign n117 = ~pi22 & n116;
  assign n118 = ~pi23 & n117;
  assign n119 = ~pi25 & n118;
  assign n120 = ~pi26 & n119;
  assign n121 = ~pi27 & n120;
  assign n122 = pi28 & n121;
  assign n123 = pi14 & n101;
  assign n124 = ~pi15 & n123;
  assign n125 = ~pi22 & n124;
  assign n126 = ~pi26 & n125;
  assign n127 = ~pi27 & n126;
  assign n128 = ~pi28 & n127;
  assign n129 = pi32 & n128;
  assign n130 = ~pi33 & n129;
  assign n131 = pi34 & n130;
  assign n132 = ~pi13 & pi14;
  assign n133 = ~pi15 & n132;
  assign n134 = ~pi16 & n133;
  assign n135 = ~pi22 & n134;
  assign n136 = ~pi26 & n135;
  assign n137 = ~pi27 & n136;
  assign n138 = ~pi28 & n137;
  assign n139 = pi32 & n138;
  assign n140 = ~pi33 & n139;
  assign n141 = pi34 & n140;
  assign n142 = pi21 & n64;
  assign n143 = ~pi22 & n142;
  assign n144 = ~pi26 & n143;
  assign n145 = ~pi27 & n144;
  assign n146 = pi28 & n145;
  assign n147 = ~pi33 & n146;
  assign n148 = pi34 & n147;
  assign n149 = pi21 & n74;
  assign n150 = ~pi22 & n149;
  assign n151 = ~pi26 & n150;
  assign n152 = ~pi27 & n151;
  assign n153 = pi28 & n152;
  assign n154 = ~pi33 & n153;
  assign n155 = pi34 & n154;
  assign n156 = pi21 & n102;
  assign n157 = ~pi22 & n156;
  assign n158 = ~pi26 & n157;
  assign n159 = ~pi27 & n158;
  assign n160 = pi28 & n159;
  assign n161 = ~pi33 & n160;
  assign n162 = pi34 & n161;
  assign n163 = ~pi23 & n65;
  assign n164 = pi24 & n163;
  assign n165 = ~pi26 & n164;
  assign n166 = ~pi27 & n165;
  assign n167 = ~pi28 & n166;
  assign n168 = pi32 & n167;
  assign n169 = pi33 & n168;
  assign n170 = pi21 & n113;
  assign n171 = ~pi22 & n170;
  assign n172 = ~pi26 & n171;
  assign n173 = ~pi27 & n172;
  assign n174 = pi28 & n173;
  assign n175 = ~pi33 & n174;
  assign n176 = pi34 & n175;
  assign n177 = ~pi23 & n75;
  assign n178 = pi24 & n177;
  assign n179 = ~pi26 & n178;
  assign n180 = ~pi27 & n179;
  assign n181 = ~pi28 & n180;
  assign n182 = pi32 & n181;
  assign n183 = pi33 & n182;
  assign n184 = pi24 & ~pi27;
  assign n185 = ~pi28 & n184;
  assign n186 = ~pi29 & n185;
  assign n187 = ~pi30 & n186;
  assign n188 = ~pi31 & n187;
  assign n189 = pi32 & n188;
  assign n190 = ~pi33 & n189;
  assign n191 = pi34 & n190;
  assign n192 = ~pi23 & pi24;
  assign n193 = ~pi25 & n192;
  assign n194 = ~pi27 & n193;
  assign n195 = ~pi28 & n194;
  assign n196 = ~pi29 & n195;
  assign n197 = ~pi30 & n196;
  assign n198 = ~pi31 & n197;
  assign n199 = pi32 & n198;
  assign n200 = ~pi33 & n199;
  assign n201 = ~pi22 & ~pi23;
  assign n202 = pi24 & n201;
  assign n203 = ~pi27 & n202;
  assign n204 = ~pi28 & n203;
  assign n205 = ~pi29 & n204;
  assign n206 = ~pi30 & n205;
  assign n207 = ~pi31 & n206;
  assign n208 = pi32 & n207;
  assign n209 = pi33 & n208;
  assign n210 = pi14 & ~pi27;
  assign n211 = ~pi28 & n210;
  assign n212 = ~pi29 & n211;
  assign n213 = ~pi30 & n212;
  assign n214 = ~pi31 & n213;
  assign n215 = pi32 & n214;
  assign n216 = ~pi33 & n215;
  assign n217 = pi34 & n216;
  assign n218 = ~pi23 & n125;
  assign n219 = ~pi26 & n218;
  assign n220 = ~pi27 & n219;
  assign n221 = ~pi28 & n220;
  assign n222 = pi32 & n221;
  assign n223 = pi33 & n222;
  assign n224 = ~pi23 & n135;
  assign n225 = ~pi26 & n224;
  assign n226 = ~pi27 & n225;
  assign n227 = ~pi28 & n226;
  assign n228 = pi32 & n227;
  assign n229 = pi33 & n228;
  assign n230 = ~pi23 & n143;
  assign n231 = ~pi26 & n230;
  assign n232 = ~pi27 & n231;
  assign n233 = pi28 & n232;
  assign n234 = pi33 & n233;
  assign n235 = ~pi23 & n150;
  assign n236 = ~pi26 & n235;
  assign n237 = ~pi27 & n236;
  assign n238 = pi28 & n237;
  assign n239 = pi33 & n238;
  assign n240 = ~pi25 & n164;
  assign n241 = ~pi26 & n240;
  assign n242 = ~pi27 & n241;
  assign n243 = pi32 & n242;
  assign n244 = pi14 & ~pi22;
  assign n245 = ~pi23 & n244;
  assign n246 = ~pi27 & n245;
  assign n247 = ~pi28 & n246;
  assign n248 = ~pi29 & n247;
  assign n249 = ~pi30 & n248;
  assign n250 = ~pi31 & n249;
  assign n251 = pi32 & n250;
  assign n252 = pi33 & n251;
  assign n253 = ~pi25 & n178;
  assign n254 = ~pi26 & n253;
  assign n255 = ~pi27 & n254;
  assign n256 = pi32 & n255;
  assign n257 = pi21 & ~pi27;
  assign n258 = pi28 & n257;
  assign n259 = ~pi29 & n258;
  assign n260 = ~pi30 & n259;
  assign n261 = ~pi31 & n260;
  assign n262 = ~pi33 & n261;
  assign n263 = pi34 & n262;
  assign n264 = ~pi23 & n157;
  assign n265 = ~pi26 & n264;
  assign n266 = ~pi27 & n265;
  assign n267 = pi28 & n266;
  assign n268 = pi33 & n267;
  assign n269 = ~pi25 & n230;
  assign n270 = ~pi26 & n269;
  assign n271 = ~pi27 & n270;
  assign n272 = pi28 & n271;
  assign n273 = ~pi23 & n171;
  assign n274 = ~pi26 & n273;
  assign n275 = ~pi27 & n274;
  assign n276 = pi28 & n275;
  assign n277 = pi33 & n276;
  assign n278 = ~pi25 & n235;
  assign n279 = ~pi26 & n278;
  assign n280 = ~pi27 & n279;
  assign n281 = pi28 & n280;
  assign n282 = pi21 & ~pi23;
  assign n283 = ~pi25 & n282;
  assign n284 = ~pi27 & n283;
  assign n285 = pi28 & n284;
  assign n286 = ~pi29 & n285;
  assign n287 = ~pi30 & n286;
  assign n288 = ~pi31 & n287;
  assign n289 = ~pi33 & n288;
  assign n290 = ~pi25 & n264;
  assign n291 = ~pi26 & n290;
  assign n292 = ~pi27 & n291;
  assign n293 = pi28 & n292;
  assign n294 = pi21 & ~pi22;
  assign n295 = ~pi23 & n294;
  assign n296 = ~pi27 & n295;
  assign n297 = pi28 & n296;
  assign n298 = ~pi29 & n297;
  assign n299 = ~pi30 & n298;
  assign n300 = ~pi31 & n299;
  assign n301 = pi33 & n300;
  assign n302 = ~pi25 & n273;
  assign n303 = ~pi26 & n302;
  assign n304 = ~pi27 & n303;
  assign n305 = pi28 & n304;
  assign n306 = ~pi33 & pi34;
  assign n307 = ~pi23 & pi33;
  assign n308 = ~n306 & ~n307;
  assign n309 = pi13 & pi14;
  assign n310 = pi08 & pi31;
  assign n311 = ~pi02 & ~pi04;
  assign n312 = ~pi01 & ~pi06;
  assign n313 = ~pi05 & n312;
  assign n314 = n311 & n313;
  assign n315 = pi29 & ~n314;
  assign n316 = ~n310 & ~n315;
  assign n317 = pi35 & n316;
  assign n318 = ~pi07 & n317;
  assign n319 = ~pi09 & pi30;
  assign n320 = pi07 & n319;
  assign n321 = ~n318 & ~n320;
  assign n322 = ~pi28 & ~n321;
  assign n323 = pi07 & ~pi09;
  assign n324 = pi20 & pi30;
  assign n325 = n323 & n324;
  assign n326 = pi19 & ~pi20;
  assign n327 = pi28 & n326;
  assign n328 = ~n325 & ~n327;
  assign n329 = ~n322 & n328;
  assign n330 = ~n309 & ~n329;
  assign n331 = ~pi11 & ~pi18;
  assign n332 = pi03 & ~pi17;
  assign n333 = pi10 & ~n332;
  assign n334 = ~n331 & n333;
  assign n335 = ~pi13 & ~n334;
  assign n336 = pi13 & ~pi14;
  assign n337 = ~n335 & ~n336;
  assign n338 = ~n310 & ~n337;
  assign n339 = pi35 & n338;
  assign n340 = ~pi09 & n339;
  assign n341 = ~pi07 & n340;
  assign n342 = ~pi06 & n341;
  assign n343 = ~pi05 & n342;
  assign n344 = ~pi04 & n343;
  assign n345 = ~pi02 & n344;
  assign n346 = ~n331 & ~n332;
  assign n347 = ~pi13 & ~n346;
  assign n348 = ~n336 & ~n347;
  assign n349 = pi30 & ~n348;
  assign n350 = pi10 & n349;
  assign n351 = pi07 & n350;
  assign n352 = ~n345 & ~n351;
  assign n353 = ~pi28 & ~n352;
  assign n354 = pi07 & pi13;
  assign n355 = pi10 & pi30;
  assign n356 = n354 & n355;
  assign n357 = pi24 & pi32;
  assign n358 = ~n356 & ~n357;
  assign n359 = ~pi14 & ~n358;
  assign n360 = pi30 & ~n346;
  assign n361 = pi10 & n360;
  assign n362 = pi07 & n361;
  assign n363 = pi14 & pi32;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~pi13 & ~n364;
  assign n366 = ~n359 & ~n365;
  assign n367 = pi20 & ~n366;
  assign n368 = ~n353 & ~n367;
  assign n369 = ~n330 & n368;
  assign n370 = ~n308 & ~n369;
  assign n371 = ~pi30 & ~pi34;
  assign n372 = pi07 & ~n371;
  assign n373 = pi20 & pi28;
  assign n374 = ~pi01 & ~n373;
  assign n375 = ~pi06 & n374;
  assign n376 = ~pi05 & n375;
  assign n377 = ~pi04 & n376;
  assign n378 = ~pi20 & ~pi29;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~n372 & ~n379;
  assign n381 = ~pi25 & n380;
  assign n382 = ~pi04 & ~pi05;
  assign n383 = ~pi06 & ~pi28;
  assign n384 = n382 & n383;
  assign n385 = pi33 & ~pi34;
  assign n386 = ~pi01 & ~pi30;
  assign n387 = n385 & n386;
  assign n388 = n384 & n387;
  assign n389 = ~n381 & ~n388;
  assign n390 = ~pi02 & ~n389;
  assign n391 = ~pi07 & ~pi28;
  assign n392 = ~pi25 & ~pi29;
  assign n393 = n391 & n392;
  assign n394 = ~n390 & ~n393;
  assign n395 = ~n310 & ~n394;
  assign n396 = pi25 & ~pi33;
  assign n397 = ~pi29 & ~n396;
  assign n398 = ~pi30 & n397;
  assign n399 = ~pi34 & n398;
  assign n400 = ~pi28 & n399;
  assign n401 = ~pi08 & n400;
  assign n402 = ~n395 & ~n401;
  assign n403 = pi35 & ~n402;
  assign n404 = pi00 & ~pi20;
  assign n405 = pi28 & n404;
  assign n406 = ~n320 & ~n405;
  assign n407 = ~pi25 & ~n406;
  assign n408 = ~n403 & ~n407;
  assign n409 = ~n309 & ~n408;
  assign n410 = ~pi28 & ~n396;
  assign n411 = ~pi02 & n410;
  assign n412 = ~pi20 & ~pi25;
  assign n413 = pi28 & n412;
  assign n414 = ~n411 & ~n413;
  assign n415 = ~pi34 & ~n414;
  assign n416 = ~pi07 & pi28;
  assign n417 = n412 & n416;
  assign n418 = ~n415 & ~n417;
  assign n419 = ~n310 & ~n418;
  assign n420 = pi35 & n419;
  assign n421 = ~pi06 & n420;
  assign n422 = ~pi05 & n421;
  assign n423 = ~pi04 & n422;
  assign n424 = pi02 & pi28;
  assign n425 = n412 & n424;
  assign n426 = ~n423 & ~n425;
  assign n427 = ~pi09 & ~n426;
  assign n428 = pi07 & ~pi25;
  assign n429 = n355 & n428;
  assign n430 = ~n427 & ~n429;
  assign n431 = ~n348 & ~n430;
  assign n432 = ~pi10 & ~n426;
  assign n433 = ~pi09 & n432;
  assign n434 = ~pi25 & n363;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~pi13 & ~n435;
  assign n437 = ~n431 & ~n436;
  assign n438 = ~n409 & n437;
  assign n439 = ~pi23 & ~n438;
  assign n440 = ~n370 & ~n439;
  assign n441 = ~pi16 & ~n440;
  assign n442 = ~pi20 & pi28;
  assign n443 = ~pi09 & ~n309;
  assign n444 = pi10 & ~n348;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~n442 & ~n445;
  assign n447 = pi30 & n446;
  assign n448 = pi07 & n447;
  assign n449 = ~pi05 & ~pi06;
  assign n450 = n311 & n449;
  assign n451 = pi29 & ~n450;
  assign n452 = ~n310 & ~n451;
  assign n453 = pi35 & n452;
  assign n454 = ~pi28 & n453;
  assign n455 = ~pi07 & n454;
  assign n456 = ~n327 & ~n455;
  assign n457 = ~n309 & ~n456;
  assign n458 = ~pi14 & pi24;
  assign n459 = ~n132 & ~n458;
  assign n460 = pi32 & ~n459;
  assign n461 = pi20 & n460;
  assign n462 = ~n457 & ~n461;
  assign n463 = ~n448 & n462;
  assign n464 = ~n308 & ~n463;
  assign n465 = ~pi02 & ~pi28;
  assign n466 = ~n442 & ~n465;
  assign n467 = ~pi06 & ~n466;
  assign n468 = ~pi05 & n467;
  assign n469 = ~pi04 & n468;
  assign n470 = ~n378 & ~n469;
  assign n471 = ~n372 & ~n470;
  assign n472 = ~pi28 & ~pi29;
  assign n473 = ~pi07 & n472;
  assign n474 = ~n471 & ~n473;
  assign n475 = ~pi25 & ~n474;
  assign n476 = ~pi28 & pi33;
  assign n477 = n371 & n476;
  assign n478 = n450 & n477;
  assign n479 = ~n475 & ~n478;
  assign n480 = ~n310 & ~n479;
  assign n481 = ~n401 & ~n480;
  assign n482 = pi35 & ~n481;
  assign n483 = ~n407 & ~n482;
  assign n484 = ~n309 & ~n483;
  assign n485 = ~pi13 & n363;
  assign n486 = ~n351 & ~n485;
  assign n487 = ~pi25 & ~n486;
  assign n488 = ~n484 & ~n487;
  assign n489 = ~pi23 & ~n488;
  assign n490 = ~n464 & ~n489;
  assign n491 = ~pi12 & ~n490;
  assign n492 = ~n441 & ~n491;
  assign n493 = ~pi26 & ~n492;
  assign n494 = ~pi15 & n493;
  assign n495 = pi07 & pi34;
  assign n496 = pi35 & ~n495;
  assign n497 = ~pi28 & n496;
  assign n498 = ~pi14 & ~pi24;
  assign n499 = pi32 & ~n498;
  assign n500 = pi20 & n499;
  assign n501 = ~n327 & ~n500;
  assign n502 = ~n497 & n501;
  assign n503 = ~pi29 & ~n502;
  assign n504 = ~pi30 & n503;
  assign n505 = ~pi23 & n504;
  assign n506 = ~pi31 & n505;
  assign n507 = pi33 & n506;
  assign n508 = ~n494 & ~n507;
  assign n509 = ~pi22 & ~n508;
  assign n510 = ~pi23 & ~pi25;
  assign n511 = ~pi34 & ~n510;
  assign n512 = ~n501 & ~n511;
  assign n513 = ~pi07 & pi34;
  assign n514 = ~pi34 & n510;
  assign n515 = ~n513 & ~n514;
  assign n516 = pi35 & ~n515;
  assign n517 = n363 & n510;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~pi28 & ~n518;
  assign n520 = ~n512 & ~n519;
  assign n521 = ~pi29 & ~n520;
  assign n522 = ~pi30 & n521;
  assign n523 = ~pi31 & n522;
  assign n524 = ~pi33 & n523;
  assign n525 = ~n509 & ~n524;
  assign n526 = ~pi27 & ~n525;
  assign n527 = ~n52 & ~n62;
  assign n528 = ~n72 & ~n82;
  assign n529 = n527 & n528;
  assign n530 = ~n91 & ~n100;
  assign n531 = ~n122 & ~n131;
  assign n532 = ~n111 & n531;
  assign n533 = n530 & n532;
  assign n534 = n529 & n533;
  assign n535 = ~n141 & ~n148;
  assign n536 = ~n155 & ~n162;
  assign n537 = n535 & n536;
  assign n538 = ~n169 & ~n176;
  assign n539 = ~n191 & ~n200;
  assign n540 = ~n183 & n539;
  assign n541 = n538 & n540;
  assign n542 = n537 & n541;
  assign n543 = n534 & n542;
  assign n544 = ~n209 & ~n217;
  assign n545 = ~n223 & ~n229;
  assign n546 = n544 & n545;
  assign n547 = ~n234 & ~n239;
  assign n548 = ~n252 & ~n256;
  assign n549 = ~n243 & n548;
  assign n550 = n547 & n549;
  assign n551 = n546 & n550;
  assign n552 = ~n263 & ~n268;
  assign n553 = ~n272 & ~n277;
  assign n554 = n552 & n553;
  assign n555 = ~n281 & ~n289;
  assign n556 = ~n301 & ~n305;
  assign n557 = ~n293 & n556;
  assign n558 = n555 & n557;
  assign n559 = n554 & n558;
  assign n560 = n551 & n559;
  assign n561 = n543 & n560;
  assign po0 = n526 | ~n561;
  assign n563 = pi20 & n64;
  assign n564 = ~pi21 & n563;
  assign n565 = ~pi22 & n564;
  assign n566 = ~pi23 & n565;
  assign n567 = ~pi25 & n566;
  assign n568 = ~pi26 & n567;
  assign n569 = ~pi27 & n568;
  assign n570 = pi28 & n569;
  assign n571 = pi20 & n74;
  assign n572 = ~pi21 & n571;
  assign n573 = ~pi22 & n572;
  assign n574 = ~pi23 & n573;
  assign n575 = ~pi25 & n574;
  assign n576 = ~pi26 & n575;
  assign n577 = ~pi27 & n576;
  assign n578 = pi28 & n577;
  assign n579 = pi20 & n102;
  assign n580 = ~pi21 & n579;
  assign n581 = ~pi22 & n580;
  assign n582 = ~pi23 & n581;
  assign n583 = ~pi25 & n582;
  assign n584 = ~pi26 & n583;
  assign n585 = ~pi27 & n584;
  assign n586 = pi28 & n585;
  assign n587 = pi20 & n113;
  assign n588 = ~pi21 & n587;
  assign n589 = ~pi22 & n588;
  assign n590 = ~pi23 & n589;
  assign n591 = ~pi25 & n590;
  assign n592 = ~pi26 & n591;
  assign n593 = ~pi27 & n592;
  assign n594 = pi28 & n593;
  assign n595 = pi12 & pi16;
  assign n596 = ~pi19 & pi28;
  assign n597 = pi30 & ~n596;
  assign n598 = pi07 & n597;
  assign n599 = pi19 & n357;
  assign n600 = ~n373 & ~n599;
  assign n601 = ~n598 & n600;
  assign n602 = ~n308 & ~n601;
  assign n603 = pi07 & ~pi23;
  assign n604 = ~pi25 & pi30;
  assign n605 = n603 & n604;
  assign n606 = ~n602 & ~n605;
  assign n607 = ~n595 & ~n606;
  assign n608 = ~pi19 & ~pi23;
  assign n609 = ~pi16 & n608;
  assign n610 = ~pi25 & n424;
  assign n611 = n609 & n610;
  assign n612 = ~n607 & ~n611;
  assign n613 = ~n309 & ~n612;
  assign n614 = pi25 & ~n476;
  assign n615 = pi24 & ~n614;
  assign n616 = pi32 & n615;
  assign n617 = ~pi08 & ~pi34;
  assign n618 = pi30 & ~pi31;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~n396 & ~n619;
  assign n621 = ~pi08 & pi33;
  assign n622 = ~pi07 & n621;
  assign n623 = ~n620 & ~n622;
  assign n624 = ~pi28 & ~n623;
  assign n625 = ~n310 & ~n495;
  assign n626 = ~pi25 & n625;
  assign n627 = ~pi19 & n626;
  assign n628 = ~pi00 & n627;
  assign n629 = ~n624 & ~n628;
  assign n630 = ~pi29 & ~n629;
  assign n631 = pi36 & n630;
  assign n632 = ~pi32 & n631;
  assign n633 = ~n616 & ~n632;
  assign n634 = ~pi13 & ~n633;
  assign n635 = ~pi14 & n630;
  assign n636 = pi36 & n635;
  assign n637 = ~n634 & ~n636;
  assign n638 = ~pi23 & ~n637;
  assign n639 = ~pi13 & ~pi32;
  assign n640 = pi14 & ~n639;
  assign n641 = ~pi07 & ~pi08;
  assign n642 = ~n618 & ~n641;
  assign n643 = ~n640 & ~n642;
  assign n644 = ~pi29 & n643;
  assign n645 = pi36 & n644;
  assign n646 = ~pi13 & n357;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~pi33 & ~n647;
  assign n649 = pi34 & n648;
  assign n650 = ~pi28 & n649;
  assign n651 = ~n638 & ~n650;
  assign n652 = ~n595 & ~n651;
  assign n653 = ~pi00 & ~pi19;
  assign n654 = ~pi25 & pi28;
  assign n655 = n653 & n654;
  assign n656 = ~pi02 & pi33;
  assign n657 = ~pi28 & n656;
  assign n658 = ~n655 & ~n657;
  assign n659 = ~pi09 & ~n334;
  assign n660 = pi01 & ~n659;
  assign n661 = ~pi16 & ~n660;
  assign n662 = pi12 & ~n661;
  assign n663 = ~n640 & ~n662;
  assign n664 = ~pi09 & pi13;
  assign n665 = ~pi14 & ~pi16;
  assign n666 = n664 & n665;
  assign n667 = ~n663 & ~n666;
  assign n668 = ~n658 & ~n667;
  assign n669 = ~n495 & n668;
  assign n670 = ~pi02 & ~n667;
  assign n671 = ~pi34 & n670;
  assign n672 = ~pi28 & n671;
  assign n673 = ~pi25 & n672;
  assign n674 = ~n669 & ~n673;
  assign n675 = ~pi23 & ~n674;
  assign n676 = ~pi33 & ~n667;
  assign n677 = ~pi02 & n676;
  assign n678 = pi34 & n677;
  assign n679 = ~pi28 & n678;
  assign n680 = ~pi07 & n679;
  assign n681 = ~n675 & ~n680;
  assign n682 = ~n310 & ~n681;
  assign n683 = pi36 & n682;
  assign n684 = ~pi06 & n683;
  assign n685 = ~pi05 & n684;
  assign n686 = ~pi04 & n685;
  assign n687 = ~n652 & ~n686;
  assign n688 = ~n613 & n687;
  assign n689 = ~pi26 & ~n688;
  assign n690 = ~pi15 & n689;
  assign n691 = ~n363 & ~n495;
  assign n692 = pi36 & n691;
  assign n693 = ~pi28 & n692;
  assign n694 = n600 & ~n693;
  assign n695 = ~pi30 & ~n694;
  assign n696 = ~pi29 & n695;
  assign n697 = pi33 & n696;
  assign n698 = ~pi31 & n697;
  assign n699 = ~pi23 & n698;
  assign n700 = ~n690 & ~n699;
  assign n701 = ~pi22 & ~n700;
  assign n702 = ~pi25 & ~pi34;
  assign n703 = ~pi23 & n702;
  assign n704 = ~n513 & ~n703;
  assign n705 = ~n363 & ~n704;
  assign n706 = pi36 & n705;
  assign n707 = ~pi28 & n706;
  assign n708 = ~n511 & ~n600;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~pi30 & ~n709;
  assign n711 = ~pi29 & n710;
  assign n712 = ~pi33 & n711;
  assign n713 = ~pi31 & n712;
  assign n714 = ~n701 & ~n713;
  assign n715 = ~pi27 & ~n714;
  assign n716 = ~n62 & ~n72;
  assign n717 = ~n52 & n716;
  assign n718 = ~n82 & ~n148;
  assign n719 = n536 & n718;
  assign n720 = n717 & n719;
  assign n721 = ~n183 & ~n191;
  assign n722 = n538 & n721;
  assign n723 = ~n570 & ~n578;
  assign n724 = ~n200 & ~n209;
  assign n725 = n723 & n724;
  assign n726 = n722 & n725;
  assign n727 = n720 & n726;
  assign n728 = ~n234 & ~n594;
  assign n729 = ~n586 & n728;
  assign n730 = ~n239 & ~n243;
  assign n731 = ~n256 & ~n263;
  assign n732 = n730 & n731;
  assign n733 = n729 & n732;
  assign n734 = ~n268 & ~n272;
  assign n735 = ~n277 & ~n281;
  assign n736 = n734 & n735;
  assign n737 = ~n289 & ~n293;
  assign n738 = n556 & n737;
  assign n739 = n736 & n738;
  assign n740 = n733 & n739;
  assign n741 = n727 & n740;
  assign po1 = n715 | ~n741;
  assign n743 = ~pi19 & ~pi20;
  assign n744 = pi28 & ~n743;
  assign n745 = ~pi21 & n744;
  assign n746 = ~pi30 & ~pi31;
  assign n747 = ~pi29 & n746;
  assign n748 = ~pi15 & ~n309;
  assign n749 = ~pi26 & ~n595;
  assign n750 = n748 & n749;
  assign n751 = ~n747 & ~n750;
  assign n752 = ~pi13 & ~n331;
  assign n753 = n333 & n752;
  assign n754 = ~pi09 & ~n753;
  assign n755 = pi01 & pi12;
  assign n756 = ~n754 & n755;
  assign n757 = ~pi06 & ~n756;
  assign n758 = ~pi05 & n757;
  assign n759 = ~pi04 & n758;
  assign n760 = ~pi02 & n759;
  assign n761 = pi29 & ~n760;
  assign n762 = ~n357 & ~n761;
  assign n763 = ~n310 & n762;
  assign n764 = ~pi07 & n763;
  assign n765 = pi37 & n764;
  assign n766 = ~n751 & ~n765;
  assign n767 = ~pi28 & ~n766;
  assign n768 = ~n363 & ~n751;
  assign n769 = pi21 & ~n768;
  assign n770 = ~n767 & ~n769;
  assign n771 = ~n745 & n770;
  assign n772 = ~n308 & ~n771;
  assign n773 = ~pi21 & pi28;
  assign n774 = ~pi33 & ~n773;
  assign n775 = pi34 & n774;
  assign n776 = ~n510 & ~n775;
  assign n777 = pi22 & ~n776;
  assign n778 = ~pi25 & ~n750;
  assign n779 = ~pi23 & n778;
  assign n780 = ~n777 & ~n779;
  assign n781 = ~n747 & ~n780;
  assign n782 = pi13 & n773;
  assign n783 = ~pi32 & ~n782;
  assign n784 = pi14 & ~n783;
  assign n785 = ~pi15 & ~pi22;
  assign n786 = n749 & n785;
  assign n787 = pi28 & ~n786;
  assign n788 = pi10 & n346;
  assign n789 = ~pi13 & n788;
  assign n790 = ~pi09 & ~n789;
  assign n791 = pi12 & ~n790;
  assign n792 = pi02 & ~n791;
  assign n793 = ~pi29 & ~n792;
  assign n794 = ~n760 & ~n793;
  assign n795 = ~n357 & ~n794;
  assign n796 = ~n310 & n795;
  assign n797 = ~n372 & n796;
  assign n798 = ~pi29 & ~n42;
  assign n799 = ~pi06 & ~n755;
  assign n800 = ~pi05 & n799;
  assign n801 = ~pi04 & n800;
  assign n802 = ~pi02 & n801;
  assign n803 = ~n798 & ~n802;
  assign n804 = ~pi13 & n346;
  assign n805 = pi10 & ~n804;
  assign n806 = ~n803 & ~n805;
  assign n807 = ~n357 & n806;
  assign n808 = ~n310 & n807;
  assign n809 = ~pi34 & n808;
  assign n810 = pi09 & n809;
  assign n811 = ~n797 & ~n810;
  assign n812 = pi37 & ~n811;
  assign n813 = ~n787 & ~n812;
  assign n814 = ~pi21 & ~n813;
  assign n815 = ~n372 & n763;
  assign n816 = pi29 & ~n802;
  assign n817 = ~n805 & ~n816;
  assign n818 = ~n357 & n817;
  assign n819 = ~n310 & n818;
  assign n820 = ~pi34 & n819;
  assign n821 = pi09 & n820;
  assign n822 = ~n815 & ~n821;
  assign n823 = ~pi28 & ~n822;
  assign n824 = pi37 & n823;
  assign n825 = ~n814 & ~n824;
  assign n826 = ~n784 & n825;
  assign n827 = ~pi25 & ~n826;
  assign n828 = pi22 & ~n773;
  assign n829 = pi09 & ~n805;
  assign n830 = pi30 & ~n829;
  assign n831 = ~n755 & ~n830;
  assign n832 = ~pi30 & ~n753;
  assign n833 = ~pi09 & n832;
  assign n834 = ~n831 & ~n833;
  assign n835 = ~pi06 & ~n834;
  assign n836 = ~pi05 & n835;
  assign n837 = ~pi04 & n836;
  assign n838 = ~pi02 & n837;
  assign n839 = ~pi29 & ~n830;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n357 & ~n840;
  assign n842 = ~n310 & n841;
  assign n843 = ~pi28 & n842;
  assign n844 = pi37 & n843;
  assign n845 = ~pi34 & n844;
  assign n846 = ~n828 & ~n845;
  assign n847 = pi33 & ~n846;
  assign n848 = ~n827 & ~n847;
  assign n849 = ~pi23 & ~n848;
  assign n850 = ~n781 & ~n849;
  assign n851 = ~n772 & n850;
  assign n852 = ~pi27 & ~n851;
  assign n853 = ~n100 & ~n111;
  assign n854 = ~n91 & n853;
  assign n855 = ~n141 & ~n570;
  assign n856 = n531 & n855;
  assign n857 = n854 & n856;
  assign n858 = ~n217 & ~n586;
  assign n859 = ~n578 & n858;
  assign n860 = ~n223 & ~n594;
  assign n861 = ~n229 & ~n252;
  assign n862 = n860 & n861;
  assign n863 = n859 & n862;
  assign n864 = n857 & n863;
  assign po2 = n852 | ~n864;
endmodule



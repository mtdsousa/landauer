// Benchmark "vda" written by ABC on Sun Apr 22 21:43:15 2018

module vda ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38;
  wire n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n309, n310, n311, n312, n313, n314, n315, n316,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n341, n342,
    n343, n344, n345, n346, n347, n348, n350, n351, n352, n353, n354, n355,
    n356, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n412, n413, n414, n417, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n681, n682, n683, n684, n685, n686, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n769, n770, n771, n772, n773, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n952, n953, n955, n956, n957, n958, n959, n960,
    n961, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978;
  assign n57 = pi01 & pi04;
  assign n58 = pi07 & n57;
  assign n59 = ~pi08 & n58;
  assign n60 = pi09 & n59;
  assign n61 = ~pi11 & n60;
  assign n62 = pi12 & n61;
  assign n63 = pi13 & n62;
  assign n64 = pi14 & n63;
  assign n65 = pi15 & n64;
  assign n66 = ~pi16 & n65;
  assign n67 = ~pi02 & pi04;
  assign n68 = pi07 & n67;
  assign n69 = ~pi08 & n68;
  assign n70 = pi09 & n69;
  assign n71 = ~pi11 & n70;
  assign n72 = pi12 & n71;
  assign n73 = pi13 & n72;
  assign n74 = pi14 & n73;
  assign n75 = pi15 & n74;
  assign n76 = ~pi16 & n75;
  assign n77 = pi04 & ~pi05;
  assign n78 = pi07 & n77;
  assign n79 = ~pi08 & n78;
  assign n80 = pi09 & n79;
  assign n81 = ~pi11 & n80;
  assign n82 = pi12 & n81;
  assign n83 = pi13 & n82;
  assign n84 = pi14 & n83;
  assign n85 = pi15 & n84;
  assign n86 = ~pi16 & n85;
  assign n87 = pi00 & pi04;
  assign n88 = pi11 & n87;
  assign n89 = ~pi12 & n88;
  assign n90 = ~pi13 & n89;
  assign n91 = pi14 & n90;
  assign n92 = ~pi15 & n91;
  assign n93 = ~pi16 & n92;
  assign n94 = ~pi11 & n57;
  assign n95 = ~pi12 & n94;
  assign n96 = ~pi13 & n95;
  assign n97 = ~pi14 & n96;
  assign n98 = pi15 & n97;
  assign n99 = pi16 & n98;
  assign n100 = ~pi11 & n77;
  assign n101 = ~pi12 & n100;
  assign n102 = ~pi13 & n101;
  assign n103 = ~pi14 & n102;
  assign n104 = pi15 & n103;
  assign n105 = pi16 & n104;
  assign n106 = pi02 & ~pi11;
  assign n107 = ~pi12 & n106;
  assign n108 = ~pi13 & n107;
  assign n109 = ~pi14 & n108;
  assign n110 = ~pi15 & n109;
  assign n111 = pi16 & n110;
  assign n112 = pi05 & ~pi11;
  assign n113 = ~pi12 & n112;
  assign n114 = pi13 & n113;
  assign n115 = ~pi14 & n114;
  assign n116 = pi15 & n115;
  assign n117 = ~pi16 & n116;
  assign n118 = pi06 & pi11;
  assign n119 = ~pi12 & n118;
  assign n120 = ~pi13 & n119;
  assign n121 = pi14 & n120;
  assign n122 = pi15 & n121;
  assign n123 = pi16 & n122;
  assign n124 = ~pi05 & ~pi11;
  assign n125 = ~pi12 & n124;
  assign n126 = pi13 & n125;
  assign n127 = ~pi14 & n126;
  assign n128 = pi15 & n127;
  assign n129 = ~pi16 & n128;
  assign n130 = ~pi11 & ~pi12;
  assign n131 = ~pi13 & n130;
  assign n132 = pi14 & n131;
  assign n133 = ~pi15 & n132;
  assign n134 = pi16 & n133;
  assign n135 = ~pi14 & n131;
  assign n136 = pi15 & n135;
  assign n137 = ~pi16 & n136;
  assign n138 = pi13 & n130;
  assign n139 = ~pi14 & n138;
  assign n140 = ~pi15 & n139;
  assign n141 = ~pi16 & n140;
  assign n142 = pi06 & ~pi11;
  assign n143 = pi12 & n142;
  assign n144 = ~pi13 & n143;
  assign n145 = pi14 & n144;
  assign n146 = ~pi15 & n145;
  assign n147 = ~pi16 & n146;
  assign n148 = pi11 & ~pi12;
  assign n149 = ~pi13 & n148;
  assign n150 = ~pi14 & n149;
  assign n151 = pi15 & n150;
  assign n152 = ~pi16 & n151;
  assign n153 = ~pi01 & pi05;
  assign n154 = ~pi11 & n153;
  assign n155 = ~pi12 & n154;
  assign n156 = ~pi13 & n155;
  assign n157 = ~pi14 & n156;
  assign n158 = pi15 & n157;
  assign n159 = pi16 & n158;
  assign n160 = ~pi12 & n142;
  assign n161 = pi13 & n160;
  assign n162 = pi14 & n161;
  assign n163 = pi15 & n162;
  assign n164 = pi16 & n163;
  assign n165 = ~pi06 & pi11;
  assign n166 = ~pi12 & n165;
  assign n167 = ~pi13 & n166;
  assign n168 = pi14 & n167;
  assign n169 = pi15 & n168;
  assign n170 = pi16 & n169;
  assign n171 = pi15 & n132;
  assign n172 = ~pi16 & n171;
  assign n173 = ~pi16 & n133;
  assign n174 = pi14 & n138;
  assign n175 = ~pi15 & n174;
  assign n176 = ~pi16 & n175;
  assign n177 = pi08 & ~pi11;
  assign n178 = ~pi12 & n177;
  assign n179 = pi13 & n178;
  assign n180 = ~pi14 & n179;
  assign n181 = pi15 & n180;
  assign n182 = pi16 & n181;
  assign n183 = ~pi11 & pi12;
  assign n184 = ~pi13 & n183;
  assign n185 = ~pi14 & n184;
  assign n186 = ~pi15 & n185;
  assign n187 = ~pi16 & n186;
  assign n188 = pi14 & n149;
  assign n189 = pi15 & n188;
  assign n190 = ~pi16 & n189;
  assign n191 = pi14 & n184;
  assign n192 = pi15 & n191;
  assign n193 = pi16 & n192;
  assign n194 = pi16 & n175;
  assign n195 = ~pi06 & ~pi11;
  assign n196 = pi12 & n195;
  assign n197 = pi13 & n196;
  assign n198 = ~pi14 & n197;
  assign n199 = pi15 & n198;
  assign n200 = pi16 & n199;
  assign n201 = pi11 & pi12;
  assign n202 = pi13 & n201;
  assign n203 = ~pi14 & n202;
  assign n204 = pi15 & n203;
  assign n205 = pi16 & n204;
  assign n206 = ~pi15 & n188;
  assign n207 = pi16 & n206;
  assign n208 = ~pi15 & n203;
  assign n209 = ~pi16 & n208;
  assign n210 = ~pi13 & n196;
  assign n211 = pi14 & n210;
  assign n212 = pi15 & n211;
  assign n213 = ~pi16 & n212;
  assign n214 = ~pi13 & n201;
  assign n215 = ~pi14 & n214;
  assign n216 = pi15 & n215;
  assign n217 = pi16 & n216;
  assign n218 = pi14 & n214;
  assign n219 = ~pi15 & n218;
  assign n220 = ~pi16 & n219;
  assign n221 = ~n217 & ~n220;
  assign n222 = ~n209 & ~n213;
  assign n223 = n221 & n222;
  assign n224 = ~n205 & ~n207;
  assign n225 = ~n194 & ~n200;
  assign n226 = n224 & n225;
  assign n227 = n223 & n226;
  assign n228 = ~n190 & ~n193;
  assign n229 = ~n182 & ~n187;
  assign n230 = n228 & n229;
  assign n231 = ~n173 & ~n176;
  assign n232 = ~n170 & ~n172;
  assign n233 = n231 & n232;
  assign n234 = n230 & n233;
  assign n235 = n227 & n234;
  assign n236 = ~n159 & ~n164;
  assign n237 = ~n147 & ~n152;
  assign n238 = n236 & n237;
  assign n239 = ~n137 & ~n141;
  assign n240 = ~n129 & ~n134;
  assign n241 = n239 & n240;
  assign n242 = n238 & n241;
  assign n243 = ~n117 & ~n123;
  assign n244 = ~n105 & ~n111;
  assign n245 = n243 & n244;
  assign n246 = ~n93 & ~n99;
  assign n247 = ~n66 & ~n76;
  assign n248 = ~n86 & n247;
  assign n249 = n246 & n248;
  assign n250 = n245 & n249;
  assign n251 = n242 & n250;
  assign po00 = ~n235 | ~n251;
  assign n253 = pi00 & ~pi04;
  assign n254 = ~pi05 & n253;
  assign n255 = pi11 & n254;
  assign n256 = ~pi12 & n255;
  assign n257 = ~pi13 & n256;
  assign n258 = pi14 & n257;
  assign n259 = ~pi15 & n258;
  assign n260 = ~pi16 & n259;
  assign n261 = pi01 & ~pi04;
  assign n262 = ~pi08 & n261;
  assign n263 = ~pi11 & n262;
  assign n264 = pi12 & n263;
  assign n265 = pi13 & n264;
  assign n266 = pi14 & n265;
  assign n267 = pi15 & n266;
  assign n268 = ~pi16 & n267;
  assign n269 = ~pi02 & ~pi04;
  assign n270 = ~pi08 & n269;
  assign n271 = ~pi11 & n270;
  assign n272 = pi12 & n271;
  assign n273 = pi13 & n272;
  assign n274 = pi14 & n273;
  assign n275 = pi15 & n274;
  assign n276 = ~pi16 & n275;
  assign n277 = ~pi04 & ~pi05;
  assign n278 = ~pi08 & n277;
  assign n279 = ~pi11 & n278;
  assign n280 = pi12 & n279;
  assign n281 = pi13 & n280;
  assign n282 = pi14 & n281;
  assign n283 = pi15 & n282;
  assign n284 = ~pi16 & n283;
  assign n285 = ~pi12 & n277;
  assign n286 = ~pi13 & n285;
  assign n287 = ~pi14 & n286;
  assign n288 = pi15 & n287;
  assign n289 = pi16 & n288;
  assign n290 = ~pi07 & ~pi08;
  assign n291 = ~pi11 & n290;
  assign n292 = pi12 & n291;
  assign n293 = pi13 & n292;
  assign n294 = pi14 & n293;
  assign n295 = ~pi16 & n294;
  assign n296 = ~pi07 & ~pi11;
  assign n297 = pi12 & n296;
  assign n298 = pi13 & n297;
  assign n299 = pi14 & n298;
  assign n300 = ~pi15 & n299;
  assign n301 = ~pi16 & n300;
  assign n302 = ~pi15 & n135;
  assign n303 = ~pi16 & n302;
  assign n304 = pi13 & n148;
  assign n305 = pi14 & n304;
  assign n306 = pi15 & n305;
  assign n307 = ~pi16 & n306;
  assign po35 = pi16 & n151;
  assign n309 = ~n284 & ~n289;
  assign n310 = ~n260 & ~n268;
  assign n311 = ~n276 & n310;
  assign n312 = n309 & n311;
  assign n313 = ~n307 & ~po35;
  assign n314 = ~n295 & ~n301;
  assign n315 = ~n303 & n314;
  assign n316 = n313 & n315;
  assign po01 = ~n312 | ~n316;
  assign n318 = ~n213 & ~n217;
  assign n319 = ~n220 & n318;
  assign n320 = ~n209 & n224;
  assign n321 = n319 & n320;
  assign n322 = ~n193 & ~n194;
  assign n323 = ~n200 & n322;
  assign n324 = ~n187 & ~n190;
  assign n325 = ~n176 & ~n182;
  assign n326 = n324 & n325;
  assign n327 = n323 & n326;
  assign n328 = n321 & n327;
  assign n329 = ~n173 & n232;
  assign n330 = ~n152 & ~n159;
  assign n331 = ~n134 & ~n137;
  assign n332 = n330 & n331;
  assign n333 = n329 & n332;
  assign n334 = ~n99 & ~n105;
  assign n335 = ~n111 & n334;
  assign n336 = ~n86 & ~n93;
  assign n337 = n247 & n336;
  assign n338 = n335 & n337;
  assign n339 = n333 & n338;
  assign po02 = ~n328 | ~n339;
  assign n341 = ~pi14 & n304;
  assign n342 = ~pi15 & n341;
  assign n343 = pi16 & n342;
  assign n344 = pi16 & n306;
  assign n345 = pi13 & n183;
  assign n346 = ~pi14 & n345;
  assign n347 = ~pi15 & n346;
  assign n348 = pi16 & n347;
  assign po11 = pi16 & n140;
  assign n350 = pi16 & n219;
  assign n351 = pi15 & n185;
  assign n352 = ~pi16 & n351;
  assign n353 = ~n343 & ~n344;
  assign n354 = ~n348 & n353;
  assign n355 = ~po11 & ~n350;
  assign n356 = ~n352 & n355;
  assign po03 = ~n354 | ~n356;
  assign n358 = ~pi03 & ~pi08;
  assign n359 = ~pi11 & n358;
  assign n360 = ~pi12 & n359;
  assign n361 = pi13 & n360;
  assign n362 = ~pi14 & n361;
  assign n363 = pi15 & n362;
  assign n364 = pi16 & n363;
  assign n365 = ~pi10 & ~pi11;
  assign n366 = ~pi12 & n365;
  assign n367 = ~pi13 & n366;
  assign n368 = pi14 & n367;
  assign n369 = pi15 & n368;
  assign po10 = pi16 & n369;
  assign n371 = pi03 & ~pi08;
  assign n372 = ~pi11 & n371;
  assign n373 = ~pi12 & n372;
  assign n374 = pi13 & n373;
  assign n375 = ~pi14 & n374;
  assign n376 = pi15 & n375;
  assign n377 = pi16 & n376;
  assign n378 = pi06 & pi10;
  assign n379 = ~pi11 & n378;
  assign n380 = pi12 & n379;
  assign n381 = ~pi13 & n380;
  assign n382 = pi14 & n381;
  assign n383 = pi15 & n382;
  assign n384 = ~pi16 & n383;
  assign n385 = pi06 & pi08;
  assign n386 = ~pi11 & n385;
  assign n387 = pi12 & n386;
  assign n388 = ~pi13 & n387;
  assign n389 = pi14 & n388;
  assign n390 = pi15 & n389;
  assign n391 = ~pi16 & n390;
  assign n392 = pi02 & pi06;
  assign n393 = ~pi11 & n392;
  assign n394 = pi12 & n393;
  assign n395 = ~pi13 & n394;
  assign n396 = pi14 & n395;
  assign n397 = pi15 & n396;
  assign n398 = ~pi16 & n397;
  assign n399 = ~n164 & ~n352;
  assign n400 = ~n141 & ~n147;
  assign n401 = n399 & n400;
  assign n402 = ~n123 & ~n348;
  assign n403 = n355 & n402;
  assign n404 = n401 & n403;
  assign n405 = ~n364 & ~po10;
  assign n406 = ~n377 & ~n384;
  assign n407 = n405 & n406;
  assign n408 = ~n391 & ~n398;
  assign n409 = n353 & n408;
  assign n410 = n407 & n409;
  assign po04 = ~n404 | ~n410;
  assign n412 = ~n147 & ~n164;
  assign n413 = ~n352 & n412;
  assign n414 = n403 & n413;
  assign po07 = ~n410 | ~n414;
  assign po08 = n172 | n173;
  assign n417 = ~po11 & ~po10;
  assign po09 = ~n412 | ~n417;
  assign n419 = ~pi01 & pi02;
  assign n420 = pi05 & n419;
  assign n421 = pi07 & n420;
  assign n422 = ~pi08 & n421;
  assign n423 = ~pi11 & n422;
  assign n424 = pi12 & n423;
  assign n425 = pi13 & n424;
  assign n426 = pi14 & n425;
  assign n427 = pi15 & n426;
  assign n428 = ~pi16 & n427;
  assign n429 = pi10 & ~pi11;
  assign n430 = ~pi12 & n429;
  assign n431 = ~pi13 & n430;
  assign n432 = pi14 & n431;
  assign n433 = pi15 & n432;
  assign n434 = pi16 & n433;
  assign n435 = ~pi00 & pi11;
  assign n436 = ~pi13 & n435;
  assign n437 = pi14 & n436;
  assign n438 = ~pi15 & n437;
  assign n439 = ~pi16 & n342;
  assign n440 = ~pi15 & n150;
  assign po34 = pi16 & n440;
  assign n442 = ~pi15 & n191;
  assign n443 = pi16 & n442;
  assign n444 = ~pi15 & n215;
  assign n445 = pi16 & n444;
  assign n446 = ~pi16 & n215;
  assign n447 = pi14 & n202;
  assign n448 = ~pi15 & n447;
  assign n449 = ~pi16 & n448;
  assign n450 = pi15 & n214;
  assign n451 = ~pi16 & n450;
  assign n452 = pi16 & n351;
  assign po38 = pi16 & n208;
  assign n454 = ~pi16 & n440;
  assign n455 = ~pi16 & n174;
  assign n456 = ~n207 & ~n209;
  assign n457 = n221 & n456;
  assign n458 = ~n170 & ~n190;
  assign n459 = ~n152 & ~n350;
  assign n460 = ~n159 & n459;
  assign n461 = n458 & n460;
  assign n462 = n457 & n461;
  assign n463 = ~n123 & ~n455;
  assign n464 = ~po35 & ~n454;
  assign n465 = ~n344 & n464;
  assign n466 = n463 & n465;
  assign n467 = ~n452 & ~po38;
  assign n468 = ~n449 & ~n451;
  assign n469 = ~n307 & n468;
  assign n470 = n467 & n469;
  assign n471 = n466 & n470;
  assign n472 = n462 & n471;
  assign n473 = ~n445 & ~n446;
  assign n474 = ~po34 & ~n443;
  assign n475 = n473 & n474;
  assign n476 = ~n301 & ~n439;
  assign n477 = ~n295 & ~n434;
  assign n478 = ~n438 & n477;
  assign n479 = n476 & n478;
  assign n480 = n475 & n479;
  assign n481 = ~n86 & ~n268;
  assign n482 = ~n276 & n481;
  assign n483 = n309 & n482;
  assign n484 = pi12 & pi13;
  assign n485 = pi15 & ~pi16;
  assign n486 = ~pi14 & n485;
  assign n487 = n484 & n486;
  assign n488 = ~n428 & ~n487;
  assign n489 = ~n260 & n488;
  assign n490 = n247 & n489;
  assign n491 = n483 & n490;
  assign n492 = n480 & n491;
  assign po12 = ~n472 | ~n492;
  assign n494 = ~pi02 & pi06;
  assign n495 = ~pi08 & n494;
  assign n496 = ~pi10 & n495;
  assign n497 = ~pi11 & n496;
  assign n498 = pi12 & n497;
  assign n499 = ~pi13 & n498;
  assign n500 = pi14 & n499;
  assign n501 = pi15 & n500;
  assign n502 = ~pi16 & n501;
  assign n503 = ~pi09 & n58;
  assign n504 = ~pi11 & n503;
  assign n505 = pi12 & n504;
  assign n506 = pi13 & n505;
  assign n507 = pi14 & n506;
  assign n508 = pi15 & n507;
  assign n509 = ~pi09 & n68;
  assign n510 = ~pi11 & n509;
  assign n511 = pi12 & n510;
  assign n512 = pi13 & n511;
  assign n513 = pi14 & n512;
  assign n514 = pi15 & n513;
  assign n515 = ~pi09 & n78;
  assign n516 = ~pi11 & n515;
  assign n517 = pi12 & n516;
  assign n518 = pi13 & n517;
  assign n519 = pi14 & n518;
  assign n520 = pi15 & n519;
  assign n521 = ~pi15 & n211;
  assign n522 = ~pi16 & n521;
  assign n523 = pi07 & ~pi11;
  assign n524 = pi12 & n523;
  assign n525 = pi13 & n524;
  assign n526 = pi14 & n525;
  assign n527 = ~pi15 & n526;
  assign n528 = ~pi16 & n527;
  assign n529 = ~pi15 & n304;
  assign n530 = pi16 & n529;
  assign n531 = pi13 & n143;
  assign n532 = pi15 & n531;
  assign n533 = pi16 & n532;
  assign n534 = pi13 & n195;
  assign n535 = pi14 & n534;
  assign n536 = pi15 & n535;
  assign n537 = pi16 & n536;
  assign n538 = ~pi16 & n347;
  assign n539 = ~pi14 & n183;
  assign n540 = ~pi15 & n539;
  assign n541 = pi16 & n540;
  assign n542 = pi15 & n341;
  assign n543 = ~pi16 & n542;
  assign n544 = pi12 & n177;
  assign n545 = pi13 & n544;
  assign n546 = pi14 & n545;
  assign n547 = pi15 & n546;
  assign n548 = ~pi16 & n547;
  assign n549 = ~pi12 & pi13;
  assign n550 = pi14 & n549;
  assign n551 = ~pi15 & n550;
  assign n552 = ~pi16 & n551;
  assign n553 = ~n364 & ~n548;
  assign n554 = ~n446 & ~n543;
  assign n555 = n553 & n554;
  assign n556 = ~n538 & ~n541;
  assign n557 = ~n533 & ~n537;
  assign n558 = n556 & n557;
  assign n559 = n555 & n558;
  assign n560 = ~n528 & ~n530;
  assign n561 = ~n434 & ~n522;
  assign n562 = n560 & n561;
  assign n563 = ~n514 & ~n520;
  assign n564 = ~n428 & ~n502;
  assign n565 = ~n508 & n564;
  assign n566 = n563 & n565;
  assign n567 = n562 & n566;
  assign n568 = n559 & n567;
  assign n569 = ~n200 & ~n209;
  assign n570 = n318 & n569;
  assign n571 = ~n187 & ~n193;
  assign n572 = ~n170 & ~n352;
  assign n573 = n571 & n572;
  assign n574 = n570 & n573;
  assign n575 = ~n129 & ~n350;
  assign n576 = n412 & n575;
  assign n577 = ~po35 & ~n344;
  assign n578 = ~n451 & ~n552;
  assign n579 = ~po38 & n578;
  assign n580 = n577 & n579;
  assign n581 = n576 & n580;
  assign n582 = n574 & n581;
  assign po13 = ~n568 | ~n582;
  assign n584 = pi05 & n261;
  assign n585 = ~pi11 & n584;
  assign n586 = ~pi12 & n585;
  assign n587 = ~pi13 & n586;
  assign n588 = ~pi14 & n587;
  assign n589 = pi15 & n588;
  assign n590 = pi16 & n589;
  assign n591 = pi05 & n253;
  assign n592 = pi11 & n591;
  assign n593 = ~pi12 & n592;
  assign n594 = ~pi13 & n593;
  assign n595 = pi14 & n594;
  assign n596 = ~pi16 & n595;
  assign n597 = pi15 & n346;
  assign n598 = ~pi16 & n597;
  assign n599 = pi16 & n542;
  assign n600 = ~n205 & ~n220;
  assign n601 = ~n194 & n228;
  assign n602 = n600 & n601;
  assign n603 = ~n170 & ~n182;
  assign n604 = ~n129 & ~po11;
  assign n605 = ~n141 & n604;
  assign n606 = n603 & n605;
  assign n607 = n602 & n606;
  assign n608 = ~n117 & ~n454;
  assign n609 = ~n455 & n608;
  assign n610 = n402 & n609;
  assign n611 = ~po35 & ~po38;
  assign n612 = n408 & ~n552;
  assign n613 = n611 & n612;
  assign n614 = n610 & n613;
  assign n615 = n607 & n614;
  assign n616 = ~po10 & ~n599;
  assign n617 = ~n452 & n616;
  assign n618 = n406 & n617;
  assign n619 = ~n443 & ~n548;
  assign n620 = ~n537 & ~n598;
  assign n621 = ~n538 & n620;
  assign n622 = n619 & n621;
  assign n623 = n618 & n622;
  assign n624 = n564 & ~n590;
  assign n625 = ~n508 & ~n596;
  assign n626 = ~n514 & n625;
  assign n627 = n624 & n626;
  assign n628 = ~n439 & ~n533;
  assign n629 = ~n520 & ~n522;
  assign n630 = ~n528 & n629;
  assign n631 = n628 & n630;
  assign n632 = n627 & n631;
  assign n633 = n623 & n632;
  assign po14 = ~n615 | ~n633;
  assign n635 = pi15 & n218;
  assign n636 = ~n200 & ~n205;
  assign n637 = ~n207 & n636;
  assign n638 = n319 & n637;
  assign n639 = ~n173 & ~n182;
  assign n640 = ~n190 & n639;
  assign n641 = ~n159 & ~n350;
  assign n642 = ~n172 & n641;
  assign n643 = n640 & n642;
  assign n644 = n638 & n643;
  assign n645 = ~n129 & ~n454;
  assign n646 = ~n134 & n645;
  assign n647 = ~po35 & n408;
  assign n648 = n646 & n647;
  assign n649 = ~n307 & ~n452;
  assign n650 = ~n364 & ~n451;
  assign n651 = n649 & n650;
  assign n652 = ~n377 & ~n635;
  assign n653 = ~n384 & n652;
  assign n654 = n651 & n653;
  assign n655 = n648 & n654;
  assign n656 = n644 & n655;
  assign n657 = ~n105 & ~n548;
  assign n658 = ~n599 & n657;
  assign n659 = ~n445 & ~n449;
  assign n660 = ~n99 & n659;
  assign n661 = n658 & n660;
  assign n662 = ~n301 & ~n530;
  assign n663 = n557 & n662;
  assign n664 = ~n93 & ~n598;
  assign n665 = ~n543 & n664;
  assign n666 = n663 & n665;
  assign n667 = n661 & n666;
  assign n668 = ~n268 & ~n520;
  assign n669 = ~n276 & n668;
  assign n670 = ~n260 & ~n502;
  assign n671 = ~n508 & ~n514;
  assign n672 = n670 & n671;
  assign n673 = n669 & n672;
  assign n674 = ~n295 & ~n528;
  assign n675 = ~n438 & n674;
  assign n676 = n309 & ~n522;
  assign n677 = n675 & n676;
  assign n678 = n673 & n677;
  assign n679 = n667 & n678;
  assign po15 = ~n656 | ~n679;
  assign n681 = pi07 & pi09;
  assign n682 = ~pi11 & n681;
  assign n683 = pi12 & n682;
  assign n684 = pi13 & n683;
  assign n685 = pi14 & n684;
  assign n686 = ~pi15 & n685;
  assign po36 = ~pi16 & n686;
  assign n688 = pi14 & n345;
  assign n689 = pi15 & n688;
  assign n690 = pi16 & n689;
  assign n691 = ~n213 & ~n220;
  assign n692 = ~n200 & ~n207;
  assign n693 = ~n209 & n692;
  assign n694 = n691 & n693;
  assign n695 = ~n190 & ~n194;
  assign n696 = ~n152 & ~n352;
  assign n697 = ~n172 & n696;
  assign n698 = n695 & n697;
  assign n699 = n694 & n698;
  assign n700 = ~n398 & ~n552;
  assign n701 = ~po38 & n700;
  assign n702 = n609 & n701;
  assign n703 = ~n137 & ~n350;
  assign n704 = ~n134 & n604;
  assign n705 = n703 & n704;
  assign n706 = n702 & n705;
  assign n707 = n699 & n706;
  assign n708 = ~n384 & ~n391;
  assign n709 = ~n111 & ~n635;
  assign n710 = ~n377 & n709;
  assign n711 = n708 & n710;
  assign n712 = ~n445 & n474;
  assign n713 = ~n548 & ~n690;
  assign n714 = ~n599 & n713;
  assign n715 = n712 & n714;
  assign n716 = n711 & n715;
  assign n717 = ~n541 & ~n543;
  assign n718 = ~n520 & ~po36;
  assign n719 = ~n434 & n718;
  assign n720 = n717 & n719;
  assign n721 = ~pi02 & ~pi06;
  assign n722 = ~pi08 & ~pi11;
  assign n723 = n721 & n722;
  assign n724 = pi13 & pi14;
  assign n725 = pi15 & pi16;
  assign n726 = n724 & n725;
  assign n727 = n723 & n726;
  assign n728 = ~n502 & ~n727;
  assign n729 = ~n590 & n728;
  assign n730 = n626 & n729;
  assign n731 = n720 & n730;
  assign n732 = n716 & n731;
  assign po16 = ~n707 | ~n732;
  assign n734 = ~n172 & ~n352;
  assign n735 = n330 & n734;
  assign n736 = ~n117 & ~n343;
  assign n737 = ~n455 & n736;
  assign n738 = n239 & n737;
  assign n739 = n735 & n738;
  assign n740 = ~n173 & ~n187;
  assign n741 = ~n190 & n740;
  assign n742 = n225 & n741;
  assign n743 = ~n205 & ~n209;
  assign n744 = n691 & n743;
  assign n745 = n742 & n744;
  assign n746 = n739 & n745;
  assign n747 = ~n552 & ~n635;
  assign n748 = ~n364 & ~n452;
  assign n749 = n747 & n748;
  assign n750 = ~n548 & ~n599;
  assign n751 = ~n445 & ~n538;
  assign n752 = ~n446 & n751;
  assign n753 = n750 & n752;
  assign n754 = n749 & n753;
  assign n755 = ~n76 & ~n86;
  assign n756 = ~n303 & ~n439;
  assign n757 = n755 & n756;
  assign n758 = ~n66 & ~n596;
  assign n759 = ~pi02 & n130;
  assign n760 = ~pi14 & ~pi15;
  assign n761 = ~pi13 & n760;
  assign n762 = n759 & n761;
  assign n763 = ~n428 & ~n762;
  assign n764 = ~n590 & n763;
  assign n765 = n758 & n764;
  assign n766 = n757 & n765;
  assign n767 = n754 & n766;
  assign po17 = ~n746 | ~n767;
  assign n769 = ~n307 & ~n449;
  assign n770 = ~n301 & ~n303;
  assign n771 = n769 & n770;
  assign n772 = ~n284 & ~n295;
  assign n773 = n311 & n772;
  assign po18 = ~n771 | ~n773;
  assign n775 = ~n276 & ~n284;
  assign n776 = n310 & n775;
  assign n777 = ~n295 & ~po36;
  assign n778 = n770 & n777;
  assign n779 = n776 & n778;
  assign n780 = ~n449 & ~n690;
  assign n781 = ~n307 & ~po38;
  assign n782 = n780 & n781;
  assign n783 = ~n123 & ~n454;
  assign n784 = ~n147 & n783;
  assign n785 = n782 & n784;
  assign n786 = n779 & n785;
  assign n787 = n456 & n636;
  assign n788 = n319 & n787;
  assign n789 = n229 & n322;
  assign n790 = ~n170 & ~n176;
  assign n791 = n236 & n790;
  assign n792 = n789 & n791;
  assign n793 = n788 & n792;
  assign po19 = ~n786 | ~n793;
  assign n795 = ~n200 & n228;
  assign n796 = n229 & n231;
  assign n797 = n795 & n796;
  assign n798 = n321 & n797;
  assign n799 = ~n172 & n412;
  assign n800 = n239 & n604;
  assign n801 = n799 & n800;
  assign n802 = ~n117 & n611;
  assign n803 = ~po34 & ~po36;
  assign n804 = ~n111 & ~po10;
  assign n805 = n803 & n804;
  assign n806 = n802 & n805;
  assign n807 = n801 & n806;
  assign po20 = ~n798 | ~n807;
  assign n809 = ~n111 & ~n690;
  assign n810 = ~n105 & n246;
  assign n811 = n809 & n810;
  assign n812 = ~n137 & ~n159;
  assign n813 = ~n134 & n783;
  assign n814 = n812 & n813;
  assign n815 = n811 & n814;
  assign n816 = ~n207 & n225;
  assign n817 = n691 & n816;
  assign n818 = ~n176 & ~n187;
  assign n819 = n329 & n818;
  assign n820 = n817 & n819;
  assign po21 = ~n815 | ~n820;
  assign n822 = ~po10 & ~n690;
  assign n823 = n803 & n822;
  assign n824 = n608 & n611;
  assign n825 = n823 & n824;
  assign n826 = ~n123 & ~po11;
  assign n827 = ~n129 & ~n141;
  assign n828 = n826 & n827;
  assign n829 = ~n147 & ~n159;
  assign n830 = ~n164 & n829;
  assign n831 = n828 & n830;
  assign n832 = n825 & n831;
  assign n833 = n229 & n790;
  assign n834 = n601 & n833;
  assign n835 = n788 & n834;
  assign po22 = ~n832 | ~n835;
  assign n837 = ~n217 & n228;
  assign n838 = ~n164 & ~n173;
  assign n839 = ~n182 & n838;
  assign n840 = n837 & n839;
  assign n841 = ~n111 & ~n141;
  assign n842 = ~n147 & n841;
  assign n843 = ~n307 & ~po10;
  assign n844 = n334 & n843;
  assign n845 = n842 & n844;
  assign n846 = n840 & n845;
  assign n847 = ~n93 & ~po34;
  assign n848 = ~n449 & n847;
  assign n849 = n778 & n848;
  assign n850 = ~n268 & ~n276;
  assign n851 = ~n284 & n850;
  assign n852 = ~n66 & ~n260;
  assign n853 = n755 & n852;
  assign n854 = n851 & n853;
  assign n855 = n849 & n854;
  assign po23 = ~n846 | ~n855;
  assign n857 = n323 & n833;
  assign n858 = n321 & n857;
  assign n859 = ~n343 & ~n398;
  assign n860 = ~n344 & n859;
  assign n861 = ~n364 & ~n377;
  assign n862 = n708 & n861;
  assign n863 = n860 & n862;
  assign n864 = n236 & ~n352;
  assign n865 = ~n147 & n402;
  assign n866 = n864 & n865;
  assign n867 = n863 & n866;
  assign po24 = ~n858 | ~n867;
  assign n869 = n400 & n575;
  assign n870 = ~n348 & ~po11;
  assign n871 = n736 & n870;
  assign n872 = n869 & n871;
  assign n873 = n406 & n408;
  assign n874 = n248 & n405;
  assign n875 = n873 & n874;
  assign n876 = n872 & n875;
  assign n877 = ~n193 & ~n200;
  assign n878 = n224 & n877;
  assign n879 = n223 & n878;
  assign n880 = ~n164 & n330;
  assign n881 = n734 & n880;
  assign n882 = n796 & n881;
  assign n883 = n879 & n882;
  assign po25 = ~n876 | ~n883;
  assign n885 = ~n200 & ~n213;
  assign n886 = ~n220 & n885;
  assign n887 = ~n176 & ~n193;
  assign n888 = ~n194 & n887;
  assign n889 = n886 & n888;
  assign n890 = ~n134 & ~n350;
  assign n891 = ~n141 & n890;
  assign n892 = n329 & n891;
  assign n893 = n889 & n892;
  assign n894 = ~n343 & n405;
  assign n895 = n810 & n894;
  assign n896 = ~n129 & n870;
  assign n897 = ~n117 & ~n344;
  assign n898 = ~n123 & n897;
  assign n899 = n896 & n898;
  assign n900 = n895 & n899;
  assign po26 = ~n893 | ~n900;
  assign n902 = ~n86 & ~n364;
  assign n903 = n247 & n902;
  assign n904 = n873 & n903;
  assign n905 = n353 & n402;
  assign n906 = ~n159 & n237;
  assign n907 = n905 & n906;
  assign n908 = n904 & n907;
  assign n909 = n399 & n790;
  assign n910 = n789 & n909;
  assign n911 = n788 & n910;
  assign po27 = ~n908 | ~n911;
  assign n913 = n248 & n810;
  assign n914 = ~n398 & n708;
  assign n915 = ~n377 & n804;
  assign n916 = n914 & n915;
  assign n917 = n913 & n916;
  assign n918 = ~n207 & ~n217;
  assign n919 = ~n190 & n229;
  assign n920 = n918 & n919;
  assign n921 = ~n141 & ~n350;
  assign n922 = ~n147 & n921;
  assign n923 = ~n173 & n399;
  assign n924 = n922 & n923;
  assign n925 = n920 & n924;
  assign po28 = ~n917 | ~n925;
  assign n927 = ~n123 & ~n344;
  assign n928 = ~n137 & n927;
  assign n929 = ~n86 & ~n111;
  assign n930 = n247 & n929;
  assign n931 = n928 & n930;
  assign n932 = ~n164 & ~n170;
  assign n933 = ~n176 & n932;
  assign n934 = n906 & n933;
  assign n935 = n931 & n934;
  assign n936 = n323 & n919;
  assign n937 = n321 & n936;
  assign po29 = ~n935 | ~n937;
  assign n939 = n222 & n637;
  assign n940 = ~n173 & ~n194;
  assign n941 = ~n172 & n572;
  assign n942 = n940 & n941;
  assign n943 = n939 & n942;
  assign n944 = ~n384 & n861;
  assign n945 = ~n343 & n408;
  assign n946 = n944 & n945;
  assign n947 = ~n348 & ~n350;
  assign n948 = ~n147 & n947;
  assign n949 = n236 & n948;
  assign n950 = n946 & n949;
  assign po30 = ~n943 | ~n950;
  assign n952 = n221 & n325;
  assign n953 = n810 & n890;
  assign po31 = ~n952 | ~n953;
  assign n955 = ~n134 & ~n352;
  assign n956 = ~n344 & ~n348;
  assign n957 = n955 & n956;
  assign n958 = n952 & n957;
  assign n959 = n708 & n859;
  assign n960 = n810 & n861;
  assign n961 = n959 & n960;
  assign po32 = ~n958 | ~n961;
  assign n963 = ~n209 & ~n217;
  assign n964 = ~n220 & n963;
  assign n965 = ~n182 & ~n194;
  assign n966 = ~n205 & n965;
  assign n967 = n964 & n966;
  assign n968 = ~n129 & ~n159;
  assign n969 = ~n352 & n968;
  assign n970 = ~n170 & ~n173;
  assign n971 = ~n176 & n970;
  assign n972 = n969 & n971;
  assign n973 = n967 & n972;
  assign n974 = n810 & n944;
  assign n975 = ~n117 & ~n348;
  assign n976 = ~po11 & n975;
  assign n977 = n945 & n976;
  assign n978 = n974 & n977;
  assign po33 = ~n973 | ~n978;
  assign po37 = n454 | n690;
  assign po05 = po02;
  assign po06 = po02;
endmodule



// Benchmark "i6" written by ABC on Sun Apr 22 21:43:05 2018

module i6 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66;
  wire n206, n207, n208, n209, n210, n211, n212, n214, n215, n216, n217,
    n218, n219, n220, n222, n223, n224, n225, n226, n227, n228, n230, n231,
    n232, n233, n234, n235, n236, n238, n239, n240, n241, n242, n243, n244,
    n246, n247, n248, n249, n250, n251, n252, n254, n255, n256, n257, n258,
    n259, n260, n262, n263, n264, n265, n266, n267, n268, n270, n271, n272,
    n273, n274, n275, n276, n278, n279, n280, n281, n282, n283, n284, n286,
    n287, n288, n289, n290, n291, n292, n294, n295, n296, n297, n298, n299,
    n300, n302, n303, n304, n305, n306, n307, n308, n310, n311, n312, n313,
    n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n326, n327,
    n328, n329, n330, n331, n332, n334, n335, n336, n337, n338, n339, n340,
    n342, n343, n344, n345, n346, n347, n348, n350, n351, n352, n353, n354,
    n355, n356, n358, n359, n360, n361, n362, n363, n364, n366, n367, n368,
    n369, n370, n371, n372, n374, n375, n376, n377, n378, n379, n380, n382,
    n383, n384, n385, n386, n387, n388, n390, n391, n392, n393, n394, n395,
    n396, n398, n399, n400, n401, n402, n403, n404, n406, n407, n408, n409,
    n410, n411, n412, n414, n415, n416, n417, n418, n419, n420, n422, n423,
    n424, n425, n426, n427, n428, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896;
  assign n206 = ~pi001 & pi002;
  assign n207 = ~pi000 & n206;
  assign n208 = ~pi001 & pi030;
  assign n209 = pi000 & n208;
  assign n210 = pi001 & ~pi030;
  assign n211 = pi000 & n210;
  assign n212 = ~n207 & ~n209;
  assign po00 = n211 | ~n212;
  assign n214 = ~pi001 & pi003;
  assign n215 = ~pi000 & n214;
  assign n216 = ~pi001 & pi031;
  assign n217 = pi000 & n216;
  assign n218 = pi001 & ~pi031;
  assign n219 = pi000 & n218;
  assign n220 = ~n215 & ~n217;
  assign po01 = n219 | ~n220;
  assign n222 = ~pi001 & pi004;
  assign n223 = ~pi000 & n222;
  assign n224 = ~pi001 & pi032;
  assign n225 = pi000 & n224;
  assign n226 = pi001 & ~pi032;
  assign n227 = pi000 & n226;
  assign n228 = ~n223 & ~n225;
  assign po02 = n227 | ~n228;
  assign n230 = ~pi001 & pi005;
  assign n231 = ~pi000 & n230;
  assign n232 = ~pi001 & pi033;
  assign n233 = pi000 & n232;
  assign n234 = pi001 & ~pi033;
  assign n235 = pi000 & n234;
  assign n236 = ~n231 & ~n233;
  assign po03 = n235 | ~n236;
  assign n238 = ~pi001 & pi006;
  assign n239 = ~pi000 & n238;
  assign n240 = ~pi001 & pi034;
  assign n241 = pi000 & n240;
  assign n242 = pi001 & ~pi034;
  assign n243 = pi000 & n242;
  assign n244 = ~n239 & ~n241;
  assign po04 = n243 | ~n244;
  assign n246 = ~pi001 & pi007;
  assign n247 = ~pi000 & n246;
  assign n248 = ~pi001 & pi035;
  assign n249 = pi000 & n248;
  assign n250 = pi001 & ~pi035;
  assign n251 = pi000 & n250;
  assign n252 = ~n247 & ~n249;
  assign po05 = n251 | ~n252;
  assign n254 = ~pi001 & pi008;
  assign n255 = ~pi000 & n254;
  assign n256 = ~pi001 & pi036;
  assign n257 = pi000 & n256;
  assign n258 = pi001 & ~pi036;
  assign n259 = pi000 & n258;
  assign n260 = ~n255 & ~n257;
  assign po06 = n259 | ~n260;
  assign n262 = ~pi001 & pi009;
  assign n263 = ~pi000 & n262;
  assign n264 = ~pi001 & pi037;
  assign n265 = pi000 & n264;
  assign n266 = pi001 & ~pi037;
  assign n267 = pi000 & n266;
  assign n268 = ~n263 & ~n265;
  assign po07 = n267 | ~n268;
  assign n270 = ~pi001 & pi010;
  assign n271 = ~pi000 & n270;
  assign n272 = ~pi001 & pi038;
  assign n273 = pi000 & n272;
  assign n274 = pi001 & ~pi038;
  assign n275 = pi000 & n274;
  assign n276 = ~n271 & ~n273;
  assign po08 = n275 | ~n276;
  assign n278 = ~pi001 & pi011;
  assign n279 = ~pi000 & n278;
  assign n280 = ~pi001 & pi039;
  assign n281 = pi000 & n280;
  assign n282 = pi001 & ~pi039;
  assign n283 = pi000 & n282;
  assign n284 = ~n279 & ~n281;
  assign po09 = n283 | ~n284;
  assign n286 = ~pi001 & pi012;
  assign n287 = ~pi000 & n286;
  assign n288 = ~pi001 & pi040;
  assign n289 = pi000 & n288;
  assign n290 = pi001 & ~pi040;
  assign n291 = pi000 & n290;
  assign n292 = ~n287 & ~n289;
  assign po10 = n291 | ~n292;
  assign n294 = ~pi001 & pi013;
  assign n295 = ~pi000 & n294;
  assign n296 = ~pi001 & pi041;
  assign n297 = pi000 & n296;
  assign n298 = pi001 & ~pi041;
  assign n299 = pi000 & n298;
  assign n300 = ~n295 & ~n297;
  assign po11 = n299 | ~n300;
  assign n302 = ~pi001 & pi014;
  assign n303 = ~pi000 & n302;
  assign n304 = ~pi001 & pi042;
  assign n305 = pi000 & n304;
  assign n306 = pi001 & ~pi042;
  assign n307 = pi000 & n306;
  assign n308 = ~n303 & ~n305;
  assign po12 = n307 | ~n308;
  assign n310 = ~pi001 & pi015;
  assign n311 = ~pi000 & n310;
  assign n312 = ~pi001 & pi043;
  assign n313 = pi000 & n312;
  assign n314 = pi001 & ~pi043;
  assign n315 = pi000 & n314;
  assign n316 = ~n311 & ~n313;
  assign po13 = n315 | ~n316;
  assign n318 = ~pi001 & pi016;
  assign n319 = ~pi000 & n318;
  assign n320 = ~pi001 & pi044;
  assign n321 = pi000 & n320;
  assign n322 = pi001 & ~pi044;
  assign n323 = pi000 & n322;
  assign n324 = ~n319 & ~n321;
  assign po14 = n323 | ~n324;
  assign n326 = ~pi001 & pi017;
  assign n327 = ~pi000 & n326;
  assign n328 = ~pi001 & pi045;
  assign n329 = pi000 & n328;
  assign n330 = pi001 & ~pi045;
  assign n331 = pi000 & n330;
  assign n332 = ~n327 & ~n329;
  assign po15 = n331 | ~n332;
  assign n334 = ~pi001 & pi018;
  assign n335 = ~pi000 & n334;
  assign n336 = ~pi001 & pi046;
  assign n337 = pi000 & n336;
  assign n338 = pi001 & ~pi046;
  assign n339 = pi000 & n338;
  assign n340 = ~n335 & ~n337;
  assign po16 = n339 | ~n340;
  assign n342 = ~pi001 & pi019;
  assign n343 = ~pi000 & n342;
  assign n344 = ~pi001 & pi047;
  assign n345 = pi000 & n344;
  assign n346 = pi001 & ~pi047;
  assign n347 = pi000 & n346;
  assign n348 = ~n343 & ~n345;
  assign po17 = n347 | ~n348;
  assign n350 = ~pi001 & pi020;
  assign n351 = ~pi000 & n350;
  assign n352 = ~pi001 & pi048;
  assign n353 = pi000 & n352;
  assign n354 = pi001 & ~pi048;
  assign n355 = pi000 & n354;
  assign n356 = ~n351 & ~n353;
  assign po18 = n355 | ~n356;
  assign n358 = ~pi001 & pi021;
  assign n359 = ~pi000 & n358;
  assign n360 = ~pi001 & pi049;
  assign n361 = pi000 & n360;
  assign n362 = pi001 & ~pi049;
  assign n363 = pi000 & n362;
  assign n364 = ~n359 & ~n361;
  assign po19 = n363 | ~n364;
  assign n366 = ~pi001 & pi022;
  assign n367 = ~pi000 & n366;
  assign n368 = ~pi001 & pi050;
  assign n369 = pi000 & n368;
  assign n370 = pi001 & ~pi050;
  assign n371 = pi000 & n370;
  assign n372 = ~n367 & ~n369;
  assign po20 = n371 | ~n372;
  assign n374 = ~pi001 & pi023;
  assign n375 = ~pi000 & n374;
  assign n376 = ~pi001 & pi051;
  assign n377 = pi000 & n376;
  assign n378 = pi001 & ~pi051;
  assign n379 = pi000 & n378;
  assign n380 = ~n375 & ~n377;
  assign po21 = n379 | ~n380;
  assign n382 = ~pi001 & pi024;
  assign n383 = ~pi000 & n382;
  assign n384 = ~pi001 & pi052;
  assign n385 = pi000 & n384;
  assign n386 = pi001 & ~pi052;
  assign n387 = pi000 & n386;
  assign n388 = ~n383 & ~n385;
  assign po22 = n387 | ~n388;
  assign n390 = ~pi001 & pi025;
  assign n391 = ~pi000 & n390;
  assign n392 = ~pi001 & pi053;
  assign n393 = pi000 & n392;
  assign n394 = pi001 & ~pi053;
  assign n395 = pi000 & n394;
  assign n396 = ~n391 & ~n393;
  assign po23 = n395 | ~n396;
  assign n398 = ~pi001 & pi026;
  assign n399 = ~pi000 & n398;
  assign n400 = ~pi001 & pi054;
  assign n401 = pi000 & n400;
  assign n402 = pi001 & ~pi054;
  assign n403 = pi000 & n402;
  assign n404 = ~n399 & ~n401;
  assign po24 = n403 | ~n404;
  assign n406 = ~pi001 & pi027;
  assign n407 = ~pi000 & n406;
  assign n408 = ~pi001 & pi055;
  assign n409 = pi000 & n408;
  assign n410 = pi001 & ~pi055;
  assign n411 = pi000 & n410;
  assign n412 = ~n407 & ~n409;
  assign po25 = n411 | ~n412;
  assign n414 = ~pi001 & pi028;
  assign n415 = ~pi000 & n414;
  assign n416 = ~pi001 & pi056;
  assign n417 = pi000 & n416;
  assign n418 = pi001 & ~pi056;
  assign n419 = pi000 & n418;
  assign n420 = ~n415 & ~n417;
  assign po26 = n419 | ~n420;
  assign n422 = ~pi001 & pi029;
  assign n423 = ~pi000 & n422;
  assign n424 = ~pi001 & pi057;
  assign n425 = pi000 & n424;
  assign n426 = pi001 & ~pi057;
  assign n427 = pi000 & n426;
  assign n428 = ~n423 & ~n425;
  assign po27 = n427 | ~n428;
  assign n430 = ~pi000 & pi058;
  assign n431 = ~pi001 & n430;
  assign n432 = pi059 & n431;
  assign n433 = pi000 & pi091;
  assign n434 = ~pi001 & n433;
  assign n435 = pi059 & n434;
  assign n436 = pi000 & ~pi091;
  assign n437 = pi001 & n436;
  assign n438 = pi059 & n437;
  assign n439 = pi001 & ~pi059;
  assign n440 = ~n432 & ~n435;
  assign n441 = ~n438 & ~n439;
  assign po28 = ~n440 | ~n441;
  assign n443 = ~pi000 & pi060;
  assign n444 = ~pi001 & n443;
  assign n445 = pi059 & n444;
  assign n446 = pi000 & pi092;
  assign n447 = ~pi001 & n446;
  assign n448 = pi059 & n447;
  assign n449 = pi000 & ~pi092;
  assign n450 = pi001 & n449;
  assign n451 = pi059 & n450;
  assign n452 = ~n445 & ~n448;
  assign n453 = ~n439 & ~n451;
  assign po29 = ~n452 | ~n453;
  assign n455 = ~pi000 & pi061;
  assign n456 = ~pi001 & n455;
  assign n457 = pi059 & n456;
  assign n458 = pi000 & pi093;
  assign n459 = ~pi001 & n458;
  assign n460 = pi059 & n459;
  assign n461 = pi000 & ~pi093;
  assign n462 = pi001 & n461;
  assign n463 = pi059 & n462;
  assign n464 = ~n457 & ~n460;
  assign n465 = ~n439 & ~n463;
  assign po30 = ~n464 | ~n465;
  assign n467 = ~pi000 & pi062;
  assign n468 = ~pi001 & n467;
  assign n469 = pi059 & n468;
  assign n470 = pi000 & pi094;
  assign n471 = ~pi001 & n470;
  assign n472 = pi059 & n471;
  assign n473 = pi000 & ~pi094;
  assign n474 = pi001 & n473;
  assign n475 = pi059 & n474;
  assign n476 = ~n469 & ~n472;
  assign n477 = ~n439 & ~n475;
  assign po31 = ~n476 | ~n477;
  assign n479 = ~pi000 & pi063;
  assign n480 = ~pi001 & n479;
  assign n481 = pi059 & n480;
  assign n482 = pi000 & pi095;
  assign n483 = ~pi001 & n482;
  assign n484 = pi059 & n483;
  assign n485 = pi000 & ~pi095;
  assign n486 = pi001 & n485;
  assign n487 = pi059 & n486;
  assign n488 = ~n481 & ~n484;
  assign n489 = ~n439 & ~n487;
  assign po32 = ~n488 | ~n489;
  assign n491 = ~pi000 & pi064;
  assign n492 = ~pi001 & n491;
  assign n493 = pi059 & n492;
  assign n494 = pi000 & pi096;
  assign n495 = ~pi001 & n494;
  assign n496 = pi059 & n495;
  assign n497 = pi000 & ~pi096;
  assign n498 = pi001 & n497;
  assign n499 = pi059 & n498;
  assign n500 = ~n493 & ~n496;
  assign n501 = ~n439 & ~n499;
  assign po33 = ~n500 | ~n501;
  assign n503 = ~pi000 & pi065;
  assign n504 = ~pi001 & n503;
  assign n505 = pi059 & n504;
  assign n506 = pi000 & pi097;
  assign n507 = ~pi001 & n506;
  assign n508 = pi059 & n507;
  assign n509 = pi000 & ~pi097;
  assign n510 = pi001 & n509;
  assign n511 = pi059 & n510;
  assign n512 = ~n505 & ~n508;
  assign n513 = ~n439 & ~n511;
  assign po34 = ~n512 | ~n513;
  assign n515 = ~pi000 & pi066;
  assign n516 = ~pi001 & n515;
  assign n517 = pi059 & n516;
  assign n518 = pi000 & pi098;
  assign n519 = ~pi001 & n518;
  assign n520 = pi059 & n519;
  assign n521 = pi000 & ~pi098;
  assign n522 = pi001 & n521;
  assign n523 = pi059 & n522;
  assign n524 = ~n517 & ~n520;
  assign n525 = ~n439 & ~n523;
  assign po35 = ~n524 | ~n525;
  assign n527 = ~pi000 & pi067;
  assign n528 = ~pi001 & n527;
  assign n529 = pi059 & n528;
  assign n530 = pi000 & pi099;
  assign n531 = ~pi001 & n530;
  assign n532 = pi059 & n531;
  assign n533 = pi000 & ~pi099;
  assign n534 = pi001 & n533;
  assign n535 = pi059 & n534;
  assign n536 = ~n529 & ~n532;
  assign n537 = ~n439 & ~n535;
  assign po36 = ~n536 | ~n537;
  assign n539 = ~pi000 & pi068;
  assign n540 = ~pi001 & n539;
  assign n541 = pi059 & n540;
  assign n542 = pi000 & pi100;
  assign n543 = ~pi001 & n542;
  assign n544 = pi059 & n543;
  assign n545 = pi000 & ~pi100;
  assign n546 = pi001 & n545;
  assign n547 = pi059 & n546;
  assign n548 = ~n541 & ~n544;
  assign n549 = ~n439 & ~n547;
  assign po37 = ~n548 | ~n549;
  assign n551 = ~pi000 & pi069;
  assign n552 = ~pi001 & n551;
  assign n553 = pi059 & n552;
  assign n554 = pi000 & pi101;
  assign n555 = ~pi001 & n554;
  assign n556 = pi059 & n555;
  assign n557 = pi000 & ~pi101;
  assign n558 = pi001 & n557;
  assign n559 = pi059 & n558;
  assign n560 = ~n553 & ~n556;
  assign n561 = ~n439 & ~n559;
  assign po38 = ~n560 | ~n561;
  assign n563 = ~pi000 & pi070;
  assign n564 = ~pi001 & n563;
  assign n565 = pi059 & n564;
  assign n566 = pi000 & pi102;
  assign n567 = ~pi001 & n566;
  assign n568 = pi059 & n567;
  assign n569 = pi000 & ~pi102;
  assign n570 = pi001 & n569;
  assign n571 = pi059 & n570;
  assign n572 = ~n565 & ~n568;
  assign n573 = ~n439 & ~n571;
  assign po39 = ~n572 | ~n573;
  assign n575 = ~pi000 & pi071;
  assign n576 = ~pi001 & n575;
  assign n577 = pi059 & n576;
  assign n578 = pi000 & pi103;
  assign n579 = ~pi001 & n578;
  assign n580 = pi059 & n579;
  assign n581 = pi000 & ~pi103;
  assign n582 = pi001 & n581;
  assign n583 = pi059 & n582;
  assign n584 = ~n577 & ~n580;
  assign n585 = ~n439 & ~n583;
  assign po40 = ~n584 | ~n585;
  assign n587 = ~pi000 & pi072;
  assign n588 = ~pi001 & n587;
  assign n589 = pi059 & n588;
  assign n590 = pi000 & pi104;
  assign n591 = ~pi001 & n590;
  assign n592 = pi059 & n591;
  assign n593 = pi000 & ~pi104;
  assign n594 = pi001 & n593;
  assign n595 = pi059 & n594;
  assign n596 = ~n589 & ~n592;
  assign n597 = ~n439 & ~n595;
  assign po41 = ~n596 | ~n597;
  assign n599 = ~pi000 & pi073;
  assign n600 = ~pi001 & n599;
  assign n601 = pi059 & n600;
  assign n602 = pi000 & pi105;
  assign n603 = ~pi001 & n602;
  assign n604 = pi059 & n603;
  assign n605 = pi000 & ~pi105;
  assign n606 = pi001 & n605;
  assign n607 = pi059 & n606;
  assign n608 = ~n601 & ~n604;
  assign n609 = ~n439 & ~n607;
  assign po42 = ~n608 | ~n609;
  assign n611 = ~pi000 & pi074;
  assign n612 = ~pi001 & n611;
  assign n613 = pi059 & n612;
  assign n614 = pi000 & pi106;
  assign n615 = ~pi001 & n614;
  assign n616 = pi059 & n615;
  assign n617 = pi000 & ~pi106;
  assign n618 = pi001 & n617;
  assign n619 = pi059 & n618;
  assign n620 = ~n613 & ~n616;
  assign n621 = ~n439 & ~n619;
  assign po43 = ~n620 | ~n621;
  assign n623 = ~pi000 & pi075;
  assign n624 = ~pi001 & n623;
  assign n625 = pi059 & n624;
  assign n626 = pi000 & pi107;
  assign n627 = ~pi001 & n626;
  assign n628 = pi059 & n627;
  assign n629 = pi000 & ~pi107;
  assign n630 = pi001 & n629;
  assign n631 = pi059 & n630;
  assign n632 = ~n625 & ~n628;
  assign n633 = ~n439 & ~n631;
  assign po44 = ~n632 | ~n633;
  assign n635 = ~pi000 & pi076;
  assign n636 = ~pi001 & n635;
  assign n637 = pi059 & n636;
  assign n638 = pi000 & pi108;
  assign n639 = ~pi001 & n638;
  assign n640 = pi059 & n639;
  assign n641 = pi000 & ~pi108;
  assign n642 = pi001 & n641;
  assign n643 = pi059 & n642;
  assign n644 = ~n637 & ~n640;
  assign n645 = ~n439 & ~n643;
  assign po45 = ~n644 | ~n645;
  assign n647 = ~pi000 & pi077;
  assign n648 = ~pi001 & n647;
  assign n649 = pi059 & n648;
  assign n650 = pi000 & pi109;
  assign n651 = ~pi001 & n650;
  assign n652 = pi059 & n651;
  assign n653 = pi000 & ~pi109;
  assign n654 = pi001 & n653;
  assign n655 = pi059 & n654;
  assign n656 = ~n649 & ~n652;
  assign n657 = ~n439 & ~n655;
  assign po46 = ~n656 | ~n657;
  assign n659 = ~pi000 & pi078;
  assign n660 = ~pi001 & n659;
  assign n661 = pi059 & n660;
  assign n662 = pi000 & pi110;
  assign n663 = ~pi001 & n662;
  assign n664 = pi059 & n663;
  assign n665 = pi000 & ~pi110;
  assign n666 = pi001 & n665;
  assign n667 = pi059 & n666;
  assign n668 = ~n661 & ~n664;
  assign n669 = ~n439 & ~n667;
  assign po47 = ~n668 | ~n669;
  assign n671 = ~pi000 & pi079;
  assign n672 = ~pi001 & n671;
  assign n673 = pi059 & n672;
  assign n674 = pi000 & pi111;
  assign n675 = ~pi001 & n674;
  assign n676 = pi059 & n675;
  assign n677 = pi000 & ~pi111;
  assign n678 = pi001 & n677;
  assign n679 = pi059 & n678;
  assign n680 = ~n673 & ~n676;
  assign n681 = ~n439 & ~n679;
  assign po48 = ~n680 | ~n681;
  assign n683 = ~pi000 & pi080;
  assign n684 = ~pi001 & n683;
  assign n685 = pi059 & n684;
  assign n686 = pi000 & pi112;
  assign n687 = ~pi001 & n686;
  assign n688 = pi059 & n687;
  assign n689 = pi000 & ~pi112;
  assign n690 = pi001 & n689;
  assign n691 = pi059 & n690;
  assign n692 = ~n685 & ~n688;
  assign n693 = ~n439 & ~n691;
  assign po49 = ~n692 | ~n693;
  assign n695 = ~pi000 & pi081;
  assign n696 = ~pi001 & n695;
  assign n697 = pi059 & n696;
  assign n698 = pi000 & pi113;
  assign n699 = ~pi001 & n698;
  assign n700 = pi059 & n699;
  assign n701 = pi000 & ~pi113;
  assign n702 = pi001 & n701;
  assign n703 = pi059 & n702;
  assign n704 = ~n697 & ~n700;
  assign n705 = ~n439 & ~n703;
  assign po50 = ~n704 | ~n705;
  assign n707 = ~pi000 & pi082;
  assign n708 = ~pi001 & n707;
  assign n709 = pi059 & n708;
  assign n710 = pi000 & pi114;
  assign n711 = ~pi001 & n710;
  assign n712 = pi059 & n711;
  assign n713 = pi000 & ~pi114;
  assign n714 = pi001 & n713;
  assign n715 = pi059 & n714;
  assign n716 = ~n709 & ~n712;
  assign n717 = ~n439 & ~n715;
  assign po51 = ~n716 | ~n717;
  assign n719 = ~pi000 & pi083;
  assign n720 = ~pi001 & n719;
  assign n721 = pi059 & n720;
  assign n722 = pi000 & pi115;
  assign n723 = ~pi001 & n722;
  assign n724 = pi059 & n723;
  assign n725 = pi000 & ~pi115;
  assign n726 = pi001 & n725;
  assign n727 = pi059 & n726;
  assign n728 = ~n721 & ~n724;
  assign n729 = ~n439 & ~n727;
  assign po52 = ~n728 | ~n729;
  assign n731 = ~pi000 & pi084;
  assign n732 = ~pi001 & n731;
  assign n733 = pi059 & n732;
  assign n734 = pi000 & pi116;
  assign n735 = ~pi001 & n734;
  assign n736 = pi059 & n735;
  assign n737 = pi000 & ~pi116;
  assign n738 = pi001 & n737;
  assign n739 = pi059 & n738;
  assign n740 = ~n733 & ~n736;
  assign n741 = ~n439 & ~n739;
  assign po53 = ~n740 | ~n741;
  assign n743 = ~pi000 & pi085;
  assign n744 = ~pi001 & n743;
  assign n745 = pi059 & n744;
  assign n746 = pi000 & pi117;
  assign n747 = ~pi001 & n746;
  assign n748 = pi059 & n747;
  assign n749 = pi000 & ~pi117;
  assign n750 = pi001 & n749;
  assign n751 = pi059 & n750;
  assign n752 = ~n745 & ~n748;
  assign n753 = ~n439 & ~n751;
  assign po54 = ~n752 | ~n753;
  assign n755 = ~pi000 & pi086;
  assign n756 = ~pi001 & n755;
  assign n757 = pi059 & n756;
  assign n758 = pi000 & pi118;
  assign n759 = ~pi001 & n758;
  assign n760 = pi059 & n759;
  assign n761 = pi000 & ~pi118;
  assign n762 = pi001 & n761;
  assign n763 = pi059 & n762;
  assign n764 = ~n757 & ~n760;
  assign n765 = ~n439 & ~n763;
  assign po55 = ~n764 | ~n765;
  assign n767 = ~pi000 & pi087;
  assign n768 = ~pi001 & n767;
  assign n769 = pi059 & n768;
  assign n770 = pi000 & pi119;
  assign n771 = ~pi001 & n770;
  assign n772 = pi059 & n771;
  assign n773 = pi000 & ~pi119;
  assign n774 = pi001 & n773;
  assign n775 = pi059 & n774;
  assign n776 = ~n769 & ~n772;
  assign n777 = ~n439 & ~n775;
  assign po56 = ~n776 | ~n777;
  assign n779 = ~pi000 & pi088;
  assign n780 = ~pi001 & n779;
  assign n781 = pi059 & n780;
  assign n782 = pi000 & pi120;
  assign n783 = ~pi001 & n782;
  assign n784 = pi059 & n783;
  assign n785 = pi000 & ~pi120;
  assign n786 = pi001 & n785;
  assign n787 = pi059 & n786;
  assign n788 = ~n781 & ~n784;
  assign n789 = ~n439 & ~n787;
  assign po57 = ~n788 | ~n789;
  assign n791 = ~pi000 & pi089;
  assign n792 = ~pi001 & n791;
  assign n793 = pi059 & n792;
  assign n794 = pi000 & pi121;
  assign n795 = ~pi001 & n794;
  assign n796 = pi059 & n795;
  assign n797 = pi000 & ~pi121;
  assign n798 = pi001 & n797;
  assign n799 = pi059 & n798;
  assign n800 = ~n793 & ~n796;
  assign n801 = ~n439 & ~n799;
  assign po58 = ~n800 | ~n801;
  assign n803 = ~pi000 & pi090;
  assign n804 = ~pi001 & n803;
  assign n805 = pi059 & n804;
  assign n806 = pi000 & pi122;
  assign n807 = ~pi001 & n806;
  assign n808 = pi059 & n807;
  assign n809 = pi000 & ~pi122;
  assign n810 = pi001 & n809;
  assign n811 = pi059 & n810;
  assign n812 = ~n805 & ~n808;
  assign n813 = ~n439 & ~n811;
  assign po59 = ~n812 | ~n813;
  assign n815 = ~pi000 & pi123;
  assign n816 = ~pi001 & n815;
  assign n817 = pi124 & n816;
  assign n818 = pi000 & pi131;
  assign n819 = ~pi001 & n818;
  assign n820 = pi124 & n819;
  assign n821 = pi001 & n818;
  assign n822 = pi124 & n821;
  assign n823 = ~n817 & ~n820;
  assign po60 = n822 | ~n823;
  assign n825 = ~pi000 & pi125;
  assign n826 = ~pi001 & n825;
  assign n827 = pi124 & n826;
  assign n828 = pi000 & pi132;
  assign n829 = ~pi001 & n828;
  assign n830 = pi124 & n829;
  assign n831 = pi000 & ~pi132;
  assign n832 = pi001 & n831;
  assign n833 = pi124 & n832;
  assign n834 = pi001 & ~pi124;
  assign n835 = ~n827 & ~n830;
  assign n836 = ~n833 & ~n834;
  assign po61 = ~n835 | ~n836;
  assign n838 = ~pi000 & pi126;
  assign n839 = ~pi001 & n838;
  assign n840 = pi124 & n839;
  assign n841 = pi000 & pi133;
  assign n842 = ~pi001 & n841;
  assign n843 = pi124 & n842;
  assign n844 = pi000 & ~pi133;
  assign n845 = pi001 & n844;
  assign n846 = pi124 & n845;
  assign n847 = ~n840 & ~n843;
  assign n848 = ~n834 & ~n846;
  assign po62 = ~n847 | ~n848;
  assign n850 = ~pi000 & pi127;
  assign n851 = ~pi001 & n850;
  assign n852 = pi124 & n851;
  assign n853 = pi000 & pi134;
  assign n854 = ~pi001 & n853;
  assign n855 = pi124 & n854;
  assign n856 = pi000 & ~pi134;
  assign n857 = pi001 & n856;
  assign n858 = pi124 & n857;
  assign n859 = ~n852 & ~n855;
  assign n860 = ~n834 & ~n858;
  assign po63 = ~n859 | ~n860;
  assign n862 = ~pi000 & pi128;
  assign n863 = ~pi001 & n862;
  assign n864 = pi124 & n863;
  assign n865 = pi000 & pi135;
  assign n866 = ~pi001 & n865;
  assign n867 = pi124 & n866;
  assign n868 = pi000 & ~pi135;
  assign n869 = pi001 & n868;
  assign n870 = pi124 & n869;
  assign n871 = ~n864 & ~n867;
  assign n872 = ~n834 & ~n870;
  assign po64 = ~n871 | ~n872;
  assign n874 = ~pi000 & pi129;
  assign n875 = ~pi001 & n874;
  assign n876 = pi124 & n875;
  assign n877 = pi000 & pi136;
  assign n878 = ~pi001 & n877;
  assign n879 = pi124 & n878;
  assign n880 = pi000 & ~pi136;
  assign n881 = pi001 & n880;
  assign n882 = pi124 & n881;
  assign n883 = ~n876 & ~n879;
  assign n884 = ~n834 & ~n882;
  assign po65 = ~n883 | ~n884;
  assign n886 = ~pi000 & pi130;
  assign n887 = ~pi001 & n886;
  assign n888 = pi124 & n887;
  assign n889 = pi000 & pi137;
  assign n890 = ~pi001 & n889;
  assign n891 = pi124 & n890;
  assign n892 = pi000 & ~pi137;
  assign n893 = pi001 & n892;
  assign n894 = pi124 & n893;
  assign n895 = ~n888 & ~n891;
  assign n896 = ~n834 & ~n894;
  assign po66 = ~n895 | ~n896;
endmodule



module cavlc_best_speed (
        pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9, 
        po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10);
input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744;
assign w0 = ~pi4 & ~pi7;
assign w1 = ~pi1 & pi2;
assign w2 = pi0 & ~pi9;
assign w3 = w1 & w2;
assign w4 = ~pi0 & pi9;
assign w5 = pi1 & ~pi8;
assign w6 = (~pi8 & w4) | (~pi8 & w5) | (w4 & w5);
assign w7 = ~w3 & ~w6;
assign w8 = pi3 & ~pi5;
assign w9 = ~pi8 & ~w8;
assign w10 = (~pi8 & w7) | (~pi8 & w9) | (w7 & w9);
assign w11 = ~pi5 & ~w7;
assign w12 = ~pi0 & ~pi9;
assign w13 = pi0 & pi9;
assign w14 = ~w12 & ~w13;
assign w15 = pi2 & pi5;
assign w16 = pi1 & w15;
assign w17 = ~w14 & w16;
assign w18 = ~pi1 & ~pi2;
assign w19 = w4 & w18;
assign w20 = pi5 & pi6;
assign w21 = (pi6 & w19) | (pi6 & w20) | (w19 & w20);
assign w22 = ~w17 & ~w21;
assign w23 = ~w11 & w22;
assign w24 = pi3 & ~w23;
assign w25 = ~pi2 & ~pi3;
assign w26 = pi1 & w25;
assign w27 = ~w14 & w26;
assign w28 = pi2 & pi6;
assign w29 = (pi6 & w2) | (pi6 & w28) | (w2 & w28);
assign w30 = pi5 & w29;
assign w31 = (pi5 & w27) | (pi5 & w30) | (w27 & w30);
assign w32 = ~pi2 & ~pi9;
assign w33 = pi1 & w32;
assign w34 = pi2 & pi9;
assign w35 = pi6 & w34;
assign w36 = (pi6 & w33) | (pi6 & w35) | (w33 & w35);
assign w37 = ~pi0 & ~pi3;
assign w38 = w36 & w37;
assign w39 = ~w31 & ~w38;
assign w40 = ~w10 & ~w39;
assign w41 = (~w10 & w24) | (~w10 & w40) | (w24 & w40);
assign w42 = ~pi5 & ~pi8;
assign w43 = ~pi2 & pi6;
assign w44 = ~pi3 & ~pi9;
assign w45 = (~pi9 & w43) | (~pi9 & w44) | (w43 & w44);
assign w46 = pi1 & ~w34;
assign w47 = (~w34 & ~w45) | (~w34 & w46) | (~w45 & w46);
assign w48 = w42 & ~w47;
assign w49 = ~pi5 & w5;
assign w50 = ~pi8 & ~pi9;
assign w51 = ~pi2 & w50;
assign w52 = ~pi5 & pi9;
assign w53 = pi2 & w52;
assign w54 = ~w51 & ~w53;
assign w55 = ~pi1 & ~pi3;
assign w56 = ~w49 & ~w55;
assign w57 = (~w49 & w54) | (~w49 & w56) | (w54 & w56);
assign w58 = ~pi0 & ~w57;
assign w59 = ~w48 & ~w58;
assign w60 = w0 & ~w59;
assign w61 = (w0 & w41) | (w0 & w60) | (w41 & w60);
assign w62 = pi6 & ~pi9;
assign w63 = ~pi5 & w62;
assign w64 = pi4 & pi9;
assign w65 = ~w20 & w64;
assign w66 = ~w63 & ~w65;
assign w67 = ~pi8 & ~w66;
assign w68 = pi6 & pi8;
assign w69 = pi4 & w68;
assign w70 = ~pi6 & w50;
assign w71 = ~w69 & ~w70;
assign w72 = pi5 & ~w71;
assign w73 = ~w67 & ~w72;
assign w74 = ~pi0 & ~pi1;
assign w75 = w25 & w74;
assign w76 = ~pi7 & w75;
assign w77 = ~w73 & w76;
assign w78 = pi1 & pi9;
assign w79 = ~pi0 & w78;
assign w80 = ~pi1 & ~pi9;
assign w81 = ~pi5 & w80;
assign w82 = (~pi5 & w79) | (~pi5 & w81) | (w79 & w81);
assign w83 = ~pi3 & w82;
assign w84 = pi0 & w80;
assign w85 = ~pi7 & w78;
assign w86 = (~pi7 & w84) | (~pi7 & w85) | (w84 & w85);
assign w87 = ~pi2 & w86;
assign w88 = (~pi2 & w83) | (~pi2 & w87) | (w83 & w87);
assign w89 = ~pi8 & w88;
assign w90 = pi3 & w2;
assign w91 = ~pi3 & pi9;
assign w92 = ~pi0 & ~pi5;
assign w93 = ~w91 & ~w92;
assign w94 = ~w90 & w93;
assign w95 = ~pi2 & ~w94;
assign w96 = pi0 & ~pi1;
assign w97 = w44 & w96;
assign w98 = pi3 & pi9;
assign w99 = pi1 & w98;
assign w100 = ~w97 & ~w99;
assign w101 = ~pi7 & ~pi8;
assign w102 = w100 & w101;
assign w103 = ~w95 & w102;
assign w104 = pi0 & ~pi2;
assign w105 = ~pi5 & pi8;
assign w106 = ~pi7 & pi9;
assign w107 = (pi9 & w105) | (pi9 & w106) | (w105 & w106);
assign w108 = pi1 & w107;
assign w109 = pi1 & ~pi7;
assign w110 = ~pi5 & ~pi9;
assign w111 = ~w109 & w110;
assign w112 = w104 & w111;
assign w113 = (w104 & w108) | (w104 & w112) | (w108 & w112);
assign w114 = ~pi5 & pi7;
assign w115 = pi8 & ~pi9;
assign w116 = w114 & w115;
assign w117 = ~pi0 & pi2;
assign w118 = ~pi1 & w117;
assign w119 = w116 & w118;
assign w120 = ~pi3 & w119;
assign w121 = (~pi3 & w113) | (~pi3 & w120) | (w113 & w120);
assign w122 = ~w103 & ~w121;
assign w123 = ~w89 & w122;
assign w124 = ~pi4 & ~pi6;
assign w125 = ~w77 & ~w124;
assign w126 = (~w77 & w123) | (~w77 & w125) | (w123 & w125);
assign w127 = ~w61 & w126;
assign w128 = pi0 & ~pi8;
assign w129 = pi1 & pi8;
assign w130 = ~w128 & ~w129;
assign w131 = ~pi9 & ~w130;
assign w132 = pi1 & w128;
assign w133 = ~pi2 & w132;
assign w134 = (~pi2 & w131) | (~pi2 & w133) | (w131 & w133);
assign w135 = w80 & w117;
assign w136 = ~pi7 & ~w135;
assign w137 = ~pi1 & ~pi8;
assign w138 = w117 & w137;
assign w139 = pi7 & w138;
assign w140 = ~w135 & ~w139;
assign w141 = (~w134 & w136) | (~w134 & w140) | (w136 & w140);
assign w142 = ~pi3 & ~pi5;
assign w143 = w124 & w142;
assign w144 = ~w141 & w143;
assign w145 = ~pi8 & pi9;
assign w146 = ~pi0 & pi5;
assign w147 = w145 & w146;
assign w148 = pi6 & w145;
assign w149 = ~pi6 & pi8;
assign w150 = ~pi5 & w149;
assign w151 = ~w148 & ~w150;
assign w152 = ~pi0 & ~w147;
assign w153 = (~w147 & w151) | (~w147 & w152) | (w151 & w152);
assign w154 = ~pi2 & ~w153;
assign w155 = ~pi6 & ~pi8;
assign w156 = ~pi0 & pi6;
assign w157 = pi2 & pi8;
assign w158 = (pi8 & w156) | (pi8 & w157) | (w156 & w157);
assign w159 = pi5 & ~w155;
assign w160 = (~w155 & ~w158) | (~w155 & w159) | (~w158 & w159);
assign w161 = ~pi9 & ~w160;
assign w162 = pi1 & w161;
assign w163 = (pi1 & w154) | (pi1 & w162) | (w154 & w162);
assign w164 = ~pi3 & w0;
assign w165 = pi2 & ~pi6;
assign w166 = w115 & w165;
assign w167 = ~pi3 & w166;
assign w168 = w0 & w167;
assign w169 = (w163 & w164) | (w163 & w168) | (w164 & w168);
assign w170 = ~pi7 & w55;
assign w171 = pi0 & pi8;
assign w172 = pi5 & w171;
assign w173 = pi6 & ~w128;
assign w174 = ~w172 & ~w173;
assign w175 = pi9 & ~w174;
assign w176 = ~pi0 & pi8;
assign w177 = ~w50 & ~w176;
assign w178 = ~pi5 & ~w177;
assign w179 = pi2 & w178;
assign w180 = (pi2 & w175) | (pi2 & w179) | (w175 & w179);
assign w181 = ~pi8 & w32;
assign w182 = w146 & w181;
assign w183 = ~pi4 & w182;
assign w184 = (~pi4 & w180) | (~pi4 & w183) | (w180 & w183);
assign w185 = ~pi6 & ~pi9;
assign w186 = pi8 & w185;
assign w187 = pi6 & pi9;
assign w188 = pi4 & w187;
assign w189 = (pi4 & w186) | (pi4 & w188) | (w186 & w188);
assign w190 = pi5 & ~pi8;
assign w191 = w185 & w190;
assign w192 = ~pi2 & w191;
assign w193 = (~pi2 & w189) | (~pi2 & w192) | (w189 & w192);
assign w194 = ~pi0 & w193;
assign w195 = w170 & w194;
assign w196 = (w170 & w184) | (w170 & w195) | (w184 & w195);
assign w197 = ~w169 & ~w196;
assign w198 = ~w144 & w197;
assign w199 = ~pi1 & w105;
assign w200 = ~pi2 & pi8;
assign w201 = pi1 & pi5;
assign w202 = ~w200 & w201;
assign w203 = ~w199 & ~w202;
assign w204 = pi2 & w190;
assign w205 = ~pi1 & ~pi5;
assign w206 = ~pi3 & w205;
assign w207 = (~pi3 & w204) | (~pi3 & w206) | (w204 & w206);
assign w208 = w203 & ~w207;
assign w209 = pi0 & ~w208;
assign w210 = ~pi1 & pi8;
assign w211 = (~pi3 & w142) | (~pi3 & w210) | (w142 & w210);
assign w212 = ~pi0 & w42;
assign w213 = (~pi0 & w211) | (~pi0 & w212) | (w211 & w212);
assign w214 = ~pi2 & w213;
assign w215 = ~pi6 & ~w214;
assign w216 = ~w209 & w215;
assign w217 = ~pi0 & w5;
assign w218 = ~pi1 & pi6;
assign w219 = ~w176 & w218;
assign w220 = ~w217 & ~w219;
assign w221 = ~pi2 & ~w220;
assign w222 = (pi8 & w200) | (pi8 & w218) | (w200 & w218);
assign w223 = pi1 & ~pi2;
assign w224 = pi3 & w223;
assign w225 = (pi3 & w222) | (pi3 & w224) | (w222 & w224);
assign w226 = ~pi5 & w225;
assign w227 = (~pi5 & w221) | (~pi5 & w226) | (w221 & w226);
assign w228 = ~pi9 & ~w227;
assign w229 = ~w216 & w228;
assign w230 = pi5 & w5;
assign w231 = pi2 & pi3;
assign w232 = pi9 & ~w231;
assign w233 = (pi9 & ~w230) | (pi9 & w232) | (~w230 & w232);
assign w234 = pi1 & pi3;
assign w235 = (pi2 & w15) | (pi2 & w234) | (w15 & w234);
assign w236 = pi3 & pi5;
assign w237 = ~w235 & ~w236;
assign w238 = ~pi2 & ~pi8;
assign w239 = ~pi1 & pi3;
assign w240 = w238 & w239;
assign w241 = pi0 & w201;
assign w242 = (pi0 & w240) | (pi0 & w241) | (w240 & w241);
assign w243 = w237 & ~w242;
assign w244 = ~pi6 & w233;
assign w245 = (w233 & w243) | (w233 & w244) | (w243 & w244);
assign w246 = ~pi7 & ~w245;
assign w247 = ~pi4 & w246;
assign w248 = ~w229 & w247;
assign w249 = w198 & ~w248;
assign w250 = pi0 & ~pi4;
assign w251 = ~pi2 & pi3;
assign w252 = ~pi1 & pi9;
assign w253 = ~w251 & ~w252;
assign w254 = (~pi5 & w105) | (~pi5 & w253) | (w105 & w253);
assign w255 = pi3 & pi6;
assign w256 = (pi3 & ~w145) | (pi3 & w255) | (~w145 & w255);
assign w257 = pi2 & ~w256;
assign w258 = w254 & ~w257;
assign w259 = w50 & w223;
assign w260 = ~pi3 & w252;
assign w261 = ~w259 & ~w260;
assign w262 = pi1 & ~pi9;
assign w263 = ~pi3 & ~pi6;
assign w264 = ~w262 & w263;
assign w265 = pi2 & ~pi9;
assign w266 = ~w218 & w265;
assign w267 = ~w264 & ~w266;
assign w268 = pi8 & ~w267;
assign w269 = w261 & ~w268;
assign w270 = w258 & w269;
assign w271 = pi8 & pi9;
assign w272 = pi3 & w271;
assign w273 = (pi3 & w51) | (pi3 & w272) | (w51 & w272);
assign w274 = pi2 & w271;
assign w275 = ~pi1 & w274;
assign w276 = (~pi1 & w273) | (~pi1 & w275) | (w273 & w275);
assign w277 = ~pi2 & ~pi5;
assign w278 = w50 & w277;
assign w279 = ~pi6 & w278;
assign w280 = (~pi6 & w276) | (~pi6 & w279) | (w276 & w279);
assign w281 = w250 & w280;
assign w282 = (w250 & w270) | (w250 & w281) | (w270 & w281);
assign w283 = pi6 & ~pi8;
assign w284 = ~w271 & ~w283;
assign w285 = ~pi5 & ~w284;
assign w286 = ~pi3 & w18;
assign w287 = pi4 & ~w286;
assign w288 = (pi4 & w285) | (pi4 & w287) | (w285 & w287);
assign w289 = ~pi0 & ~w288;
assign w290 = pi2 & ~w149;
assign w291 = pi3 & pi8;
assign w292 = (~pi1 & w1) | (~pi1 & w291) | (w1 & w291);
assign w293 = ~w290 & ~w292;
assign w294 = pi5 & ~w293;
assign w295 = ~w43 & ~w145;
assign w296 = ~pi1 & ~w295;
assign w297 = ~pi2 & pi9;
assign w298 = (~pi2 & w283) | (~pi2 & w297) | (w283 & w297);
assign w299 = pi3 & w298;
assign w300 = (pi3 & w296) | (pi3 & w299) | (w296 & w299);
assign w301 = ~w294 & ~w300;
assign w302 = ~pi2 & pi5;
assign w303 = pi2 & ~pi5;
assign w304 = ~w302 & ~w303;
assign w305 = pi1 & w115;
assign w306 = ~w304 & w305;
assign w307 = ~pi5 & pi6;
assign w308 = w137 & w307;
assign w309 = pi1 & ~w42;
assign w310 = ~w308 & ~w309;
assign w311 = w44 & ~w310;
assign w312 = ~w306 & ~w311;
assign w313 = w301 & w312;
assign w314 = w98 & w155;
assign w315 = ~pi4 & ~w314;
assign w316 = ~pi8 & w187;
assign w317 = ~pi3 & w185;
assign w318 = (~pi3 & w316) | (~pi3 & w317) | (w316 & w317);
assign w319 = pi1 & w318;
assign w320 = w315 & ~w319;
assign w321 = w289 & ~w320;
assign w322 = (w289 & ~w313) | (w289 & w321) | (~w313 & w321);
assign w323 = ~w282 & ~w322;
assign w324 = w124 & ~w146;
assign w325 = ~pi3 & w324;
assign w326 = ~w50 & ~w271;
assign w327 = ~pi5 & ~w34;
assign w328 = (~w34 & w326) | (~w34 & w327) | (w326 & w327);
assign w329 = pi1 & ~w328;
assign w330 = ~pi9 & ~w5;
assign w331 = pi2 & w145;
assign w332 = (pi2 & w330) | (pi2 & w331) | (w330 & w331);
assign w333 = w325 & w332;
assign w334 = (w325 & w329) | (w325 & w333) | (w329 & w333);
assign w335 = pi7 & ~w214;
assign w336 = ~w209 & w335;
assign w337 = ~pi2 & w143;
assign w338 = w336 & w337;
assign w339 = ~w334 & w338;
assign w340 = w323 & w339;
assign w341 = w214 & w337;
assign w342 = (w209 & w337) | (w209 & w341) | (w337 & w341);
assign w343 = pi7 & ~w342;
assign w344 = w334 & ~w343;
assign w345 = (~w323 & ~w343) | (~w323 & w344) | (~w343 & w344);
assign w346 = ~w340 & ~w345;
assign w347 = ~w115 & w231;
assign w348 = ~pi5 & w347;
assign w349 = (~pi2 & w50) | (~pi2 & w277) | (w50 & w277);
assign w350 = ~pi3 & w34;
assign w351 = (~pi3 & w349) | (~pi3 & w350) | (w349 & w350);
assign w352 = ~w15 & ~w91;
assign w353 = pi8 & ~w352;
assign w354 = ~w351 & ~w353;
assign w355 = (pi6 & w20) | (pi6 & ~w347) | (w20 & ~w347);
assign w356 = (~w348 & w354) | (~w348 & w355) | (w354 & w355);
assign w357 = w62 & w142;
assign w358 = pi6 & w142;
assign w359 = w137 & ~w142;
assign w360 = ~w358 & ~w359;
assign w361 = ~pi9 & ~w360;
assign w362 = (~w356 & w357) | (~w356 & w361) | (w357 & w361);
assign w363 = pi0 & pi1;
assign w364 = (w241 & ~w347) | (w241 & w363) | (~w347 & w363);
assign w365 = pi1 & pi6;
assign w366 = pi1 & w20;
assign w367 = (~w347 & w365) | (~w347 & w366) | (w365 & w366);
assign w368 = pi0 & w367;
assign w369 = (w354 & w364) | (w354 & w368) | (w364 & w368);
assign w370 = (pi0 & w362) | (pi0 & w369) | (w362 & w369);
assign w371 = ~w91 & ~w149;
assign w372 = ~pi2 & ~w371;
assign w373 = ~w115 & ~w263;
assign w374 = pi1 & ~w373;
assign w375 = (pi1 & w372) | (pi1 & w374) | (w372 & w374);
assign w376 = w62 & w375;
assign w377 = ~pi1 & w373;
assign w378 = ~w372 & w377;
assign w379 = ~pi5 & w378;
assign w380 = (~pi5 & w376) | (~pi5 & w379) | (w376 & w379);
assign w381 = ~pi6 & w378;
assign w382 = pi5 & pi8;
assign w383 = (~pi9 & w32) | (~pi9 & w382) | (w32 & w382);
assign w384 = ~pi6 & w238;
assign w385 = (~pi6 & w383) | (~pi6 & w384) | (w383 & w384);
assign w386 = pi9 & w165;
assign w387 = ~pi5 & w43;
assign w388 = (~pi5 & w386) | (~pi5 & w387) | (w386 & w387);
assign w389 = ~w385 & ~w388;
assign w390 = pi3 & ~w389;
assign w391 = ~w381 & ~w390;
assign w392 = ~w380 & w391;
assign w393 = ~pi4 & ~w392;
assign w394 = (~pi4 & w370) | (~pi4 & w393) | (w370 & w393);
assign w395 = ~pi5 & ~pi6;
assign w396 = w271 & w395;
assign w397 = ~pi3 & w20;
assign w398 = (~pi3 & w396) | (~pi3 & w397) | (w396 & w397);
assign w399 = ~pi2 & pi4;
assign w400 = w398 & w399;
assign w401 = pi6 & ~w25;
assign w402 = ~pi4 & w231;
assign w403 = (~pi4 & w401) | (~pi4 & w402) | (w401 & w402);
assign w404 = ~pi1 & w403;
assign w405 = (~pi1 & w400) | (~pi1 & w404) | (w400 & w404);
assign w406 = ~pi5 & w403;
assign w407 = (~pi5 & w400) | (~pi5 & w406) | (w400 & w406);
assign w408 = ~pi6 & pi9;
assign w409 = w382 & w408;
assign w410 = ~pi9 & w42;
assign w411 = ~w409 & ~w410;
assign w412 = pi2 & ~w411;
assign w413 = pi6 & w42;
assign w414 = (pi3 & w8) | (pi3 & w149) | (w8 & w149);
assign w415 = ~w413 & ~w414;
assign w416 = pi1 & ~w415;
assign w417 = (pi1 & w412) | (pi1 & w416) | (w412 & w416);
assign w418 = ~w407 & ~w417;
assign w419 = pi4 & ~w405;
assign w420 = (~w405 & w418) | (~w405 & w419) | (w418 & w419);
assign w421 = ~pi0 & ~w420;
assign w422 = ~w394 & ~w421;
assign w423 = ~pi7 & ~w422;
assign w424 = pi2 & ~pi4;
assign w425 = ~w74 & w424;
assign w426 = pi3 & ~pi4;
assign w427 = ~pi3 & pi4;
assign w428 = ~w426 & ~w427;
assign w429 = ~pi2 & ~w428;
assign w430 = w74 & w429;
assign w431 = ~w425 & ~w430;
assign w432 = ~pi7 & ~w431;
assign w433 = w20 & w432;
assign w434 = ~pi2 & w74;
assign w435 = ~pi4 & ~w434;
assign w436 = pi3 & w435;
assign w437 = w427 & w434;
assign w438 = ~w436 & ~w437;
assign w439 = ~pi7 & ~w438;
assign w440 = w20 & w439;
assign w441 = ~w20 & ~w427;
assign w442 = (~w20 & ~w434) | (~w20 & w441) | (~w434 & w441);
assign w443 = ~pi7 & ~w442;
assign w444 = pi2 & w262;
assign w445 = ~pi8 & w80;
assign w446 = pi0 & w78;
assign w447 = (pi0 & w445) | (pi0 & w446) | (w445 & w446);
assign w448 = ~w444 & ~w447;
assign w449 = pi8 & w252;
assign w450 = ~pi0 & w262;
assign w451 = (~pi0 & w449) | (~pi0 & w450) | (w449 & w450);
assign w452 = ~pi6 & w451;
assign w453 = w448 & ~w452;
assign w454 = ~pi5 & ~w453;
assign w455 = w43 & w171;
assign w456 = w5 & ~w117;
assign w457 = ~w455 & ~w456;
assign w458 = pi9 & ~w457;
assign w459 = pi0 & pi5;
assign w460 = ~w176 & ~w459;
assign w461 = pi3 & w262;
assign w462 = ~w460 & w461;
assign w463 = (pi3 & w458) | (pi3 & w462) | (w458 & w462);
assign w464 = (pi3 & w454) | (pi3 & w463) | (w454 & w463);
assign w465 = ~w14 & w302;
assign w466 = (pi9 & w187) | (pi9 & w303) | (w187 & w303);
assign w467 = ~pi0 & w466;
assign w468 = ~w465 & ~w467;
assign w469 = ~pi8 & ~w468;
assign w470 = pi2 & ~w50;
assign w471 = pi0 & w271;
assign w472 = ~w470 & ~w471;
assign w473 = pi1 & ~pi6;
assign w474 = (pi1 & w472) | (pi1 & w473) | (w472 & w473);
assign w475 = ~w469 & w474;
assign w476 = w34 & w176;
assign w477 = pi0 & ~w382;
assign w478 = ~pi9 & w283;
assign w479 = (~pi9 & w477) | (~pi9 & w478) | (w477 & w478);
assign w480 = pi2 & ~w476;
assign w481 = (~w476 & ~w479) | (~w476 & w480) | (~w479 & w480);
assign w482 = ~pi1 & w481;
assign w483 = ~w475 & ~w482;
assign w484 = ~w464 & ~w483;
assign w485 = ~pi7 & ~w484;
assign w486 = (~pi9 & w32) | (~pi9 & w205) | (w32 & w205);
assign w487 = ~pi6 & w486;
assign w488 = pi5 & pi9;
assign w489 = w363 & w488;
assign w490 = (pi0 & w487) | (pi0 & w489) | (w487 & w489);
assign w491 = ~w110 & w117;
assign w492 = pi8 & w491;
assign w493 = (pi8 & w490) | (pi8 & w492) | (w490 & w492);
assign w494 = ~pi1 & w50;
assign w495 = pi2 & w4;
assign w496 = ~w494 & ~w495;
assign w497 = pi5 & ~w496;
assign w498 = ~w51 & ~w274;
assign w499 = pi6 & ~w498;
assign w500 = ~w497 & ~w499;
assign w501 = ~w493 & w500;
assign w502 = ~pi7 & ~w501;
assign w503 = ~pi3 & ~pi4;
assign w504 = ~pi0 & pi1;
assign w505 = w32 & w504;
assign w506 = pi1 & w297;
assign w507 = w171 & w506;
assign w508 = w74 & w265;
assign w509 = pi7 & w508;
assign w510 = (pi7 & w507) | (pi7 & w509) | (w507 & w509);
assign w511 = ~w505 & ~w510;
assign w512 = w395 & w503;
assign w513 = pi7 & w32;
assign w514 = ~pi0 & w1;
assign w515 = ~w513 & ~w514;
assign w516 = ~pi3 & ~pi8;
assign w517 = w395 & w516;
assign w518 = ~pi4 & w517;
assign w519 = ~w515 & w518;
assign w520 = (~w511 & w512) | (~w511 & w519) | (w512 & w519);
assign w521 = (w502 & w503) | (w502 & w520) | (w503 & w520);
assign w522 = (~pi4 & w485) | (~pi4 & w521) | (w485 & w521);
assign w523 = ~w443 & ~w522;
assign w524 = pi0 & pi3;
assign w525 = ~pi2 & ~w524;
assign w526 = ~w326 & ~w525;
assign w527 = pi5 & w231;
assign w528 = (pi5 & w526) | (pi5 & w527) | (w526 & w527);
assign w529 = pi3 & w50;
assign w530 = pi0 & pi2;
assign w531 = w529 & w530;
assign w532 = ~pi1 & ~w531;
assign w533 = ~w528 & w532;
assign w534 = pi3 & ~pi9;
assign w535 = w302 & w534;
assign w536 = ~w236 & ~w265;
assign w537 = ~pi0 & ~w536;
assign w538 = pi5 & w251;
assign w539 = ~pi8 & w538;
assign w540 = (~pi8 & w537) | (~pi8 & w539) | (w537 & w539);
assign w541 = ~w535 & ~w540;
assign w542 = ~w265 & ~w297;
assign w543 = pi0 & ~w542;
assign w544 = pi5 & ~pi9;
assign w545 = ~pi0 & w544;
assign w546 = pi8 & w545;
assign w547 = (pi8 & w543) | (pi8 & w546) | (w543 & w546);
assign w548 = w15 & w145;
assign w549 = ~pi3 & w548;
assign w550 = (~pi3 & w547) | (~pi3 & w549) | (w547 & w549);
assign w551 = w541 & ~w550;
assign w552 = ~pi1 & ~w533;
assign w553 = (~w533 & ~w551) | (~w533 & w552) | (~w551 & w552);
assign w554 = ~pi6 & ~pi7;
assign w555 = pi4 & ~w142;
assign w556 = (pi4 & ~w434) | (pi4 & w555) | (~w434 & w555);
assign w557 = w554 & ~w556;
assign w558 = pi5 & w271;
assign w559 = ~pi4 & ~w231;
assign w560 = (~pi4 & ~w558) | (~pi4 & w559) | (~w558 & w559);
assign w561 = ~w556 & ~w560;
assign w562 = w554 & w561;
assign w563 = (w553 & w557) | (w553 & w562) | (w557 & w562);
assign w564 = ~pi0 & w32;
assign w565 = ~w350 & ~w564;
assign w566 = ~pi8 & ~w565;
assign w567 = pi0 & w115;
assign w568 = ~w470 & ~w567;
assign w569 = pi6 & ~w568;
assign w570 = ~w566 & ~w569;
assign w571 = w156 & ~w326;
assign w572 = ~w12 & ~w145;
assign w573 = ~pi2 & ~pi6;
assign w574 = ~w572 & w573;
assign w575 = ~w571 & ~w574;
assign w576 = pi3 & ~w575;
assign w577 = w570 & ~w576;
assign w578 = ~pi1 & ~w577;
assign w579 = w62 & w200;
assign w580 = ~pi3 & w157;
assign w581 = ~pi2 & w283;
assign w582 = ~w580 & ~w581;
assign w583 = ~pi3 & pi8;
assign w584 = ~w43 & ~w583;
assign w585 = pi0 & ~w584;
assign w586 = w582 & ~w585;
assign w587 = ~pi9 & ~w579;
assign w588 = (~w579 & w586) | (~w579 & w587) | (w586 & w587);
assign w589 = ~pi3 & w50;
assign w590 = ~pi0 & ~pi2;
assign w591 = w271 & w590;
assign w592 = pi2 & ~w271;
assign w593 = ~w591 & ~w592;
assign w594 = ~pi3 & ~w589;
assign w595 = (~w589 & w593) | (~w589 & w594) | (w593 & w594);
assign w596 = ~w44 & ~w157;
assign w597 = pi0 & ~w596;
assign w598 = ~pi6 & w597;
assign w599 = (~pi6 & ~w595) | (~pi6 & w598) | (~w595 & w598);
assign w600 = w588 & ~w599;
assign w601 = pi1 & ~w600;
assign w602 = ~w578 & ~w601;
assign w603 = ~pi2 & pi7;
assign w604 = w567 & w603;
assign w605 = ~w115 & ~w145;
assign w606 = w117 & ~w605;
assign w607 = ~w604 & ~w606;
assign w608 = ~pi1 & w143;
assign w609 = ~w607 & w608;
assign w610 = ~pi5 & ~pi7;
assign w611 = ~pi4 & w610;
assign w612 = ~w609 & ~w611;
assign w613 = w251 & w283;
assign w614 = ~pi9 & w613;
assign w615 = ~pi4 & w614;
assign w616 = w610 & w615;
assign w617 = ~w609 & ~w616;
assign w618 = (w602 & w612) | (w602 & w617) | (w612 & w617);
assign w619 = ~w563 & w618;
assign w620 = pi0 & pi6;
assign w621 = (pi6 & ~w271) | (pi6 & w620) | (~w271 & w620);
assign w622 = (~pi1 & w176) | (~pi1 & w252) | (w176 & w252);
assign w623 = w621 & ~w622;
assign w624 = pi3 & w424;
assign w625 = (w426 & w623) | (w426 & w624) | (w623 & w624);
assign w626 = ~pi1 & ~w2;
assign w627 = pi8 & ~w363;
assign w628 = ~w626 & ~w627;
assign w629 = ~pi6 & ~w628;
assign w630 = w625 & ~w629;
assign w631 = w437 & w610;
assign w632 = (w610 & w630) | (w610 & w631) | (w630 & w631);
assign w633 = w291 & w302;
assign w634 = ~pi3 & w303;
assign w635 = ~w633 & ~w634;
assign w636 = pi1 & ~w635;
assign w637 = ~w205 & ~w459;
assign w638 = pi8 & w251;
assign w639 = ~w637 & w638;
assign w640 = pi9 & w639;
assign w641 = (pi9 & w636) | (pi9 & w640) | (w636 & w640);
assign w642 = pi3 & w252;
assign w643 = w302 & w642;
assign w644 = ~w78 & ~w80;
assign w645 = pi2 & ~w644;
assign w646 = ~pi2 & w262;
assign w647 = ~pi5 & w34;
assign w648 = (~pi5 & w646) | (~pi5 & w647) | (w646 & w647);
assign w649 = ~w645 & ~w648;
assign w650 = pi3 & ~w643;
assign w651 = (~w643 & w649) | (~w643 & w650) | (w649 & w650);
assign w652 = w80 & w302;
assign w653 = ~pi3 & w78;
assign w654 = ~w652 & ~w653;
assign w655 = ~pi0 & ~w654;
assign w656 = ~pi8 & w655;
assign w657 = (~pi8 & ~w651) | (~pi8 & w656) | (~w651 & w656);
assign w658 = ~w641 & ~w657;
assign w659 = ~pi1 & pi5;
assign w660 = w251 & w659;
assign w661 = pi1 & pi2;
assign w662 = w142 & ~w661;
assign w663 = ~pi2 & w659;
assign w664 = ~w662 & ~w663;
assign w665 = ~pi0 & ~w660;
assign w666 = (~w660 & w664) | (~w660 & w665) | (w664 & w665);
assign w667 = pi8 & ~w666;
assign w668 = ~pi0 & w105;
assign w669 = ~pi3 & pi5;
assign w670 = pi1 & w669;
assign w671 = (pi1 & w668) | (pi1 & w670) | (w668 & w670);
assign w672 = pi2 & w671;
assign w673 = ~pi9 & w672;
assign w674 = (~pi9 & w667) | (~pi9 & w673) | (w667 & w673);
assign w675 = ~pi7 & w674;
assign w676 = (~pi7 & ~w658) | (~pi7 & w675) | (~w658 & w675);
assign w677 = pi2 & ~w605;
assign w678 = ~pi1 & w51;
assign w679 = (~pi1 & w677) | (~pi1 & w678) | (w677 & w678);
assign w680 = ~pi2 & w115;
assign w681 = w96 & w680;
assign w682 = pi0 & ~w681;
assign w683 = w145 & w223;
assign w684 = ~pi0 & w683;
assign w685 = ~w681 & ~w684;
assign w686 = (~w679 & w682) | (~w679 & w685) | (w682 & w685);
assign w687 = w142 & ~w686;
assign w688 = w124 & w687;
assign w689 = (w124 & w676) | (w124 & w688) | (w676 & w688);
assign w690 = ~w632 & ~w689;
assign w691 = ~pi1 & ~w50;
assign w692 = pi0 & ~pi6;
assign w693 = ~pi5 & w692;
assign w694 = ~pi7 & ~w231;
assign w695 = (~pi7 & ~w693) | (~pi7 & w694) | (~w693 & w694);
assign w696 = ~w691 & ~w695;
assign w697 = ~pi3 & pi6;
assign w698 = ~pi4 & ~w697;
assign w699 = ~pi2 & ~pi4;
assign w700 = (~pi2 & w55) | (~pi2 & w699) | (w55 & w699);
assign w701 = ~w698 & ~w700;
assign w702 = (~pi7 & ~w25) | (~pi7 & w109) | (~w25 & w109);
assign w703 = pi2 & ~pi3;
assign w704 = ~pi0 & ~pi7;
assign w705 = (~pi0 & w703) | (~pi0 & w704) | (w703 & w704);
assign w706 = ~w702 & ~w705;
assign w707 = ~w20 & ~w706;
assign w708 = ~w701 & w707;
assign w709 = ~w696 & w708;
assign w710 = pi5 & ~w50;
assign w711 = (pi2 & w274) | (pi2 & w710) | (w274 & w710);
assign w712 = pi2 & w239;
assign w713 = (w1 & ~w711) | (w1 & w712) | (~w711 & w712);
assign w714 = (~pi1 & w239) | (~pi1 & ~w711) | (w239 & ~w711);
assign w715 = ~w395 & w427;
assign w716 = (pi8 & w68) | (pi8 & w488) | (w68 & w488);
assign w717 = pi0 & ~w187;
assign w718 = (~w187 & ~w716) | (~w187 & w717) | (~w716 & w717);
assign w719 = ~pi3 & ~w715;
assign w720 = (~w715 & ~w718) | (~w715 & w719) | (~w718 & w719);
assign w721 = w714 & ~w720;
assign w722 = ~w713 & ~w721;
assign w723 = (pi8 & w187) | (pi8 & w583) | (w187 & w583);
assign w724 = ~pi0 & w723;
assign w725 = ~pi3 & ~w110;
assign w726 = ~pi2 & w725;
assign w727 = (~pi2 & w724) | (~pi2 & w726) | (w724 & w726);
assign w728 = pi1 & ~w727;
assign w729 = (~pi6 & w155) | (~pi6 & ~w488) | (w155 & ~w488);
assign w730 = ~pi3 & ~w729;
assign w731 = w8 & ~w271;
assign w732 = w165 & w731;
assign w733 = ~w730 & ~w732;
assign w734 = w728 & w733;
assign w735 = w722 & ~w734;
assign w736 = w709 & ~w735;
assign w737 = pi0 & ~w691;
assign w738 = pi1 & ~w271;
assign w739 = ~w737 & ~w738;
assign w740 = pi2 & ~w739;
assign w741 = w426 & w740;
assign w742 = ~w437 & ~w741;
assign w743 = w610 & ~w742;
assign w744 = ~pi6 & w743;
assign one = 1;
assign po00 = ~w127;
assign po01 = ~w249;
assign po02 = ~w346;
assign po03 = w423;
assign po04 = w433;
assign po05 = w440;
assign po06 = w523;
assign po07 = w619;
assign po08 = w690;
assign po09 = w736;
assign po10 = w744;
endmodule

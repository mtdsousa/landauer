module dec_best_speed (
        pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, 
        po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255);
input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419;
assign w0 = ~pi4 & ~pi5;
assign w1 = ~pi6 & pi7;
assign w2 = w0 & w1;
assign w3 = ~pi0 & ~pi1;
assign w4 = ~pi2 & w3;
assign w5 = w2 & w4;
assign w6 = ~pi3 & w5;
assign w7 = pi0 & ~pi1;
assign w8 = ~pi2 & w7;
assign w9 = w2 & w8;
assign w10 = ~pi3 & w9;
assign w11 = ~pi0 & pi1;
assign w12 = ~pi2 & w11;
assign w13 = w2 & w12;
assign w14 = ~pi3 & w13;
assign w15 = pi0 & pi1;
assign w16 = ~pi2 & w15;
assign w17 = w2 & w16;
assign w18 = ~pi3 & w17;
assign w19 = pi2 & w3;
assign w20 = w2 & w19;
assign w21 = ~pi3 & w20;
assign w22 = pi2 & w7;
assign w23 = w2 & w22;
assign w24 = ~pi3 & w23;
assign w25 = pi2 & w11;
assign w26 = w2 & w25;
assign w27 = ~pi3 & w26;
assign w28 = pi2 & w15;
assign w29 = w2 & w28;
assign w30 = ~pi3 & w29;
assign w31 = pi3 & w5;
assign w32 = pi3 & w9;
assign w33 = pi3 & w13;
assign w34 = pi3 & w17;
assign w35 = pi3 & w20;
assign w36 = pi3 & w23;
assign w37 = pi3 & w26;
assign w38 = pi3 & w29;
assign w39 = pi4 & ~pi5;
assign w40 = w1 & w39;
assign w41 = w4 & w40;
assign w42 = ~pi3 & w41;
assign w43 = w8 & w40;
assign w44 = ~pi3 & w43;
assign w45 = w12 & w40;
assign w46 = ~pi3 & w45;
assign w47 = w16 & w40;
assign w48 = ~pi3 & w47;
assign w49 = w19 & w40;
assign w50 = ~pi3 & w49;
assign w51 = w22 & w40;
assign w52 = ~pi3 & w51;
assign w53 = w25 & w40;
assign w54 = ~pi3 & w53;
assign w55 = w28 & w40;
assign w56 = ~pi3 & w55;
assign w57 = pi3 & w41;
assign w58 = pi3 & w43;
assign w59 = pi3 & w45;
assign w60 = pi3 & w47;
assign w61 = pi3 & w49;
assign w62 = pi3 & w51;
assign w63 = pi3 & w53;
assign w64 = pi3 & w55;
assign w65 = ~pi4 & pi5;
assign w66 = w1 & w65;
assign w67 = w4 & w66;
assign w68 = ~pi3 & w67;
assign w69 = w8 & w66;
assign w70 = ~pi3 & w69;
assign w71 = w12 & w66;
assign w72 = ~pi3 & w71;
assign w73 = w16 & w66;
assign w74 = ~pi3 & w73;
assign w75 = w19 & w66;
assign w76 = ~pi3 & w75;
assign w77 = w22 & w66;
assign w78 = ~pi3 & w77;
assign w79 = w25 & w66;
assign w80 = ~pi3 & w79;
assign w81 = w28 & w66;
assign w82 = ~pi3 & w81;
assign w83 = pi3 & w67;
assign w84 = pi3 & w69;
assign w85 = pi3 & w71;
assign w86 = pi3 & w73;
assign w87 = pi3 & w75;
assign w88 = pi3 & w77;
assign w89 = pi3 & w79;
assign w90 = pi3 & w81;
assign w91 = pi4 & pi5;
assign w92 = w1 & w91;
assign w93 = w4 & w92;
assign w94 = ~pi3 & w93;
assign w95 = w8 & w92;
assign w96 = ~pi3 & w95;
assign w97 = w12 & w92;
assign w98 = ~pi3 & w97;
assign w99 = w16 & w92;
assign w100 = ~pi3 & w99;
assign w101 = w19 & w92;
assign w102 = ~pi3 & w101;
assign w103 = w22 & w92;
assign w104 = ~pi3 & w103;
assign w105 = w25 & w92;
assign w106 = ~pi3 & w105;
assign w107 = w28 & w92;
assign w108 = ~pi3 & w107;
assign w109 = pi3 & w93;
assign w110 = pi3 & w95;
assign w111 = pi3 & w97;
assign w112 = pi3 & w99;
assign w113 = pi3 & w101;
assign w114 = pi3 & w103;
assign w115 = pi3 & w105;
assign w116 = pi3 & w107;
assign w117 = pi6 & pi7;
assign w118 = w0 & w117;
assign w119 = w4 & w118;
assign w120 = ~pi3 & w119;
assign w121 = w8 & w118;
assign w122 = ~pi3 & w121;
assign w123 = w12 & w118;
assign w124 = ~pi3 & w123;
assign w125 = w16 & w118;
assign w126 = ~pi3 & w125;
assign w127 = w19 & w118;
assign w128 = ~pi3 & w127;
assign w129 = w22 & w118;
assign w130 = ~pi3 & w129;
assign w131 = w25 & w118;
assign w132 = ~pi3 & w131;
assign w133 = w28 & w118;
assign w134 = ~pi3 & w133;
assign w135 = pi3 & w119;
assign w136 = pi3 & w121;
assign w137 = pi3 & w123;
assign w138 = pi3 & w125;
assign w139 = pi3 & w127;
assign w140 = pi3 & w129;
assign w141 = pi3 & w131;
assign w142 = pi3 & w133;
assign w143 = w39 & w117;
assign w144 = w4 & w143;
assign w145 = ~pi3 & w144;
assign w146 = w8 & w143;
assign w147 = ~pi3 & w146;
assign w148 = w12 & w143;
assign w149 = ~pi3 & w148;
assign w150 = w16 & w143;
assign w151 = ~pi3 & w150;
assign w152 = w19 & w143;
assign w153 = ~pi3 & w152;
assign w154 = w22 & w143;
assign w155 = ~pi3 & w154;
assign w156 = w25 & w143;
assign w157 = ~pi3 & w156;
assign w158 = w28 & w143;
assign w159 = ~pi3 & w158;
assign w160 = pi3 & w144;
assign w161 = pi3 & w146;
assign w162 = pi3 & w148;
assign w163 = pi3 & w150;
assign w164 = pi3 & w152;
assign w165 = pi3 & w154;
assign w166 = pi3 & w156;
assign w167 = pi3 & w158;
assign w168 = w65 & w117;
assign w169 = w4 & w168;
assign w170 = ~pi3 & w169;
assign w171 = w8 & w168;
assign w172 = ~pi3 & w171;
assign w173 = w12 & w168;
assign w174 = ~pi3 & w173;
assign w175 = w16 & w168;
assign w176 = ~pi3 & w175;
assign w177 = w19 & w168;
assign w178 = ~pi3 & w177;
assign w179 = w22 & w168;
assign w180 = ~pi3 & w179;
assign w181 = w25 & w168;
assign w182 = ~pi3 & w181;
assign w183 = w28 & w168;
assign w184 = ~pi3 & w183;
assign w185 = pi3 & w169;
assign w186 = pi3 & w171;
assign w187 = pi3 & w173;
assign w188 = pi3 & w175;
assign w189 = pi3 & w177;
assign w190 = pi3 & w179;
assign w191 = pi3 & w181;
assign w192 = pi3 & w183;
assign w193 = w91 & w117;
assign w194 = w4 & w193;
assign w195 = ~pi3 & w194;
assign w196 = w8 & w193;
assign w197 = ~pi3 & w196;
assign w198 = w12 & w193;
assign w199 = ~pi3 & w198;
assign w200 = w16 & w193;
assign w201 = ~pi3 & w200;
assign w202 = w19 & w193;
assign w203 = ~pi3 & w202;
assign w204 = w22 & w193;
assign w205 = ~pi3 & w204;
assign w206 = w25 & w193;
assign w207 = ~pi3 & w206;
assign w208 = w28 & w193;
assign w209 = ~pi3 & w208;
assign w210 = pi3 & w194;
assign w211 = pi3 & w196;
assign w212 = pi3 & w198;
assign w213 = pi3 & w200;
assign w214 = pi3 & w202;
assign w215 = pi3 & w204;
assign w216 = pi3 & w206;
assign w217 = pi3 & w208;
assign w218 = ~pi6 & ~pi7;
assign w219 = w0 & w218;
assign w220 = w4 & w219;
assign w221 = ~pi3 & w220;
assign w222 = w8 & w219;
assign w223 = ~pi3 & w222;
assign w224 = w12 & w219;
assign w225 = ~pi3 & w224;
assign w226 = w16 & w219;
assign w227 = ~pi3 & w226;
assign w228 = w19 & w219;
assign w229 = ~pi3 & w228;
assign w230 = w22 & w219;
assign w231 = ~pi3 & w230;
assign w232 = w25 & w219;
assign w233 = ~pi3 & w232;
assign w234 = w28 & w219;
assign w235 = ~pi3 & w234;
assign w236 = pi3 & w220;
assign w237 = pi3 & w222;
assign w238 = pi3 & w224;
assign w239 = pi3 & w226;
assign w240 = pi3 & w228;
assign w241 = pi3 & w230;
assign w242 = pi3 & w232;
assign w243 = pi3 & w234;
assign w244 = w39 & w218;
assign w245 = w4 & w244;
assign w246 = ~pi3 & w245;
assign w247 = w8 & w244;
assign w248 = ~pi3 & w247;
assign w249 = w12 & w244;
assign w250 = ~pi3 & w249;
assign w251 = w16 & w244;
assign w252 = ~pi3 & w251;
assign w253 = w19 & w244;
assign w254 = ~pi3 & w253;
assign w255 = w22 & w244;
assign w256 = ~pi3 & w255;
assign w257 = w25 & w244;
assign w258 = ~pi3 & w257;
assign w259 = w28 & w244;
assign w260 = ~pi3 & w259;
assign w261 = pi3 & w245;
assign w262 = pi3 & w247;
assign w263 = pi3 & w249;
assign w264 = pi3 & w251;
assign w265 = pi3 & w253;
assign w266 = pi3 & w255;
assign w267 = pi3 & w257;
assign w268 = pi3 & w259;
assign w269 = w65 & w218;
assign w270 = w4 & w269;
assign w271 = ~pi3 & w270;
assign w272 = w8 & w269;
assign w273 = ~pi3 & w272;
assign w274 = w12 & w269;
assign w275 = ~pi3 & w274;
assign w276 = w16 & w269;
assign w277 = ~pi3 & w276;
assign w278 = w19 & w269;
assign w279 = ~pi3 & w278;
assign w280 = w22 & w269;
assign w281 = ~pi3 & w280;
assign w282 = w25 & w269;
assign w283 = ~pi3 & w282;
assign w284 = w28 & w269;
assign w285 = ~pi3 & w284;
assign w286 = pi3 & w270;
assign w287 = pi3 & w272;
assign w288 = pi3 & w274;
assign w289 = pi3 & w276;
assign w290 = pi3 & w278;
assign w291 = pi3 & w280;
assign w292 = pi3 & w282;
assign w293 = pi3 & w284;
assign w294 = w91 & w218;
assign w295 = w4 & w294;
assign w296 = ~pi3 & w295;
assign w297 = w8 & w294;
assign w298 = ~pi3 & w297;
assign w299 = w12 & w294;
assign w300 = ~pi3 & w299;
assign w301 = w16 & w294;
assign w302 = ~pi3 & w301;
assign w303 = w19 & w294;
assign w304 = ~pi3 & w303;
assign w305 = w22 & w294;
assign w306 = ~pi3 & w305;
assign w307 = w25 & w294;
assign w308 = ~pi3 & w307;
assign w309 = w28 & w294;
assign w310 = ~pi3 & w309;
assign w311 = pi3 & w295;
assign w312 = pi3 & w297;
assign w313 = pi3 & w299;
assign w314 = pi3 & w301;
assign w315 = pi3 & w303;
assign w316 = pi3 & w305;
assign w317 = pi3 & w307;
assign w318 = pi3 & w309;
assign w319 = pi6 & ~pi7;
assign w320 = w0 & w319;
assign w321 = w4 & w320;
assign w322 = ~pi3 & w321;
assign w323 = w8 & w320;
assign w324 = ~pi3 & w323;
assign w325 = w12 & w320;
assign w326 = ~pi3 & w325;
assign w327 = w16 & w320;
assign w328 = ~pi3 & w327;
assign w329 = w19 & w320;
assign w330 = ~pi3 & w329;
assign w331 = w22 & w320;
assign w332 = ~pi3 & w331;
assign w333 = w25 & w320;
assign w334 = ~pi3 & w333;
assign w335 = w28 & w320;
assign w336 = ~pi3 & w335;
assign w337 = pi3 & w321;
assign w338 = pi3 & w323;
assign w339 = pi3 & w325;
assign w340 = pi3 & w327;
assign w341 = pi3 & w329;
assign w342 = pi3 & w331;
assign w343 = pi3 & w333;
assign w344 = pi3 & w335;
assign w345 = w39 & w319;
assign w346 = w4 & w345;
assign w347 = ~pi3 & w346;
assign w348 = w8 & w345;
assign w349 = ~pi3 & w348;
assign w350 = w12 & w345;
assign w351 = ~pi3 & w350;
assign w352 = w16 & w345;
assign w353 = ~pi3 & w352;
assign w354 = w19 & w345;
assign w355 = ~pi3 & w354;
assign w356 = w22 & w345;
assign w357 = ~pi3 & w356;
assign w358 = w25 & w345;
assign w359 = ~pi3 & w358;
assign w360 = w28 & w345;
assign w361 = ~pi3 & w360;
assign w362 = pi3 & w346;
assign w363 = pi3 & w348;
assign w364 = pi3 & w350;
assign w365 = pi3 & w352;
assign w366 = pi3 & w354;
assign w367 = pi3 & w356;
assign w368 = pi3 & w358;
assign w369 = pi3 & w360;
assign w370 = w65 & w319;
assign w371 = w4 & w370;
assign w372 = ~pi3 & w371;
assign w373 = w8 & w370;
assign w374 = ~pi3 & w373;
assign w375 = w12 & w370;
assign w376 = ~pi3 & w375;
assign w377 = w16 & w370;
assign w378 = ~pi3 & w377;
assign w379 = w19 & w370;
assign w380 = ~pi3 & w379;
assign w381 = w22 & w370;
assign w382 = ~pi3 & w381;
assign w383 = w25 & w370;
assign w384 = ~pi3 & w383;
assign w385 = w28 & w370;
assign w386 = ~pi3 & w385;
assign w387 = pi3 & w371;
assign w388 = pi3 & w373;
assign w389 = pi3 & w375;
assign w390 = pi3 & w377;
assign w391 = pi3 & w379;
assign w392 = pi3 & w381;
assign w393 = pi3 & w383;
assign w394 = pi3 & w385;
assign w395 = w91 & w319;
assign w396 = w4 & w395;
assign w397 = ~pi3 & w396;
assign w398 = w8 & w395;
assign w399 = ~pi3 & w398;
assign w400 = w12 & w395;
assign w401 = ~pi3 & w400;
assign w402 = w16 & w395;
assign w403 = ~pi3 & w402;
assign w404 = w19 & w395;
assign w405 = ~pi3 & w404;
assign w406 = w22 & w395;
assign w407 = ~pi3 & w406;
assign w408 = w25 & w395;
assign w409 = ~pi3 & w408;
assign w410 = w28 & w395;
assign w411 = ~pi3 & w410;
assign w412 = pi3 & w396;
assign w413 = pi3 & w398;
assign w414 = pi3 & w400;
assign w415 = pi3 & w402;
assign w416 = pi3 & w404;
assign w417 = pi3 & w406;
assign w418 = pi3 & w408;
assign w419 = pi3 & w410;
assign one = 1;
assign po000 = w6;
assign po001 = w10;
assign po002 = w14;
assign po003 = w18;
assign po004 = w21;
assign po005 = w24;
assign po006 = w27;
assign po007 = w30;
assign po008 = w31;
assign po009 = w32;
assign po010 = w33;
assign po011 = w34;
assign po012 = w35;
assign po013 = w36;
assign po014 = w37;
assign po015 = w38;
assign po016 = w42;
assign po017 = w44;
assign po018 = w46;
assign po019 = w48;
assign po020 = w50;
assign po021 = w52;
assign po022 = w54;
assign po023 = w56;
assign po024 = w57;
assign po025 = w58;
assign po026 = w59;
assign po027 = w60;
assign po028 = w61;
assign po029 = w62;
assign po030 = w63;
assign po031 = w64;
assign po032 = w68;
assign po033 = w70;
assign po034 = w72;
assign po035 = w74;
assign po036 = w76;
assign po037 = w78;
assign po038 = w80;
assign po039 = w82;
assign po040 = w83;
assign po041 = w84;
assign po042 = w85;
assign po043 = w86;
assign po044 = w87;
assign po045 = w88;
assign po046 = w89;
assign po047 = w90;
assign po048 = w94;
assign po049 = w96;
assign po050 = w98;
assign po051 = w100;
assign po052 = w102;
assign po053 = w104;
assign po054 = w106;
assign po055 = w108;
assign po056 = w109;
assign po057 = w110;
assign po058 = w111;
assign po059 = w112;
assign po060 = w113;
assign po061 = w114;
assign po062 = w115;
assign po063 = w116;
assign po064 = w120;
assign po065 = w122;
assign po066 = w124;
assign po067 = w126;
assign po068 = w128;
assign po069 = w130;
assign po070 = w132;
assign po071 = w134;
assign po072 = w135;
assign po073 = w136;
assign po074 = w137;
assign po075 = w138;
assign po076 = w139;
assign po077 = w140;
assign po078 = w141;
assign po079 = w142;
assign po080 = w145;
assign po081 = w147;
assign po082 = w149;
assign po083 = w151;
assign po084 = w153;
assign po085 = w155;
assign po086 = w157;
assign po087 = w159;
assign po088 = w160;
assign po089 = w161;
assign po090 = w162;
assign po091 = w163;
assign po092 = w164;
assign po093 = w165;
assign po094 = w166;
assign po095 = w167;
assign po096 = w170;
assign po097 = w172;
assign po098 = w174;
assign po099 = w176;
assign po100 = w178;
assign po101 = w180;
assign po102 = w182;
assign po103 = w184;
assign po104 = w185;
assign po105 = w186;
assign po106 = w187;
assign po107 = w188;
assign po108 = w189;
assign po109 = w190;
assign po110 = w191;
assign po111 = w192;
assign po112 = w195;
assign po113 = w197;
assign po114 = w199;
assign po115 = w201;
assign po116 = w203;
assign po117 = w205;
assign po118 = w207;
assign po119 = w209;
assign po120 = w210;
assign po121 = w211;
assign po122 = w212;
assign po123 = w213;
assign po124 = w214;
assign po125 = w215;
assign po126 = w216;
assign po127 = w217;
assign po128 = w221;
assign po129 = w223;
assign po130 = w225;
assign po131 = w227;
assign po132 = w229;
assign po133 = w231;
assign po134 = w233;
assign po135 = w235;
assign po136 = w236;
assign po137 = w237;
assign po138 = w238;
assign po139 = w239;
assign po140 = w240;
assign po141 = w241;
assign po142 = w242;
assign po143 = w243;
assign po144 = w246;
assign po145 = w248;
assign po146 = w250;
assign po147 = w252;
assign po148 = w254;
assign po149 = w256;
assign po150 = w258;
assign po151 = w260;
assign po152 = w261;
assign po153 = w262;
assign po154 = w263;
assign po155 = w264;
assign po156 = w265;
assign po157 = w266;
assign po158 = w267;
assign po159 = w268;
assign po160 = w271;
assign po161 = w273;
assign po162 = w275;
assign po163 = w277;
assign po164 = w279;
assign po165 = w281;
assign po166 = w283;
assign po167 = w285;
assign po168 = w286;
assign po169 = w287;
assign po170 = w288;
assign po171 = w289;
assign po172 = w290;
assign po173 = w291;
assign po174 = w292;
assign po175 = w293;
assign po176 = w296;
assign po177 = w298;
assign po178 = w300;
assign po179 = w302;
assign po180 = w304;
assign po181 = w306;
assign po182 = w308;
assign po183 = w310;
assign po184 = w311;
assign po185 = w312;
assign po186 = w313;
assign po187 = w314;
assign po188 = w315;
assign po189 = w316;
assign po190 = w317;
assign po191 = w318;
assign po192 = w322;
assign po193 = w324;
assign po194 = w326;
assign po195 = w328;
assign po196 = w330;
assign po197 = w332;
assign po198 = w334;
assign po199 = w336;
assign po200 = w337;
assign po201 = w338;
assign po202 = w339;
assign po203 = w340;
assign po204 = w341;
assign po205 = w342;
assign po206 = w343;
assign po207 = w344;
assign po208 = w347;
assign po209 = w349;
assign po210 = w351;
assign po211 = w353;
assign po212 = w355;
assign po213 = w357;
assign po214 = w359;
assign po215 = w361;
assign po216 = w362;
assign po217 = w363;
assign po218 = w364;
assign po219 = w365;
assign po220 = w366;
assign po221 = w367;
assign po222 = w368;
assign po223 = w369;
assign po224 = w372;
assign po225 = w374;
assign po226 = w376;
assign po227 = w378;
assign po228 = w380;
assign po229 = w382;
assign po230 = w384;
assign po231 = w386;
assign po232 = w387;
assign po233 = w388;
assign po234 = w389;
assign po235 = w390;
assign po236 = w391;
assign po237 = w392;
assign po238 = w393;
assign po239 = w394;
assign po240 = w397;
assign po241 = w399;
assign po242 = w401;
assign po243 = w403;
assign po244 = w405;
assign po245 = w407;
assign po246 = w409;
assign po247 = w411;
assign po248 = w412;
assign po249 = w413;
assign po250 = w414;
assign po251 = w415;
assign po252 = w416;
assign po253 = w417;
assign po254 = w418;
assign po255 = w419;
endmodule
